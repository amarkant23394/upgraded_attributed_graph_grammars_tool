module test_final(IN_1_0_l,IN_2_0_l,IN_3_0_l,IN_4_0_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_8_r,blif_reset_net_8_r,N1371_0_r,N1508_0_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r);
input IN_1_0_l,IN_2_0_l,IN_3_0_l,IN_4_0_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_8_r,blif_reset_net_8_r;
output N1371_0_r,N1508_0_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r;
wire N1371_0_l,N1508_0_l,n3_0_l,n4_0_l,N6147_3_l,n3_3_l,N6138_3_l,n_42_8_l,G199_8_l,N3_8_l,n3_8_l,N1372_10_l,N1508_10_l,n5_10_l,n6_10_l,n3_0_r,n4_0_r,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n6_4_r,n7_4_r,n8_4_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,N3_8_r,n1_8_r,n3_8_r,N6150_9_r,n3_9_r;
nor I_0(N1371_0_l,IN_2_0_l,n4_0_l);
nor I_1(N1508_0_l,n3_0_l,n4_0_l);
nor I_2(n3_0_l,IN_3_0_l,IN_4_0_l);
not I_3(n4_0_l,IN_1_0_l);
nor I_4(N6147_3_l,IN_3_3_l,n3_3_l);
not I_5(n3_3_l,N6138_3_l);
nor I_6(N6138_3_l,IN_1_3_l,IN_2_3_l);
nor I_7(n_42_8_l,IN_1_8_l,IN_3_8_l);
DFFARX1 I_8(N3_8_l,blif_clk_net_8_r,n1_8_r,G199_8_l,);
and I_9(N3_8_l,IN_6_8_l,n3_8_l);
nand I_10(n3_8_l,IN_2_8_l,IN_3_8_l);
not I_11(N1372_10_l,n6_10_l);
nor I_12(N1508_10_l,n5_10_l,n6_10_l);
nor I_13(n5_10_l,IN_3_10_l,IN_4_10_l);
nand I_14(n6_10_l,IN_1_10_l,IN_2_10_l);
nor I_15(N1371_0_r,n4_0_r,n_42_8_l);
nor I_16(N1508_0_r,n3_0_r,n4_0_r);
nor I_17(n3_0_r,N1371_0_l,N1508_0_l);
not I_18(n4_0_r,N1372_10_l);
nor I_19(N6147_2_r,n5_2_r,n6_2_r);
nor I_20(n5_2_r,n7_2_r,N1508_10_l);
not I_21(n6_2_r,N6138_2_r);
nor I_22(N6138_2_r,n_42_8_l,N6147_3_l);
nor I_23(n7_2_r,N1372_10_l,G199_8_l);
nor I_24(N6147_3_r,n3_3_r,N6147_3_l);
not I_25(n3_3_r,N6138_3_r);
nor I_26(N6138_3_r,G199_8_l,N1508_0_l);
not I_27(N1372_4_r,n7_4_r);
nor I_28(N1508_4_r,n6_4_r,n7_4_r);
nor I_29(n6_4_r,n8_4_r,N6147_3_l);
nand I_30(n7_4_r,N1508_10_l,G199_8_l);
and I_31(n8_4_r,G199_8_l,N1372_10_l);
nor I_32(N1507_6_r,n8_6_r,n9_6_r);
and I_33(N1508_6_r,n6_6_r,n_42_8_l);
nor I_34(n6_6_r,n7_6_r,n8_6_r);
not I_35(n7_6_r,N1508_10_l);
nor I_36(n8_6_r,n9_6_r,N6147_3_l);
and I_37(n9_6_r,N1508_10_l,n_42_8_l);
nor I_38(n_42_8_r,N1371_0_l,n_42_8_l);
DFFARX1 I_39(N3_8_r,blif_clk_net_8_r,n1_8_r,G199_8_r,);
and I_40(N3_8_r,n3_8_r,N1508_0_l);
not I_41(n1_8_r,blif_reset_net_8_r);
nand I_42(n3_8_r,N1371_0_l,N6147_3_l);
not I_43(N6150_9_r,N1371_0_l);
nor I_44(N6147_9_r,N6150_9_r,n3_9_r);
nor I_45(N6134_9_r,n3_9_r,N1372_10_l);
nor I_46(n3_9_r,N1508_0_l,N1371_0_l);
buf I_47(I_BUFF_1_9_r,N1508_0_l);
endmodule


