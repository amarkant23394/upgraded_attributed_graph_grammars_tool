module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,IN_1_3_l_7,IN_2_3_l_7,IN_3_3_l_7,IN_1_4_l_7,IN_2_4_l_7,IN_3_4_l_7,IN_4_4_l_7,IN_5_4_l_7,blif_clk_net_5_r_4,blif_reset_net_5_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,IN_1_3_l_7,IN_2_3_l_7,IN_3_3_l_7,IN_1_4_l_7,IN_2_4_l_7,IN_3_4_l_7,IN_4_4_l_7,IN_5_4_l_7,blif_clk_net_5_r_4,blif_reset_net_5_r_4;
output N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4;
wire N1371_0_r_7,N1508_0_r_7,N6147_2_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,N1507_6_r_7,N1508_6_r_7,n_431_5_r_7,n19_7,n20_7,n21_7,n22_7,n23_7,n24_7,n25_7,n26_7,n27_7,n28_7,n29_7,n30_7,n31_7,n32_7,N1371_0_r_4,n_102_5_r_4,n_431_5_r_4,n4_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4;
nor I_0(N1371_0_r_7,n22_7,n24_7);
nor I_1(N1508_0_r_7,n24_7,n28_7);
nor I_2(N6147_2_r_7,n21_7,n26_7);
nand I_3(n_429_or_0_5_r_7,n19_7,n24_7);
DFFARX1 I_4(n_431_5_r_7,blif_clk_net_5_r_4,n4_4,G78_5_r_7,);
nand I_5(n_576_5_r_7,N1371_0_r_7,n19_7);
not I_6(n_102_5_r_7,n22_7);
nand I_7(n_547_5_r_7,n20_7,n21_7);
nor I_8(N1507_6_r_7,n22_7,n27_7);
nor I_9(N1508_6_r_7,IN_3_1_l_7,n27_7);
nand I_10(n_431_5_r_7,n24_7,n25_7);
nor I_11(n19_7,IN_1_3_l_7,n30_7);
nor I_12(n20_7,n22_7,n23_7);
not I_13(n21_7,n29_7);
nor I_14(n22_7,n29_7,n31_7);
not I_15(n23_7,n27_7);
not I_16(n24_7,N1508_6_r_7);
nand I_17(n25_7,N1507_6_r_7,n19_7);
or I_18(n26_7,n19_7,n23_7);
nand I_19(n27_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_20(n28_7,n19_7,n21_7);
nand I_21(n29_7,IN_1_4_l_7,IN_2_4_l_7);
or I_22(n30_7,IN_2_3_l_7,IN_3_3_l_7);
nor I_23(n31_7,IN_5_4_l_7,n32_7);
and I_24(n32_7,IN_3_4_l_7,IN_4_4_l_7);
nor I_25(N1371_0_r_4,n25_4,n29_4);
nor I_26(N1508_0_r_4,n25_4,n32_4);
nor I_27(N6147_2_r_4,n24_4,n31_4);
or I_28(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_29(n_431_5_r_4,blif_clk_net_5_r_4,n4_4,G78_5_r_4,);
nand I_30(n_576_5_r_4,n22_4,n23_4);
nand I_31(n_102_5_r_4,n34_4,n35_4);
nand I_32(n_547_5_r_4,n26_4,n27_4);
nor I_33(N1507_6_r_4,n27_4,n30_4);
nor I_34(N1508_6_r_4,n30_4,n33_4);
nand I_35(n_431_5_r_4,n_102_5_r_4,n28_4);
not I_36(n4_4,blif_reset_net_5_r_4);
nor I_37(n22_4,n24_4,n25_4);
nor I_38(n23_4,n37_4,N6147_2_r_7);
not I_39(n24_4,n_102_5_r_4);
nand I_40(n25_4,n_576_5_r_7,n_102_5_r_7);
nor I_41(n26_4,n23_4,n24_4);
not I_42(n27_4,n25_4);
nand I_43(n28_4,n23_4,n29_4);
nor I_44(n29_4,n25_4,G78_5_r_7);
not I_45(n30_4,n29_4);
nor I_46(n31_4,N1371_0_r_4,n32_4);
nor I_47(n32_4,n23_4,n29_4);
nand I_48(n33_4,n23_4,n24_4);
nor I_49(n34_4,N1508_0_r_7,G78_5_r_7);
or I_50(n35_4,n36_4,n_429_or_0_5_r_7);
nor I_51(n36_4,N1508_0_r_7,n_547_5_r_7);
or I_52(n37_4,N6147_2_r_7,n_429_or_0_5_r_7);
endmodule


