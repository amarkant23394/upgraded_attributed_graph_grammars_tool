module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_7_r_3,n10_3,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
not I_41(N1372_1_r_3,n40_3);
nor I_42(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_43(N1507_6_r_3,n31_3,n42_3);
nor I_44(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_45(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_46(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_47(n_573_7_r_3,n30_3,n31_3);
nor I_48(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_49(n_569_7_r_3,n30_3,n32_3);
nor I_50(n_452_7_r_3,n35_3,N1508_6_r_1);
not I_51(N6147_9_r_3,n32_3);
nor I_52(N6134_9_r_3,n36_3,n37_3);
not I_53(I_BUFF_1_9_r_3,n45_3);
nor I_54(n4_7_r_3,I_BUFF_1_9_r_3,N1508_6_r_1);
not I_55(n10_3,blif_reset_net_7_r_3);
not I_56(n30_3,n39_3);
not I_57(n31_3,n35_3);
nand I_58(n32_3,n41_3,n_573_7_r_1);
nor I_59(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_60(n34_3,n46_3,G42_7_r_1);
nor I_61(n35_3,n43_3,n44_3);
not I_62(n36_3,n34_3);
nor I_63(n37_3,N6147_9_r_3,N1508_6_r_1);
or I_64(n38_3,n_572_7_r_3,n34_3);
nor I_65(n39_3,n44_3,N1508_0_r_1);
nand I_66(n40_3,n39_3,N1508_6_r_1);
nand I_67(n41_3,N1507_6_r_1,G42_7_r_1);
nor I_68(n42_3,n34_3,n45_3);
not I_69(n43_3,N1507_6_r_1);
nor I_70(n44_3,n_549_7_r_1,n_572_7_r_1);
nand I_71(n45_3,n49_3,n50_3);
and I_72(n46_3,n47_3,n_572_7_r_1);
nand I_73(n47_3,n41_3,n48_3);
not I_74(n48_3,n_573_7_r_1);
nor I_75(n49_3,N6147_9_r_1,N1508_6_r_1);
or I_76(n50_3,n51_3,n_569_7_r_1);
nor I_77(n51_3,N1508_0_r_1,N6134_9_r_1);
endmodule


