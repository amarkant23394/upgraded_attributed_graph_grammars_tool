module test_I3214(I2945,I3058,I3137,I1294_clk,I1301_rst,I3214);
input I2945,I3058,I3137,I1294_clk,I1301_rst;
output I3214;
wire I2568,I2600_rst,I3154,I3246_rst,I3560,I2583,I3263;
DFFARX1 I_0 (I2945,I1294_clk,I2600_rst,I2568);
not I_1(I2600_rst,I1301_rst);
or I_2(I3154,I3137,I3058);
not I_3(I3246_rst,I1301_rst);
nand I_4(I3560,I3263,I2583);
DFFARX1 I_5 (I3154,I1294_clk,I2600_rst,I2583);
DFFARX1 I_6 (I3560,I1294_clk,I3246_rst,I3214);
not I_7(I3263,I2568);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule