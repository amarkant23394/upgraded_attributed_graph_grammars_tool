module test_I5833(I4515,I1477,I1470,I4530,I5833);
input I4515,I1477,I1470,I4530;
output I5833;
wire I5751,I5768,I4524,I4595,I5785,I4742,I5802;
not I_0(I5751,I1477);
nand I_1(I5768,I4530,I4515);
nor I_2(I4524,I4742,I4595);
DFFARX1 I_3(I1470,,,I4595,);
and I_4(I5785,I5768,I4524);
DFFARX1 I_5(I1470,,,I4742,);
DFFARX1 I_6(I5785,I1470,I5751,,,I5802,);
DFFARX1 I_7(I5802,I1470,I5751,,,I5833,);
endmodule


