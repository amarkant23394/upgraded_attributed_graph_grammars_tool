module test_I5719(I4629,I1477,I4518,I1470,I5719);
input I4629,I1477,I4518,I1470;
output I5719;
wire I6265,I6248,I5864,I5751,I6203,I4595,I4527,I4536,I4515,I5915;
and I_0(I6265,I5915,I6248);
nand I_1(I6248,I6203,I5864);
nor I_2(I5864,I4536,I4515);
not I_3(I5751,I1477);
DFFARX1 I_4(I4518,I1470,I5751,,,I6203,);
DFFARX1 I_5(I1470,,,I4595,);
or I_6(I4527,I4629,I4595);
nor I_7(I4536,I4595);
not I_8(I4515,I4629);
DFFARX1 I_9(I4527,I1470,I5751,,,I5915,);
DFFARX1 I_10(I6265,I1470,I5751,,,I5719,);
endmodule


