module test_I16804(I1477,I14957,I12602,I15109,I15016,I1470,I15519,I16804);
input I1477,I14957,I12602,I15109,I15016,I1470,I15519;
output I16804;
wire I14948,I14951,I14965,I16903,I14945,I16835,I16852,I16818,I15372,I16934,I16869,I15126,I15245,I16886;
DFFARX1 I_0(I15519,I1470,I14965,,,I14948,);
nand I_1(I16804,I16934,I16903);
nand I_2(I14951,I15016,I15245);
not I_3(I14965,I1477);
nor I_4(I16903,I16886,I16869);
nand I_5(I14945,I15372,I15126);
nand I_6(I16835,I14948);
and I_7(I16852,I16835,I14957);
not I_8(I16818,I1477);
DFFARX1 I_9(I12602,I1470,I14965,,,I15372,);
DFFARX1 I_10(I14945,I1470,I16818,,,I16934,);
DFFARX1 I_11(I16852,I1470,I16818,,,I16869,);
not I_12(I15126,I15109);
nor I_13(I15245,I15126);
nor I_14(I16886,I14951,I14948);
endmodule


