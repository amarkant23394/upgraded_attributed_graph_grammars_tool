module test_I6872(I1477,I1470,I6872);
input I1477,I1470;
output I6872;
wire I5625,I5067,I6907,I7269,I5105,I5642;
DFFARX1 I_0(I1470,I5105,,,I5625,);
DFFARX1 I_1(I7269,I1470,I6907,,,I6872,);
DFFARX1 I_2(I5642,I1470,I5105,,,I5067,);
not I_3(I6907,I1477);
DFFARX1 I_4(I5067,I1470,I6907,,,I7269,);
not I_5(I5105,I1477);
not I_6(I5642,I5625);
endmodule


