module test_I12524(I10349,I1477,I10538,I1470,I12524);
input I10349,I1477,I10538,I1470;
output I12524;
wire I10038,I12425,I12442,I11973;
nand I_0(I10038,I10349,I10538);
DFFARX1 I_1(I10038,I1470,I11973,,,I12425,);
not I_2(I12524,I12442);
not I_3(I12442,I12425);
not I_4(I11973,I1477);
endmodule


