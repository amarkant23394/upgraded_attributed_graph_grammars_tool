module test_I3747(I1733,I1477,I1423,I1279,I1470,I1586,I1383,I3747);
input I1733,I1477,I1423,I1279,I1470,I1586,I1383;
output I3747;
wire I1518,I3388,I1750,I1504,I1880,I1603,I1897,I1767;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
or I_2(I1750,I1733,I1279);
nand I_3(I1504,I1767,I1897);
DFFARX1 I_4(I1383,I1470,I1518,,,I1880,);
nand I_5(I1603,I1586,I1423);
DFFARX1 I_6(I1504,I1470,I3388,,,I3747,);
nor I_7(I1897,I1880,I1603);
DFFARX1 I_8(I1750,I1470,I1518,,,I1767,);
endmodule


