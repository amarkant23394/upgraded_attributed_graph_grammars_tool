module test_final(G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,n_452_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15,n4_1_l_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n_452_1_r_15,blif_clk_net_1_r_9,n5_9,G42_1_r_15,);
and I_1(n_572_1_r_15,n17_15,n19_15);
nand I_2(n_573_1_r_15,n15_15,n18_15);
nor I_3(n_549_1_r_15,n21_15,n22_15);
nand I_4(n_569_1_r_15,n15_15,n20_15);
nor I_5(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_6(G42_1_l_15,blif_clk_net_1_r_9,n5_9,ACVQN2_3_r_15,);
nor I_7(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_8(N1_4_r_15,blif_clk_net_1_r_9,n5_9,G199_4_r_15,);
DFFARX1 I_9(n_573_1_l_15,blif_clk_net_1_r_9,n5_9,G214_4_r_15,);
nor I_10(n4_1_l_15,G18_1_l_15,IN_1_1_l_15);
DFFARX1 I_11(n4_1_l_15,blif_clk_net_1_r_9,n5_9,G42_1_l_15,);
not I_12(n15_15,G42_1_l_15);
DFFARX1 I_13(IN_1_3_l_15,blif_clk_net_1_r_9,n5_9,n17_internal_15,);
not I_14(n17_15,n17_internal_15);
DFFARX1 I_15(IN_2_3_l_15,blif_clk_net_1_r_9,n5_9,n30_15,);
nor I_16(n_572_1_l_15,G15_1_l_15,IN_7_1_l_15);
DFFARX1 I_17(n_572_1_l_15,blif_clk_net_1_r_9,n5_9,n14_internal_15,);
not I_18(n14_15,n14_internal_15);
nand I_19(N1_4_r_15,n25_15,n26_15);
or I_20(n_573_1_l_15,IN_5_1_l_15,IN_9_1_l_15);
nor I_21(n18_15,IN_9_1_l_15,IN_10_1_l_15);
nand I_22(n19_15,n27_15,n28_15);
nand I_23(n20_15,IN_4_3_l_15,n30_15);
not I_24(n21_15,n20_15);
and I_25(n22_15,n17_15,n_572_1_l_15);
nor I_26(n23_15,G18_1_l_15,IN_5_1_l_15);
or I_27(n24_15,IN_9_1_l_15,IN_10_1_l_15);
or I_28(n25_15,G18_1_l_15,n_573_1_l_15);
nand I_29(n26_15,n19_15,n23_15);
not I_30(n27_15,IN_10_1_l_15);
nand I_31(n28_15,IN_4_1_l_15,n29_15);
not I_32(n29_15,G15_1_l_15);
DFFARX1 I_33(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_34(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_35(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_36(n_549_1_r_9,n17_9,n18_9);
or I_37(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_38(n_452_1_r_9,n26_9,n25_9);
nor I_39(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_40(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_41(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_42(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_43(N3_2_l_9,n22_9,G199_4_r_15);
not I_44(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_45(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_46(n16_9,n27_9);
DFFARX1 I_47(n_573_1_r_15,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_48(n15_9,n26_9);
DFFARX1 I_49(n_572_1_r_15,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_50(n29_9,n29_internal_9);
and I_51(N1_4_l_9,n24_9,n_572_1_r_15);
DFFARX1 I_52(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_53(G214_4_r_15,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_54(n28_9,n28_internal_9);
nor I_55(n4_1_r_9,n27_9,n26_9);
nor I_56(N3_2_r_9,n15_9,n21_9);
nor I_57(N1_4_r_9,n16_9,n21_9);
nor I_58(n_42_2_l_9,n_549_1_r_15,n_266_and_0_3_r_15);
not I_59(n17_9,n_452_1_r_9);
nand I_60(n18_9,n27_9,n15_9);
nor I_61(n19_9,n29_9,n20_9);
not I_62(n20_9,G42_1_r_15);
and I_63(n21_9,n23_9,G42_1_r_15);
nand I_64(n22_9,n_266_and_0_3_r_15,G42_1_r_15);
nor I_65(n23_9,n29_9,n28_9);
nand I_66(n24_9,n_569_1_r_15,ACVQN2_3_r_15);
endmodule


