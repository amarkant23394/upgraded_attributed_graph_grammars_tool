module test_I15109(I1477,I10627,I1470,I10630,I12636,I15109);
input I1477,I10627,I1470,I10630,I12636;
output I15109;
wire I12619,I12670,I12783,I12584,I12735,I12653;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
DFFARX1 I_2(I12735,I1470,I12619,,,I12783,);
and I_3(I12584,I12670,I12783);
not I_4(I15109,I12584);
DFFARX1 I_5(I10630,I1470,I12619,,,I12735,);
and I_6(I12653,I12636,I10627);
endmodule


