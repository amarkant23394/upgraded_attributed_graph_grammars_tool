module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_8_r_6,n9_6,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N1371_0_r_6,n30_6,n33_6);
nor I_36(N1508_0_r_6,n33_6,n44_6);
not I_37(N1372_1_r_6,n41_6);
nor I_38(N1508_1_r_6,n40_6,n41_6);
nor I_39(N1507_6_r_6,n39_6,n45_6);
nor I_40(N1508_6_r_6,n37_6,n38_6);
nor I_41(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_42(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_43(N6147_9_r_6,n32_6,n33_6);
nor I_44(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_45(I_BUFF_1_9_r_6,n37_6);
not I_46(N1372_10_r_6,n43_6);
nor I_47(N1508_10_r_6,n42_6,n43_6);
nor I_48(N3_8_r_6,n36_6,N1371_0_r_4);
not I_49(n9_6,blif_reset_net_8_r_6);
nor I_50(n30_6,n53_6,n_549_7_r_4);
not I_51(n31_6,n36_6);
nor I_52(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_53(n33_6,N1371_0_r_4);
not I_54(n34_6,n35_6);
nand I_55(n35_6,n49_6,N1507_6_r_4);
nand I_56(n36_6,n51_6,n_569_7_r_4);
nand I_57(n37_6,n54_6,N1507_6_r_4);
or I_58(n38_6,n35_6,n39_6);
nor I_59(n39_6,n40_6,n45_6);
and I_60(n40_6,n46_6,n47_6);
nand I_61(n41_6,n30_6,n31_6);
nor I_62(n42_6,n34_6,n40_6);
nand I_63(n43_6,n30_6,N1371_0_r_4);
nor I_64(n44_6,n31_6,n40_6);
nor I_65(n45_6,n35_6,n36_6);
nor I_66(n46_6,N1371_0_r_4,n_572_7_r_4);
or I_67(n47_6,n48_6,n_549_7_r_4);
nor I_68(n48_6,N6134_9_r_4,N1508_6_r_4);
and I_69(n49_6,n50_6,n_452_7_r_4);
nand I_70(n50_6,n51_6,n52_6);
nand I_71(n51_6,G42_7_r_4,n_572_7_r_4);
not I_72(n52_6,n_569_7_r_4);
nor I_73(n53_6,N1508_6_r_4,G42_7_r_4);
or I_74(n54_6,N1508_6_r_4,G42_7_r_4);
endmodule


