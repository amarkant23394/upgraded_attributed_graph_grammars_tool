module test_I7782(I3957,I1477,I6442,I1470,I6623,I3972,I7782);
input I3957,I1477,I6442,I1470,I6623,I3972;
output I7782;
wire I6781,I7765,I6722,I6640,I6329,I6688,I6312,I6705,I6291,I6303,I7748;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
nor I_1(I7765,I7748,I6303);
or I_2(I6722,I6705,I6640);
and I_3(I6640,I6442,I6623);
not I_4(I6329,I1477);
DFFARX1 I_5(I1470,I6329,,,I6688,);
and I_6(I7782,I7765,I6312);
DFFARX1 I_7(I6722,I1470,I6329,,,I6312,);
and I_8(I6705,I6688,I3972);
DFFARX1 I_9(I6705,I1470,I6329,,,I6291,);
DFFARX1 I_10(I6781,I1470,I6329,,,I6303,);
not I_11(I7748,I6291);
endmodule


