module test_I9559(I8202,I1477,I8561,I1470,I9559);
input I8202,I1477,I8561,I1470;
output I9559;
wire I9508,I9542,I8216,I8199,I8184,I9525,I9491;
nand I_0(I9508,I8199,I8202);
DFFARX1 I_1(I9525,I1470,I9491,,,I9542,);
not I_2(I8216,I1477);
DFFARX1 I_3(I1470,I8216,,,I8199,);
not I_4(I9559,I9542);
DFFARX1 I_5(I8561,I1470,I8216,,,I8184,);
and I_6(I9525,I9508,I8184);
not I_7(I9491,I1477);
endmodule


