module test_I1535(I1455,I1535);
input I1455;
output I1535;
wire ;
not I_0(I1535,I1455);
endmodule


