module test_I17628(I13908,I13761,I1470,I15611,I16007,I17628);
input I13908,I13761,I1470,I15611,I16007;
output I17628;
wire I15713,I17611,I13743,I15730,I15832,I15576,I14162,I15628,I16052,I13749,I15573,I17594,I15591,I16069;
not I_0(I15713,I13761);
nor I_1(I17611,I17594,I15591);
DFFARX1 I_2(I1470,,,I13743,);
and I_3(I17628,I17611,I15573);
not I_4(I15730,I15713);
nand I_5(I15832,I15628,I13749);
DFFARX1 I_6(I16007,I1470,I15611,,,I15576,);
DFFARX1 I_7(I1470,,,I14162,);
not I_8(I15628,I13743);
DFFARX1 I_9(I1470,I15611,,,I16052,);
nand I_10(I13749,I14162,I13908);
nand I_11(I15573,I15832,I15730);
not I_12(I17594,I15576);
nor I_13(I15591,I16069,I15832);
not I_14(I16069,I16052);
endmodule


