module test_final(IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_5_r_0,blif_reset_net_5_r_0,N1371_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0);
input IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_5_r_0,blif_reset_net_5_r_0;
output N1371_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0;
wire N1371_0_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_102_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4,n_431_5_r_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,N1508_0_r_0,n_102_5_r_0,N3_8_l_0,n5_0,n40_0,n4_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0;
nor I_0(N1371_0_r_4,n25_4,n29_4);
nor I_1(N1508_0_r_4,n25_4,n32_4);
nor I_2(N6147_2_r_4,n24_4,n31_4);
or I_3(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_4(n_431_5_r_4,blif_clk_net_5_r_0,n5_0,G78_5_r_4,);
nand I_5(n_576_5_r_4,n22_4,n23_4);
nand I_6(n_102_5_r_4,n34_4,n35_4);
nand I_7(n_547_5_r_4,n26_4,n27_4);
nor I_8(N1507_6_r_4,n27_4,n30_4);
nor I_9(N1508_6_r_4,n30_4,n33_4);
nand I_10(n_431_5_r_4,n_102_5_r_4,n28_4);
nor I_11(n22_4,n24_4,n25_4);
nor I_12(n23_4,IN_1_3_l_4,n37_4);
not I_13(n24_4,n_102_5_r_4);
nand I_14(n25_4,IN_1_1_l_4,IN_2_1_l_4);
nor I_15(n26_4,n23_4,n24_4);
not I_16(n27_4,n25_4);
nand I_17(n28_4,n23_4,n29_4);
nor I_18(n29_4,IN_3_1_l_4,n25_4);
not I_19(n30_4,n29_4);
nor I_20(n31_4,N1371_0_r_4,n32_4);
nor I_21(n32_4,n23_4,n29_4);
nand I_22(n33_4,n23_4,n24_4);
nor I_23(n34_4,IN_1_2_l_4,IN_2_2_l_4);
or I_24(n35_4,IN_5_2_l_4,n36_4);
nor I_25(n36_4,IN_3_2_l_4,IN_4_2_l_4);
or I_26(n37_4,IN_2_3_l_4,IN_3_3_l_4);
nor I_27(N1371_0_r_0,n24_0,n25_0);
not I_28(N1508_0_r_0,n25_0);
nor I_29(N6147_2_r_0,n28_0,n29_0);
nand I_30(n_429_or_0_5_r_0,n4_0,n25_0);
DFFARX1 I_31(n4_0,blif_clk_net_5_r_0,n5_0,G78_5_r_0,);
nand I_32(n_576_5_r_0,n23_0,n24_0);
not I_33(n_102_5_r_0,n40_0);
nand I_34(n_547_5_r_0,n26_0,n27_0);
nor I_35(N1507_6_r_0,n_102_5_r_0,n37_0);
nor I_36(N1508_6_r_0,n25_0,n33_0);
and I_37(N3_8_l_0,n32_0,n_429_or_0_5_r_4);
not I_38(n5_0,blif_reset_net_5_r_0);
DFFARX1 I_39(N3_8_l_0,blif_clk_net_5_r_0,n5_0,n40_0,);
not I_40(n4_0,n31_0);
nor I_41(n23_0,n40_0,n25_0);
and I_42(n24_0,n4_0,n39_0);
nand I_43(n25_0,N1508_0_r_4,n_547_5_r_4);
nor I_44(n26_0,n40_0,n24_0);
nor I_45(n27_0,G78_5_r_4,n_576_5_r_4);
nor I_46(n28_0,n25_0,N6147_2_r_4);
nand I_47(n29_0,n_102_5_r_0,n30_0);
nand I_48(n30_0,n27_0,n31_0);
nand I_49(n31_0,N1508_6_r_4,n_429_or_0_5_r_4);
nand I_50(n32_0,N6147_2_r_4,G78_5_r_4);
nand I_51(n33_0,n34_0,n35_0);
nand I_52(n34_0,n_102_5_r_0,n36_0);
not I_53(n35_0,N6147_2_r_4);
not I_54(n36_0,n27_0);
nor I_55(n37_0,n36_0,n38_0);
nand I_56(n38_0,N1508_0_r_0,n35_0);
or I_57(n39_0,N1507_6_r_4,N1508_0_r_4);
endmodule


