module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_7_r_3,n10_3,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_7_r_3,n10_3,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
not I_40(N1372_1_r_3,n40_3);
nor I_41(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_42(N1507_6_r_3,n31_3,n42_3);
nor I_43(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_44(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_45(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_46(n_573_7_r_3,n30_3,n31_3);
nor I_47(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_48(n_569_7_r_3,n30_3,n32_3);
nor I_49(n_452_7_r_3,n35_3,N1371_0_r_16);
not I_50(N6147_9_r_3,n32_3);
nor I_51(N6134_9_r_3,n36_3,n37_3);
not I_52(I_BUFF_1_9_r_3,n45_3);
nor I_53(n4_7_r_3,I_BUFF_1_9_r_3,N1371_0_r_16);
not I_54(n10_3,blif_reset_net_7_r_3);
not I_55(n30_3,n39_3);
not I_56(n31_3,n35_3);
nand I_57(n32_3,n41_3,n_569_7_r_16);
nor I_58(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_59(n34_3,n46_3,N1372_1_r_16);
nor I_60(n35_3,n43_3,n44_3);
not I_61(n36_3,n34_3);
nor I_62(n37_3,N6147_9_r_3,N1371_0_r_16);
or I_63(n38_3,n_572_7_r_3,n34_3);
nor I_64(n39_3,n44_3,N1507_6_r_16);
nand I_65(n40_3,n39_3,N1371_0_r_16);
nand I_66(n41_3,G42_7_r_16,n_572_7_r_16);
nor I_67(n42_3,n34_3,n45_3);
not I_68(n43_3,N1371_0_r_16);
nor I_69(n44_3,N1508_0_r_16,N1508_6_r_16);
nand I_70(n45_3,n49_3,n50_3);
and I_71(n46_3,n47_3,N6147_2_r_16);
nand I_72(n47_3,n41_3,n48_3);
not I_73(n48_3,n_569_7_r_16);
nor I_74(n49_3,N1508_1_r_16,n_452_7_r_16);
or I_75(n50_3,n51_3,N1372_1_r_16);
nor I_76(n51_3,n_573_7_r_16,N1508_0_r_16);
endmodule


