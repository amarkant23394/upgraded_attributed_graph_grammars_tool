module test_I5385(I3422,I1477,I3521,I3846,I1470,I3365,I5300,I5385);
input I3422,I1477,I3521,I3846,I1470,I3365,I5300;
output I5385;
wire I5266,I3388,I5351,I3362,I5334,I3380,I5317,I5249,I5105;
not I_0(I5266,I5249);
not I_1(I3388,I1477);
DFFARX1 I_2(I5334,I1470,I5105,,,I5351,);
DFFARX1 I_3(I3422,I1470,I3388,,,I3362,);
nor I_4(I5385,I5351,I5266);
or I_5(I5334,I5317,I3362);
nand I_6(I3380,I3521,I3846);
and I_7(I5317,I5300,I3365);
not I_8(I5249,I3380);
not I_9(I5105,I1477);
endmodule


