module test_I8090(I1477,I1470,I4068,I8090);
input I1477,I1470,I4068;
output I8090;
wire I3975,I3966,I3954,I7570,I6309,I6442,I6329,I6493,I4034,I6459;
nor I_0(I3975,I4034);
or I_1(I3966,I4068,I4034);
DFFARX1 I_2(I6309,I1470,I7570,,,I8090,);
not I_3(I3954,I4068);
not I_4(I7570,I1477);
nand I_5(I6309,I6493,I6459);
nor I_6(I6442,I3975,I3954);
not I_7(I6329,I1477);
DFFARX1 I_8(I3966,I1470,I6329,,,I6493,);
DFFARX1 I_9(I1470,,,I4034,);
not I_10(I6459,I6442);
endmodule


