module test_I16798(I1477,I14945,I15109,I15016,I14942,I1470,I15519,I15245,I16798);
input I1477,I14945,I15109,I15016,I14942,I1470,I15519,I15245;
output I16798;
wire I14948,I14951,I14965,I17047,I17013,I17030,I16968,I14939,I16818,I15341,I14930,I16934,I16951,I16886;
DFFARX1 I_0(I15519,I1470,I14965,,,I14948,);
nand I_1(I14951,I15016,I15245);
not I_2(I14965,I1477);
DFFARX1 I_3(I17030,I1470,I16818,,,I17047,);
nand I_4(I17013,I14942,I14939);
and I_5(I17030,I17013,I14930);
nor I_6(I16968,I16886,I16951);
DFFARX1 I_7(I15016,I1470,I14965,,,I14939,);
not I_8(I16818,I1477);
nand I_9(I16798,I17047,I16968);
DFFARX1 I_10(I1470,I14965,,,I15341,);
and I_11(I14930,I15109,I15341);
DFFARX1 I_12(I14945,I1470,I16818,,,I16934,);
not I_13(I16951,I16934);
nor I_14(I16886,I14951,I14948);
endmodule


