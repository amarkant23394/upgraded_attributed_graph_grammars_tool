module test_I16229(I14667,I1477,I14520,I1470,I14588,I16229);
input I14667,I1477,I14520,I1470,I14588;
output I16229;
wire I14901,I14777,I14537,I14344,I14808,I16534,I14347,I16240,I16644,I16551,I14335,I14715,I14370;
DFFARX1 I_0(I14808,I1470,I14370,,,I14901,);
or I_1(I14777,I14667,I14588);
DFFARX1 I_2(I14520,I1470,I14370,,,I14537,);
nand I_3(I14344,I14537,I14715);
DFFARX1 I_4(I1470,I14370,,,I14808,);
DFFARX1 I_5(I14335,I1470,I16240,,,I16534,);
DFFARX1 I_6(I14777,I1470,I14370,,,I14347,);
nor I_7(I16229,I16644,I16551);
not I_8(I16240,I1477);
DFFARX1 I_9(I14347,I1470,I16240,,,I16644,);
and I_10(I16551,I16534,I14344);
and I_11(I14335,I14808,I14901);
not I_12(I14715,I14667);
not I_13(I14370,I1477);
endmodule


