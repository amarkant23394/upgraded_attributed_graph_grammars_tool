module Benchmark_testing25000(I1579,I1587,I1595,I1603,I1611,I1619,I1627,I1635,I1643,I1651,I1659,I1667,I1675,I1683,I1691,I1699,I1707,I1715,I1723,I1731,I1739,I1747,I1755,I1763,I1771,I1779,I1787,I1795,I1803,I1811,I1819,I1827,I1835,I1843,I1851,I1859,I1867,I1875,I1883,I1891,I1899,I1907,I1915,I1923,I1931,I1939,I1947,I1955,I1963,I1971,I1979,I1987,I1995,I2003,I2011,I2019,I2027,I2035,I2043,I2051,I2059,I2067,I2075,I2083,I2091,I2099,I2107,I2115,I2123,I2131,I2139,I2147,I2155,I2163,I2171,I2179,I2187,I2195,I2203,I2211,I2219,I2227,I2235,I2243,I2251,I2259,I2267,I2275,I2283,I2291,I2299,I2307,I2315,I2323,I2331,I2339,I2347,I2355,I2363,I2371,I2379,I2387,I2395,I2403,I2411,I2419,I2427,I2435,I2443,I2451,I2459,I2467,I2475,I2483,I2491,I2499,I2507,I2515,I2523,I2531,I2539,I2547,I2555,I2563,I2571,I2579,I2587,I2595,I2603,I2611,I2619,I2627,I2635,I2643,I2651,I2659,I2667,I2675,I2683,I2691,I2699,I2707,I2715,I2723,I2731,I2739,I2747,I2755,I2763,I2771,I2779,I2787,I2795,I2803,I2811,I2819,I2827,I2835,I2843,I2851,I2859,I2867,I2875,I2883,I2891,I2898,I2905,I120433,I120445,I120412,I120418,I120421,I120427,I120415,I120430,I120442,I120439,I120424,I120436,I127352,I127364,I127331,I127337,I127340,I127346,I127334,I127349,I127361,I127358,I127343,I127355,I158594,I158624,I158600,I158612,I158615,I158618,I158621,I158606,I158609,I158597,I158627,I158603,I193218,I193209,I193206,I193230,I193212,I193221,I193227,I193224,I193215,I278070,I278085,I278073,I278088,I278079,I278100,I278076,I278097,I278091,I278082,I278094,I289359,I289353,I289356,I289341,I289344,I289347,I289365,I289371,I289368,I289350,I289362,I354982,I354967,I354964,I354985,I354961,I354970,I354979,I354976,I354973,I378399,I378387,I378411,I378393,I378396,I378405,I378414,I378402,I378390,I378420,I378417,I378408,I433160,I433127,I433130,I433139,I433151,I433133,I433136,I433142,I433145,I433148,I433157,I433154,I442221,I442188,I442191,I442200,I442212,I442194,I442197,I442203,I442206,I442209,I442218,I442215,I444312,I444279,I444282,I444291,I444303,I444285,I444288,I444294,I444297,I444300,I444309,I444306);
input I1579,I1587,I1595,I1603,I1611,I1619,I1627,I1635,I1643,I1651,I1659,I1667,I1675,I1683,I1691,I1699,I1707,I1715,I1723,I1731,I1739,I1747,I1755,I1763,I1771,I1779,I1787,I1795,I1803,I1811,I1819,I1827,I1835,I1843,I1851,I1859,I1867,I1875,I1883,I1891,I1899,I1907,I1915,I1923,I1931,I1939,I1947,I1955,I1963,I1971,I1979,I1987,I1995,I2003,I2011,I2019,I2027,I2035,I2043,I2051,I2059,I2067,I2075,I2083,I2091,I2099,I2107,I2115,I2123,I2131,I2139,I2147,I2155,I2163,I2171,I2179,I2187,I2195,I2203,I2211,I2219,I2227,I2235,I2243,I2251,I2259,I2267,I2275,I2283,I2291,I2299,I2307,I2315,I2323,I2331,I2339,I2347,I2355,I2363,I2371,I2379,I2387,I2395,I2403,I2411,I2419,I2427,I2435,I2443,I2451,I2459,I2467,I2475,I2483,I2491,I2499,I2507,I2515,I2523,I2531,I2539,I2547,I2555,I2563,I2571,I2579,I2587,I2595,I2603,I2611,I2619,I2627,I2635,I2643,I2651,I2659,I2667,I2675,I2683,I2691,I2699,I2707,I2715,I2723,I2731,I2739,I2747,I2755,I2763,I2771,I2779,I2787,I2795,I2803,I2811,I2819,I2827,I2835,I2843,I2851,I2859,I2867,I2875,I2883,I2891,I2898,I2905;
output I120433,I120445,I120412,I120418,I120421,I120427,I120415,I120430,I120442,I120439,I120424,I120436,I127352,I127364,I127331,I127337,I127340,I127346,I127334,I127349,I127361,I127358,I127343,I127355,I158594,I158624,I158600,I158612,I158615,I158618,I158621,I158606,I158609,I158597,I158627,I158603,I193218,I193209,I193206,I193230,I193212,I193221,I193227,I193224,I193215,I278070,I278085,I278073,I278088,I278079,I278100,I278076,I278097,I278091,I278082,I278094,I289359,I289353,I289356,I289341,I289344,I289347,I289365,I289371,I289368,I289350,I289362,I354982,I354967,I354964,I354985,I354961,I354970,I354979,I354976,I354973,I378399,I378387,I378411,I378393,I378396,I378405,I378414,I378402,I378390,I378420,I378417,I378408,I433160,I433127,I433130,I433139,I433151,I433133,I433136,I433142,I433145,I433148,I433157,I433154,I442221,I442188,I442191,I442200,I442212,I442194,I442197,I442203,I442206,I442209,I442218,I442215,I444312,I444279,I444282,I444291,I444303,I444285,I444288,I444294,I444297,I444300,I444309,I444306;
wire I1579,I1587,I1595,I1603,I1611,I1619,I1627,I1635,I1643,I1651,I1659,I1667,I1675,I1683,I1691,I1699,I1707,I1715,I1723,I1731,I1739,I1747,I1755,I1763,I1771,I1779,I1787,I1795,I1803,I1811,I1819,I1827,I1835,I1843,I1851,I1859,I1867,I1875,I1883,I1891,I1899,I1907,I1915,I1923,I1931,I1939,I1947,I1955,I1963,I1971,I1979,I1987,I1995,I2003,I2011,I2019,I2027,I2035,I2043,I2051,I2059,I2067,I2075,I2083,I2091,I2099,I2107,I2115,I2123,I2131,I2139,I2147,I2155,I2163,I2171,I2179,I2187,I2195,I2203,I2211,I2219,I2227,I2235,I2243,I2251,I2259,I2267,I2275,I2283,I2291,I2299,I2307,I2315,I2323,I2331,I2339,I2347,I2355,I2363,I2371,I2379,I2387,I2395,I2403,I2411,I2419,I2427,I2435,I2443,I2451,I2459,I2467,I2475,I2483,I2491,I2499,I2507,I2515,I2523,I2531,I2539,I2547,I2555,I2563,I2571,I2579,I2587,I2595,I2603,I2611,I2619,I2627,I2635,I2643,I2651,I2659,I2667,I2675,I2683,I2691,I2699,I2707,I2715,I2723,I2731,I2739,I2747,I2755,I2763,I2771,I2779,I2787,I2795,I2803,I2811,I2819,I2827,I2835,I2843,I2851,I2859,I2867,I2875,I2883,I2891,I2898,I2905,I2946,I2963,I275784,I275793,I2980,I2997,I275787,I3014,I275790,I3031,I3048,I2914,I275796,I2929,I3093,I275802,I275778,I3110,I275805,I3127,I275781,I3144,I3161,I2911,I3192,I3209,I2923,I3240,I2920,I3271,I3288,I2926,I3319,I3336,I275775,I3353,I3370,I275799,I3387,I3404,I2908,I3435,I3452,I2917,I2935,I2932,I2938,I3558,I3575,I435245,I435251,I3592,I3609,I435221,I3626,I435242,I3643,I3660,I3526,I435224,I3541,I3705,I435233,I435227,I3722,I3739,I435248,I435239,I3756,I3773,I3523,I3804,I3821,I3535,I3852,I3532,I3883,I3900,I3538,I3931,I3948,I435218,I435236,I3965,I3982,I435230,I3999,I4016,I3520,I4047,I4064,I3529,I3547,I3544,I3550,I4170,I4187,I145680,I145686,I4204,I4221,I145674,I4238,I145701,I4255,I4272,I4138,I145683,I4153,I4317,I145704,I145707,I4334,I145692,I4351,I145677,I145698,I4368,I4385,I4135,I4416,I4433,I4147,I4464,I4144,I4495,I4512,I4150,I4543,I4560,I145695,I4577,I4594,I145689,I4611,I4628,I4132,I4659,I4676,I4141,I4159,I4156,I4162,I4782,I4799,I154520,I154526,I4816,I4833,I154514,I4850,I154541,I4867,I4884,I4750,I154523,I4765,I4929,I154544,I154547,I4946,I154532,I4963,I154517,I154538,I4980,I4997,I4747,I5028,I5045,I4759,I5076,I4756,I5107,I5124,I4762,I5155,I5172,I154535,I5189,I5206,I154529,I5223,I5240,I4744,I5271,I5288,I4753,I4771,I4768,I4774,I5394,I5411,I360920,I5428,I5445,I360923,I5462,I360932,I5479,I5496,I5362,I360917,I5377,I5541,I360914,I5558,I360926,I5575,I360911,I5592,I5609,I5359,I5640,I5657,I5371,I5688,I5368,I5719,I5736,I5374,I5767,I5784,I5801,I5818,I360935,I360929,I5835,I5852,I5356,I5883,I5900,I5365,I5383,I5380,I5386,I6006,I6023,I23206,I23224,I6040,I6057,I23215,I6074,I23209,I6091,I6108,I5974,I23212,I5989,I6153,I23227,I6170,I23218,I6187,I23221,I6204,I6221,I5971,I6252,I6269,I5983,I6300,I5980,I6331,I6348,I5986,I6379,I6396,I6413,I23230,I6430,I23233,I6447,I6464,I5968,I6495,I6512,I5977,I5995,I5992,I5998,I6618,I6635,I115380,I115386,I6652,I6669,I115392,I6686,I115383,I6703,I6720,I6586,I115407,I6601,I6765,I115404,I115389,I6782,I115413,I6799,I115401,I115410,I6816,I6833,I6583,I6864,I6881,I6595,I6912,I6592,I6943,I6960,I6598,I6991,I7008,I115395,I7025,I7042,I115398,I7059,I7076,I6580,I7107,I7124,I6589,I6607,I6604,I6610,I7230,I7247,I272724,I272733,I7264,I7281,I272727,I7298,I272730,I7315,I7332,I7198,I272736,I7213,I7377,I272742,I272718,I7394,I272745,I7411,I272721,I7428,I7445,I7195,I7476,I7493,I7207,I7524,I7204,I7555,I7572,I7210,I7603,I7620,I272715,I7637,I7654,I272739,I7671,I7688,I7192,I7719,I7736,I7201,I7219,I7216,I7222,I7842,I7859,I184166,I184151,I7876,I7893,I184148,I7910,I184160,I7927,I7944,I7810,I7825,I7989,I184157,I184169,I8006,I184154,I8023,I184163,I8040,I8057,I7807,I8088,I8105,I7819,I8136,I7816,I8167,I8184,I7822,I8215,I8232,I8249,I8266,I184145,I8283,I8300,I7804,I8331,I8348,I7813,I7831,I7828,I7834,I8454,I8471,I252069,I252078,I8488,I8505,I252072,I8522,I252075,I8539,I8556,I8422,I252081,I8437,I8601,I252087,I252063,I8618,I252090,I8635,I252066,I8652,I8669,I8419,I8700,I8717,I8431,I8748,I8428,I8779,I8796,I8434,I8827,I8844,I252060,I8861,I8878,I252084,I8895,I8912,I8416,I8943,I8960,I8425,I8443,I8440,I8446,I9066,I9083,I403343,I403358,I9100,I9117,I9134,I403349,I9151,I9168,I9034,I403355,I9049,I9213,I403346,I9230,I9247,I403352,I403361,I9264,I9281,I9031,I9312,I9329,I9043,I9360,I9040,I9391,I9408,I9046,I9439,I9456,I403364,I9473,I9490,I403367,I9507,I9524,I9028,I9555,I9572,I9037,I9055,I9052,I9058,I9678,I9695,I227651,I227657,I9712,I9729,I227675,I9746,I227654,I9763,I9780,I9646,I227663,I9661,I9825,I227666,I227660,I9842,I227672,I9859,I9876,I9893,I9643,I9924,I9941,I9655,I9972,I9652,I10003,I10020,I9658,I10051,I10068,I227648,I227669,I10085,I10102,I10119,I10136,I9640,I10167,I10184,I9649,I9667,I9664,I9670,I10290,I10307,I343665,I10324,I10341,I343668,I10358,I343677,I10375,I10392,I10258,I343662,I10273,I10437,I343659,I10454,I343671,I10471,I343656,I10488,I10505,I10255,I10536,I10553,I10267,I10584,I10264,I10615,I10632,I10270,I10663,I10680,I10697,I10714,I343680,I343674,I10731,I10748,I10252,I10779,I10796,I10261,I10279,I10276,I10282,I10902,I10919,I21778,I21796,I10936,I10953,I21787,I10970,I21781,I10987,I11004,I10870,I21784,I10885,I11049,I21799,I11066,I21790,I11083,I21793,I11100,I11117,I10867,I11148,I11165,I10879,I11196,I10876,I11227,I11244,I10882,I11275,I11292,I11309,I21802,I11326,I21805,I11343,I11360,I10864,I11391,I11408,I10873,I10891,I10888,I10894,I11514,I11531,I191833,I191818,I11548,I11565,I191815,I11582,I191827,I11599,I11616,I11482,I11497,I11661,I191824,I191836,I11678,I191821,I11695,I191830,I11712,I11729,I11479,I11760,I11777,I11491,I11808,I11488,I11839,I11856,I11494,I11887,I11904,I11921,I11938,I191812,I11955,I11972,I11476,I12003,I12020,I11485,I11503,I11500,I11506,I12126,I12143,I324030,I12160,I12177,I324033,I12194,I324042,I12211,I12228,I12094,I324027,I12109,I12273,I324024,I12290,I324036,I12307,I324021,I12324,I12341,I12091,I12372,I12389,I12103,I12420,I12100,I12451,I12468,I12106,I12499,I12516,I12533,I12550,I324045,I324039,I12567,I12584,I12088,I12615,I12632,I12097,I12115,I12112,I12118,I12738,I12755,I341285,I12772,I12789,I341288,I12806,I341297,I12823,I12840,I12706,I341282,I12721,I12885,I341279,I12902,I341291,I12919,I341276,I12936,I12953,I12703,I12984,I13001,I12715,I13032,I12712,I13063,I13080,I12718,I13111,I13128,I13145,I13162,I341300,I341294,I13179,I13196,I12700,I13227,I13244,I12709,I12727,I12724,I12730,I13350,I13367,I44913,I44934,I13384,I13401,I44898,I13418,I44901,I13435,I13452,I13318,I44931,I13333,I13497,I44904,I44910,I13514,I44928,I13531,I44916,I44925,I13548,I13565,I13315,I13596,I13613,I13327,I13644,I13324,I13675,I13692,I13330,I13723,I13740,I44907,I13757,I44919,I13774,I44922,I13791,I13808,I13312,I13839,I13856,I13321,I13339,I13336,I13342,I13959,I13976,I400632,I13993,I400635,I400638,I14010,I14027,I14044,I14061,I400626,I14078,I14095,I14112,I400644,I14129,I400623,I14146,I14163,I14180,I13927,I14211,I14228,I14245,I14262,I400641,I14279,I14296,I14313,I13924,I14344,I13951,I14375,I400647,I400629,I14392,I14409,I14426,I14443,I13942,I14474,I14491,I13930,I13948,I14536,I14553,I13933,I14584,I13939,I13945,I13936,I14673,I14690,I229919,I14707,I229895,I229907,I14724,I14741,I14758,I14775,I14792,I229892,I14809,I14826,I229916,I229898,I14843,I229910,I14860,I14877,I14894,I14641,I14925,I14942,I229901,I14959,I14976,I229904,I14993,I15010,I15027,I14638,I15058,I14665,I15089,I15106,I229913,I15123,I15140,I15157,I14656,I15188,I15205,I14644,I14662,I15250,I15267,I14647,I15298,I14653,I14659,I14650,I15387,I15404,I438018,I15421,I438009,I438012,I15438,I15455,I15472,I15489,I438006,I15506,I438033,I15523,I15540,I438024,I15557,I438021,I15574,I15591,I15608,I15355,I15639,I15656,I438030,I15673,I15690,I438036,I438027,I15707,I15724,I15741,I15352,I15772,I15379,I15803,I438015,I438039,I15820,I15837,I15854,I15871,I15370,I15902,I15919,I15358,I15376,I15964,I15981,I15361,I16012,I15367,I15373,I15364,I16101,I16118,I149086,I16135,I149098,I149104,I16152,I16169,I16186,I16203,I149077,I16220,I149101,I16237,I16254,I149083,I149074,I16271,I149092,I16288,I16305,I16322,I16069,I16353,I16370,I149095,I16387,I16404,I149080,I16421,I16438,I16455,I16066,I16486,I16093,I16517,I16534,I149107,I16551,I149089,I16568,I16585,I16084,I16616,I16633,I16072,I16090,I16678,I16695,I16075,I16726,I16081,I16087,I16078,I16815,I16832,I353795,I16849,I353783,I353774,I16866,I16883,I16900,I16917,I16934,I353789,I16951,I16968,I353771,I353780,I16985,I353786,I17002,I17019,I17036,I16783,I17067,I17084,I17101,I17118,I17135,I17152,I17169,I16780,I17200,I16807,I17231,I353777,I17248,I353792,I17265,I17282,I17299,I16798,I17330,I17347,I16786,I16804,I17392,I17409,I16789,I17440,I16795,I16801,I16792,I17529,I17546,I383585,I17563,I383567,I383558,I17580,I17597,I17614,I17631,I383579,I17648,I383588,I17665,I17682,I383555,I17699,I383561,I17716,I17733,I17750,I17497,I17781,I17798,I383564,I17815,I17832,I383582,I383573,I17849,I17866,I17883,I17494,I17914,I17521,I17945,I383570,I17962,I17979,I383576,I17996,I18013,I17512,I18044,I18061,I17500,I17518,I18106,I18123,I17503,I18154,I17509,I17515,I17506,I18243,I18260,I45680,I18277,I45701,I18294,I18311,I18328,I18345,I45695,I18362,I45707,I18379,I18396,I45683,I45698,I18413,I45692,I18430,I18447,I18464,I18211,I18495,I18512,I45704,I18529,I18546,I45686,I45710,I18563,I18580,I18597,I18208,I18628,I18235,I18659,I45689,I18676,I45713,I18693,I45716,I18710,I18727,I18226,I18758,I18775,I18214,I18232,I18820,I18837,I18217,I18868,I18223,I18229,I18220,I18957,I18974,I200882,I18991,I200888,I200873,I19008,I19025,I19042,I19059,I19076,I200891,I19093,I19110,I200885,I200879,I19127,I200876,I19144,I19161,I19178,I18925,I19209,I19226,I19243,I19260,I200897,I19277,I19294,I19311,I18922,I19342,I18949,I19373,I200894,I19390,I19407,I19424,I19441,I18940,I19472,I19489,I18928,I18946,I19534,I19551,I18931,I19582,I18937,I18943,I18934,I19671,I19688,I382939,I19705,I382921,I382912,I19722,I19739,I19756,I19773,I382933,I19790,I382942,I19807,I19824,I382909,I19841,I382915,I19858,I19875,I19892,I19639,I19923,I19940,I382918,I19957,I19974,I382936,I382927,I19991,I20008,I20025,I19636,I20056,I19663,I20087,I382924,I20104,I20121,I382930,I20138,I20155,I19654,I20186,I20203,I19642,I19660,I20248,I20265,I19645,I20296,I19651,I19657,I19648,I20385,I20402,I321520,I20419,I321535,I321505,I20436,I20453,I20470,I20487,I321517,I20504,I321508,I20521,I20538,I321529,I321532,I20555,I321511,I20572,I20589,I20606,I20353,I20637,I20654,I321514,I20671,I20688,I20705,I20722,I20739,I20350,I20770,I20377,I20801,I321526,I20818,I321523,I20835,I20852,I20869,I20368,I20900,I20917,I20356,I20374,I20962,I20979,I20359,I21010,I20365,I20371,I20362,I21099,I21116,I143697,I21133,I143703,I143688,I21150,I21167,I21184,I21201,I143715,I21218,I143685,I21235,I21252,I143694,I143706,I21269,I143691,I21286,I21303,I21320,I21067,I21351,I21368,I143709,I21385,I21402,I143700,I21419,I21436,I21453,I21064,I21484,I21091,I21515,I143718,I21532,I143712,I21549,I21566,I21583,I21082,I21614,I21631,I21070,I21088,I21676,I21693,I21073,I21724,I21079,I21085,I21076,I21813,I21830,I328210,I21847,I328198,I328189,I21864,I21881,I21898,I21915,I21932,I328204,I21949,I21966,I328186,I328195,I21983,I328201,I22000,I22017,I22034,I22065,I22082,I22099,I22116,I22133,I22150,I22167,I22198,I22229,I328192,I22246,I328207,I22263,I22280,I22297,I22328,I22345,I22390,I22407,I22438,I22527,I22544,I116021,I22561,I116027,I116012,I22578,I22595,I22612,I22629,I116039,I22646,I116009,I22663,I22680,I116018,I116030,I22697,I116015,I22714,I22731,I22748,I22495,I22779,I22796,I116033,I22813,I22830,I116024,I22847,I22864,I22881,I22492,I22912,I22519,I22943,I116042,I22960,I116036,I22977,I22994,I23011,I22510,I23042,I23059,I22498,I22516,I23104,I23121,I22501,I23152,I22507,I22513,I22504,I23241,I23258,I48808,I23275,I48829,I23292,I23309,I23326,I23343,I48823,I23360,I48835,I23377,I23394,I48811,I48826,I23411,I48820,I23428,I23445,I23462,I23493,I23510,I48832,I23527,I23544,I48814,I48838,I23561,I23578,I23595,I23626,I23657,I48817,I23674,I48841,I23691,I48844,I23708,I23725,I23756,I23773,I23818,I23835,I23866,I23955,I23972,I179105,I23989,I179102,I179114,I24006,I24023,I24040,I24057,I179123,I24074,I179120,I24091,I24108,I179099,I179096,I24125,I179117,I24142,I24159,I24176,I23923,I24207,I24224,I179108,I24241,I24258,I179126,I24275,I24292,I24309,I23920,I24340,I23947,I24371,I24388,I179111,I24405,I24422,I24439,I23938,I24470,I24487,I23926,I23944,I24532,I24549,I23929,I24580,I23935,I23941,I23932,I24669,I24686,I363309,I24703,I363318,I363315,I24720,I24737,I24754,I24771,I363324,I24788,I363303,I24805,I24822,I363291,I363297,I24839,I363294,I24856,I24873,I24890,I24637,I24921,I24938,I24955,I24972,I363321,I363306,I24989,I25006,I25023,I24634,I25054,I24661,I25085,I363300,I25102,I25119,I363312,I25136,I25153,I24652,I25184,I25201,I24640,I24658,I25246,I25263,I24643,I25294,I24649,I24655,I24646,I25383,I25400,I97202,I25417,I97193,I97190,I25434,I25451,I25468,I25485,I97199,I25502,I25519,I25536,I97214,I25553,I97205,I25570,I25587,I25604,I25351,I25635,I25652,I25669,I25686,I97217,I97196,I25703,I25720,I25737,I25348,I25768,I25375,I25799,I25816,I97211,I25833,I97208,I25850,I25867,I25366,I25898,I25915,I25354,I25372,I25960,I25977,I25357,I26008,I25363,I25369,I25360,I26097,I26114,I165406,I26131,I165418,I165424,I26148,I26165,I26182,I26199,I165397,I26216,I165421,I26233,I26250,I165403,I165394,I26267,I165412,I26284,I26301,I26318,I26065,I26349,I26366,I165415,I26383,I26400,I165400,I26417,I26434,I26451,I26062,I26482,I26089,I26513,I26530,I165427,I26547,I165409,I26564,I26581,I26080,I26612,I26629,I26068,I26086,I26674,I26691,I26071,I26722,I26077,I26083,I26074,I26811,I26828,I434533,I26845,I434524,I434527,I26862,I26879,I26896,I26913,I434521,I26930,I434548,I26947,I26964,I434539,I26981,I434536,I26998,I27015,I27032,I26779,I27063,I27080,I434545,I27097,I27114,I434551,I434542,I27131,I27148,I27165,I26776,I27196,I26803,I27227,I434530,I434554,I27244,I27261,I27278,I27295,I26794,I27326,I27343,I26782,I26800,I27388,I27405,I26785,I27436,I26791,I26797,I26788,I27525,I27542,I27559,I27576,I27593,I27610,I27627,I27644,I27661,I27678,I27695,I27712,I27729,I27746,I27493,I27777,I27794,I27811,I27828,I27845,I27862,I27879,I27490,I27910,I27517,I27941,I27958,I27975,I27992,I28009,I27508,I28040,I28057,I27496,I27514,I28102,I28119,I27499,I28150,I27505,I27511,I27502,I28239,I28256,I65752,I28273,I65743,I65740,I28290,I28307,I28324,I28341,I65749,I28358,I28375,I28392,I65764,I28409,I65755,I28426,I28443,I28460,I28207,I28491,I28508,I28525,I28542,I65767,I65746,I28559,I28576,I28593,I28204,I28624,I28231,I28655,I28672,I65761,I28689,I65758,I28706,I28723,I28222,I28754,I28771,I28210,I28228,I28816,I28833,I28213,I28864,I28219,I28225,I28216,I28953,I28970,I162686,I28987,I162698,I162704,I29004,I29021,I29038,I29055,I162677,I29072,I162701,I29089,I29106,I162683,I162674,I29123,I162692,I29140,I29157,I29174,I28921,I29205,I29222,I162695,I29239,I29256,I162680,I29273,I29290,I29307,I28918,I29338,I28945,I29369,I29386,I162707,I29403,I162689,I29420,I29437,I28936,I29468,I29485,I28924,I28942,I29530,I29547,I28927,I29578,I28933,I28939,I28930,I29667,I29684,I300321,I29701,I300336,I300306,I29718,I29735,I29752,I29769,I300318,I29786,I300309,I29803,I29820,I300330,I300333,I29837,I300312,I29854,I29871,I29888,I29635,I29919,I29936,I300315,I29953,I29970,I29987,I30004,I30021,I29632,I30052,I29659,I30083,I300327,I30100,I300324,I30117,I30134,I30151,I29650,I30182,I30199,I29638,I29656,I30244,I30261,I29641,I30292,I29647,I29653,I29644,I30381,I30398,I339515,I30415,I339503,I339494,I30432,I30449,I30466,I30483,I30500,I339509,I30517,I30534,I339491,I339500,I30551,I339506,I30568,I30585,I30602,I30349,I30633,I30650,I30667,I30684,I30701,I30718,I30735,I30346,I30766,I30373,I30797,I339497,I30814,I339512,I30831,I30848,I30865,I30364,I30896,I30913,I30352,I30370,I30958,I30975,I30355,I31006,I30361,I30367,I30358,I31095,I31112,I245190,I31129,I245184,I245196,I31146,I31163,I31180,I31197,I245202,I31214,I245178,I31231,I31248,I245187,I245175,I31265,I245181,I31282,I31299,I31316,I31063,I31347,I31364,I245205,I31381,I31398,I31415,I31432,I31449,I31060,I31480,I31087,I31511,I245193,I31528,I245199,I31545,I31562,I31579,I31078,I31610,I31627,I31066,I31084,I31672,I31689,I31069,I31720,I31075,I31081,I31072,I31809,I31826,I51936,I31843,I51957,I31860,I31877,I31894,I31911,I51951,I31928,I51963,I31945,I31962,I51939,I51954,I31979,I51948,I31996,I32013,I32030,I31777,I32061,I32078,I51960,I32095,I32112,I51942,I51966,I32129,I32146,I32163,I31774,I32194,I31801,I32225,I51945,I32242,I51969,I32259,I51972,I32276,I32293,I31792,I32324,I32341,I31780,I31798,I32386,I32403,I31783,I32434,I31789,I31795,I31786,I32523,I32540,I241365,I32557,I241359,I241371,I32574,I32591,I32608,I32625,I241377,I32642,I241353,I32659,I32676,I241362,I241350,I32693,I241356,I32710,I32727,I32744,I32491,I32775,I32792,I241380,I32809,I32826,I32843,I32860,I32877,I32488,I32908,I32515,I32939,I241368,I32956,I241374,I32973,I32990,I33007,I32506,I33038,I33055,I32494,I32512,I33100,I33117,I32497,I33148,I32503,I32509,I32500,I33237,I33254,I88396,I33271,I88387,I88384,I33288,I33305,I33322,I33339,I88393,I33356,I33373,I33390,I88408,I33407,I88399,I33424,I33441,I33458,I33205,I33489,I33506,I33523,I33540,I88411,I88390,I33557,I33574,I33591,I33202,I33622,I33229,I33653,I33670,I88405,I33687,I88402,I33704,I33721,I33220,I33752,I33769,I33208,I33226,I33814,I33831,I33211,I33862,I33217,I33223,I33214,I33951,I33968,I359150,I33985,I359138,I359129,I34002,I34019,I34036,I34053,I34070,I359144,I34087,I34104,I359126,I359135,I34121,I359141,I34138,I34155,I34172,I33919,I34203,I34220,I34237,I34254,I34271,I34288,I34305,I33916,I34336,I33943,I34367,I359132,I34384,I359147,I34401,I34418,I34435,I33934,I34466,I34483,I33922,I33940,I34528,I34545,I33925,I34576,I33931,I33937,I33928,I34665,I34682,I107215,I34699,I107221,I107206,I34716,I34733,I34750,I34767,I107233,I34784,I107203,I34801,I34818,I107212,I107224,I34835,I107209,I34852,I34869,I34886,I34633,I34917,I34934,I107227,I34951,I34968,I107218,I34985,I35002,I35019,I34630,I35050,I34657,I35081,I107236,I35098,I107230,I35115,I35132,I35149,I34648,I35180,I35197,I34636,I34654,I35242,I35259,I34639,I35290,I34645,I34651,I34642,I35379,I35396,I252840,I35413,I252834,I252846,I35430,I35447,I35464,I35481,I252852,I35498,I252828,I35515,I35532,I252837,I252825,I35549,I252831,I35566,I35583,I35600,I35347,I35631,I35648,I252855,I35665,I35682,I35699,I35716,I35733,I35344,I35764,I35371,I35795,I252843,I35812,I252849,I35829,I35846,I35863,I35362,I35894,I35911,I35350,I35368,I35956,I35973,I35353,I36004,I35359,I35365,I35356,I36093,I36110,I236775,I36127,I236769,I236781,I36144,I36161,I36178,I36195,I236787,I36212,I236763,I36229,I36246,I236772,I236760,I36263,I236766,I36280,I36297,I36314,I36061,I36345,I36362,I236790,I36379,I36396,I36413,I36430,I36447,I36058,I36478,I36085,I36509,I236778,I36526,I236784,I36543,I36560,I36577,I36076,I36608,I36625,I36064,I36082,I36670,I36687,I36067,I36718,I36073,I36079,I36070,I36807,I36824,I330590,I36841,I330578,I330569,I36858,I36875,I36892,I36909,I36926,I330584,I36943,I36960,I330566,I330575,I36977,I330581,I36994,I37011,I37028,I36775,I37059,I37076,I37093,I37110,I37127,I37144,I37161,I36772,I37192,I36799,I37223,I330572,I37240,I330587,I37257,I37274,I37291,I36790,I37322,I37339,I36778,I36796,I37384,I37401,I36781,I37432,I36787,I36793,I36784,I37521,I37538,I164726,I37555,I164738,I164744,I37572,I37589,I37606,I37623,I164717,I37640,I164741,I37657,I37674,I164723,I164714,I37691,I164732,I37708,I37725,I37742,I37489,I37773,I37790,I164735,I37807,I37824,I164720,I37841,I37858,I37875,I37486,I37906,I37513,I37937,I37954,I164747,I37971,I164729,I37988,I38005,I37504,I38036,I38053,I37492,I37510,I38098,I38115,I37495,I38146,I37501,I37507,I37498,I38235,I38252,I324640,I38269,I324628,I324619,I38286,I38303,I38320,I38337,I38354,I324634,I38371,I38388,I324616,I324625,I38405,I324631,I38422,I38439,I38456,I38203,I38487,I38504,I38521,I38538,I38555,I38572,I38589,I38200,I38620,I38227,I38651,I324622,I38668,I324637,I38685,I38702,I38719,I38218,I38750,I38767,I38206,I38224,I38812,I38829,I38209,I38860,I38215,I38221,I38212,I38949,I38966,I309093,I38983,I309108,I309078,I39000,I39017,I39034,I39051,I309090,I39068,I309081,I39085,I39102,I309102,I309105,I39119,I309084,I39136,I39153,I39170,I38917,I39201,I39218,I309087,I39235,I39252,I39269,I39286,I39303,I38914,I39334,I38941,I39365,I309099,I39382,I309096,I39399,I39416,I39433,I38932,I39464,I39481,I38920,I38938,I39526,I39543,I38923,I39574,I38929,I38935,I38926,I39663,I39680,I373249,I39697,I373231,I373222,I39714,I39731,I39748,I39765,I373243,I39782,I373252,I39799,I39816,I373219,I39833,I373225,I39850,I39867,I39884,I39631,I39915,I39932,I373228,I39949,I39966,I373246,I373237,I39983,I40000,I40017,I39628,I40048,I39655,I40079,I373234,I40096,I40113,I373240,I40130,I40147,I39646,I40178,I40195,I39634,I39652,I40240,I40257,I39637,I40288,I39643,I39649,I39640,I40377,I40394,I199488,I40411,I199494,I199479,I40428,I40445,I40462,I40479,I40496,I199497,I40513,I40530,I199491,I199485,I40547,I199482,I40564,I40581,I40598,I40345,I40629,I40646,I40663,I40680,I199503,I40697,I40714,I40731,I40342,I40762,I40369,I40793,I199500,I40810,I40827,I40844,I40861,I40360,I40892,I40909,I40348,I40366,I40954,I40971,I40351,I41002,I40357,I40363,I40354,I41091,I41108,I211967,I41125,I211943,I211955,I41142,I41159,I41176,I41193,I41210,I211940,I41227,I41244,I211964,I211946,I41261,I211958,I41278,I41295,I41312,I41059,I41343,I41360,I211949,I41377,I41394,I211952,I41411,I41428,I41445,I41056,I41476,I41083,I41507,I41524,I211961,I41541,I41558,I41575,I41074,I41606,I41623,I41062,I41080,I41668,I41685,I41065,I41716,I41071,I41077,I41068,I41814,I41831,I41848,I41874,I41882,I41899,I41770,I41930,I41947,I41964,I41981,I41998,I42015,I41776,I42046,I42063,I42080,I42097,I42114,I41773,I41797,I42159,I42176,I42202,I41779,I41806,I42238,I42255,I42272,I41791,I42303,I41794,I42334,I42351,I41785,I42382,I42399,I41803,I41800,I42444,I42461,I41788,I42492,I42509,I42526,I41782,I42596,I42613,I282660,I282690,I42630,I282675,I42656,I42664,I42681,I282666,I42552,I42712,I42729,I282687,I42746,I282681,I42763,I42780,I282669,I282672,I42797,I42558,I42828,I42845,I282663,I42862,I42879,I42896,I42555,I42579,I42941,I42958,I282684,I42984,I42561,I42588,I43020,I43037,I43054,I42573,I43085,I42576,I43116,I282678,I43133,I42567,I43164,I43181,I42585,I42582,I43226,I43243,I42570,I43274,I43291,I43308,I42564,I43378,I43395,I203721,I203727,I43412,I203724,I43438,I43446,I43463,I203739,I43334,I43494,I203715,I43511,I203718,I43528,I203712,I43545,I43562,I43579,I43340,I43610,I43627,I43644,I43661,I43678,I43337,I43361,I43723,I43740,I203730,I43766,I43343,I43370,I43802,I43819,I43836,I43355,I43867,I43358,I43898,I203733,I203736,I43915,I43349,I43946,I43963,I43367,I43364,I44008,I44025,I43352,I44056,I44073,I44090,I43346,I44160,I44177,I188342,I188339,I44194,I188336,I44220,I44228,I44245,I188333,I44116,I44276,I188327,I44293,I44310,I44327,I44344,I188351,I188330,I44361,I44122,I44392,I44409,I44426,I44443,I44460,I44119,I44143,I44505,I44522,I188345,I44548,I44125,I44152,I44584,I44601,I44618,I44137,I44649,I44140,I44680,I188348,I44697,I44131,I44728,I44745,I44149,I44146,I44790,I44807,I44134,I44838,I44855,I44872,I44128,I44942,I44959,I218681,I218687,I44976,I218684,I45002,I45010,I45027,I218699,I45058,I218675,I45075,I218678,I45092,I218672,I45109,I45126,I45143,I45174,I45191,I45208,I45225,I45242,I45287,I45304,I218690,I45330,I45366,I45383,I45400,I45431,I45462,I218693,I218696,I45479,I45510,I45527,I45572,I45589,I45620,I45637,I45654,I45724,I45741,I45758,I45784,I45792,I45809,I45840,I45857,I45874,I45891,I45908,I45925,I45956,I45973,I45990,I46007,I46024,I46069,I46086,I46112,I46148,I46165,I46182,I46213,I46244,I46261,I46292,I46309,I46354,I46371,I46402,I46419,I46436,I46506,I46523,I91544,I91535,I46540,I91529,I46566,I46574,I46591,I91553,I46462,I46622,I91547,I46639,I91538,I46656,I46673,I46690,I91532,I46707,I46468,I46738,I46755,I91550,I46772,I46789,I46806,I46465,I46489,I46851,I46868,I91541,I46894,I46471,I46498,I46930,I46947,I46964,I46483,I46995,I46486,I47026,I91556,I47043,I46477,I47074,I47091,I46495,I46492,I47136,I47153,I46480,I47184,I47201,I47218,I46474,I47288,I47305,I47322,I47348,I47356,I47373,I47244,I47404,I47421,I47438,I47455,I47472,I47489,I47250,I47520,I47537,I47554,I47571,I47588,I47247,I47271,I47633,I47650,I47676,I47253,I47280,I47712,I47729,I47746,I47265,I47777,I47268,I47808,I47825,I47259,I47856,I47873,I47277,I47274,I47918,I47935,I47262,I47966,I47983,I48000,I47256,I48070,I48087,I306894,I306912,I48104,I306900,I48130,I48138,I48155,I306885,I48026,I48186,I306915,I48203,I306909,I48220,I306891,I48237,I48254,I306888,I48271,I48032,I48302,I48319,I48336,I48353,I48370,I48029,I48053,I48415,I48432,I306903,I48458,I48035,I48062,I48494,I48511,I48528,I48047,I48559,I48050,I48590,I306897,I306906,I48607,I48041,I48638,I48655,I48059,I48056,I48700,I48717,I48044,I48748,I48765,I48782,I48038,I48852,I48869,I356154,I356157,I48886,I356166,I48912,I48920,I48937,I356160,I48968,I356151,I48985,I49002,I49019,I49036,I356175,I49053,I49084,I49101,I356163,I49118,I49135,I49152,I49197,I49214,I356169,I49240,I49276,I49293,I49310,I49341,I49372,I356172,I49389,I49420,I49437,I49482,I49499,I49530,I49547,I49564,I49634,I49651,I277305,I277335,I49668,I277320,I49694,I49702,I49719,I277311,I49590,I49750,I49767,I277332,I49784,I277326,I49801,I49818,I277314,I277317,I49835,I49596,I49866,I49883,I277308,I49900,I49917,I49934,I49593,I49617,I49979,I49996,I277329,I50022,I49599,I49626,I50058,I50075,I50092,I49611,I50123,I49614,I50154,I277323,I50171,I49605,I50202,I50219,I49623,I49620,I50264,I50281,I49608,I50312,I50329,I50346,I49602,I50416,I50433,I368899,I368890,I50450,I368902,I50476,I50484,I50501,I368914,I50372,I50532,I368908,I50549,I368893,I50566,I368911,I50583,I50600,I368917,I368887,I50617,I50378,I50648,I50665,I368884,I50682,I50699,I50716,I50375,I50399,I50761,I50778,I50804,I50381,I50408,I50840,I50857,I50874,I50393,I50905,I50396,I50936,I368905,I368896,I50953,I50387,I50984,I51001,I50405,I50402,I51046,I51063,I50390,I51094,I51111,I51128,I50384,I51198,I51215,I347229,I347232,I51232,I347241,I51258,I51266,I51283,I347235,I51154,I51314,I347226,I51331,I51348,I51365,I51382,I347250,I51399,I51160,I51430,I51447,I347238,I51464,I51481,I51498,I51157,I51181,I51543,I51560,I347244,I51586,I51163,I51190,I51622,I51639,I51656,I51175,I51687,I51178,I51718,I347247,I51735,I51169,I51766,I51783,I51187,I51184,I51828,I51845,I51172,I51876,I51893,I51910,I51166,I51980,I51997,I177649,I177634,I52014,I52040,I52048,I52065,I177640,I52096,I177658,I52113,I177661,I52130,I177646,I52147,I52164,I177664,I52181,I52212,I52229,I177643,I52246,I52263,I52280,I52325,I52342,I177637,I52368,I52404,I52421,I52438,I52469,I52500,I177652,I177655,I52517,I52548,I52565,I52610,I52627,I52658,I52675,I52692,I52762,I52779,I101545,I101566,I52796,I101575,I52822,I52830,I52847,I101569,I52718,I52878,I101560,I52895,I101563,I52912,I101551,I52929,I52946,I101548,I52963,I52724,I52994,I53011,I101542,I53028,I53045,I53062,I52721,I52745,I53107,I53124,I101557,I101554,I53150,I52727,I52754,I53186,I53203,I53220,I52739,I53251,I52742,I53282,I101572,I53299,I52733,I53330,I53347,I52751,I52748,I53392,I53409,I52736,I53440,I53457,I53474,I52730,I53544,I53561,I108464,I108485,I53578,I108494,I53604,I53612,I53629,I108488,I53500,I53660,I108479,I53677,I108482,I53694,I108470,I53711,I53728,I108467,I53745,I53506,I53776,I53793,I108461,I53810,I53827,I53844,I53503,I53527,I53889,I53906,I108476,I108473,I53932,I53509,I53536,I53968,I53985,I54002,I53521,I54033,I53524,I54064,I108491,I54081,I53515,I54112,I54129,I53533,I53530,I54174,I54191,I53518,I54222,I54239,I54256,I53512,I54326,I54343,I70158,I70149,I54360,I70143,I54386,I54394,I54411,I70167,I54282,I54442,I70161,I54459,I70152,I54476,I54493,I54510,I70146,I54527,I54288,I54558,I54575,I70164,I54592,I54609,I54626,I54285,I54309,I54671,I54688,I70155,I54714,I54291,I54318,I54750,I54767,I54784,I54303,I54815,I54306,I54846,I70170,I54863,I54297,I54894,I54911,I54315,I54312,I54956,I54973,I54300,I55004,I55021,I55038,I54294,I55108,I55125,I105319,I105340,I55142,I105349,I55168,I55176,I55193,I105343,I55064,I55224,I105334,I55241,I105337,I55258,I105325,I55275,I55292,I105322,I55309,I55070,I55340,I55357,I105316,I55374,I55391,I55408,I55067,I55091,I55453,I55470,I105331,I105328,I55496,I55073,I55100,I55532,I55549,I55566,I55085,I55597,I55088,I55628,I105346,I55645,I55079,I55676,I55693,I55097,I55094,I55738,I55755,I55082,I55786,I55803,I55820,I55076,I55890,I55907,I314204,I314222,I55924,I314210,I55950,I55958,I55975,I314195,I55846,I56006,I314225,I56023,I314219,I56040,I314201,I56057,I56074,I314198,I56091,I55852,I56122,I56139,I56156,I56173,I56190,I55849,I55873,I56235,I56252,I314213,I56278,I55855,I55882,I56314,I56331,I56348,I55867,I56379,I55870,I56410,I314207,I314216,I56427,I55861,I56458,I56475,I55879,I55876,I56520,I56537,I55864,I56568,I56585,I56602,I55858,I56672,I56689,I68900,I68891,I56706,I68885,I56732,I56740,I56757,I68909,I56628,I56788,I68903,I56805,I68894,I56822,I56839,I56856,I68888,I56873,I56634,I56904,I56921,I68906,I56938,I56955,I56972,I56631,I56655,I57017,I57034,I68897,I57060,I56637,I56664,I57096,I57113,I57130,I56649,I57161,I56652,I57192,I68912,I57209,I56643,I57240,I57257,I56661,I56658,I57302,I57319,I56646,I57350,I57367,I57384,I56640,I57454,I57471,I179842,I179827,I57488,I57514,I57522,I57539,I179833,I57410,I57570,I179851,I57587,I179854,I57604,I179839,I57621,I57638,I179857,I57655,I57416,I57686,I57703,I179836,I57720,I57737,I57754,I57413,I57437,I57799,I57816,I179830,I57842,I57419,I57446,I57878,I57895,I57912,I57431,I57943,I57434,I57974,I179845,I179848,I57991,I57425,I58022,I58039,I57443,I57440,I58084,I58101,I57428,I58132,I58149,I58166,I57422,I58227,I58244,I202270,I58261,I202288,I58278,I58295,I202285,I58312,I58329,I58207,I58360,I202291,I58192,I58216,I58405,I202279,I58422,I202267,I58439,I58456,I58473,I58195,I58504,I58213,I58535,I202273,I58552,I202276,I58569,I58219,I58600,I58617,I58634,I202282,I58651,I58668,I58685,I58702,I58201,I58733,I58204,I58764,I58210,I58795,I58198,I58856,I58873,I396549,I396558,I58890,I396552,I58907,I58924,I396543,I58941,I58958,I58836,I58989,I58821,I58845,I59034,I59051,I396546,I59068,I59085,I59102,I58824,I59133,I58842,I59164,I59181,I396567,I59198,I58848,I59229,I396564,I59246,I396555,I59263,I396561,I59280,I59297,I59314,I59331,I58830,I59362,I58833,I59393,I58839,I59424,I58827,I59485,I59502,I298847,I298862,I59519,I298853,I59536,I59553,I298859,I59570,I59587,I59465,I59618,I298871,I59450,I59474,I59663,I298868,I59680,I298856,I59697,I59714,I59731,I59453,I59762,I59471,I59793,I298844,I59810,I298874,I59827,I59477,I59858,I298850,I59875,I298865,I59892,I59909,I59926,I59943,I59960,I59459,I59991,I59462,I60022,I59468,I60053,I59456,I60114,I60131,I397229,I397238,I60148,I397232,I60165,I60182,I397223,I60199,I60216,I60094,I60247,I60079,I60103,I60292,I60309,I397226,I60326,I60343,I60360,I60082,I60391,I60100,I60422,I60439,I397247,I60456,I60106,I60487,I397244,I60504,I397235,I60521,I397241,I60538,I60555,I60572,I60589,I60088,I60620,I60091,I60651,I60097,I60682,I60085,I60743,I60760,I271188,I60777,I271197,I60794,I60811,I271185,I60828,I60845,I60723,I60876,I271206,I60708,I60732,I60921,I271212,I60938,I271215,I271203,I60955,I60972,I60989,I60711,I61020,I60729,I61051,I271209,I61068,I61085,I60735,I61116,I271191,I271194,I61133,I61150,I271200,I61167,I61184,I61201,I61218,I60717,I61249,I60720,I61280,I60726,I61311,I60714,I61372,I61389,I61406,I61423,I61440,I61457,I61474,I61352,I61505,I61337,I61361,I61550,I61567,I61584,I61601,I61618,I61340,I61649,I61358,I61680,I61697,I61714,I61364,I61745,I61762,I61779,I61796,I61813,I61830,I61847,I61346,I61878,I61349,I61909,I61355,I61940,I61343,I62001,I62018,I379694,I379679,I62035,I379709,I62052,I62069,I379706,I62086,I62103,I61981,I62134,I379700,I61966,I61990,I62179,I379697,I62196,I379682,I62213,I62230,I62247,I61969,I62278,I61987,I62309,I62326,I379685,I62343,I61993,I62374,I379712,I379688,I62391,I62408,I379703,I379691,I62425,I62442,I62459,I62476,I61975,I62507,I61978,I62538,I61984,I62569,I61972,I62630,I62647,I62664,I62681,I62698,I62715,I62732,I62610,I62763,I62595,I62619,I62808,I62825,I62842,I62859,I62876,I62598,I62907,I62616,I62938,I62955,I62972,I62622,I63003,I63020,I63037,I63054,I63071,I63088,I63105,I62604,I63136,I62607,I63167,I62613,I63198,I62601,I63259,I63276,I132378,I132375,I63293,I132363,I63310,I63327,I132390,I63344,I63361,I63239,I63392,I132381,I63224,I63248,I63437,I132366,I63454,I132384,I63471,I63488,I63505,I63227,I63536,I63245,I63567,I132372,I63584,I132369,I63601,I63251,I63632,I132396,I63649,I63666,I132387,I132393,I63683,I63700,I63717,I63734,I63233,I63765,I63236,I63796,I63242,I63827,I63230,I63888,I63905,I244413,I63922,I244422,I63939,I63956,I244410,I63973,I63990,I63868,I64021,I244431,I63853,I63877,I64066,I244437,I64083,I244440,I244428,I64100,I64117,I64134,I63856,I64165,I63874,I64196,I244434,I64213,I64230,I63880,I64261,I244416,I244419,I64278,I64295,I244425,I64312,I64329,I64346,I64363,I63862,I64394,I63865,I64425,I63871,I64456,I63859,I64517,I64534,I285689,I285704,I64551,I285695,I64568,I64585,I285701,I64602,I64619,I64497,I64650,I285713,I64482,I64506,I64695,I285710,I64712,I285698,I64729,I64746,I64763,I64485,I64794,I64503,I64825,I285686,I64842,I285716,I64859,I64509,I64890,I285692,I64907,I285707,I64924,I64941,I64958,I64975,I64992,I64491,I65023,I64494,I65054,I64500,I65085,I64488,I65146,I65163,I398589,I398598,I65180,I398592,I65197,I65214,I398583,I65231,I65248,I65126,I65279,I65111,I65135,I65324,I65341,I398586,I65358,I65375,I65392,I65114,I65423,I65132,I65454,I65471,I398607,I65488,I65138,I65519,I398604,I65536,I398595,I65553,I398601,I65570,I65587,I65604,I65621,I65120,I65652,I65123,I65683,I65129,I65714,I65117,I65775,I65792,I317853,I317868,I65809,I317859,I65826,I65843,I317865,I65860,I65877,I65908,I317877,I65953,I317874,I65970,I317862,I65987,I66004,I66021,I66052,I66083,I317850,I66100,I317880,I66117,I66148,I317856,I66165,I317871,I66182,I66199,I66216,I66233,I66250,I66281,I66312,I66343,I66404,I66421,I234468,I66438,I234477,I66455,I66472,I234465,I66489,I66506,I66384,I66537,I234486,I66369,I66393,I66582,I234492,I66599,I234495,I234483,I66616,I66633,I66650,I66372,I66681,I66390,I66712,I234489,I66729,I66746,I66396,I66777,I234471,I234474,I66794,I66811,I234480,I66828,I66845,I66862,I66879,I66378,I66910,I66381,I66941,I66387,I66972,I66375,I67033,I67050,I125459,I125456,I67067,I125444,I67084,I67101,I125471,I67118,I67135,I67013,I67166,I125462,I66998,I67022,I67211,I125447,I67228,I125465,I67245,I67262,I67279,I67001,I67310,I67019,I67341,I125453,I67358,I125450,I67375,I67025,I67406,I125477,I67423,I67440,I125468,I125474,I67457,I67474,I67491,I67508,I67007,I67539,I67010,I67570,I67016,I67601,I67004,I67662,I67679,I67696,I67713,I67730,I67747,I67764,I67642,I67795,I67627,I67651,I67840,I67857,I67874,I67891,I67908,I67630,I67939,I67648,I67970,I67987,I68004,I67654,I68035,I68052,I68069,I68086,I68103,I68120,I68137,I67636,I68168,I67639,I68199,I67645,I68230,I67633,I68291,I68308,I412926,I412929,I68325,I412947,I68342,I68359,I412920,I68376,I68393,I68271,I68424,I412917,I68256,I68280,I68469,I412914,I68486,I412944,I412923,I68503,I68520,I68537,I68259,I68568,I68277,I68599,I412935,I68616,I412941,I68633,I68283,I68664,I412932,I68681,I68698,I412938,I68715,I68732,I68749,I68766,I68265,I68797,I68268,I68828,I68274,I68859,I68262,I68920,I68937,I404709,I404718,I68954,I404712,I68971,I68988,I404703,I69005,I69022,I69053,I69098,I69115,I404706,I69132,I69149,I69166,I69197,I69228,I69245,I404727,I69262,I69293,I404724,I69310,I404715,I69327,I404721,I69344,I69361,I69378,I69395,I69426,I69457,I69488,I69549,I69566,I328781,I328793,I69583,I328784,I69600,I69617,I328796,I69634,I69651,I69529,I69682,I328805,I69514,I69538,I69727,I69744,I328787,I69761,I69778,I69795,I69517,I69826,I69535,I69857,I69874,I328802,I69891,I69541,I69922,I328799,I69939,I328790,I69956,I69973,I69990,I70007,I70024,I69523,I70055,I69526,I70086,I69532,I70117,I69520,I70178,I70195,I226176,I226155,I70212,I226170,I70229,I70246,I226152,I70263,I70280,I70311,I226167,I70356,I226158,I70373,I226164,I70390,I70407,I70424,I70455,I70486,I226173,I70503,I70520,I70551,I226161,I70568,I70585,I226179,I70602,I70619,I70636,I70653,I70684,I70715,I70746,I70807,I70824,I232173,I70841,I232182,I70858,I70875,I232170,I70892,I70909,I70787,I70940,I232191,I70772,I70796,I70985,I232197,I71002,I232200,I232188,I71019,I71036,I71053,I70775,I71084,I70793,I71115,I232194,I71132,I71149,I70799,I71180,I232176,I232179,I71197,I71214,I232185,I71231,I71248,I71265,I71282,I70781,I71313,I70784,I71344,I70790,I71375,I70778,I71436,I71453,I111621,I111618,I71470,I111606,I71487,I71504,I111633,I71521,I71538,I71416,I71569,I111624,I71401,I71425,I71614,I111609,I71631,I111627,I71648,I71665,I71682,I71404,I71713,I71422,I71744,I111615,I71761,I111612,I71778,I71428,I71809,I111639,I71826,I71843,I111630,I111636,I71860,I71877,I71894,I71911,I71410,I71942,I71413,I71973,I71419,I72004,I71407,I72065,I72082,I151132,I151123,I72099,I151117,I72116,I72133,I151129,I72150,I72167,I72045,I72198,I151141,I72030,I72054,I72243,I151138,I72260,I151147,I151120,I72277,I72294,I72311,I72033,I72342,I72051,I72373,I151126,I72390,I151114,I72407,I72057,I72438,I151144,I151135,I72455,I72472,I72489,I72506,I72523,I72540,I72039,I72571,I72042,I72602,I72048,I72633,I72036,I72694,I72711,I331161,I331173,I72728,I331164,I72745,I72762,I331176,I72779,I72796,I72674,I72827,I331185,I72659,I72683,I72872,I72889,I331167,I72906,I72923,I72940,I72662,I72971,I72680,I73002,I73019,I331182,I73036,I72686,I73067,I331179,I73084,I331170,I73101,I73118,I73135,I73152,I73169,I72668,I73200,I72671,I73231,I72677,I73262,I72665,I73323,I73340,I129862,I129859,I73357,I129847,I73374,I73391,I129874,I73408,I73425,I73303,I73456,I129865,I73288,I73312,I73501,I129850,I73518,I129868,I73535,I73552,I73569,I73291,I73600,I73309,I73631,I129856,I73648,I129853,I73665,I73315,I73696,I129880,I73713,I73730,I129871,I129877,I73747,I73764,I73781,I73798,I73297,I73829,I73300,I73860,I73306,I73891,I73294,I73952,I73969,I127975,I127972,I73986,I127960,I74003,I74020,I127987,I74037,I74054,I73932,I74085,I127978,I73917,I73941,I74130,I127963,I74147,I127981,I74164,I74181,I74198,I73920,I74229,I73938,I74260,I127969,I74277,I127966,I74294,I73944,I74325,I127993,I74342,I74359,I127984,I127990,I74376,I74393,I74410,I74427,I73926,I74458,I73929,I74489,I73935,I74520,I73923,I74581,I74598,I332946,I332958,I74615,I332949,I74632,I74649,I332961,I74666,I74683,I74561,I74714,I332970,I74546,I74570,I74759,I74776,I332952,I74793,I74810,I74827,I74549,I74858,I74567,I74889,I74906,I332967,I74923,I74573,I74954,I332964,I74971,I332955,I74988,I75005,I75022,I75039,I75056,I74555,I75087,I74558,I75118,I74564,I75149,I74552,I75210,I75227,I75244,I75261,I75278,I75295,I75312,I75190,I75343,I75175,I75199,I75388,I75405,I75422,I75439,I75456,I75178,I75487,I75196,I75518,I75535,I75552,I75202,I75583,I75600,I75617,I75634,I75651,I75668,I75685,I75184,I75716,I75187,I75747,I75193,I75778,I75181,I75839,I75856,I150452,I150443,I75873,I150437,I75890,I75907,I150449,I75924,I75941,I75819,I75972,I150461,I75804,I75828,I76017,I150458,I76034,I150467,I150440,I76051,I76068,I76085,I75807,I76116,I75825,I76147,I150446,I76164,I150434,I76181,I75831,I76212,I150464,I150455,I76229,I76246,I76263,I76280,I76297,I76314,I75813,I76345,I75816,I76376,I75822,I76407,I75810,I76468,I76485,I375818,I375803,I76502,I375833,I76519,I76536,I375830,I76553,I76570,I76448,I76601,I375824,I76433,I76457,I76646,I375821,I76663,I375806,I76680,I76697,I76714,I76436,I76745,I76454,I76776,I76793,I375809,I76810,I76460,I76841,I375836,I375812,I76858,I76875,I375827,I375815,I76892,I76909,I76926,I76943,I76442,I76974,I76445,I77005,I76451,I77036,I76439,I77097,I77114,I380340,I380325,I77131,I380355,I77148,I77165,I380352,I77182,I77199,I77077,I77230,I380346,I77062,I77086,I77275,I380343,I77292,I380328,I77309,I77326,I77343,I77065,I77374,I77083,I77405,I77422,I380331,I77439,I77089,I77470,I380358,I380334,I77487,I77504,I380349,I380337,I77521,I77538,I77555,I77572,I77071,I77603,I77074,I77634,I77080,I77665,I77068,I77726,I77743,I195997,I77760,I196015,I77777,I77794,I196012,I77811,I77828,I77706,I77859,I196018,I77691,I77715,I77904,I196006,I77921,I195994,I77938,I77955,I77972,I77694,I78003,I77712,I78034,I196000,I78051,I196003,I78068,I77718,I78099,I78116,I78133,I196009,I78150,I78167,I78184,I78201,I77700,I78232,I77703,I78263,I77709,I78294,I77697,I78355,I78372,I190421,I78389,I190439,I78406,I78423,I190436,I78440,I78457,I78335,I78488,I190442,I78320,I78344,I78533,I190430,I78550,I190418,I78567,I78584,I78601,I78323,I78632,I78341,I78663,I190424,I78680,I190427,I78697,I78347,I78728,I78745,I78762,I190433,I78779,I78796,I78813,I78830,I78329,I78861,I78332,I78892,I78338,I78923,I78326,I78984,I79001,I79018,I79035,I79052,I79069,I79086,I78964,I79117,I78949,I78973,I79162,I79179,I79196,I79213,I79230,I78952,I79261,I78970,I79292,I79309,I79326,I78976,I79357,I79374,I79391,I79408,I79425,I79442,I79459,I78958,I79490,I78961,I79521,I78967,I79552,I78955,I79613,I79630,I413623,I413626,I79647,I413644,I79664,I79681,I413617,I79698,I79715,I79593,I79746,I413614,I79578,I79602,I79791,I413611,I79808,I413641,I413620,I79825,I79842,I79859,I79581,I79890,I79599,I79921,I413632,I79938,I413638,I79955,I79605,I79986,I413629,I80003,I80020,I413635,I80037,I80054,I80071,I80088,I79587,I80119,I79590,I80150,I79596,I80181,I79584,I80242,I80259,I254358,I80276,I254367,I80293,I80310,I254355,I80327,I80344,I80222,I80375,I254376,I80207,I80231,I80420,I254382,I80437,I254385,I254373,I80454,I80471,I80488,I80210,I80519,I80228,I80550,I254379,I80567,I80584,I80234,I80615,I254361,I254364,I80632,I80649,I254370,I80666,I80683,I80700,I80717,I80216,I80748,I80219,I80779,I80225,I80810,I80213,I80871,I80888,I220940,I220919,I80905,I220934,I80922,I80939,I220916,I80956,I80973,I80851,I81004,I220931,I80836,I80860,I81049,I220922,I81066,I220928,I81083,I81100,I81117,I80839,I81148,I80857,I81179,I220937,I81196,I81213,I80863,I81244,I220925,I81261,I81278,I220943,I81295,I81312,I81329,I81346,I80845,I81377,I80848,I81408,I80854,I81439,I80842,I81500,I81517,I81534,I81551,I81568,I81585,I81602,I81480,I81633,I81465,I81489,I81678,I81695,I81712,I81729,I81746,I81468,I81777,I81486,I81808,I81825,I81842,I81492,I81873,I81890,I81907,I81924,I81941,I81958,I81975,I81474,I82006,I81477,I82037,I81483,I82068,I81471,I82129,I82146,I298116,I298131,I82163,I298122,I82180,I82197,I298128,I82214,I82231,I82109,I82262,I298140,I82094,I82118,I82307,I298137,I82324,I298125,I82341,I82358,I82375,I82097,I82406,I82115,I82437,I298113,I82454,I298143,I82471,I82121,I82502,I298119,I82519,I298134,I82536,I82553,I82570,I82587,I82604,I82103,I82635,I82106,I82666,I82112,I82697,I82100,I82758,I82775,I82792,I82809,I82826,I82843,I82860,I82738,I82891,I82723,I82747,I82936,I82953,I82970,I82987,I83004,I82726,I83035,I82744,I83066,I83083,I83100,I82750,I83131,I83148,I83165,I83182,I83199,I83216,I83233,I82732,I83264,I82735,I83295,I82741,I83326,I82729,I83387,I83404,I102186,I102183,I83421,I102171,I83438,I83455,I102198,I83472,I83489,I83367,I83520,I102189,I83352,I83376,I83565,I102174,I83582,I102192,I83599,I83616,I83633,I83355,I83664,I83373,I83695,I102180,I83712,I102177,I83729,I83379,I83760,I102204,I83777,I83794,I102195,I102201,I83811,I83828,I83845,I83862,I83361,I83893,I83364,I83924,I83370,I83955,I83358,I84016,I84033,I147732,I147723,I84050,I147717,I84067,I84084,I147729,I84101,I84118,I83996,I84149,I147741,I83981,I84005,I84194,I147738,I84211,I147747,I147720,I84228,I84245,I84262,I83984,I84293,I84002,I84324,I147726,I84341,I147714,I84358,I84008,I84389,I147744,I147735,I84406,I84423,I84440,I84457,I84474,I84491,I83990,I84522,I83993,I84553,I83999,I84584,I83987,I84645,I84662,I406069,I406078,I84679,I406072,I84696,I84713,I406063,I84730,I84747,I84625,I84778,I84610,I84634,I84823,I84840,I406066,I84857,I84874,I84891,I84613,I84922,I84631,I84953,I84970,I406087,I84987,I84637,I85018,I406084,I85035,I406075,I85052,I406081,I85069,I85086,I85103,I85120,I84619,I85151,I84622,I85182,I84628,I85213,I84616,I85274,I85291,I308350,I308365,I85308,I308356,I85325,I85342,I308362,I85359,I85376,I85254,I85407,I308374,I85239,I85263,I85452,I308371,I85469,I308359,I85486,I85503,I85520,I85242,I85551,I85260,I85582,I308347,I85599,I308377,I85616,I85266,I85647,I308353,I85664,I308368,I85681,I85698,I85715,I85732,I85749,I85248,I85780,I85251,I85811,I85257,I85842,I85245,I85903,I85920,I287151,I287166,I85937,I287157,I85954,I85971,I287163,I85988,I86005,I85883,I86036,I287175,I85868,I85892,I86081,I287172,I86098,I287160,I86115,I86132,I86149,I85871,I86180,I85889,I86211,I287148,I86228,I287178,I86245,I85895,I86276,I287154,I86293,I287169,I86310,I86327,I86344,I86361,I86378,I85877,I86409,I85880,I86440,I85886,I86471,I85874,I86532,I86549,I243648,I86566,I243657,I86583,I86600,I243645,I86617,I86634,I86512,I86665,I243666,I86497,I86521,I86710,I243672,I86727,I243675,I243663,I86744,I86761,I86778,I86500,I86809,I86518,I86840,I243669,I86857,I86874,I86524,I86905,I243651,I243654,I86922,I86939,I243660,I86956,I86973,I86990,I87007,I86506,I87038,I86509,I87069,I86515,I87100,I86503,I87161,I87178,I226924,I226903,I87195,I226918,I87212,I87229,I226900,I87246,I87263,I87141,I87294,I226915,I87126,I87150,I87339,I226906,I87356,I226912,I87373,I87390,I87407,I87129,I87438,I87147,I87469,I226921,I87486,I87503,I87153,I87534,I226909,I87551,I87568,I226927,I87585,I87602,I87619,I87636,I87135,I87667,I87138,I87698,I87144,I87729,I87132,I87790,I87807,I274248,I87824,I274257,I87841,I87858,I274245,I87875,I87892,I87770,I87923,I274266,I87755,I87779,I87968,I274272,I87985,I274275,I274263,I88002,I88019,I88036,I87758,I88067,I87776,I88098,I274269,I88115,I88132,I87782,I88163,I274251,I274254,I88180,I88197,I274260,I88214,I88231,I88248,I88265,I87764,I88296,I87767,I88327,I87773,I88358,I87761,I88419,I88436,I332351,I332363,I88453,I332354,I88470,I88487,I332366,I88504,I88521,I88552,I332375,I88597,I88614,I332357,I88631,I88648,I88665,I88696,I88727,I88744,I332372,I88761,I88792,I332369,I88809,I332360,I88826,I88843,I88860,I88877,I88894,I88925,I88956,I88987,I89048,I89065,I89082,I89099,I89116,I89133,I89150,I89028,I89181,I89013,I89037,I89226,I89243,I89260,I89277,I89294,I89016,I89325,I89034,I89356,I89373,I89390,I89040,I89421,I89438,I89455,I89472,I89489,I89506,I89523,I89022,I89554,I89025,I89585,I89031,I89616,I89019,I89677,I89694,I162012,I162003,I89711,I161997,I89728,I89745,I162009,I89762,I89779,I89657,I89810,I162021,I89642,I89666,I89855,I162018,I89872,I162027,I162000,I89889,I89906,I89923,I89645,I89954,I89663,I89985,I162006,I90002,I161994,I90019,I89669,I90050,I162024,I162015,I90067,I90084,I90101,I90118,I90135,I90152,I89651,I90183,I89654,I90214,I89660,I90245,I89648,I90306,I90323,I90340,I90357,I90374,I90391,I90408,I90286,I90439,I90271,I90295,I90484,I90501,I90518,I90535,I90552,I90274,I90583,I90292,I90614,I90631,I90648,I90298,I90679,I90696,I90713,I90730,I90747,I90764,I90781,I90280,I90812,I90283,I90843,I90289,I90874,I90277,I90935,I90952,I90969,I90986,I91003,I91020,I91037,I90915,I91068,I90900,I90924,I91113,I91130,I91147,I91164,I91181,I90903,I91212,I90921,I91243,I91260,I91277,I90927,I91308,I91325,I91342,I91359,I91376,I91393,I91410,I90909,I91441,I90912,I91472,I90918,I91503,I90906,I91564,I91581,I423381,I423384,I91598,I423402,I91615,I91632,I423375,I91649,I91666,I91697,I423372,I91742,I423369,I91759,I423399,I423378,I91776,I91793,I91810,I91841,I91872,I423390,I91889,I423396,I91906,I91937,I423387,I91954,I91971,I423393,I91988,I92005,I92022,I92039,I92070,I92101,I92132,I92193,I92210,I210468,I210447,I92227,I210462,I92244,I92261,I210444,I92278,I92295,I92173,I92326,I210459,I92158,I92182,I92371,I210450,I92388,I210456,I92405,I92422,I92439,I92161,I92470,I92179,I92501,I210465,I92518,I92535,I92185,I92566,I210453,I92583,I92600,I210471,I92617,I92634,I92651,I92668,I92167,I92699,I92170,I92730,I92176,I92761,I92164,I92822,I92839,I295923,I295938,I92856,I295929,I92873,I92890,I295935,I92907,I92924,I92802,I92955,I295947,I92787,I92811,I93000,I295944,I93017,I295932,I93034,I93051,I93068,I92790,I93099,I92808,I93130,I295920,I93147,I295950,I93164,I92814,I93195,I295926,I93212,I295941,I93229,I93246,I93263,I93280,I93297,I92796,I93328,I92799,I93359,I92805,I93390,I92793,I93451,I93468,I322236,I322248,I93485,I322239,I93502,I93519,I322251,I93536,I93553,I93431,I93584,I322260,I93416,I93440,I93629,I93646,I322242,I93663,I93680,I93697,I93419,I93728,I93437,I93759,I93776,I322257,I93793,I93443,I93824,I322254,I93841,I322245,I93858,I93875,I93892,I93909,I93926,I93425,I93957,I93428,I93988,I93434,I94019,I93422,I94080,I94097,I411532,I411535,I94114,I411553,I94131,I94148,I411526,I94165,I94182,I94060,I94213,I411523,I94045,I94069,I94258,I411520,I94275,I411550,I411529,I94292,I94309,I94326,I94048,I94357,I94066,I94388,I411541,I94405,I411547,I94422,I94072,I94453,I411538,I94470,I94487,I411544,I94504,I94521,I94538,I94555,I94054,I94586,I94057,I94617,I94063,I94648,I94051,I94709,I94726,I167452,I167443,I94743,I167437,I94760,I94777,I167449,I94794,I94811,I94689,I94842,I167461,I94674,I94698,I94887,I167458,I94904,I167467,I167440,I94921,I94938,I94955,I94677,I94986,I94695,I95017,I167446,I95034,I167434,I95051,I94701,I95082,I167464,I167455,I95099,I95116,I95133,I95150,I95167,I95184,I94683,I95215,I94686,I95246,I94692,I95277,I94680,I95338,I95355,I268893,I95372,I268902,I95389,I95406,I268890,I95423,I95440,I95318,I95471,I268911,I95303,I95327,I95516,I268917,I95533,I268920,I268908,I95550,I95567,I95584,I95306,I95615,I95324,I95646,I268914,I95663,I95680,I95330,I95711,I268896,I268899,I95728,I95745,I268905,I95762,I95779,I95796,I95813,I95312,I95844,I95315,I95875,I95321,I95906,I95309,I95967,I95984,I147052,I147043,I96001,I147037,I96018,I96035,I147049,I96052,I96069,I95947,I96100,I147061,I95932,I95956,I96145,I147058,I96162,I147067,I147040,I96179,I96196,I96213,I95935,I96244,I95953,I96275,I147046,I96292,I147034,I96309,I95959,I96340,I147064,I147055,I96357,I96374,I96391,I96408,I96425,I96442,I95941,I96473,I95944,I96504,I95950,I96535,I95938,I96596,I96613,I96630,I96647,I96664,I96681,I96698,I96576,I96729,I96561,I96585,I96774,I96791,I96808,I96825,I96842,I96564,I96873,I96582,I96904,I96921,I96938,I96588,I96969,I96986,I97003,I97020,I97037,I97054,I97071,I96570,I97102,I96573,I97133,I96579,I97164,I96567,I97225,I97242,I137410,I137407,I97259,I137395,I97276,I97293,I137422,I97310,I97327,I97358,I137413,I97403,I137398,I97420,I137416,I97437,I97454,I97471,I97502,I97533,I137404,I97550,I137401,I97567,I97598,I137428,I97615,I97632,I137419,I137425,I97649,I97666,I97683,I97700,I97731,I97762,I97793,I97851,I97868,I223184,I223172,I97885,I97902,I223163,I97919,I223187,I97936,I97953,I223169,I97828,I97984,I97837,I98015,I223166,I98032,I223175,I98049,I98066,I97819,I98097,I98114,I97843,I98145,I223160,I223178,I98162,I223181,I98179,I98196,I98213,I98230,I98247,I98264,I98281,I97825,I97840,I98326,I97822,I98357,I98374,I97834,I98405,I97831,I98463,I98480,I221688,I221676,I98497,I98514,I221667,I98531,I221691,I98548,I98565,I221673,I98440,I98596,I98449,I98627,I221670,I98644,I221679,I98661,I98678,I98431,I98709,I98726,I98455,I98757,I221664,I221682,I98774,I221685,I98791,I98808,I98825,I98842,I98859,I98876,I98893,I98437,I98452,I98938,I98434,I98969,I98986,I98446,I99017,I98443,I99075,I99092,I214956,I214944,I99109,I99126,I214935,I99143,I214959,I99160,I99177,I214941,I99052,I99208,I99061,I99239,I214938,I99256,I214947,I99273,I99290,I99043,I99321,I99338,I99067,I99369,I214932,I214950,I99386,I214953,I99403,I99420,I99437,I99454,I99471,I99488,I99505,I99049,I99064,I99550,I99046,I99581,I99598,I99058,I99629,I99055,I99696,I99713,I182757,I182754,I99730,I182766,I182763,I99747,I99764,I99781,I182751,I182760,I99798,I99815,I99832,I99849,I99866,I99676,I99897,I182769,I99914,I99931,I182775,I99948,I99965,I99688,I99996,I182772,I99655,I100027,I100044,I99661,I99664,I100089,I100106,I100123,I99670,I99658,I100168,I100185,I99673,I99685,I99682,I100244,I99667,I99679,I100325,I100342,I438730,I438703,I100359,I438733,I438712,I100376,I100393,I100410,I438721,I438706,I100427,I438724,I100444,I100461,I100478,I100495,I100305,I100526,I438727,I100543,I438709,I100560,I438715,I100577,I100594,I100317,I100625,I438718,I100284,I100656,I100673,I100290,I100293,I100718,I100735,I438736,I100752,I100299,I100287,I100797,I100814,I100302,I100314,I100311,I100873,I100296,I100308,I100954,I100971,I100988,I101005,I101022,I101039,I101056,I101073,I101090,I101107,I101124,I100934,I101155,I101172,I101189,I101206,I101223,I100946,I101254,I100913,I101285,I101302,I100919,I100922,I101347,I101364,I101381,I100928,I100916,I101426,I101443,I100931,I100943,I100940,I101502,I100925,I100937,I101583,I101600,I101617,I101634,I101651,I101668,I101685,I101702,I101719,I101736,I101753,I101784,I101801,I101818,I101835,I101852,I101883,I101914,I101931,I101976,I101993,I102010,I102055,I102072,I102131,I102212,I102229,I422002,I421975,I102246,I422005,I421984,I102263,I102280,I102297,I421993,I421978,I102314,I421996,I102331,I102348,I102365,I102382,I102413,I421999,I102430,I421981,I102447,I421987,I102464,I102481,I102512,I421990,I102543,I102560,I102605,I102622,I422008,I102639,I102684,I102701,I102760,I102841,I102858,I102875,I102892,I102909,I102926,I102943,I102960,I102977,I102994,I103011,I102821,I103042,I103059,I103076,I103093,I103110,I102833,I103141,I102800,I103172,I103189,I102806,I102809,I103234,I103251,I103268,I102815,I102803,I103313,I103330,I102818,I102830,I102827,I103389,I102812,I102824,I103470,I103487,I103504,I103521,I103538,I103555,I103572,I103589,I103606,I103623,I103640,I103450,I103671,I103688,I103705,I103722,I103739,I103462,I103770,I103429,I103801,I103818,I103435,I103438,I103863,I103880,I103897,I103444,I103432,I103942,I103959,I103447,I103459,I103456,I104018,I103441,I103453,I104099,I104116,I368112,I368097,I104133,I368100,I368118,I104150,I104167,I104184,I368091,I368085,I104201,I368088,I104218,I104235,I104252,I104269,I104079,I104300,I368109,I104317,I368106,I104334,I368115,I104351,I104368,I104091,I104399,I368094,I368103,I104058,I104430,I104447,I104064,I104067,I104492,I104509,I104526,I104073,I104061,I104571,I104588,I104076,I104088,I104085,I104647,I104070,I104082,I104728,I104745,I215686,I215701,I104762,I215695,I215698,I104779,I104796,I104813,I215683,I215692,I104830,I104847,I104864,I104881,I104898,I104708,I104929,I215680,I104946,I104963,I215689,I215707,I104980,I104997,I104720,I105028,I215704,I104687,I105059,I105076,I104693,I104696,I105121,I105138,I105155,I104702,I104690,I105200,I105217,I104705,I104717,I104714,I105276,I104699,I104711,I105357,I105374,I419214,I419187,I105391,I419217,I419196,I105408,I105425,I105442,I419205,I419190,I105459,I419208,I105476,I105493,I105510,I105527,I105558,I419211,I105575,I419193,I105592,I419199,I105609,I105626,I105657,I419202,I105688,I105705,I105750,I105767,I419220,I105784,I105829,I105846,I105905,I105986,I106003,I106020,I106037,I106054,I106071,I106088,I106105,I106122,I106139,I106156,I105966,I106187,I106204,I106221,I106238,I106255,I105978,I106286,I105945,I106317,I106334,I105951,I105954,I106379,I106396,I106413,I105960,I105948,I106458,I106475,I105963,I105975,I105972,I106534,I105957,I105969,I106615,I106632,I225410,I225425,I106649,I225419,I225422,I106666,I106683,I106700,I225407,I225416,I106717,I106734,I106751,I106768,I106785,I106595,I106816,I225404,I106833,I106850,I225413,I225431,I106867,I106884,I106607,I106915,I225428,I106574,I106946,I106963,I106580,I106583,I107008,I107025,I107042,I106589,I106577,I107087,I107104,I106592,I106604,I106601,I107163,I106586,I106598,I107244,I107261,I185545,I185542,I107278,I185554,I185551,I107295,I107312,I107329,I185539,I185548,I107346,I107363,I107380,I107397,I107414,I107445,I185557,I107462,I107479,I185563,I107496,I107513,I107544,I185560,I107575,I107592,I107637,I107654,I107671,I107716,I107733,I107792,I107873,I107890,I280368,I280383,I107907,I280389,I280371,I107924,I107941,I107958,I280374,I280386,I107975,I107992,I108009,I108026,I108043,I107853,I108074,I280377,I280365,I108091,I108108,I280392,I280395,I108125,I108142,I107865,I108173,I280380,I107832,I108204,I108221,I107838,I107841,I108266,I108283,I108300,I107847,I107835,I108345,I108362,I107850,I107862,I107859,I108421,I107844,I107856,I108502,I108519,I108536,I108553,I108570,I108587,I108604,I108621,I108638,I108655,I108672,I108703,I108720,I108737,I108754,I108771,I108802,I108833,I108850,I108895,I108912,I108929,I108974,I108991,I109050,I109131,I109148,I417820,I417793,I109165,I417823,I417802,I109182,I109199,I109216,I417811,I417796,I109233,I417814,I109250,I109267,I109284,I109301,I109111,I109332,I417817,I109349,I417799,I109366,I417805,I109383,I109400,I109123,I109431,I417808,I109090,I109462,I109479,I109096,I109099,I109524,I109541,I417826,I109558,I109105,I109093,I109603,I109620,I109108,I109120,I109117,I109679,I109102,I109114,I109760,I109777,I109794,I109811,I109828,I109845,I109862,I109879,I109896,I109913,I109930,I109740,I109961,I109978,I109995,I110012,I110029,I109752,I110060,I109719,I110091,I110108,I109725,I109728,I110153,I110170,I110187,I109734,I109722,I110232,I110249,I109737,I109749,I109746,I110308,I109731,I109743,I110389,I110406,I397909,I397918,I110423,I397912,I397927,I110440,I110457,I110474,I397924,I110491,I397903,I110508,I110525,I110542,I110559,I110369,I110590,I397906,I110607,I110624,I397915,I110641,I110658,I110381,I110689,I397921,I110348,I110720,I110737,I110354,I110357,I110782,I110799,I110816,I110363,I110351,I110861,I110878,I110366,I110378,I110375,I110937,I110360,I110372,I111018,I111035,I111052,I111069,I111086,I111103,I111120,I111137,I111154,I111171,I111188,I110998,I111219,I111236,I111253,I111270,I111287,I111010,I111318,I110977,I111349,I111366,I110983,I110986,I111411,I111428,I111445,I110992,I110980,I111490,I111507,I110995,I111007,I111004,I111566,I110989,I111001,I111647,I111664,I111681,I111698,I111715,I111732,I111749,I111766,I111783,I111800,I111817,I111848,I111865,I111882,I111899,I111916,I111947,I111978,I111995,I112040,I112057,I112074,I112119,I112136,I112195,I112276,I112293,I112310,I112327,I112344,I112361,I112378,I112395,I112412,I112429,I112446,I112256,I112477,I112494,I112511,I112528,I112545,I112268,I112576,I112235,I112607,I112624,I112241,I112244,I112669,I112686,I112703,I112250,I112238,I112748,I112765,I112253,I112265,I112262,I112824,I112247,I112259,I112905,I112922,I405389,I405398,I112939,I405392,I405407,I112956,I112973,I112990,I405404,I113007,I405383,I113024,I113041,I113058,I113075,I112885,I113106,I405386,I113123,I113140,I405395,I113157,I113174,I112897,I113205,I405401,I112864,I113236,I113253,I112870,I112873,I113298,I113315,I113332,I112879,I112867,I113377,I113394,I112882,I112894,I112891,I113453,I112876,I112888,I113534,I113551,I276543,I276558,I113568,I276564,I276546,I113585,I113602,I113619,I276549,I276561,I113636,I113653,I113670,I113687,I113704,I113514,I113735,I276552,I276540,I113752,I113769,I276567,I276570,I113786,I113803,I113526,I113834,I276555,I113493,I113865,I113882,I113499,I113502,I113927,I113944,I113961,I113508,I113496,I114006,I114023,I113511,I113523,I113520,I114082,I113505,I113517,I114163,I114180,I186939,I186936,I114197,I186948,I186945,I114214,I114231,I114248,I186933,I186942,I114265,I114282,I114299,I114316,I114333,I114143,I114364,I186951,I114381,I114398,I186957,I114415,I114432,I114155,I114463,I186954,I114122,I114494,I114511,I114128,I114131,I114556,I114573,I114590,I114137,I114125,I114635,I114652,I114140,I114152,I114149,I114711,I114134,I114146,I114792,I114809,I114826,I114843,I114860,I114877,I114894,I114911,I114928,I114945,I114962,I114772,I114993,I115010,I115027,I115044,I115061,I114784,I115092,I114751,I115123,I115140,I114757,I114760,I115185,I115202,I115219,I114766,I114754,I115264,I115281,I114769,I114781,I114778,I115340,I114763,I114775,I115421,I115438,I170843,I170861,I115455,I170864,I170858,I115472,I115489,I115506,I170852,I170834,I115523,I170840,I115540,I115557,I115574,I115591,I115622,I170846,I170867,I115639,I170837,I115656,I170849,I115673,I115690,I115721,I170855,I115752,I115769,I115814,I115831,I115848,I115893,I115910,I115969,I116050,I116067,I173563,I173581,I116084,I173584,I173578,I116101,I116118,I116135,I173572,I173554,I116152,I173560,I116169,I116186,I116203,I116220,I116251,I173566,I173587,I116268,I173557,I116285,I173569,I116302,I116319,I116350,I173575,I116381,I116398,I116443,I116460,I116477,I116522,I116539,I116598,I116679,I116696,I279603,I279618,I116713,I279624,I279606,I116730,I116747,I116764,I279609,I279621,I116781,I116798,I116815,I116832,I116849,I116659,I116880,I279612,I279600,I116897,I116914,I279627,I279630,I116931,I116948,I116671,I116979,I279615,I116638,I117010,I117027,I116644,I116647,I117072,I117089,I117106,I116653,I116641,I117151,I117168,I116656,I116668,I116665,I117227,I116650,I116662,I117308,I117325,I117342,I117359,I117376,I117393,I117410,I117427,I117444,I117461,I117478,I117288,I117509,I117526,I117543,I117560,I117577,I117300,I117608,I117267,I117639,I117656,I117273,I117276,I117701,I117718,I117735,I117282,I117270,I117780,I117797,I117285,I117297,I117294,I117856,I117279,I117291,I117937,I117954,I117971,I117988,I118005,I118022,I118039,I118056,I118073,I118090,I118107,I117917,I118138,I118155,I118172,I118189,I118206,I117929,I118237,I117896,I118268,I118285,I117902,I117905,I118330,I118347,I118364,I117911,I117899,I118409,I118426,I117914,I117926,I117923,I118485,I117908,I117920,I118566,I118583,I433851,I433824,I118600,I433854,I433833,I118617,I118634,I118651,I433842,I433827,I118668,I433845,I118685,I118702,I118719,I118736,I118546,I118767,I433848,I118784,I433830,I118801,I433836,I118818,I118835,I118558,I118866,I433839,I118525,I118897,I118914,I118531,I118534,I118959,I118976,I433857,I118993,I118540,I118528,I119038,I119055,I118543,I118555,I118552,I119114,I118537,I118549,I119195,I119212,I119229,I119246,I119263,I119280,I119297,I119314,I119331,I119348,I119365,I119175,I119396,I119413,I119430,I119447,I119464,I119187,I119495,I119154,I119526,I119543,I119160,I119163,I119588,I119605,I119622,I119169,I119157,I119667,I119684,I119172,I119184,I119181,I119743,I119166,I119178,I119824,I119841,I119858,I119875,I119892,I119909,I119926,I119943,I119960,I119977,I119994,I119804,I120025,I120042,I120059,I120076,I120093,I119816,I120124,I119783,I120155,I120172,I119789,I119792,I120217,I120234,I120251,I119798,I119786,I120296,I120313,I119801,I119813,I119810,I120372,I119795,I119807,I120453,I120470,I120487,I120504,I120521,I120538,I120555,I120572,I120589,I120606,I120623,I120654,I120671,I120688,I120705,I120722,I120753,I120784,I120801,I120846,I120863,I120880,I120925,I120942,I121001,I121082,I121099,I249768,I249783,I121116,I249789,I249771,I121133,I121150,I121167,I249774,I249786,I121184,I121201,I121218,I121235,I121252,I121062,I121283,I249777,I249765,I121300,I121317,I249792,I249795,I121334,I121351,I121074,I121382,I249780,I121041,I121413,I121430,I121047,I121050,I121475,I121492,I121509,I121056,I121044,I121554,I121571,I121059,I121071,I121068,I121630,I121053,I121065,I121711,I121728,I235998,I236013,I121745,I236019,I236001,I121762,I121779,I121796,I236004,I236016,I121813,I121830,I121847,I121864,I121881,I121691,I121912,I236007,I235995,I121929,I121946,I236022,I236025,I121963,I121980,I121703,I122011,I236010,I121670,I122042,I122059,I121676,I121679,I122104,I122121,I122138,I121685,I121673,I122183,I122200,I121688,I121700,I121697,I122259,I121682,I121694,I122340,I122357,I231408,I231423,I122374,I231429,I231411,I122391,I122408,I122425,I231414,I231426,I122442,I122459,I122476,I122493,I122510,I122320,I122541,I231417,I231405,I122558,I122575,I231432,I231435,I122592,I122609,I122332,I122640,I231420,I122299,I122671,I122688,I122305,I122308,I122733,I122750,I122767,I122314,I122302,I122812,I122829,I122317,I122329,I122326,I122888,I122311,I122323,I122969,I122986,I189727,I189724,I123003,I189736,I189733,I123020,I123037,I123054,I189721,I189730,I123071,I123088,I123105,I123122,I123139,I122949,I123170,I189739,I123187,I123204,I189745,I123221,I123238,I122961,I123269,I189742,I122928,I123300,I123317,I122934,I122937,I123362,I123379,I123396,I122943,I122931,I123441,I123458,I122946,I122958,I122955,I123517,I122940,I122952,I123598,I123615,I123632,I123649,I123666,I123683,I123700,I123717,I123734,I123751,I123768,I123578,I123799,I123816,I123833,I123850,I123867,I123590,I123898,I123557,I123929,I123946,I123563,I123566,I123991,I124008,I124025,I123572,I123560,I124070,I124087,I123575,I123587,I123584,I124146,I123569,I123581,I124227,I124244,I271953,I271968,I124261,I271974,I271956,I124278,I124295,I124312,I271959,I271971,I124329,I124346,I124363,I124380,I124397,I124207,I124428,I271962,I271950,I124445,I124462,I271977,I271980,I124479,I124496,I124219,I124527,I271965,I124186,I124558,I124575,I124192,I124195,I124620,I124637,I124654,I124201,I124189,I124699,I124716,I124204,I124216,I124213,I124775,I124198,I124210,I124856,I124873,I124890,I124907,I124924,I124941,I124958,I124975,I124992,I125009,I125026,I124836,I125057,I125074,I125091,I125108,I125125,I124848,I125156,I124815,I125187,I125204,I124821,I124824,I125249,I125266,I125283,I124830,I124818,I125328,I125345,I124833,I124845,I124842,I125404,I124827,I124839,I125485,I125502,I164043,I164061,I125519,I164064,I164058,I125536,I125553,I125570,I164052,I164034,I125587,I164040,I125604,I125621,I125638,I125655,I125686,I164046,I164067,I125703,I164037,I125720,I164049,I125737,I125754,I125785,I164055,I125816,I125833,I125878,I125895,I125912,I125957,I125974,I126033,I126114,I126131,I168803,I168821,I126148,I168824,I168818,I126165,I126182,I126199,I168812,I168794,I126216,I168800,I126233,I126250,I126267,I126284,I126094,I126315,I168806,I168827,I126332,I168797,I126349,I168809,I126366,I126383,I126106,I126414,I168815,I126073,I126445,I126462,I126079,I126082,I126507,I126524,I126541,I126088,I126076,I126586,I126603,I126091,I126103,I126100,I126662,I126085,I126097,I126743,I126760,I126777,I126794,I126811,I126828,I126845,I126862,I126879,I126896,I126913,I126723,I126944,I126961,I126978,I126995,I127012,I126735,I127043,I126702,I127074,I127091,I126708,I126711,I127136,I127153,I127170,I126717,I126705,I127215,I127232,I126720,I126732,I126729,I127291,I126714,I126726,I127372,I127389,I159963,I159981,I127406,I159984,I159978,I127423,I127440,I127457,I159972,I159954,I127474,I159960,I127491,I127508,I127525,I127542,I127573,I159966,I159987,I127590,I159957,I127607,I159969,I127624,I127641,I127672,I159975,I127703,I127720,I127765,I127782,I127799,I127844,I127861,I127920,I128001,I128018,I232938,I232953,I128035,I232959,I232941,I128052,I128069,I128086,I232944,I232956,I128103,I128120,I128137,I128154,I128171,I128202,I232947,I232935,I128219,I128236,I232962,I232965,I128253,I128270,I128301,I232950,I128332,I128349,I128394,I128411,I128428,I128473,I128490,I128549,I128630,I128647,I128664,I128681,I128698,I128715,I128732,I128749,I128766,I128783,I128800,I128610,I128831,I128848,I128865,I128882,I128899,I128622,I128930,I128589,I128961,I128978,I128595,I128598,I129023,I129040,I129057,I128604,I128592,I129102,I129119,I128607,I128619,I128616,I129178,I128601,I128613,I129259,I129276,I129293,I129310,I129327,I129344,I129361,I129378,I129395,I129412,I129429,I129239,I129460,I129477,I129494,I129511,I129528,I129251,I129559,I129218,I129590,I129607,I129224,I129227,I129652,I129669,I129686,I129233,I129221,I129731,I129748,I129236,I129248,I129245,I129807,I129230,I129242,I129888,I129905,I129922,I129939,I129956,I129973,I129990,I130007,I130024,I130041,I130058,I130089,I130106,I130123,I130140,I130157,I130188,I130219,I130236,I130281,I130298,I130315,I130360,I130377,I130436,I130517,I130534,I247473,I247488,I130551,I247494,I247476,I130568,I130585,I130602,I247479,I247491,I130619,I130636,I130653,I130670,I130687,I130497,I130718,I247482,I247470,I130735,I130752,I247497,I247500,I130769,I130786,I130509,I130817,I247485,I130476,I130848,I130865,I130482,I130485,I130910,I130927,I130944,I130491,I130479,I130989,I131006,I130494,I130506,I130503,I131065,I130488,I130500,I131146,I131163,I410850,I410823,I131180,I410853,I410832,I131197,I131214,I131231,I410841,I410826,I131248,I410844,I131265,I131282,I131299,I131316,I131126,I131347,I410847,I131364,I410829,I131381,I410835,I131398,I131415,I131138,I131446,I410838,I131105,I131477,I131494,I131111,I131114,I131539,I131556,I410856,I131573,I131120,I131108,I131618,I131635,I131123,I131135,I131132,I131694,I131117,I131129,I131775,I131792,I131809,I131826,I131843,I131860,I131877,I131894,I131911,I131928,I131945,I131755,I131976,I131993,I132010,I132027,I132044,I131767,I132075,I131734,I132106,I132123,I131740,I131743,I132168,I132185,I132202,I131749,I131737,I132247,I132264,I131752,I131764,I131761,I132323,I131746,I131758,I132404,I132421,I132438,I132455,I132472,I132489,I132506,I132523,I132540,I132557,I132574,I132605,I132622,I132639,I132656,I132673,I132704,I132735,I132752,I132797,I132814,I132831,I132876,I132893,I132952,I133033,I133050,I157243,I157261,I133067,I157264,I157258,I133084,I133101,I133118,I157252,I157234,I133135,I157240,I133152,I133169,I133186,I133203,I133013,I133234,I157246,I157267,I133251,I157237,I133268,I157249,I133285,I133302,I133025,I133333,I157255,I132992,I133364,I133381,I132998,I133001,I133426,I133443,I133460,I133007,I132995,I133505,I133522,I133010,I133022,I133019,I133581,I133004,I133016,I133662,I133679,I246708,I246723,I133696,I246729,I246711,I133713,I133730,I133747,I246714,I246726,I133764,I133781,I133798,I133815,I133832,I133642,I133863,I246717,I246705,I133880,I133897,I246732,I246735,I133914,I133931,I133654,I133962,I246720,I133621,I133993,I134010,I133627,I133630,I134055,I134072,I134089,I133636,I133624,I134134,I134151,I133639,I133651,I133648,I134210,I133633,I133645,I134291,I134308,I409469,I409478,I134325,I409472,I409487,I134342,I134359,I134376,I409484,I134393,I409463,I134410,I134427,I134444,I134461,I134271,I134492,I409466,I134509,I134526,I409475,I134543,I134560,I134283,I134591,I409481,I134250,I134622,I134639,I134256,I134259,I134684,I134701,I134718,I134265,I134253,I134763,I134780,I134268,I134280,I134277,I134839,I134262,I134274,I134920,I134937,I283428,I283443,I134954,I283449,I283431,I134971,I134988,I135005,I283434,I283446,I135022,I135039,I135056,I135073,I135090,I134900,I135121,I283437,I283425,I135138,I135155,I283452,I283455,I135172,I135189,I134912,I135220,I283440,I134879,I135251,I135268,I134885,I134888,I135313,I135330,I135347,I134894,I134882,I135392,I135409,I134897,I134909,I134906,I135468,I134891,I134903,I135549,I135566,I135583,I135600,I135617,I135634,I135651,I135668,I135685,I135702,I135719,I135529,I135750,I135767,I135784,I135801,I135818,I135541,I135849,I135508,I135880,I135897,I135514,I135517,I135942,I135959,I135976,I135523,I135511,I136021,I136038,I135526,I135538,I135535,I136097,I135520,I135532,I136178,I136195,I237528,I237543,I136212,I237549,I237531,I136229,I136246,I136263,I237534,I237546,I136280,I136297,I136314,I136331,I136348,I136158,I136379,I237537,I237525,I136396,I136413,I237552,I237555,I136430,I136447,I136170,I136478,I237540,I136137,I136509,I136526,I136143,I136146,I136571,I136588,I136605,I136152,I136140,I136650,I136667,I136155,I136167,I136164,I136726,I136149,I136161,I136807,I136824,I136841,I136858,I136875,I136892,I136909,I136926,I136943,I136960,I136977,I136787,I137008,I137025,I137042,I137059,I137076,I136799,I137107,I136766,I137138,I137155,I136772,I136775,I137200,I137217,I137234,I136781,I136769,I137279,I137296,I136784,I136796,I136793,I137355,I136778,I136790,I137436,I137453,I137470,I137487,I137504,I137521,I137538,I137555,I137572,I137589,I137606,I137637,I137654,I137671,I137688,I137705,I137736,I137767,I137784,I137829,I137846,I137863,I137908,I137925,I137984,I138065,I138082,I211198,I211213,I138099,I211207,I211210,I138116,I138133,I138150,I211195,I211204,I138167,I138184,I138201,I138218,I138235,I138045,I138266,I211192,I138283,I138300,I211201,I211219,I138317,I138334,I138057,I138365,I211216,I138024,I138396,I138413,I138030,I138033,I138458,I138475,I138492,I138039,I138027,I138537,I138554,I138042,I138054,I138051,I138613,I138036,I138048,I138694,I138711,I138728,I138745,I138762,I138779,I138796,I138813,I138830,I138847,I138864,I138674,I138895,I138912,I138929,I138946,I138963,I138686,I138994,I138653,I139025,I139042,I138659,I138662,I139087,I139104,I139121,I138668,I138656,I139166,I139183,I138671,I138683,I138680,I139242,I138665,I138677,I139323,I139340,I259713,I259728,I139357,I259734,I259716,I139374,I139391,I139408,I259719,I259731,I139425,I139442,I139459,I139476,I139493,I139303,I139524,I259722,I259710,I139541,I139558,I259737,I259740,I139575,I139592,I139315,I139623,I259725,I139282,I139654,I139671,I139288,I139291,I139716,I139733,I139750,I139297,I139285,I139795,I139812,I139300,I139312,I139309,I139871,I139294,I139306,I139952,I139969,I242118,I242133,I139986,I242139,I242121,I140003,I140020,I140037,I242124,I242136,I140054,I140071,I140088,I140105,I140122,I139932,I140153,I242127,I242115,I140170,I140187,I242142,I242145,I140204,I140221,I139944,I140252,I242130,I139911,I140283,I140300,I139917,I139920,I140345,I140362,I140379,I139926,I139914,I140424,I140441,I139929,I139941,I139938,I140500,I139923,I139935,I140581,I140598,I140615,I140632,I140649,I140666,I140683,I140700,I140717,I140734,I140751,I140561,I140782,I140799,I140816,I140833,I140850,I140573,I140881,I140540,I140912,I140929,I140546,I140549,I140974,I140991,I141008,I140555,I140543,I141053,I141070,I140558,I140570,I140567,I141129,I140552,I140564,I141210,I141227,I141244,I141261,I141278,I141295,I141312,I141329,I141346,I141363,I141380,I141190,I141411,I141428,I141445,I141462,I141479,I141202,I141510,I141169,I141541,I141558,I141175,I141178,I141603,I141620,I141637,I141184,I141172,I141682,I141699,I141187,I141199,I141196,I141758,I141181,I141193,I141839,I141856,I406749,I406758,I141873,I406752,I406767,I141890,I141907,I141924,I406764,I141941,I406743,I141958,I141975,I141992,I142009,I141819,I142040,I406746,I142057,I142074,I406755,I142091,I142108,I141831,I142139,I406761,I141798,I142170,I142187,I141804,I141807,I142232,I142249,I142266,I141813,I141801,I142311,I142328,I141816,I141828,I141825,I142387,I141810,I141822,I142468,I142485,I428275,I428248,I142502,I428278,I428257,I142519,I142536,I142553,I428266,I428251,I142570,I428269,I142587,I142604,I142621,I142638,I142448,I142669,I428272,I142686,I428254,I142703,I428260,I142720,I142737,I142460,I142768,I428263,I142427,I142799,I142816,I142433,I142436,I142861,I142878,I428281,I142895,I142442,I142430,I142940,I142957,I142445,I142457,I142454,I143016,I142439,I142451,I143097,I143114,I143131,I143148,I143165,I143182,I143199,I143216,I143233,I143250,I143267,I143077,I143298,I143315,I143332,I143349,I143366,I143089,I143397,I143056,I143428,I143445,I143062,I143065,I143490,I143507,I143524,I143071,I143059,I143569,I143586,I143074,I143086,I143083,I143645,I143068,I143080,I143726,I143743,I385520,I385496,I143760,I385526,I385508,I143777,I143794,I143811,I385514,I385523,I143828,I385499,I143845,I143862,I143879,I143896,I143927,I385505,I143944,I143961,I385493,I143978,I143995,I144026,I385511,I385517,I144057,I144074,I144119,I144136,I385502,I144153,I144198,I144215,I144274,I144355,I144372,I323426,I323435,I144389,I144406,I323441,I144423,I323447,I144440,I144457,I323429,I144314,I144488,I144344,I144519,I323438,I144536,I323444,I144553,I144570,I144587,I144320,I144332,I144632,I144335,I144663,I144680,I323432,I144697,I144714,I144731,I144748,I144338,I144341,I144793,I323450,I144810,I144827,I144844,I144861,I144326,I144892,I144329,I144923,I144317,I144954,I144347,I144323,I145035,I145052,I235248,I235251,I145069,I145086,I235233,I145103,I235260,I145120,I145137,I235245,I144994,I145168,I145024,I145199,I235257,I145216,I235236,I235239,I145233,I145250,I145267,I145000,I145012,I145312,I145015,I145343,I145360,I145377,I235242,I145394,I145411,I145428,I145018,I145021,I145473,I235230,I145490,I235254,I145507,I145524,I145541,I145006,I145572,I145009,I145603,I144997,I145634,I145027,I145003,I145715,I145732,I424066,I424084,I145749,I145766,I424099,I145783,I424069,I145800,I145817,I424072,I145848,I145879,I424093,I145896,I424081,I424096,I145913,I145930,I145947,I145992,I146023,I146040,I424087,I146057,I146074,I146091,I146108,I146153,I146170,I424075,I146187,I424090,I424078,I146204,I146221,I146252,I146283,I146314,I146395,I146412,I146429,I146446,I146463,I146480,I146497,I146354,I146528,I146384,I146559,I146576,I146593,I146610,I146627,I146360,I146372,I146672,I146375,I146703,I146720,I146737,I146754,I146771,I146788,I146378,I146381,I146833,I146850,I146867,I146884,I146901,I146366,I146932,I146369,I146963,I146357,I146994,I146387,I146363,I147075,I147092,I147109,I147126,I147143,I147160,I147177,I147208,I147239,I147256,I147273,I147290,I147307,I147352,I147383,I147400,I147417,I147434,I147451,I147468,I147513,I147530,I147547,I147564,I147581,I147612,I147643,I147674,I147755,I147772,I441491,I441509,I147789,I147806,I441524,I147823,I441494,I147840,I147857,I441497,I147888,I147919,I441518,I147936,I441506,I441521,I147953,I147970,I147987,I148032,I148063,I148080,I441512,I148097,I148114,I148131,I148148,I148193,I148210,I441500,I148227,I441515,I441503,I148244,I148261,I148292,I148323,I148354,I148435,I148452,I229165,I229144,I148469,I148486,I229147,I148503,I229171,I148520,I148537,I229162,I148394,I148568,I148424,I148599,I229159,I148616,I229153,I148633,I148650,I148667,I148400,I148412,I148712,I148415,I148743,I148760,I229156,I148777,I148794,I148811,I148828,I148418,I148421,I148873,I229150,I148890,I148907,I229168,I148924,I148941,I148406,I148972,I148409,I149003,I148397,I149034,I148427,I148403,I149115,I149132,I278853,I278856,I149149,I149166,I278838,I149183,I278865,I149200,I149217,I278850,I149248,I149279,I278862,I149296,I278841,I278844,I149313,I149330,I149347,I149392,I149423,I149440,I149457,I278847,I149474,I149491,I149508,I149553,I278835,I149570,I278859,I149587,I149604,I149621,I149652,I149683,I149714,I149795,I149812,I239838,I239841,I149829,I149846,I239823,I149863,I239850,I149880,I149897,I239835,I149754,I149928,I149784,I149959,I239847,I149976,I239826,I239829,I149993,I150010,I150027,I149760,I149772,I150072,I149775,I150103,I150120,I150137,I239832,I150154,I150171,I150188,I149778,I149781,I150233,I239820,I150250,I239844,I150267,I150284,I150301,I149766,I150332,I149769,I150363,I149757,I150394,I149787,I149763,I150475,I150492,I268143,I268146,I150509,I150526,I268128,I150543,I268155,I150560,I150577,I268140,I150608,I150639,I268152,I150656,I268131,I268134,I150673,I150690,I150707,I150752,I150783,I150800,I150817,I268137,I150834,I150851,I150868,I150913,I268125,I150930,I268149,I150947,I150964,I150981,I151012,I151043,I151074,I151155,I151172,I353176,I353185,I151189,I151206,I353191,I151223,I353197,I151240,I151257,I353179,I151288,I151319,I353188,I151336,I353194,I151353,I151370,I151387,I151432,I151463,I151480,I353182,I151497,I151514,I151531,I151548,I151593,I353200,I151610,I151627,I151644,I151661,I151692,I151723,I151754,I151835,I151852,I421278,I421296,I151869,I151886,I421311,I151903,I421281,I151920,I151937,I421284,I151794,I151968,I151824,I151999,I421305,I152016,I421293,I421308,I152033,I152050,I152067,I151800,I151812,I152112,I151815,I152143,I152160,I421299,I152177,I152194,I152211,I152228,I151818,I151821,I152273,I152290,I421287,I152307,I421302,I421290,I152324,I152341,I151806,I152372,I151809,I152403,I151797,I152434,I151827,I151803,I152515,I152532,I362696,I362705,I152549,I152566,I362711,I152583,I362717,I152600,I152617,I362699,I152474,I152648,I152504,I152679,I362708,I152696,I362714,I152713,I152730,I152747,I152480,I152492,I152792,I152495,I152823,I152840,I362702,I152857,I152874,I152891,I152908,I152498,I152501,I152953,I362720,I152970,I152987,I153004,I153021,I152486,I153052,I152489,I153083,I152477,I153114,I152507,I152483,I153195,I153212,I153229,I153246,I153263,I153280,I153297,I153154,I153328,I153184,I153359,I153376,I153393,I153410,I153427,I153160,I153172,I153472,I153175,I153503,I153520,I153537,I153554,I153571,I153588,I153178,I153181,I153633,I153650,I153667,I153684,I153701,I153166,I153732,I153169,I153763,I153157,I153794,I153187,I153163,I153875,I153892,I153909,I153926,I153943,I153960,I153977,I153834,I154008,I153864,I154039,I154056,I154073,I154090,I154107,I153840,I153852,I154152,I153855,I154183,I154200,I154217,I154234,I154251,I154268,I153858,I153861,I154313,I154330,I154347,I154364,I154381,I153846,I154412,I153849,I154443,I153837,I154474,I153867,I153843,I154555,I154572,I154589,I154606,I154623,I154640,I154657,I154688,I154719,I154736,I154753,I154770,I154787,I154832,I154863,I154880,I154897,I154914,I154931,I154948,I154993,I155010,I155027,I155044,I155061,I155092,I155123,I155154,I155235,I155252,I395192,I155269,I155286,I395204,I155303,I395183,I155320,I155337,I395186,I155194,I155368,I155224,I155399,I395201,I155416,I395195,I395189,I155433,I155450,I155467,I155200,I155212,I155512,I155215,I155543,I155560,I155577,I155594,I155611,I155628,I155218,I155221,I155673,I395198,I155690,I155707,I395207,I155724,I155741,I155206,I155772,I155209,I155803,I155197,I155834,I155227,I155203,I155915,I155932,I407432,I155949,I155966,I407444,I155983,I407423,I156000,I156017,I407426,I155874,I156048,I155904,I156079,I407441,I156096,I407435,I407429,I156113,I156130,I156147,I155880,I155892,I156192,I155895,I156223,I156240,I156257,I156274,I156291,I156308,I155898,I155901,I156353,I407438,I156370,I156387,I407447,I156404,I156421,I155886,I156452,I155889,I156483,I155877,I156514,I155907,I155883,I156595,I156612,I156629,I156646,I156663,I156680,I156697,I156554,I156728,I156584,I156759,I156776,I156793,I156810,I156827,I156560,I156572,I156872,I156575,I156903,I156920,I156937,I156954,I156971,I156988,I156578,I156581,I157033,I157050,I157067,I157084,I157101,I156566,I157132,I156569,I157163,I156557,I157194,I156587,I156563,I157275,I157292,I206725,I206704,I157309,I157326,I206707,I157343,I206731,I157360,I157377,I206722,I157408,I157439,I206719,I157456,I206713,I157473,I157490,I157507,I157552,I157583,I157600,I206716,I157617,I157634,I157651,I157668,I157713,I206710,I157730,I157747,I206728,I157764,I157781,I157812,I157843,I157874,I157955,I157972,I358531,I358540,I157989,I158006,I358546,I158023,I358552,I158040,I158057,I358534,I157914,I158088,I157944,I158119,I358543,I158136,I358549,I158153,I158170,I158187,I157920,I157932,I158232,I157935,I158263,I158280,I358537,I158297,I158314,I158331,I158348,I157938,I157941,I158393,I358555,I158410,I158427,I158444,I158461,I157926,I158492,I157929,I158523,I157917,I158554,I157947,I157923,I158635,I158652,I351391,I351400,I158669,I158686,I351406,I158703,I351412,I158720,I158737,I351394,I158768,I158799,I351403,I158816,I351409,I158833,I158850,I158867,I158912,I158943,I158960,I351397,I158977,I158994,I159011,I159028,I159073,I351415,I159090,I159107,I159124,I159141,I159172,I159203,I159234,I159315,I159332,I214205,I214184,I159349,I159366,I214187,I159383,I214211,I159400,I159417,I214202,I159274,I159448,I159304,I159479,I214199,I159496,I214193,I159513,I159530,I159547,I159280,I159292,I159592,I159295,I159623,I159640,I214196,I159657,I159674,I159691,I159708,I159298,I159301,I159753,I214190,I159770,I159787,I214208,I159804,I159821,I159286,I159852,I159289,I159883,I159277,I159914,I159307,I159283,I159995,I160012,I160029,I160046,I160063,I160080,I160097,I160128,I160159,I160176,I160193,I160210,I160227,I160272,I160303,I160320,I160337,I160354,I160371,I160388,I160433,I160450,I160467,I160484,I160501,I160532,I160563,I160594,I160675,I160692,I160709,I160726,I160743,I160760,I160777,I160634,I160808,I160664,I160839,I160856,I160873,I160890,I160907,I160640,I160652,I160952,I160655,I160983,I161000,I161017,I161034,I161051,I161068,I160658,I160661,I161113,I161130,I161147,I161164,I161181,I160646,I161212,I160649,I161243,I160637,I161274,I160667,I160643,I161355,I161372,I304722,I304698,I161389,I161406,I161423,I304716,I161440,I161457,I304704,I161314,I161488,I161344,I161519,I304707,I161536,I304701,I304692,I161553,I161570,I161587,I161320,I161332,I161632,I161335,I161663,I161680,I304719,I161697,I304713,I161714,I161731,I161748,I161338,I161341,I161793,I304710,I161810,I161827,I304695,I161844,I161861,I161326,I161892,I161329,I161923,I161317,I161954,I161347,I161323,I162035,I162052,I415005,I415023,I162069,I162086,I415038,I162103,I415008,I162120,I162137,I415011,I162168,I162199,I415032,I162216,I415020,I415035,I162233,I162250,I162267,I162312,I162343,I162360,I415026,I162377,I162394,I162411,I162428,I162473,I162490,I415014,I162507,I415029,I415017,I162524,I162541,I162572,I162603,I162634,I162715,I162732,I217197,I217176,I162749,I162766,I217179,I162783,I217203,I162800,I162817,I217194,I162848,I162879,I217191,I162896,I217185,I162913,I162930,I162947,I162992,I163023,I163040,I217188,I163057,I163074,I163091,I163108,I163153,I217182,I163170,I163187,I217200,I163204,I163221,I163252,I163283,I163314,I163395,I163412,I250548,I250551,I163429,I163446,I250533,I163463,I250560,I163480,I163497,I250545,I163354,I163528,I163384,I163559,I250557,I163576,I250536,I250539,I163593,I163610,I163627,I163360,I163372,I163672,I163375,I163703,I163720,I163737,I250542,I163754,I163771,I163788,I163378,I163381,I163833,I250530,I163850,I250554,I163867,I163884,I163901,I163366,I163932,I163369,I163963,I163357,I163994,I163387,I163363,I164075,I164092,I360316,I360325,I164109,I164126,I360331,I164143,I360337,I164160,I164177,I360319,I164208,I164239,I360328,I164256,I360334,I164273,I164290,I164307,I164352,I164383,I164400,I360322,I164417,I164434,I164451,I164468,I164513,I360340,I164530,I164547,I164564,I164581,I164612,I164643,I164674,I164755,I164772,I164789,I164806,I164823,I164840,I164857,I164888,I164919,I164936,I164953,I164970,I164987,I165032,I165063,I165080,I165097,I165114,I165131,I165148,I165193,I165210,I165227,I165244,I165261,I165292,I165323,I165354,I165435,I165452,I165469,I165486,I165503,I165520,I165537,I165568,I165599,I165616,I165633,I165650,I165667,I165712,I165743,I165760,I165777,I165794,I165811,I165828,I165873,I165890,I165907,I165924,I165941,I165972,I166003,I166034,I166115,I166132,I416399,I416417,I166149,I166166,I416432,I166183,I416402,I166200,I166217,I416405,I166074,I166248,I166104,I166279,I416426,I166296,I416414,I416429,I166313,I166330,I166347,I166080,I166092,I166392,I166095,I166423,I166440,I416420,I166457,I166474,I166491,I166508,I166098,I166101,I166553,I166570,I416408,I166587,I416423,I416411,I166604,I166621,I166086,I166652,I166089,I166683,I166077,I166714,I166107,I166083,I166795,I166812,I166829,I166846,I166863,I166880,I166897,I166754,I166928,I166784,I166959,I166976,I166993,I167010,I167027,I166760,I166772,I167072,I166775,I167103,I167120,I167137,I167154,I167171,I167188,I166778,I166781,I167233,I167250,I167267,I167284,I167301,I166766,I167332,I166769,I167363,I166757,I167394,I166787,I166763,I167475,I167492,I208969,I208948,I167509,I167526,I208951,I167543,I208975,I167560,I167577,I208966,I167608,I167639,I208963,I167656,I208957,I167673,I167690,I167707,I167752,I167783,I167800,I208960,I167817,I167834,I167851,I167868,I167913,I208954,I167930,I167947,I208972,I167964,I167981,I168012,I168043,I168074,I168155,I168172,I357341,I357350,I168189,I168206,I357356,I168223,I357362,I168240,I168257,I357344,I168114,I168288,I168144,I168319,I357353,I168336,I357359,I168353,I168370,I168387,I168120,I168132,I168432,I168135,I168463,I168480,I357347,I168497,I168514,I168531,I168548,I168138,I168141,I168593,I357365,I168610,I168627,I168644,I168661,I168126,I168692,I168129,I168723,I168117,I168754,I168147,I168123,I168835,I168852,I388723,I388750,I168869,I168886,I388726,I168903,I388741,I168920,I168937,I388747,I168968,I168999,I388738,I169016,I388735,I388729,I169033,I169050,I169067,I169112,I169143,I169160,I169177,I388753,I169194,I169211,I169228,I169273,I169290,I388744,I169307,I388756,I388732,I169324,I169341,I169372,I169403,I169434,I169515,I169532,I366505,I366499,I169549,I169566,I366511,I169583,I366514,I169600,I169617,I366517,I169474,I169648,I169504,I169679,I366502,I169696,I366493,I366490,I169713,I169730,I169747,I169480,I169492,I169792,I169495,I169823,I169840,I366487,I169857,I366496,I169874,I169891,I169908,I169498,I169501,I169953,I366520,I169970,I169987,I366508,I170004,I170021,I169486,I170052,I169489,I170083,I169477,I170114,I169507,I169483,I170195,I170212,I445673,I445691,I170229,I170246,I445706,I170263,I445676,I170280,I170297,I445679,I170154,I170328,I170184,I170359,I445700,I170376,I445688,I445703,I170393,I170410,I170427,I170160,I170172,I170472,I170175,I170503,I170520,I445694,I170537,I170554,I170571,I170588,I170178,I170181,I170633,I170650,I445682,I170667,I445697,I445685,I170684,I170701,I170166,I170732,I170169,I170763,I170157,I170794,I170187,I170163,I170875,I170892,I260493,I260496,I170909,I170926,I260478,I170943,I260505,I170960,I170977,I260490,I171008,I171039,I260502,I171056,I260481,I260484,I171073,I171090,I171107,I171152,I171183,I171200,I171217,I260487,I171234,I171251,I171268,I171313,I260475,I171330,I260499,I171347,I171364,I171381,I171412,I171443,I171474,I171555,I171572,I253608,I253611,I171589,I171606,I253593,I171623,I253620,I171640,I171657,I253605,I171514,I171688,I171544,I171719,I253617,I171736,I253596,I253599,I171753,I171770,I171787,I171520,I171532,I171832,I171535,I171863,I171880,I171897,I253602,I171914,I171931,I171948,I171538,I171541,I171993,I253590,I172010,I253614,I172027,I172044,I172061,I171526,I172092,I171529,I172123,I171517,I172154,I171547,I171523,I172235,I172252,I261258,I261261,I172269,I172286,I261243,I172303,I261270,I172320,I172337,I261255,I172194,I172368,I172224,I172399,I261267,I172416,I261246,I261249,I172433,I172450,I172467,I172200,I172212,I172512,I172215,I172543,I172560,I172577,I261252,I172594,I172611,I172628,I172218,I172221,I172673,I261240,I172690,I261264,I172707,I172724,I172741,I172206,I172772,I172209,I172803,I172197,I172834,I172227,I172203,I172915,I172932,I172949,I172966,I172983,I173000,I173017,I172874,I173048,I172904,I173079,I173096,I173113,I173130,I173147,I172880,I172892,I173192,I172895,I173223,I173240,I173257,I173274,I173291,I173308,I172898,I172901,I173353,I173370,I173387,I173404,I173421,I172886,I173452,I172889,I173483,I172877,I173514,I172907,I172883,I173595,I173612,I334136,I334145,I173629,I173646,I334151,I173663,I334157,I173680,I173697,I334139,I173728,I173759,I334148,I173776,I334154,I173793,I173810,I173827,I173872,I173903,I173920,I334142,I173937,I173954,I173971,I173988,I174033,I334160,I174050,I174067,I174084,I174101,I174132,I174163,I174194,I174275,I174292,I174309,I174326,I174343,I174360,I174377,I174234,I174408,I174264,I174439,I174456,I174473,I174490,I174507,I174240,I174252,I174552,I174255,I174583,I174600,I174617,I174634,I174651,I174668,I174258,I174261,I174713,I174730,I174747,I174764,I174781,I174246,I174812,I174249,I174843,I174237,I174874,I174267,I174243,I174955,I174972,I392599,I392626,I174989,I175006,I392602,I175023,I392617,I175040,I175057,I392623,I174914,I175088,I174944,I175119,I392614,I175136,I392611,I392605,I175153,I175170,I175187,I174920,I174932,I175232,I174935,I175263,I175280,I175297,I392629,I175314,I175331,I175348,I174938,I174941,I175393,I175410,I392620,I175427,I392632,I392608,I175444,I175461,I174926,I175492,I174929,I175523,I174917,I175554,I174947,I174923,I175635,I175652,I239073,I239076,I175669,I175686,I239058,I175703,I239085,I175720,I175737,I239070,I175594,I175768,I175624,I175799,I239082,I175816,I239061,I239064,I175833,I175850,I175867,I175600,I175612,I175912,I175615,I175943,I175960,I175977,I239067,I175994,I176011,I176028,I175618,I175621,I176073,I239055,I176090,I239079,I176107,I176124,I176141,I175606,I176172,I175609,I176203,I175597,I176234,I175627,I175603,I176315,I176332,I176349,I176366,I176383,I176400,I176417,I176274,I176448,I176304,I176479,I176496,I176513,I176530,I176547,I176280,I176292,I176592,I176295,I176623,I176640,I176657,I176674,I176691,I176708,I176298,I176301,I176753,I176770,I176787,I176804,I176821,I176286,I176852,I176289,I176883,I176277,I176914,I176307,I176283,I176995,I177012,I245958,I245961,I177029,I177046,I245943,I177063,I245970,I177080,I177097,I245955,I176954,I177128,I176984,I177159,I245967,I177176,I245946,I245949,I177193,I177210,I177227,I176960,I176972,I177272,I176975,I177303,I177320,I177337,I245952,I177354,I177371,I177388,I176978,I176981,I177433,I245940,I177450,I245964,I177467,I177484,I177501,I176966,I177532,I176969,I177563,I176957,I177594,I176987,I176963,I177672,I177689,I177706,I177732,I177740,I177757,I177774,I177791,I177808,I177825,I177842,I177859,I177876,I177893,I177910,I177927,I177944,I177961,I177992,I178009,I178040,I178066,I178088,I178119,I178150,I178167,I178184,I178215,I178232,I178263,I178294,I178311,I178403,I178420,I267366,I267384,I178437,I267378,I178463,I178471,I267372,I178488,I178505,I267390,I178522,I178539,I267387,I178556,I178573,I267360,I267363,I178590,I178607,I178624,I178641,I178658,I267369,I178675,I178692,I178374,I178723,I178740,I178386,I178771,I267375,I178797,I178365,I178819,I178395,I178850,I178392,I178881,I178898,I267381,I178915,I178368,I178946,I178963,I178383,I178994,I178371,I179025,I179042,I178380,I178377,I178389,I179134,I179151,I425466,I425478,I179168,I425475,I179194,I179202,I425481,I179219,I179236,I425493,I179253,I425484,I179270,I425460,I179287,I179304,I425487,I179321,I179338,I179355,I179372,I179389,I425463,I179406,I179423,I179454,I179471,I179502,I425469,I425472,I179528,I179550,I179581,I179612,I179629,I425490,I179646,I179677,I179694,I179725,I179756,I179773,I179865,I179882,I317128,I317143,I179899,I317119,I179925,I179933,I317125,I179950,I179967,I317146,I179984,I317122,I180001,I317149,I180018,I180035,I317131,I317134,I180052,I180069,I180086,I180103,I180120,I180137,I180154,I180185,I180202,I180233,I180259,I180281,I180312,I180343,I180360,I317140,I317137,I180377,I180408,I180425,I180456,I180487,I180504,I180596,I180613,I180630,I180656,I180664,I180681,I180698,I180715,I180732,I180749,I180766,I180783,I180800,I180817,I180834,I180851,I180868,I180885,I180567,I180916,I180933,I180579,I180964,I180990,I180558,I181012,I180588,I181043,I180585,I181074,I181091,I181108,I180561,I181139,I181156,I180576,I181187,I180564,I181218,I181235,I180573,I180570,I180582,I181327,I181344,I249006,I249024,I181361,I249018,I181387,I181395,I249012,I181412,I181429,I249030,I181446,I181463,I249027,I181480,I181497,I249000,I249003,I181514,I181531,I181548,I181565,I181582,I249009,I181599,I181616,I181298,I181647,I181664,I181310,I181695,I249015,I181721,I181289,I181743,I181319,I181774,I181316,I181805,I181822,I249021,I181839,I181292,I181870,I181887,I181307,I181918,I181295,I181949,I181966,I181304,I181301,I181313,I182058,I182075,I318590,I318605,I182092,I318581,I182118,I182126,I318587,I182143,I182160,I318608,I182177,I318584,I182194,I318611,I182211,I182228,I318593,I318596,I182245,I182262,I182279,I182296,I182313,I182330,I182347,I182029,I182378,I182395,I182041,I182426,I182452,I182020,I182474,I182050,I182505,I182047,I182536,I182553,I318602,I318599,I182570,I182023,I182601,I182618,I182038,I182649,I182026,I182680,I182697,I182035,I182032,I182044,I182783,I182800,I294479,I294461,I182817,I294470,I182843,I182851,I182868,I294464,I182885,I182902,I294488,I182919,I294467,I182936,I182953,I182984,I183001,I294473,I183018,I294458,I183035,I183052,I183069,I294485,I183086,I183103,I183120,I183151,I183168,I183185,I294476,I294482,I183216,I183233,I183264,I183281,I183298,I183329,I183360,I183405,I183422,I183480,I183497,I265833,I265830,I183514,I265836,I183540,I183548,I183565,I265842,I183582,I183599,I183616,I265839,I183633,I183650,I183460,I183681,I183698,I265860,I183715,I265848,I183732,I183749,I183766,I265851,I183783,I265845,I183800,I183817,I183451,I183848,I183865,I183882,I265854,I265857,I183448,I183913,I183930,I183472,I183961,I183978,I183995,I183454,I184026,I183463,I184057,I183469,I183466,I184102,I184119,I183457,I184177,I184194,I269658,I269655,I184211,I269661,I184237,I184245,I184262,I269667,I184279,I184296,I184313,I269664,I184330,I184347,I184378,I184395,I269685,I184412,I269673,I184429,I184446,I184463,I269676,I184480,I269670,I184497,I184514,I184545,I184562,I184579,I269679,I269682,I184610,I184627,I184658,I184675,I184692,I184723,I184754,I184799,I184816,I184874,I184891,I428954,I428945,I184908,I428948,I184934,I184942,I184959,I428963,I184976,I184993,I428975,I185010,I428972,I428966,I185027,I185044,I184854,I185075,I185092,I428969,I185109,I428951,I185126,I185143,I185160,I428960,I185177,I428957,I185194,I185211,I184845,I185242,I185259,I185276,I428978,I184842,I185307,I185324,I184866,I185355,I185372,I185389,I184848,I185420,I184857,I185451,I184863,I184860,I185496,I185513,I184851,I185571,I185588,I185605,I185631,I185639,I185656,I185673,I185690,I185707,I185724,I185741,I185772,I185789,I185806,I185823,I185840,I185857,I185874,I185891,I185908,I185939,I185956,I185973,I186004,I186021,I186052,I186069,I186086,I186117,I186148,I186193,I186210,I186268,I186285,I186302,I186328,I186336,I186353,I186370,I186387,I186404,I186421,I186438,I186248,I186469,I186486,I186503,I186520,I186537,I186554,I186571,I186588,I186605,I186239,I186636,I186653,I186670,I186236,I186701,I186718,I186260,I186749,I186766,I186783,I186242,I186814,I186251,I186845,I186257,I186254,I186890,I186907,I186245,I186965,I186982,I255123,I255120,I186999,I255126,I187025,I187033,I187050,I255132,I187067,I187084,I187101,I255129,I187118,I187135,I187166,I187183,I255150,I187200,I255138,I187217,I187234,I187251,I255141,I187268,I255135,I187285,I187302,I187333,I187350,I187367,I255144,I255147,I187398,I187415,I187446,I187463,I187480,I187511,I187542,I187587,I187604,I187662,I187679,I187696,I187722,I187730,I187747,I187764,I187781,I187798,I187815,I187832,I187642,I187863,I187880,I187897,I187914,I187931,I187948,I187965,I187982,I187999,I187633,I188030,I188047,I188064,I187630,I188095,I188112,I187654,I188143,I188160,I188177,I187636,I188208,I187645,I188239,I187651,I187648,I188284,I188301,I187639,I188359,I188376,I213463,I213436,I188393,I213448,I188419,I188427,I188444,I213454,I188461,I188478,I213451,I188495,I213445,I188512,I188529,I188560,I188577,I213460,I188594,I213439,I188611,I188628,I188645,I213457,I188662,I213442,I188679,I188696,I188727,I188744,I188761,I188792,I188809,I188840,I188857,I188874,I188905,I188936,I188981,I188998,I189056,I189073,I275013,I275010,I189090,I275016,I189116,I189124,I189141,I275022,I189158,I189175,I189192,I275019,I189209,I189226,I189036,I189257,I189274,I275040,I189291,I275028,I189308,I189325,I189342,I275031,I189359,I275025,I189376,I189393,I189027,I189424,I189441,I189458,I275034,I275037,I189024,I189489,I189506,I189048,I189537,I189554,I189571,I189030,I189602,I189039,I189633,I189045,I189042,I189678,I189695,I189033,I189753,I189770,I316409,I316391,I189787,I316400,I189813,I189821,I189838,I316394,I189855,I189872,I316418,I189889,I316397,I189906,I189923,I189954,I189971,I316403,I189988,I316388,I190005,I190022,I190039,I316415,I190056,I190073,I190090,I190121,I190138,I190155,I316406,I316412,I190186,I190203,I190234,I190251,I190268,I190299,I190330,I190375,I190392,I190450,I190467,I190484,I190510,I190518,I190535,I190552,I190569,I190586,I190603,I190620,I190651,I190668,I190685,I190702,I190719,I190736,I190753,I190770,I190787,I190818,I190835,I190852,I190883,I190900,I190931,I190948,I190965,I190996,I191027,I191072,I191089,I191147,I191164,I233703,I233700,I191181,I233706,I191207,I191215,I191232,I233712,I191249,I191266,I191283,I233709,I191300,I191317,I191127,I191348,I191365,I233730,I191382,I233718,I191399,I191416,I191433,I233721,I191450,I233715,I191467,I191484,I191118,I191515,I191532,I191549,I233724,I233727,I191115,I191580,I191597,I191139,I191628,I191645,I191662,I191121,I191693,I191130,I191724,I191136,I191133,I191769,I191786,I191124,I191844,I191861,I350201,I350213,I191878,I350204,I191904,I191912,I191929,I350216,I191946,I191963,I350222,I191980,I350207,I350210,I191997,I192014,I192045,I192062,I350219,I192079,I192096,I192113,I192130,I350225,I192147,I192164,I192181,I192212,I192229,I192246,I192277,I192294,I192325,I192342,I192359,I192390,I192421,I192466,I192483,I192541,I192558,I192575,I192601,I192609,I192626,I192643,I192660,I192677,I192694,I192711,I192521,I192742,I192759,I192776,I192793,I192810,I192827,I192844,I192861,I192878,I192512,I192909,I192926,I192943,I192509,I192974,I192991,I192533,I193022,I193039,I193056,I192515,I193087,I192524,I193118,I192530,I192527,I193163,I193180,I192518,I193238,I193255,I220195,I220168,I193272,I220180,I193298,I193306,I193323,I220186,I193340,I193357,I220183,I193374,I220177,I193391,I193408,I193439,I193456,I220192,I193473,I220171,I193490,I193507,I193524,I220189,I193541,I220174,I193558,I193575,I193606,I193623,I193640,I193671,I193688,I193719,I193736,I193753,I193784,I193815,I193860,I193877,I193935,I193952,I362101,I362113,I193969,I362104,I193995,I194003,I194020,I362116,I194037,I194054,I362122,I194071,I362107,I362110,I194088,I194105,I193915,I194136,I194153,I362119,I194170,I194187,I194204,I194221,I362125,I194238,I194255,I194272,I193906,I194303,I194320,I194337,I193903,I194368,I194385,I193927,I194416,I194433,I194450,I193909,I194481,I193918,I194512,I193924,I193921,I194557,I194574,I193912,I194632,I194649,I343061,I343073,I194666,I343064,I194692,I194700,I194717,I343076,I194734,I194751,I343082,I194768,I343067,I343070,I194785,I194802,I194612,I194833,I194850,I343079,I194867,I194884,I194901,I194918,I343085,I194935,I194952,I194969,I194603,I195000,I195017,I195034,I194600,I195065,I195082,I194624,I195113,I195130,I195147,I194606,I195178,I194615,I195209,I194621,I194618,I195254,I195271,I194609,I195329,I195346,I284976,I284958,I195363,I284967,I195389,I195397,I195414,I284961,I195431,I195448,I284985,I195465,I284964,I195482,I195499,I195309,I195530,I195547,I284970,I195564,I284955,I195581,I195598,I195615,I284982,I195632,I195649,I195666,I195300,I195697,I195714,I195731,I284973,I284979,I195297,I195762,I195779,I195321,I195810,I195827,I195844,I195303,I195875,I195312,I195906,I195318,I195315,I195951,I195968,I195306,I196026,I196043,I314947,I314929,I196060,I314938,I196086,I196094,I196111,I314932,I196128,I196145,I314956,I196162,I314935,I196179,I196196,I196227,I196244,I314941,I196261,I314926,I196278,I196295,I196312,I314953,I196329,I196346,I196363,I196394,I196411,I196428,I314944,I314950,I196459,I196476,I196507,I196524,I196541,I196572,I196603,I196648,I196665,I196723,I196740,I196757,I196783,I196791,I196808,I196825,I196842,I196859,I196876,I196893,I196703,I196924,I196941,I196958,I196975,I196992,I197009,I197026,I197043,I197060,I196694,I197091,I197108,I197125,I196691,I197156,I197173,I196715,I197204,I197221,I197238,I196697,I197269,I196706,I197300,I196712,I196709,I197345,I197362,I196700,I197420,I197437,I197454,I197480,I197488,I197505,I197522,I197539,I197556,I197573,I197590,I197400,I197621,I197638,I197655,I197672,I197689,I197706,I197723,I197740,I197757,I197391,I197788,I197805,I197822,I197388,I197853,I197870,I197412,I197901,I197918,I197935,I197394,I197966,I197403,I197997,I197409,I197406,I198042,I198059,I197397,I198117,I198134,I369683,I369695,I198151,I369689,I198177,I198185,I198202,I198219,I198236,I369704,I198253,I369692,I369713,I198270,I198287,I198097,I198318,I198335,I369698,I198352,I369707,I198369,I198386,I198403,I369716,I369710,I198420,I369686,I198437,I198454,I198088,I198485,I198502,I198519,I369701,I198085,I198550,I198567,I198109,I198598,I198615,I198632,I198091,I198663,I198100,I198694,I198106,I198103,I198739,I198756,I198094,I198814,I198831,I258948,I258945,I198848,I258951,I198874,I198882,I198899,I258957,I198916,I198933,I198950,I258954,I198967,I198984,I198794,I199015,I199032,I258975,I199049,I258963,I199066,I199083,I199100,I258966,I199117,I258960,I199134,I199151,I198785,I199182,I199199,I199216,I258969,I258972,I198782,I199247,I199264,I198806,I199295,I199312,I199329,I198788,I199360,I198797,I199391,I198803,I198800,I199436,I199453,I198791,I199511,I199528,I431045,I431036,I199545,I431039,I199571,I199579,I199596,I431054,I199613,I199630,I431066,I199647,I431063,I431057,I199664,I199681,I199712,I199729,I431060,I199746,I431042,I199763,I199780,I199797,I431051,I199814,I431048,I199831,I199848,I199879,I199896,I199913,I431069,I199944,I199961,I199992,I200009,I200026,I200057,I200088,I200133,I200150,I200208,I200225,I326996,I327008,I200242,I326999,I200268,I200276,I200293,I327011,I200310,I200327,I327017,I200344,I327002,I327005,I200361,I200378,I200188,I200409,I200426,I327014,I200443,I200460,I200477,I200494,I327020,I200511,I200528,I200545,I200179,I200576,I200593,I200610,I200176,I200641,I200658,I200200,I200689,I200706,I200723,I200182,I200754,I200191,I200785,I200197,I200194,I200830,I200847,I200185,I200905,I200922,I200939,I200965,I200973,I200990,I201007,I201024,I201041,I201058,I201075,I201106,I201123,I201140,I201157,I201174,I201191,I201208,I201225,I201242,I201273,I201290,I201307,I201338,I201355,I201386,I201403,I201420,I201451,I201482,I201527,I201544,I201602,I201619,I256653,I256650,I201636,I256656,I201662,I201670,I201687,I256662,I201704,I201721,I201738,I256659,I201755,I201772,I201582,I201803,I201820,I256680,I201837,I256668,I201854,I201871,I201888,I256671,I201905,I256665,I201922,I201939,I201573,I201970,I201987,I202004,I256674,I256677,I201570,I202035,I202052,I201594,I202083,I202100,I202117,I201576,I202148,I201585,I202179,I201591,I201588,I202224,I202241,I201579,I202299,I202316,I322831,I322843,I202333,I322834,I202359,I202367,I202384,I322846,I202401,I202418,I322852,I202435,I322837,I322840,I202452,I202469,I202500,I202517,I322849,I202534,I202551,I202568,I202585,I322855,I202602,I202619,I202636,I202667,I202684,I202701,I202732,I202749,I202780,I202797,I202814,I202845,I202876,I202921,I202938,I202999,I203016,I203033,I203059,I203067,I203084,I203101,I203118,I203135,I203152,I203169,I203186,I203203,I203220,I203237,I203254,I203271,I203288,I202991,I203319,I203336,I203353,I203370,I202973,I203401,I203418,I202967,I203449,I203475,I203483,I202970,I202964,I202982,I203542,I203559,I203576,I203593,I202985,I203624,I202988,I203655,I202979,I203686,I202976,I203747,I203764,I281151,I281136,I203781,I281130,I203807,I203815,I203832,I281133,I203849,I203866,I281160,I281154,I203883,I203900,I203917,I281157,I203934,I203951,I203968,I281145,I203985,I204002,I204019,I204036,I204067,I281139,I204084,I204101,I204118,I204149,I281142,I204166,I204197,I204223,I204231,I204290,I204307,I281148,I204324,I204341,I204372,I204403,I204434,I204495,I204512,I204529,I204555,I204563,I204580,I204597,I204614,I204631,I204648,I204665,I204682,I204699,I204716,I204733,I204750,I204767,I204784,I204487,I204815,I204832,I204849,I204866,I204469,I204897,I204914,I204463,I204945,I204971,I204979,I204466,I204460,I204478,I205038,I205055,I205072,I205089,I204481,I205120,I204484,I205151,I204475,I205182,I204472,I205243,I205260,I205277,I205303,I205311,I205328,I205345,I205362,I205379,I205396,I205413,I205430,I205447,I205464,I205481,I205498,I205515,I205532,I205235,I205563,I205580,I205597,I205614,I205217,I205645,I205662,I205211,I205693,I205719,I205727,I205214,I205208,I205226,I205786,I205803,I205820,I205837,I205229,I205868,I205232,I205899,I205223,I205930,I205220,I205991,I206008,I381635,I381617,I206025,I381641,I206051,I206059,I206076,I381644,I206093,I206110,I381650,I381632,I206127,I206144,I206161,I381626,I206178,I206195,I206212,I381623,I206229,I381638,I206246,I206263,I206280,I205983,I206311,I381620,I206328,I206345,I206362,I205965,I206393,I206410,I205959,I206441,I381647,I206467,I206475,I205962,I205956,I205974,I206534,I381629,I206551,I206568,I206585,I205977,I206616,I205980,I206647,I205971,I206678,I205968,I206739,I206756,I206773,I206799,I206807,I206824,I206841,I206858,I206875,I206892,I206909,I206926,I206943,I206960,I206977,I206994,I207011,I207028,I207059,I207076,I207093,I207110,I207141,I207158,I207189,I207215,I207223,I207282,I207299,I207316,I207333,I207364,I207395,I207426,I207487,I207504,I207521,I207547,I207555,I207572,I207589,I207606,I207623,I207640,I207657,I207674,I207691,I207708,I207725,I207742,I207759,I207776,I207479,I207807,I207824,I207841,I207858,I207461,I207889,I207906,I207455,I207937,I207963,I207971,I207458,I207452,I207470,I208030,I208047,I208064,I208081,I207473,I208112,I207476,I208143,I207467,I208174,I207464,I208235,I208252,I390033,I390015,I208269,I390039,I208295,I208303,I208320,I390042,I208337,I208354,I390048,I390030,I208371,I208388,I208405,I390024,I208422,I208439,I208456,I390021,I208473,I390036,I208490,I208507,I208524,I208227,I208555,I390018,I208572,I208589,I208606,I208209,I208637,I208654,I208203,I208685,I390045,I208711,I208719,I208206,I208200,I208218,I208778,I390027,I208795,I208812,I208829,I208221,I208860,I208224,I208891,I208215,I208922,I208212,I208983,I209000,I209017,I209043,I209051,I209068,I209085,I209102,I209119,I209136,I209153,I209170,I209187,I209204,I209221,I209238,I209255,I209272,I209303,I209320,I209337,I209354,I209385,I209402,I209433,I209459,I209467,I209526,I209543,I209560,I209577,I209608,I209639,I209670,I209731,I209748,I301774,I301771,I209765,I301768,I209791,I209799,I209816,I301777,I209833,I209850,I301795,I209867,I209884,I209901,I301798,I209918,I209935,I209952,I301783,I209969,I301789,I209986,I210003,I210020,I209723,I210051,I210068,I210085,I210102,I209705,I210133,I210150,I209699,I210181,I210207,I210215,I209702,I209696,I209714,I210274,I301780,I301786,I210291,I301792,I210308,I210325,I209717,I210356,I209720,I210387,I209711,I210418,I209708,I210479,I210496,I210513,I210539,I210547,I210564,I210581,I210598,I210615,I210632,I210649,I210666,I210683,I210700,I210717,I210734,I210751,I210768,I210799,I210816,I210833,I210850,I210881,I210898,I210929,I210955,I210963,I211022,I211039,I211056,I211073,I211104,I211135,I211166,I211227,I211244,I266616,I266601,I211261,I266595,I211287,I211295,I211312,I266598,I211329,I211346,I266625,I266619,I211363,I211380,I211397,I266622,I211414,I211431,I211448,I266610,I211465,I211482,I211499,I211516,I211547,I266604,I211564,I211581,I211598,I211629,I266607,I211646,I211677,I211703,I211711,I211770,I211787,I266613,I211804,I211821,I211852,I211883,I211914,I211975,I211992,I212009,I212035,I212043,I212060,I212077,I212094,I212111,I212128,I212145,I212162,I212179,I212196,I212213,I212230,I212247,I212264,I212295,I212312,I212329,I212346,I212377,I212394,I212425,I212451,I212459,I212518,I212535,I212552,I212569,I212600,I212631,I212662,I212723,I212740,I212757,I212783,I212791,I212808,I212825,I212842,I212859,I212876,I212893,I212910,I212927,I212944,I212961,I212978,I212995,I213012,I212715,I213043,I213060,I213077,I213094,I212697,I213125,I213142,I212691,I213173,I213199,I213207,I212694,I212688,I212706,I213266,I213283,I213300,I213317,I212709,I213348,I212712,I213379,I212703,I213410,I212700,I213471,I213488,I213505,I213531,I213539,I213556,I213573,I213590,I213607,I213624,I213641,I213658,I213675,I213692,I213709,I213726,I213743,I213760,I213791,I213808,I213825,I213842,I213873,I213890,I213921,I213947,I213955,I214014,I214031,I214048,I214065,I214096,I214127,I214158,I214219,I214236,I214253,I214279,I214287,I214304,I214321,I214338,I214355,I214372,I214389,I214406,I214423,I214440,I214457,I214474,I214491,I214508,I214539,I214556,I214573,I214590,I214621,I214638,I214669,I214695,I214703,I214762,I214779,I214796,I214813,I214844,I214875,I214906,I214967,I214984,I215001,I215027,I215035,I215052,I215069,I215086,I215103,I215120,I215137,I215154,I215171,I215188,I215205,I215222,I215239,I215256,I215287,I215304,I215321,I215338,I215369,I215386,I215417,I215443,I215451,I215510,I215527,I215544,I215561,I215592,I215623,I215654,I215715,I215732,I215749,I215775,I215783,I215800,I215817,I215834,I215851,I215868,I215885,I215902,I215919,I215936,I215953,I215970,I215987,I216004,I216035,I216052,I216069,I216086,I216117,I216134,I216165,I216191,I216199,I216258,I216275,I216292,I216309,I216340,I216371,I216402,I216463,I216480,I380989,I380971,I216497,I380995,I216523,I216531,I216548,I380998,I216565,I216582,I381004,I380986,I216599,I216616,I216633,I380980,I216650,I216667,I216684,I380977,I216701,I380992,I216718,I216735,I216752,I216455,I216783,I380974,I216800,I216817,I216834,I216437,I216865,I216882,I216431,I216913,I381001,I216939,I216947,I216434,I216428,I216446,I217006,I380983,I217023,I217040,I217057,I216449,I217088,I216452,I217119,I216443,I217150,I216440,I217211,I217228,I217245,I217271,I217279,I217296,I217313,I217330,I217347,I217364,I217381,I217398,I217415,I217432,I217449,I217466,I217483,I217500,I217531,I217548,I217565,I217582,I217613,I217630,I217661,I217687,I217695,I217754,I217771,I217788,I217805,I217836,I217867,I217898,I217959,I217976,I345444,I345441,I217993,I345450,I218019,I218027,I218044,I345447,I218061,I218078,I345456,I218095,I218112,I218129,I218146,I218163,I218180,I218197,I218214,I218231,I218248,I217951,I218279,I345459,I218296,I218313,I218330,I217933,I218361,I345453,I218378,I217927,I218409,I345465,I218435,I218443,I217930,I217924,I217942,I218502,I345462,I218519,I218536,I218553,I217945,I218584,I217948,I218615,I217939,I218646,I217936,I218707,I218724,I393263,I393245,I218741,I393269,I218767,I218775,I218792,I393272,I218809,I218826,I393278,I393260,I218843,I218860,I218877,I393254,I218894,I218911,I218928,I393251,I218945,I393266,I218962,I218979,I218996,I219027,I393248,I219044,I219061,I219078,I219109,I219126,I219157,I393275,I219183,I219191,I219250,I393257,I219267,I219284,I219301,I219332,I219363,I219394,I219455,I219472,I219489,I219515,I219523,I219540,I219557,I219574,I219591,I219608,I219625,I219642,I219659,I219676,I219693,I219710,I219727,I219744,I219447,I219775,I219792,I219809,I219826,I219429,I219857,I219874,I219423,I219905,I219931,I219939,I219426,I219420,I219438,I219998,I220015,I220032,I220049,I219441,I220080,I219444,I220111,I219435,I220142,I219432,I220203,I220220,I320049,I320046,I220237,I320043,I220263,I220271,I220288,I320052,I220305,I220322,I320070,I220339,I220356,I220373,I320073,I220390,I220407,I220424,I320058,I220441,I320064,I220458,I220475,I220492,I220523,I220540,I220557,I220574,I220605,I220622,I220653,I220679,I220687,I220746,I320055,I320061,I220763,I320067,I220780,I220797,I220828,I220859,I220890,I220951,I220968,I393909,I393891,I220985,I393915,I221011,I221019,I221036,I393918,I221053,I221070,I393924,I393906,I221087,I221104,I221121,I393900,I221138,I221155,I221172,I393897,I221189,I393912,I221206,I221223,I221240,I221271,I393894,I221288,I221305,I221322,I221353,I221370,I221401,I393921,I221427,I221435,I221494,I393903,I221511,I221528,I221545,I221576,I221607,I221638,I221699,I221716,I221733,I221759,I221767,I221784,I221801,I221818,I221835,I221852,I221869,I221886,I221903,I221920,I221937,I221954,I221971,I221988,I222019,I222036,I222053,I222070,I222101,I222118,I222149,I222175,I222183,I222242,I222259,I222276,I222293,I222324,I222355,I222386,I222447,I222464,I222481,I222507,I222515,I222532,I222549,I222566,I222583,I222600,I222617,I222634,I222651,I222668,I222685,I222702,I222719,I222736,I222439,I222767,I222784,I222801,I222818,I222421,I222849,I222866,I222415,I222897,I222923,I222931,I222418,I222412,I222430,I222990,I223007,I223024,I223041,I222433,I223072,I222436,I223103,I222427,I223134,I222424,I223195,I223212,I382281,I382263,I223229,I382287,I223255,I223263,I223280,I382290,I223297,I223314,I382296,I382278,I223331,I223348,I223365,I382272,I223382,I223399,I223416,I382269,I223433,I382284,I223450,I223467,I223484,I223515,I382266,I223532,I223549,I223566,I223597,I223614,I223645,I382293,I223671,I223679,I223738,I382275,I223755,I223772,I223789,I223820,I223851,I223882,I223943,I223960,I223977,I224003,I224011,I224028,I224045,I224062,I224079,I224096,I224113,I224130,I224147,I224164,I224181,I224198,I224215,I224232,I223935,I224263,I224280,I224297,I224314,I223917,I224345,I224362,I223911,I224393,I224419,I224427,I223914,I223908,I223926,I224486,I224503,I224520,I224537,I223929,I224568,I223932,I224599,I223923,I224630,I223920,I224691,I224708,I311277,I311274,I224725,I311271,I224751,I224759,I224776,I311280,I224793,I224810,I311298,I224827,I224844,I224861,I311301,I224878,I224895,I224912,I311286,I224929,I311292,I224946,I224963,I224980,I224683,I225011,I225028,I225045,I225062,I224665,I225093,I225110,I224659,I225141,I225167,I225175,I224662,I224656,I224674,I225234,I311283,I311289,I225251,I311295,I225268,I225285,I224677,I225316,I224680,I225347,I224671,I225378,I224668,I225439,I225456,I225473,I225499,I225507,I225524,I225541,I225558,I225575,I225592,I225609,I225626,I225643,I225660,I225677,I225694,I225711,I225728,I225759,I225776,I225793,I225810,I225841,I225858,I225889,I225915,I225923,I225982,I225999,I226016,I226033,I226064,I226095,I226126,I226187,I226204,I329974,I329971,I226221,I329980,I226247,I226255,I226272,I329977,I226289,I226306,I329986,I226323,I226340,I226357,I226374,I226391,I226408,I226425,I226442,I226459,I226476,I226507,I329989,I226524,I226541,I226558,I226589,I329983,I226606,I226637,I329995,I226663,I226671,I226730,I329992,I226747,I226764,I226781,I226812,I226843,I226874,I226935,I226952,I389387,I389369,I226969,I389393,I226995,I227003,I227020,I389396,I227037,I227054,I389402,I389384,I227071,I227088,I227105,I389378,I227122,I227139,I227156,I389375,I227173,I389390,I227190,I227207,I227224,I227255,I389372,I227272,I227289,I227306,I227337,I227354,I227385,I389399,I227411,I227419,I227478,I389381,I227495,I227512,I227529,I227560,I227591,I227622,I227683,I227700,I288616,I288613,I227717,I288610,I227743,I227751,I227768,I288619,I227785,I227802,I288637,I227819,I227836,I227853,I288640,I227870,I227887,I227904,I288625,I227921,I288631,I227938,I227955,I227972,I228003,I228020,I228037,I228054,I228085,I228102,I228133,I228159,I228167,I228226,I288622,I288628,I228243,I288634,I228260,I228277,I228308,I228339,I228370,I228431,I228448,I312008,I312005,I228465,I312002,I228491,I228499,I228516,I312011,I228533,I228550,I312029,I228567,I228584,I228601,I312032,I228618,I228635,I228652,I312017,I228669,I312023,I228686,I228703,I228720,I228423,I228751,I228768,I228785,I228802,I228405,I228833,I228850,I228399,I228881,I228907,I228915,I228402,I228396,I228414,I228974,I312014,I312020,I228991,I312026,I229008,I229025,I228417,I229056,I228420,I229087,I228411,I229118,I228408,I229179,I229196,I310546,I310543,I229213,I310540,I229239,I229247,I229264,I310549,I229281,I229298,I310567,I229315,I229332,I229349,I310570,I229366,I229383,I229400,I310555,I229417,I310561,I229434,I229451,I229468,I229499,I229516,I229533,I229550,I229581,I229598,I229629,I229655,I229663,I229722,I310552,I310558,I229739,I310564,I229756,I229773,I229804,I229835,I229866,I229927,I229944,I281916,I281901,I229961,I281895,I229987,I229995,I230012,I281898,I230029,I230046,I281925,I281919,I230063,I230080,I230097,I281922,I230114,I230131,I230148,I281910,I230165,I230182,I230199,I230216,I230247,I281904,I230264,I230281,I230298,I230329,I281907,I230346,I230377,I230403,I230411,I230470,I230487,I281913,I230504,I230521,I230552,I230583,I230614,I230678,I230695,I230712,I230729,I230746,I230763,I230780,I230797,I230640,I230828,I230845,I230862,I230879,I230896,I230913,I230930,I230655,I230961,I230978,I230643,I230658,I231023,I231040,I231057,I231074,I231091,I231108,I230649,I231139,I231156,I231173,I231190,I231207,I230670,I231238,I230646,I231269,I230667,I230661,I231314,I231331,I230652,I231362,I231379,I230664,I231443,I231460,I231477,I231494,I231511,I231528,I231545,I231562,I231593,I231610,I231627,I231644,I231661,I231678,I231695,I231726,I231743,I231788,I231805,I231822,I231839,I231856,I231873,I231904,I231921,I231938,I231955,I231972,I232003,I232034,I232079,I232096,I232127,I232144,I232208,I232225,I326404,I326401,I232242,I232259,I326410,I232276,I232293,I326422,I232310,I232327,I326419,I232358,I232375,I232392,I326425,I232409,I326413,I232426,I232443,I232460,I232491,I232508,I232553,I232570,I232587,I326407,I232604,I232621,I232638,I232669,I326416,I232686,I232703,I232720,I232737,I232768,I232799,I232844,I232861,I232892,I232909,I232973,I232990,I233007,I233024,I233041,I233058,I233075,I233092,I233123,I233140,I233157,I233174,I233191,I233208,I233225,I233256,I233273,I233318,I233335,I233352,I233369,I233386,I233403,I233434,I233451,I233468,I233485,I233502,I233533,I233564,I233609,I233626,I233657,I233674,I233738,I233755,I437333,I437330,I233772,I233789,I437318,I233806,I233823,I437339,I233840,I233857,I437309,I233888,I233905,I233922,I437327,I233939,I437342,I437324,I233956,I233973,I233990,I234021,I234038,I234083,I234100,I437336,I234117,I437315,I234134,I234151,I234168,I234199,I437321,I234216,I437312,I234233,I234250,I234267,I234298,I234329,I234374,I234391,I234422,I234439,I234503,I234520,I234537,I234554,I234571,I234588,I234605,I234622,I234653,I234670,I234687,I234704,I234721,I234738,I234755,I234786,I234803,I234848,I234865,I234882,I234899,I234916,I234933,I234964,I234981,I234998,I235015,I235032,I235063,I235094,I235139,I235156,I235187,I235204,I235268,I235285,I361509,I361506,I235302,I235319,I361515,I235336,I235353,I361527,I235370,I235387,I361524,I235418,I235435,I235452,I361530,I235469,I361518,I235486,I235503,I235520,I235551,I235568,I235613,I235630,I235647,I361512,I235664,I235681,I235698,I235729,I361521,I235746,I235763,I235780,I235797,I235828,I235859,I235904,I235921,I235952,I235969,I236033,I236050,I236067,I236084,I236101,I236118,I236135,I236152,I236183,I236200,I236217,I236234,I236251,I236268,I236285,I236316,I236333,I236378,I236395,I236412,I236429,I236446,I236463,I236494,I236511,I236528,I236545,I236562,I236593,I236624,I236669,I236686,I236717,I236734,I236798,I236815,I335329,I335326,I236832,I236849,I335335,I236866,I236883,I335347,I236900,I236917,I335344,I236948,I236965,I236982,I335350,I236999,I335338,I237016,I237033,I237050,I237081,I237098,I237143,I237160,I237177,I335332,I237194,I237211,I237228,I237259,I335341,I237276,I237293,I237310,I237327,I237358,I237389,I237434,I237451,I237482,I237499,I237563,I237580,I237597,I237614,I237631,I237648,I237665,I237682,I237713,I237730,I237747,I237764,I237781,I237798,I237815,I237846,I237863,I237908,I237925,I237942,I237959,I237976,I237993,I238024,I238041,I238058,I238075,I238092,I238123,I238154,I238199,I238216,I238247,I238264,I238328,I238345,I395872,I395884,I238362,I238379,I395866,I238396,I238413,I395878,I238430,I238447,I238290,I238478,I238495,I238512,I395863,I238529,I395881,I395875,I238546,I238563,I238580,I238305,I238611,I238628,I238293,I238308,I238673,I238690,I395887,I238707,I238724,I238741,I238758,I238299,I238789,I238806,I238823,I395869,I238840,I238857,I238320,I238888,I238296,I238919,I238317,I238311,I238964,I238981,I238302,I239012,I239029,I238314,I239093,I239110,I367289,I367304,I239127,I239144,I367313,I239161,I239178,I367301,I239195,I239212,I367298,I239243,I239260,I239277,I367292,I239294,I367310,I239311,I239328,I239345,I239376,I239393,I239438,I239455,I367316,I239472,I367319,I239489,I239506,I239523,I239554,I367286,I239571,I239588,I367295,I367307,I239605,I239622,I239653,I239684,I239729,I239746,I239777,I239794,I239858,I239875,I239892,I239909,I239926,I239943,I239960,I239977,I240008,I240025,I240042,I240059,I240076,I240093,I240110,I240141,I240158,I240203,I240220,I240237,I240254,I240271,I240288,I240319,I240336,I240353,I240370,I240387,I240418,I240449,I240494,I240511,I240542,I240559,I240623,I240640,I240657,I240674,I240691,I240708,I240725,I240742,I240585,I240773,I240790,I240807,I240824,I240841,I240858,I240875,I240600,I240906,I240923,I240588,I240603,I240968,I240985,I241002,I241019,I241036,I241053,I240594,I241084,I241101,I241118,I241135,I241152,I240615,I241183,I240591,I241214,I240612,I240606,I241259,I241276,I240597,I241307,I241324,I240609,I241388,I241405,I346634,I346631,I241422,I241439,I346640,I241456,I241473,I346652,I241490,I241507,I346649,I241538,I241555,I241572,I346655,I241589,I346643,I241606,I241623,I241640,I241671,I241688,I241733,I241750,I241767,I346637,I241784,I241801,I241818,I241849,I346646,I241866,I241883,I241900,I241917,I241948,I241979,I242024,I242041,I242072,I242089,I242153,I242170,I242187,I242204,I242221,I242238,I242255,I242272,I242303,I242320,I242337,I242354,I242371,I242388,I242405,I242436,I242453,I242498,I242515,I242532,I242549,I242566,I242583,I242614,I242631,I242648,I242665,I242682,I242713,I242744,I242789,I242806,I242837,I242854,I242918,I242935,I242952,I242969,I242986,I243003,I243020,I243037,I242880,I243068,I243085,I243102,I243119,I243136,I243153,I243170,I242895,I243201,I243218,I242883,I242898,I243263,I243280,I243297,I243314,I243331,I243348,I242889,I243379,I243396,I243413,I243430,I243447,I242910,I243478,I242886,I243509,I242907,I242901,I243554,I243571,I242892,I243602,I243619,I242904,I243683,I243700,I402672,I402684,I243717,I243734,I402666,I243751,I243768,I402678,I243785,I243802,I243833,I243850,I243867,I402663,I243884,I402681,I402675,I243901,I243918,I243935,I243966,I243983,I244028,I244045,I402687,I244062,I244079,I244096,I244113,I244144,I244161,I244178,I402669,I244195,I244212,I244243,I244274,I244319,I244336,I244367,I244384,I244448,I244465,I244482,I244499,I244516,I244533,I244550,I244567,I244598,I244615,I244632,I244649,I244666,I244683,I244700,I244731,I244748,I244793,I244810,I244827,I244844,I244861,I244878,I244909,I244926,I244943,I244960,I244977,I245008,I245039,I245084,I245101,I245132,I245149,I245213,I245230,I245247,I245264,I245281,I245298,I245315,I245332,I245363,I245380,I245397,I245414,I245431,I245448,I245465,I245496,I245513,I245558,I245575,I245592,I245609,I245626,I245643,I245674,I245691,I245708,I245725,I245742,I245773,I245804,I245849,I245866,I245897,I245914,I245978,I245995,I246012,I246029,I246046,I246063,I246080,I246097,I246128,I246145,I246162,I246179,I246196,I246213,I246230,I246261,I246278,I246323,I246340,I246357,I246374,I246391,I246408,I246439,I246456,I246473,I246490,I246507,I246538,I246569,I246614,I246631,I246662,I246679,I246743,I246760,I372576,I372579,I246777,I246794,I372573,I246811,I246828,I372591,I246845,I246862,I372600,I246893,I246910,I246927,I372585,I246944,I372582,I246961,I246978,I246995,I247026,I247043,I247088,I247105,I247122,I247139,I247156,I247173,I247204,I372603,I372588,I247221,I372597,I247238,I372606,I372594,I247255,I247272,I247303,I247334,I247379,I247396,I247427,I247444,I247508,I247525,I247542,I247559,I247576,I247593,I247610,I247627,I247658,I247675,I247692,I247709,I247726,I247743,I247760,I247791,I247808,I247853,I247870,I247887,I247904,I247921,I247938,I247969,I247986,I248003,I248020,I248037,I248068,I248099,I248144,I248161,I248192,I248209,I248273,I248290,I248307,I248324,I248341,I248358,I248375,I248392,I248235,I248423,I248440,I248457,I248474,I248491,I248508,I248525,I248250,I248556,I248573,I248238,I248253,I248618,I248635,I248652,I248669,I248686,I248703,I248244,I248734,I248751,I248768,I248785,I248802,I248265,I248833,I248241,I248864,I248262,I248256,I248909,I248926,I248247,I248957,I248974,I248259,I249038,I249055,I350799,I350796,I249072,I249089,I350805,I249106,I249123,I350817,I249140,I249157,I350814,I249188,I249205,I249222,I350820,I249239,I350808,I249256,I249273,I249290,I249321,I249338,I249383,I249400,I249417,I350802,I249434,I249451,I249468,I249499,I350811,I249516,I249533,I249550,I249567,I249598,I249629,I249674,I249691,I249722,I249739,I249803,I249820,I399952,I399964,I249837,I249854,I399946,I249871,I249888,I399958,I249905,I249922,I249953,I249970,I249987,I399943,I250004,I399961,I399955,I250021,I250038,I250055,I250086,I250103,I250148,I250165,I399967,I250182,I250199,I250216,I250233,I250264,I250281,I250298,I399949,I250315,I250332,I250363,I250394,I250439,I250456,I250487,I250504,I250568,I250585,I250602,I250619,I250636,I250653,I250670,I250687,I250718,I250735,I250752,I250769,I250786,I250803,I250820,I250851,I250868,I250913,I250930,I250947,I250964,I250981,I250998,I251029,I251046,I251063,I251080,I251097,I251128,I251159,I251204,I251221,I251252,I251269,I251333,I251350,I349609,I349606,I251367,I251384,I349615,I251401,I251418,I349627,I251435,I251452,I349624,I251295,I251483,I251500,I251517,I349630,I251534,I349618,I251551,I251568,I251585,I251310,I251616,I251633,I251298,I251313,I251678,I251695,I251712,I349612,I251729,I251746,I251763,I251304,I251794,I349621,I251811,I251828,I251845,I251862,I251325,I251893,I251301,I251924,I251322,I251316,I251969,I251986,I251307,I252017,I252034,I251319,I252098,I252115,I252132,I252149,I252166,I252183,I252200,I252217,I252248,I252265,I252282,I252299,I252316,I252333,I252350,I252381,I252398,I252443,I252460,I252477,I252494,I252511,I252528,I252559,I252576,I252593,I252610,I252627,I252658,I252689,I252734,I252751,I252782,I252799,I252863,I252880,I306154,I306172,I252897,I252914,I306157,I252931,I252948,I306166,I252965,I252982,I306178,I253013,I253030,I253047,I306175,I253064,I306181,I253081,I253098,I253115,I253146,I253163,I253208,I253225,I306160,I253242,I306163,I253259,I253276,I253293,I253324,I306184,I253341,I253358,I306169,I253375,I253392,I253423,I253454,I253499,I253516,I253547,I253564,I253628,I253645,I376452,I376455,I253662,I253679,I376449,I253696,I253713,I376467,I253730,I253747,I376476,I253778,I253795,I253812,I376461,I253829,I376458,I253846,I253863,I253880,I253911,I253928,I253973,I253990,I254007,I254024,I254041,I254058,I254089,I376479,I376464,I254106,I376473,I254123,I376482,I376470,I254140,I254157,I254188,I254219,I254264,I254281,I254312,I254329,I254393,I254410,I414332,I414329,I254427,I254444,I414317,I254461,I254478,I414338,I254495,I254512,I414308,I254543,I254560,I254577,I414326,I254594,I414341,I414323,I254611,I254628,I254645,I254676,I254693,I254738,I254755,I414335,I254772,I414314,I254789,I254806,I254823,I254854,I414320,I254871,I414311,I254888,I254905,I254922,I254953,I254984,I255029,I255046,I255077,I255094,I255158,I255175,I255192,I255209,I255226,I255243,I255260,I255277,I255308,I255325,I255342,I255359,I255376,I255393,I255410,I255441,I255458,I255503,I255520,I255537,I255554,I255571,I255588,I255619,I255636,I255653,I255670,I255687,I255718,I255749,I255794,I255811,I255842,I255859,I255923,I255940,I255957,I255974,I255991,I256008,I256025,I256042,I255885,I256073,I256090,I256107,I256124,I256141,I256158,I256175,I255900,I256206,I256223,I255888,I255903,I256268,I256285,I256302,I256319,I256336,I256353,I255894,I256384,I256401,I256418,I256435,I256452,I255915,I256483,I255891,I256514,I255912,I255906,I256559,I256576,I255897,I256607,I256624,I255909,I256688,I256705,I340684,I340681,I256722,I256739,I340690,I256756,I256773,I340702,I256790,I256807,I340699,I256838,I256855,I256872,I340705,I256889,I340693,I256906,I256923,I256940,I256971,I256988,I257033,I257050,I257067,I340687,I257084,I257101,I257118,I257149,I340696,I257166,I257183,I257200,I257217,I257248,I257279,I257324,I257341,I257372,I257389,I257453,I257470,I435939,I435936,I257487,I257504,I435924,I257521,I257538,I435945,I257555,I257572,I435915,I257415,I257603,I257620,I257637,I435933,I257654,I435948,I435930,I257671,I257688,I257705,I257430,I257736,I257753,I257418,I257433,I257798,I257815,I435942,I257832,I435921,I257849,I257866,I257883,I257424,I257914,I435927,I257931,I435918,I257948,I257965,I257982,I257445,I258013,I257421,I258044,I257442,I257436,I258089,I258106,I257427,I258137,I258154,I257439,I258218,I258235,I408792,I408804,I258252,I258269,I408786,I258286,I258303,I408798,I258320,I258337,I258180,I258368,I258385,I258402,I408783,I258419,I408801,I408795,I258436,I258453,I258470,I258195,I258501,I258518,I258183,I258198,I258563,I258580,I408807,I258597,I258614,I258631,I258648,I258189,I258679,I258696,I258713,I408789,I258730,I258747,I258210,I258778,I258186,I258809,I258207,I258201,I258854,I258871,I258192,I258902,I258919,I258204,I258983,I259000,I259017,I259034,I259051,I259068,I259085,I259102,I259133,I259150,I259167,I259184,I259201,I259218,I259235,I259266,I259283,I259328,I259345,I259362,I259379,I259396,I259413,I259444,I259461,I259478,I259495,I259512,I259543,I259574,I259619,I259636,I259667,I259684,I259748,I259765,I291534,I291552,I259782,I259799,I291537,I259816,I259833,I291546,I259850,I259867,I291558,I259898,I259915,I259932,I291555,I259949,I291561,I259966,I259983,I260000,I260031,I260048,I260093,I260110,I291540,I260127,I291543,I260144,I260161,I260178,I260209,I291564,I260226,I260243,I291549,I260260,I260277,I260308,I260339,I260384,I260401,I260432,I260449,I260513,I260530,I260547,I260564,I260581,I260598,I260615,I260632,I260663,I260680,I260697,I260714,I260731,I260748,I260765,I260796,I260813,I260858,I260875,I260892,I260909,I260926,I260943,I260974,I260991,I261008,I261025,I261042,I261073,I261104,I261149,I261166,I261197,I261214,I261278,I261295,I261312,I261329,I261346,I261363,I261380,I261397,I261428,I261445,I261462,I261479,I261496,I261513,I261530,I261561,I261578,I261623,I261640,I261657,I261674,I261691,I261708,I261739,I261756,I261773,I261790,I261807,I261838,I261869,I261914,I261931,I261962,I261979,I262043,I262060,I262077,I262094,I262111,I262128,I262145,I262162,I262005,I262193,I262210,I262227,I262244,I262261,I262278,I262295,I262020,I262326,I262343,I262008,I262023,I262388,I262405,I262422,I262439,I262456,I262473,I262014,I262504,I262521,I262538,I262555,I262572,I262035,I262603,I262011,I262634,I262032,I262026,I262679,I262696,I262017,I262727,I262744,I262029,I262808,I262825,I436636,I436633,I262842,I262859,I436621,I262876,I262893,I436642,I262910,I262927,I436612,I262770,I262958,I262975,I262992,I436630,I263009,I436645,I436627,I263026,I263043,I263060,I262785,I263091,I263108,I262773,I262788,I263153,I263170,I436639,I263187,I436618,I263204,I263221,I263238,I262779,I263269,I436624,I263286,I436615,I263303,I263320,I263337,I262800,I263368,I262776,I263399,I262797,I262791,I263444,I263461,I262782,I263492,I263509,I262794,I263573,I263590,I263607,I263624,I263641,I263658,I263675,I263692,I263535,I263723,I263740,I263757,I263774,I263791,I263808,I263825,I263550,I263856,I263873,I263538,I263553,I263918,I263935,I263952,I263969,I263986,I264003,I263544,I264034,I264051,I264068,I264085,I264102,I263565,I264133,I263541,I264164,I263562,I263556,I264209,I264226,I263547,I264257,I264274,I263559,I264338,I264355,I264372,I264389,I264406,I264423,I264440,I264457,I264300,I264488,I264505,I264522,I264539,I264556,I264573,I264590,I264315,I264621,I264638,I264303,I264318,I264683,I264700,I264717,I264734,I264751,I264768,I264309,I264799,I264816,I264833,I264850,I264867,I264330,I264898,I264306,I264929,I264327,I264321,I264974,I264991,I264312,I265022,I265039,I264324,I265103,I265120,I319312,I319330,I265137,I265154,I319315,I265171,I265188,I319324,I265205,I265222,I319336,I265065,I265253,I265270,I265287,I319333,I265304,I319339,I265321,I265338,I265355,I265080,I265386,I265403,I265068,I265083,I265448,I265465,I319318,I265482,I319321,I265499,I265516,I265533,I265074,I265564,I319342,I265581,I265598,I319327,I265615,I265632,I265095,I265663,I265071,I265694,I265092,I265086,I265739,I265756,I265077,I265787,I265804,I265089,I265868,I265885,I313464,I313482,I265902,I265919,I313467,I265936,I265953,I313476,I265970,I265987,I313488,I266018,I266035,I266052,I313485,I266069,I313491,I266086,I266103,I266120,I266151,I266168,I266213,I266230,I313470,I266247,I313473,I266264,I266281,I266298,I266329,I313494,I266346,I266363,I313479,I266380,I266397,I266428,I266459,I266504,I266521,I266552,I266569,I266633,I266650,I338304,I338301,I266667,I266684,I338310,I266701,I266718,I338322,I266735,I266752,I338319,I266783,I266800,I266817,I338325,I266834,I338313,I266851,I266868,I266885,I266916,I266933,I266978,I266995,I267012,I338307,I267029,I267046,I267063,I267094,I338316,I267111,I267128,I267145,I267162,I267193,I267224,I267269,I267286,I267317,I267334,I267398,I267415,I370485,I370500,I267432,I267449,I370509,I267466,I267483,I370497,I267500,I267517,I370494,I267548,I267565,I267582,I370488,I267599,I370506,I267616,I267633,I267650,I267681,I267698,I267743,I267760,I370512,I267777,I370515,I267794,I267811,I267828,I267859,I370482,I267876,I267893,I370491,I370503,I267910,I267927,I267958,I267989,I268034,I268051,I268082,I268099,I268163,I268180,I268197,I268214,I268231,I268248,I268265,I268282,I268313,I268330,I268347,I268364,I268381,I268398,I268415,I268446,I268463,I268508,I268525,I268542,I268559,I268576,I268593,I268624,I268641,I268658,I268675,I268692,I268723,I268754,I268799,I268816,I268847,I268864,I268928,I268945,I410152,I410164,I268962,I268979,I410146,I268996,I269013,I410158,I269030,I269047,I269078,I269095,I269112,I410143,I269129,I410161,I410155,I269146,I269163,I269180,I269211,I269228,I269273,I269290,I410167,I269307,I269324,I269341,I269358,I269389,I269406,I269423,I410149,I269440,I269457,I269488,I269519,I269564,I269581,I269612,I269629,I269693,I269710,I344849,I344846,I269727,I269744,I344855,I269761,I269778,I344867,I269795,I269812,I344864,I269843,I269860,I269877,I344870,I269894,I344858,I269911,I269928,I269945,I269976,I269993,I270038,I270055,I270072,I344852,I270089,I270106,I270123,I270154,I344861,I270171,I270188,I270205,I270222,I270253,I270284,I270329,I270346,I270377,I270394,I270458,I270475,I270492,I270509,I270526,I270543,I270560,I270577,I270420,I270608,I270625,I270642,I270659,I270676,I270693,I270710,I270435,I270741,I270758,I270423,I270438,I270803,I270820,I270837,I270854,I270871,I270888,I270429,I270919,I270936,I270953,I270970,I270987,I270450,I271018,I270426,I271049,I270447,I270441,I271094,I271111,I270432,I271142,I271159,I270444,I271223,I271240,I271257,I271274,I271291,I271308,I271325,I271342,I271373,I271390,I271407,I271424,I271441,I271458,I271475,I271506,I271523,I271568,I271585,I271602,I271619,I271636,I271653,I271684,I271701,I271718,I271735,I271752,I271783,I271814,I271859,I271876,I271907,I271924,I271988,I272005,I344254,I344251,I272022,I272039,I344260,I272056,I272073,I344272,I272090,I272107,I344269,I272138,I272155,I272172,I344275,I272189,I344263,I272206,I272223,I272240,I272271,I272288,I272333,I272350,I272367,I344257,I272384,I272401,I272418,I272449,I344266,I272466,I272483,I272500,I272517,I272548,I272579,I272624,I272641,I272672,I272689,I272753,I272770,I272787,I272804,I272821,I272838,I272855,I272872,I272903,I272920,I272937,I272954,I272971,I272988,I273005,I273036,I273053,I273098,I273115,I273132,I273149,I273166,I273183,I273214,I273231,I273248,I273265,I273282,I273313,I273344,I273389,I273406,I273437,I273454,I273518,I273535,I420605,I420602,I273552,I273569,I420590,I273586,I273603,I420611,I273620,I273637,I420581,I273480,I273668,I273685,I273702,I420599,I273719,I420614,I420596,I273736,I273753,I273770,I273495,I273801,I273818,I273483,I273498,I273863,I273880,I420608,I273897,I420587,I273914,I273931,I273948,I273489,I273979,I420593,I273996,I420584,I274013,I274030,I274047,I273510,I274078,I273486,I274109,I273507,I273501,I274154,I274171,I273492,I274202,I274219,I273504,I274283,I274300,I293727,I293745,I274317,I274334,I293730,I274351,I274368,I293739,I274385,I274402,I293751,I274433,I274450,I274467,I293748,I274484,I293754,I274501,I274518,I274535,I274566,I274583,I274628,I274645,I293733,I274662,I293736,I274679,I274696,I274713,I274744,I293757,I274761,I274778,I293742,I274795,I274812,I274843,I274874,I274919,I274936,I274967,I274984,I275048,I275065,I275082,I275099,I275116,I275133,I275150,I275167,I275198,I275215,I275232,I275249,I275266,I275283,I275300,I275331,I275348,I275393,I275410,I275427,I275444,I275461,I275478,I275509,I275526,I275543,I275560,I275577,I275608,I275639,I275684,I275701,I275732,I275749,I275813,I275830,I275847,I275864,I275881,I275898,I275915,I275932,I275963,I275980,I275997,I276014,I276031,I276048,I276065,I276096,I276113,I276158,I276175,I276192,I276209,I276226,I276243,I276274,I276291,I276308,I276325,I276342,I276373,I276404,I276449,I276466,I276497,I276514,I276578,I276595,I276612,I276629,I276646,I276663,I276680,I276697,I276728,I276745,I276762,I276779,I276796,I276813,I276830,I276861,I276878,I276923,I276940,I276957,I276974,I276991,I277008,I277039,I277056,I277073,I277090,I277107,I277138,I277169,I277214,I277231,I277262,I277279,I277343,I277360,I277377,I277394,I277411,I277428,I277445,I277462,I277493,I277510,I277527,I277544,I277561,I277578,I277595,I277626,I277643,I277688,I277705,I277722,I277739,I277756,I277773,I277804,I277821,I277838,I277855,I277872,I277903,I277934,I277979,I277996,I278027,I278044,I278108,I278125,I278142,I278159,I278176,I278193,I278210,I278227,I278258,I278275,I278292,I278309,I278326,I278343,I278360,I278391,I278408,I278453,I278470,I278487,I278504,I278521,I278538,I278569,I278586,I278603,I278620,I278637,I278668,I278699,I278744,I278761,I278792,I278809,I278873,I278890,I307616,I307634,I278907,I278924,I307619,I278941,I278958,I307628,I278975,I278992,I307640,I279023,I279040,I279057,I307637,I279074,I307643,I279091,I279108,I279125,I279156,I279173,I279218,I279235,I307622,I279252,I307625,I279269,I279286,I279303,I279334,I307646,I279351,I279368,I307631,I279385,I279402,I279433,I279464,I279509,I279526,I279557,I279574,I279638,I279655,I315657,I315675,I279672,I279689,I315660,I279706,I279723,I315669,I279740,I279757,I315681,I279788,I279805,I279822,I315678,I279839,I315684,I279856,I279873,I279890,I279921,I279938,I279983,I280000,I315663,I280017,I315666,I280034,I280051,I280068,I280099,I315687,I280116,I280133,I315672,I280150,I280167,I280198,I280229,I280274,I280291,I280322,I280339,I280403,I280420,I349014,I349011,I280437,I280454,I349020,I280471,I280488,I349032,I280505,I280522,I349029,I280553,I280570,I280587,I349035,I280604,I349023,I280621,I280638,I280655,I280686,I280703,I280748,I280765,I280782,I349017,I280799,I280816,I280833,I280864,I349026,I280881,I280898,I280915,I280932,I280963,I280994,I281039,I281056,I281087,I281104,I281168,I281185,I422696,I422693,I281202,I281219,I422681,I281236,I281253,I422702,I281270,I281287,I422672,I281318,I281335,I281352,I422690,I281369,I422705,I422687,I281386,I281403,I281420,I281451,I281468,I281513,I281530,I422699,I281547,I422678,I281564,I281581,I281598,I281629,I422684,I281646,I422675,I281663,I281680,I281697,I281728,I281759,I281804,I281821,I281852,I281869,I281933,I281950,I281967,I281984,I282001,I282018,I282035,I282052,I282083,I282100,I282117,I282134,I282151,I282168,I282185,I282216,I282233,I282278,I282295,I282312,I282329,I282346,I282363,I282394,I282411,I282428,I282445,I282462,I282493,I282524,I282569,I282586,I282617,I282634,I282698,I282715,I282732,I282749,I282766,I282783,I282800,I282817,I282848,I282865,I282882,I282899,I282916,I282933,I282950,I282981,I282998,I283043,I283060,I283077,I283094,I283111,I283128,I283159,I283176,I283193,I283210,I283227,I283258,I283289,I283334,I283351,I283382,I283399,I283463,I283480,I424787,I424784,I283497,I283514,I424772,I283531,I283548,I424793,I283565,I283582,I424763,I283613,I283630,I283647,I424781,I283664,I424796,I424778,I283681,I283698,I283715,I283746,I283763,I283808,I283825,I424790,I283842,I424769,I283859,I283876,I283893,I283924,I424775,I283941,I424766,I283958,I283975,I283992,I284023,I284054,I284099,I284116,I284147,I284164,I284228,I284245,I284262,I284279,I284296,I284313,I284330,I284347,I284190,I284378,I284395,I284412,I284429,I284446,I284463,I284480,I284205,I284511,I284528,I284193,I284208,I284573,I284590,I284607,I284624,I284641,I284658,I284199,I284689,I284706,I284723,I284740,I284757,I284220,I284788,I284196,I284819,I284217,I284211,I284864,I284881,I284202,I284912,I284929,I284214,I284993,I285010,I285027,I285044,I285061,I285078,I285095,I285112,I285129,I285146,I285163,I285180,I285197,I285214,I285231,I285248,I285293,I285310,I285327,I285358,I285375,I285392,I285409,I285454,I285485,I285502,I285519,I285550,I285567,I285598,I285629,I285660,I285724,I285741,I401303,I401318,I285758,I285775,I401309,I285792,I285809,I285826,I401306,I285843,I401327,I285860,I401324,I285877,I285894,I285911,I401321,I401315,I285928,I401312,I285945,I285962,I285979,I286024,I286041,I286058,I286089,I286106,I286123,I286140,I286185,I286216,I286233,I286250,I286281,I286298,I286329,I286360,I286391,I286455,I286472,I357960,I357945,I286489,I286506,I286523,I286540,I357939,I286557,I357942,I286574,I357936,I286591,I357951,I286608,I286625,I286642,I357948,I286659,I286676,I286693,I286710,I286435,I286429,I286755,I286772,I286789,I286432,I286820,I357954,I286837,I357957,I286854,I286871,I286417,I286420,I286916,I286423,I286947,I286964,I286981,I286441,I287012,I287029,I286447,I287060,I286444,I287091,I286426,I287122,I286438,I287186,I287203,I287220,I287237,I287254,I287271,I287288,I287305,I287322,I287339,I287356,I287373,I287390,I287407,I287424,I287441,I287486,I287503,I287520,I287551,I287568,I287585,I287602,I287647,I287678,I287695,I287712,I287743,I287760,I287791,I287822,I287853,I287917,I287934,I287951,I287968,I287985,I288002,I288019,I288036,I288053,I288070,I288087,I288104,I288121,I288138,I288155,I288172,I287897,I287891,I288217,I288234,I288251,I287894,I288282,I288299,I288316,I288333,I287879,I287882,I288378,I287885,I288409,I288426,I288443,I287903,I288474,I288491,I287909,I288522,I287906,I288553,I287888,I288584,I287900,I288648,I288665,I288682,I288699,I288716,I288733,I288750,I288767,I288784,I288801,I288818,I288835,I288852,I288869,I288886,I288903,I288948,I288965,I288982,I289013,I289030,I289047,I289064,I289109,I289140,I289157,I289174,I289205,I289222,I289253,I289284,I289315,I289379,I289396,I289413,I289430,I289447,I289464,I289481,I289498,I289515,I289532,I289549,I289566,I289583,I289600,I289617,I289634,I289679,I289696,I289713,I289744,I289761,I289778,I289795,I289840,I289871,I289888,I289905,I289936,I289953,I289984,I290015,I290046,I290110,I290127,I290144,I290161,I290178,I290195,I290212,I290229,I290246,I290263,I290280,I290297,I290314,I290331,I290348,I290365,I290090,I290084,I290410,I290427,I290444,I290087,I290475,I290492,I290509,I290526,I290072,I290075,I290571,I290078,I290602,I290619,I290636,I290096,I290667,I290684,I290102,I290715,I290099,I290746,I290081,I290777,I290093,I290841,I290858,I290875,I290892,I290909,I290926,I290943,I290960,I290977,I290994,I291011,I291028,I291045,I291062,I291079,I291096,I290821,I290815,I291141,I291158,I291175,I290818,I291206,I291223,I291240,I291257,I290803,I290806,I291302,I290809,I291333,I291350,I291367,I290827,I291398,I291415,I290833,I291446,I290830,I291477,I290812,I291508,I290824,I291572,I291589,I373868,I373874,I291606,I291623,I373898,I291640,I291657,I373865,I291674,I373871,I291691,I373880,I291708,I373895,I291725,I291742,I291759,I373886,I373883,I291776,I291793,I291810,I291827,I291872,I291889,I291906,I291937,I373877,I373889,I291954,I291971,I291988,I292033,I292064,I373892,I292081,I292098,I292129,I292146,I292177,I292208,I292239,I292303,I292320,I292337,I292354,I292371,I292388,I292405,I292422,I292439,I292456,I292473,I292490,I292507,I292524,I292541,I292558,I292283,I292277,I292603,I292620,I292637,I292280,I292668,I292685,I292702,I292719,I292265,I292268,I292764,I292271,I292795,I292812,I292829,I292289,I292860,I292877,I292295,I292908,I292292,I292939,I292274,I292970,I292286,I293034,I293051,I419884,I419890,I293068,I293085,I293102,I293119,I419905,I293136,I419917,I293153,I419887,I419899,I293170,I419908,I293187,I293204,I293221,I419914,I419896,I293238,I293255,I293272,I293289,I293014,I293008,I293334,I293351,I293368,I293011,I293399,I419902,I419911,I293416,I419893,I293433,I293450,I292996,I292999,I293495,I293002,I293526,I293543,I293560,I293020,I293591,I293608,I293026,I293639,I293023,I293670,I293005,I293701,I293017,I293765,I293782,I293799,I293816,I293833,I293850,I293867,I293884,I293901,I293918,I293935,I293952,I293969,I293986,I294003,I294020,I294065,I294082,I294099,I294130,I294147,I294164,I294181,I294226,I294257,I294274,I294291,I294322,I294339,I294370,I294401,I294432,I294496,I294513,I294530,I294547,I294564,I294581,I294598,I294615,I294632,I294649,I294666,I294683,I294700,I294717,I294734,I294751,I294796,I294813,I294830,I294861,I294878,I294895,I294912,I294957,I294988,I295005,I295022,I295053,I295070,I295101,I295132,I295163,I295227,I295244,I295261,I295278,I295295,I295312,I295329,I295346,I295363,I295380,I295397,I295414,I295431,I295448,I295465,I295482,I295207,I295201,I295527,I295544,I295561,I295204,I295592,I295609,I295626,I295643,I295189,I295192,I295688,I295195,I295719,I295736,I295753,I295213,I295784,I295801,I295219,I295832,I295216,I295863,I295198,I295894,I295210,I295958,I295975,I295992,I296009,I296026,I296043,I296060,I296077,I296094,I296111,I296128,I296145,I296162,I296179,I296196,I296213,I296258,I296275,I296292,I296323,I296340,I296357,I296374,I296419,I296450,I296467,I296484,I296515,I296532,I296563,I296594,I296625,I296689,I296706,I296723,I296740,I296757,I296774,I296791,I296808,I296825,I296842,I296859,I296876,I296893,I296910,I296927,I296944,I296669,I296663,I296989,I297006,I297023,I296666,I297054,I297071,I297088,I297105,I296651,I296654,I297150,I296657,I297181,I297198,I297215,I296675,I297246,I297263,I296681,I297294,I296678,I297325,I296660,I297356,I296672,I297420,I297437,I297454,I297471,I297488,I297505,I297522,I297539,I297556,I297573,I297590,I297607,I297624,I297641,I297658,I297675,I297400,I297394,I297720,I297737,I297754,I297397,I297785,I297802,I297819,I297836,I297382,I297385,I297881,I297388,I297912,I297929,I297946,I297406,I297977,I297994,I297412,I298025,I297409,I298056,I297391,I298087,I297403,I298151,I298168,I298185,I298202,I298219,I298236,I298253,I298270,I298287,I298304,I298321,I298338,I298355,I298372,I298389,I298406,I298451,I298468,I298485,I298516,I298533,I298550,I298567,I298612,I298643,I298660,I298677,I298708,I298725,I298756,I298787,I298818,I298882,I298899,I298916,I298933,I298950,I298967,I298984,I299001,I299018,I299035,I299052,I299069,I299086,I299103,I299120,I299137,I299182,I299199,I299216,I299247,I299264,I299281,I299298,I299343,I299374,I299391,I299408,I299439,I299456,I299487,I299518,I299549,I299613,I299630,I299647,I299664,I299681,I299698,I299715,I299732,I299749,I299766,I299783,I299800,I299817,I299834,I299851,I299868,I299593,I299587,I299913,I299930,I299947,I299590,I299978,I299995,I300012,I300029,I299575,I299578,I300074,I299581,I300105,I300122,I300139,I299599,I300170,I300187,I299605,I300218,I299602,I300249,I299584,I300280,I299596,I300344,I300361,I325830,I325815,I300378,I300395,I300412,I300429,I325809,I300446,I325812,I300463,I325806,I300480,I325821,I300497,I300514,I300531,I325818,I300548,I300565,I300582,I300599,I300644,I300661,I300678,I300709,I325824,I300726,I325827,I300743,I300760,I300805,I300836,I300853,I300870,I300901,I300918,I300949,I300980,I301011,I301075,I301092,I301109,I301126,I301143,I301160,I301177,I301194,I301211,I301228,I301245,I301262,I301279,I301296,I301313,I301330,I301055,I301049,I301375,I301392,I301409,I301052,I301440,I301457,I301474,I301491,I301037,I301040,I301536,I301043,I301567,I301584,I301601,I301061,I301632,I301649,I301067,I301680,I301064,I301711,I301046,I301742,I301058,I301806,I301823,I301840,I301857,I301874,I301891,I301908,I301925,I301942,I301959,I301976,I301993,I302010,I302027,I302044,I302061,I302106,I302123,I302140,I302171,I302188,I302205,I302222,I302267,I302298,I302315,I302332,I302363,I302380,I302411,I302442,I302473,I302537,I302554,I390664,I390670,I302571,I302588,I390694,I302605,I302622,I390661,I302639,I390667,I302656,I390676,I302673,I390691,I302690,I302707,I302724,I390682,I390679,I302741,I302758,I302775,I302792,I302517,I302511,I302837,I302854,I302871,I302514,I302902,I390673,I390685,I302919,I302936,I302953,I302499,I302502,I302998,I302505,I303029,I390688,I303046,I303063,I302523,I303094,I303111,I302529,I303142,I302526,I303173,I302508,I303204,I302520,I303268,I303285,I386142,I386148,I303302,I303319,I386172,I303336,I303353,I386139,I303370,I386145,I303387,I386154,I303404,I386169,I303421,I303438,I303455,I386160,I386157,I303472,I303489,I303506,I303523,I303248,I303242,I303568,I303585,I303602,I303245,I303633,I386151,I386163,I303650,I303667,I303684,I303230,I303233,I303729,I303236,I303760,I386166,I303777,I303794,I303254,I303825,I303842,I303260,I303873,I303257,I303904,I303239,I303935,I303251,I303999,I304016,I444976,I444982,I304033,I304050,I304067,I304084,I444997,I304101,I445009,I304118,I444979,I444991,I304135,I445000,I304152,I304169,I304186,I445006,I444988,I304203,I304220,I304237,I304254,I303979,I303973,I304299,I304316,I304333,I303976,I304364,I444994,I445003,I304381,I444985,I304398,I304415,I303961,I303964,I304460,I303967,I304491,I304508,I304525,I303985,I304556,I304573,I303991,I304604,I303988,I304635,I303970,I304666,I303982,I304730,I304747,I442885,I442891,I304764,I304781,I304798,I304815,I442906,I304832,I442918,I304849,I442888,I442900,I304866,I442909,I304883,I304900,I304917,I442915,I442897,I304934,I304951,I304968,I304985,I305030,I305047,I305064,I305095,I442903,I442912,I305112,I442894,I305129,I305146,I305191,I305222,I305239,I305256,I305287,I305304,I305335,I305366,I305397,I305461,I305478,I305495,I305512,I305529,I305546,I305563,I305580,I305597,I305614,I305631,I305648,I305665,I305682,I305699,I305716,I305441,I305435,I305761,I305778,I305795,I305438,I305826,I305843,I305860,I305877,I305423,I305426,I305922,I305429,I305953,I305970,I305987,I305447,I306018,I306035,I305453,I306066,I305450,I306097,I305432,I306128,I305444,I306192,I306209,I306226,I306243,I306260,I306277,I306294,I306311,I306328,I306345,I306362,I306379,I306396,I306413,I306430,I306447,I306492,I306509,I306526,I306557,I306574,I306591,I306608,I306653,I306684,I306701,I306718,I306749,I306766,I306797,I306828,I306859,I306923,I306940,I386788,I386794,I306957,I306974,I386818,I306991,I307008,I386785,I307025,I386791,I307042,I386800,I307059,I386815,I307076,I307093,I307110,I386806,I386803,I307127,I307144,I307161,I307178,I307223,I307240,I307257,I307288,I386797,I386809,I307305,I307322,I307339,I307384,I307415,I386812,I307432,I307449,I307480,I307497,I307528,I307559,I307590,I307654,I307671,I307688,I307705,I307722,I307739,I307756,I307773,I307790,I307807,I307824,I307841,I307858,I307875,I307892,I307909,I307954,I307971,I307988,I308019,I308036,I308053,I308070,I308115,I308146,I308163,I308180,I308211,I308228,I308259,I308290,I308321,I308385,I308402,I354390,I354375,I308419,I308436,I308453,I308470,I354369,I308487,I354372,I308504,I354366,I308521,I354381,I308538,I308555,I308572,I354378,I308589,I308606,I308623,I308640,I308685,I308702,I308719,I308750,I354384,I308767,I354387,I308784,I308801,I308846,I308877,I308894,I308911,I308942,I308959,I308990,I309021,I309052,I309116,I309133,I309150,I309167,I309184,I309201,I309218,I309235,I309252,I309269,I309286,I309303,I309320,I309337,I309354,I309371,I309416,I309433,I309450,I309481,I309498,I309515,I309532,I309577,I309608,I309625,I309642,I309673,I309690,I309721,I309752,I309783,I309847,I309864,I309881,I309898,I309915,I309932,I309949,I309966,I309983,I310000,I310017,I310034,I310051,I310068,I310085,I310102,I309827,I309821,I310147,I310164,I310181,I309824,I310212,I310229,I310246,I310263,I309809,I309812,I310308,I309815,I310339,I310356,I310373,I309833,I310404,I310421,I309839,I310452,I309836,I310483,I309818,I310514,I309830,I310578,I310595,I310612,I310629,I310646,I310663,I310680,I310697,I310714,I310731,I310748,I310765,I310782,I310799,I310816,I310833,I310878,I310895,I310912,I310943,I310960,I310977,I310994,I311039,I311070,I311087,I311104,I311135,I311152,I311183,I311214,I311245,I311309,I311326,I311343,I311360,I311377,I311394,I311411,I311428,I311445,I311462,I311479,I311496,I311513,I311530,I311547,I311564,I311609,I311626,I311643,I311674,I311691,I311708,I311725,I311770,I311801,I311818,I311835,I311866,I311883,I311914,I311945,I311976,I312040,I312057,I408103,I408118,I312074,I312091,I408109,I312108,I312125,I312142,I408106,I312159,I408127,I312176,I408124,I312193,I312210,I312227,I408121,I408115,I312244,I408112,I312261,I312278,I312295,I312340,I312357,I312374,I312405,I312422,I312439,I312456,I312501,I312532,I312549,I312566,I312597,I312614,I312645,I312676,I312707,I312771,I312788,I412217,I412223,I312805,I312822,I312839,I312856,I412238,I312873,I412250,I312890,I412220,I412232,I312907,I412241,I312924,I312941,I312958,I412247,I412229,I312975,I312992,I313009,I313026,I312751,I312745,I313071,I313088,I313105,I312748,I313136,I412235,I412244,I313153,I412226,I313170,I313187,I312733,I312736,I313232,I312739,I313263,I313280,I313297,I312757,I313328,I313345,I312763,I313376,I312760,I313407,I312742,I313438,I312754,I313502,I313519,I313536,I313553,I313570,I313587,I313604,I313621,I313638,I313655,I313672,I313689,I313706,I313723,I313740,I313757,I313802,I313819,I313836,I313867,I313884,I313901,I313918,I313963,I313994,I314011,I314028,I314059,I314076,I314107,I314138,I314169,I314233,I314250,I314267,I314284,I314301,I314318,I314335,I314352,I314369,I314386,I314403,I314420,I314437,I314454,I314471,I314488,I314533,I314550,I314567,I314598,I314615,I314632,I314649,I314694,I314725,I314742,I314759,I314790,I314807,I314838,I314869,I314900,I314964,I314981,I387434,I387440,I314998,I315015,I387464,I315032,I315049,I387431,I315066,I387437,I315083,I387446,I315100,I387461,I315117,I315134,I315151,I387452,I387449,I315168,I315185,I315202,I315219,I315264,I315281,I315298,I315329,I387443,I387455,I315346,I315363,I315380,I315425,I315456,I387458,I315473,I315490,I315521,I315538,I315569,I315600,I315631,I315695,I315712,I377098,I377104,I315729,I315746,I377128,I315763,I315780,I377095,I315797,I377101,I315814,I377110,I315831,I377125,I315848,I315865,I315882,I377116,I377113,I315899,I315916,I315933,I315950,I315995,I316012,I316029,I316060,I377107,I377119,I316077,I316094,I316111,I316156,I316187,I377122,I316204,I316221,I316252,I316269,I316300,I316331,I316362,I316426,I316443,I316460,I316477,I316494,I316511,I316528,I316545,I316562,I316579,I316596,I316613,I316630,I316647,I316664,I316681,I316726,I316743,I316760,I316791,I316808,I316825,I316842,I316887,I316918,I316935,I316952,I316983,I317000,I317031,I317062,I317093,I317157,I317174,I317191,I317208,I317225,I317242,I317259,I317276,I317293,I317310,I317327,I317344,I317361,I317378,I317395,I317412,I317457,I317474,I317491,I317522,I317539,I317556,I317573,I317618,I317649,I317666,I317683,I317714,I317731,I317762,I317793,I317824,I317888,I317905,I317922,I317939,I317956,I317973,I317990,I318007,I318024,I318041,I318058,I318075,I318092,I318109,I318126,I318143,I318188,I318205,I318222,I318253,I318270,I318287,I318304,I318349,I318380,I318397,I318414,I318445,I318462,I318493,I318524,I318555,I318619,I318636,I418490,I418496,I318653,I318670,I318687,I318704,I418511,I318721,I418523,I318738,I418493,I418505,I318755,I418514,I318772,I318789,I318806,I418520,I418502,I318823,I318840,I318857,I318874,I318919,I318936,I318953,I318984,I418508,I418517,I319001,I418499,I319018,I319035,I319080,I319111,I319128,I319145,I319176,I319193,I319224,I319255,I319286,I319350,I319367,I431733,I431739,I319384,I319401,I319418,I319435,I431754,I319452,I431766,I319469,I431736,I431748,I319486,I431757,I319503,I319520,I319537,I431763,I431745,I319554,I319571,I319588,I319605,I319650,I319667,I319684,I319715,I431751,I431760,I319732,I431742,I319749,I319766,I319811,I319842,I319859,I319876,I319907,I319924,I319955,I319986,I320017,I320081,I320098,I320115,I320132,I320149,I320166,I320183,I320200,I320217,I320234,I320251,I320268,I320285,I320302,I320319,I320336,I320381,I320398,I320415,I320446,I320463,I320480,I320497,I320542,I320573,I320590,I320607,I320638,I320655,I320686,I320717,I320748,I320812,I320829,I320846,I320863,I320880,I320897,I320914,I320931,I320948,I320965,I320982,I320999,I321016,I321033,I321050,I321067,I320792,I320786,I321112,I321129,I321146,I320789,I321177,I321194,I321211,I321228,I320774,I320777,I321273,I320780,I321304,I321321,I321338,I320798,I321369,I321386,I320804,I321417,I320801,I321448,I320783,I321479,I320795,I321543,I321560,I321577,I321594,I321611,I321628,I321645,I321662,I321679,I321696,I321713,I321730,I321747,I321764,I321781,I321798,I321843,I321860,I321877,I321908,I321925,I321942,I321959,I322004,I322035,I322052,I322069,I322100,I322117,I322148,I322179,I322210,I322268,I322285,I322302,I322319,I322336,I322353,I322370,I322387,I322404,I322421,I322438,I322469,I322486,I322503,I322520,I322537,I322554,I322571,I322616,I322647,I322664,I322695,I322712,I322743,I322788,I322805,I322863,I322880,I322897,I322914,I322931,I322948,I322965,I322982,I322999,I323016,I323033,I323064,I323081,I323098,I323115,I323132,I323149,I323166,I323211,I323242,I323259,I323290,I323307,I323338,I323383,I323400,I323458,I323475,I323492,I323509,I323526,I323543,I323560,I323577,I323594,I323611,I323628,I323659,I323676,I323693,I323710,I323727,I323744,I323761,I323806,I323837,I323854,I323885,I323902,I323933,I323978,I323995,I324053,I324070,I324087,I324104,I324121,I324138,I324155,I324172,I324189,I324206,I324223,I324254,I324271,I324288,I324305,I324322,I324339,I324356,I324401,I324432,I324449,I324480,I324497,I324528,I324573,I324590,I324648,I324665,I324682,I324699,I324716,I324733,I324750,I324767,I324784,I324801,I324818,I324849,I324866,I324883,I324900,I324917,I324934,I324951,I324996,I325027,I325044,I325075,I325092,I325123,I325168,I325185,I325243,I325260,I325277,I325294,I325311,I325328,I325345,I325362,I325379,I325396,I325413,I325232,I325444,I325461,I325478,I325495,I325512,I325529,I325546,I325217,I325214,I325591,I325235,I325622,I325639,I325211,I325670,I325687,I325220,I325718,I325229,I325226,I325763,I325780,I325223,I325838,I325855,I325872,I325889,I325906,I325923,I325940,I325957,I325974,I325991,I326008,I326039,I326056,I326073,I326090,I326107,I326124,I326141,I326186,I326217,I326234,I326265,I326282,I326313,I326358,I326375,I326433,I326450,I402004,I402001,I326467,I401992,I401989,I326484,I326501,I326518,I401986,I401998,I326535,I326552,I326569,I326586,I326603,I326634,I326651,I326668,I326685,I326702,I401983,I326719,I326736,I326781,I326812,I401995,I402007,I326829,I326860,I326877,I326908,I326953,I326970,I327028,I327045,I327062,I327079,I327096,I327113,I327130,I327147,I327164,I327181,I327198,I327229,I327246,I327263,I327280,I327297,I327314,I327331,I327376,I327407,I327424,I327455,I327472,I327503,I327548,I327565,I327623,I327640,I327657,I327674,I327691,I327708,I327725,I327742,I327759,I327776,I327793,I327612,I327824,I327841,I327858,I327875,I327892,I327909,I327926,I327597,I327594,I327971,I327615,I328002,I328019,I327591,I328050,I328067,I327600,I328098,I327609,I327606,I328143,I328160,I327603,I328218,I328235,I328252,I328269,I328286,I328303,I328320,I328337,I328354,I328371,I328388,I328419,I328436,I328453,I328470,I328487,I328504,I328521,I328566,I328597,I328614,I328645,I328662,I328693,I328738,I328755,I328813,I328830,I388107,I388104,I328847,I388089,I388083,I328864,I328881,I328898,I388110,I388077,I328915,I328932,I328949,I328966,I328983,I329014,I388101,I388092,I329031,I388095,I329048,I329065,I329082,I388098,I388080,I329099,I329116,I329161,I329192,I329209,I329240,I388086,I329257,I329288,I329333,I329350,I329408,I329425,I429648,I429645,I329442,I429651,I429669,I329459,I329476,I329493,I429660,I429654,I329510,I429675,I329527,I329544,I329561,I329578,I329397,I329609,I429642,I429666,I329626,I429672,I329643,I329660,I329677,I329694,I329711,I329382,I329379,I329756,I329400,I329787,I429657,I329804,I329376,I329835,I429663,I329852,I329385,I329883,I329394,I329391,I329928,I329945,I329388,I330003,I330020,I330037,I330054,I330071,I330088,I330105,I330122,I330139,I330156,I330173,I330204,I330221,I330238,I330255,I330272,I330289,I330306,I330351,I330382,I330399,I330430,I330447,I330478,I330523,I330540,I330598,I330615,I330632,I330649,I330666,I330683,I330700,I330717,I330734,I330751,I330768,I330799,I330816,I330833,I330850,I330867,I330884,I330901,I330946,I330977,I330994,I331025,I331042,I331073,I331118,I331135,I331193,I331210,I331227,I331244,I331261,I331278,I331295,I331312,I331329,I331346,I331363,I331394,I331411,I331428,I331445,I331462,I331479,I331496,I331541,I331572,I331589,I331620,I331637,I331668,I331713,I331730,I331788,I331805,I331822,I331839,I331856,I331873,I331890,I331907,I331924,I331941,I331958,I331777,I331989,I332006,I332023,I332040,I332057,I332074,I332091,I331762,I331759,I332136,I331780,I332167,I332184,I331756,I332215,I332232,I331765,I332263,I331774,I331771,I332308,I332325,I331768,I332383,I332400,I332417,I332434,I332451,I332468,I332485,I332502,I332519,I332536,I332553,I332584,I332601,I332618,I332635,I332652,I332669,I332686,I332731,I332762,I332779,I332810,I332827,I332858,I332903,I332920,I332978,I332995,I333012,I333029,I333046,I333063,I333080,I333097,I333114,I333131,I333148,I333179,I333196,I333213,I333230,I333247,I333264,I333281,I333326,I333357,I333374,I333405,I333422,I333453,I333498,I333515,I333573,I333590,I399284,I399281,I333607,I399272,I399269,I333624,I333641,I333658,I399266,I399278,I333675,I333692,I333709,I333726,I333743,I333562,I333774,I333791,I333808,I333825,I333842,I399263,I333859,I333876,I333547,I333544,I333921,I333565,I333952,I399275,I399287,I333969,I333541,I334000,I334017,I333550,I334048,I333559,I333556,I334093,I334110,I333553,I334168,I334185,I334202,I334219,I334236,I334253,I334270,I334287,I334304,I334321,I334338,I334369,I334386,I334403,I334420,I334437,I334454,I334471,I334516,I334547,I334564,I334595,I334612,I334643,I334688,I334705,I334763,I334780,I365688,I365691,I334797,I365703,I365709,I334814,I334831,I334848,I365694,I334865,I334882,I334899,I334916,I334933,I334752,I334964,I365712,I365706,I334981,I365721,I334998,I335015,I335032,I365715,I365697,I335049,I335066,I334737,I334734,I335111,I334755,I335142,I365718,I335159,I334731,I335190,I365700,I335207,I334740,I335238,I334749,I334746,I335283,I335300,I334743,I335358,I335375,I335392,I335409,I335426,I335443,I335460,I335477,I335494,I335511,I335528,I335559,I335576,I335593,I335610,I335627,I335644,I335661,I335706,I335737,I335754,I335785,I335802,I335833,I335878,I335895,I335953,I335970,I335987,I336004,I336021,I336038,I336055,I336072,I336089,I336106,I336123,I335942,I336154,I336171,I336188,I336205,I336222,I336239,I336256,I335927,I335924,I336301,I335945,I336332,I336349,I335921,I336380,I336397,I335930,I336428,I335939,I335936,I336473,I336490,I335933,I336548,I336565,I336582,I336599,I336616,I336633,I336650,I336667,I336684,I336701,I336718,I336537,I336749,I336766,I336783,I336800,I336817,I336834,I336851,I336522,I336519,I336896,I336540,I336927,I336944,I336516,I336975,I336992,I336525,I337023,I336534,I336531,I337068,I337085,I336528,I337143,I337160,I337177,I337194,I337211,I337228,I337245,I337262,I337279,I337296,I337313,I337132,I337344,I337361,I337378,I337395,I337412,I337429,I337446,I337117,I337114,I337491,I337135,I337522,I337539,I337111,I337570,I337587,I337120,I337618,I337129,I337126,I337663,I337680,I337123,I337738,I337755,I426163,I426160,I337772,I426166,I426184,I337789,I337806,I337823,I426175,I426169,I337840,I426190,I337857,I337874,I337891,I337908,I337727,I337939,I426157,I426181,I337956,I426187,I337973,I337990,I338007,I338024,I338041,I337712,I337709,I338086,I337730,I338117,I426172,I338134,I337706,I338165,I426178,I338182,I337715,I338213,I337724,I337721,I338258,I338275,I337718,I338333,I338350,I439406,I439403,I338367,I439409,I439427,I338384,I338401,I338418,I439418,I439412,I338435,I439433,I338452,I338469,I338486,I338503,I338534,I439400,I439424,I338551,I439430,I338568,I338585,I338602,I338619,I338636,I338681,I338712,I439415,I338729,I338760,I439421,I338777,I338808,I338853,I338870,I338928,I338945,I338962,I338979,I338996,I339013,I339030,I339047,I339064,I339081,I339098,I338917,I339129,I339146,I339163,I339180,I339197,I339214,I339231,I338902,I338899,I339276,I338920,I339307,I339324,I338896,I339355,I339372,I338905,I339403,I338914,I338911,I339448,I339465,I338908,I339523,I339540,I339557,I339574,I339591,I339608,I339625,I339642,I339659,I339676,I339693,I339724,I339741,I339758,I339775,I339792,I339809,I339826,I339871,I339902,I339919,I339950,I339967,I339998,I340043,I340060,I340118,I340135,I440800,I440797,I340152,I440803,I440821,I340169,I340186,I340203,I440812,I440806,I340220,I440827,I340237,I340254,I340271,I340288,I340107,I340319,I440794,I440818,I340336,I440824,I340353,I340370,I340387,I340404,I340421,I340092,I340089,I340466,I340110,I340497,I440809,I340514,I340086,I340545,I440815,I340562,I340095,I340593,I340104,I340101,I340638,I340655,I340098,I340713,I340730,I340747,I340764,I340781,I340798,I340815,I340832,I340849,I340866,I340883,I340914,I340931,I340948,I340965,I340982,I340999,I341016,I341061,I341092,I341109,I341140,I341157,I341188,I341233,I341250,I341308,I341325,I341342,I341359,I341376,I341393,I341410,I341427,I341444,I341461,I341478,I341509,I341526,I341543,I341560,I341577,I341594,I341611,I341656,I341687,I341704,I341735,I341752,I341783,I341828,I341845,I341903,I341920,I341937,I341954,I341971,I341988,I342005,I342022,I342039,I342056,I342073,I341892,I342104,I342121,I342138,I342155,I342172,I342189,I342206,I341877,I341874,I342251,I341895,I342282,I342299,I341871,I342330,I342347,I341880,I342378,I341889,I341886,I342423,I342440,I341883,I342498,I342515,I342532,I342549,I342566,I342583,I342600,I342617,I342634,I342651,I342668,I342487,I342699,I342716,I342733,I342750,I342767,I342784,I342801,I342472,I342469,I342846,I342490,I342877,I342894,I342466,I342925,I342942,I342475,I342973,I342484,I342481,I343018,I343035,I342478,I343093,I343110,I343127,I343144,I343161,I343178,I343195,I343212,I343229,I343246,I343263,I343294,I343311,I343328,I343345,I343362,I343379,I343396,I343441,I343472,I343489,I343520,I343537,I343568,I343613,I343630,I343688,I343705,I343722,I343739,I343756,I343773,I343790,I343807,I343824,I343841,I343858,I343889,I343906,I343923,I343940,I343957,I343974,I343991,I344036,I344067,I344084,I344115,I344132,I344163,I344208,I344225,I344283,I344300,I344317,I344334,I344351,I344368,I344385,I344402,I344419,I344436,I344453,I344484,I344501,I344518,I344535,I344552,I344569,I344586,I344631,I344662,I344679,I344710,I344727,I344758,I344803,I344820,I344878,I344895,I344912,I344929,I344946,I344963,I344980,I344997,I345014,I345031,I345048,I345079,I345096,I345113,I345130,I345147,I345164,I345181,I345226,I345257,I345274,I345305,I345322,I345353,I345398,I345415,I345473,I345490,I345507,I345524,I345541,I345558,I345575,I345592,I345609,I345626,I345643,I345674,I345691,I345708,I345725,I345742,I345759,I345776,I345821,I345852,I345869,I345900,I345917,I345948,I345993,I346010,I346068,I346085,I346102,I346119,I346136,I346153,I346170,I346187,I346204,I346221,I346238,I346057,I346269,I346286,I346303,I346320,I346337,I346354,I346371,I346042,I346039,I346416,I346060,I346447,I346464,I346036,I346495,I346512,I346045,I346543,I346054,I346051,I346588,I346605,I346048,I346663,I346680,I346697,I346714,I346731,I346748,I346765,I346782,I346799,I346816,I346833,I346864,I346881,I346898,I346915,I346932,I346949,I346966,I347011,I347042,I347059,I347090,I347107,I347138,I347183,I347200,I347258,I347275,I347292,I347309,I347326,I347343,I347360,I347377,I347394,I347411,I347428,I347459,I347476,I347493,I347510,I347527,I347544,I347561,I347606,I347637,I347654,I347685,I347702,I347733,I347778,I347795,I347853,I347870,I347887,I347904,I347921,I347938,I347955,I347972,I347989,I348006,I348023,I347842,I348054,I348071,I348088,I348105,I348122,I348139,I348156,I347827,I347824,I348201,I347845,I348232,I348249,I347821,I348280,I348297,I347830,I348328,I347839,I347836,I348373,I348390,I347833,I348448,I348465,I348482,I348499,I348516,I348533,I348550,I348567,I348584,I348601,I348618,I348437,I348649,I348666,I348683,I348700,I348717,I348734,I348751,I348422,I348419,I348796,I348440,I348827,I348844,I348416,I348875,I348892,I348425,I348923,I348434,I348431,I348968,I348985,I348428,I349043,I349060,I349077,I349094,I349111,I349128,I349145,I349162,I349179,I349196,I349213,I349244,I349261,I349278,I349295,I349312,I349329,I349346,I349391,I349422,I349439,I349470,I349487,I349518,I349563,I349580,I349638,I349655,I426860,I426857,I349672,I426863,I426881,I349689,I349706,I349723,I426872,I426866,I349740,I426887,I349757,I349774,I349791,I349808,I349839,I426854,I426878,I349856,I426884,I349873,I349890,I349907,I349924,I349941,I349986,I350017,I426869,I350034,I350065,I426875,I350082,I350113,I350158,I350175,I350233,I350250,I350267,I350284,I350301,I350318,I350335,I350352,I350369,I350386,I350403,I350434,I350451,I350468,I350485,I350502,I350519,I350536,I350581,I350612,I350629,I350660,I350677,I350708,I350753,I350770,I350828,I350845,I350862,I350879,I350896,I350913,I350930,I350947,I350964,I350981,I350998,I351029,I351046,I351063,I351080,I351097,I351114,I351131,I351176,I351207,I351224,I351255,I351272,I351303,I351348,I351365,I351423,I351440,I375187,I375184,I351457,I375169,I375163,I351474,I351491,I351508,I375190,I375157,I351525,I351542,I351559,I351576,I351593,I351624,I375181,I375172,I351641,I375175,I351658,I351675,I351692,I375178,I375160,I351709,I351726,I351771,I351802,I351819,I351850,I375166,I351867,I351898,I351943,I351960,I352018,I352035,I352052,I352069,I352086,I352103,I352120,I352137,I352154,I352171,I352188,I352007,I352219,I352236,I352253,I352270,I352287,I352304,I352321,I351992,I351989,I352366,I352010,I352397,I352414,I351986,I352445,I352462,I351995,I352493,I352004,I352001,I352538,I352555,I351998,I352613,I352630,I352647,I352664,I352681,I352698,I352715,I352732,I352749,I352766,I352783,I352602,I352814,I352831,I352848,I352865,I352882,I352899,I352916,I352587,I352584,I352961,I352605,I352992,I353009,I352581,I353040,I353057,I352590,I353088,I352599,I352596,I353133,I353150,I352593,I353208,I353225,I443588,I443585,I353242,I443591,I443609,I353259,I353276,I353293,I443600,I443594,I353310,I443615,I353327,I353344,I353361,I353378,I353409,I443582,I443606,I353426,I443612,I353443,I353460,I353477,I353494,I353511,I353556,I353587,I443597,I353604,I353635,I443603,I353652,I353683,I353728,I353745,I353803,I353820,I353837,I353854,I353871,I353888,I353905,I353922,I353939,I353956,I353973,I354004,I354021,I354038,I354055,I354072,I354089,I354106,I354151,I354182,I354199,I354230,I354247,I354278,I354323,I354340,I354398,I354415,I354432,I354449,I354466,I354483,I354500,I354517,I354534,I354551,I354568,I354599,I354616,I354633,I354650,I354667,I354684,I354701,I354746,I354777,I354794,I354825,I354842,I354873,I354918,I354935,I354993,I355010,I355027,I355044,I355061,I355078,I355095,I355112,I355129,I355146,I355163,I355194,I355211,I355228,I355245,I355262,I355279,I355296,I355341,I355372,I355389,I355420,I355437,I355468,I355513,I355530,I355588,I355605,I432436,I432433,I355622,I432439,I432457,I355639,I355656,I355673,I432448,I432442,I355690,I432463,I355707,I355724,I355741,I355758,I355577,I355789,I432430,I432454,I355806,I432460,I355823,I355840,I355857,I355874,I355891,I355562,I355559,I355936,I355580,I355967,I432445,I355984,I355556,I356015,I432451,I356032,I355565,I356063,I355574,I355571,I356108,I356125,I355568,I356183,I356200,I356217,I356234,I356251,I356268,I356285,I356302,I356319,I356336,I356353,I356384,I356401,I356418,I356435,I356452,I356469,I356486,I356531,I356562,I356579,I356610,I356627,I356658,I356703,I356720,I356778,I356795,I356812,I356829,I356846,I356863,I356880,I356897,I356914,I356931,I356948,I356767,I356979,I356996,I357013,I357030,I357047,I357064,I357081,I356752,I356749,I357126,I356770,I357157,I357174,I356746,I357205,I357222,I356755,I357253,I356764,I356761,I357298,I357315,I356758,I357373,I357390,I357407,I357424,I357441,I357458,I357475,I357492,I357509,I357526,I357543,I357574,I357591,I357608,I357625,I357642,I357659,I357676,I357721,I357752,I357769,I357800,I357817,I357848,I357893,I357910,I357968,I357985,I358002,I358019,I358036,I358053,I358070,I358087,I358104,I358121,I358138,I358169,I358186,I358203,I358220,I358237,I358254,I358271,I358316,I358347,I358364,I358395,I358412,I358443,I358488,I358505,I358563,I358580,I358597,I358614,I358631,I358648,I358665,I358682,I358699,I358716,I358733,I358764,I358781,I358798,I358815,I358832,I358849,I358866,I358911,I358942,I358959,I358990,I359007,I359038,I359083,I359100,I359158,I359175,I359192,I359209,I359226,I359243,I359260,I359277,I359294,I359311,I359328,I359359,I359376,I359393,I359410,I359427,I359444,I359461,I359506,I359537,I359554,I359585,I359602,I359633,I359678,I359695,I359753,I359770,I359787,I359804,I359821,I359838,I359855,I359872,I359889,I359906,I359923,I359742,I359954,I359971,I359988,I360005,I360022,I360039,I360056,I359727,I359724,I360101,I359745,I360132,I360149,I359721,I360180,I360197,I359730,I360228,I359739,I359736,I360273,I360290,I359733,I360348,I360365,I360382,I360399,I360416,I360433,I360450,I360467,I360484,I360501,I360518,I360549,I360566,I360583,I360600,I360617,I360634,I360651,I360696,I360727,I360744,I360775,I360792,I360823,I360868,I360885,I360943,I360960,I360977,I360994,I361011,I361028,I361045,I361062,I361079,I361096,I361113,I361144,I361161,I361178,I361195,I361212,I361229,I361246,I361291,I361322,I361339,I361370,I361387,I361418,I361463,I361480,I361538,I361555,I361572,I361589,I361606,I361623,I361640,I361657,I361674,I361691,I361708,I361739,I361756,I361773,I361790,I361807,I361824,I361841,I361886,I361917,I361934,I361965,I361982,I362013,I362058,I362075,I362133,I362150,I362167,I362184,I362201,I362218,I362235,I362252,I362269,I362286,I362303,I362334,I362351,I362368,I362385,I362402,I362419,I362436,I362481,I362512,I362529,I362560,I362577,I362608,I362653,I362670,I362728,I362745,I362762,I362779,I362796,I362813,I362830,I362847,I362864,I362881,I362898,I362929,I362946,I362963,I362980,I362997,I363014,I363031,I363076,I363107,I363124,I363155,I363172,I363203,I363248,I363265,I363332,I363349,I363366,I363383,I363400,I363417,I363434,I363451,I363468,I363485,I363502,I363533,I363550,I363567,I363598,I363615,I363632,I363649,I363680,I363711,I363737,I363745,I363762,I363779,I363796,I363827,I363844,I363861,I363892,I363909,I363954,I363999,I364016,I364033,I364064,I364131,I364148,I364165,I364182,I364199,I364216,I364233,I364250,I364267,I364284,I364301,I364093,I364332,I364349,I364366,I364105,I364397,I364414,I364431,I364448,I364111,I364479,I364102,I364510,I364536,I364544,I364561,I364578,I364595,I364120,I364626,I364643,I364660,I364090,I364691,I364708,I364108,I364123,I364753,I364096,I364117,I364798,I364815,I364832,I364099,I364863,I364114,I364930,I364947,I364964,I364981,I364998,I365015,I365032,I365049,I365066,I365083,I365100,I364892,I365131,I365148,I365165,I364904,I365196,I365213,I365230,I365247,I364910,I365278,I364901,I365309,I365335,I365343,I365360,I365377,I365394,I364919,I365425,I365442,I365459,I364889,I365490,I365507,I364907,I364922,I365552,I364895,I364916,I365597,I365614,I365631,I364898,I365662,I364913,I365729,I365746,I365763,I365780,I365797,I365814,I365831,I365848,I365865,I365882,I365899,I365930,I365947,I365964,I365995,I366012,I366029,I366046,I366077,I366108,I366134,I366142,I366159,I366176,I366193,I366224,I366241,I366258,I366289,I366306,I366351,I366396,I366413,I366430,I366461,I366528,I366545,I430369,I430351,I366562,I430366,I430360,I366579,I366596,I366613,I366630,I430345,I430372,I366647,I366664,I366681,I430342,I366698,I430363,I366729,I366746,I430354,I366763,I430357,I366794,I366811,I366828,I366845,I366876,I366907,I430348,I366933,I366941,I366958,I366975,I366992,I367023,I367040,I430339,I367057,I367088,I367105,I367150,I367195,I367212,I367229,I367260,I367327,I367344,I367361,I367378,I367395,I367412,I367429,I367446,I367463,I367480,I367497,I367528,I367545,I367562,I367593,I367610,I367627,I367644,I367675,I367706,I367732,I367740,I367757,I367774,I367791,I367822,I367839,I367856,I367887,I367904,I367949,I367994,I368011,I368028,I368059,I368126,I368143,I368160,I368177,I368194,I368211,I368228,I368245,I368262,I368279,I368296,I368327,I368344,I368361,I368392,I368409,I368426,I368443,I368474,I368505,I368531,I368539,I368556,I368573,I368590,I368621,I368638,I368655,I368686,I368703,I368748,I368793,I368810,I368827,I368858,I368925,I368942,I440127,I440109,I368959,I440124,I440118,I368976,I368993,I369010,I369027,I440103,I440130,I369044,I369061,I369078,I440100,I369095,I440121,I369126,I369143,I440112,I369160,I440115,I369191,I369208,I369225,I369242,I369273,I369304,I440106,I369330,I369338,I369355,I369372,I369389,I369420,I369437,I440097,I369454,I369485,I369502,I369547,I369592,I369609,I369626,I369657,I369724,I369741,I369758,I369775,I369792,I369809,I369826,I369843,I369860,I369877,I369894,I369925,I369942,I369959,I369990,I370007,I370024,I370041,I370072,I370103,I370129,I370137,I370154,I370171,I370188,I370219,I370236,I370253,I370284,I370301,I370346,I370391,I370408,I370425,I370456,I370523,I370540,I370557,I370574,I370591,I370608,I370625,I370642,I370659,I370676,I370693,I370724,I370741,I370758,I370789,I370806,I370823,I370840,I370871,I370902,I370928,I370936,I370953,I370970,I370987,I371018,I371035,I371052,I371083,I371100,I371145,I371190,I371207,I371224,I371255,I371322,I371339,I371356,I371373,I371390,I371407,I371424,I371441,I371467,I371475,I371492,I371509,I371293,I371540,I371557,I371574,I371281,I371305,I371619,I371636,I371653,I371670,I371687,I371287,I371718,I371735,I371290,I371299,I371308,I371296,I371808,I371825,I371284,I371856,I371314,I371311,I371901,I371302,I371968,I371985,I372002,I372019,I372036,I372053,I372070,I372087,I372113,I372121,I372138,I372155,I371939,I372186,I372203,I372220,I371927,I371951,I372265,I372282,I372299,I372316,I372333,I371933,I372364,I372381,I371936,I371945,I371954,I371942,I372454,I372471,I371930,I372502,I371960,I371957,I372547,I371948,I372614,I372631,I372648,I372665,I372682,I372699,I372716,I372733,I372759,I372767,I372784,I372801,I372832,I372849,I372866,I372911,I372928,I372945,I372962,I372979,I373010,I373027,I373100,I373117,I373148,I373193,I373260,I373277,I373294,I373311,I373328,I373345,I373362,I373379,I373405,I373413,I373430,I373447,I373478,I373495,I373512,I373557,I373574,I373591,I373608,I373625,I373656,I373673,I373746,I373763,I373794,I373839,I373906,I373923,I373940,I373957,I373974,I373991,I374008,I374025,I374051,I374059,I374076,I374093,I374124,I374141,I374158,I374203,I374220,I374237,I374254,I374271,I374302,I374319,I374392,I374409,I374440,I374485,I374552,I374569,I374586,I374603,I374620,I374637,I374654,I374671,I374697,I374705,I374722,I374739,I374523,I374770,I374787,I374804,I374511,I374535,I374849,I374866,I374883,I374900,I374917,I374517,I374948,I374965,I374520,I374529,I374538,I374526,I375038,I375055,I374514,I375086,I374544,I374541,I375131,I374532,I375198,I375215,I375232,I375249,I375266,I375283,I375300,I375317,I375343,I375351,I375368,I375385,I375416,I375433,I375450,I375495,I375512,I375529,I375546,I375563,I375594,I375611,I375684,I375701,I375732,I375777,I375844,I375861,I375878,I375895,I375912,I375929,I375946,I375963,I375989,I375997,I376014,I376031,I376062,I376079,I376096,I376141,I376158,I376175,I376192,I376209,I376240,I376257,I376330,I376347,I376378,I376423,I376490,I376507,I376524,I376541,I376558,I376575,I376592,I376609,I376635,I376643,I376660,I376677,I376708,I376725,I376742,I376787,I376804,I376821,I376838,I376855,I376886,I376903,I376976,I376993,I377024,I377069,I377136,I377153,I377170,I377187,I377204,I377221,I377238,I377255,I377281,I377289,I377306,I377323,I377354,I377371,I377388,I377433,I377450,I377467,I377484,I377501,I377532,I377549,I377622,I377639,I377670,I377715,I377782,I377799,I377816,I377833,I377850,I377867,I377884,I377901,I377927,I377935,I377952,I377969,I377753,I378000,I378017,I378034,I377741,I377765,I378079,I378096,I378113,I378130,I378147,I377747,I378178,I378195,I377750,I377759,I377768,I377756,I378268,I378285,I377744,I378316,I377774,I377771,I378361,I377762,I378428,I378445,I415735,I415708,I378462,I415705,I415723,I378479,I378496,I378513,I378530,I415726,I415711,I378547,I415729,I378573,I378581,I415702,I378598,I378615,I378646,I415720,I378663,I415717,I378680,I378725,I415714,I378742,I415732,I378759,I378776,I378793,I378824,I378841,I378914,I378931,I378962,I379007,I379074,I379091,I379108,I379125,I379142,I379159,I379176,I379193,I379219,I379227,I379244,I379261,I379045,I379292,I379309,I379326,I379033,I379057,I379371,I379388,I379405,I379422,I379439,I379039,I379470,I379487,I379042,I379051,I379060,I379048,I379560,I379577,I379036,I379608,I379066,I379063,I379653,I379054,I379720,I379737,I379754,I379771,I379788,I379805,I379822,I379839,I379865,I379873,I379890,I379907,I379938,I379955,I379972,I380017,I380034,I380051,I380068,I380085,I380116,I380133,I380206,I380223,I380254,I380299,I380366,I380383,I404032,I404029,I380400,I404038,I404041,I380417,I380434,I380451,I380468,I404035,I380485,I404026,I380511,I380519,I404023,I380536,I380553,I380584,I380601,I380618,I380663,I404044,I380680,I404047,I380697,I380714,I380731,I380762,I380779,I380852,I380869,I380900,I380945,I381012,I381029,I381046,I381063,I381080,I381097,I381114,I381131,I381157,I381165,I381182,I381199,I381230,I381247,I381264,I381309,I381326,I381343,I381360,I381377,I381408,I381425,I381498,I381515,I381546,I381591,I381658,I381675,I417129,I417102,I381692,I417099,I417117,I381709,I381726,I381743,I381760,I417120,I417105,I381777,I417123,I381803,I381811,I417096,I381828,I381845,I381876,I417114,I381893,I417111,I381910,I381955,I417108,I381972,I417126,I381989,I382006,I382023,I382054,I382071,I382144,I382161,I382192,I382237,I382304,I382321,I382338,I382355,I382372,I382389,I382406,I382423,I382449,I382457,I382474,I382491,I382522,I382539,I382556,I382601,I382618,I382635,I382652,I382669,I382700,I382717,I382790,I382807,I382838,I382883,I382950,I382967,I382984,I383001,I383018,I383035,I383052,I383069,I383095,I383103,I383120,I383137,I383168,I383185,I383202,I383247,I383264,I383281,I383298,I383315,I383346,I383363,I383436,I383453,I383484,I383529,I383596,I383613,I383630,I383647,I383664,I383681,I383698,I383715,I383741,I383749,I383766,I383783,I383814,I383831,I383848,I383893,I383910,I383927,I383944,I383961,I383992,I384009,I384082,I384099,I384130,I384175,I384242,I384259,I384276,I384293,I384310,I384327,I384344,I384361,I384387,I384395,I384412,I384429,I384213,I384460,I384477,I384494,I384201,I384225,I384539,I384556,I384573,I384590,I384607,I384207,I384638,I384655,I384210,I384219,I384228,I384216,I384728,I384745,I384204,I384776,I384234,I384231,I384821,I384222,I384888,I384905,I384922,I384939,I384956,I384973,I384990,I385007,I385033,I385041,I385058,I385075,I384859,I385106,I385123,I385140,I384847,I384871,I385185,I385202,I385219,I385236,I385253,I384853,I385284,I385301,I384856,I384865,I384874,I384862,I385374,I385391,I384850,I385422,I384880,I384877,I385467,I384868,I385534,I385551,I427584,I427557,I385568,I427554,I427572,I385585,I385602,I385619,I385636,I427575,I427560,I385653,I427578,I385679,I385687,I427551,I385704,I385721,I385752,I427569,I385769,I427566,I385786,I385831,I427563,I385848,I427581,I385865,I385882,I385899,I385930,I385947,I386020,I386037,I386068,I386113,I386180,I386197,I386214,I386231,I386248,I386265,I386282,I386299,I386325,I386333,I386350,I386367,I386398,I386415,I386432,I386477,I386494,I386511,I386528,I386545,I386576,I386593,I386666,I386683,I386714,I386759,I386826,I386843,I386860,I386877,I386894,I386911,I386928,I386945,I386971,I386979,I386996,I387013,I387044,I387061,I387078,I387123,I387140,I387157,I387174,I387191,I387222,I387239,I387312,I387329,I387360,I387405,I387472,I387489,I387506,I387523,I387540,I387557,I387574,I387591,I387617,I387625,I387642,I387659,I387690,I387707,I387724,I387769,I387786,I387803,I387820,I387837,I387868,I387885,I387958,I387975,I388006,I388051,I388118,I388135,I388152,I388169,I388186,I388203,I388220,I388237,I388263,I388271,I388288,I388305,I388336,I388353,I388370,I388415,I388432,I388449,I388466,I388483,I388514,I388531,I388604,I388621,I388652,I388697,I388764,I388781,I388798,I388815,I388832,I388849,I388866,I388883,I388909,I388917,I388934,I388951,I388982,I388999,I389016,I389061,I389078,I389095,I389112,I389129,I389160,I389177,I389250,I389267,I389298,I389343,I389410,I389427,I389444,I389461,I389478,I389495,I389512,I389529,I389555,I389563,I389580,I389597,I389628,I389645,I389662,I389707,I389724,I389741,I389758,I389775,I389806,I389823,I389896,I389913,I389944,I389989,I390056,I390073,I390090,I390107,I390124,I390141,I390158,I390175,I390201,I390209,I390226,I390243,I390274,I390291,I390308,I390353,I390370,I390387,I390404,I390421,I390452,I390469,I390542,I390559,I390590,I390635,I390702,I390719,I390736,I390753,I390770,I390787,I390804,I390821,I390847,I390855,I390872,I390889,I390920,I390937,I390954,I390999,I391016,I391033,I391050,I391067,I391098,I391115,I391188,I391205,I391236,I391281,I391348,I391365,I391382,I391399,I391416,I391433,I391450,I391467,I391493,I391501,I391518,I391535,I391319,I391566,I391583,I391600,I391307,I391331,I391645,I391662,I391679,I391696,I391713,I391313,I391744,I391761,I391316,I391325,I391334,I391322,I391834,I391851,I391310,I391882,I391340,I391337,I391927,I391328,I391994,I392011,I392028,I392045,I392062,I392079,I392096,I392113,I392139,I392147,I392164,I392181,I391965,I392212,I392229,I392246,I391953,I391977,I392291,I392308,I392325,I392342,I392359,I391959,I392390,I392407,I391962,I391971,I391980,I391968,I392480,I392497,I391956,I392528,I391986,I391983,I392573,I391974,I392640,I392657,I392674,I392691,I392708,I392725,I392742,I392759,I392785,I392793,I392810,I392827,I392858,I392875,I392892,I392937,I392954,I392971,I392988,I393005,I393036,I393053,I393126,I393143,I393174,I393219,I393286,I393303,I393320,I393337,I393354,I393371,I393388,I393405,I393431,I393439,I393456,I393473,I393504,I393521,I393538,I393583,I393600,I393617,I393634,I393651,I393682,I393699,I393772,I393789,I393820,I393865,I393932,I393949,I393966,I393983,I394000,I394017,I394034,I394051,I394077,I394085,I394102,I394119,I394150,I394167,I394184,I394229,I394246,I394263,I394280,I394297,I394328,I394345,I394418,I394435,I394466,I394511,I394578,I394595,I394612,I394629,I394646,I394663,I394680,I394697,I394723,I394731,I394748,I394765,I394549,I394796,I394813,I394830,I394537,I394561,I394875,I394892,I394909,I394926,I394943,I394543,I394974,I394991,I394546,I394555,I394564,I394552,I395064,I395081,I394540,I395112,I394570,I394567,I395157,I394558,I395215,I395232,I395249,I395266,I395283,I395300,I395317,I395334,I395351,I395368,I395385,I395402,I395419,I395436,I395453,I395470,I395529,I395546,I395577,I395594,I395625,I395656,I395673,I395690,I395707,I395724,I395741,I395758,I395789,I395806,I395837,I395895,I395912,I395929,I395946,I395963,I395980,I395997,I396014,I396031,I396048,I396065,I396082,I396099,I396116,I396133,I396150,I396209,I396226,I396257,I396274,I396305,I396336,I396353,I396370,I396387,I396404,I396421,I396438,I396469,I396486,I396517,I396575,I396592,I396609,I396626,I396643,I396660,I396677,I396694,I396711,I396728,I396745,I396762,I396779,I396796,I396813,I396830,I396889,I396906,I396937,I396954,I396985,I397016,I397033,I397050,I397067,I397084,I397101,I397118,I397149,I397166,I397197,I397255,I397272,I397289,I397306,I397323,I397340,I397357,I397374,I397391,I397408,I397425,I397442,I397459,I397476,I397493,I397510,I397569,I397586,I397617,I397634,I397665,I397696,I397713,I397730,I397747,I397764,I397781,I397798,I397829,I397846,I397877,I397935,I397952,I397969,I397986,I398003,I398020,I398037,I398054,I398071,I398088,I398105,I398122,I398139,I398156,I398173,I398190,I398249,I398266,I398297,I398314,I398345,I398376,I398393,I398410,I398427,I398444,I398461,I398478,I398509,I398526,I398557,I398615,I398632,I398649,I398666,I398683,I398700,I398717,I398734,I398751,I398768,I398785,I398802,I398819,I398836,I398853,I398870,I398929,I398946,I398977,I398994,I399025,I399056,I399073,I399090,I399107,I399124,I399141,I399158,I399189,I399206,I399237,I399295,I399312,I399329,I399346,I399363,I399380,I399397,I399414,I399431,I399448,I399465,I399482,I399499,I399516,I399533,I399550,I399609,I399626,I399657,I399674,I399705,I399736,I399753,I399770,I399787,I399804,I399821,I399838,I399869,I399886,I399917,I399975,I399992,I400009,I400026,I400043,I400060,I400077,I400094,I400111,I400128,I400145,I400162,I400179,I400196,I400213,I400230,I400289,I400306,I400337,I400354,I400385,I400416,I400433,I400450,I400467,I400484,I400501,I400518,I400549,I400566,I400597,I400655,I400672,I400689,I400706,I400723,I400740,I400757,I400774,I400791,I400808,I400825,I400842,I400859,I400876,I400893,I400910,I400969,I400986,I401017,I401034,I401065,I401096,I401113,I401130,I401147,I401164,I401181,I401198,I401229,I401246,I401277,I401335,I401352,I401369,I401386,I401403,I401420,I401437,I401454,I401471,I401488,I401505,I401522,I401539,I401556,I401573,I401590,I401649,I401666,I401697,I401714,I401745,I401776,I401793,I401810,I401827,I401844,I401861,I401878,I401909,I401926,I401957,I402015,I402032,I402049,I402066,I402083,I402100,I402117,I402134,I402151,I402168,I402185,I402202,I402219,I402236,I402253,I402270,I402329,I402346,I402377,I402394,I402425,I402456,I402473,I402490,I402507,I402524,I402541,I402558,I402589,I402606,I402637,I402695,I402712,I402729,I402746,I402763,I402780,I402797,I402814,I402831,I402848,I402865,I402882,I402899,I402916,I402933,I402950,I403009,I403026,I403057,I403074,I403105,I403136,I403153,I403170,I403187,I403204,I403221,I403238,I403269,I403286,I403317,I403375,I403392,I403409,I403426,I403443,I403460,I403477,I403494,I403511,I403528,I403545,I403562,I403579,I403596,I403613,I403630,I403689,I403706,I403737,I403754,I403785,I403816,I403833,I403850,I403867,I403884,I403901,I403918,I403949,I403966,I403997,I404055,I404072,I404089,I404106,I404123,I404140,I404157,I404174,I404191,I404208,I404225,I404242,I404259,I404276,I404293,I404310,I404369,I404386,I404417,I404434,I404465,I404496,I404513,I404530,I404547,I404564,I404581,I404598,I404629,I404646,I404677,I404735,I404752,I404769,I404786,I404803,I404820,I404837,I404854,I404871,I404888,I404905,I404922,I404939,I404956,I404973,I404990,I405049,I405066,I405097,I405114,I405145,I405176,I405193,I405210,I405227,I405244,I405261,I405278,I405309,I405326,I405357,I405415,I405432,I405449,I405466,I405483,I405500,I405517,I405534,I405551,I405568,I405585,I405602,I405619,I405636,I405653,I405670,I405729,I405746,I405777,I405794,I405825,I405856,I405873,I405890,I405907,I405924,I405941,I405958,I405989,I406006,I406037,I406095,I406112,I406129,I406146,I406163,I406180,I406197,I406214,I406231,I406248,I406265,I406282,I406299,I406316,I406333,I406350,I406409,I406426,I406457,I406474,I406505,I406536,I406553,I406570,I406587,I406604,I406621,I406638,I406669,I406686,I406717,I406775,I406792,I406809,I406826,I406843,I406860,I406877,I406894,I406911,I406928,I406945,I406962,I406979,I406996,I407013,I407030,I407089,I407106,I407137,I407154,I407185,I407216,I407233,I407250,I407267,I407284,I407301,I407318,I407349,I407366,I407397,I407455,I407472,I407489,I407506,I407523,I407540,I407557,I407574,I407591,I407608,I407625,I407642,I407659,I407676,I407693,I407710,I407769,I407786,I407817,I407834,I407865,I407896,I407913,I407930,I407947,I407964,I407981,I407998,I408029,I408046,I408077,I408135,I408152,I408169,I408186,I408203,I408220,I408237,I408254,I408271,I408288,I408305,I408322,I408339,I408356,I408373,I408390,I408449,I408466,I408497,I408514,I408545,I408576,I408593,I408610,I408627,I408644,I408661,I408678,I408709,I408726,I408757,I408815,I408832,I408849,I408866,I408883,I408900,I408917,I408934,I408951,I408968,I408985,I409002,I409019,I409036,I409053,I409070,I409129,I409146,I409177,I409194,I409225,I409256,I409273,I409290,I409307,I409324,I409341,I409358,I409389,I409406,I409437,I409495,I409512,I409529,I409546,I409563,I409580,I409597,I409614,I409631,I409648,I409665,I409682,I409699,I409716,I409733,I409750,I409809,I409826,I409857,I409874,I409905,I409936,I409953,I409970,I409987,I410004,I410021,I410038,I410069,I410086,I410117,I410175,I410192,I410209,I410226,I410243,I410260,I410277,I410294,I410311,I410328,I410345,I410362,I410379,I410396,I410413,I410430,I410489,I410506,I410537,I410554,I410585,I410616,I410633,I410650,I410667,I410684,I410701,I410718,I410749,I410766,I410797,I410864,I410881,I410898,I410924,I410932,I410949,I410966,I410983,I411000,I411017,I411034,I411051,I411068,I411085,I411102,I411119,I411136,I411153,I411184,I411201,I411218,I411263,I411308,I411325,I411370,I411387,I411418,I411435,I411466,I411561,I411578,I411595,I411621,I411629,I411646,I411663,I411680,I411697,I411714,I411731,I411748,I411765,I411782,I411799,I411816,I411833,I411850,I411881,I411898,I411915,I411960,I412005,I412022,I412067,I412084,I412115,I412132,I412163,I412258,I412275,I412292,I412318,I412326,I412343,I412360,I412377,I412394,I412411,I412428,I412445,I412462,I412479,I412496,I412513,I412530,I412547,I412578,I412595,I412612,I412657,I412702,I412719,I412764,I412781,I412812,I412829,I412860,I412955,I412972,I412989,I413015,I413023,I413040,I413057,I413074,I413091,I413108,I413125,I413142,I413159,I413176,I413193,I413210,I413227,I413244,I413275,I413292,I413309,I413354,I413399,I413416,I413461,I413478,I413509,I413526,I413557,I413652,I413669,I413686,I413712,I413720,I413737,I413754,I413771,I413788,I413805,I413822,I413839,I413856,I413873,I413890,I413907,I413924,I413941,I413972,I413989,I414006,I414051,I414096,I414113,I414158,I414175,I414206,I414223,I414254,I414349,I414366,I414383,I414409,I414417,I414434,I414451,I414468,I414485,I414502,I414519,I414536,I414553,I414570,I414587,I414604,I414621,I414638,I414669,I414686,I414703,I414748,I414793,I414810,I414855,I414872,I414903,I414920,I414951,I415046,I415063,I415080,I415106,I415114,I415131,I415148,I415165,I415182,I415199,I415216,I415233,I415250,I415267,I415284,I415301,I415318,I415335,I415366,I415383,I415400,I415445,I415490,I415507,I415552,I415569,I415600,I415617,I415648,I415743,I415760,I415777,I415803,I415811,I415828,I415845,I415862,I415879,I415896,I415913,I415930,I415947,I415964,I415981,I415998,I416015,I416032,I416063,I416080,I416097,I416142,I416187,I416204,I416249,I416266,I416297,I416314,I416345,I416440,I416457,I416474,I416500,I416508,I416525,I416542,I416559,I416576,I416593,I416610,I416627,I416644,I416661,I416678,I416695,I416712,I416729,I416760,I416777,I416794,I416839,I416884,I416901,I416946,I416963,I416994,I417011,I417042,I417137,I417154,I417171,I417197,I417205,I417222,I417239,I417256,I417273,I417290,I417307,I417324,I417341,I417358,I417375,I417392,I417409,I417426,I417457,I417474,I417491,I417536,I417581,I417598,I417643,I417660,I417691,I417708,I417739,I417834,I417851,I417868,I417894,I417902,I417919,I417936,I417953,I417970,I417987,I418004,I418021,I418038,I418055,I418072,I418089,I418106,I418123,I418154,I418171,I418188,I418233,I418278,I418295,I418340,I418357,I418388,I418405,I418436,I418531,I418548,I418565,I418591,I418599,I418616,I418633,I418650,I418667,I418684,I418701,I418718,I418735,I418752,I418769,I418786,I418803,I418820,I418851,I418868,I418885,I418930,I418975,I418992,I419037,I419054,I419085,I419102,I419133,I419228,I419245,I419262,I419288,I419296,I419313,I419330,I419347,I419364,I419381,I419398,I419415,I419432,I419449,I419466,I419483,I419500,I419517,I419548,I419565,I419582,I419627,I419672,I419689,I419734,I419751,I419782,I419799,I419830,I419925,I419942,I419959,I419985,I419993,I420010,I420027,I420044,I420061,I420078,I420095,I420112,I420129,I420146,I420163,I420180,I420197,I420214,I420245,I420262,I420279,I420324,I420369,I420386,I420431,I420448,I420479,I420496,I420527,I420622,I420639,I420656,I420682,I420690,I420707,I420724,I420741,I420758,I420775,I420792,I420809,I420826,I420843,I420860,I420877,I420894,I420911,I420942,I420959,I420976,I421021,I421066,I421083,I421128,I421145,I421176,I421193,I421224,I421319,I421336,I421353,I421379,I421387,I421404,I421421,I421438,I421455,I421472,I421489,I421506,I421523,I421540,I421557,I421574,I421591,I421608,I421639,I421656,I421673,I421718,I421763,I421780,I421825,I421842,I421873,I421890,I421921,I422016,I422033,I422050,I422076,I422084,I422101,I422118,I422135,I422152,I422169,I422186,I422203,I422220,I422237,I422254,I422271,I422288,I422305,I422336,I422353,I422370,I422415,I422460,I422477,I422522,I422539,I422570,I422587,I422618,I422713,I422730,I422747,I422773,I422781,I422798,I422815,I422832,I422849,I422866,I422883,I422900,I422917,I422934,I422951,I422968,I422985,I423002,I423033,I423050,I423067,I423112,I423157,I423174,I423219,I423236,I423267,I423284,I423315,I423410,I423427,I423444,I423470,I423478,I423495,I423512,I423529,I423546,I423563,I423580,I423597,I423614,I423631,I423648,I423665,I423682,I423699,I423730,I423747,I423764,I423809,I423854,I423871,I423916,I423933,I423964,I423981,I424012,I424107,I424124,I424141,I424167,I424175,I424192,I424209,I424226,I424243,I424260,I424277,I424294,I424311,I424328,I424345,I424362,I424379,I424396,I424427,I424444,I424461,I424506,I424551,I424568,I424613,I424630,I424661,I424678,I424709,I424804,I424821,I424838,I424864,I424872,I424889,I424906,I424923,I424940,I424957,I424974,I424991,I425008,I425025,I425042,I425059,I425076,I425093,I425124,I425141,I425158,I425203,I425248,I425265,I425310,I425327,I425358,I425375,I425406,I425501,I425518,I425535,I425561,I425569,I425586,I425603,I425620,I425637,I425654,I425671,I425688,I425705,I425722,I425739,I425756,I425773,I425790,I425821,I425838,I425855,I425900,I425945,I425962,I426007,I426024,I426055,I426072,I426103,I426198,I426215,I426232,I426258,I426266,I426283,I426300,I426317,I426334,I426351,I426368,I426385,I426402,I426419,I426436,I426453,I426470,I426487,I426518,I426535,I426552,I426597,I426642,I426659,I426704,I426721,I426752,I426769,I426800,I426895,I426912,I426929,I426955,I426963,I426980,I426997,I427014,I427031,I427048,I427065,I427082,I427099,I427116,I427133,I427150,I427167,I427184,I427215,I427232,I427249,I427294,I427339,I427356,I427401,I427418,I427449,I427466,I427497,I427592,I427609,I427626,I427652,I427660,I427677,I427694,I427711,I427728,I427745,I427762,I427779,I427796,I427813,I427830,I427847,I427864,I427881,I427912,I427929,I427946,I427991,I428036,I428053,I428098,I428115,I428146,I428163,I428194,I428289,I428306,I428323,I428349,I428357,I428374,I428391,I428408,I428425,I428442,I428459,I428476,I428493,I428510,I428527,I428544,I428561,I428578,I428609,I428626,I428643,I428688,I428733,I428750,I428795,I428812,I428843,I428860,I428891,I428986,I429003,I429020,I429046,I429054,I429071,I429088,I429105,I429122,I429139,I429156,I429173,I429190,I429207,I429224,I429241,I429258,I429275,I429306,I429323,I429340,I429385,I429430,I429447,I429492,I429509,I429540,I429557,I429588,I429683,I429700,I429717,I429743,I429751,I429768,I429785,I429802,I429819,I429836,I429853,I429870,I429887,I429904,I429921,I429938,I429955,I429972,I430003,I430020,I430037,I430082,I430127,I430144,I430189,I430206,I430237,I430254,I430285,I430380,I430397,I430414,I430440,I430448,I430465,I430482,I430499,I430516,I430533,I430550,I430567,I430584,I430601,I430618,I430635,I430652,I430669,I430700,I430717,I430734,I430779,I430824,I430841,I430886,I430903,I430934,I430951,I430982,I431077,I431094,I431111,I431137,I431145,I431162,I431179,I431196,I431213,I431230,I431247,I431264,I431281,I431298,I431315,I431332,I431349,I431366,I431397,I431414,I431431,I431476,I431521,I431538,I431583,I431600,I431631,I431648,I431679,I431774,I431791,I431808,I431834,I431842,I431859,I431876,I431893,I431910,I431927,I431944,I431961,I431978,I431995,I432012,I432029,I432046,I432063,I432094,I432111,I432128,I432173,I432218,I432235,I432280,I432297,I432328,I432345,I432376,I432471,I432488,I432505,I432531,I432539,I432556,I432573,I432590,I432607,I432624,I432641,I432658,I432675,I432692,I432709,I432726,I432743,I432760,I432791,I432808,I432825,I432870,I432915,I432932,I432977,I432994,I433025,I433042,I433073,I433168,I433185,I433202,I433228,I433236,I433253,I433270,I433287,I433304,I433321,I433338,I433355,I433372,I433389,I433406,I433423,I433440,I433457,I433488,I433505,I433522,I433567,I433612,I433629,I433674,I433691,I433722,I433739,I433770,I433865,I433882,I433899,I433925,I433933,I433950,I433967,I433984,I434001,I434018,I434035,I434052,I434069,I434086,I434103,I434120,I434137,I434154,I434185,I434202,I434219,I434264,I434309,I434326,I434371,I434388,I434419,I434436,I434467,I434562,I434579,I434596,I434622,I434630,I434647,I434664,I434681,I434698,I434715,I434732,I434749,I434766,I434783,I434800,I434817,I434834,I434851,I434882,I434899,I434916,I434961,I435006,I435023,I435068,I435085,I435116,I435133,I435164,I435259,I435276,I435293,I435319,I435327,I435344,I435361,I435378,I435395,I435412,I435429,I435446,I435463,I435480,I435497,I435514,I435531,I435548,I435579,I435596,I435613,I435658,I435703,I435720,I435765,I435782,I435813,I435830,I435861,I435956,I435973,I435990,I436016,I436024,I436041,I436058,I436075,I436092,I436109,I436126,I436143,I436160,I436177,I436194,I436211,I436228,I436245,I436276,I436293,I436310,I436355,I436400,I436417,I436462,I436479,I436510,I436527,I436558,I436653,I436670,I436687,I436713,I436721,I436738,I436755,I436772,I436789,I436806,I436823,I436840,I436857,I436874,I436891,I436908,I436925,I436942,I436973,I436990,I437007,I437052,I437097,I437114,I437159,I437176,I437207,I437224,I437255,I437350,I437367,I437384,I437410,I437418,I437435,I437452,I437469,I437486,I437503,I437520,I437537,I437554,I437571,I437588,I437605,I437622,I437639,I437670,I437687,I437704,I437749,I437794,I437811,I437856,I437873,I437904,I437921,I437952,I438047,I438064,I438081,I438107,I438115,I438132,I438149,I438166,I438183,I438200,I438217,I438234,I438251,I438268,I438285,I438302,I438319,I438336,I438367,I438384,I438401,I438446,I438491,I438508,I438553,I438570,I438601,I438618,I438649,I438744,I438761,I438778,I438804,I438812,I438829,I438846,I438863,I438880,I438897,I438914,I438931,I438948,I438965,I438982,I438999,I439016,I439033,I439064,I439081,I439098,I439143,I439188,I439205,I439250,I439267,I439298,I439315,I439346,I439441,I439458,I439475,I439501,I439509,I439526,I439543,I439560,I439577,I439594,I439611,I439628,I439645,I439662,I439679,I439696,I439713,I439730,I439761,I439778,I439795,I439840,I439885,I439902,I439947,I439964,I439995,I440012,I440043,I440138,I440155,I440172,I440198,I440206,I440223,I440240,I440257,I440274,I440291,I440308,I440325,I440342,I440359,I440376,I440393,I440410,I440427,I440458,I440475,I440492,I440537,I440582,I440599,I440644,I440661,I440692,I440709,I440740,I440835,I440852,I440869,I440895,I440903,I440920,I440937,I440954,I440971,I440988,I441005,I441022,I441039,I441056,I441073,I441090,I441107,I441124,I441155,I441172,I441189,I441234,I441279,I441296,I441341,I441358,I441389,I441406,I441437,I441532,I441549,I441566,I441592,I441600,I441617,I441634,I441651,I441668,I441685,I441702,I441719,I441736,I441753,I441770,I441787,I441804,I441821,I441852,I441869,I441886,I441931,I441976,I441993,I442038,I442055,I442086,I442103,I442134,I442229,I442246,I442263,I442289,I442297,I442314,I442331,I442348,I442365,I442382,I442399,I442416,I442433,I442450,I442467,I442484,I442501,I442518,I442549,I442566,I442583,I442628,I442673,I442690,I442735,I442752,I442783,I442800,I442831,I442926,I442943,I442960,I442986,I442994,I443011,I443028,I443045,I443062,I443079,I443096,I443113,I443130,I443147,I443164,I443181,I443198,I443215,I443246,I443263,I443280,I443325,I443370,I443387,I443432,I443449,I443480,I443497,I443528,I443623,I443640,I443657,I443683,I443691,I443708,I443725,I443742,I443759,I443776,I443793,I443810,I443827,I443844,I443861,I443878,I443895,I443912,I443943,I443960,I443977,I444022,I444067,I444084,I444129,I444146,I444177,I444194,I444225,I444320,I444337,I444354,I444380,I444388,I444405,I444422,I444439,I444456,I444473,I444490,I444507,I444524,I444541,I444558,I444575,I444592,I444609,I444640,I444657,I444674,I444719,I444764,I444781,I444826,I444843,I444874,I444891,I444922,I445017,I445034,I445051,I445077,I445085,I445102,I445119,I445136,I445153,I445170,I445187,I445204,I445221,I445238,I445255,I445272,I445289,I445306,I445337,I445354,I445371,I445416,I445461,I445478,I445523,I445540,I445571,I445588,I445619,I445714,I445731,I445748,I445774,I445782,I445799,I445816,I445833,I445850,I445867,I445884,I445901,I445918,I445935,I445952,I445969,I445986,I446003,I446034,I446051,I446068,I446113,I446158,I446175,I446220,I446237,I446268,I446285,I446316;
not I_0 (I2946,I2905);
or I_1 (I2963,I275784,I275793);
nor I_2 (I2980,I275784,I275793);
nor I_3 (I2997,I2980,I275787);
nand I_4 (I3014,I2963,I275790);
not I_5 (I3031,I3014);
nor I_6 (I3048,I2997,I3031);
or I_7 (I2914,I3014,I275796);
nor I_8 (I2929,I3031,I275796);
and I_9 (I3093,I275802,I275778);
nor I_10 (I3110,I3093,I275805);
nand I_11 (I3127,I275781,I275781);
nor I_12 (I3144,I3127,I3110);
not I_13 (I3161,I3144);
nor I_14 (I2911,I3161,I3048);
nor I_15 (I3192,I3161,I275796);
nor I_16 (I3209,I3144,I275796);
nand I_17 (I2923,I2997,I3209);
nor I_18 (I3240,I3144,I3127);
nand I_19 (I2920,I3240,I275796);
not I_20 (I3271,I3127);
nor I_21 (I3288,I3031,I3271);
DFFARX1 I_22 (I3288,I2898,I2946,I2926,);
nor I_23 (I3319,I3271,I3014);
nor I_24 (I3336,I275775,I275778);
or I_25 (I3353,I3336,I275775);
nor I_26 (I3370,I275784,I275799);
nand I_27 (I3387,I3370,I3353);
not I_28 (I3404,I3387);
nor I_29 (I2908,I3161,I3404);
nand I_30 (I3435,I3404,I3319);
nand I_31 (I3452,I3161,I3435);
DFFARX1 I_32 (I3452,I2898,I2946,I2917,);
nor I_33 (I2935,I3404,I3192);
or I_34 (I2932,I3404,I2997);
nand I_35 (I2938,I3127,I3387);
not I_36 (I3558,I2905);
or I_37 (I3575,I435245,I435251);
nor I_38 (I3592,I435245,I435251);
nor I_39 (I3609,I3592,I435221);
nand I_40 (I3626,I3575,I435242);
not I_41 (I3643,I3626);
nor I_42 (I3660,I3609,I3643);
or I_43 (I3526,I3626,I435224);
nor I_44 (I3541,I3643,I435224);
and I_45 (I3705,I435233,I435227);
nor I_46 (I3722,I3705,I435221);
nand I_47 (I3739,I435248,I435239);
nor I_48 (I3756,I3739,I3722);
not I_49 (I3773,I3756);
nor I_50 (I3523,I3773,I3660);
nor I_51 (I3804,I3773,I435224);
nor I_52 (I3821,I3756,I435224);
nand I_53 (I3535,I3609,I3821);
nor I_54 (I3852,I3756,I3739);
nand I_55 (I3532,I3852,I435224);
not I_56 (I3883,I3739);
nor I_57 (I3900,I3643,I3883);
DFFARX1 I_58 (I3900,I2898,I3558,I3538,);
nor I_59 (I3931,I3883,I3626);
nor I_60 (I3948,I435218,I435236);
or I_61 (I3965,I3948,I435224);
nor I_62 (I3982,I435230,I435218);
nand I_63 (I3999,I3982,I3965);
not I_64 (I4016,I3999);
nor I_65 (I3520,I3773,I4016);
nand I_66 (I4047,I4016,I3931);
nand I_67 (I4064,I3773,I4047);
DFFARX1 I_68 (I4064,I2898,I3558,I3529,);
nor I_69 (I3547,I4016,I3804);
or I_70 (I3544,I4016,I3609);
nand I_71 (I3550,I3739,I3999);
not I_72 (I4170,I2905);
or I_73 (I4187,I145680,I145686);
nor I_74 (I4204,I145680,I145686);
nor I_75 (I4221,I4204,I145674);
nand I_76 (I4238,I4187,I145701);
not I_77 (I4255,I4238);
nor I_78 (I4272,I4221,I4255);
or I_79 (I4138,I4238,I145683);
nor I_80 (I4153,I4255,I145683);
and I_81 (I4317,I145704,I145707);
nor I_82 (I4334,I4317,I145692);
nand I_83 (I4351,I145677,I145698);
nor I_84 (I4368,I4351,I4334);
not I_85 (I4385,I4368);
nor I_86 (I4135,I4385,I4272);
nor I_87 (I4416,I4385,I145683);
nor I_88 (I4433,I4368,I145683);
nand I_89 (I4147,I4221,I4433);
nor I_90 (I4464,I4368,I4351);
nand I_91 (I4144,I4464,I145683);
not I_92 (I4495,I4351);
nor I_93 (I4512,I4255,I4495);
DFFARX1 I_94 (I4512,I2898,I4170,I4150,);
nor I_95 (I4543,I4495,I4238);
nor I_96 (I4560,I145674,I145695);
or I_97 (I4577,I4560,I145677);
nor I_98 (I4594,I145689,I145680);
nand I_99 (I4611,I4594,I4577);
not I_100 (I4628,I4611);
nor I_101 (I4132,I4385,I4628);
nand I_102 (I4659,I4628,I4543);
nand I_103 (I4676,I4385,I4659);
DFFARX1 I_104 (I4676,I2898,I4170,I4141,);
nor I_105 (I4159,I4628,I4416);
or I_106 (I4156,I4628,I4221);
nand I_107 (I4162,I4351,I4611);
not I_108 (I4782,I2905);
or I_109 (I4799,I154520,I154526);
nor I_110 (I4816,I154520,I154526);
nor I_111 (I4833,I4816,I154514);
nand I_112 (I4850,I4799,I154541);
not I_113 (I4867,I4850);
nor I_114 (I4884,I4833,I4867);
or I_115 (I4750,I4850,I154523);
nor I_116 (I4765,I4867,I154523);
and I_117 (I4929,I154544,I154547);
nor I_118 (I4946,I4929,I154532);
nand I_119 (I4963,I154517,I154538);
nor I_120 (I4980,I4963,I4946);
not I_121 (I4997,I4980);
nor I_122 (I4747,I4997,I4884);
nor I_123 (I5028,I4997,I154523);
nor I_124 (I5045,I4980,I154523);
nand I_125 (I4759,I4833,I5045);
nor I_126 (I5076,I4980,I4963);
nand I_127 (I4756,I5076,I154523);
not I_128 (I5107,I4963);
nor I_129 (I5124,I4867,I5107);
DFFARX1 I_130 (I5124,I2898,I4782,I4762,);
nor I_131 (I5155,I5107,I4850);
nor I_132 (I5172,I154514,I154535);
or I_133 (I5189,I5172,I154517);
nor I_134 (I5206,I154529,I154520);
nand I_135 (I5223,I5206,I5189);
not I_136 (I5240,I5223);
nor I_137 (I4744,I4997,I5240);
nand I_138 (I5271,I5240,I5155);
nand I_139 (I5288,I4997,I5271);
DFFARX1 I_140 (I5288,I2898,I4782,I4753,);
nor I_141 (I4771,I5240,I5028);
or I_142 (I4768,I5240,I4833);
nand I_143 (I4774,I4963,I5223);
not I_144 (I5394,I2905);
or I_145 (I5411,I360920,I360920);
nor I_146 (I5428,I360920,I360920);
nor I_147 (I5445,I5428,I360923);
nand I_148 (I5462,I5411,I360932);
not I_149 (I5479,I5462);
nor I_150 (I5496,I5445,I5479);
or I_151 (I5362,I5462,I360917);
nor I_152 (I5377,I5479,I360917);
and I_153 (I5541,I360914,I360923);
nor I_154 (I5558,I5541,I360926);
nand I_155 (I5575,I360914,I360911);
nor I_156 (I5592,I5575,I5558);
not I_157 (I5609,I5592);
nor I_158 (I5359,I5609,I5496);
nor I_159 (I5640,I5609,I360917);
nor I_160 (I5657,I5592,I360917);
nand I_161 (I5371,I5445,I5657);
nor I_162 (I5688,I5592,I5575);
nand I_163 (I5368,I5688,I360917);
not I_164 (I5719,I5575);
nor I_165 (I5736,I5479,I5719);
DFFARX1 I_166 (I5736,I2898,I5394,I5374,);
nor I_167 (I5767,I5719,I5462);
nor I_168 (I5784,I360917,I360911);
or I_169 (I5801,I5784,I360926);
nor I_170 (I5818,I360935,I360929);
nand I_171 (I5835,I5818,I5801);
not I_172 (I5852,I5835);
nor I_173 (I5356,I5609,I5852);
nand I_174 (I5883,I5852,I5767);
nand I_175 (I5900,I5609,I5883);
DFFARX1 I_176 (I5900,I2898,I5394,I5365,);
nor I_177 (I5383,I5852,I5640);
or I_178 (I5380,I5852,I5445);
nand I_179 (I5386,I5575,I5835);
not I_180 (I6006,I2905);
or I_181 (I6023,I23206,I23224);
nor I_182 (I6040,I23206,I23224);
nor I_183 (I6057,I6040,I23215);
nand I_184 (I6074,I6023,I23209);
not I_185 (I6091,I6074);
nor I_186 (I6108,I6057,I6091);
or I_187 (I5974,I6074,I23212);
nor I_188 (I5989,I6091,I23212);
and I_189 (I6153,I23227,I23209);
nor I_190 (I6170,I6153,I23218);
nand I_191 (I6187,I23221,I23215);
nor I_192 (I6204,I6187,I6170);
not I_193 (I6221,I6204);
nor I_194 (I5971,I6221,I6108);
nor I_195 (I6252,I6221,I23212);
nor I_196 (I6269,I6204,I23212);
nand I_197 (I5983,I6057,I6269);
nor I_198 (I6300,I6204,I6187);
nand I_199 (I5980,I6300,I23212);
not I_200 (I6331,I6187);
nor I_201 (I6348,I6091,I6331);
DFFARX1 I_202 (I6348,I2898,I6006,I5986,);
nor I_203 (I6379,I6331,I6074);
nor I_204 (I6396,I23212,I23218);
or I_205 (I6413,I6396,I23230);
nor I_206 (I6430,I23206,I23233);
nand I_207 (I6447,I6430,I6413);
not I_208 (I6464,I6447);
nor I_209 (I5968,I6221,I6464);
nand I_210 (I6495,I6464,I6379);
nand I_211 (I6512,I6221,I6495);
DFFARX1 I_212 (I6512,I2898,I6006,I5977,);
nor I_213 (I5995,I6464,I6252);
or I_214 (I5992,I6464,I6057);
nand I_215 (I5998,I6187,I6447);
not I_216 (I6618,I2905);
or I_217 (I6635,I115380,I115386);
nor I_218 (I6652,I115380,I115386);
nor I_219 (I6669,I6652,I115392);
nand I_220 (I6686,I6635,I115383);
not I_221 (I6703,I6686);
nor I_222 (I6720,I6669,I6703);
or I_223 (I6586,I6686,I115407);
nor I_224 (I6601,I6703,I115407);
and I_225 (I6765,I115404,I115389);
nor I_226 (I6782,I6765,I115413);
nand I_227 (I6799,I115401,I115410);
nor I_228 (I6816,I6799,I6782);
not I_229 (I6833,I6816);
nor I_230 (I6583,I6833,I6720);
nor I_231 (I6864,I6833,I115407);
nor I_232 (I6881,I6816,I115407);
nand I_233 (I6595,I6669,I6881);
nor I_234 (I6912,I6816,I6799);
nand I_235 (I6592,I6912,I115407);
not I_236 (I6943,I6799);
nor I_237 (I6960,I6703,I6943);
DFFARX1 I_238 (I6960,I2898,I6618,I6598,);
nor I_239 (I6991,I6943,I6686);
nor I_240 (I7008,I115395,I115383);
or I_241 (I7025,I7008,I115386);
nor I_242 (I7042,I115398,I115380);
nand I_243 (I7059,I7042,I7025);
not I_244 (I7076,I7059);
nor I_245 (I6580,I6833,I7076);
nand I_246 (I7107,I7076,I6991);
nand I_247 (I7124,I6833,I7107);
DFFARX1 I_248 (I7124,I2898,I6618,I6589,);
nor I_249 (I6607,I7076,I6864);
or I_250 (I6604,I7076,I6669);
nand I_251 (I6610,I6799,I7059);
not I_252 (I7230,I2905);
or I_253 (I7247,I272724,I272733);
nor I_254 (I7264,I272724,I272733);
nor I_255 (I7281,I7264,I272727);
nand I_256 (I7298,I7247,I272730);
not I_257 (I7315,I7298);
nor I_258 (I7332,I7281,I7315);
or I_259 (I7198,I7298,I272736);
nor I_260 (I7213,I7315,I272736);
and I_261 (I7377,I272742,I272718);
nor I_262 (I7394,I7377,I272745);
nand I_263 (I7411,I272721,I272721);
nor I_264 (I7428,I7411,I7394);
not I_265 (I7445,I7428);
nor I_266 (I7195,I7445,I7332);
nor I_267 (I7476,I7445,I272736);
nor I_268 (I7493,I7428,I272736);
nand I_269 (I7207,I7281,I7493);
nor I_270 (I7524,I7428,I7411);
nand I_271 (I7204,I7524,I272736);
not I_272 (I7555,I7411);
nor I_273 (I7572,I7315,I7555);
DFFARX1 I_274 (I7572,I2898,I7230,I7210,);
nor I_275 (I7603,I7555,I7298);
nor I_276 (I7620,I272715,I272718);
or I_277 (I7637,I7620,I272715);
nor I_278 (I7654,I272724,I272739);
nand I_279 (I7671,I7654,I7637);
not I_280 (I7688,I7671);
nor I_281 (I7192,I7445,I7688);
nand I_282 (I7719,I7688,I7603);
nand I_283 (I7736,I7445,I7719);
DFFARX1 I_284 (I7736,I2898,I7230,I7201,);
nor I_285 (I7219,I7688,I7476);
or I_286 (I7216,I7688,I7281);
nand I_287 (I7222,I7411,I7671);
not I_288 (I7842,I2905);
or I_289 (I7859,I184166,I184151);
nor I_290 (I7876,I184166,I184151);
nor I_291 (I7893,I7876,I184148);
nand I_292 (I7910,I7859,I184160);
not I_293 (I7927,I7910);
nor I_294 (I7944,I7893,I7927);
or I_295 (I7810,I7910,I184148);
nor I_296 (I7825,I7927,I184148);
and I_297 (I7989,I184157,I184169);
nor I_298 (I8006,I7989,I184154);
nand I_299 (I8023,I184163,I184160);
nor I_300 (I8040,I8023,I8006);
not I_301 (I8057,I8040);
nor I_302 (I7807,I8057,I7944);
nor I_303 (I8088,I8057,I184148);
nor I_304 (I8105,I8040,I184148);
nand I_305 (I7819,I7893,I8105);
nor I_306 (I8136,I8040,I8023);
nand I_307 (I7816,I8136,I184148);
not I_308 (I8167,I8023);
nor I_309 (I8184,I7927,I8167);
DFFARX1 I_310 (I8184,I2898,I7842,I7822,);
nor I_311 (I8215,I8167,I7910);
nor I_312 (I8232,I184151,I184157);
or I_313 (I8249,I8232,I184154);
nor I_314 (I8266,I184145,I184145);
nand I_315 (I8283,I8266,I8249);
not I_316 (I8300,I8283);
nor I_317 (I7804,I8057,I8300);
nand I_318 (I8331,I8300,I8215);
nand I_319 (I8348,I8057,I8331);
DFFARX1 I_320 (I8348,I2898,I7842,I7813,);
nor I_321 (I7831,I8300,I8088);
or I_322 (I7828,I8300,I7893);
nand I_323 (I7834,I8023,I8283);
not I_324 (I8454,I2905);
or I_325 (I8471,I252069,I252078);
nor I_326 (I8488,I252069,I252078);
nor I_327 (I8505,I8488,I252072);
nand I_328 (I8522,I8471,I252075);
not I_329 (I8539,I8522);
nor I_330 (I8556,I8505,I8539);
or I_331 (I8422,I8522,I252081);
nor I_332 (I8437,I8539,I252081);
and I_333 (I8601,I252087,I252063);
nor I_334 (I8618,I8601,I252090);
nand I_335 (I8635,I252066,I252066);
nor I_336 (I8652,I8635,I8618);
not I_337 (I8669,I8652);
nor I_338 (I8419,I8669,I8556);
nor I_339 (I8700,I8669,I252081);
nor I_340 (I8717,I8652,I252081);
nand I_341 (I8431,I8505,I8717);
nor I_342 (I8748,I8652,I8635);
nand I_343 (I8428,I8748,I252081);
not I_344 (I8779,I8635);
nor I_345 (I8796,I8539,I8779);
DFFARX1 I_346 (I8796,I2898,I8454,I8434,);
nor I_347 (I8827,I8779,I8522);
nor I_348 (I8844,I252060,I252063);
or I_349 (I8861,I8844,I252060);
nor I_350 (I8878,I252069,I252084);
nand I_351 (I8895,I8878,I8861);
not I_352 (I8912,I8895);
nor I_353 (I8416,I8669,I8912);
nand I_354 (I8943,I8912,I8827);
nand I_355 (I8960,I8669,I8943);
DFFARX1 I_356 (I8960,I2898,I8454,I8425,);
nor I_357 (I8443,I8912,I8700);
or I_358 (I8440,I8912,I8505);
nand I_359 (I8446,I8635,I8895);
not I_360 (I9066,I2905);
or I_361 (I9083,I403343,I403358);
nor I_362 (I9100,I403343,I403358);
nor I_363 (I9117,I9100,I403358);
nand I_364 (I9134,I9083,I403349);
not I_365 (I9151,I9134);
nor I_366 (I9168,I9117,I9151);
or I_367 (I9034,I9134,I403355);
nor I_368 (I9049,I9151,I403355);
and I_369 (I9213,I403346,I403346);
nor I_370 (I9230,I9213,I403343);
nand I_371 (I9247,I403352,I403361);
nor I_372 (I9264,I9247,I9230);
not I_373 (I9281,I9264);
nor I_374 (I9031,I9281,I9168);
nor I_375 (I9312,I9281,I403355);
nor I_376 (I9329,I9264,I403355);
nand I_377 (I9043,I9117,I9329);
nor I_378 (I9360,I9264,I9247);
nand I_379 (I9040,I9360,I403355);
not I_380 (I9391,I9247);
nor I_381 (I9408,I9151,I9391);
DFFARX1 I_382 (I9408,I2898,I9066,I9046,);
nor I_383 (I9439,I9391,I9134);
nor I_384 (I9456,I403349,I403364);
or I_385 (I9473,I9456,I403355);
nor I_386 (I9490,I403352,I403367);
nand I_387 (I9507,I9490,I9473);
not I_388 (I9524,I9507);
nor I_389 (I9028,I9281,I9524);
nand I_390 (I9555,I9524,I9439);
nand I_391 (I9572,I9281,I9555);
DFFARX1 I_392 (I9572,I2898,I9066,I9037,);
nor I_393 (I9055,I9524,I9312);
or I_394 (I9052,I9524,I9117);
nand I_395 (I9058,I9247,I9507);
not I_396 (I9678,I2905);
or I_397 (I9695,I227651,I227657);
nor I_398 (I9712,I227651,I227657);
nor I_399 (I9729,I9712,I227675);
nand I_400 (I9746,I9695,I227654);
not I_401 (I9763,I9746);
nor I_402 (I9780,I9729,I9763);
or I_403 (I9646,I9746,I227663);
nor I_404 (I9661,I9763,I227663);
and I_405 (I9825,I227666,I227660);
nor I_406 (I9842,I9825,I227672);
nand I_407 (I9859,I227660,I227651);
nor I_408 (I9876,I9859,I9842);
not I_409 (I9893,I9876);
nor I_410 (I9643,I9893,I9780);
nor I_411 (I9924,I9893,I227663);
nor I_412 (I9941,I9876,I227663);
nand I_413 (I9655,I9729,I9941);
nor I_414 (I9972,I9876,I9859);
nand I_415 (I9652,I9972,I227663);
not I_416 (I10003,I9859);
nor I_417 (I10020,I9763,I10003);
DFFARX1 I_418 (I10020,I2898,I9678,I9658,);
nor I_419 (I10051,I10003,I9746);
nor I_420 (I10068,I227648,I227669);
or I_421 (I10085,I10068,I227654);
nor I_422 (I10102,I227657,I227648);
nand I_423 (I10119,I10102,I10085);
not I_424 (I10136,I10119);
nor I_425 (I9640,I9893,I10136);
nand I_426 (I10167,I10136,I10051);
nand I_427 (I10184,I9893,I10167);
DFFARX1 I_428 (I10184,I2898,I9678,I9649,);
nor I_429 (I9667,I10136,I9924);
or I_430 (I9664,I10136,I9729);
nand I_431 (I9670,I9859,I10119);
not I_432 (I10290,I2905);
or I_433 (I10307,I343665,I343665);
nor I_434 (I10324,I343665,I343665);
nor I_435 (I10341,I10324,I343668);
nand I_436 (I10358,I10307,I343677);
not I_437 (I10375,I10358);
nor I_438 (I10392,I10341,I10375);
or I_439 (I10258,I10358,I343662);
nor I_440 (I10273,I10375,I343662);
and I_441 (I10437,I343659,I343668);
nor I_442 (I10454,I10437,I343671);
nand I_443 (I10471,I343659,I343656);
nor I_444 (I10488,I10471,I10454);
not I_445 (I10505,I10488);
nor I_446 (I10255,I10505,I10392);
nor I_447 (I10536,I10505,I343662);
nor I_448 (I10553,I10488,I343662);
nand I_449 (I10267,I10341,I10553);
nor I_450 (I10584,I10488,I10471);
nand I_451 (I10264,I10584,I343662);
not I_452 (I10615,I10471);
nor I_453 (I10632,I10375,I10615);
DFFARX1 I_454 (I10632,I2898,I10290,I10270,);
nor I_455 (I10663,I10615,I10358);
nor I_456 (I10680,I343662,I343656);
or I_457 (I10697,I10680,I343671);
nor I_458 (I10714,I343680,I343674);
nand I_459 (I10731,I10714,I10697);
not I_460 (I10748,I10731);
nor I_461 (I10252,I10505,I10748);
nand I_462 (I10779,I10748,I10663);
nand I_463 (I10796,I10505,I10779);
DFFARX1 I_464 (I10796,I2898,I10290,I10261,);
nor I_465 (I10279,I10748,I10536);
or I_466 (I10276,I10748,I10341);
nand I_467 (I10282,I10471,I10731);
not I_468 (I10902,I2905);
or I_469 (I10919,I21778,I21796);
nor I_470 (I10936,I21778,I21796);
nor I_471 (I10953,I10936,I21787);
nand I_472 (I10970,I10919,I21781);
not I_473 (I10987,I10970);
nor I_474 (I11004,I10953,I10987);
or I_475 (I10870,I10970,I21784);
nor I_476 (I10885,I10987,I21784);
and I_477 (I11049,I21799,I21781);
nor I_478 (I11066,I11049,I21790);
nand I_479 (I11083,I21793,I21787);
nor I_480 (I11100,I11083,I11066);
not I_481 (I11117,I11100);
nor I_482 (I10867,I11117,I11004);
nor I_483 (I11148,I11117,I21784);
nor I_484 (I11165,I11100,I21784);
nand I_485 (I10879,I10953,I11165);
nor I_486 (I11196,I11100,I11083);
nand I_487 (I10876,I11196,I21784);
not I_488 (I11227,I11083);
nor I_489 (I11244,I10987,I11227);
DFFARX1 I_490 (I11244,I2898,I10902,I10882,);
nor I_491 (I11275,I11227,I10970);
nor I_492 (I11292,I21784,I21790);
or I_493 (I11309,I11292,I21802);
nor I_494 (I11326,I21778,I21805);
nand I_495 (I11343,I11326,I11309);
not I_496 (I11360,I11343);
nor I_497 (I10864,I11117,I11360);
nand I_498 (I11391,I11360,I11275);
nand I_499 (I11408,I11117,I11391);
DFFARX1 I_500 (I11408,I2898,I10902,I10873,);
nor I_501 (I10891,I11360,I11148);
or I_502 (I10888,I11360,I10953);
nand I_503 (I10894,I11083,I11343);
not I_504 (I11514,I2905);
or I_505 (I11531,I191833,I191818);
nor I_506 (I11548,I191833,I191818);
nor I_507 (I11565,I11548,I191815);
nand I_508 (I11582,I11531,I191827);
not I_509 (I11599,I11582);
nor I_510 (I11616,I11565,I11599);
or I_511 (I11482,I11582,I191815);
nor I_512 (I11497,I11599,I191815);
and I_513 (I11661,I191824,I191836);
nor I_514 (I11678,I11661,I191821);
nand I_515 (I11695,I191830,I191827);
nor I_516 (I11712,I11695,I11678);
not I_517 (I11729,I11712);
nor I_518 (I11479,I11729,I11616);
nor I_519 (I11760,I11729,I191815);
nor I_520 (I11777,I11712,I191815);
nand I_521 (I11491,I11565,I11777);
nor I_522 (I11808,I11712,I11695);
nand I_523 (I11488,I11808,I191815);
not I_524 (I11839,I11695);
nor I_525 (I11856,I11599,I11839);
DFFARX1 I_526 (I11856,I2898,I11514,I11494,);
nor I_527 (I11887,I11839,I11582);
nor I_528 (I11904,I191818,I191824);
or I_529 (I11921,I11904,I191821);
nor I_530 (I11938,I191812,I191812);
nand I_531 (I11955,I11938,I11921);
not I_532 (I11972,I11955);
nor I_533 (I11476,I11729,I11972);
nand I_534 (I12003,I11972,I11887);
nand I_535 (I12020,I11729,I12003);
DFFARX1 I_536 (I12020,I2898,I11514,I11485,);
nor I_537 (I11503,I11972,I11760);
or I_538 (I11500,I11972,I11565);
nand I_539 (I11506,I11695,I11955);
not I_540 (I12126,I2905);
or I_541 (I12143,I324030,I324030);
nor I_542 (I12160,I324030,I324030);
nor I_543 (I12177,I12160,I324033);
nand I_544 (I12194,I12143,I324042);
not I_545 (I12211,I12194);
nor I_546 (I12228,I12177,I12211);
or I_547 (I12094,I12194,I324027);
nor I_548 (I12109,I12211,I324027);
and I_549 (I12273,I324024,I324033);
nor I_550 (I12290,I12273,I324036);
nand I_551 (I12307,I324024,I324021);
nor I_552 (I12324,I12307,I12290);
not I_553 (I12341,I12324);
nor I_554 (I12091,I12341,I12228);
nor I_555 (I12372,I12341,I324027);
nor I_556 (I12389,I12324,I324027);
nand I_557 (I12103,I12177,I12389);
nor I_558 (I12420,I12324,I12307);
nand I_559 (I12100,I12420,I324027);
not I_560 (I12451,I12307);
nor I_561 (I12468,I12211,I12451);
DFFARX1 I_562 (I12468,I2898,I12126,I12106,);
nor I_563 (I12499,I12451,I12194);
nor I_564 (I12516,I324027,I324021);
or I_565 (I12533,I12516,I324036);
nor I_566 (I12550,I324045,I324039);
nand I_567 (I12567,I12550,I12533);
not I_568 (I12584,I12567);
nor I_569 (I12088,I12341,I12584);
nand I_570 (I12615,I12584,I12499);
nand I_571 (I12632,I12341,I12615);
DFFARX1 I_572 (I12632,I2898,I12126,I12097,);
nor I_573 (I12115,I12584,I12372);
or I_574 (I12112,I12584,I12177);
nand I_575 (I12118,I12307,I12567);
not I_576 (I12738,I2905);
or I_577 (I12755,I341285,I341285);
nor I_578 (I12772,I341285,I341285);
nor I_579 (I12789,I12772,I341288);
nand I_580 (I12806,I12755,I341297);
not I_581 (I12823,I12806);
nor I_582 (I12840,I12789,I12823);
or I_583 (I12706,I12806,I341282);
nor I_584 (I12721,I12823,I341282);
and I_585 (I12885,I341279,I341288);
nor I_586 (I12902,I12885,I341291);
nand I_587 (I12919,I341279,I341276);
nor I_588 (I12936,I12919,I12902);
not I_589 (I12953,I12936);
nor I_590 (I12703,I12953,I12840);
nor I_591 (I12984,I12953,I341282);
nor I_592 (I13001,I12936,I341282);
nand I_593 (I12715,I12789,I13001);
nor I_594 (I13032,I12936,I12919);
nand I_595 (I12712,I13032,I341282);
not I_596 (I13063,I12919);
nor I_597 (I13080,I12823,I13063);
DFFARX1 I_598 (I13080,I2898,I12738,I12718,);
nor I_599 (I13111,I13063,I12806);
nor I_600 (I13128,I341282,I341276);
or I_601 (I13145,I13128,I341291);
nor I_602 (I13162,I341300,I341294);
nand I_603 (I13179,I13162,I13145);
not I_604 (I13196,I13179);
nor I_605 (I12700,I12953,I13196);
nand I_606 (I13227,I13196,I13111);
nand I_607 (I13244,I12953,I13227);
DFFARX1 I_608 (I13244,I2898,I12738,I12709,);
nor I_609 (I12727,I13196,I12984);
or I_610 (I12724,I13196,I12789);
nand I_611 (I12730,I12919,I13179);
not I_612 (I13350,I2905);
or I_613 (I13367,I44913,I44934);
nor I_614 (I13384,I44913,I44934);
nor I_615 (I13401,I13384,I44898);
nand I_616 (I13418,I13367,I44901);
not I_617 (I13435,I13418);
nor I_618 (I13452,I13401,I13435);
or I_619 (I13318,I13418,I44931);
nor I_620 (I13333,I13435,I44931);
and I_621 (I13497,I44904,I44910);
nor I_622 (I13514,I13497,I44928);
nand I_623 (I13531,I44916,I44925);
nor I_624 (I13548,I13531,I13514);
not I_625 (I13565,I13548);
nor I_626 (I13315,I13565,I13452);
nor I_627 (I13596,I13565,I44931);
nor I_628 (I13613,I13548,I44931);
nand I_629 (I13327,I13401,I13613);
nor I_630 (I13644,I13548,I13531);
nand I_631 (I13324,I13644,I44931);
not I_632 (I13675,I13531);
nor I_633 (I13692,I13435,I13675);
DFFARX1 I_634 (I13692,I2898,I13350,I13330,);
nor I_635 (I13723,I13675,I13418);
nor I_636 (I13740,I44907,I44901);
or I_637 (I13757,I13740,I44919);
nor I_638 (I13774,I44922,I44898);
nand I_639 (I13791,I13774,I13757);
not I_640 (I13808,I13791);
nor I_641 (I13312,I13565,I13808);
nand I_642 (I13839,I13808,I13723);
nand I_643 (I13856,I13565,I13839);
DFFARX1 I_644 (I13856,I2898,I13350,I13321,);
nor I_645 (I13339,I13808,I13596);
or I_646 (I13336,I13808,I13401);
nand I_647 (I13342,I13531,I13791);
not I_648 (I13959,I2905);
not I_649 (I13976,I400632);
nand I_650 (I13993,I400635,I400638);
nand I_651 (I14010,I13993,I400632);
not I_652 (I14027,I14010);
nand I_653 (I14044,I13993,I13976);
and I_654 (I14061,I14044,I400626);
nand I_655 (I14078,I14061,I400632);
not I_656 (I14095,I14078);
or I_657 (I14112,I400626,I400644);
nor I_658 (I14129,I14112,I400623);
not I_659 (I14146,I14129);
nor I_660 (I14163,I14010,I14146);
nor I_661 (I14180,I14095,I14163);
nor I_662 (I13927,I14180,I14163);
nand I_663 (I14211,I14146,I14078);
not I_664 (I14228,I400623);
nand I_665 (I14245,I14211,I14228);
nand I_666 (I14262,I400635,I400641);
not I_667 (I14279,I14262);
nand I_668 (I14296,I14279,I400623);
nor I_669 (I14313,I14279,I14027);
nor I_670 (I13924,I14262,I14245);
nand I_671 (I14344,I14027,I14262);
nand I_672 (I13951,I14296,I14344);
nor I_673 (I14375,I400647,I400629);
not I_674 (I14392,I400638);
nor I_675 (I14409,I14392,I400629);
nor I_676 (I14426,I14409,I400623);
and I_677 (I14443,I14279,I14426);
nor I_678 (I13942,I14443,I14129);
not I_679 (I14474,I14409);
or I_680 (I14491,I14474,I14180);
nor I_681 (I13930,I14010,I14491);
nor I_682 (I13948,I14313,I14474);
nor I_683 (I14536,I14375,I14392);
nor I_684 (I14553,I14279,I14536);
DFFARX1 I_685 (I14553,I2898,I13959,I13933,);
nor I_686 (I14584,I14536,I14095);
not I_687 (I13939,I14584);
or I_688 (I13945,I14536,I14129);
nor I_689 (I13936,I14409,I14536);
not I_690 (I14673,I2905);
not I_691 (I14690,I229919);
nand I_692 (I14707,I229895,I229907);
nand I_693 (I14724,I14707,I229919);
not I_694 (I14741,I14724);
nand I_695 (I14758,I14707,I14690);
and I_696 (I14775,I14758,I229895);
nand I_697 (I14792,I14775,I229892);
not I_698 (I14809,I14792);
or I_699 (I14826,I229916,I229898);
nor I_700 (I14843,I14826,I229910);
not I_701 (I14860,I14843);
nor I_702 (I14877,I14724,I14860);
nor I_703 (I14894,I14809,I14877);
nor I_704 (I14641,I14894,I14877);
nand I_705 (I14925,I14860,I14792);
not I_706 (I14942,I229901);
nand I_707 (I14959,I14925,I14942);
nand I_708 (I14976,I229892,I229904);
not I_709 (I14993,I14976);
nand I_710 (I15010,I14993,I229901);
nor I_711 (I15027,I14993,I14741);
nor I_712 (I14638,I14976,I14959);
nand I_713 (I15058,I14741,I14976);
nand I_714 (I14665,I15010,I15058);
nor I_715 (I15089,I229904,I229901);
not I_716 (I15106,I229913);
nor I_717 (I15123,I15106,I229898);
nor I_718 (I15140,I15123,I229901);
and I_719 (I15157,I14993,I15140);
nor I_720 (I14656,I15157,I14843);
not I_721 (I15188,I15123);
or I_722 (I15205,I15188,I14894);
nor I_723 (I14644,I14724,I15205);
nor I_724 (I14662,I15027,I15188);
nor I_725 (I15250,I15089,I15106);
nor I_726 (I15267,I14993,I15250);
DFFARX1 I_727 (I15267,I2898,I14673,I14647,);
nor I_728 (I15298,I15250,I14809);
not I_729 (I14653,I15298);
or I_730 (I14659,I15250,I14843);
nor I_731 (I14650,I15123,I15250);
not I_732 (I15387,I2905);
not I_733 (I15404,I438018);
nand I_734 (I15421,I438009,I438012);
nand I_735 (I15438,I15421,I438018);
not I_736 (I15455,I15438);
nand I_737 (I15472,I15421,I15404);
and I_738 (I15489,I15472,I438006);
nand I_739 (I15506,I15489,I438033);
not I_740 (I15523,I15506);
or I_741 (I15540,I438024,I438009);
nor I_742 (I15557,I15540,I438021);
not I_743 (I15574,I15557);
nor I_744 (I15591,I15438,I15574);
nor I_745 (I15608,I15523,I15591);
nor I_746 (I15355,I15608,I15591);
nand I_747 (I15639,I15574,I15506);
not I_748 (I15656,I438030);
nand I_749 (I15673,I15639,I15656);
nand I_750 (I15690,I438036,I438027);
not I_751 (I15707,I15690);
nand I_752 (I15724,I15707,I438030);
nor I_753 (I15741,I15707,I15455);
nor I_754 (I15352,I15690,I15673);
nand I_755 (I15772,I15455,I15690);
nand I_756 (I15379,I15724,I15772);
nor I_757 (I15803,I438015,I438039);
not I_758 (I15820,I438012);
nor I_759 (I15837,I15820,I438006);
nor I_760 (I15854,I15837,I438030);
and I_761 (I15871,I15707,I15854);
nor I_762 (I15370,I15871,I15557);
not I_763 (I15902,I15837);
or I_764 (I15919,I15902,I15608);
nor I_765 (I15358,I15438,I15919);
nor I_766 (I15376,I15741,I15902);
nor I_767 (I15964,I15803,I15820);
nor I_768 (I15981,I15707,I15964);
DFFARX1 I_769 (I15981,I2898,I15387,I15361,);
nor I_770 (I16012,I15964,I15523);
not I_771 (I15367,I16012);
or I_772 (I15373,I15964,I15557);
nor I_773 (I15364,I15837,I15964);
not I_774 (I16101,I2905);
not I_775 (I16118,I149086);
nand I_776 (I16135,I149098,I149104);
nand I_777 (I16152,I16135,I149086);
not I_778 (I16169,I16152);
nand I_779 (I16186,I16135,I16118);
and I_780 (I16203,I16186,I149077);
nand I_781 (I16220,I16203,I149101);
not I_782 (I16237,I16220);
or I_783 (I16254,I149083,I149074);
nor I_784 (I16271,I16254,I149092);
not I_785 (I16288,I16271);
nor I_786 (I16305,I16152,I16288);
nor I_787 (I16322,I16237,I16305);
nor I_788 (I16069,I16322,I16305);
nand I_789 (I16353,I16288,I16220);
not I_790 (I16370,I149095);
nand I_791 (I16387,I16353,I16370);
nand I_792 (I16404,I149080,I149077);
not I_793 (I16421,I16404);
nand I_794 (I16438,I16421,I149095);
nor I_795 (I16455,I16421,I16169);
nor I_796 (I16066,I16404,I16387);
nand I_797 (I16486,I16169,I16404);
nand I_798 (I16093,I16438,I16486);
nor I_799 (I16517,I149074,I149080);
not I_800 (I16534,I149107);
nor I_801 (I16551,I16534,I149089);
nor I_802 (I16568,I16551,I149095);
and I_803 (I16585,I16421,I16568);
nor I_804 (I16084,I16585,I16271);
not I_805 (I16616,I16551);
or I_806 (I16633,I16616,I16322);
nor I_807 (I16072,I16152,I16633);
nor I_808 (I16090,I16455,I16616);
nor I_809 (I16678,I16517,I16534);
nor I_810 (I16695,I16421,I16678);
DFFARX1 I_811 (I16695,I2898,I16101,I16075,);
nor I_812 (I16726,I16678,I16237);
not I_813 (I16081,I16726);
or I_814 (I16087,I16678,I16271);
nor I_815 (I16078,I16551,I16678);
not I_816 (I16815,I2905);
not I_817 (I16832,I353795);
nand I_818 (I16849,I353783,I353774);
nand I_819 (I16866,I16849,I353795);
not I_820 (I16883,I16866);
nand I_821 (I16900,I16849,I16832);
and I_822 (I16917,I16900,I353783);
nand I_823 (I16934,I16917,I353789);
not I_824 (I16951,I16934);
or I_825 (I16968,I353771,I353780);
nor I_826 (I16985,I16968,I353786);
not I_827 (I17002,I16985);
nor I_828 (I17019,I16866,I17002);
nor I_829 (I17036,I16951,I17019);
nor I_830 (I16783,I17036,I17019);
nand I_831 (I17067,I17002,I16934);
not I_832 (I17084,I353780);
nand I_833 (I17101,I17067,I17084);
nand I_834 (I17118,I353774,I353771);
not I_835 (I17135,I17118);
nand I_836 (I17152,I17135,I353780);
nor I_837 (I17169,I17135,I16883);
nor I_838 (I16780,I17118,I17101);
nand I_839 (I17200,I16883,I17118);
nand I_840 (I16807,I17152,I17200);
nor I_841 (I17231,I353786,I353777);
not I_842 (I17248,I353792);
nor I_843 (I17265,I17248,I353777);
nor I_844 (I17282,I17265,I353780);
and I_845 (I17299,I17135,I17282);
nor I_846 (I16798,I17299,I16985);
not I_847 (I17330,I17265);
or I_848 (I17347,I17330,I17036);
nor I_849 (I16786,I16866,I17347);
nor I_850 (I16804,I17169,I17330);
nor I_851 (I17392,I17231,I17248);
nor I_852 (I17409,I17135,I17392);
DFFARX1 I_853 (I17409,I2898,I16815,I16789,);
nor I_854 (I17440,I17392,I16951);
not I_855 (I16795,I17440);
or I_856 (I16801,I17392,I16985);
nor I_857 (I16792,I17265,I17392);
not I_858 (I17529,I2905);
not I_859 (I17546,I383585);
nand I_860 (I17563,I383567,I383558);
nand I_861 (I17580,I17563,I383585);
not I_862 (I17597,I17580);
nand I_863 (I17614,I17563,I17546);
and I_864 (I17631,I17614,I383579);
nand I_865 (I17648,I17631,I383588);
not I_866 (I17665,I17648);
or I_867 (I17682,I383555,I383555);
nor I_868 (I17699,I17682,I383561);
not I_869 (I17716,I17699);
nor I_870 (I17733,I17580,I17716);
nor I_871 (I17750,I17665,I17733);
nor I_872 (I17497,I17750,I17733);
nand I_873 (I17781,I17716,I17648);
not I_874 (I17798,I383564);
nand I_875 (I17815,I17781,I17798);
nand I_876 (I17832,I383582,I383573);
not I_877 (I17849,I17832);
nand I_878 (I17866,I17849,I383564);
nor I_879 (I17883,I17849,I17597);
nor I_880 (I17494,I17832,I17815);
nand I_881 (I17914,I17597,I17832);
nand I_882 (I17521,I17866,I17914);
nor I_883 (I17945,I383558,I383570);
not I_884 (I17962,I383561);
nor I_885 (I17979,I17962,I383576);
nor I_886 (I17996,I17979,I383564);
and I_887 (I18013,I17849,I17996);
nor I_888 (I17512,I18013,I17699);
not I_889 (I18044,I17979);
or I_890 (I18061,I18044,I17750);
nor I_891 (I17500,I17580,I18061);
nor I_892 (I17518,I17883,I18044);
nor I_893 (I18106,I17945,I17962);
nor I_894 (I18123,I17849,I18106);
DFFARX1 I_895 (I18123,I2898,I17529,I17503,);
nor I_896 (I18154,I18106,I17665);
not I_897 (I17509,I18154);
or I_898 (I17515,I18106,I17699);
nor I_899 (I17506,I17979,I18106);
not I_900 (I18243,I2905);
not I_901 (I18260,I45680);
nand I_902 (I18277,I45701,I45680);
nand I_903 (I18294,I18277,I45680);
not I_904 (I18311,I18294);
nand I_905 (I18328,I18277,I18260);
and I_906 (I18345,I18328,I45695);
nand I_907 (I18362,I18345,I45707);
not I_908 (I18379,I18362);
or I_909 (I18396,I45683,I45698);
nor I_910 (I18413,I18396,I45692);
not I_911 (I18430,I18413);
nor I_912 (I18447,I18294,I18430);
nor I_913 (I18464,I18379,I18447);
nor I_914 (I18211,I18464,I18447);
nand I_915 (I18495,I18430,I18362);
not I_916 (I18512,I45704);
nand I_917 (I18529,I18495,I18512);
nand I_918 (I18546,I45686,I45710);
not I_919 (I18563,I18546);
nand I_920 (I18580,I18563,I45704);
nor I_921 (I18597,I18563,I18311);
nor I_922 (I18208,I18546,I18529);
nand I_923 (I18628,I18311,I18546);
nand I_924 (I18235,I18580,I18628);
nor I_925 (I18659,I45689,I45683);
not I_926 (I18676,I45713);
nor I_927 (I18693,I18676,I45716);
nor I_928 (I18710,I18693,I45704);
and I_929 (I18727,I18563,I18710);
nor I_930 (I18226,I18727,I18413);
not I_931 (I18758,I18693);
or I_932 (I18775,I18758,I18464);
nor I_933 (I18214,I18294,I18775);
nor I_934 (I18232,I18597,I18758);
nor I_935 (I18820,I18659,I18676);
nor I_936 (I18837,I18563,I18820);
DFFARX1 I_937 (I18837,I2898,I18243,I18217,);
nor I_938 (I18868,I18820,I18379);
not I_939 (I18223,I18868);
or I_940 (I18229,I18820,I18413);
nor I_941 (I18220,I18693,I18820);
not I_942 (I18957,I2905);
not I_943 (I18974,I200882);
nand I_944 (I18991,I200888,I200873);
nand I_945 (I19008,I18991,I200882);
not I_946 (I19025,I19008);
nand I_947 (I19042,I18991,I18974);
and I_948 (I19059,I19042,I200873);
nand I_949 (I19076,I19059,I200891);
not I_950 (I19093,I19076);
or I_951 (I19110,I200885,I200879);
nor I_952 (I19127,I19110,I200876);
not I_953 (I19144,I19127);
nor I_954 (I19161,I19008,I19144);
nor I_955 (I19178,I19093,I19161);
nor I_956 (I18925,I19178,I19161);
nand I_957 (I19209,I19144,I19076);
not I_958 (I19226,I200876);
nand I_959 (I19243,I19209,I19226);
nand I_960 (I19260,I200879,I200897);
not I_961 (I19277,I19260);
nand I_962 (I19294,I19277,I200876);
nor I_963 (I19311,I19277,I19025);
nor I_964 (I18922,I19260,I19243);
nand I_965 (I19342,I19025,I19260);
nand I_966 (I18949,I19294,I19342);
nor I_967 (I19373,I200882,I200894);
not I_968 (I19390,I200888);
nor I_969 (I19407,I19390,I200885);
nor I_970 (I19424,I19407,I200876);
and I_971 (I19441,I19277,I19424);
nor I_972 (I18940,I19441,I19127);
not I_973 (I19472,I19407);
or I_974 (I19489,I19472,I19178);
nor I_975 (I18928,I19008,I19489);
nor I_976 (I18946,I19311,I19472);
nor I_977 (I19534,I19373,I19390);
nor I_978 (I19551,I19277,I19534);
DFFARX1 I_979 (I19551,I2898,I18957,I18931,);
nor I_980 (I19582,I19534,I19093);
not I_981 (I18937,I19582);
or I_982 (I18943,I19534,I19127);
nor I_983 (I18934,I19407,I19534);
not I_984 (I19671,I2905);
not I_985 (I19688,I382939);
nand I_986 (I19705,I382921,I382912);
nand I_987 (I19722,I19705,I382939);
not I_988 (I19739,I19722);
nand I_989 (I19756,I19705,I19688);
and I_990 (I19773,I19756,I382933);
nand I_991 (I19790,I19773,I382942);
not I_992 (I19807,I19790);
or I_993 (I19824,I382909,I382909);
nor I_994 (I19841,I19824,I382915);
not I_995 (I19858,I19841);
nor I_996 (I19875,I19722,I19858);
nor I_997 (I19892,I19807,I19875);
nor I_998 (I19639,I19892,I19875);
nand I_999 (I19923,I19858,I19790);
not I_1000 (I19940,I382918);
nand I_1001 (I19957,I19923,I19940);
nand I_1002 (I19974,I382936,I382927);
not I_1003 (I19991,I19974);
nand I_1004 (I20008,I19991,I382918);
nor I_1005 (I20025,I19991,I19739);
nor I_1006 (I19636,I19974,I19957);
nand I_1007 (I20056,I19739,I19974);
nand I_1008 (I19663,I20008,I20056);
nor I_1009 (I20087,I382912,I382924);
not I_1010 (I20104,I382915);
nor I_1011 (I20121,I20104,I382930);
nor I_1012 (I20138,I20121,I382918);
and I_1013 (I20155,I19991,I20138);
nor I_1014 (I19654,I20155,I19841);
not I_1015 (I20186,I20121);
or I_1016 (I20203,I20186,I19892);
nor I_1017 (I19642,I19722,I20203);
nor I_1018 (I19660,I20025,I20186);
nor I_1019 (I20248,I20087,I20104);
nor I_1020 (I20265,I19991,I20248);
DFFARX1 I_1021 (I20265,I2898,I19671,I19645,);
nor I_1022 (I20296,I20248,I19807);
not I_1023 (I19651,I20296);
or I_1024 (I19657,I20248,I19841);
nor I_1025 (I19648,I20121,I20248);
not I_1026 (I20385,I2905);
not I_1027 (I20402,I321520);
nand I_1028 (I20419,I321535,I321505);
nand I_1029 (I20436,I20419,I321520);
not I_1030 (I20453,I20436);
nand I_1031 (I20470,I20419,I20402);
and I_1032 (I20487,I20470,I321517);
nand I_1033 (I20504,I20487,I321508);
not I_1034 (I20521,I20504);
or I_1035 (I20538,I321529,I321532);
nor I_1036 (I20555,I20538,I321511);
not I_1037 (I20572,I20555);
nor I_1038 (I20589,I20436,I20572);
nor I_1039 (I20606,I20521,I20589);
nor I_1040 (I20353,I20606,I20589);
nand I_1041 (I20637,I20572,I20504);
not I_1042 (I20654,I321514);
nand I_1043 (I20671,I20637,I20654);
nand I_1044 (I20688,I321505,I321508);
not I_1045 (I20705,I20688);
nand I_1046 (I20722,I20705,I321514);
nor I_1047 (I20739,I20705,I20453);
nor I_1048 (I20350,I20688,I20671);
nand I_1049 (I20770,I20453,I20688);
nand I_1050 (I20377,I20722,I20770);
nor I_1051 (I20801,I321514,I321526);
not I_1052 (I20818,I321523);
nor I_1053 (I20835,I20818,I321511);
nor I_1054 (I20852,I20835,I321514);
and I_1055 (I20869,I20705,I20852);
nor I_1056 (I20368,I20869,I20555);
not I_1057 (I20900,I20835);
or I_1058 (I20917,I20900,I20606);
nor I_1059 (I20356,I20436,I20917);
nor I_1060 (I20374,I20739,I20900);
nor I_1061 (I20962,I20801,I20818);
nor I_1062 (I20979,I20705,I20962);
DFFARX1 I_1063 (I20979,I2898,I20385,I20359,);
nor I_1064 (I21010,I20962,I20521);
not I_1065 (I20365,I21010);
or I_1066 (I20371,I20962,I20555);
nor I_1067 (I20362,I20835,I20962);
not I_1068 (I21099,I2905);
not I_1069 (I21116,I143697);
nand I_1070 (I21133,I143703,I143688);
nand I_1071 (I21150,I21133,I143697);
not I_1072 (I21167,I21150);
nand I_1073 (I21184,I21133,I21116);
and I_1074 (I21201,I21184,I143715);
nand I_1075 (I21218,I21201,I143685);
not I_1076 (I21235,I21218);
or I_1077 (I21252,I143694,I143706);
nor I_1078 (I21269,I21252,I143691);
not I_1079 (I21286,I21269);
nor I_1080 (I21303,I21150,I21286);
nor I_1081 (I21320,I21235,I21303);
nor I_1082 (I21067,I21320,I21303);
nand I_1083 (I21351,I21286,I21218);
not I_1084 (I21368,I143709);
nand I_1085 (I21385,I21351,I21368);
nand I_1086 (I21402,I143700,I143688);
not I_1087 (I21419,I21402);
nand I_1088 (I21436,I21419,I143709);
nor I_1089 (I21453,I21419,I21167);
nor I_1090 (I21064,I21402,I21385);
nand I_1091 (I21484,I21167,I21402);
nand I_1092 (I21091,I21436,I21484);
nor I_1093 (I21515,I143718,I143691);
not I_1094 (I21532,I143712);
nor I_1095 (I21549,I21532,I143685);
nor I_1096 (I21566,I21549,I143709);
and I_1097 (I21583,I21419,I21566);
nor I_1098 (I21082,I21583,I21269);
not I_1099 (I21614,I21549);
or I_1100 (I21631,I21614,I21320);
nor I_1101 (I21070,I21150,I21631);
nor I_1102 (I21088,I21453,I21614);
nor I_1103 (I21676,I21515,I21532);
nor I_1104 (I21693,I21419,I21676);
DFFARX1 I_1105 (I21693,I2898,I21099,I21073,);
nor I_1106 (I21724,I21676,I21235);
not I_1107 (I21079,I21724);
or I_1108 (I21085,I21676,I21269);
nor I_1109 (I21076,I21549,I21676);
not I_1110 (I21813,I2905);
not I_1111 (I21830,I328210);
nand I_1112 (I21847,I328198,I328189);
nand I_1113 (I21864,I21847,I328210);
not I_1114 (I21881,I21864);
nand I_1115 (I21898,I21847,I21830);
and I_1116 (I21915,I21898,I328198);
nand I_1117 (I21932,I21915,I328204);
not I_1118 (I21949,I21932);
or I_1119 (I21966,I328186,I328195);
nor I_1120 (I21983,I21966,I328201);
not I_1121 (I22000,I21983);
nor I_1122 (I22017,I21864,I22000);
nor I_1123 (I22034,I21949,I22017);
nor I_1124 (I21781,I22034,I22017);
nand I_1125 (I22065,I22000,I21932);
not I_1126 (I22082,I328195);
nand I_1127 (I22099,I22065,I22082);
nand I_1128 (I22116,I328189,I328186);
not I_1129 (I22133,I22116);
nand I_1130 (I22150,I22133,I328195);
nor I_1131 (I22167,I22133,I21881);
nor I_1132 (I21778,I22116,I22099);
nand I_1133 (I22198,I21881,I22116);
nand I_1134 (I21805,I22150,I22198);
nor I_1135 (I22229,I328201,I328192);
not I_1136 (I22246,I328207);
nor I_1137 (I22263,I22246,I328192);
nor I_1138 (I22280,I22263,I328195);
and I_1139 (I22297,I22133,I22280);
nor I_1140 (I21796,I22297,I21983);
not I_1141 (I22328,I22263);
or I_1142 (I22345,I22328,I22034);
nor I_1143 (I21784,I21864,I22345);
nor I_1144 (I21802,I22167,I22328);
nor I_1145 (I22390,I22229,I22246);
nor I_1146 (I22407,I22133,I22390);
DFFARX1 I_1147 (I22407,I2898,I21813,I21787,);
nor I_1148 (I22438,I22390,I21949);
not I_1149 (I21793,I22438);
or I_1150 (I21799,I22390,I21983);
nor I_1151 (I21790,I22263,I22390);
not I_1152 (I22527,I2905);
not I_1153 (I22544,I116021);
nand I_1154 (I22561,I116027,I116012);
nand I_1155 (I22578,I22561,I116021);
not I_1156 (I22595,I22578);
nand I_1157 (I22612,I22561,I22544);
and I_1158 (I22629,I22612,I116039);
nand I_1159 (I22646,I22629,I116009);
not I_1160 (I22663,I22646);
or I_1161 (I22680,I116018,I116030);
nor I_1162 (I22697,I22680,I116015);
not I_1163 (I22714,I22697);
nor I_1164 (I22731,I22578,I22714);
nor I_1165 (I22748,I22663,I22731);
nor I_1166 (I22495,I22748,I22731);
nand I_1167 (I22779,I22714,I22646);
not I_1168 (I22796,I116033);
nand I_1169 (I22813,I22779,I22796);
nand I_1170 (I22830,I116024,I116012);
not I_1171 (I22847,I22830);
nand I_1172 (I22864,I22847,I116033);
nor I_1173 (I22881,I22847,I22595);
nor I_1174 (I22492,I22830,I22813);
nand I_1175 (I22912,I22595,I22830);
nand I_1176 (I22519,I22864,I22912);
nor I_1177 (I22943,I116042,I116015);
not I_1178 (I22960,I116036);
nor I_1179 (I22977,I22960,I116009);
nor I_1180 (I22994,I22977,I116033);
and I_1181 (I23011,I22847,I22994);
nor I_1182 (I22510,I23011,I22697);
not I_1183 (I23042,I22977);
or I_1184 (I23059,I23042,I22748);
nor I_1185 (I22498,I22578,I23059);
nor I_1186 (I22516,I22881,I23042);
nor I_1187 (I23104,I22943,I22960);
nor I_1188 (I23121,I22847,I23104);
DFFARX1 I_1189 (I23121,I2898,I22527,I22501,);
nor I_1190 (I23152,I23104,I22663);
not I_1191 (I22507,I23152);
or I_1192 (I22513,I23104,I22697);
nor I_1193 (I22504,I22977,I23104);
not I_1194 (I23241,I2905);
not I_1195 (I23258,I48808);
nand I_1196 (I23275,I48829,I48808);
nand I_1197 (I23292,I23275,I48808);
not I_1198 (I23309,I23292);
nand I_1199 (I23326,I23275,I23258);
and I_1200 (I23343,I23326,I48823);
nand I_1201 (I23360,I23343,I48835);
not I_1202 (I23377,I23360);
or I_1203 (I23394,I48811,I48826);
nor I_1204 (I23411,I23394,I48820);
not I_1205 (I23428,I23411);
nor I_1206 (I23445,I23292,I23428);
nor I_1207 (I23462,I23377,I23445);
nor I_1208 (I23209,I23462,I23445);
nand I_1209 (I23493,I23428,I23360);
not I_1210 (I23510,I48832);
nand I_1211 (I23527,I23493,I23510);
nand I_1212 (I23544,I48814,I48838);
not I_1213 (I23561,I23544);
nand I_1214 (I23578,I23561,I48832);
nor I_1215 (I23595,I23561,I23309);
nor I_1216 (I23206,I23544,I23527);
nand I_1217 (I23626,I23309,I23544);
nand I_1218 (I23233,I23578,I23626);
nor I_1219 (I23657,I48817,I48811);
not I_1220 (I23674,I48841);
nor I_1221 (I23691,I23674,I48844);
nor I_1222 (I23708,I23691,I48832);
and I_1223 (I23725,I23561,I23708);
nor I_1224 (I23224,I23725,I23411);
not I_1225 (I23756,I23691);
or I_1226 (I23773,I23756,I23462);
nor I_1227 (I23212,I23292,I23773);
nor I_1228 (I23230,I23595,I23756);
nor I_1229 (I23818,I23657,I23674);
nor I_1230 (I23835,I23561,I23818);
DFFARX1 I_1231 (I23835,I2898,I23241,I23215,);
nor I_1232 (I23866,I23818,I23377);
not I_1233 (I23221,I23866);
or I_1234 (I23227,I23818,I23411);
nor I_1235 (I23218,I23691,I23818);
not I_1236 (I23955,I2905);
not I_1237 (I23972,I179105);
nand I_1238 (I23989,I179102,I179114);
nand I_1239 (I24006,I23989,I179105);
not I_1240 (I24023,I24006);
nand I_1241 (I24040,I23989,I23972);
and I_1242 (I24057,I24040,I179123);
nand I_1243 (I24074,I24057,I179120);
not I_1244 (I24091,I24074);
or I_1245 (I24108,I179099,I179096);
nor I_1246 (I24125,I24108,I179117);
not I_1247 (I24142,I24125);
nor I_1248 (I24159,I24006,I24142);
nor I_1249 (I24176,I24091,I24159);
nor I_1250 (I23923,I24176,I24159);
nand I_1251 (I24207,I24142,I24074);
not I_1252 (I24224,I179108);
nand I_1253 (I24241,I24207,I24224);
nand I_1254 (I24258,I179102,I179126);
not I_1255 (I24275,I24258);
nand I_1256 (I24292,I24275,I179108);
nor I_1257 (I24309,I24275,I24023);
nor I_1258 (I23920,I24258,I24241);
nand I_1259 (I24340,I24023,I24258);
nand I_1260 (I23947,I24292,I24340);
nor I_1261 (I24371,I179096,I179099);
not I_1262 (I24388,I179111);
nor I_1263 (I24405,I24388,I179105);
nor I_1264 (I24422,I24405,I179108);
and I_1265 (I24439,I24275,I24422);
nor I_1266 (I23938,I24439,I24125);
not I_1267 (I24470,I24405);
or I_1268 (I24487,I24470,I24176);
nor I_1269 (I23926,I24006,I24487);
nor I_1270 (I23944,I24309,I24470);
nor I_1271 (I24532,I24371,I24388);
nor I_1272 (I24549,I24275,I24532);
DFFARX1 I_1273 (I24549,I2898,I23955,I23929,);
nor I_1274 (I24580,I24532,I24091);
not I_1275 (I23935,I24580);
or I_1276 (I23941,I24532,I24125);
nor I_1277 (I23932,I24405,I24532);
not I_1278 (I24669,I2905);
not I_1279 (I24686,I363309);
nand I_1280 (I24703,I363318,I363315);
nand I_1281 (I24720,I24703,I363309);
not I_1282 (I24737,I24720);
nand I_1283 (I24754,I24703,I24686);
and I_1284 (I24771,I24754,I363324);
nand I_1285 (I24788,I24771,I363303);
not I_1286 (I24805,I24788);
or I_1287 (I24822,I363291,I363297);
nor I_1288 (I24839,I24822,I363294);
not I_1289 (I24856,I24839);
nor I_1290 (I24873,I24720,I24856);
nor I_1291 (I24890,I24805,I24873);
nor I_1292 (I24637,I24890,I24873);
nand I_1293 (I24921,I24856,I24788);
not I_1294 (I24938,I363294);
nand I_1295 (I24955,I24921,I24938);
nand I_1296 (I24972,I363321,I363306);
not I_1297 (I24989,I24972);
nand I_1298 (I25006,I24989,I363294);
nor I_1299 (I25023,I24989,I24737);
nor I_1300 (I24634,I24972,I24955);
nand I_1301 (I25054,I24737,I24972);
nand I_1302 (I24661,I25006,I25054);
nor I_1303 (I25085,I363300,I363297);
not I_1304 (I25102,I363291);
nor I_1305 (I25119,I25102,I363312);
nor I_1306 (I25136,I25119,I363294);
and I_1307 (I25153,I24989,I25136);
nor I_1308 (I24652,I25153,I24839);
not I_1309 (I25184,I25119);
or I_1310 (I25201,I25184,I24890);
nor I_1311 (I24640,I24720,I25201);
nor I_1312 (I24658,I25023,I25184);
nor I_1313 (I25246,I25085,I25102);
nor I_1314 (I25263,I24989,I25246);
DFFARX1 I_1315 (I25263,I2898,I24669,I24643,);
nor I_1316 (I25294,I25246,I24805);
not I_1317 (I24649,I25294);
or I_1318 (I24655,I25246,I24839);
nor I_1319 (I24646,I25119,I25246);
not I_1320 (I25383,I2905);
not I_1321 (I25400,I97202);
nand I_1322 (I25417,I97193,I97190);
nand I_1323 (I25434,I25417,I97202);
not I_1324 (I25451,I25434);
nand I_1325 (I25468,I25417,I25400);
and I_1326 (I25485,I25468,I97199);
nand I_1327 (I25502,I25485,I97199);
not I_1328 (I25519,I25502);
or I_1329 (I25536,I97202,I97214);
nor I_1330 (I25553,I25536,I97205);
not I_1331 (I25570,I25553);
nor I_1332 (I25587,I25434,I25570);
nor I_1333 (I25604,I25519,I25587);
nor I_1334 (I25351,I25604,I25587);
nand I_1335 (I25635,I25570,I25502);
not I_1336 (I25652,I97193);
nand I_1337 (I25669,I25635,I25652);
nand I_1338 (I25686,I97217,I97196);
not I_1339 (I25703,I25686);
nand I_1340 (I25720,I25703,I97193);
nor I_1341 (I25737,I25703,I25451);
nor I_1342 (I25348,I25686,I25669);
nand I_1343 (I25768,I25451,I25686);
nand I_1344 (I25375,I25720,I25768);
nor I_1345 (I25799,I97196,I97190);
not I_1346 (I25816,I97211);
nor I_1347 (I25833,I25816,I97208);
nor I_1348 (I25850,I25833,I97193);
and I_1349 (I25867,I25703,I25850);
nor I_1350 (I25366,I25867,I25553);
not I_1351 (I25898,I25833);
or I_1352 (I25915,I25898,I25604);
nor I_1353 (I25354,I25434,I25915);
nor I_1354 (I25372,I25737,I25898);
nor I_1355 (I25960,I25799,I25816);
nor I_1356 (I25977,I25703,I25960);
DFFARX1 I_1357 (I25977,I2898,I25383,I25357,);
nor I_1358 (I26008,I25960,I25519);
not I_1359 (I25363,I26008);
or I_1360 (I25369,I25960,I25553);
nor I_1361 (I25360,I25833,I25960);
not I_1362 (I26097,I2905);
not I_1363 (I26114,I165406);
nand I_1364 (I26131,I165418,I165424);
nand I_1365 (I26148,I26131,I165406);
not I_1366 (I26165,I26148);
nand I_1367 (I26182,I26131,I26114);
and I_1368 (I26199,I26182,I165397);
nand I_1369 (I26216,I26199,I165421);
not I_1370 (I26233,I26216);
or I_1371 (I26250,I165403,I165394);
nor I_1372 (I26267,I26250,I165412);
not I_1373 (I26284,I26267);
nor I_1374 (I26301,I26148,I26284);
nor I_1375 (I26318,I26233,I26301);
nor I_1376 (I26065,I26318,I26301);
nand I_1377 (I26349,I26284,I26216);
not I_1378 (I26366,I165415);
nand I_1379 (I26383,I26349,I26366);
nand I_1380 (I26400,I165400,I165397);
not I_1381 (I26417,I26400);
nand I_1382 (I26434,I26417,I165415);
nor I_1383 (I26451,I26417,I26165);
nor I_1384 (I26062,I26400,I26383);
nand I_1385 (I26482,I26165,I26400);
nand I_1386 (I26089,I26434,I26482);
nor I_1387 (I26513,I165394,I165400);
not I_1388 (I26530,I165427);
nor I_1389 (I26547,I26530,I165409);
nor I_1390 (I26564,I26547,I165415);
and I_1391 (I26581,I26417,I26564);
nor I_1392 (I26080,I26581,I26267);
not I_1393 (I26612,I26547);
or I_1394 (I26629,I26612,I26318);
nor I_1395 (I26068,I26148,I26629);
nor I_1396 (I26086,I26451,I26612);
nor I_1397 (I26674,I26513,I26530);
nor I_1398 (I26691,I26417,I26674);
DFFARX1 I_1399 (I26691,I2898,I26097,I26071,);
nor I_1400 (I26722,I26674,I26233);
not I_1401 (I26077,I26722);
or I_1402 (I26083,I26674,I26267);
nor I_1403 (I26074,I26547,I26674);
not I_1404 (I26811,I2905);
not I_1405 (I26828,I434533);
nand I_1406 (I26845,I434524,I434527);
nand I_1407 (I26862,I26845,I434533);
not I_1408 (I26879,I26862);
nand I_1409 (I26896,I26845,I26828);
and I_1410 (I26913,I26896,I434521);
nand I_1411 (I26930,I26913,I434548);
not I_1412 (I26947,I26930);
or I_1413 (I26964,I434539,I434524);
nor I_1414 (I26981,I26964,I434536);
not I_1415 (I26998,I26981);
nor I_1416 (I27015,I26862,I26998);
nor I_1417 (I27032,I26947,I27015);
nor I_1418 (I26779,I27032,I27015);
nand I_1419 (I27063,I26998,I26930);
not I_1420 (I27080,I434545);
nand I_1421 (I27097,I27063,I27080);
nand I_1422 (I27114,I434551,I434542);
not I_1423 (I27131,I27114);
nand I_1424 (I27148,I27131,I434545);
nor I_1425 (I27165,I27131,I26879);
nor I_1426 (I26776,I27114,I27097);
nand I_1427 (I27196,I26879,I27114);
nand I_1428 (I26803,I27148,I27196);
nor I_1429 (I27227,I434530,I434554);
not I_1430 (I27244,I434527);
nor I_1431 (I27261,I27244,I434521);
nor I_1432 (I27278,I27261,I434545);
and I_1433 (I27295,I27131,I27278);
nor I_1434 (I26794,I27295,I26981);
not I_1435 (I27326,I27261);
or I_1436 (I27343,I27326,I27032);
nor I_1437 (I26782,I26862,I27343);
nor I_1438 (I26800,I27165,I27326);
nor I_1439 (I27388,I27227,I27244);
nor I_1440 (I27405,I27131,I27388);
DFFARX1 I_1441 (I27405,I2898,I26811,I26785,);
nor I_1442 (I27436,I27388,I26947);
not I_1443 (I26791,I27436);
or I_1444 (I26797,I27388,I26981);
nor I_1445 (I26788,I27261,I27388);
not I_1446 (I27525,I2905);
not I_1447 (I27542,I5371);
nand I_1448 (I27559,I5362,I5356);
nand I_1449 (I27576,I27559,I5371);
not I_1450 (I27593,I27576);
nand I_1451 (I27610,I27559,I27542);
and I_1452 (I27627,I27610,I5365);
nand I_1453 (I27644,I27627,I5368);
not I_1454 (I27661,I27644);
or I_1455 (I27678,I5377,I5359);
nor I_1456 (I27695,I27678,I5380);
not I_1457 (I27712,I27695);
nor I_1458 (I27729,I27576,I27712);
nor I_1459 (I27746,I27661,I27729);
nor I_1460 (I27493,I27746,I27729);
nand I_1461 (I27777,I27712,I27644);
not I_1462 (I27794,I5359);
nand I_1463 (I27811,I27777,I27794);
nand I_1464 (I27828,I5383,I5362);
not I_1465 (I27845,I27828);
nand I_1466 (I27862,I27845,I5359);
nor I_1467 (I27879,I27845,I27593);
nor I_1468 (I27490,I27828,I27811);
nand I_1469 (I27910,I27593,I27828);
nand I_1470 (I27517,I27862,I27910);
nor I_1471 (I27941,I5356,I5365);
not I_1472 (I27958,I5374);
nor I_1473 (I27975,I27958,I5386);
nor I_1474 (I27992,I27975,I5359);
and I_1475 (I28009,I27845,I27992);
nor I_1476 (I27508,I28009,I27695);
not I_1477 (I28040,I27975);
or I_1478 (I28057,I28040,I27746);
nor I_1479 (I27496,I27576,I28057);
nor I_1480 (I27514,I27879,I28040);
nor I_1481 (I28102,I27941,I27958);
nor I_1482 (I28119,I27845,I28102);
DFFARX1 I_1483 (I28119,I2898,I27525,I27499,);
nor I_1484 (I28150,I28102,I27661);
not I_1485 (I27505,I28150);
or I_1486 (I27511,I28102,I27695);
nor I_1487 (I27502,I27975,I28102);
not I_1488 (I28239,I2905);
not I_1489 (I28256,I65752);
nand I_1490 (I28273,I65743,I65740);
nand I_1491 (I28290,I28273,I65752);
not I_1492 (I28307,I28290);
nand I_1493 (I28324,I28273,I28256);
and I_1494 (I28341,I28324,I65749);
nand I_1495 (I28358,I28341,I65749);
not I_1496 (I28375,I28358);
or I_1497 (I28392,I65752,I65764);
nor I_1498 (I28409,I28392,I65755);
not I_1499 (I28426,I28409);
nor I_1500 (I28443,I28290,I28426);
nor I_1501 (I28460,I28375,I28443);
nor I_1502 (I28207,I28460,I28443);
nand I_1503 (I28491,I28426,I28358);
not I_1504 (I28508,I65743);
nand I_1505 (I28525,I28491,I28508);
nand I_1506 (I28542,I65767,I65746);
not I_1507 (I28559,I28542);
nand I_1508 (I28576,I28559,I65743);
nor I_1509 (I28593,I28559,I28307);
nor I_1510 (I28204,I28542,I28525);
nand I_1511 (I28624,I28307,I28542);
nand I_1512 (I28231,I28576,I28624);
nor I_1513 (I28655,I65746,I65740);
not I_1514 (I28672,I65761);
nor I_1515 (I28689,I28672,I65758);
nor I_1516 (I28706,I28689,I65743);
and I_1517 (I28723,I28559,I28706);
nor I_1518 (I28222,I28723,I28409);
not I_1519 (I28754,I28689);
or I_1520 (I28771,I28754,I28460);
nor I_1521 (I28210,I28290,I28771);
nor I_1522 (I28228,I28593,I28754);
nor I_1523 (I28816,I28655,I28672);
nor I_1524 (I28833,I28559,I28816);
DFFARX1 I_1525 (I28833,I2898,I28239,I28213,);
nor I_1526 (I28864,I28816,I28375);
not I_1527 (I28219,I28864);
or I_1528 (I28225,I28816,I28409);
nor I_1529 (I28216,I28689,I28816);
not I_1530 (I28953,I2905);
not I_1531 (I28970,I162686);
nand I_1532 (I28987,I162698,I162704);
nand I_1533 (I29004,I28987,I162686);
not I_1534 (I29021,I29004);
nand I_1535 (I29038,I28987,I28970);
and I_1536 (I29055,I29038,I162677);
nand I_1537 (I29072,I29055,I162701);
not I_1538 (I29089,I29072);
or I_1539 (I29106,I162683,I162674);
nor I_1540 (I29123,I29106,I162692);
not I_1541 (I29140,I29123);
nor I_1542 (I29157,I29004,I29140);
nor I_1543 (I29174,I29089,I29157);
nor I_1544 (I28921,I29174,I29157);
nand I_1545 (I29205,I29140,I29072);
not I_1546 (I29222,I162695);
nand I_1547 (I29239,I29205,I29222);
nand I_1548 (I29256,I162680,I162677);
not I_1549 (I29273,I29256);
nand I_1550 (I29290,I29273,I162695);
nor I_1551 (I29307,I29273,I29021);
nor I_1552 (I28918,I29256,I29239);
nand I_1553 (I29338,I29021,I29256);
nand I_1554 (I28945,I29290,I29338);
nor I_1555 (I29369,I162674,I162680);
not I_1556 (I29386,I162707);
nor I_1557 (I29403,I29386,I162689);
nor I_1558 (I29420,I29403,I162695);
and I_1559 (I29437,I29273,I29420);
nor I_1560 (I28936,I29437,I29123);
not I_1561 (I29468,I29403);
or I_1562 (I29485,I29468,I29174);
nor I_1563 (I28924,I29004,I29485);
nor I_1564 (I28942,I29307,I29468);
nor I_1565 (I29530,I29369,I29386);
nor I_1566 (I29547,I29273,I29530);
DFFARX1 I_1567 (I29547,I2898,I28953,I28927,);
nor I_1568 (I29578,I29530,I29089);
not I_1569 (I28933,I29578);
or I_1570 (I28939,I29530,I29123);
nor I_1571 (I28930,I29403,I29530);
not I_1572 (I29667,I2905);
not I_1573 (I29684,I300321);
nand I_1574 (I29701,I300336,I300306);
nand I_1575 (I29718,I29701,I300321);
not I_1576 (I29735,I29718);
nand I_1577 (I29752,I29701,I29684);
and I_1578 (I29769,I29752,I300318);
nand I_1579 (I29786,I29769,I300309);
not I_1580 (I29803,I29786);
or I_1581 (I29820,I300330,I300333);
nor I_1582 (I29837,I29820,I300312);
not I_1583 (I29854,I29837);
nor I_1584 (I29871,I29718,I29854);
nor I_1585 (I29888,I29803,I29871);
nor I_1586 (I29635,I29888,I29871);
nand I_1587 (I29919,I29854,I29786);
not I_1588 (I29936,I300315);
nand I_1589 (I29953,I29919,I29936);
nand I_1590 (I29970,I300306,I300309);
not I_1591 (I29987,I29970);
nand I_1592 (I30004,I29987,I300315);
nor I_1593 (I30021,I29987,I29735);
nor I_1594 (I29632,I29970,I29953);
nand I_1595 (I30052,I29735,I29970);
nand I_1596 (I29659,I30004,I30052);
nor I_1597 (I30083,I300315,I300327);
not I_1598 (I30100,I300324);
nor I_1599 (I30117,I30100,I300312);
nor I_1600 (I30134,I30117,I300315);
and I_1601 (I30151,I29987,I30134);
nor I_1602 (I29650,I30151,I29837);
not I_1603 (I30182,I30117);
or I_1604 (I30199,I30182,I29888);
nor I_1605 (I29638,I29718,I30199);
nor I_1606 (I29656,I30021,I30182);
nor I_1607 (I30244,I30083,I30100);
nor I_1608 (I30261,I29987,I30244);
DFFARX1 I_1609 (I30261,I2898,I29667,I29641,);
nor I_1610 (I30292,I30244,I29803);
not I_1611 (I29647,I30292);
or I_1612 (I29653,I30244,I29837);
nor I_1613 (I29644,I30117,I30244);
not I_1614 (I30381,I2905);
not I_1615 (I30398,I339515);
nand I_1616 (I30415,I339503,I339494);
nand I_1617 (I30432,I30415,I339515);
not I_1618 (I30449,I30432);
nand I_1619 (I30466,I30415,I30398);
and I_1620 (I30483,I30466,I339503);
nand I_1621 (I30500,I30483,I339509);
not I_1622 (I30517,I30500);
or I_1623 (I30534,I339491,I339500);
nor I_1624 (I30551,I30534,I339506);
not I_1625 (I30568,I30551);
nor I_1626 (I30585,I30432,I30568);
nor I_1627 (I30602,I30517,I30585);
nor I_1628 (I30349,I30602,I30585);
nand I_1629 (I30633,I30568,I30500);
not I_1630 (I30650,I339500);
nand I_1631 (I30667,I30633,I30650);
nand I_1632 (I30684,I339494,I339491);
not I_1633 (I30701,I30684);
nand I_1634 (I30718,I30701,I339500);
nor I_1635 (I30735,I30701,I30449);
nor I_1636 (I30346,I30684,I30667);
nand I_1637 (I30766,I30449,I30684);
nand I_1638 (I30373,I30718,I30766);
nor I_1639 (I30797,I339506,I339497);
not I_1640 (I30814,I339512);
nor I_1641 (I30831,I30814,I339497);
nor I_1642 (I30848,I30831,I339500);
and I_1643 (I30865,I30701,I30848);
nor I_1644 (I30364,I30865,I30551);
not I_1645 (I30896,I30831);
or I_1646 (I30913,I30896,I30602);
nor I_1647 (I30352,I30432,I30913);
nor I_1648 (I30370,I30735,I30896);
nor I_1649 (I30958,I30797,I30814);
nor I_1650 (I30975,I30701,I30958);
DFFARX1 I_1651 (I30975,I2898,I30381,I30355,);
nor I_1652 (I31006,I30958,I30517);
not I_1653 (I30361,I31006);
or I_1654 (I30367,I30958,I30551);
nor I_1655 (I30358,I30831,I30958);
not I_1656 (I31095,I2905);
not I_1657 (I31112,I245190);
nand I_1658 (I31129,I245184,I245196);
nand I_1659 (I31146,I31129,I245190);
not I_1660 (I31163,I31146);
nand I_1661 (I31180,I31129,I31112);
and I_1662 (I31197,I31180,I245202);
nand I_1663 (I31214,I31197,I245178);
not I_1664 (I31231,I31214);
or I_1665 (I31248,I245187,I245175);
nor I_1666 (I31265,I31248,I245181);
not I_1667 (I31282,I31265);
nor I_1668 (I31299,I31146,I31282);
nor I_1669 (I31316,I31231,I31299);
nor I_1670 (I31063,I31316,I31299);
nand I_1671 (I31347,I31282,I31214);
not I_1672 (I31364,I245205);
nand I_1673 (I31381,I31347,I31364);
nand I_1674 (I31398,I245175,I245178);
not I_1675 (I31415,I31398);
nand I_1676 (I31432,I31415,I245205);
nor I_1677 (I31449,I31415,I31163);
nor I_1678 (I31060,I31398,I31381);
nand I_1679 (I31480,I31163,I31398);
nand I_1680 (I31087,I31432,I31480);
nor I_1681 (I31511,I245181,I245193);
not I_1682 (I31528,I245199);
nor I_1683 (I31545,I31528,I245184);
nor I_1684 (I31562,I31545,I245205);
and I_1685 (I31579,I31415,I31562);
nor I_1686 (I31078,I31579,I31265);
not I_1687 (I31610,I31545);
or I_1688 (I31627,I31610,I31316);
nor I_1689 (I31066,I31146,I31627);
nor I_1690 (I31084,I31449,I31610);
nor I_1691 (I31672,I31511,I31528);
nor I_1692 (I31689,I31415,I31672);
DFFARX1 I_1693 (I31689,I2898,I31095,I31069,);
nor I_1694 (I31720,I31672,I31231);
not I_1695 (I31075,I31720);
or I_1696 (I31081,I31672,I31265);
nor I_1697 (I31072,I31545,I31672);
not I_1698 (I31809,I2905);
not I_1699 (I31826,I51936);
nand I_1700 (I31843,I51957,I51936);
nand I_1701 (I31860,I31843,I51936);
not I_1702 (I31877,I31860);
nand I_1703 (I31894,I31843,I31826);
and I_1704 (I31911,I31894,I51951);
nand I_1705 (I31928,I31911,I51963);
not I_1706 (I31945,I31928);
or I_1707 (I31962,I51939,I51954);
nor I_1708 (I31979,I31962,I51948);
not I_1709 (I31996,I31979);
nor I_1710 (I32013,I31860,I31996);
nor I_1711 (I32030,I31945,I32013);
nor I_1712 (I31777,I32030,I32013);
nand I_1713 (I32061,I31996,I31928);
not I_1714 (I32078,I51960);
nand I_1715 (I32095,I32061,I32078);
nand I_1716 (I32112,I51942,I51966);
not I_1717 (I32129,I32112);
nand I_1718 (I32146,I32129,I51960);
nor I_1719 (I32163,I32129,I31877);
nor I_1720 (I31774,I32112,I32095);
nand I_1721 (I32194,I31877,I32112);
nand I_1722 (I31801,I32146,I32194);
nor I_1723 (I32225,I51945,I51939);
not I_1724 (I32242,I51969);
nor I_1725 (I32259,I32242,I51972);
nor I_1726 (I32276,I32259,I51960);
and I_1727 (I32293,I32129,I32276);
nor I_1728 (I31792,I32293,I31979);
not I_1729 (I32324,I32259);
or I_1730 (I32341,I32324,I32030);
nor I_1731 (I31780,I31860,I32341);
nor I_1732 (I31798,I32163,I32324);
nor I_1733 (I32386,I32225,I32242);
nor I_1734 (I32403,I32129,I32386);
DFFARX1 I_1735 (I32403,I2898,I31809,I31783,);
nor I_1736 (I32434,I32386,I31945);
not I_1737 (I31789,I32434);
or I_1738 (I31795,I32386,I31979);
nor I_1739 (I31786,I32259,I32386);
not I_1740 (I32523,I2905);
not I_1741 (I32540,I241365);
nand I_1742 (I32557,I241359,I241371);
nand I_1743 (I32574,I32557,I241365);
not I_1744 (I32591,I32574);
nand I_1745 (I32608,I32557,I32540);
and I_1746 (I32625,I32608,I241377);
nand I_1747 (I32642,I32625,I241353);
not I_1748 (I32659,I32642);
or I_1749 (I32676,I241362,I241350);
nor I_1750 (I32693,I32676,I241356);
not I_1751 (I32710,I32693);
nor I_1752 (I32727,I32574,I32710);
nor I_1753 (I32744,I32659,I32727);
nor I_1754 (I32491,I32744,I32727);
nand I_1755 (I32775,I32710,I32642);
not I_1756 (I32792,I241380);
nand I_1757 (I32809,I32775,I32792);
nand I_1758 (I32826,I241350,I241353);
not I_1759 (I32843,I32826);
nand I_1760 (I32860,I32843,I241380);
nor I_1761 (I32877,I32843,I32591);
nor I_1762 (I32488,I32826,I32809);
nand I_1763 (I32908,I32591,I32826);
nand I_1764 (I32515,I32860,I32908);
nor I_1765 (I32939,I241356,I241368);
not I_1766 (I32956,I241374);
nor I_1767 (I32973,I32956,I241359);
nor I_1768 (I32990,I32973,I241380);
and I_1769 (I33007,I32843,I32990);
nor I_1770 (I32506,I33007,I32693);
not I_1771 (I33038,I32973);
or I_1772 (I33055,I33038,I32744);
nor I_1773 (I32494,I32574,I33055);
nor I_1774 (I32512,I32877,I33038);
nor I_1775 (I33100,I32939,I32956);
nor I_1776 (I33117,I32843,I33100);
DFFARX1 I_1777 (I33117,I2898,I32523,I32497,);
nor I_1778 (I33148,I33100,I32659);
not I_1779 (I32503,I33148);
or I_1780 (I32509,I33100,I32693);
nor I_1781 (I32500,I32973,I33100);
not I_1782 (I33237,I2905);
not I_1783 (I33254,I88396);
nand I_1784 (I33271,I88387,I88384);
nand I_1785 (I33288,I33271,I88396);
not I_1786 (I33305,I33288);
nand I_1787 (I33322,I33271,I33254);
and I_1788 (I33339,I33322,I88393);
nand I_1789 (I33356,I33339,I88393);
not I_1790 (I33373,I33356);
or I_1791 (I33390,I88396,I88408);
nor I_1792 (I33407,I33390,I88399);
not I_1793 (I33424,I33407);
nor I_1794 (I33441,I33288,I33424);
nor I_1795 (I33458,I33373,I33441);
nor I_1796 (I33205,I33458,I33441);
nand I_1797 (I33489,I33424,I33356);
not I_1798 (I33506,I88387);
nand I_1799 (I33523,I33489,I33506);
nand I_1800 (I33540,I88411,I88390);
not I_1801 (I33557,I33540);
nand I_1802 (I33574,I33557,I88387);
nor I_1803 (I33591,I33557,I33305);
nor I_1804 (I33202,I33540,I33523);
nand I_1805 (I33622,I33305,I33540);
nand I_1806 (I33229,I33574,I33622);
nor I_1807 (I33653,I88390,I88384);
not I_1808 (I33670,I88405);
nor I_1809 (I33687,I33670,I88402);
nor I_1810 (I33704,I33687,I88387);
and I_1811 (I33721,I33557,I33704);
nor I_1812 (I33220,I33721,I33407);
not I_1813 (I33752,I33687);
or I_1814 (I33769,I33752,I33458);
nor I_1815 (I33208,I33288,I33769);
nor I_1816 (I33226,I33591,I33752);
nor I_1817 (I33814,I33653,I33670);
nor I_1818 (I33831,I33557,I33814);
DFFARX1 I_1819 (I33831,I2898,I33237,I33211,);
nor I_1820 (I33862,I33814,I33373);
not I_1821 (I33217,I33862);
or I_1822 (I33223,I33814,I33407);
nor I_1823 (I33214,I33687,I33814);
not I_1824 (I33951,I2905);
not I_1825 (I33968,I359150);
nand I_1826 (I33985,I359138,I359129);
nand I_1827 (I34002,I33985,I359150);
not I_1828 (I34019,I34002);
nand I_1829 (I34036,I33985,I33968);
and I_1830 (I34053,I34036,I359138);
nand I_1831 (I34070,I34053,I359144);
not I_1832 (I34087,I34070);
or I_1833 (I34104,I359126,I359135);
nor I_1834 (I34121,I34104,I359141);
not I_1835 (I34138,I34121);
nor I_1836 (I34155,I34002,I34138);
nor I_1837 (I34172,I34087,I34155);
nor I_1838 (I33919,I34172,I34155);
nand I_1839 (I34203,I34138,I34070);
not I_1840 (I34220,I359135);
nand I_1841 (I34237,I34203,I34220);
nand I_1842 (I34254,I359129,I359126);
not I_1843 (I34271,I34254);
nand I_1844 (I34288,I34271,I359135);
nor I_1845 (I34305,I34271,I34019);
nor I_1846 (I33916,I34254,I34237);
nand I_1847 (I34336,I34019,I34254);
nand I_1848 (I33943,I34288,I34336);
nor I_1849 (I34367,I359141,I359132);
not I_1850 (I34384,I359147);
nor I_1851 (I34401,I34384,I359132);
nor I_1852 (I34418,I34401,I359135);
and I_1853 (I34435,I34271,I34418);
nor I_1854 (I33934,I34435,I34121);
not I_1855 (I34466,I34401);
or I_1856 (I34483,I34466,I34172);
nor I_1857 (I33922,I34002,I34483);
nor I_1858 (I33940,I34305,I34466);
nor I_1859 (I34528,I34367,I34384);
nor I_1860 (I34545,I34271,I34528);
DFFARX1 I_1861 (I34545,I2898,I33951,I33925,);
nor I_1862 (I34576,I34528,I34087);
not I_1863 (I33931,I34576);
or I_1864 (I33937,I34528,I34121);
nor I_1865 (I33928,I34401,I34528);
not I_1866 (I34665,I2905);
not I_1867 (I34682,I107215);
nand I_1868 (I34699,I107221,I107206);
nand I_1869 (I34716,I34699,I107215);
not I_1870 (I34733,I34716);
nand I_1871 (I34750,I34699,I34682);
and I_1872 (I34767,I34750,I107233);
nand I_1873 (I34784,I34767,I107203);
not I_1874 (I34801,I34784);
or I_1875 (I34818,I107212,I107224);
nor I_1876 (I34835,I34818,I107209);
not I_1877 (I34852,I34835);
nor I_1878 (I34869,I34716,I34852);
nor I_1879 (I34886,I34801,I34869);
nor I_1880 (I34633,I34886,I34869);
nand I_1881 (I34917,I34852,I34784);
not I_1882 (I34934,I107227);
nand I_1883 (I34951,I34917,I34934);
nand I_1884 (I34968,I107218,I107206);
not I_1885 (I34985,I34968);
nand I_1886 (I35002,I34985,I107227);
nor I_1887 (I35019,I34985,I34733);
nor I_1888 (I34630,I34968,I34951);
nand I_1889 (I35050,I34733,I34968);
nand I_1890 (I34657,I35002,I35050);
nor I_1891 (I35081,I107236,I107209);
not I_1892 (I35098,I107230);
nor I_1893 (I35115,I35098,I107203);
nor I_1894 (I35132,I35115,I107227);
and I_1895 (I35149,I34985,I35132);
nor I_1896 (I34648,I35149,I34835);
not I_1897 (I35180,I35115);
or I_1898 (I35197,I35180,I34886);
nor I_1899 (I34636,I34716,I35197);
nor I_1900 (I34654,I35019,I35180);
nor I_1901 (I35242,I35081,I35098);
nor I_1902 (I35259,I34985,I35242);
DFFARX1 I_1903 (I35259,I2898,I34665,I34639,);
nor I_1904 (I35290,I35242,I34801);
not I_1905 (I34645,I35290);
or I_1906 (I34651,I35242,I34835);
nor I_1907 (I34642,I35115,I35242);
not I_1908 (I35379,I2905);
not I_1909 (I35396,I252840);
nand I_1910 (I35413,I252834,I252846);
nand I_1911 (I35430,I35413,I252840);
not I_1912 (I35447,I35430);
nand I_1913 (I35464,I35413,I35396);
and I_1914 (I35481,I35464,I252852);
nand I_1915 (I35498,I35481,I252828);
not I_1916 (I35515,I35498);
or I_1917 (I35532,I252837,I252825);
nor I_1918 (I35549,I35532,I252831);
not I_1919 (I35566,I35549);
nor I_1920 (I35583,I35430,I35566);
nor I_1921 (I35600,I35515,I35583);
nor I_1922 (I35347,I35600,I35583);
nand I_1923 (I35631,I35566,I35498);
not I_1924 (I35648,I252855);
nand I_1925 (I35665,I35631,I35648);
nand I_1926 (I35682,I252825,I252828);
not I_1927 (I35699,I35682);
nand I_1928 (I35716,I35699,I252855);
nor I_1929 (I35733,I35699,I35447);
nor I_1930 (I35344,I35682,I35665);
nand I_1931 (I35764,I35447,I35682);
nand I_1932 (I35371,I35716,I35764);
nor I_1933 (I35795,I252831,I252843);
not I_1934 (I35812,I252849);
nor I_1935 (I35829,I35812,I252834);
nor I_1936 (I35846,I35829,I252855);
and I_1937 (I35863,I35699,I35846);
nor I_1938 (I35362,I35863,I35549);
not I_1939 (I35894,I35829);
or I_1940 (I35911,I35894,I35600);
nor I_1941 (I35350,I35430,I35911);
nor I_1942 (I35368,I35733,I35894);
nor I_1943 (I35956,I35795,I35812);
nor I_1944 (I35973,I35699,I35956);
DFFARX1 I_1945 (I35973,I2898,I35379,I35353,);
nor I_1946 (I36004,I35956,I35515);
not I_1947 (I35359,I36004);
or I_1948 (I35365,I35956,I35549);
nor I_1949 (I35356,I35829,I35956);
not I_1950 (I36093,I2905);
not I_1951 (I36110,I236775);
nand I_1952 (I36127,I236769,I236781);
nand I_1953 (I36144,I36127,I236775);
not I_1954 (I36161,I36144);
nand I_1955 (I36178,I36127,I36110);
and I_1956 (I36195,I36178,I236787);
nand I_1957 (I36212,I36195,I236763);
not I_1958 (I36229,I36212);
or I_1959 (I36246,I236772,I236760);
nor I_1960 (I36263,I36246,I236766);
not I_1961 (I36280,I36263);
nor I_1962 (I36297,I36144,I36280);
nor I_1963 (I36314,I36229,I36297);
nor I_1964 (I36061,I36314,I36297);
nand I_1965 (I36345,I36280,I36212);
not I_1966 (I36362,I236790);
nand I_1967 (I36379,I36345,I36362);
nand I_1968 (I36396,I236760,I236763);
not I_1969 (I36413,I36396);
nand I_1970 (I36430,I36413,I236790);
nor I_1971 (I36447,I36413,I36161);
nor I_1972 (I36058,I36396,I36379);
nand I_1973 (I36478,I36161,I36396);
nand I_1974 (I36085,I36430,I36478);
nor I_1975 (I36509,I236766,I236778);
not I_1976 (I36526,I236784);
nor I_1977 (I36543,I36526,I236769);
nor I_1978 (I36560,I36543,I236790);
and I_1979 (I36577,I36413,I36560);
nor I_1980 (I36076,I36577,I36263);
not I_1981 (I36608,I36543);
or I_1982 (I36625,I36608,I36314);
nor I_1983 (I36064,I36144,I36625);
nor I_1984 (I36082,I36447,I36608);
nor I_1985 (I36670,I36509,I36526);
nor I_1986 (I36687,I36413,I36670);
DFFARX1 I_1987 (I36687,I2898,I36093,I36067,);
nor I_1988 (I36718,I36670,I36229);
not I_1989 (I36073,I36718);
or I_1990 (I36079,I36670,I36263);
nor I_1991 (I36070,I36543,I36670);
not I_1992 (I36807,I2905);
not I_1993 (I36824,I330590);
nand I_1994 (I36841,I330578,I330569);
nand I_1995 (I36858,I36841,I330590);
not I_1996 (I36875,I36858);
nand I_1997 (I36892,I36841,I36824);
and I_1998 (I36909,I36892,I330578);
nand I_1999 (I36926,I36909,I330584);
not I_2000 (I36943,I36926);
or I_2001 (I36960,I330566,I330575);
nor I_2002 (I36977,I36960,I330581);
not I_2003 (I36994,I36977);
nor I_2004 (I37011,I36858,I36994);
nor I_2005 (I37028,I36943,I37011);
nor I_2006 (I36775,I37028,I37011);
nand I_2007 (I37059,I36994,I36926);
not I_2008 (I37076,I330575);
nand I_2009 (I37093,I37059,I37076);
nand I_2010 (I37110,I330569,I330566);
not I_2011 (I37127,I37110);
nand I_2012 (I37144,I37127,I330575);
nor I_2013 (I37161,I37127,I36875);
nor I_2014 (I36772,I37110,I37093);
nand I_2015 (I37192,I36875,I37110);
nand I_2016 (I36799,I37144,I37192);
nor I_2017 (I37223,I330581,I330572);
not I_2018 (I37240,I330587);
nor I_2019 (I37257,I37240,I330572);
nor I_2020 (I37274,I37257,I330575);
and I_2021 (I37291,I37127,I37274);
nor I_2022 (I36790,I37291,I36977);
not I_2023 (I37322,I37257);
or I_2024 (I37339,I37322,I37028);
nor I_2025 (I36778,I36858,I37339);
nor I_2026 (I36796,I37161,I37322);
nor I_2027 (I37384,I37223,I37240);
nor I_2028 (I37401,I37127,I37384);
DFFARX1 I_2029 (I37401,I2898,I36807,I36781,);
nor I_2030 (I37432,I37384,I36943);
not I_2031 (I36787,I37432);
or I_2032 (I36793,I37384,I36977);
nor I_2033 (I36784,I37257,I37384);
not I_2034 (I37521,I2905);
not I_2035 (I37538,I164726);
nand I_2036 (I37555,I164738,I164744);
nand I_2037 (I37572,I37555,I164726);
not I_2038 (I37589,I37572);
nand I_2039 (I37606,I37555,I37538);
and I_2040 (I37623,I37606,I164717);
nand I_2041 (I37640,I37623,I164741);
not I_2042 (I37657,I37640);
or I_2043 (I37674,I164723,I164714);
nor I_2044 (I37691,I37674,I164732);
not I_2045 (I37708,I37691);
nor I_2046 (I37725,I37572,I37708);
nor I_2047 (I37742,I37657,I37725);
nor I_2048 (I37489,I37742,I37725);
nand I_2049 (I37773,I37708,I37640);
not I_2050 (I37790,I164735);
nand I_2051 (I37807,I37773,I37790);
nand I_2052 (I37824,I164720,I164717);
not I_2053 (I37841,I37824);
nand I_2054 (I37858,I37841,I164735);
nor I_2055 (I37875,I37841,I37589);
nor I_2056 (I37486,I37824,I37807);
nand I_2057 (I37906,I37589,I37824);
nand I_2058 (I37513,I37858,I37906);
nor I_2059 (I37937,I164714,I164720);
not I_2060 (I37954,I164747);
nor I_2061 (I37971,I37954,I164729);
nor I_2062 (I37988,I37971,I164735);
and I_2063 (I38005,I37841,I37988);
nor I_2064 (I37504,I38005,I37691);
not I_2065 (I38036,I37971);
or I_2066 (I38053,I38036,I37742);
nor I_2067 (I37492,I37572,I38053);
nor I_2068 (I37510,I37875,I38036);
nor I_2069 (I38098,I37937,I37954);
nor I_2070 (I38115,I37841,I38098);
DFFARX1 I_2071 (I38115,I2898,I37521,I37495,);
nor I_2072 (I38146,I38098,I37657);
not I_2073 (I37501,I38146);
or I_2074 (I37507,I38098,I37691);
nor I_2075 (I37498,I37971,I38098);
not I_2076 (I38235,I2905);
not I_2077 (I38252,I324640);
nand I_2078 (I38269,I324628,I324619);
nand I_2079 (I38286,I38269,I324640);
not I_2080 (I38303,I38286);
nand I_2081 (I38320,I38269,I38252);
and I_2082 (I38337,I38320,I324628);
nand I_2083 (I38354,I38337,I324634);
not I_2084 (I38371,I38354);
or I_2085 (I38388,I324616,I324625);
nor I_2086 (I38405,I38388,I324631);
not I_2087 (I38422,I38405);
nor I_2088 (I38439,I38286,I38422);
nor I_2089 (I38456,I38371,I38439);
nor I_2090 (I38203,I38456,I38439);
nand I_2091 (I38487,I38422,I38354);
not I_2092 (I38504,I324625);
nand I_2093 (I38521,I38487,I38504);
nand I_2094 (I38538,I324619,I324616);
not I_2095 (I38555,I38538);
nand I_2096 (I38572,I38555,I324625);
nor I_2097 (I38589,I38555,I38303);
nor I_2098 (I38200,I38538,I38521);
nand I_2099 (I38620,I38303,I38538);
nand I_2100 (I38227,I38572,I38620);
nor I_2101 (I38651,I324631,I324622);
not I_2102 (I38668,I324637);
nor I_2103 (I38685,I38668,I324622);
nor I_2104 (I38702,I38685,I324625);
and I_2105 (I38719,I38555,I38702);
nor I_2106 (I38218,I38719,I38405);
not I_2107 (I38750,I38685);
or I_2108 (I38767,I38750,I38456);
nor I_2109 (I38206,I38286,I38767);
nor I_2110 (I38224,I38589,I38750);
nor I_2111 (I38812,I38651,I38668);
nor I_2112 (I38829,I38555,I38812);
DFFARX1 I_2113 (I38829,I2898,I38235,I38209,);
nor I_2114 (I38860,I38812,I38371);
not I_2115 (I38215,I38860);
or I_2116 (I38221,I38812,I38405);
nor I_2117 (I38212,I38685,I38812);
not I_2118 (I38949,I2905);
not I_2119 (I38966,I309093);
nand I_2120 (I38983,I309108,I309078);
nand I_2121 (I39000,I38983,I309093);
not I_2122 (I39017,I39000);
nand I_2123 (I39034,I38983,I38966);
and I_2124 (I39051,I39034,I309090);
nand I_2125 (I39068,I39051,I309081);
not I_2126 (I39085,I39068);
or I_2127 (I39102,I309102,I309105);
nor I_2128 (I39119,I39102,I309084);
not I_2129 (I39136,I39119);
nor I_2130 (I39153,I39000,I39136);
nor I_2131 (I39170,I39085,I39153);
nor I_2132 (I38917,I39170,I39153);
nand I_2133 (I39201,I39136,I39068);
not I_2134 (I39218,I309087);
nand I_2135 (I39235,I39201,I39218);
nand I_2136 (I39252,I309078,I309081);
not I_2137 (I39269,I39252);
nand I_2138 (I39286,I39269,I309087);
nor I_2139 (I39303,I39269,I39017);
nor I_2140 (I38914,I39252,I39235);
nand I_2141 (I39334,I39017,I39252);
nand I_2142 (I38941,I39286,I39334);
nor I_2143 (I39365,I309087,I309099);
not I_2144 (I39382,I309096);
nor I_2145 (I39399,I39382,I309084);
nor I_2146 (I39416,I39399,I309087);
and I_2147 (I39433,I39269,I39416);
nor I_2148 (I38932,I39433,I39119);
not I_2149 (I39464,I39399);
or I_2150 (I39481,I39464,I39170);
nor I_2151 (I38920,I39000,I39481);
nor I_2152 (I38938,I39303,I39464);
nor I_2153 (I39526,I39365,I39382);
nor I_2154 (I39543,I39269,I39526);
DFFARX1 I_2155 (I39543,I2898,I38949,I38923,);
nor I_2156 (I39574,I39526,I39085);
not I_2157 (I38929,I39574);
or I_2158 (I38935,I39526,I39119);
nor I_2159 (I38926,I39399,I39526);
not I_2160 (I39663,I2905);
not I_2161 (I39680,I373249);
nand I_2162 (I39697,I373231,I373222);
nand I_2163 (I39714,I39697,I373249);
not I_2164 (I39731,I39714);
nand I_2165 (I39748,I39697,I39680);
and I_2166 (I39765,I39748,I373243);
nand I_2167 (I39782,I39765,I373252);
not I_2168 (I39799,I39782);
or I_2169 (I39816,I373219,I373219);
nor I_2170 (I39833,I39816,I373225);
not I_2171 (I39850,I39833);
nor I_2172 (I39867,I39714,I39850);
nor I_2173 (I39884,I39799,I39867);
nor I_2174 (I39631,I39884,I39867);
nand I_2175 (I39915,I39850,I39782);
not I_2176 (I39932,I373228);
nand I_2177 (I39949,I39915,I39932);
nand I_2178 (I39966,I373246,I373237);
not I_2179 (I39983,I39966);
nand I_2180 (I40000,I39983,I373228);
nor I_2181 (I40017,I39983,I39731);
nor I_2182 (I39628,I39966,I39949);
nand I_2183 (I40048,I39731,I39966);
nand I_2184 (I39655,I40000,I40048);
nor I_2185 (I40079,I373222,I373234);
not I_2186 (I40096,I373225);
nor I_2187 (I40113,I40096,I373240);
nor I_2188 (I40130,I40113,I373228);
and I_2189 (I40147,I39983,I40130);
nor I_2190 (I39646,I40147,I39833);
not I_2191 (I40178,I40113);
or I_2192 (I40195,I40178,I39884);
nor I_2193 (I39634,I39714,I40195);
nor I_2194 (I39652,I40017,I40178);
nor I_2195 (I40240,I40079,I40096);
nor I_2196 (I40257,I39983,I40240);
DFFARX1 I_2197 (I40257,I2898,I39663,I39637,);
nor I_2198 (I40288,I40240,I39799);
not I_2199 (I39643,I40288);
or I_2200 (I39649,I40240,I39833);
nor I_2201 (I39640,I40113,I40240);
not I_2202 (I40377,I2905);
not I_2203 (I40394,I199488);
nand I_2204 (I40411,I199494,I199479);
nand I_2205 (I40428,I40411,I199488);
not I_2206 (I40445,I40428);
nand I_2207 (I40462,I40411,I40394);
and I_2208 (I40479,I40462,I199479);
nand I_2209 (I40496,I40479,I199497);
not I_2210 (I40513,I40496);
or I_2211 (I40530,I199491,I199485);
nor I_2212 (I40547,I40530,I199482);
not I_2213 (I40564,I40547);
nor I_2214 (I40581,I40428,I40564);
nor I_2215 (I40598,I40513,I40581);
nor I_2216 (I40345,I40598,I40581);
nand I_2217 (I40629,I40564,I40496);
not I_2218 (I40646,I199482);
nand I_2219 (I40663,I40629,I40646);
nand I_2220 (I40680,I199485,I199503);
not I_2221 (I40697,I40680);
nand I_2222 (I40714,I40697,I199482);
nor I_2223 (I40731,I40697,I40445);
nor I_2224 (I40342,I40680,I40663);
nand I_2225 (I40762,I40445,I40680);
nand I_2226 (I40369,I40714,I40762);
nor I_2227 (I40793,I199488,I199500);
not I_2228 (I40810,I199494);
nor I_2229 (I40827,I40810,I199491);
nor I_2230 (I40844,I40827,I199482);
and I_2231 (I40861,I40697,I40844);
nor I_2232 (I40360,I40861,I40547);
not I_2233 (I40892,I40827);
or I_2234 (I40909,I40892,I40598);
nor I_2235 (I40348,I40428,I40909);
nor I_2236 (I40366,I40731,I40892);
nor I_2237 (I40954,I40793,I40810);
nor I_2238 (I40971,I40697,I40954);
DFFARX1 I_2239 (I40971,I2898,I40377,I40351,);
nor I_2240 (I41002,I40954,I40513);
not I_2241 (I40357,I41002);
or I_2242 (I40363,I40954,I40547);
nor I_2243 (I40354,I40827,I40954);
not I_2244 (I41091,I2905);
not I_2245 (I41108,I211967);
nand I_2246 (I41125,I211943,I211955);
nand I_2247 (I41142,I41125,I211967);
not I_2248 (I41159,I41142);
nand I_2249 (I41176,I41125,I41108);
and I_2250 (I41193,I41176,I211943);
nand I_2251 (I41210,I41193,I211940);
not I_2252 (I41227,I41210);
or I_2253 (I41244,I211964,I211946);
nor I_2254 (I41261,I41244,I211958);
not I_2255 (I41278,I41261);
nor I_2256 (I41295,I41142,I41278);
nor I_2257 (I41312,I41227,I41295);
nor I_2258 (I41059,I41312,I41295);
nand I_2259 (I41343,I41278,I41210);
not I_2260 (I41360,I211949);
nand I_2261 (I41377,I41343,I41360);
nand I_2262 (I41394,I211940,I211952);
not I_2263 (I41411,I41394);
nand I_2264 (I41428,I41411,I211949);
nor I_2265 (I41445,I41411,I41159);
nor I_2266 (I41056,I41394,I41377);
nand I_2267 (I41476,I41159,I41394);
nand I_2268 (I41083,I41428,I41476);
nor I_2269 (I41507,I211952,I211949);
not I_2270 (I41524,I211961);
nor I_2271 (I41541,I41524,I211946);
nor I_2272 (I41558,I41541,I211949);
and I_2273 (I41575,I41411,I41558);
nor I_2274 (I41074,I41575,I41261);
not I_2275 (I41606,I41541);
or I_2276 (I41623,I41606,I41312);
nor I_2277 (I41062,I41142,I41623);
nor I_2278 (I41080,I41445,I41606);
nor I_2279 (I41668,I41507,I41524);
nor I_2280 (I41685,I41411,I41668);
DFFARX1 I_2281 (I41685,I2898,I41091,I41065,);
nor I_2282 (I41716,I41668,I41227);
not I_2283 (I41071,I41716);
or I_2284 (I41077,I41668,I41261);
nor I_2285 (I41068,I41541,I41668);
not I_2286 (I41814,I2905);
nand I_2287 (I41831,I16786,I16780);
and I_2288 (I41848,I41831,I16792);
DFFARX1 I_2289 (I41848,I2898,I41814,I41874,);
not I_2290 (I41882,I41874);
nor I_2291 (I41899,I16801,I16780);
nor I_2292 (I41770,I41882,I41899);
not I_2293 (I41930,I16786);
or I_2294 (I41947,I16792,I16786);
nor I_2295 (I41964,I16783,I16792);
not I_2296 (I41981,I41964);
nor I_2297 (I41998,I16798,I16807);
nand I_2298 (I42015,I41981,I41998);
not I_2299 (I41776,I42015);
not I_2300 (I42046,I16798);
nand I_2301 (I42063,I42046,I16780);
nand I_2302 (I42080,I41930,I42063);
not I_2303 (I42097,I42080);
nor I_2304 (I42114,I42097,I41998);
nor I_2305 (I41773,I41882,I42114);
or I_2306 (I41797,I42097,I41899);
or I_2307 (I42159,I16798,I16807);
nor I_2308 (I42176,I16789,I16783);
DFFARX1 I_2309 (I42176,I2898,I41814,I42202,);
nor I_2310 (I41779,I42202,I42015);
nor I_2311 (I41806,I42202,I41899);
not I_2312 (I42238,I42202);
nor I_2313 (I42255,I16789,I16783);
nor I_2314 (I42272,I42202,I42255);
DFFARX1 I_2315 (I42272,I2898,I41814,I41791,);
nor I_2316 (I42303,I41882,I42255);
nor I_2317 (I41794,I42255,I41947);
nand I_2318 (I42334,I16789,I16804);
nor I_2319 (I42351,I42334,I16795);
nor I_2320 (I41785,I42351,I41964);
not I_2321 (I42382,I42351);
nand I_2322 (I42399,I42382,I41964);
nand I_2323 (I41803,I42382,I42080);
nor I_2324 (I41800,I42351,I42303);
not I_2325 (I42444,I42334);
nand I_2326 (I42461,I42444,I42399);
nor I_2327 (I41788,I42238,I42461);
nand I_2328 (I42492,I42334,I42159);
nand I_2329 (I42509,I42382,I42492);
nand I_2330 (I42526,I42509,I41930);
nor I_2331 (I41782,I41981,I42526);
not I_2332 (I42596,I2905);
nand I_2333 (I42613,I282660,I282690);
and I_2334 (I42630,I42613,I282675);
DFFARX1 I_2335 (I42630,I2898,I42596,I42656,);
not I_2336 (I42664,I42656);
nor I_2337 (I42681,I282666,I282690);
nor I_2338 (I42552,I42664,I42681);
not I_2339 (I42712,I282666);
or I_2340 (I42729,I282687,I282666);
nor I_2341 (I42746,I282681,I282687);
not I_2342 (I42763,I42746);
nor I_2343 (I42780,I282669,I282672);
nand I_2344 (I42797,I42763,I42780);
not I_2345 (I42558,I42797);
not I_2346 (I42828,I282669);
nand I_2347 (I42845,I42828,I282663);
nand I_2348 (I42862,I42712,I42845);
not I_2349 (I42879,I42862);
nor I_2350 (I42896,I42879,I42780);
nor I_2351 (I42555,I42664,I42896);
or I_2352 (I42579,I42879,I42681);
or I_2353 (I42941,I282669,I282672);
nor I_2354 (I42958,I282660,I282684);
DFFARX1 I_2355 (I42958,I2898,I42596,I42984,);
nor I_2356 (I42561,I42984,I42797);
nor I_2357 (I42588,I42984,I42681);
not I_2358 (I43020,I42984);
nor I_2359 (I43037,I282660,I282681);
nor I_2360 (I43054,I42984,I43037);
DFFARX1 I_2361 (I43054,I2898,I42596,I42573,);
nor I_2362 (I43085,I42664,I43037);
nor I_2363 (I42576,I43037,I42729);
nand I_2364 (I43116,I282663,I282678);
nor I_2365 (I43133,I43116,I282669);
nor I_2366 (I42567,I43133,I42746);
not I_2367 (I43164,I43133);
nand I_2368 (I43181,I43164,I42746);
nand I_2369 (I42585,I43164,I42862);
nor I_2370 (I42582,I43133,I43085);
not I_2371 (I43226,I43116);
nand I_2372 (I43243,I43226,I43181);
nor I_2373 (I42570,I43020,I43243);
nand I_2374 (I43274,I43116,I42941);
nand I_2375 (I43291,I43164,I43274);
nand I_2376 (I43308,I43291,I42712);
nor I_2377 (I42564,I42763,I43308);
not I_2378 (I43378,I2905);
nand I_2379 (I43395,I203721,I203727);
and I_2380 (I43412,I43395,I203724);
DFFARX1 I_2381 (I43412,I2898,I43378,I43438,);
not I_2382 (I43446,I43438);
nor I_2383 (I43463,I203739,I203727);
nor I_2384 (I43334,I43446,I43463);
not I_2385 (I43494,I203715);
or I_2386 (I43511,I203718,I203715);
nor I_2387 (I43528,I203712,I203718);
not I_2388 (I43545,I43528);
nor I_2389 (I43562,I203724,I203718);
nand I_2390 (I43579,I43545,I43562);
not I_2391 (I43340,I43579);
not I_2392 (I43610,I203724);
nand I_2393 (I43627,I43610,I203715);
nand I_2394 (I43644,I43494,I43627);
not I_2395 (I43661,I43644);
nor I_2396 (I43678,I43661,I43562);
nor I_2397 (I43337,I43446,I43678);
or I_2398 (I43361,I43661,I43463);
or I_2399 (I43723,I203724,I203718);
nor I_2400 (I43740,I203712,I203730);
DFFARX1 I_2401 (I43740,I2898,I43378,I43766,);
nor I_2402 (I43343,I43766,I43579);
nor I_2403 (I43370,I43766,I43463);
not I_2404 (I43802,I43766);
nor I_2405 (I43819,I203712,I203712);
nor I_2406 (I43836,I43766,I43819);
DFFARX1 I_2407 (I43836,I2898,I43378,I43355,);
nor I_2408 (I43867,I43446,I43819);
nor I_2409 (I43358,I43819,I43511);
nand I_2410 (I43898,I203733,I203736);
nor I_2411 (I43915,I43898,I203721);
nor I_2412 (I43349,I43915,I43528);
not I_2413 (I43946,I43915);
nand I_2414 (I43963,I43946,I43528);
nand I_2415 (I43367,I43946,I43644);
nor I_2416 (I43364,I43915,I43867);
not I_2417 (I44008,I43898);
nand I_2418 (I44025,I44008,I43963);
nor I_2419 (I43352,I43802,I44025);
nand I_2420 (I44056,I43898,I43723);
nand I_2421 (I44073,I43946,I44056);
nand I_2422 (I44090,I44073,I43494);
nor I_2423 (I43346,I43545,I44090);
not I_2424 (I44160,I2905);
nand I_2425 (I44177,I188342,I188339);
and I_2426 (I44194,I44177,I188336);
DFFARX1 I_2427 (I44194,I2898,I44160,I44220,);
not I_2428 (I44228,I44220);
nor I_2429 (I44245,I188333,I188339);
nor I_2430 (I44116,I44228,I44245);
not I_2431 (I44276,I188327);
or I_2432 (I44293,I188342,I188327);
nor I_2433 (I44310,I188336,I188342);
not I_2434 (I44327,I44310);
nor I_2435 (I44344,I188351,I188330);
nand I_2436 (I44361,I44327,I44344);
not I_2437 (I44122,I44361);
not I_2438 (I44392,I188351);
nand I_2439 (I44409,I44392,I188327);
nand I_2440 (I44426,I44276,I44409);
not I_2441 (I44443,I44426);
nor I_2442 (I44460,I44443,I44344);
nor I_2443 (I44119,I44228,I44460);
or I_2444 (I44143,I44443,I44245);
or I_2445 (I44505,I188351,I188330);
nor I_2446 (I44522,I188330,I188345);
DFFARX1 I_2447 (I44522,I2898,I44160,I44548,);
nor I_2448 (I44125,I44548,I44361);
nor I_2449 (I44152,I44548,I44245);
not I_2450 (I44584,I44548);
nor I_2451 (I44601,I188330,I188336);
nor I_2452 (I44618,I44548,I44601);
DFFARX1 I_2453 (I44618,I2898,I44160,I44137,);
nor I_2454 (I44649,I44228,I44601);
nor I_2455 (I44140,I44601,I44293);
nand I_2456 (I44680,I188348,I188339);
nor I_2457 (I44697,I44680,I188333);
nor I_2458 (I44131,I44697,I44310);
not I_2459 (I44728,I44697);
nand I_2460 (I44745,I44728,I44310);
nand I_2461 (I44149,I44728,I44426);
nor I_2462 (I44146,I44697,I44649);
not I_2463 (I44790,I44680);
nand I_2464 (I44807,I44790,I44745);
nor I_2465 (I44134,I44584,I44807);
nand I_2466 (I44838,I44680,I44505);
nand I_2467 (I44855,I44728,I44838);
nand I_2468 (I44872,I44855,I44276);
nor I_2469 (I44128,I44327,I44872);
not I_2470 (I44942,I2905);
nand I_2471 (I44959,I218681,I218687);
and I_2472 (I44976,I44959,I218684);
DFFARX1 I_2473 (I44976,I2898,I44942,I45002,);
not I_2474 (I45010,I45002);
nor I_2475 (I45027,I218699,I218687);
nor I_2476 (I44898,I45010,I45027);
not I_2477 (I45058,I218675);
or I_2478 (I45075,I218678,I218675);
nor I_2479 (I45092,I218672,I218678);
not I_2480 (I45109,I45092);
nor I_2481 (I45126,I218684,I218678);
nand I_2482 (I45143,I45109,I45126);
not I_2483 (I44904,I45143);
not I_2484 (I45174,I218684);
nand I_2485 (I45191,I45174,I218675);
nand I_2486 (I45208,I45058,I45191);
not I_2487 (I45225,I45208);
nor I_2488 (I45242,I45225,I45126);
nor I_2489 (I44901,I45010,I45242);
or I_2490 (I44925,I45225,I45027);
or I_2491 (I45287,I218684,I218678);
nor I_2492 (I45304,I218672,I218690);
DFFARX1 I_2493 (I45304,I2898,I44942,I45330,);
nor I_2494 (I44907,I45330,I45143);
nor I_2495 (I44934,I45330,I45027);
not I_2496 (I45366,I45330);
nor I_2497 (I45383,I218672,I218672);
nor I_2498 (I45400,I45330,I45383);
DFFARX1 I_2499 (I45400,I2898,I44942,I44919,);
nor I_2500 (I45431,I45010,I45383);
nor I_2501 (I44922,I45383,I45075);
nand I_2502 (I45462,I218693,I218696);
nor I_2503 (I45479,I45462,I218681);
nor I_2504 (I44913,I45479,I45092);
not I_2505 (I45510,I45479);
nand I_2506 (I45527,I45510,I45092);
nand I_2507 (I44931,I45510,I45208);
nor I_2508 (I44928,I45479,I45431);
not I_2509 (I45572,I45462);
nand I_2510 (I45589,I45572,I45527);
nor I_2511 (I44916,I45366,I45589);
nand I_2512 (I45620,I45462,I45287);
nand I_2513 (I45637,I45510,I45620);
nand I_2514 (I45654,I45637,I45058);
nor I_2515 (I44910,I45109,I45654);
not I_2516 (I45724,I2905);
nand I_2517 (I45741,I22498,I22492);
and I_2518 (I45758,I45741,I22504);
DFFARX1 I_2519 (I45758,I2898,I45724,I45784,);
not I_2520 (I45792,I45784);
nor I_2521 (I45809,I22513,I22492);
nor I_2522 (I45680,I45792,I45809);
not I_2523 (I45840,I22498);
or I_2524 (I45857,I22504,I22498);
nor I_2525 (I45874,I22495,I22504);
not I_2526 (I45891,I45874);
nor I_2527 (I45908,I22510,I22519);
nand I_2528 (I45925,I45891,I45908);
not I_2529 (I45686,I45925);
not I_2530 (I45956,I22510);
nand I_2531 (I45973,I45956,I22492);
nand I_2532 (I45990,I45840,I45973);
not I_2533 (I46007,I45990);
nor I_2534 (I46024,I46007,I45908);
nor I_2535 (I45683,I45792,I46024);
or I_2536 (I45707,I46007,I45809);
or I_2537 (I46069,I22510,I22519);
nor I_2538 (I46086,I22501,I22495);
DFFARX1 I_2539 (I46086,I2898,I45724,I46112,);
nor I_2540 (I45689,I46112,I45925);
nor I_2541 (I45716,I46112,I45809);
not I_2542 (I46148,I46112);
nor I_2543 (I46165,I22501,I22495);
nor I_2544 (I46182,I46112,I46165);
DFFARX1 I_2545 (I46182,I2898,I45724,I45701,);
nor I_2546 (I46213,I45792,I46165);
nor I_2547 (I45704,I46165,I45857);
nand I_2548 (I46244,I22501,I22516);
nor I_2549 (I46261,I46244,I22507);
nor I_2550 (I45695,I46261,I45874);
not I_2551 (I46292,I46261);
nand I_2552 (I46309,I46292,I45874);
nand I_2553 (I45713,I46292,I45990);
nor I_2554 (I45710,I46261,I46213);
not I_2555 (I46354,I46244);
nand I_2556 (I46371,I46354,I46309);
nor I_2557 (I45698,I46148,I46371);
nand I_2558 (I46402,I46244,I46069);
nand I_2559 (I46419,I46292,I46402);
nand I_2560 (I46436,I46419,I45840);
nor I_2561 (I45692,I45891,I46436);
not I_2562 (I46506,I2905);
nand I_2563 (I46523,I91544,I91535);
and I_2564 (I46540,I46523,I91529);
DFFARX1 I_2565 (I46540,I2898,I46506,I46566,);
not I_2566 (I46574,I46566);
nor I_2567 (I46591,I91553,I91535);
nor I_2568 (I46462,I46574,I46591);
not I_2569 (I46622,I91547);
or I_2570 (I46639,I91538,I91547);
nor I_2571 (I46656,I91535,I91538);
not I_2572 (I46673,I46656);
nor I_2573 (I46690,I91538,I91532);
nand I_2574 (I46707,I46673,I46690);
not I_2575 (I46468,I46707);
not I_2576 (I46738,I91538);
nand I_2577 (I46755,I46738,I91550);
nand I_2578 (I46772,I46622,I46755);
not I_2579 (I46789,I46772);
nor I_2580 (I46806,I46789,I46690);
nor I_2581 (I46465,I46574,I46806);
or I_2582 (I46489,I46789,I46591);
or I_2583 (I46851,I91538,I91532);
nor I_2584 (I46868,I91541,I91529);
DFFARX1 I_2585 (I46868,I2898,I46506,I46894,);
nor I_2586 (I46471,I46894,I46707);
nor I_2587 (I46498,I46894,I46591);
not I_2588 (I46930,I46894);
nor I_2589 (I46947,I91541,I91535);
nor I_2590 (I46964,I46894,I46947);
DFFARX1 I_2591 (I46964,I2898,I46506,I46483,);
nor I_2592 (I46995,I46574,I46947);
nor I_2593 (I46486,I46947,I46639);
nand I_2594 (I47026,I91541,I91556);
nor I_2595 (I47043,I47026,I91532);
nor I_2596 (I46477,I47043,I46656);
not I_2597 (I47074,I47043);
nand I_2598 (I47091,I47074,I46656);
nand I_2599 (I46495,I47074,I46772);
nor I_2600 (I46492,I47043,I46995);
not I_2601 (I47136,I47026);
nand I_2602 (I47153,I47136,I47091);
nor I_2603 (I46480,I46930,I47153);
nand I_2604 (I47184,I47026,I46851);
nand I_2605 (I47201,I47074,I47184);
nand I_2606 (I47218,I47201,I46622);
nor I_2607 (I46474,I46673,I47218);
not I_2608 (I47288,I2905);
nand I_2609 (I47305,I20356,I20350);
and I_2610 (I47322,I47305,I20362);
DFFARX1 I_2611 (I47322,I2898,I47288,I47348,);
not I_2612 (I47356,I47348);
nor I_2613 (I47373,I20371,I20350);
nor I_2614 (I47244,I47356,I47373);
not I_2615 (I47404,I20356);
or I_2616 (I47421,I20362,I20356);
nor I_2617 (I47438,I20353,I20362);
not I_2618 (I47455,I47438);
nor I_2619 (I47472,I20368,I20377);
nand I_2620 (I47489,I47455,I47472);
not I_2621 (I47250,I47489);
not I_2622 (I47520,I20368);
nand I_2623 (I47537,I47520,I20350);
nand I_2624 (I47554,I47404,I47537);
not I_2625 (I47571,I47554);
nor I_2626 (I47588,I47571,I47472);
nor I_2627 (I47247,I47356,I47588);
or I_2628 (I47271,I47571,I47373);
or I_2629 (I47633,I20368,I20377);
nor I_2630 (I47650,I20359,I20353);
DFFARX1 I_2631 (I47650,I2898,I47288,I47676,);
nor I_2632 (I47253,I47676,I47489);
nor I_2633 (I47280,I47676,I47373);
not I_2634 (I47712,I47676);
nor I_2635 (I47729,I20359,I20353);
nor I_2636 (I47746,I47676,I47729);
DFFARX1 I_2637 (I47746,I2898,I47288,I47265,);
nor I_2638 (I47777,I47356,I47729);
nor I_2639 (I47268,I47729,I47421);
nand I_2640 (I47808,I20359,I20374);
nor I_2641 (I47825,I47808,I20365);
nor I_2642 (I47259,I47825,I47438);
not I_2643 (I47856,I47825);
nand I_2644 (I47873,I47856,I47438);
nand I_2645 (I47277,I47856,I47554);
nor I_2646 (I47274,I47825,I47777);
not I_2647 (I47918,I47808);
nand I_2648 (I47935,I47918,I47873);
nor I_2649 (I47262,I47712,I47935);
nand I_2650 (I47966,I47808,I47633);
nand I_2651 (I47983,I47856,I47966);
nand I_2652 (I48000,I47983,I47404);
nor I_2653 (I47256,I47455,I48000);
not I_2654 (I48070,I2905);
nand I_2655 (I48087,I306894,I306912);
and I_2656 (I48104,I48087,I306900);
DFFARX1 I_2657 (I48104,I2898,I48070,I48130,);
not I_2658 (I48138,I48130);
nor I_2659 (I48155,I306885,I306912);
nor I_2660 (I48026,I48138,I48155);
not I_2661 (I48186,I306915);
or I_2662 (I48203,I306909,I306915);
nor I_2663 (I48220,I306891,I306909);
not I_2664 (I48237,I48220);
nor I_2665 (I48254,I306894,I306888);
nand I_2666 (I48271,I48237,I48254);
not I_2667 (I48032,I48271);
not I_2668 (I48302,I306894);
nand I_2669 (I48319,I48302,I306888);
nand I_2670 (I48336,I48186,I48319);
not I_2671 (I48353,I48336);
nor I_2672 (I48370,I48353,I48254);
nor I_2673 (I48029,I48138,I48370);
or I_2674 (I48053,I48353,I48155);
or I_2675 (I48415,I306894,I306888);
nor I_2676 (I48432,I306903,I306891);
DFFARX1 I_2677 (I48432,I2898,I48070,I48458,);
nor I_2678 (I48035,I48458,I48271);
nor I_2679 (I48062,I48458,I48155);
not I_2680 (I48494,I48458);
nor I_2681 (I48511,I306903,I306891);
nor I_2682 (I48528,I48458,I48511);
DFFARX1 I_2683 (I48528,I2898,I48070,I48047,);
nor I_2684 (I48559,I48138,I48511);
nor I_2685 (I48050,I48511,I48203);
nand I_2686 (I48590,I306897,I306906);
nor I_2687 (I48607,I48590,I306885);
nor I_2688 (I48041,I48607,I48220);
not I_2689 (I48638,I48607);
nand I_2690 (I48655,I48638,I48220);
nand I_2691 (I48059,I48638,I48336);
nor I_2692 (I48056,I48607,I48559);
not I_2693 (I48700,I48590);
nand I_2694 (I48717,I48700,I48655);
nor I_2695 (I48044,I48494,I48717);
nand I_2696 (I48748,I48590,I48415);
nand I_2697 (I48765,I48638,I48748);
nand I_2698 (I48782,I48765,I48186);
nor I_2699 (I48038,I48237,I48782);
not I_2700 (I48852,I2905);
nand I_2701 (I48869,I356154,I356157);
and I_2702 (I48886,I48869,I356166);
DFFARX1 I_2703 (I48886,I2898,I48852,I48912,);
not I_2704 (I48920,I48912);
nor I_2705 (I48937,I356160,I356157);
nor I_2706 (I48808,I48920,I48937);
not I_2707 (I48968,I356151);
or I_2708 (I48985,I356157,I356151);
nor I_2709 (I49002,I356166,I356157);
not I_2710 (I49019,I49002);
nor I_2711 (I49036,I356160,I356175);
nand I_2712 (I49053,I49019,I49036);
not I_2713 (I48814,I49053);
not I_2714 (I49084,I356160);
nand I_2715 (I49101,I49084,I356163);
nand I_2716 (I49118,I48968,I49101);
not I_2717 (I49135,I49118);
nor I_2718 (I49152,I49135,I49036);
nor I_2719 (I48811,I48920,I49152);
or I_2720 (I48835,I49135,I48937);
or I_2721 (I49197,I356160,I356175);
nor I_2722 (I49214,I356169,I356163);
DFFARX1 I_2723 (I49214,I2898,I48852,I49240,);
nor I_2724 (I48817,I49240,I49053);
nor I_2725 (I48844,I49240,I48937);
not I_2726 (I49276,I49240);
nor I_2727 (I49293,I356169,I356166);
nor I_2728 (I49310,I49240,I49293);
DFFARX1 I_2729 (I49310,I2898,I48852,I48829,);
nor I_2730 (I49341,I48920,I49293);
nor I_2731 (I48832,I49293,I48985);
nand I_2732 (I49372,I356154,I356172);
nor I_2733 (I49389,I49372,I356151);
nor I_2734 (I48823,I49389,I49002);
not I_2735 (I49420,I49389);
nand I_2736 (I49437,I49420,I49002);
nand I_2737 (I48841,I49420,I49118);
nor I_2738 (I48838,I49389,I49341);
not I_2739 (I49482,I49372);
nand I_2740 (I49499,I49482,I49437);
nor I_2741 (I48826,I49276,I49499);
nand I_2742 (I49530,I49372,I49197);
nand I_2743 (I49547,I49420,I49530);
nand I_2744 (I49564,I49547,I48968);
nor I_2745 (I48820,I49019,I49564);
not I_2746 (I49634,I2905);
nand I_2747 (I49651,I277305,I277335);
and I_2748 (I49668,I49651,I277320);
DFFARX1 I_2749 (I49668,I2898,I49634,I49694,);
not I_2750 (I49702,I49694);
nor I_2751 (I49719,I277311,I277335);
nor I_2752 (I49590,I49702,I49719);
not I_2753 (I49750,I277311);
or I_2754 (I49767,I277332,I277311);
nor I_2755 (I49784,I277326,I277332);
not I_2756 (I49801,I49784);
nor I_2757 (I49818,I277314,I277317);
nand I_2758 (I49835,I49801,I49818);
not I_2759 (I49596,I49835);
not I_2760 (I49866,I277314);
nand I_2761 (I49883,I49866,I277308);
nand I_2762 (I49900,I49750,I49883);
not I_2763 (I49917,I49900);
nor I_2764 (I49934,I49917,I49818);
nor I_2765 (I49593,I49702,I49934);
or I_2766 (I49617,I49917,I49719);
or I_2767 (I49979,I277314,I277317);
nor I_2768 (I49996,I277305,I277329);
DFFARX1 I_2769 (I49996,I2898,I49634,I50022,);
nor I_2770 (I49599,I50022,I49835);
nor I_2771 (I49626,I50022,I49719);
not I_2772 (I50058,I50022);
nor I_2773 (I50075,I277305,I277326);
nor I_2774 (I50092,I50022,I50075);
DFFARX1 I_2775 (I50092,I2898,I49634,I49611,);
nor I_2776 (I50123,I49702,I50075);
nor I_2777 (I49614,I50075,I49767);
nand I_2778 (I50154,I277308,I277323);
nor I_2779 (I50171,I50154,I277314);
nor I_2780 (I49605,I50171,I49784);
not I_2781 (I50202,I50171);
nand I_2782 (I50219,I50202,I49784);
nand I_2783 (I49623,I50202,I49900);
nor I_2784 (I49620,I50171,I50123);
not I_2785 (I50264,I50154);
nand I_2786 (I50281,I50264,I50219);
nor I_2787 (I49608,I50058,I50281);
nand I_2788 (I50312,I50154,I49979);
nand I_2789 (I50329,I50202,I50312);
nand I_2790 (I50346,I50329,I49750);
nor I_2791 (I49602,I49801,I50346);
not I_2792 (I50416,I2905);
nand I_2793 (I50433,I368899,I368890);
and I_2794 (I50450,I50433,I368902);
DFFARX1 I_2795 (I50450,I2898,I50416,I50476,);
not I_2796 (I50484,I50476);
nor I_2797 (I50501,I368914,I368890);
nor I_2798 (I50372,I50484,I50501);
not I_2799 (I50532,I368908);
or I_2800 (I50549,I368893,I368908);
nor I_2801 (I50566,I368911,I368893);
not I_2802 (I50583,I50566);
nor I_2803 (I50600,I368917,I368887);
nand I_2804 (I50617,I50583,I50600);
not I_2805 (I50378,I50617);
not I_2806 (I50648,I368917);
nand I_2807 (I50665,I50648,I368884);
nand I_2808 (I50682,I50532,I50665);
not I_2809 (I50699,I50682);
nor I_2810 (I50716,I50699,I50600);
nor I_2811 (I50375,I50484,I50716);
or I_2812 (I50399,I50699,I50501);
or I_2813 (I50761,I368917,I368887);
nor I_2814 (I50778,I368887,I368884);
DFFARX1 I_2815 (I50778,I2898,I50416,I50804,);
nor I_2816 (I50381,I50804,I50617);
nor I_2817 (I50408,I50804,I50501);
not I_2818 (I50840,I50804);
nor I_2819 (I50857,I368887,I368911);
nor I_2820 (I50874,I50804,I50857);
DFFARX1 I_2821 (I50874,I2898,I50416,I50393,);
nor I_2822 (I50905,I50484,I50857);
nor I_2823 (I50396,I50857,I50549);
nand I_2824 (I50936,I368905,I368896);
nor I_2825 (I50953,I50936,I368890);
nor I_2826 (I50387,I50953,I50566);
not I_2827 (I50984,I50953);
nand I_2828 (I51001,I50984,I50566);
nand I_2829 (I50405,I50984,I50682);
nor I_2830 (I50402,I50953,I50905);
not I_2831 (I51046,I50936);
nand I_2832 (I51063,I51046,I51001);
nor I_2833 (I50390,I50840,I51063);
nand I_2834 (I51094,I50936,I50761);
nand I_2835 (I51111,I50984,I51094);
nand I_2836 (I51128,I51111,I50532);
nor I_2837 (I50384,I50583,I51128);
not I_2838 (I51198,I2905);
nand I_2839 (I51215,I347229,I347232);
and I_2840 (I51232,I51215,I347241);
DFFARX1 I_2841 (I51232,I2898,I51198,I51258,);
not I_2842 (I51266,I51258);
nor I_2843 (I51283,I347235,I347232);
nor I_2844 (I51154,I51266,I51283);
not I_2845 (I51314,I347226);
or I_2846 (I51331,I347232,I347226);
nor I_2847 (I51348,I347241,I347232);
not I_2848 (I51365,I51348);
nor I_2849 (I51382,I347235,I347250);
nand I_2850 (I51399,I51365,I51382);
not I_2851 (I51160,I51399);
not I_2852 (I51430,I347235);
nand I_2853 (I51447,I51430,I347238);
nand I_2854 (I51464,I51314,I51447);
not I_2855 (I51481,I51464);
nor I_2856 (I51498,I51481,I51382);
nor I_2857 (I51157,I51266,I51498);
or I_2858 (I51181,I51481,I51283);
or I_2859 (I51543,I347235,I347250);
nor I_2860 (I51560,I347244,I347238);
DFFARX1 I_2861 (I51560,I2898,I51198,I51586,);
nor I_2862 (I51163,I51586,I51399);
nor I_2863 (I51190,I51586,I51283);
not I_2864 (I51622,I51586);
nor I_2865 (I51639,I347244,I347241);
nor I_2866 (I51656,I51586,I51639);
DFFARX1 I_2867 (I51656,I2898,I51198,I51175,);
nor I_2868 (I51687,I51266,I51639);
nor I_2869 (I51178,I51639,I51331);
nand I_2870 (I51718,I347229,I347247);
nor I_2871 (I51735,I51718,I347226);
nor I_2872 (I51169,I51735,I51348);
not I_2873 (I51766,I51735);
nand I_2874 (I51783,I51766,I51348);
nand I_2875 (I51187,I51766,I51464);
nor I_2876 (I51184,I51735,I51687);
not I_2877 (I51828,I51718);
nand I_2878 (I51845,I51828,I51783);
nor I_2879 (I51172,I51622,I51845);
nand I_2880 (I51876,I51718,I51543);
nand I_2881 (I51893,I51766,I51876);
nand I_2882 (I51910,I51893,I51314);
nor I_2883 (I51166,I51365,I51910);
not I_2884 (I51980,I2905);
nand I_2885 (I51997,I177649,I177634);
and I_2886 (I52014,I51997,I177634);
DFFARX1 I_2887 (I52014,I2898,I51980,I52040,);
not I_2888 (I52048,I52040);
nor I_2889 (I52065,I177640,I177634);
nor I_2890 (I51936,I52048,I52065);
not I_2891 (I52096,I177658);
or I_2892 (I52113,I177661,I177658);
nor I_2893 (I52130,I177646,I177661);
not I_2894 (I52147,I52130);
nor I_2895 (I52164,I177640,I177664);
nand I_2896 (I52181,I52147,I52164);
not I_2897 (I51942,I52181);
not I_2898 (I52212,I177640);
nand I_2899 (I52229,I52212,I177643);
nand I_2900 (I52246,I52096,I52229);
not I_2901 (I52263,I52246);
nor I_2902 (I52280,I52263,I52164);
nor I_2903 (I51939,I52048,I52280);
or I_2904 (I51963,I52263,I52065);
or I_2905 (I52325,I177640,I177664);
nor I_2906 (I52342,I177637,I177637);
DFFARX1 I_2907 (I52342,I2898,I51980,I52368,);
nor I_2908 (I51945,I52368,I52181);
nor I_2909 (I51972,I52368,I52065);
not I_2910 (I52404,I52368);
nor I_2911 (I52421,I177637,I177646);
nor I_2912 (I52438,I52368,I52421);
DFFARX1 I_2913 (I52438,I2898,I51980,I51957,);
nor I_2914 (I52469,I52048,I52421);
nor I_2915 (I51960,I52421,I52113);
nand I_2916 (I52500,I177652,I177655);
nor I_2917 (I52517,I52500,I177643);
nor I_2918 (I51951,I52517,I52130);
not I_2919 (I52548,I52517);
nand I_2920 (I52565,I52548,I52130);
nand I_2921 (I51969,I52548,I52246);
nor I_2922 (I51966,I52517,I52469);
not I_2923 (I52610,I52500);
nand I_2924 (I52627,I52610,I52565);
nor I_2925 (I51954,I52404,I52627);
nand I_2926 (I52658,I52500,I52325);
nand I_2927 (I52675,I52548,I52658);
nand I_2928 (I52692,I52675,I52096);
nor I_2929 (I51948,I52147,I52692);
not I_2930 (I52762,I2905);
nand I_2931 (I52779,I101545,I101566);
and I_2932 (I52796,I52779,I101575);
DFFARX1 I_2933 (I52796,I2898,I52762,I52822,);
not I_2934 (I52830,I52822);
nor I_2935 (I52847,I101569,I101566);
nor I_2936 (I52718,I52830,I52847);
not I_2937 (I52878,I101560);
or I_2938 (I52895,I101563,I101560);
nor I_2939 (I52912,I101551,I101563);
not I_2940 (I52929,I52912);
nor I_2941 (I52946,I101548,I101545);
nand I_2942 (I52963,I52929,I52946);
not I_2943 (I52724,I52963);
not I_2944 (I52994,I101548);
nand I_2945 (I53011,I52994,I101542);
nand I_2946 (I53028,I52878,I53011);
not I_2947 (I53045,I53028);
nor I_2948 (I53062,I53045,I52946);
nor I_2949 (I52721,I52830,I53062);
or I_2950 (I52745,I53045,I52847);
or I_2951 (I53107,I101548,I101545);
nor I_2952 (I53124,I101557,I101554);
DFFARX1 I_2953 (I53124,I2898,I52762,I53150,);
nor I_2954 (I52727,I53150,I52963);
nor I_2955 (I52754,I53150,I52847);
not I_2956 (I53186,I53150);
nor I_2957 (I53203,I101557,I101551);
nor I_2958 (I53220,I53150,I53203);
DFFARX1 I_2959 (I53220,I2898,I52762,I52739,);
nor I_2960 (I53251,I52830,I53203);
nor I_2961 (I52742,I53203,I52895);
nand I_2962 (I53282,I101572,I101542);
nor I_2963 (I53299,I53282,I101548);
nor I_2964 (I52733,I53299,I52912);
not I_2965 (I53330,I53299);
nand I_2966 (I53347,I53330,I52912);
nand I_2967 (I52751,I53330,I53028);
nor I_2968 (I52748,I53299,I53251);
not I_2969 (I53392,I53282);
nand I_2970 (I53409,I53392,I53347);
nor I_2971 (I52736,I53186,I53409);
nand I_2972 (I53440,I53282,I53107);
nand I_2973 (I53457,I53330,I53440);
nand I_2974 (I53474,I53457,I52878);
nor I_2975 (I52730,I52929,I53474);
not I_2976 (I53544,I2905);
nand I_2977 (I53561,I108464,I108485);
and I_2978 (I53578,I53561,I108494);
DFFARX1 I_2979 (I53578,I2898,I53544,I53604,);
not I_2980 (I53612,I53604);
nor I_2981 (I53629,I108488,I108485);
nor I_2982 (I53500,I53612,I53629);
not I_2983 (I53660,I108479);
or I_2984 (I53677,I108482,I108479);
nor I_2985 (I53694,I108470,I108482);
not I_2986 (I53711,I53694);
nor I_2987 (I53728,I108467,I108464);
nand I_2988 (I53745,I53711,I53728);
not I_2989 (I53506,I53745);
not I_2990 (I53776,I108467);
nand I_2991 (I53793,I53776,I108461);
nand I_2992 (I53810,I53660,I53793);
not I_2993 (I53827,I53810);
nor I_2994 (I53844,I53827,I53728);
nor I_2995 (I53503,I53612,I53844);
or I_2996 (I53527,I53827,I53629);
or I_2997 (I53889,I108467,I108464);
nor I_2998 (I53906,I108476,I108473);
DFFARX1 I_2999 (I53906,I2898,I53544,I53932,);
nor I_3000 (I53509,I53932,I53745);
nor I_3001 (I53536,I53932,I53629);
not I_3002 (I53968,I53932);
nor I_3003 (I53985,I108476,I108470);
nor I_3004 (I54002,I53932,I53985);
DFFARX1 I_3005 (I54002,I2898,I53544,I53521,);
nor I_3006 (I54033,I53612,I53985);
nor I_3007 (I53524,I53985,I53677);
nand I_3008 (I54064,I108491,I108461);
nor I_3009 (I54081,I54064,I108467);
nor I_3010 (I53515,I54081,I53694);
not I_3011 (I54112,I54081);
nand I_3012 (I54129,I54112,I53694);
nand I_3013 (I53533,I54112,I53810);
nor I_3014 (I53530,I54081,I54033);
not I_3015 (I54174,I54064);
nand I_3016 (I54191,I54174,I54129);
nor I_3017 (I53518,I53968,I54191);
nand I_3018 (I54222,I54064,I53889);
nand I_3019 (I54239,I54112,I54222);
nand I_3020 (I54256,I54239,I53660);
nor I_3021 (I53512,I53711,I54256);
not I_3022 (I54326,I2905);
nand I_3023 (I54343,I70158,I70149);
and I_3024 (I54360,I54343,I70143);
DFFARX1 I_3025 (I54360,I2898,I54326,I54386,);
not I_3026 (I54394,I54386);
nor I_3027 (I54411,I70167,I70149);
nor I_3028 (I54282,I54394,I54411);
not I_3029 (I54442,I70161);
or I_3030 (I54459,I70152,I70161);
nor I_3031 (I54476,I70149,I70152);
not I_3032 (I54493,I54476);
nor I_3033 (I54510,I70152,I70146);
nand I_3034 (I54527,I54493,I54510);
not I_3035 (I54288,I54527);
not I_3036 (I54558,I70152);
nand I_3037 (I54575,I54558,I70164);
nand I_3038 (I54592,I54442,I54575);
not I_3039 (I54609,I54592);
nor I_3040 (I54626,I54609,I54510);
nor I_3041 (I54285,I54394,I54626);
or I_3042 (I54309,I54609,I54411);
or I_3043 (I54671,I70152,I70146);
nor I_3044 (I54688,I70155,I70143);
DFFARX1 I_3045 (I54688,I2898,I54326,I54714,);
nor I_3046 (I54291,I54714,I54527);
nor I_3047 (I54318,I54714,I54411);
not I_3048 (I54750,I54714);
nor I_3049 (I54767,I70155,I70149);
nor I_3050 (I54784,I54714,I54767);
DFFARX1 I_3051 (I54784,I2898,I54326,I54303,);
nor I_3052 (I54815,I54394,I54767);
nor I_3053 (I54306,I54767,I54459);
nand I_3054 (I54846,I70155,I70170);
nor I_3055 (I54863,I54846,I70146);
nor I_3056 (I54297,I54863,I54476);
not I_3057 (I54894,I54863);
nand I_3058 (I54911,I54894,I54476);
nand I_3059 (I54315,I54894,I54592);
nor I_3060 (I54312,I54863,I54815);
not I_3061 (I54956,I54846);
nand I_3062 (I54973,I54956,I54911);
nor I_3063 (I54300,I54750,I54973);
nand I_3064 (I55004,I54846,I54671);
nand I_3065 (I55021,I54894,I55004);
nand I_3066 (I55038,I55021,I54442);
nor I_3067 (I54294,I54493,I55038);
not I_3068 (I55108,I2905);
nand I_3069 (I55125,I105319,I105340);
and I_3070 (I55142,I55125,I105349);
DFFARX1 I_3071 (I55142,I2898,I55108,I55168,);
not I_3072 (I55176,I55168);
nor I_3073 (I55193,I105343,I105340);
nor I_3074 (I55064,I55176,I55193);
not I_3075 (I55224,I105334);
or I_3076 (I55241,I105337,I105334);
nor I_3077 (I55258,I105325,I105337);
not I_3078 (I55275,I55258);
nor I_3079 (I55292,I105322,I105319);
nand I_3080 (I55309,I55275,I55292);
not I_3081 (I55070,I55309);
not I_3082 (I55340,I105322);
nand I_3083 (I55357,I55340,I105316);
nand I_3084 (I55374,I55224,I55357);
not I_3085 (I55391,I55374);
nor I_3086 (I55408,I55391,I55292);
nor I_3087 (I55067,I55176,I55408);
or I_3088 (I55091,I55391,I55193);
or I_3089 (I55453,I105322,I105319);
nor I_3090 (I55470,I105331,I105328);
DFFARX1 I_3091 (I55470,I2898,I55108,I55496,);
nor I_3092 (I55073,I55496,I55309);
nor I_3093 (I55100,I55496,I55193);
not I_3094 (I55532,I55496);
nor I_3095 (I55549,I105331,I105325);
nor I_3096 (I55566,I55496,I55549);
DFFARX1 I_3097 (I55566,I2898,I55108,I55085,);
nor I_3098 (I55597,I55176,I55549);
nor I_3099 (I55088,I55549,I55241);
nand I_3100 (I55628,I105346,I105316);
nor I_3101 (I55645,I55628,I105322);
nor I_3102 (I55079,I55645,I55258);
not I_3103 (I55676,I55645);
nand I_3104 (I55693,I55676,I55258);
nand I_3105 (I55097,I55676,I55374);
nor I_3106 (I55094,I55645,I55597);
not I_3107 (I55738,I55628);
nand I_3108 (I55755,I55738,I55693);
nor I_3109 (I55082,I55532,I55755);
nand I_3110 (I55786,I55628,I55453);
nand I_3111 (I55803,I55676,I55786);
nand I_3112 (I55820,I55803,I55224);
nor I_3113 (I55076,I55275,I55820);
not I_3114 (I55890,I2905);
nand I_3115 (I55907,I314204,I314222);
and I_3116 (I55924,I55907,I314210);
DFFARX1 I_3117 (I55924,I2898,I55890,I55950,);
not I_3118 (I55958,I55950);
nor I_3119 (I55975,I314195,I314222);
nor I_3120 (I55846,I55958,I55975);
not I_3121 (I56006,I314225);
or I_3122 (I56023,I314219,I314225);
nor I_3123 (I56040,I314201,I314219);
not I_3124 (I56057,I56040);
nor I_3125 (I56074,I314204,I314198);
nand I_3126 (I56091,I56057,I56074);
not I_3127 (I55852,I56091);
not I_3128 (I56122,I314204);
nand I_3129 (I56139,I56122,I314198);
nand I_3130 (I56156,I56006,I56139);
not I_3131 (I56173,I56156);
nor I_3132 (I56190,I56173,I56074);
nor I_3133 (I55849,I55958,I56190);
or I_3134 (I55873,I56173,I55975);
or I_3135 (I56235,I314204,I314198);
nor I_3136 (I56252,I314213,I314201);
DFFARX1 I_3137 (I56252,I2898,I55890,I56278,);
nor I_3138 (I55855,I56278,I56091);
nor I_3139 (I55882,I56278,I55975);
not I_3140 (I56314,I56278);
nor I_3141 (I56331,I314213,I314201);
nor I_3142 (I56348,I56278,I56331);
DFFARX1 I_3143 (I56348,I2898,I55890,I55867,);
nor I_3144 (I56379,I55958,I56331);
nor I_3145 (I55870,I56331,I56023);
nand I_3146 (I56410,I314207,I314216);
nor I_3147 (I56427,I56410,I314195);
nor I_3148 (I55861,I56427,I56040);
not I_3149 (I56458,I56427);
nand I_3150 (I56475,I56458,I56040);
nand I_3151 (I55879,I56458,I56156);
nor I_3152 (I55876,I56427,I56379);
not I_3153 (I56520,I56410);
nand I_3154 (I56537,I56520,I56475);
nor I_3155 (I55864,I56314,I56537);
nand I_3156 (I56568,I56410,I56235);
nand I_3157 (I56585,I56458,I56568);
nand I_3158 (I56602,I56585,I56006);
nor I_3159 (I55858,I56057,I56602);
not I_3160 (I56672,I2905);
nand I_3161 (I56689,I68900,I68891);
and I_3162 (I56706,I56689,I68885);
DFFARX1 I_3163 (I56706,I2898,I56672,I56732,);
not I_3164 (I56740,I56732);
nor I_3165 (I56757,I68909,I68891);
nor I_3166 (I56628,I56740,I56757);
not I_3167 (I56788,I68903);
or I_3168 (I56805,I68894,I68903);
nor I_3169 (I56822,I68891,I68894);
not I_3170 (I56839,I56822);
nor I_3171 (I56856,I68894,I68888);
nand I_3172 (I56873,I56839,I56856);
not I_3173 (I56634,I56873);
not I_3174 (I56904,I68894);
nand I_3175 (I56921,I56904,I68906);
nand I_3176 (I56938,I56788,I56921);
not I_3177 (I56955,I56938);
nor I_3178 (I56972,I56955,I56856);
nor I_3179 (I56631,I56740,I56972);
or I_3180 (I56655,I56955,I56757);
or I_3181 (I57017,I68894,I68888);
nor I_3182 (I57034,I68897,I68885);
DFFARX1 I_3183 (I57034,I2898,I56672,I57060,);
nor I_3184 (I56637,I57060,I56873);
nor I_3185 (I56664,I57060,I56757);
not I_3186 (I57096,I57060);
nor I_3187 (I57113,I68897,I68891);
nor I_3188 (I57130,I57060,I57113);
DFFARX1 I_3189 (I57130,I2898,I56672,I56649,);
nor I_3190 (I57161,I56740,I57113);
nor I_3191 (I56652,I57113,I56805);
nand I_3192 (I57192,I68897,I68912);
nor I_3193 (I57209,I57192,I68888);
nor I_3194 (I56643,I57209,I56822);
not I_3195 (I57240,I57209);
nand I_3196 (I57257,I57240,I56822);
nand I_3197 (I56661,I57240,I56938);
nor I_3198 (I56658,I57209,I57161);
not I_3199 (I57302,I57192);
nand I_3200 (I57319,I57302,I57257);
nor I_3201 (I56646,I57096,I57319);
nand I_3202 (I57350,I57192,I57017);
nand I_3203 (I57367,I57240,I57350);
nand I_3204 (I57384,I57367,I56788);
nor I_3205 (I56640,I56839,I57384);
not I_3206 (I57454,I2905);
nand I_3207 (I57471,I179842,I179827);
and I_3208 (I57488,I57471,I179827);
DFFARX1 I_3209 (I57488,I2898,I57454,I57514,);
not I_3210 (I57522,I57514);
nor I_3211 (I57539,I179833,I179827);
nor I_3212 (I57410,I57522,I57539);
not I_3213 (I57570,I179851);
or I_3214 (I57587,I179854,I179851);
nor I_3215 (I57604,I179839,I179854);
not I_3216 (I57621,I57604);
nor I_3217 (I57638,I179833,I179857);
nand I_3218 (I57655,I57621,I57638);
not I_3219 (I57416,I57655);
not I_3220 (I57686,I179833);
nand I_3221 (I57703,I57686,I179836);
nand I_3222 (I57720,I57570,I57703);
not I_3223 (I57737,I57720);
nor I_3224 (I57754,I57737,I57638);
nor I_3225 (I57413,I57522,I57754);
or I_3226 (I57437,I57737,I57539);
or I_3227 (I57799,I179833,I179857);
nor I_3228 (I57816,I179830,I179830);
DFFARX1 I_3229 (I57816,I2898,I57454,I57842,);
nor I_3230 (I57419,I57842,I57655);
nor I_3231 (I57446,I57842,I57539);
not I_3232 (I57878,I57842);
nor I_3233 (I57895,I179830,I179839);
nor I_3234 (I57912,I57842,I57895);
DFFARX1 I_3235 (I57912,I2898,I57454,I57431,);
nor I_3236 (I57943,I57522,I57895);
nor I_3237 (I57434,I57895,I57587);
nand I_3238 (I57974,I179845,I179848);
nor I_3239 (I57991,I57974,I179836);
nor I_3240 (I57425,I57991,I57604);
not I_3241 (I58022,I57991);
nand I_3242 (I58039,I58022,I57604);
nand I_3243 (I57443,I58022,I57720);
nor I_3244 (I57440,I57991,I57943);
not I_3245 (I58084,I57974);
nand I_3246 (I58101,I58084,I58039);
nor I_3247 (I57428,I57878,I58101);
nand I_3248 (I58132,I57974,I57799);
nand I_3249 (I58149,I58022,I58132);
nand I_3250 (I58166,I58149,I57570);
nor I_3251 (I57422,I57621,I58166);
not I_3252 (I58227,I2905);
nor I_3253 (I58244,I202270,I202270);
nor I_3254 (I58261,I58244,I202288);
not I_3255 (I58278,I58261);
not I_3256 (I58295,I202285);
nor I_3257 (I58312,I58295,I58244);
not I_3258 (I58329,I58312);
nand I_3259 (I58207,I58278,I58329);
nand I_3260 (I58360,I58261,I202291);
not I_3261 (I58192,I58360);
nor I_3262 (I58216,I58312,I202291);
not I_3263 (I58405,I202279);
nand I_3264 (I58422,I202267,I202279);
nand I_3265 (I58439,I58422,I58405);
nand I_3266 (I58456,I58422,I202279);
not I_3267 (I58473,I58456);
nor I_3268 (I58195,I58473,I58360);
nor I_3269 (I58504,I58473,I202291);
nand I_3270 (I58213,I58278,I58456);
and I_3271 (I58535,I58439,I202273);
nand I_3272 (I58552,I58535,I202276);
not I_3273 (I58569,I58552);
nor I_3274 (I58219,I58569,I58504);
nor I_3275 (I58600,I202267,I202273);
or I_3276 (I58617,I58600,I202276);
nor I_3277 (I58634,I202282,I202282);
nand I_3278 (I58651,I58634,I58617);
not I_3279 (I58668,I58651);
nor I_3280 (I58685,I58668,I58312);
or I_3281 (I58702,I58685,I58552);
nor I_3282 (I58201,I58278,I58702);
nor I_3283 (I58733,I58668,I202291);
DFFARX1 I_3284 (I58733,I2898,I58227,I58204,);
nor I_3285 (I58764,I58668,I58552);
nor I_3286 (I58210,I58473,I58764);
nor I_3287 (I58795,I58552,I58651);
nor I_3288 (I58198,I58329,I58795);
not I_3289 (I58856,I2905);
nor I_3290 (I58873,I396549,I396558);
nor I_3291 (I58890,I58873,I396552);
not I_3292 (I58907,I58890);
not I_3293 (I58924,I396543);
nor I_3294 (I58941,I58924,I58873);
not I_3295 (I58958,I58941);
nand I_3296 (I58836,I58907,I58958);
nand I_3297 (I58989,I58890,I396549);
not I_3298 (I58821,I58989);
nor I_3299 (I58845,I58941,I396549);
not I_3300 (I59034,I396558);
nand I_3301 (I59051,I396543,I396546);
nand I_3302 (I59068,I59051,I59034);
nand I_3303 (I59085,I59051,I396558);
not I_3304 (I59102,I59085);
nor I_3305 (I58824,I59102,I58989);
nor I_3306 (I59133,I59102,I396549);
nand I_3307 (I58842,I58907,I59085);
and I_3308 (I59164,I59068,I396552);
nand I_3309 (I59181,I59164,I396567);
not I_3310 (I59198,I59181);
nor I_3311 (I58848,I59198,I59133);
nor I_3312 (I59229,I396546,I396564);
or I_3313 (I59246,I59229,I396555);
nor I_3314 (I59263,I396555,I396561);
nand I_3315 (I59280,I59263,I59246);
not I_3316 (I59297,I59280);
nor I_3317 (I59314,I59297,I58941);
or I_3318 (I59331,I59314,I59181);
nor I_3319 (I58830,I58907,I59331);
nor I_3320 (I59362,I59297,I396549);
DFFARX1 I_3321 (I59362,I2898,I58856,I58833,);
nor I_3322 (I59393,I59297,I59181);
nor I_3323 (I58839,I59102,I59393);
nor I_3324 (I59424,I59181,I59280);
nor I_3325 (I58827,I58958,I59424);
not I_3326 (I59485,I2905);
nor I_3327 (I59502,I298847,I298862);
nor I_3328 (I59519,I59502,I298853);
not I_3329 (I59536,I59519);
not I_3330 (I59553,I298859);
nor I_3331 (I59570,I59553,I59502);
not I_3332 (I59587,I59570);
nand I_3333 (I59465,I59536,I59587);
nand I_3334 (I59618,I59519,I298871);
not I_3335 (I59450,I59618);
nor I_3336 (I59474,I59570,I298871);
not I_3337 (I59663,I298868);
nand I_3338 (I59680,I298856,I298847);
nand I_3339 (I59697,I59680,I59663);
nand I_3340 (I59714,I59680,I298868);
not I_3341 (I59731,I59714);
nor I_3342 (I59453,I59731,I59618);
nor I_3343 (I59762,I59731,I298871);
nand I_3344 (I59471,I59536,I59714);
and I_3345 (I59793,I59697,I298844);
nand I_3346 (I59810,I59793,I298874);
not I_3347 (I59827,I59810);
nor I_3348 (I59477,I59827,I59762);
nor I_3349 (I59858,I298844,I298850);
or I_3350 (I59875,I59858,I298865);
nor I_3351 (I59892,I298850,I298853);
nand I_3352 (I59909,I59892,I59875);
not I_3353 (I59926,I59909);
nor I_3354 (I59943,I59926,I59570);
or I_3355 (I59960,I59943,I59810);
nor I_3356 (I59459,I59536,I59960);
nor I_3357 (I59991,I59926,I298871);
DFFARX1 I_3358 (I59991,I2898,I59485,I59462,);
nor I_3359 (I60022,I59926,I59810);
nor I_3360 (I59468,I59731,I60022);
nor I_3361 (I60053,I59810,I59909);
nor I_3362 (I59456,I59587,I60053);
not I_3363 (I60114,I2905);
nor I_3364 (I60131,I397229,I397238);
nor I_3365 (I60148,I60131,I397232);
not I_3366 (I60165,I60148);
not I_3367 (I60182,I397223);
nor I_3368 (I60199,I60182,I60131);
not I_3369 (I60216,I60199);
nand I_3370 (I60094,I60165,I60216);
nand I_3371 (I60247,I60148,I397229);
not I_3372 (I60079,I60247);
nor I_3373 (I60103,I60199,I397229);
not I_3374 (I60292,I397238);
nand I_3375 (I60309,I397223,I397226);
nand I_3376 (I60326,I60309,I60292);
nand I_3377 (I60343,I60309,I397238);
not I_3378 (I60360,I60343);
nor I_3379 (I60082,I60360,I60247);
nor I_3380 (I60391,I60360,I397229);
nand I_3381 (I60100,I60165,I60343);
and I_3382 (I60422,I60326,I397232);
nand I_3383 (I60439,I60422,I397247);
not I_3384 (I60456,I60439);
nor I_3385 (I60106,I60456,I60391);
nor I_3386 (I60487,I397226,I397244);
or I_3387 (I60504,I60487,I397235);
nor I_3388 (I60521,I397235,I397241);
nand I_3389 (I60538,I60521,I60504);
not I_3390 (I60555,I60538);
nor I_3391 (I60572,I60555,I60199);
or I_3392 (I60589,I60572,I60439);
nor I_3393 (I60088,I60165,I60589);
nor I_3394 (I60620,I60555,I397229);
DFFARX1 I_3395 (I60620,I2898,I60114,I60091,);
nor I_3396 (I60651,I60555,I60439);
nor I_3397 (I60097,I60360,I60651);
nor I_3398 (I60682,I60439,I60538);
nor I_3399 (I60085,I60216,I60682);
not I_3400 (I60743,I2905);
nor I_3401 (I60760,I271188,I271188);
nor I_3402 (I60777,I60760,I271197);
not I_3403 (I60794,I60777);
not I_3404 (I60811,I271185);
nor I_3405 (I60828,I60811,I60760);
not I_3406 (I60845,I60828);
nand I_3407 (I60723,I60794,I60845);
nand I_3408 (I60876,I60777,I271206);
not I_3409 (I60708,I60876);
nor I_3410 (I60732,I60828,I271206);
not I_3411 (I60921,I271212);
nand I_3412 (I60938,I271215,I271203);
nand I_3413 (I60955,I60938,I60921);
nand I_3414 (I60972,I60938,I271212);
not I_3415 (I60989,I60972);
nor I_3416 (I60711,I60989,I60876);
nor I_3417 (I61020,I60989,I271206);
nand I_3418 (I60729,I60794,I60972);
and I_3419 (I61051,I60955,I271209);
nand I_3420 (I61068,I61051,I271185);
not I_3421 (I61085,I61068);
nor I_3422 (I60735,I61085,I61020);
nor I_3423 (I61116,I271191,I271194);
or I_3424 (I61133,I61116,I271194);
nor I_3425 (I61150,I271200,I271191);
nand I_3426 (I61167,I61150,I61133);
not I_3427 (I61184,I61167);
nor I_3428 (I61201,I61184,I60828);
or I_3429 (I61218,I61201,I61068);
nor I_3430 (I60717,I60794,I61218);
nor I_3431 (I61249,I61184,I271206);
DFFARX1 I_3432 (I61249,I2898,I60743,I60720,);
nor I_3433 (I61280,I61184,I61068);
nor I_3434 (I60726,I60989,I61280);
nor I_3435 (I61311,I61068,I61167);
nor I_3436 (I60714,I60845,I61311);
not I_3437 (I61372,I2905);
nor I_3438 (I61389,I38218,I38212);
nor I_3439 (I61406,I61389,I38200);
not I_3440 (I61423,I61406);
not I_3441 (I61440,I38203);
nor I_3442 (I61457,I61440,I61389);
not I_3443 (I61474,I61457);
nand I_3444 (I61352,I61423,I61474);
nand I_3445 (I61505,I61406,I38206);
not I_3446 (I61337,I61505);
nor I_3447 (I61361,I61457,I38206);
not I_3448 (I61550,I38215);
nand I_3449 (I61567,I38209,I38203);
nand I_3450 (I61584,I61567,I61550);
nand I_3451 (I61601,I61567,I38215);
not I_3452 (I61618,I61601);
nor I_3453 (I61340,I61618,I61505);
nor I_3454 (I61649,I61618,I38206);
nand I_3455 (I61358,I61423,I61601);
and I_3456 (I61680,I61584,I38212);
nand I_3457 (I61697,I61680,I38209);
not I_3458 (I61714,I61697);
nor I_3459 (I61364,I61714,I61649);
nor I_3460 (I61745,I38227,I38200);
or I_3461 (I61762,I61745,I38221);
nor I_3462 (I61779,I38224,I38206);
nand I_3463 (I61796,I61779,I61762);
not I_3464 (I61813,I61796);
nor I_3465 (I61830,I61813,I61457);
or I_3466 (I61847,I61830,I61697);
nor I_3467 (I61346,I61423,I61847);
nor I_3468 (I61878,I61813,I38206);
DFFARX1 I_3469 (I61878,I2898,I61372,I61349,);
nor I_3470 (I61909,I61813,I61697);
nor I_3471 (I61355,I61618,I61909);
nor I_3472 (I61940,I61697,I61796);
nor I_3473 (I61343,I61474,I61940);
not I_3474 (I62001,I2905);
nor I_3475 (I62018,I379694,I379679);
nor I_3476 (I62035,I62018,I379709);
not I_3477 (I62052,I62035);
not I_3478 (I62069,I379706);
nor I_3479 (I62086,I62069,I62018);
not I_3480 (I62103,I62086);
nand I_3481 (I61981,I62052,I62103);
nand I_3482 (I62134,I62035,I379700);
not I_3483 (I61966,I62134);
nor I_3484 (I61990,I62086,I379700);
not I_3485 (I62179,I379697);
nand I_3486 (I62196,I379679,I379682);
nand I_3487 (I62213,I62196,I62179);
nand I_3488 (I62230,I62196,I379697);
not I_3489 (I62247,I62230);
nor I_3490 (I61969,I62247,I62134);
nor I_3491 (I62278,I62247,I379700);
nand I_3492 (I61987,I62052,I62230);
and I_3493 (I62309,I62213,I379682);
nand I_3494 (I62326,I62309,I379685);
not I_3495 (I62343,I62326);
nor I_3496 (I61993,I62343,I62278);
nor I_3497 (I62374,I379712,I379688);
or I_3498 (I62391,I62374,I379685);
nor I_3499 (I62408,I379703,I379691);
nand I_3500 (I62425,I62408,I62391);
not I_3501 (I62442,I62425);
nor I_3502 (I62459,I62442,I62086);
or I_3503 (I62476,I62459,I62326);
nor I_3504 (I61975,I62052,I62476);
nor I_3505 (I62507,I62442,I379700);
DFFARX1 I_3506 (I62507,I2898,I62001,I61978,);
nor I_3507 (I62538,I62442,I62326);
nor I_3508 (I61984,I62247,I62538);
nor I_3509 (I62569,I62326,I62425);
nor I_3510 (I61972,I62103,I62569);
not I_3511 (I62630,I2905);
nor I_3512 (I62647,I26794,I26788);
nor I_3513 (I62664,I62647,I26776);
not I_3514 (I62681,I62664);
not I_3515 (I62698,I26779);
nor I_3516 (I62715,I62698,I62647);
not I_3517 (I62732,I62715);
nand I_3518 (I62610,I62681,I62732);
nand I_3519 (I62763,I62664,I26782);
not I_3520 (I62595,I62763);
nor I_3521 (I62619,I62715,I26782);
not I_3522 (I62808,I26791);
nand I_3523 (I62825,I26785,I26779);
nand I_3524 (I62842,I62825,I62808);
nand I_3525 (I62859,I62825,I26791);
not I_3526 (I62876,I62859);
nor I_3527 (I62598,I62876,I62763);
nor I_3528 (I62907,I62876,I26782);
nand I_3529 (I62616,I62681,I62859);
and I_3530 (I62938,I62842,I26788);
nand I_3531 (I62955,I62938,I26785);
not I_3532 (I62972,I62955);
nor I_3533 (I62622,I62972,I62907);
nor I_3534 (I63003,I26803,I26776);
or I_3535 (I63020,I63003,I26797);
nor I_3536 (I63037,I26800,I26782);
nand I_3537 (I63054,I63037,I63020);
not I_3538 (I63071,I63054);
nor I_3539 (I63088,I63071,I62715);
or I_3540 (I63105,I63088,I62955);
nor I_3541 (I62604,I62681,I63105);
nor I_3542 (I63136,I63071,I26782);
DFFARX1 I_3543 (I63136,I2898,I62630,I62607,);
nor I_3544 (I63167,I63071,I62955);
nor I_3545 (I62613,I62876,I63167);
nor I_3546 (I63198,I62955,I63054);
nor I_3547 (I62601,I62732,I63198);
not I_3548 (I63259,I2905);
nor I_3549 (I63276,I132378,I132375);
nor I_3550 (I63293,I63276,I132363);
not I_3551 (I63310,I63293);
not I_3552 (I63327,I132390);
nor I_3553 (I63344,I63327,I63276);
not I_3554 (I63361,I63344);
nand I_3555 (I63239,I63310,I63361);
nand I_3556 (I63392,I63293,I132381);
not I_3557 (I63224,I63392);
nor I_3558 (I63248,I63344,I132381);
not I_3559 (I63437,I132366);
nand I_3560 (I63454,I132384,I132363);
nand I_3561 (I63471,I63454,I63437);
nand I_3562 (I63488,I63454,I132366);
not I_3563 (I63505,I63488);
nor I_3564 (I63227,I63505,I63392);
nor I_3565 (I63536,I63505,I132381);
nand I_3566 (I63245,I63310,I63488);
and I_3567 (I63567,I63471,I132372);
nand I_3568 (I63584,I63567,I132369);
not I_3569 (I63601,I63584);
nor I_3570 (I63251,I63601,I63536);
nor I_3571 (I63632,I132369,I132396);
or I_3572 (I63649,I63632,I132366);
nor I_3573 (I63666,I132387,I132393);
nand I_3574 (I63683,I63666,I63649);
not I_3575 (I63700,I63683);
nor I_3576 (I63717,I63700,I63344);
or I_3577 (I63734,I63717,I63584);
nor I_3578 (I63233,I63310,I63734);
nor I_3579 (I63765,I63700,I132381);
DFFARX1 I_3580 (I63765,I2898,I63259,I63236,);
nor I_3581 (I63796,I63700,I63584);
nor I_3582 (I63242,I63505,I63796);
nor I_3583 (I63827,I63584,I63683);
nor I_3584 (I63230,I63361,I63827);
not I_3585 (I63888,I2905);
nor I_3586 (I63905,I244413,I244413);
nor I_3587 (I63922,I63905,I244422);
not I_3588 (I63939,I63922);
not I_3589 (I63956,I244410);
nor I_3590 (I63973,I63956,I63905);
not I_3591 (I63990,I63973);
nand I_3592 (I63868,I63939,I63990);
nand I_3593 (I64021,I63922,I244431);
not I_3594 (I63853,I64021);
nor I_3595 (I63877,I63973,I244431);
not I_3596 (I64066,I244437);
nand I_3597 (I64083,I244440,I244428);
nand I_3598 (I64100,I64083,I64066);
nand I_3599 (I64117,I64083,I244437);
not I_3600 (I64134,I64117);
nor I_3601 (I63856,I64134,I64021);
nor I_3602 (I64165,I64134,I244431);
nand I_3603 (I63874,I63939,I64117);
and I_3604 (I64196,I64100,I244434);
nand I_3605 (I64213,I64196,I244410);
not I_3606 (I64230,I64213);
nor I_3607 (I63880,I64230,I64165);
nor I_3608 (I64261,I244416,I244419);
or I_3609 (I64278,I64261,I244419);
nor I_3610 (I64295,I244425,I244416);
nand I_3611 (I64312,I64295,I64278);
not I_3612 (I64329,I64312);
nor I_3613 (I64346,I64329,I63973);
or I_3614 (I64363,I64346,I64213);
nor I_3615 (I63862,I63939,I64363);
nor I_3616 (I64394,I64329,I244431);
DFFARX1 I_3617 (I64394,I2898,I63888,I63865,);
nor I_3618 (I64425,I64329,I64213);
nor I_3619 (I63871,I64134,I64425);
nor I_3620 (I64456,I64213,I64312);
nor I_3621 (I63859,I63990,I64456);
not I_3622 (I64517,I2905);
nor I_3623 (I64534,I285689,I285704);
nor I_3624 (I64551,I64534,I285695);
not I_3625 (I64568,I64551);
not I_3626 (I64585,I285701);
nor I_3627 (I64602,I64585,I64534);
not I_3628 (I64619,I64602);
nand I_3629 (I64497,I64568,I64619);
nand I_3630 (I64650,I64551,I285713);
not I_3631 (I64482,I64650);
nor I_3632 (I64506,I64602,I285713);
not I_3633 (I64695,I285710);
nand I_3634 (I64712,I285698,I285689);
nand I_3635 (I64729,I64712,I64695);
nand I_3636 (I64746,I64712,I285710);
not I_3637 (I64763,I64746);
nor I_3638 (I64485,I64763,I64650);
nor I_3639 (I64794,I64763,I285713);
nand I_3640 (I64503,I64568,I64746);
and I_3641 (I64825,I64729,I285686);
nand I_3642 (I64842,I64825,I285716);
not I_3643 (I64859,I64842);
nor I_3644 (I64509,I64859,I64794);
nor I_3645 (I64890,I285686,I285692);
or I_3646 (I64907,I64890,I285707);
nor I_3647 (I64924,I285692,I285695);
nand I_3648 (I64941,I64924,I64907);
not I_3649 (I64958,I64941);
nor I_3650 (I64975,I64958,I64602);
or I_3651 (I64992,I64975,I64842);
nor I_3652 (I64491,I64568,I64992);
nor I_3653 (I65023,I64958,I285713);
DFFARX1 I_3654 (I65023,I2898,I64517,I64494,);
nor I_3655 (I65054,I64958,I64842);
nor I_3656 (I64500,I64763,I65054);
nor I_3657 (I65085,I64842,I64941);
nor I_3658 (I64488,I64619,I65085);
not I_3659 (I65146,I2905);
nor I_3660 (I65163,I398589,I398598);
nor I_3661 (I65180,I65163,I398592);
not I_3662 (I65197,I65180);
not I_3663 (I65214,I398583);
nor I_3664 (I65231,I65214,I65163);
not I_3665 (I65248,I65231);
nand I_3666 (I65126,I65197,I65248);
nand I_3667 (I65279,I65180,I398589);
not I_3668 (I65111,I65279);
nor I_3669 (I65135,I65231,I398589);
not I_3670 (I65324,I398598);
nand I_3671 (I65341,I398583,I398586);
nand I_3672 (I65358,I65341,I65324);
nand I_3673 (I65375,I65341,I398598);
not I_3674 (I65392,I65375);
nor I_3675 (I65114,I65392,I65279);
nor I_3676 (I65423,I65392,I398589);
nand I_3677 (I65132,I65197,I65375);
and I_3678 (I65454,I65358,I398592);
nand I_3679 (I65471,I65454,I398607);
not I_3680 (I65488,I65471);
nor I_3681 (I65138,I65488,I65423);
nor I_3682 (I65519,I398586,I398604);
or I_3683 (I65536,I65519,I398595);
nor I_3684 (I65553,I398595,I398601);
nand I_3685 (I65570,I65553,I65536);
not I_3686 (I65587,I65570);
nor I_3687 (I65604,I65587,I65231);
or I_3688 (I65621,I65604,I65471);
nor I_3689 (I65120,I65197,I65621);
nor I_3690 (I65652,I65587,I398589);
DFFARX1 I_3691 (I65652,I2898,I65146,I65123,);
nor I_3692 (I65683,I65587,I65471);
nor I_3693 (I65129,I65392,I65683);
nor I_3694 (I65714,I65471,I65570);
nor I_3695 (I65117,I65248,I65714);
not I_3696 (I65775,I2905);
nor I_3697 (I65792,I317853,I317868);
nor I_3698 (I65809,I65792,I317859);
not I_3699 (I65826,I65809);
not I_3700 (I65843,I317865);
nor I_3701 (I65860,I65843,I65792);
not I_3702 (I65877,I65860);
nand I_3703 (I65755,I65826,I65877);
nand I_3704 (I65908,I65809,I317877);
not I_3705 (I65740,I65908);
nor I_3706 (I65764,I65860,I317877);
not I_3707 (I65953,I317874);
nand I_3708 (I65970,I317862,I317853);
nand I_3709 (I65987,I65970,I65953);
nand I_3710 (I66004,I65970,I317874);
not I_3711 (I66021,I66004);
nor I_3712 (I65743,I66021,I65908);
nor I_3713 (I66052,I66021,I317877);
nand I_3714 (I65761,I65826,I66004);
and I_3715 (I66083,I65987,I317850);
nand I_3716 (I66100,I66083,I317880);
not I_3717 (I66117,I66100);
nor I_3718 (I65767,I66117,I66052);
nor I_3719 (I66148,I317850,I317856);
or I_3720 (I66165,I66148,I317871);
nor I_3721 (I66182,I317856,I317859);
nand I_3722 (I66199,I66182,I66165);
not I_3723 (I66216,I66199);
nor I_3724 (I66233,I66216,I65860);
or I_3725 (I66250,I66233,I66100);
nor I_3726 (I65749,I65826,I66250);
nor I_3727 (I66281,I66216,I317877);
DFFARX1 I_3728 (I66281,I2898,I65775,I65752,);
nor I_3729 (I66312,I66216,I66100);
nor I_3730 (I65758,I66021,I66312);
nor I_3731 (I66343,I66100,I66199);
nor I_3732 (I65746,I65877,I66343);
not I_3733 (I66404,I2905);
nor I_3734 (I66421,I234468,I234468);
nor I_3735 (I66438,I66421,I234477);
not I_3736 (I66455,I66438);
not I_3737 (I66472,I234465);
nor I_3738 (I66489,I66472,I66421);
not I_3739 (I66506,I66489);
nand I_3740 (I66384,I66455,I66506);
nand I_3741 (I66537,I66438,I234486);
not I_3742 (I66369,I66537);
nor I_3743 (I66393,I66489,I234486);
not I_3744 (I66582,I234492);
nand I_3745 (I66599,I234495,I234483);
nand I_3746 (I66616,I66599,I66582);
nand I_3747 (I66633,I66599,I234492);
not I_3748 (I66650,I66633);
nor I_3749 (I66372,I66650,I66537);
nor I_3750 (I66681,I66650,I234486);
nand I_3751 (I66390,I66455,I66633);
and I_3752 (I66712,I66616,I234489);
nand I_3753 (I66729,I66712,I234465);
not I_3754 (I66746,I66729);
nor I_3755 (I66396,I66746,I66681);
nor I_3756 (I66777,I234471,I234474);
or I_3757 (I66794,I66777,I234474);
nor I_3758 (I66811,I234480,I234471);
nand I_3759 (I66828,I66811,I66794);
not I_3760 (I66845,I66828);
nor I_3761 (I66862,I66845,I66489);
or I_3762 (I66879,I66862,I66729);
nor I_3763 (I66378,I66455,I66879);
nor I_3764 (I66910,I66845,I234486);
DFFARX1 I_3765 (I66910,I2898,I66404,I66381,);
nor I_3766 (I66941,I66845,I66729);
nor I_3767 (I66387,I66650,I66941);
nor I_3768 (I66972,I66729,I66828);
nor I_3769 (I66375,I66506,I66972);
not I_3770 (I67033,I2905);
nor I_3771 (I67050,I125459,I125456);
nor I_3772 (I67067,I67050,I125444);
not I_3773 (I67084,I67067);
not I_3774 (I67101,I125471);
nor I_3775 (I67118,I67101,I67050);
not I_3776 (I67135,I67118);
nand I_3777 (I67013,I67084,I67135);
nand I_3778 (I67166,I67067,I125462);
not I_3779 (I66998,I67166);
nor I_3780 (I67022,I67118,I125462);
not I_3781 (I67211,I125447);
nand I_3782 (I67228,I125465,I125444);
nand I_3783 (I67245,I67228,I67211);
nand I_3784 (I67262,I67228,I125447);
not I_3785 (I67279,I67262);
nor I_3786 (I67001,I67279,I67166);
nor I_3787 (I67310,I67279,I125462);
nand I_3788 (I67019,I67084,I67262);
and I_3789 (I67341,I67245,I125453);
nand I_3790 (I67358,I67341,I125450);
not I_3791 (I67375,I67358);
nor I_3792 (I67025,I67375,I67310);
nor I_3793 (I67406,I125450,I125477);
or I_3794 (I67423,I67406,I125447);
nor I_3795 (I67440,I125468,I125474);
nand I_3796 (I67457,I67440,I67423);
not I_3797 (I67474,I67457);
nor I_3798 (I67491,I67474,I67118);
or I_3799 (I67508,I67491,I67358);
nor I_3800 (I67007,I67084,I67508);
nor I_3801 (I67539,I67474,I125462);
DFFARX1 I_3802 (I67539,I2898,I67033,I67010,);
nor I_3803 (I67570,I67474,I67358);
nor I_3804 (I67016,I67279,I67570);
nor I_3805 (I67601,I67358,I67457);
nor I_3806 (I67004,I67135,I67601);
not I_3807 (I67662,I2905);
nor I_3808 (I67679,I18940,I18934);
nor I_3809 (I67696,I67679,I18922);
not I_3810 (I67713,I67696);
not I_3811 (I67730,I18925);
nor I_3812 (I67747,I67730,I67679);
not I_3813 (I67764,I67747);
nand I_3814 (I67642,I67713,I67764);
nand I_3815 (I67795,I67696,I18928);
not I_3816 (I67627,I67795);
nor I_3817 (I67651,I67747,I18928);
not I_3818 (I67840,I18937);
nand I_3819 (I67857,I18931,I18925);
nand I_3820 (I67874,I67857,I67840);
nand I_3821 (I67891,I67857,I18937);
not I_3822 (I67908,I67891);
nor I_3823 (I67630,I67908,I67795);
nor I_3824 (I67939,I67908,I18928);
nand I_3825 (I67648,I67713,I67891);
and I_3826 (I67970,I67874,I18934);
nand I_3827 (I67987,I67970,I18931);
not I_3828 (I68004,I67987);
nor I_3829 (I67654,I68004,I67939);
nor I_3830 (I68035,I18949,I18922);
or I_3831 (I68052,I68035,I18943);
nor I_3832 (I68069,I18946,I18928);
nand I_3833 (I68086,I68069,I68052);
not I_3834 (I68103,I68086);
nor I_3835 (I68120,I68103,I67747);
or I_3836 (I68137,I68120,I67987);
nor I_3837 (I67636,I67713,I68137);
nor I_3838 (I68168,I68103,I18928);
DFFARX1 I_3839 (I68168,I2898,I67662,I67639,);
nor I_3840 (I68199,I68103,I67987);
nor I_3841 (I67645,I67908,I68199);
nor I_3842 (I68230,I67987,I68086);
nor I_3843 (I67633,I67764,I68230);
not I_3844 (I68291,I2905);
nor I_3845 (I68308,I412926,I412929);
nor I_3846 (I68325,I68308,I412947);
not I_3847 (I68342,I68325);
not I_3848 (I68359,I412920);
nor I_3849 (I68376,I68359,I68308);
not I_3850 (I68393,I68376);
nand I_3851 (I68271,I68342,I68393);
nand I_3852 (I68424,I68325,I412917);
not I_3853 (I68256,I68424);
nor I_3854 (I68280,I68376,I412917);
not I_3855 (I68469,I412914);
nand I_3856 (I68486,I412944,I412923);
nand I_3857 (I68503,I68486,I68469);
nand I_3858 (I68520,I68486,I412914);
not I_3859 (I68537,I68520);
nor I_3860 (I68259,I68537,I68424);
nor I_3861 (I68568,I68537,I412917);
nand I_3862 (I68277,I68342,I68520);
and I_3863 (I68599,I68503,I412935);
nand I_3864 (I68616,I68599,I412941);
not I_3865 (I68633,I68616);
nor I_3866 (I68283,I68633,I68568);
nor I_3867 (I68664,I412932,I412920);
or I_3868 (I68681,I68664,I412917);
nor I_3869 (I68698,I412914,I412938);
nand I_3870 (I68715,I68698,I68681);
not I_3871 (I68732,I68715);
nor I_3872 (I68749,I68732,I68376);
or I_3873 (I68766,I68749,I68616);
nor I_3874 (I68265,I68342,I68766);
nor I_3875 (I68797,I68732,I412917);
DFFARX1 I_3876 (I68797,I2898,I68291,I68268,);
nor I_3877 (I68828,I68732,I68616);
nor I_3878 (I68274,I68537,I68828);
nor I_3879 (I68859,I68616,I68715);
nor I_3880 (I68262,I68393,I68859);
not I_3881 (I68920,I2905);
nor I_3882 (I68937,I404709,I404718);
nor I_3883 (I68954,I68937,I404712);
not I_3884 (I68971,I68954);
not I_3885 (I68988,I404703);
nor I_3886 (I69005,I68988,I68937);
not I_3887 (I69022,I69005);
nand I_3888 (I68900,I68971,I69022);
nand I_3889 (I69053,I68954,I404709);
not I_3890 (I68885,I69053);
nor I_3891 (I68909,I69005,I404709);
not I_3892 (I69098,I404718);
nand I_3893 (I69115,I404703,I404706);
nand I_3894 (I69132,I69115,I69098);
nand I_3895 (I69149,I69115,I404718);
not I_3896 (I69166,I69149);
nor I_3897 (I68888,I69166,I69053);
nor I_3898 (I69197,I69166,I404709);
nand I_3899 (I68906,I68971,I69149);
and I_3900 (I69228,I69132,I404712);
nand I_3901 (I69245,I69228,I404727);
not I_3902 (I69262,I69245);
nor I_3903 (I68912,I69262,I69197);
nor I_3904 (I69293,I404706,I404724);
or I_3905 (I69310,I69293,I404715);
nor I_3906 (I69327,I404715,I404721);
nand I_3907 (I69344,I69327,I69310);
not I_3908 (I69361,I69344);
nor I_3909 (I69378,I69361,I69005);
or I_3910 (I69395,I69378,I69245);
nor I_3911 (I68894,I68971,I69395);
nor I_3912 (I69426,I69361,I404709);
DFFARX1 I_3913 (I69426,I2898,I68920,I68897,);
nor I_3914 (I69457,I69361,I69245);
nor I_3915 (I68903,I69166,I69457);
nor I_3916 (I69488,I69245,I69344);
nor I_3917 (I68891,I69022,I69488);
not I_3918 (I69549,I2905);
nor I_3919 (I69566,I328781,I328793);
nor I_3920 (I69583,I69566,I328784);
not I_3921 (I69600,I69583);
not I_3922 (I69617,I328796);
nor I_3923 (I69634,I69617,I69566);
not I_3924 (I69651,I69634);
nand I_3925 (I69529,I69600,I69651);
nand I_3926 (I69682,I69583,I328805);
not I_3927 (I69514,I69682);
nor I_3928 (I69538,I69634,I328805);
not I_3929 (I69727,I328793);
nand I_3930 (I69744,I328787,I328787);
nand I_3931 (I69761,I69744,I69727);
nand I_3932 (I69778,I69744,I328793);
not I_3933 (I69795,I69778);
nor I_3934 (I69517,I69795,I69682);
nor I_3935 (I69826,I69795,I328805);
nand I_3936 (I69535,I69600,I69778);
and I_3937 (I69857,I69761,I328784);
nand I_3938 (I69874,I69857,I328802);
not I_3939 (I69891,I69874);
nor I_3940 (I69541,I69891,I69826);
nor I_3941 (I69922,I328799,I328781);
or I_3942 (I69939,I69922,I328790);
nor I_3943 (I69956,I328790,I328796);
nand I_3944 (I69973,I69956,I69939);
not I_3945 (I69990,I69973);
nor I_3946 (I70007,I69990,I69634);
or I_3947 (I70024,I70007,I69874);
nor I_3948 (I69523,I69600,I70024);
nor I_3949 (I70055,I69990,I328805);
DFFARX1 I_3950 (I70055,I2898,I69549,I69526,);
nor I_3951 (I70086,I69990,I69874);
nor I_3952 (I69532,I69795,I70086);
nor I_3953 (I70117,I69874,I69973);
nor I_3954 (I69520,I69651,I70117);
not I_3955 (I70178,I2905);
nor I_3956 (I70195,I226176,I226155);
nor I_3957 (I70212,I70195,I226170);
not I_3958 (I70229,I70212);
not I_3959 (I70246,I226152);
nor I_3960 (I70263,I70246,I70195);
not I_3961 (I70280,I70263);
nand I_3962 (I70158,I70229,I70280);
nand I_3963 (I70311,I70212,I226167);
not I_3964 (I70143,I70311);
nor I_3965 (I70167,I70263,I226167);
not I_3966 (I70356,I226158);
nand I_3967 (I70373,I226164,I226155);
nand I_3968 (I70390,I70373,I70356);
nand I_3969 (I70407,I70373,I226158);
not I_3970 (I70424,I70407);
nor I_3971 (I70146,I70424,I70311);
nor I_3972 (I70455,I70424,I226167);
nand I_3973 (I70164,I70229,I70407);
and I_3974 (I70486,I70390,I226173);
nand I_3975 (I70503,I70486,I226152);
not I_3976 (I70520,I70503);
nor I_3977 (I70170,I70520,I70455);
nor I_3978 (I70551,I226161,I226158);
or I_3979 (I70568,I70551,I226164);
nor I_3980 (I70585,I226161,I226179);
nand I_3981 (I70602,I70585,I70568);
not I_3982 (I70619,I70602);
nor I_3983 (I70636,I70619,I70263);
or I_3984 (I70653,I70636,I70503);
nor I_3985 (I70152,I70229,I70653);
nor I_3986 (I70684,I70619,I226167);
DFFARX1 I_3987 (I70684,I2898,I70178,I70155,);
nor I_3988 (I70715,I70619,I70503);
nor I_3989 (I70161,I70424,I70715);
nor I_3990 (I70746,I70503,I70602);
nor I_3991 (I70149,I70280,I70746);
not I_3992 (I70807,I2905);
nor I_3993 (I70824,I232173,I232173);
nor I_3994 (I70841,I70824,I232182);
not I_3995 (I70858,I70841);
not I_3996 (I70875,I232170);
nor I_3997 (I70892,I70875,I70824);
not I_3998 (I70909,I70892);
nand I_3999 (I70787,I70858,I70909);
nand I_4000 (I70940,I70841,I232191);
not I_4001 (I70772,I70940);
nor I_4002 (I70796,I70892,I232191);
not I_4003 (I70985,I232197);
nand I_4004 (I71002,I232200,I232188);
nand I_4005 (I71019,I71002,I70985);
nand I_4006 (I71036,I71002,I232197);
not I_4007 (I71053,I71036);
nor I_4008 (I70775,I71053,I70940);
nor I_4009 (I71084,I71053,I232191);
nand I_4010 (I70793,I70858,I71036);
and I_4011 (I71115,I71019,I232194);
nand I_4012 (I71132,I71115,I232170);
not I_4013 (I71149,I71132);
nor I_4014 (I70799,I71149,I71084);
nor I_4015 (I71180,I232176,I232179);
or I_4016 (I71197,I71180,I232179);
nor I_4017 (I71214,I232185,I232176);
nand I_4018 (I71231,I71214,I71197);
not I_4019 (I71248,I71231);
nor I_4020 (I71265,I71248,I70892);
or I_4021 (I71282,I71265,I71132);
nor I_4022 (I70781,I70858,I71282);
nor I_4023 (I71313,I71248,I232191);
DFFARX1 I_4024 (I71313,I2898,I70807,I70784,);
nor I_4025 (I71344,I71248,I71132);
nor I_4026 (I70790,I71053,I71344);
nor I_4027 (I71375,I71132,I71231);
nor I_4028 (I70778,I70909,I71375);
not I_4029 (I71436,I2905);
nor I_4030 (I71453,I111621,I111618);
nor I_4031 (I71470,I71453,I111606);
not I_4032 (I71487,I71470);
not I_4033 (I71504,I111633);
nor I_4034 (I71521,I71504,I71453);
not I_4035 (I71538,I71521);
nand I_4036 (I71416,I71487,I71538);
nand I_4037 (I71569,I71470,I111624);
not I_4038 (I71401,I71569);
nor I_4039 (I71425,I71521,I111624);
not I_4040 (I71614,I111609);
nand I_4041 (I71631,I111627,I111606);
nand I_4042 (I71648,I71631,I71614);
nand I_4043 (I71665,I71631,I111609);
not I_4044 (I71682,I71665);
nor I_4045 (I71404,I71682,I71569);
nor I_4046 (I71713,I71682,I111624);
nand I_4047 (I71422,I71487,I71665);
and I_4048 (I71744,I71648,I111615);
nand I_4049 (I71761,I71744,I111612);
not I_4050 (I71778,I71761);
nor I_4051 (I71428,I71778,I71713);
nor I_4052 (I71809,I111612,I111639);
or I_4053 (I71826,I71809,I111609);
nor I_4054 (I71843,I111630,I111636);
nand I_4055 (I71860,I71843,I71826);
not I_4056 (I71877,I71860);
nor I_4057 (I71894,I71877,I71521);
or I_4058 (I71911,I71894,I71761);
nor I_4059 (I71410,I71487,I71911);
nor I_4060 (I71942,I71877,I111624);
DFFARX1 I_4061 (I71942,I2898,I71436,I71413,);
nor I_4062 (I71973,I71877,I71761);
nor I_4063 (I71419,I71682,I71973);
nor I_4064 (I72004,I71761,I71860);
nor I_4065 (I71407,I71538,I72004);
not I_4066 (I72065,I2905);
nor I_4067 (I72082,I151132,I151123);
nor I_4068 (I72099,I72082,I151117);
not I_4069 (I72116,I72099);
not I_4070 (I72133,I151129);
nor I_4071 (I72150,I72133,I72082);
not I_4072 (I72167,I72150);
nand I_4073 (I72045,I72116,I72167);
nand I_4074 (I72198,I72099,I151141);
not I_4075 (I72030,I72198);
nor I_4076 (I72054,I72150,I151141);
not I_4077 (I72243,I151138);
nand I_4078 (I72260,I151147,I151120);
nand I_4079 (I72277,I72260,I72243);
nand I_4080 (I72294,I72260,I151138);
not I_4081 (I72311,I72294);
nor I_4082 (I72033,I72311,I72198);
nor I_4083 (I72342,I72311,I151141);
nand I_4084 (I72051,I72116,I72294);
and I_4085 (I72373,I72277,I151126);
nand I_4086 (I72390,I72373,I151114);
not I_4087 (I72407,I72390);
nor I_4088 (I72057,I72407,I72342);
nor I_4089 (I72438,I151144,I151135);
or I_4090 (I72455,I72438,I151117);
nor I_4091 (I72472,I151114,I151120);
nand I_4092 (I72489,I72472,I72455);
not I_4093 (I72506,I72489);
nor I_4094 (I72523,I72506,I72150);
or I_4095 (I72540,I72523,I72390);
nor I_4096 (I72039,I72116,I72540);
nor I_4097 (I72571,I72506,I151141);
DFFARX1 I_4098 (I72571,I2898,I72065,I72042,);
nor I_4099 (I72602,I72506,I72390);
nor I_4100 (I72048,I72311,I72602);
nor I_4101 (I72633,I72390,I72489);
nor I_4102 (I72036,I72167,I72633);
not I_4103 (I72694,I2905);
nor I_4104 (I72711,I331161,I331173);
nor I_4105 (I72728,I72711,I331164);
not I_4106 (I72745,I72728);
not I_4107 (I72762,I331176);
nor I_4108 (I72779,I72762,I72711);
not I_4109 (I72796,I72779);
nand I_4110 (I72674,I72745,I72796);
nand I_4111 (I72827,I72728,I331185);
not I_4112 (I72659,I72827);
nor I_4113 (I72683,I72779,I331185);
not I_4114 (I72872,I331173);
nand I_4115 (I72889,I331167,I331167);
nand I_4116 (I72906,I72889,I72872);
nand I_4117 (I72923,I72889,I331173);
not I_4118 (I72940,I72923);
nor I_4119 (I72662,I72940,I72827);
nor I_4120 (I72971,I72940,I331185);
nand I_4121 (I72680,I72745,I72923);
and I_4122 (I73002,I72906,I331164);
nand I_4123 (I73019,I73002,I331182);
not I_4124 (I73036,I73019);
nor I_4125 (I72686,I73036,I72971);
nor I_4126 (I73067,I331179,I331161);
or I_4127 (I73084,I73067,I331170);
nor I_4128 (I73101,I331170,I331176);
nand I_4129 (I73118,I73101,I73084);
not I_4130 (I73135,I73118);
nor I_4131 (I73152,I73135,I72779);
or I_4132 (I73169,I73152,I73019);
nor I_4133 (I72668,I72745,I73169);
nor I_4134 (I73200,I73135,I331185);
DFFARX1 I_4135 (I73200,I2898,I72694,I72671,);
nor I_4136 (I73231,I73135,I73019);
nor I_4137 (I72677,I72940,I73231);
nor I_4138 (I73262,I73019,I73118);
nor I_4139 (I72665,I72796,I73262);
not I_4140 (I73323,I2905);
nor I_4141 (I73340,I129862,I129859);
nor I_4142 (I73357,I73340,I129847);
not I_4143 (I73374,I73357);
not I_4144 (I73391,I129874);
nor I_4145 (I73408,I73391,I73340);
not I_4146 (I73425,I73408);
nand I_4147 (I73303,I73374,I73425);
nand I_4148 (I73456,I73357,I129865);
not I_4149 (I73288,I73456);
nor I_4150 (I73312,I73408,I129865);
not I_4151 (I73501,I129850);
nand I_4152 (I73518,I129868,I129847);
nand I_4153 (I73535,I73518,I73501);
nand I_4154 (I73552,I73518,I129850);
not I_4155 (I73569,I73552);
nor I_4156 (I73291,I73569,I73456);
nor I_4157 (I73600,I73569,I129865);
nand I_4158 (I73309,I73374,I73552);
and I_4159 (I73631,I73535,I129856);
nand I_4160 (I73648,I73631,I129853);
not I_4161 (I73665,I73648);
nor I_4162 (I73315,I73665,I73600);
nor I_4163 (I73696,I129853,I129880);
or I_4164 (I73713,I73696,I129850);
nor I_4165 (I73730,I129871,I129877);
nand I_4166 (I73747,I73730,I73713);
not I_4167 (I73764,I73747);
nor I_4168 (I73781,I73764,I73408);
or I_4169 (I73798,I73781,I73648);
nor I_4170 (I73297,I73374,I73798);
nor I_4171 (I73829,I73764,I129865);
DFFARX1 I_4172 (I73829,I2898,I73323,I73300,);
nor I_4173 (I73860,I73764,I73648);
nor I_4174 (I73306,I73569,I73860);
nor I_4175 (I73891,I73648,I73747);
nor I_4176 (I73294,I73425,I73891);
not I_4177 (I73952,I2905);
nor I_4178 (I73969,I127975,I127972);
nor I_4179 (I73986,I73969,I127960);
not I_4180 (I74003,I73986);
not I_4181 (I74020,I127987);
nor I_4182 (I74037,I74020,I73969);
not I_4183 (I74054,I74037);
nand I_4184 (I73932,I74003,I74054);
nand I_4185 (I74085,I73986,I127978);
not I_4186 (I73917,I74085);
nor I_4187 (I73941,I74037,I127978);
not I_4188 (I74130,I127963);
nand I_4189 (I74147,I127981,I127960);
nand I_4190 (I74164,I74147,I74130);
nand I_4191 (I74181,I74147,I127963);
not I_4192 (I74198,I74181);
nor I_4193 (I73920,I74198,I74085);
nor I_4194 (I74229,I74198,I127978);
nand I_4195 (I73938,I74003,I74181);
and I_4196 (I74260,I74164,I127969);
nand I_4197 (I74277,I74260,I127966);
not I_4198 (I74294,I74277);
nor I_4199 (I73944,I74294,I74229);
nor I_4200 (I74325,I127966,I127993);
or I_4201 (I74342,I74325,I127963);
nor I_4202 (I74359,I127984,I127990);
nand I_4203 (I74376,I74359,I74342);
not I_4204 (I74393,I74376);
nor I_4205 (I74410,I74393,I74037);
or I_4206 (I74427,I74410,I74277);
nor I_4207 (I73926,I74003,I74427);
nor I_4208 (I74458,I74393,I127978);
DFFARX1 I_4209 (I74458,I2898,I73952,I73929,);
nor I_4210 (I74489,I74393,I74277);
nor I_4211 (I73935,I74198,I74489);
nor I_4212 (I74520,I74277,I74376);
nor I_4213 (I73923,I74054,I74520);
not I_4214 (I74581,I2905);
nor I_4215 (I74598,I332946,I332958);
nor I_4216 (I74615,I74598,I332949);
not I_4217 (I74632,I74615);
not I_4218 (I74649,I332961);
nor I_4219 (I74666,I74649,I74598);
not I_4220 (I74683,I74666);
nand I_4221 (I74561,I74632,I74683);
nand I_4222 (I74714,I74615,I332970);
not I_4223 (I74546,I74714);
nor I_4224 (I74570,I74666,I332970);
not I_4225 (I74759,I332958);
nand I_4226 (I74776,I332952,I332952);
nand I_4227 (I74793,I74776,I74759);
nand I_4228 (I74810,I74776,I332958);
not I_4229 (I74827,I74810);
nor I_4230 (I74549,I74827,I74714);
nor I_4231 (I74858,I74827,I332970);
nand I_4232 (I74567,I74632,I74810);
and I_4233 (I74889,I74793,I332949);
nand I_4234 (I74906,I74889,I332967);
not I_4235 (I74923,I74906);
nor I_4236 (I74573,I74923,I74858);
nor I_4237 (I74954,I332964,I332946);
or I_4238 (I74971,I74954,I332955);
nor I_4239 (I74988,I332955,I332961);
nand I_4240 (I75005,I74988,I74971);
not I_4241 (I75022,I75005);
nor I_4242 (I75039,I75022,I74666);
or I_4243 (I75056,I75039,I74906);
nor I_4244 (I74555,I74632,I75056);
nor I_4245 (I75087,I75022,I332970);
DFFARX1 I_4246 (I75087,I2898,I74581,I74558,);
nor I_4247 (I75118,I75022,I74906);
nor I_4248 (I74564,I74827,I75118);
nor I_4249 (I75149,I74906,I75005);
nor I_4250 (I74552,I74683,I75149);
not I_4251 (I75210,I2905);
nor I_4252 (I75227,I11485,I11491);
nor I_4253 (I75244,I75227,I11503);
not I_4254 (I75261,I75244);
not I_4255 (I75278,I11500);
nor I_4256 (I75295,I75278,I75227);
not I_4257 (I75312,I75295);
nand I_4258 (I75190,I75261,I75312);
nand I_4259 (I75343,I75244,I11506);
not I_4260 (I75175,I75343);
nor I_4261 (I75199,I75295,I11506);
not I_4262 (I75388,I11482);
nand I_4263 (I75405,I11494,I11476);
nand I_4264 (I75422,I75405,I75388);
nand I_4265 (I75439,I75405,I11482);
not I_4266 (I75456,I75439);
nor I_4267 (I75178,I75456,I75343);
nor I_4268 (I75487,I75456,I11506);
nand I_4269 (I75196,I75261,I75439);
and I_4270 (I75518,I75422,I11488);
nand I_4271 (I75535,I75518,I11485);
not I_4272 (I75552,I75535);
nor I_4273 (I75202,I75552,I75487);
nor I_4274 (I75583,I11482,I11479);
or I_4275 (I75600,I75583,I11479);
nor I_4276 (I75617,I11497,I11476);
nand I_4277 (I75634,I75617,I75600);
not I_4278 (I75651,I75634);
nor I_4279 (I75668,I75651,I75295);
or I_4280 (I75685,I75668,I75535);
nor I_4281 (I75184,I75261,I75685);
nor I_4282 (I75716,I75651,I11506);
DFFARX1 I_4283 (I75716,I2898,I75210,I75187,);
nor I_4284 (I75747,I75651,I75535);
nor I_4285 (I75193,I75456,I75747);
nor I_4286 (I75778,I75535,I75634);
nor I_4287 (I75181,I75312,I75778);
not I_4288 (I75839,I2905);
nor I_4289 (I75856,I150452,I150443);
nor I_4290 (I75873,I75856,I150437);
not I_4291 (I75890,I75873);
not I_4292 (I75907,I150449);
nor I_4293 (I75924,I75907,I75856);
not I_4294 (I75941,I75924);
nand I_4295 (I75819,I75890,I75941);
nand I_4296 (I75972,I75873,I150461);
not I_4297 (I75804,I75972);
nor I_4298 (I75828,I75924,I150461);
not I_4299 (I76017,I150458);
nand I_4300 (I76034,I150467,I150440);
nand I_4301 (I76051,I76034,I76017);
nand I_4302 (I76068,I76034,I150458);
not I_4303 (I76085,I76068);
nor I_4304 (I75807,I76085,I75972);
nor I_4305 (I76116,I76085,I150461);
nand I_4306 (I75825,I75890,I76068);
and I_4307 (I76147,I76051,I150446);
nand I_4308 (I76164,I76147,I150434);
not I_4309 (I76181,I76164);
nor I_4310 (I75831,I76181,I76116);
nor I_4311 (I76212,I150464,I150455);
or I_4312 (I76229,I76212,I150437);
nor I_4313 (I76246,I150434,I150440);
nand I_4314 (I76263,I76246,I76229);
not I_4315 (I76280,I76263);
nor I_4316 (I76297,I76280,I75924);
or I_4317 (I76314,I76297,I76164);
nor I_4318 (I75813,I75890,I76314);
nor I_4319 (I76345,I76280,I150461);
DFFARX1 I_4320 (I76345,I2898,I75839,I75816,);
nor I_4321 (I76376,I76280,I76164);
nor I_4322 (I75822,I76085,I76376);
nor I_4323 (I76407,I76164,I76263);
nor I_4324 (I75810,I75941,I76407);
not I_4325 (I76468,I2905);
nor I_4326 (I76485,I375818,I375803);
nor I_4327 (I76502,I76485,I375833);
not I_4328 (I76519,I76502);
not I_4329 (I76536,I375830);
nor I_4330 (I76553,I76536,I76485);
not I_4331 (I76570,I76553);
nand I_4332 (I76448,I76519,I76570);
nand I_4333 (I76601,I76502,I375824);
not I_4334 (I76433,I76601);
nor I_4335 (I76457,I76553,I375824);
not I_4336 (I76646,I375821);
nand I_4337 (I76663,I375803,I375806);
nand I_4338 (I76680,I76663,I76646);
nand I_4339 (I76697,I76663,I375821);
not I_4340 (I76714,I76697);
nor I_4341 (I76436,I76714,I76601);
nor I_4342 (I76745,I76714,I375824);
nand I_4343 (I76454,I76519,I76697);
and I_4344 (I76776,I76680,I375806);
nand I_4345 (I76793,I76776,I375809);
not I_4346 (I76810,I76793);
nor I_4347 (I76460,I76810,I76745);
nor I_4348 (I76841,I375836,I375812);
or I_4349 (I76858,I76841,I375809);
nor I_4350 (I76875,I375827,I375815);
nand I_4351 (I76892,I76875,I76858);
not I_4352 (I76909,I76892);
nor I_4353 (I76926,I76909,I76553);
or I_4354 (I76943,I76926,I76793);
nor I_4355 (I76442,I76519,I76943);
nor I_4356 (I76974,I76909,I375824);
DFFARX1 I_4357 (I76974,I2898,I76468,I76445,);
nor I_4358 (I77005,I76909,I76793);
nor I_4359 (I76451,I76714,I77005);
nor I_4360 (I77036,I76793,I76892);
nor I_4361 (I76439,I76570,I77036);
not I_4362 (I77097,I2905);
nor I_4363 (I77114,I380340,I380325);
nor I_4364 (I77131,I77114,I380355);
not I_4365 (I77148,I77131);
not I_4366 (I77165,I380352);
nor I_4367 (I77182,I77165,I77114);
not I_4368 (I77199,I77182);
nand I_4369 (I77077,I77148,I77199);
nand I_4370 (I77230,I77131,I380346);
not I_4371 (I77062,I77230);
nor I_4372 (I77086,I77182,I380346);
not I_4373 (I77275,I380343);
nand I_4374 (I77292,I380325,I380328);
nand I_4375 (I77309,I77292,I77275);
nand I_4376 (I77326,I77292,I380343);
not I_4377 (I77343,I77326);
nor I_4378 (I77065,I77343,I77230);
nor I_4379 (I77374,I77343,I380346);
nand I_4380 (I77083,I77148,I77326);
and I_4381 (I77405,I77309,I380328);
nand I_4382 (I77422,I77405,I380331);
not I_4383 (I77439,I77422);
nor I_4384 (I77089,I77439,I77374);
nor I_4385 (I77470,I380358,I380334);
or I_4386 (I77487,I77470,I380331);
nor I_4387 (I77504,I380349,I380337);
nand I_4388 (I77521,I77504,I77487);
not I_4389 (I77538,I77521);
nor I_4390 (I77555,I77538,I77182);
or I_4391 (I77572,I77555,I77422);
nor I_4392 (I77071,I77148,I77572);
nor I_4393 (I77603,I77538,I380346);
DFFARX1 I_4394 (I77603,I2898,I77097,I77074,);
nor I_4395 (I77634,I77538,I77422);
nor I_4396 (I77080,I77343,I77634);
nor I_4397 (I77665,I77422,I77521);
nor I_4398 (I77068,I77199,I77665);
not I_4399 (I77726,I2905);
nor I_4400 (I77743,I195997,I195997);
nor I_4401 (I77760,I77743,I196015);
not I_4402 (I77777,I77760);
not I_4403 (I77794,I196012);
nor I_4404 (I77811,I77794,I77743);
not I_4405 (I77828,I77811);
nand I_4406 (I77706,I77777,I77828);
nand I_4407 (I77859,I77760,I196018);
not I_4408 (I77691,I77859);
nor I_4409 (I77715,I77811,I196018);
not I_4410 (I77904,I196006);
nand I_4411 (I77921,I195994,I196006);
nand I_4412 (I77938,I77921,I77904);
nand I_4413 (I77955,I77921,I196006);
not I_4414 (I77972,I77955);
nor I_4415 (I77694,I77972,I77859);
nor I_4416 (I78003,I77972,I196018);
nand I_4417 (I77712,I77777,I77955);
and I_4418 (I78034,I77938,I196000);
nand I_4419 (I78051,I78034,I196003);
not I_4420 (I78068,I78051);
nor I_4421 (I77718,I78068,I78003);
nor I_4422 (I78099,I195994,I196000);
or I_4423 (I78116,I78099,I196003);
nor I_4424 (I78133,I196009,I196009);
nand I_4425 (I78150,I78133,I78116);
not I_4426 (I78167,I78150);
nor I_4427 (I78184,I78167,I77811);
or I_4428 (I78201,I78184,I78051);
nor I_4429 (I77700,I77777,I78201);
nor I_4430 (I78232,I78167,I196018);
DFFARX1 I_4431 (I78232,I2898,I77726,I77703,);
nor I_4432 (I78263,I78167,I78051);
nor I_4433 (I77709,I77972,I78263);
nor I_4434 (I78294,I78051,I78150);
nor I_4435 (I77697,I77828,I78294);
not I_4436 (I78355,I2905);
nor I_4437 (I78372,I190421,I190421);
nor I_4438 (I78389,I78372,I190439);
not I_4439 (I78406,I78389);
not I_4440 (I78423,I190436);
nor I_4441 (I78440,I78423,I78372);
not I_4442 (I78457,I78440);
nand I_4443 (I78335,I78406,I78457);
nand I_4444 (I78488,I78389,I190442);
not I_4445 (I78320,I78488);
nor I_4446 (I78344,I78440,I190442);
not I_4447 (I78533,I190430);
nand I_4448 (I78550,I190418,I190430);
nand I_4449 (I78567,I78550,I78533);
nand I_4450 (I78584,I78550,I190430);
not I_4451 (I78601,I78584);
nor I_4452 (I78323,I78601,I78488);
nor I_4453 (I78632,I78601,I190442);
nand I_4454 (I78341,I78406,I78584);
and I_4455 (I78663,I78567,I190424);
nand I_4456 (I78680,I78663,I190427);
not I_4457 (I78697,I78680);
nor I_4458 (I78347,I78697,I78632);
nor I_4459 (I78728,I190418,I190424);
or I_4460 (I78745,I78728,I190427);
nor I_4461 (I78762,I190433,I190433);
nand I_4462 (I78779,I78762,I78745);
not I_4463 (I78796,I78779);
nor I_4464 (I78813,I78796,I78440);
or I_4465 (I78830,I78813,I78680);
nor I_4466 (I78329,I78406,I78830);
nor I_4467 (I78861,I78796,I190442);
DFFARX1 I_4468 (I78861,I2898,I78355,I78332,);
nor I_4469 (I78892,I78796,I78680);
nor I_4470 (I78338,I78601,I78892);
nor I_4471 (I78923,I78680,I78779);
nor I_4472 (I78326,I78457,I78923);
not I_4473 (I78984,I2905);
nor I_4474 (I79001,I51157,I51175);
nor I_4475 (I79018,I79001,I51154);
not I_4476 (I79035,I79018);
not I_4477 (I79052,I51154);
nor I_4478 (I79069,I79052,I79001);
not I_4479 (I79086,I79069);
nand I_4480 (I78964,I79035,I79086);
nand I_4481 (I79117,I79018,I51163);
not I_4482 (I78949,I79117);
nor I_4483 (I78973,I79069,I51163);
not I_4484 (I79162,I51190);
nand I_4485 (I79179,I51169,I51172);
nand I_4486 (I79196,I79179,I79162);
nand I_4487 (I79213,I79179,I51190);
not I_4488 (I79230,I79213);
nor I_4489 (I78952,I79230,I79117);
nor I_4490 (I79261,I79230,I51163);
nand I_4491 (I78970,I79035,I79213);
and I_4492 (I79292,I79196,I51187);
nand I_4493 (I79309,I79292,I51178);
not I_4494 (I79326,I79309);
nor I_4495 (I78976,I79326,I79261);
nor I_4496 (I79357,I51160,I51181);
or I_4497 (I79374,I79357,I51157);
nor I_4498 (I79391,I51166,I51184);
nand I_4499 (I79408,I79391,I79374);
not I_4500 (I79425,I79408);
nor I_4501 (I79442,I79425,I79069);
or I_4502 (I79459,I79442,I79309);
nor I_4503 (I78958,I79035,I79459);
nor I_4504 (I79490,I79425,I51163);
DFFARX1 I_4505 (I79490,I2898,I78984,I78961,);
nor I_4506 (I79521,I79425,I79309);
nor I_4507 (I78967,I79230,I79521);
nor I_4508 (I79552,I79309,I79408);
nor I_4509 (I78955,I79086,I79552);
not I_4510 (I79613,I2905);
nor I_4511 (I79630,I413623,I413626);
nor I_4512 (I79647,I79630,I413644);
not I_4513 (I79664,I79647);
not I_4514 (I79681,I413617);
nor I_4515 (I79698,I79681,I79630);
not I_4516 (I79715,I79698);
nand I_4517 (I79593,I79664,I79715);
nand I_4518 (I79746,I79647,I413614);
not I_4519 (I79578,I79746);
nor I_4520 (I79602,I79698,I413614);
not I_4521 (I79791,I413611);
nand I_4522 (I79808,I413641,I413620);
nand I_4523 (I79825,I79808,I79791);
nand I_4524 (I79842,I79808,I413611);
not I_4525 (I79859,I79842);
nor I_4526 (I79581,I79859,I79746);
nor I_4527 (I79890,I79859,I413614);
nand I_4528 (I79599,I79664,I79842);
and I_4529 (I79921,I79825,I413632);
nand I_4530 (I79938,I79921,I413638);
not I_4531 (I79955,I79938);
nor I_4532 (I79605,I79955,I79890);
nor I_4533 (I79986,I413629,I413617);
or I_4534 (I80003,I79986,I413614);
nor I_4535 (I80020,I413611,I413635);
nand I_4536 (I80037,I80020,I80003);
not I_4537 (I80054,I80037);
nor I_4538 (I80071,I80054,I79698);
or I_4539 (I80088,I80071,I79938);
nor I_4540 (I79587,I79664,I80088);
nor I_4541 (I80119,I80054,I413614);
DFFARX1 I_4542 (I80119,I2898,I79613,I79590,);
nor I_4543 (I80150,I80054,I79938);
nor I_4544 (I79596,I79859,I80150);
nor I_4545 (I80181,I79938,I80037);
nor I_4546 (I79584,I79715,I80181);
not I_4547 (I80242,I2905);
nor I_4548 (I80259,I254358,I254358);
nor I_4549 (I80276,I80259,I254367);
not I_4550 (I80293,I80276);
not I_4551 (I80310,I254355);
nor I_4552 (I80327,I80310,I80259);
not I_4553 (I80344,I80327);
nand I_4554 (I80222,I80293,I80344);
nand I_4555 (I80375,I80276,I254376);
not I_4556 (I80207,I80375);
nor I_4557 (I80231,I80327,I254376);
not I_4558 (I80420,I254382);
nand I_4559 (I80437,I254385,I254373);
nand I_4560 (I80454,I80437,I80420);
nand I_4561 (I80471,I80437,I254382);
not I_4562 (I80488,I80471);
nor I_4563 (I80210,I80488,I80375);
nor I_4564 (I80519,I80488,I254376);
nand I_4565 (I80228,I80293,I80471);
and I_4566 (I80550,I80454,I254379);
nand I_4567 (I80567,I80550,I254355);
not I_4568 (I80584,I80567);
nor I_4569 (I80234,I80584,I80519);
nor I_4570 (I80615,I254361,I254364);
or I_4571 (I80632,I80615,I254364);
nor I_4572 (I80649,I254370,I254361);
nand I_4573 (I80666,I80649,I80632);
not I_4574 (I80683,I80666);
nor I_4575 (I80700,I80683,I80327);
or I_4576 (I80717,I80700,I80567);
nor I_4577 (I80216,I80293,I80717);
nor I_4578 (I80748,I80683,I254376);
DFFARX1 I_4579 (I80748,I2898,I80242,I80219,);
nor I_4580 (I80779,I80683,I80567);
nor I_4581 (I80225,I80488,I80779);
nor I_4582 (I80810,I80567,I80666);
nor I_4583 (I80213,I80344,I80810);
not I_4584 (I80871,I2905);
nor I_4585 (I80888,I220940,I220919);
nor I_4586 (I80905,I80888,I220934);
not I_4587 (I80922,I80905);
not I_4588 (I80939,I220916);
nor I_4589 (I80956,I80939,I80888);
not I_4590 (I80973,I80956);
nand I_4591 (I80851,I80922,I80973);
nand I_4592 (I81004,I80905,I220931);
not I_4593 (I80836,I81004);
nor I_4594 (I80860,I80956,I220931);
not I_4595 (I81049,I220922);
nand I_4596 (I81066,I220928,I220919);
nand I_4597 (I81083,I81066,I81049);
nand I_4598 (I81100,I81066,I220922);
not I_4599 (I81117,I81100);
nor I_4600 (I80839,I81117,I81004);
nor I_4601 (I81148,I81117,I220931);
nand I_4602 (I80857,I80922,I81100);
and I_4603 (I81179,I81083,I220937);
nand I_4604 (I81196,I81179,I220916);
not I_4605 (I81213,I81196);
nor I_4606 (I80863,I81213,I81148);
nor I_4607 (I81244,I220925,I220922);
or I_4608 (I81261,I81244,I220928);
nor I_4609 (I81278,I220925,I220943);
nand I_4610 (I81295,I81278,I81261);
not I_4611 (I81312,I81295);
nor I_4612 (I81329,I81312,I80956);
or I_4613 (I81346,I81329,I81196);
nor I_4614 (I80845,I80922,I81346);
nor I_4615 (I81377,I81312,I220931);
DFFARX1 I_4616 (I81377,I2898,I80871,I80848,);
nor I_4617 (I81408,I81312,I81196);
nor I_4618 (I80854,I81117,I81408);
nor I_4619 (I81439,I81196,I81295);
nor I_4620 (I80842,I80973,I81439);
not I_4621 (I81500,I2905);
nor I_4622 (I81517,I26080,I26074);
nor I_4623 (I81534,I81517,I26062);
not I_4624 (I81551,I81534);
not I_4625 (I81568,I26065);
nor I_4626 (I81585,I81568,I81517);
not I_4627 (I81602,I81585);
nand I_4628 (I81480,I81551,I81602);
nand I_4629 (I81633,I81534,I26068);
not I_4630 (I81465,I81633);
nor I_4631 (I81489,I81585,I26068);
not I_4632 (I81678,I26077);
nand I_4633 (I81695,I26071,I26065);
nand I_4634 (I81712,I81695,I81678);
nand I_4635 (I81729,I81695,I26077);
not I_4636 (I81746,I81729);
nor I_4637 (I81468,I81746,I81633);
nor I_4638 (I81777,I81746,I26068);
nand I_4639 (I81486,I81551,I81729);
and I_4640 (I81808,I81712,I26074);
nand I_4641 (I81825,I81808,I26071);
not I_4642 (I81842,I81825);
nor I_4643 (I81492,I81842,I81777);
nor I_4644 (I81873,I26089,I26062);
or I_4645 (I81890,I81873,I26083);
nor I_4646 (I81907,I26086,I26068);
nand I_4647 (I81924,I81907,I81890);
not I_4648 (I81941,I81924);
nor I_4649 (I81958,I81941,I81585);
or I_4650 (I81975,I81958,I81825);
nor I_4651 (I81474,I81551,I81975);
nor I_4652 (I82006,I81941,I26068);
DFFARX1 I_4653 (I82006,I2898,I81500,I81477,);
nor I_4654 (I82037,I81941,I81825);
nor I_4655 (I81483,I81746,I82037);
nor I_4656 (I82068,I81825,I81924);
nor I_4657 (I81471,I81602,I82068);
not I_4658 (I82129,I2905);
nor I_4659 (I82146,I298116,I298131);
nor I_4660 (I82163,I82146,I298122);
not I_4661 (I82180,I82163);
not I_4662 (I82197,I298128);
nor I_4663 (I82214,I82197,I82146);
not I_4664 (I82231,I82214);
nand I_4665 (I82109,I82180,I82231);
nand I_4666 (I82262,I82163,I298140);
not I_4667 (I82094,I82262);
nor I_4668 (I82118,I82214,I298140);
not I_4669 (I82307,I298137);
nand I_4670 (I82324,I298125,I298116);
nand I_4671 (I82341,I82324,I82307);
nand I_4672 (I82358,I82324,I298137);
not I_4673 (I82375,I82358);
nor I_4674 (I82097,I82375,I82262);
nor I_4675 (I82406,I82375,I298140);
nand I_4676 (I82115,I82180,I82358);
and I_4677 (I82437,I82341,I298113);
nand I_4678 (I82454,I82437,I298143);
not I_4679 (I82471,I82454);
nor I_4680 (I82121,I82471,I82406);
nor I_4681 (I82502,I298113,I298119);
or I_4682 (I82519,I82502,I298134);
nor I_4683 (I82536,I298119,I298122);
nand I_4684 (I82553,I82536,I82519);
not I_4685 (I82570,I82553);
nor I_4686 (I82587,I82570,I82214);
or I_4687 (I82604,I82587,I82454);
nor I_4688 (I82103,I82180,I82604);
nor I_4689 (I82635,I82570,I298140);
DFFARX1 I_4690 (I82635,I2898,I82129,I82106,);
nor I_4691 (I82666,I82570,I82454);
nor I_4692 (I82112,I82375,I82666);
nor I_4693 (I82697,I82454,I82553);
nor I_4694 (I82100,I82231,I82697);
not I_4695 (I82758,I2905);
nor I_4696 (I82775,I53503,I53521);
nor I_4697 (I82792,I82775,I53500);
not I_4698 (I82809,I82792);
not I_4699 (I82826,I53500);
nor I_4700 (I82843,I82826,I82775);
not I_4701 (I82860,I82843);
nand I_4702 (I82738,I82809,I82860);
nand I_4703 (I82891,I82792,I53509);
not I_4704 (I82723,I82891);
nor I_4705 (I82747,I82843,I53509);
not I_4706 (I82936,I53536);
nand I_4707 (I82953,I53515,I53518);
nand I_4708 (I82970,I82953,I82936);
nand I_4709 (I82987,I82953,I53536);
not I_4710 (I83004,I82987);
nor I_4711 (I82726,I83004,I82891);
nor I_4712 (I83035,I83004,I53509);
nand I_4713 (I82744,I82809,I82987);
and I_4714 (I83066,I82970,I53533);
nand I_4715 (I83083,I83066,I53524);
not I_4716 (I83100,I83083);
nor I_4717 (I82750,I83100,I83035);
nor I_4718 (I83131,I53506,I53527);
or I_4719 (I83148,I83131,I53503);
nor I_4720 (I83165,I53512,I53530);
nand I_4721 (I83182,I83165,I83148);
not I_4722 (I83199,I83182);
nor I_4723 (I83216,I83199,I82843);
or I_4724 (I83233,I83216,I83083);
nor I_4725 (I82732,I82809,I83233);
nor I_4726 (I83264,I83199,I53509);
DFFARX1 I_4727 (I83264,I2898,I82758,I82735,);
nor I_4728 (I83295,I83199,I83083);
nor I_4729 (I82741,I83004,I83295);
nor I_4730 (I83326,I83083,I83182);
nor I_4731 (I82729,I82860,I83326);
not I_4732 (I83387,I2905);
nor I_4733 (I83404,I102186,I102183);
nor I_4734 (I83421,I83404,I102171);
not I_4735 (I83438,I83421);
not I_4736 (I83455,I102198);
nor I_4737 (I83472,I83455,I83404);
not I_4738 (I83489,I83472);
nand I_4739 (I83367,I83438,I83489);
nand I_4740 (I83520,I83421,I102189);
not I_4741 (I83352,I83520);
nor I_4742 (I83376,I83472,I102189);
not I_4743 (I83565,I102174);
nand I_4744 (I83582,I102192,I102171);
nand I_4745 (I83599,I83582,I83565);
nand I_4746 (I83616,I83582,I102174);
not I_4747 (I83633,I83616);
nor I_4748 (I83355,I83633,I83520);
nor I_4749 (I83664,I83633,I102189);
nand I_4750 (I83373,I83438,I83616);
and I_4751 (I83695,I83599,I102180);
nand I_4752 (I83712,I83695,I102177);
not I_4753 (I83729,I83712);
nor I_4754 (I83379,I83729,I83664);
nor I_4755 (I83760,I102177,I102204);
or I_4756 (I83777,I83760,I102174);
nor I_4757 (I83794,I102195,I102201);
nand I_4758 (I83811,I83794,I83777);
not I_4759 (I83828,I83811);
nor I_4760 (I83845,I83828,I83472);
or I_4761 (I83862,I83845,I83712);
nor I_4762 (I83361,I83438,I83862);
nor I_4763 (I83893,I83828,I102189);
DFFARX1 I_4764 (I83893,I2898,I83387,I83364,);
nor I_4765 (I83924,I83828,I83712);
nor I_4766 (I83370,I83633,I83924);
nor I_4767 (I83955,I83712,I83811);
nor I_4768 (I83358,I83489,I83955);
not I_4769 (I84016,I2905);
nor I_4770 (I84033,I147732,I147723);
nor I_4771 (I84050,I84033,I147717);
not I_4772 (I84067,I84050);
not I_4773 (I84084,I147729);
nor I_4774 (I84101,I84084,I84033);
not I_4775 (I84118,I84101);
nand I_4776 (I83996,I84067,I84118);
nand I_4777 (I84149,I84050,I147741);
not I_4778 (I83981,I84149);
nor I_4779 (I84005,I84101,I147741);
not I_4780 (I84194,I147738);
nand I_4781 (I84211,I147747,I147720);
nand I_4782 (I84228,I84211,I84194);
nand I_4783 (I84245,I84211,I147738);
not I_4784 (I84262,I84245);
nor I_4785 (I83984,I84262,I84149);
nor I_4786 (I84293,I84262,I147741);
nand I_4787 (I84002,I84067,I84245);
and I_4788 (I84324,I84228,I147726);
nand I_4789 (I84341,I84324,I147714);
not I_4790 (I84358,I84341);
nor I_4791 (I84008,I84358,I84293);
nor I_4792 (I84389,I147744,I147735);
or I_4793 (I84406,I84389,I147717);
nor I_4794 (I84423,I147714,I147720);
nand I_4795 (I84440,I84423,I84406);
not I_4796 (I84457,I84440);
nor I_4797 (I84474,I84457,I84101);
or I_4798 (I84491,I84474,I84341);
nor I_4799 (I83990,I84067,I84491);
nor I_4800 (I84522,I84457,I147741);
DFFARX1 I_4801 (I84522,I2898,I84016,I83993,);
nor I_4802 (I84553,I84457,I84341);
nor I_4803 (I83999,I84262,I84553);
nor I_4804 (I84584,I84341,I84440);
nor I_4805 (I83987,I84118,I84584);
not I_4806 (I84645,I2905);
nor I_4807 (I84662,I406069,I406078);
nor I_4808 (I84679,I84662,I406072);
not I_4809 (I84696,I84679);
not I_4810 (I84713,I406063);
nor I_4811 (I84730,I84713,I84662);
not I_4812 (I84747,I84730);
nand I_4813 (I84625,I84696,I84747);
nand I_4814 (I84778,I84679,I406069);
not I_4815 (I84610,I84778);
nor I_4816 (I84634,I84730,I406069);
not I_4817 (I84823,I406078);
nand I_4818 (I84840,I406063,I406066);
nand I_4819 (I84857,I84840,I84823);
nand I_4820 (I84874,I84840,I406078);
not I_4821 (I84891,I84874);
nor I_4822 (I84613,I84891,I84778);
nor I_4823 (I84922,I84891,I406069);
nand I_4824 (I84631,I84696,I84874);
and I_4825 (I84953,I84857,I406072);
nand I_4826 (I84970,I84953,I406087);
not I_4827 (I84987,I84970);
nor I_4828 (I84637,I84987,I84922);
nor I_4829 (I85018,I406066,I406084);
or I_4830 (I85035,I85018,I406075);
nor I_4831 (I85052,I406075,I406081);
nand I_4832 (I85069,I85052,I85035);
not I_4833 (I85086,I85069);
nor I_4834 (I85103,I85086,I84730);
or I_4835 (I85120,I85103,I84970);
nor I_4836 (I84619,I84696,I85120);
nor I_4837 (I85151,I85086,I406069);
DFFARX1 I_4838 (I85151,I2898,I84645,I84622,);
nor I_4839 (I85182,I85086,I84970);
nor I_4840 (I84628,I84891,I85182);
nor I_4841 (I85213,I84970,I85069);
nor I_4842 (I84616,I84747,I85213);
not I_4843 (I85274,I2905);
nor I_4844 (I85291,I308350,I308365);
nor I_4845 (I85308,I85291,I308356);
not I_4846 (I85325,I85308);
not I_4847 (I85342,I308362);
nor I_4848 (I85359,I85342,I85291);
not I_4849 (I85376,I85359);
nand I_4850 (I85254,I85325,I85376);
nand I_4851 (I85407,I85308,I308374);
not I_4852 (I85239,I85407);
nor I_4853 (I85263,I85359,I308374);
not I_4854 (I85452,I308371);
nand I_4855 (I85469,I308359,I308350);
nand I_4856 (I85486,I85469,I85452);
nand I_4857 (I85503,I85469,I308371);
not I_4858 (I85520,I85503);
nor I_4859 (I85242,I85520,I85407);
nor I_4860 (I85551,I85520,I308374);
nand I_4861 (I85260,I85325,I85503);
and I_4862 (I85582,I85486,I308347);
nand I_4863 (I85599,I85582,I308377);
not I_4864 (I85616,I85599);
nor I_4865 (I85266,I85616,I85551);
nor I_4866 (I85647,I308347,I308353);
or I_4867 (I85664,I85647,I308368);
nor I_4868 (I85681,I308353,I308356);
nand I_4869 (I85698,I85681,I85664);
not I_4870 (I85715,I85698);
nor I_4871 (I85732,I85715,I85359);
or I_4872 (I85749,I85732,I85599);
nor I_4873 (I85248,I85325,I85749);
nor I_4874 (I85780,I85715,I308374);
DFFARX1 I_4875 (I85780,I2898,I85274,I85251,);
nor I_4876 (I85811,I85715,I85599);
nor I_4877 (I85257,I85520,I85811);
nor I_4878 (I85842,I85599,I85698);
nor I_4879 (I85245,I85376,I85842);
not I_4880 (I85903,I2905);
nor I_4881 (I85920,I287151,I287166);
nor I_4882 (I85937,I85920,I287157);
not I_4883 (I85954,I85937);
not I_4884 (I85971,I287163);
nor I_4885 (I85988,I85971,I85920);
not I_4886 (I86005,I85988);
nand I_4887 (I85883,I85954,I86005);
nand I_4888 (I86036,I85937,I287175);
not I_4889 (I85868,I86036);
nor I_4890 (I85892,I85988,I287175);
not I_4891 (I86081,I287172);
nand I_4892 (I86098,I287160,I287151);
nand I_4893 (I86115,I86098,I86081);
nand I_4894 (I86132,I86098,I287172);
not I_4895 (I86149,I86132);
nor I_4896 (I85871,I86149,I86036);
nor I_4897 (I86180,I86149,I287175);
nand I_4898 (I85889,I85954,I86132);
and I_4899 (I86211,I86115,I287148);
nand I_4900 (I86228,I86211,I287178);
not I_4901 (I86245,I86228);
nor I_4902 (I85895,I86245,I86180);
nor I_4903 (I86276,I287148,I287154);
or I_4904 (I86293,I86276,I287169);
nor I_4905 (I86310,I287154,I287157);
nand I_4906 (I86327,I86310,I86293);
not I_4907 (I86344,I86327);
nor I_4908 (I86361,I86344,I85988);
or I_4909 (I86378,I86361,I86228);
nor I_4910 (I85877,I85954,I86378);
nor I_4911 (I86409,I86344,I287175);
DFFARX1 I_4912 (I86409,I2898,I85903,I85880,);
nor I_4913 (I86440,I86344,I86228);
nor I_4914 (I85886,I86149,I86440);
nor I_4915 (I86471,I86228,I86327);
nor I_4916 (I85874,I86005,I86471);
not I_4917 (I86532,I2905);
nor I_4918 (I86549,I243648,I243648);
nor I_4919 (I86566,I86549,I243657);
not I_4920 (I86583,I86566);
not I_4921 (I86600,I243645);
nor I_4922 (I86617,I86600,I86549);
not I_4923 (I86634,I86617);
nand I_4924 (I86512,I86583,I86634);
nand I_4925 (I86665,I86566,I243666);
not I_4926 (I86497,I86665);
nor I_4927 (I86521,I86617,I243666);
not I_4928 (I86710,I243672);
nand I_4929 (I86727,I243675,I243663);
nand I_4930 (I86744,I86727,I86710);
nand I_4931 (I86761,I86727,I243672);
not I_4932 (I86778,I86761);
nor I_4933 (I86500,I86778,I86665);
nor I_4934 (I86809,I86778,I243666);
nand I_4935 (I86518,I86583,I86761);
and I_4936 (I86840,I86744,I243669);
nand I_4937 (I86857,I86840,I243645);
not I_4938 (I86874,I86857);
nor I_4939 (I86524,I86874,I86809);
nor I_4940 (I86905,I243651,I243654);
or I_4941 (I86922,I86905,I243654);
nor I_4942 (I86939,I243660,I243651);
nand I_4943 (I86956,I86939,I86922);
not I_4944 (I86973,I86956);
nor I_4945 (I86990,I86973,I86617);
or I_4946 (I87007,I86990,I86857);
nor I_4947 (I86506,I86583,I87007);
nor I_4948 (I87038,I86973,I243666);
DFFARX1 I_4949 (I87038,I2898,I86532,I86509,);
nor I_4950 (I87069,I86973,I86857);
nor I_4951 (I86515,I86778,I87069);
nor I_4952 (I87100,I86857,I86956);
nor I_4953 (I86503,I86634,I87100);
not I_4954 (I87161,I2905);
nor I_4955 (I87178,I226924,I226903);
nor I_4956 (I87195,I87178,I226918);
not I_4957 (I87212,I87195);
not I_4958 (I87229,I226900);
nor I_4959 (I87246,I87229,I87178);
not I_4960 (I87263,I87246);
nand I_4961 (I87141,I87212,I87263);
nand I_4962 (I87294,I87195,I226915);
not I_4963 (I87126,I87294);
nor I_4964 (I87150,I87246,I226915);
not I_4965 (I87339,I226906);
nand I_4966 (I87356,I226912,I226903);
nand I_4967 (I87373,I87356,I87339);
nand I_4968 (I87390,I87356,I226906);
not I_4969 (I87407,I87390);
nor I_4970 (I87129,I87407,I87294);
nor I_4971 (I87438,I87407,I226915);
nand I_4972 (I87147,I87212,I87390);
and I_4973 (I87469,I87373,I226921);
nand I_4974 (I87486,I87469,I226900);
not I_4975 (I87503,I87486);
nor I_4976 (I87153,I87503,I87438);
nor I_4977 (I87534,I226909,I226906);
or I_4978 (I87551,I87534,I226912);
nor I_4979 (I87568,I226909,I226927);
nand I_4980 (I87585,I87568,I87551);
not I_4981 (I87602,I87585);
nor I_4982 (I87619,I87602,I87246);
or I_4983 (I87636,I87619,I87486);
nor I_4984 (I87135,I87212,I87636);
nor I_4985 (I87667,I87602,I226915);
DFFARX1 I_4986 (I87667,I2898,I87161,I87138,);
nor I_4987 (I87698,I87602,I87486);
nor I_4988 (I87144,I87407,I87698);
nor I_4989 (I87729,I87486,I87585);
nor I_4990 (I87132,I87263,I87729);
not I_4991 (I87790,I2905);
nor I_4992 (I87807,I274248,I274248);
nor I_4993 (I87824,I87807,I274257);
not I_4994 (I87841,I87824);
not I_4995 (I87858,I274245);
nor I_4996 (I87875,I87858,I87807);
not I_4997 (I87892,I87875);
nand I_4998 (I87770,I87841,I87892);
nand I_4999 (I87923,I87824,I274266);
not I_5000 (I87755,I87923);
nor I_5001 (I87779,I87875,I274266);
not I_5002 (I87968,I274272);
nand I_5003 (I87985,I274275,I274263);
nand I_5004 (I88002,I87985,I87968);
nand I_5005 (I88019,I87985,I274272);
not I_5006 (I88036,I88019);
nor I_5007 (I87758,I88036,I87923);
nor I_5008 (I88067,I88036,I274266);
nand I_5009 (I87776,I87841,I88019);
and I_5010 (I88098,I88002,I274269);
nand I_5011 (I88115,I88098,I274245);
not I_5012 (I88132,I88115);
nor I_5013 (I87782,I88132,I88067);
nor I_5014 (I88163,I274251,I274254);
or I_5015 (I88180,I88163,I274254);
nor I_5016 (I88197,I274260,I274251);
nand I_5017 (I88214,I88197,I88180);
not I_5018 (I88231,I88214);
nor I_5019 (I88248,I88231,I87875);
or I_5020 (I88265,I88248,I88115);
nor I_5021 (I87764,I87841,I88265);
nor I_5022 (I88296,I88231,I274266);
DFFARX1 I_5023 (I88296,I2898,I87790,I87767,);
nor I_5024 (I88327,I88231,I88115);
nor I_5025 (I87773,I88036,I88327);
nor I_5026 (I88358,I88115,I88214);
nor I_5027 (I87761,I87892,I88358);
not I_5028 (I88419,I2905);
nor I_5029 (I88436,I332351,I332363);
nor I_5030 (I88453,I88436,I332354);
not I_5031 (I88470,I88453);
not I_5032 (I88487,I332366);
nor I_5033 (I88504,I88487,I88436);
not I_5034 (I88521,I88504);
nand I_5035 (I88399,I88470,I88521);
nand I_5036 (I88552,I88453,I332375);
not I_5037 (I88384,I88552);
nor I_5038 (I88408,I88504,I332375);
not I_5039 (I88597,I332363);
nand I_5040 (I88614,I332357,I332357);
nand I_5041 (I88631,I88614,I88597);
nand I_5042 (I88648,I88614,I332363);
not I_5043 (I88665,I88648);
nor I_5044 (I88387,I88665,I88552);
nor I_5045 (I88696,I88665,I332375);
nand I_5046 (I88405,I88470,I88648);
and I_5047 (I88727,I88631,I332354);
nand I_5048 (I88744,I88727,I332372);
not I_5049 (I88761,I88744);
nor I_5050 (I88411,I88761,I88696);
nor I_5051 (I88792,I332369,I332351);
or I_5052 (I88809,I88792,I332360);
nor I_5053 (I88826,I332360,I332366);
nand I_5054 (I88843,I88826,I88809);
not I_5055 (I88860,I88843);
nor I_5056 (I88877,I88860,I88504);
or I_5057 (I88894,I88877,I88744);
nor I_5058 (I88393,I88470,I88894);
nor I_5059 (I88925,I88860,I332375);
DFFARX1 I_5060 (I88925,I2898,I88419,I88396,);
nor I_5061 (I88956,I88860,I88744);
nor I_5062 (I88402,I88665,I88956);
nor I_5063 (I88987,I88744,I88843);
nor I_5064 (I88390,I88521,I88987);
not I_5065 (I89048,I2905);
nor I_5066 (I89065,I44119,I44137);
nor I_5067 (I89082,I89065,I44116);
not I_5068 (I89099,I89082);
not I_5069 (I89116,I44116);
nor I_5070 (I89133,I89116,I89065);
not I_5071 (I89150,I89133);
nand I_5072 (I89028,I89099,I89150);
nand I_5073 (I89181,I89082,I44125);
not I_5074 (I89013,I89181);
nor I_5075 (I89037,I89133,I44125);
not I_5076 (I89226,I44152);
nand I_5077 (I89243,I44131,I44134);
nand I_5078 (I89260,I89243,I89226);
nand I_5079 (I89277,I89243,I44152);
not I_5080 (I89294,I89277);
nor I_5081 (I89016,I89294,I89181);
nor I_5082 (I89325,I89294,I44125);
nand I_5083 (I89034,I89099,I89277);
and I_5084 (I89356,I89260,I44149);
nand I_5085 (I89373,I89356,I44140);
not I_5086 (I89390,I89373);
nor I_5087 (I89040,I89390,I89325);
nor I_5088 (I89421,I44122,I44143);
or I_5089 (I89438,I89421,I44119);
nor I_5090 (I89455,I44128,I44146);
nand I_5091 (I89472,I89455,I89438);
not I_5092 (I89489,I89472);
nor I_5093 (I89506,I89489,I89133);
or I_5094 (I89523,I89506,I89373);
nor I_5095 (I89022,I89099,I89523);
nor I_5096 (I89554,I89489,I44125);
DFFARX1 I_5097 (I89554,I2898,I89048,I89025,);
nor I_5098 (I89585,I89489,I89373);
nor I_5099 (I89031,I89294,I89585);
nor I_5100 (I89616,I89373,I89472);
nor I_5101 (I89019,I89150,I89616);
not I_5102 (I89677,I2905);
nor I_5103 (I89694,I162012,I162003);
nor I_5104 (I89711,I89694,I161997);
not I_5105 (I89728,I89711);
not I_5106 (I89745,I162009);
nor I_5107 (I89762,I89745,I89694);
not I_5108 (I89779,I89762);
nand I_5109 (I89657,I89728,I89779);
nand I_5110 (I89810,I89711,I162021);
not I_5111 (I89642,I89810);
nor I_5112 (I89666,I89762,I162021);
not I_5113 (I89855,I162018);
nand I_5114 (I89872,I162027,I162000);
nand I_5115 (I89889,I89872,I89855);
nand I_5116 (I89906,I89872,I162018);
not I_5117 (I89923,I89906);
nor I_5118 (I89645,I89923,I89810);
nor I_5119 (I89954,I89923,I162021);
nand I_5120 (I89663,I89728,I89906);
and I_5121 (I89985,I89889,I162006);
nand I_5122 (I90002,I89985,I161994);
not I_5123 (I90019,I90002);
nor I_5124 (I89669,I90019,I89954);
nor I_5125 (I90050,I162024,I162015);
or I_5126 (I90067,I90050,I161997);
nor I_5127 (I90084,I161994,I162000);
nand I_5128 (I90101,I90084,I90067);
not I_5129 (I90118,I90101);
nor I_5130 (I90135,I90118,I89762);
or I_5131 (I90152,I90135,I90002);
nor I_5132 (I89651,I89728,I90152);
nor I_5133 (I90183,I90118,I162021);
DFFARX1 I_5134 (I90183,I2898,I89677,I89654,);
nor I_5135 (I90214,I90118,I90002);
nor I_5136 (I89660,I89923,I90214);
nor I_5137 (I90245,I90002,I90101);
nor I_5138 (I89648,I89779,I90245);
not I_5139 (I90306,I2905);
nor I_5140 (I90323,I2691,I2747);
nor I_5141 (I90340,I90323,I2051);
not I_5142 (I90357,I90340);
not I_5143 (I90374,I2251);
nor I_5144 (I90391,I90374,I90323);
not I_5145 (I90408,I90391);
nand I_5146 (I90286,I90357,I90408);
nand I_5147 (I90439,I90340,I1899);
not I_5148 (I90271,I90439);
nor I_5149 (I90295,I90391,I1899);
not I_5150 (I90484,I2291);
nand I_5151 (I90501,I2203,I2259);
nand I_5152 (I90518,I90501,I90484);
nand I_5153 (I90535,I90501,I2291);
not I_5154 (I90552,I90535);
nor I_5155 (I90274,I90552,I90439);
nor I_5156 (I90583,I90552,I1899);
nand I_5157 (I90292,I90357,I90535);
and I_5158 (I90614,I90518,I2339);
nand I_5159 (I90631,I90614,I1955);
not I_5160 (I90648,I90631);
nor I_5161 (I90298,I90648,I90583);
nor I_5162 (I90679,I2843,I2267);
or I_5163 (I90696,I90679,I2283);
nor I_5164 (I90713,I2059,I2211);
nand I_5165 (I90730,I90713,I90696);
not I_5166 (I90747,I90730);
nor I_5167 (I90764,I90747,I90391);
or I_5168 (I90781,I90764,I90631);
nor I_5169 (I90280,I90357,I90781);
nor I_5170 (I90812,I90747,I1899);
DFFARX1 I_5171 (I90812,I2898,I90306,I90283,);
nor I_5172 (I90843,I90747,I90631);
nor I_5173 (I90289,I90552,I90843);
nor I_5174 (I90874,I90631,I90730);
nor I_5175 (I90277,I90408,I90874);
not I_5176 (I90935,I2905);
nor I_5177 (I90952,I40360,I40354);
nor I_5178 (I90969,I90952,I40342);
not I_5179 (I90986,I90969);
not I_5180 (I91003,I40345);
nor I_5181 (I91020,I91003,I90952);
not I_5182 (I91037,I91020);
nand I_5183 (I90915,I90986,I91037);
nand I_5184 (I91068,I90969,I40348);
not I_5185 (I90900,I91068);
nor I_5186 (I90924,I91020,I40348);
not I_5187 (I91113,I40357);
nand I_5188 (I91130,I40351,I40345);
nand I_5189 (I91147,I91130,I91113);
nand I_5190 (I91164,I91130,I40357);
not I_5191 (I91181,I91164);
nor I_5192 (I90903,I91181,I91068);
nor I_5193 (I91212,I91181,I40348);
nand I_5194 (I90921,I90986,I91164);
and I_5195 (I91243,I91147,I40354);
nand I_5196 (I91260,I91243,I40351);
not I_5197 (I91277,I91260);
nor I_5198 (I90927,I91277,I91212);
nor I_5199 (I91308,I40369,I40342);
or I_5200 (I91325,I91308,I40363);
nor I_5201 (I91342,I40366,I40348);
nand I_5202 (I91359,I91342,I91325);
not I_5203 (I91376,I91359);
nor I_5204 (I91393,I91376,I91020);
or I_5205 (I91410,I91393,I91260);
nor I_5206 (I90909,I90986,I91410);
nor I_5207 (I91441,I91376,I40348);
DFFARX1 I_5208 (I91441,I2898,I90935,I90912,);
nor I_5209 (I91472,I91376,I91260);
nor I_5210 (I90918,I91181,I91472);
nor I_5211 (I91503,I91260,I91359);
nor I_5212 (I90906,I91037,I91503);
not I_5213 (I91564,I2905);
nor I_5214 (I91581,I423381,I423384);
nor I_5215 (I91598,I91581,I423402);
not I_5216 (I91615,I91598);
not I_5217 (I91632,I423375);
nor I_5218 (I91649,I91632,I91581);
not I_5219 (I91666,I91649);
nand I_5220 (I91544,I91615,I91666);
nand I_5221 (I91697,I91598,I423372);
not I_5222 (I91529,I91697);
nor I_5223 (I91553,I91649,I423372);
not I_5224 (I91742,I423369);
nand I_5225 (I91759,I423399,I423378);
nand I_5226 (I91776,I91759,I91742);
nand I_5227 (I91793,I91759,I423369);
not I_5228 (I91810,I91793);
nor I_5229 (I91532,I91810,I91697);
nor I_5230 (I91841,I91810,I423372);
nand I_5231 (I91550,I91615,I91793);
and I_5232 (I91872,I91776,I423390);
nand I_5233 (I91889,I91872,I423396);
not I_5234 (I91906,I91889);
nor I_5235 (I91556,I91906,I91841);
nor I_5236 (I91937,I423387,I423375);
or I_5237 (I91954,I91937,I423372);
nor I_5238 (I91971,I423369,I423393);
nand I_5239 (I91988,I91971,I91954);
not I_5240 (I92005,I91988);
nor I_5241 (I92022,I92005,I91649);
or I_5242 (I92039,I92022,I91889);
nor I_5243 (I91538,I91615,I92039);
nor I_5244 (I92070,I92005,I423372);
DFFARX1 I_5245 (I92070,I2898,I91564,I91541,);
nor I_5246 (I92101,I92005,I91889);
nor I_5247 (I91547,I91810,I92101);
nor I_5248 (I92132,I91889,I91988);
nor I_5249 (I91535,I91666,I92132);
not I_5250 (I92193,I2905);
nor I_5251 (I92210,I210468,I210447);
nor I_5252 (I92227,I92210,I210462);
not I_5253 (I92244,I92227);
not I_5254 (I92261,I210444);
nor I_5255 (I92278,I92261,I92210);
not I_5256 (I92295,I92278);
nand I_5257 (I92173,I92244,I92295);
nand I_5258 (I92326,I92227,I210459);
not I_5259 (I92158,I92326);
nor I_5260 (I92182,I92278,I210459);
not I_5261 (I92371,I210450);
nand I_5262 (I92388,I210456,I210447);
nand I_5263 (I92405,I92388,I92371);
nand I_5264 (I92422,I92388,I210450);
not I_5265 (I92439,I92422);
nor I_5266 (I92161,I92439,I92326);
nor I_5267 (I92470,I92439,I210459);
nand I_5268 (I92179,I92244,I92422);
and I_5269 (I92501,I92405,I210465);
nand I_5270 (I92518,I92501,I210444);
not I_5271 (I92535,I92518);
nor I_5272 (I92185,I92535,I92470);
nor I_5273 (I92566,I210453,I210450);
or I_5274 (I92583,I92566,I210456);
nor I_5275 (I92600,I210453,I210471);
nand I_5276 (I92617,I92600,I92583);
not I_5277 (I92634,I92617);
nor I_5278 (I92651,I92634,I92278);
or I_5279 (I92668,I92651,I92518);
nor I_5280 (I92167,I92244,I92668);
nor I_5281 (I92699,I92634,I210459);
DFFARX1 I_5282 (I92699,I2898,I92193,I92170,);
nor I_5283 (I92730,I92634,I92518);
nor I_5284 (I92176,I92439,I92730);
nor I_5285 (I92761,I92518,I92617);
nor I_5286 (I92164,I92295,I92761);
not I_5287 (I92822,I2905);
nor I_5288 (I92839,I295923,I295938);
nor I_5289 (I92856,I92839,I295929);
not I_5290 (I92873,I92856);
not I_5291 (I92890,I295935);
nor I_5292 (I92907,I92890,I92839);
not I_5293 (I92924,I92907);
nand I_5294 (I92802,I92873,I92924);
nand I_5295 (I92955,I92856,I295947);
not I_5296 (I92787,I92955);
nor I_5297 (I92811,I92907,I295947);
not I_5298 (I93000,I295944);
nand I_5299 (I93017,I295932,I295923);
nand I_5300 (I93034,I93017,I93000);
nand I_5301 (I93051,I93017,I295944);
not I_5302 (I93068,I93051);
nor I_5303 (I92790,I93068,I92955);
nor I_5304 (I93099,I93068,I295947);
nand I_5305 (I92808,I92873,I93051);
and I_5306 (I93130,I93034,I295920);
nand I_5307 (I93147,I93130,I295950);
not I_5308 (I93164,I93147);
nor I_5309 (I92814,I93164,I93099);
nor I_5310 (I93195,I295920,I295926);
or I_5311 (I93212,I93195,I295941);
nor I_5312 (I93229,I295926,I295929);
nand I_5313 (I93246,I93229,I93212);
not I_5314 (I93263,I93246);
nor I_5315 (I93280,I93263,I92907);
or I_5316 (I93297,I93280,I93147);
nor I_5317 (I92796,I92873,I93297);
nor I_5318 (I93328,I93263,I295947);
DFFARX1 I_5319 (I93328,I2898,I92822,I92799,);
nor I_5320 (I93359,I93263,I93147);
nor I_5321 (I92805,I93068,I93359);
nor I_5322 (I93390,I93147,I93246);
nor I_5323 (I92793,I92924,I93390);
not I_5324 (I93451,I2905);
nor I_5325 (I93468,I322236,I322248);
nor I_5326 (I93485,I93468,I322239);
not I_5327 (I93502,I93485);
not I_5328 (I93519,I322251);
nor I_5329 (I93536,I93519,I93468);
not I_5330 (I93553,I93536);
nand I_5331 (I93431,I93502,I93553);
nand I_5332 (I93584,I93485,I322260);
not I_5333 (I93416,I93584);
nor I_5334 (I93440,I93536,I322260);
not I_5335 (I93629,I322248);
nand I_5336 (I93646,I322242,I322242);
nand I_5337 (I93663,I93646,I93629);
nand I_5338 (I93680,I93646,I322248);
not I_5339 (I93697,I93680);
nor I_5340 (I93419,I93697,I93584);
nor I_5341 (I93728,I93697,I322260);
nand I_5342 (I93437,I93502,I93680);
and I_5343 (I93759,I93663,I322239);
nand I_5344 (I93776,I93759,I322257);
not I_5345 (I93793,I93776);
nor I_5346 (I93443,I93793,I93728);
nor I_5347 (I93824,I322254,I322236);
or I_5348 (I93841,I93824,I322245);
nor I_5349 (I93858,I322245,I322251);
nand I_5350 (I93875,I93858,I93841);
not I_5351 (I93892,I93875);
nor I_5352 (I93909,I93892,I93536);
or I_5353 (I93926,I93909,I93776);
nor I_5354 (I93425,I93502,I93926);
nor I_5355 (I93957,I93892,I322260);
DFFARX1 I_5356 (I93957,I2898,I93451,I93428,);
nor I_5357 (I93988,I93892,I93776);
nor I_5358 (I93434,I93697,I93988);
nor I_5359 (I94019,I93776,I93875);
nor I_5360 (I93422,I93553,I94019);
not I_5361 (I94080,I2905);
nor I_5362 (I94097,I411532,I411535);
nor I_5363 (I94114,I94097,I411553);
not I_5364 (I94131,I94114);
not I_5365 (I94148,I411526);
nor I_5366 (I94165,I94148,I94097);
not I_5367 (I94182,I94165);
nand I_5368 (I94060,I94131,I94182);
nand I_5369 (I94213,I94114,I411523);
not I_5370 (I94045,I94213);
nor I_5371 (I94069,I94165,I411523);
not I_5372 (I94258,I411520);
nand I_5373 (I94275,I411550,I411529);
nand I_5374 (I94292,I94275,I94258);
nand I_5375 (I94309,I94275,I411520);
not I_5376 (I94326,I94309);
nor I_5377 (I94048,I94326,I94213);
nor I_5378 (I94357,I94326,I411523);
nand I_5379 (I94066,I94131,I94309);
and I_5380 (I94388,I94292,I411541);
nand I_5381 (I94405,I94388,I411547);
not I_5382 (I94422,I94405);
nor I_5383 (I94072,I94422,I94357);
nor I_5384 (I94453,I411538,I411526);
or I_5385 (I94470,I94453,I411523);
nor I_5386 (I94487,I411520,I411544);
nand I_5387 (I94504,I94487,I94470);
not I_5388 (I94521,I94504);
nor I_5389 (I94538,I94521,I94165);
or I_5390 (I94555,I94538,I94405);
nor I_5391 (I94054,I94131,I94555);
nor I_5392 (I94586,I94521,I411523);
DFFARX1 I_5393 (I94586,I2898,I94080,I94057,);
nor I_5394 (I94617,I94521,I94405);
nor I_5395 (I94063,I94326,I94617);
nor I_5396 (I94648,I94405,I94504);
nor I_5397 (I94051,I94182,I94648);
not I_5398 (I94709,I2905);
nor I_5399 (I94726,I167452,I167443);
nor I_5400 (I94743,I94726,I167437);
not I_5401 (I94760,I94743);
not I_5402 (I94777,I167449);
nor I_5403 (I94794,I94777,I94726);
not I_5404 (I94811,I94794);
nand I_5405 (I94689,I94760,I94811);
nand I_5406 (I94842,I94743,I167461);
not I_5407 (I94674,I94842);
nor I_5408 (I94698,I94794,I167461);
not I_5409 (I94887,I167458);
nand I_5410 (I94904,I167467,I167440);
nand I_5411 (I94921,I94904,I94887);
nand I_5412 (I94938,I94904,I167458);
not I_5413 (I94955,I94938);
nor I_5414 (I94677,I94955,I94842);
nor I_5415 (I94986,I94955,I167461);
nand I_5416 (I94695,I94760,I94938);
and I_5417 (I95017,I94921,I167446);
nand I_5418 (I95034,I95017,I167434);
not I_5419 (I95051,I95034);
nor I_5420 (I94701,I95051,I94986);
nor I_5421 (I95082,I167464,I167455);
or I_5422 (I95099,I95082,I167437);
nor I_5423 (I95116,I167434,I167440);
nand I_5424 (I95133,I95116,I95099);
not I_5425 (I95150,I95133);
nor I_5426 (I95167,I95150,I94794);
or I_5427 (I95184,I95167,I95034);
nor I_5428 (I94683,I94760,I95184);
nor I_5429 (I95215,I95150,I167461);
DFFARX1 I_5430 (I95215,I2898,I94709,I94686,);
nor I_5431 (I95246,I95150,I95034);
nor I_5432 (I94692,I94955,I95246);
nor I_5433 (I95277,I95034,I95133);
nor I_5434 (I94680,I94811,I95277);
not I_5435 (I95338,I2905);
nor I_5436 (I95355,I268893,I268893);
nor I_5437 (I95372,I95355,I268902);
not I_5438 (I95389,I95372);
not I_5439 (I95406,I268890);
nor I_5440 (I95423,I95406,I95355);
not I_5441 (I95440,I95423);
nand I_5442 (I95318,I95389,I95440);
nand I_5443 (I95471,I95372,I268911);
not I_5444 (I95303,I95471);
nor I_5445 (I95327,I95423,I268911);
not I_5446 (I95516,I268917);
nand I_5447 (I95533,I268920,I268908);
nand I_5448 (I95550,I95533,I95516);
nand I_5449 (I95567,I95533,I268917);
not I_5450 (I95584,I95567);
nor I_5451 (I95306,I95584,I95471);
nor I_5452 (I95615,I95584,I268911);
nand I_5453 (I95324,I95389,I95567);
and I_5454 (I95646,I95550,I268914);
nand I_5455 (I95663,I95646,I268890);
not I_5456 (I95680,I95663);
nor I_5457 (I95330,I95680,I95615);
nor I_5458 (I95711,I268896,I268899);
or I_5459 (I95728,I95711,I268899);
nor I_5460 (I95745,I268905,I268896);
nand I_5461 (I95762,I95745,I95728);
not I_5462 (I95779,I95762);
nor I_5463 (I95796,I95779,I95423);
or I_5464 (I95813,I95796,I95663);
nor I_5465 (I95312,I95389,I95813);
nor I_5466 (I95844,I95779,I268911);
DFFARX1 I_5467 (I95844,I2898,I95338,I95315,);
nor I_5468 (I95875,I95779,I95663);
nor I_5469 (I95321,I95584,I95875);
nor I_5470 (I95906,I95663,I95762);
nor I_5471 (I95309,I95440,I95906);
not I_5472 (I95967,I2905);
nor I_5473 (I95984,I147052,I147043);
nor I_5474 (I96001,I95984,I147037);
not I_5475 (I96018,I96001);
not I_5476 (I96035,I147049);
nor I_5477 (I96052,I96035,I95984);
not I_5478 (I96069,I96052);
nand I_5479 (I95947,I96018,I96069);
nand I_5480 (I96100,I96001,I147061);
not I_5481 (I95932,I96100);
nor I_5482 (I95956,I96052,I147061);
not I_5483 (I96145,I147058);
nand I_5484 (I96162,I147067,I147040);
nand I_5485 (I96179,I96162,I96145);
nand I_5486 (I96196,I96162,I147058);
not I_5487 (I96213,I96196);
nor I_5488 (I95935,I96213,I96100);
nor I_5489 (I96244,I96213,I147061);
nand I_5490 (I95953,I96018,I96196);
and I_5491 (I96275,I96179,I147046);
nand I_5492 (I96292,I96275,I147034);
not I_5493 (I96309,I96292);
nor I_5494 (I95959,I96309,I96244);
nor I_5495 (I96340,I147064,I147055);
or I_5496 (I96357,I96340,I147037);
nor I_5497 (I96374,I147034,I147040);
nand I_5498 (I96391,I96374,I96357);
not I_5499 (I96408,I96391);
nor I_5500 (I96425,I96408,I96052);
or I_5501 (I96442,I96425,I96292);
nor I_5502 (I95941,I96018,I96442);
nor I_5503 (I96473,I96408,I147061);
DFFARX1 I_5504 (I96473,I2898,I95967,I95944,);
nor I_5505 (I96504,I96408,I96292);
nor I_5506 (I95950,I96213,I96504);
nor I_5507 (I96535,I96292,I96391);
nor I_5508 (I95938,I96069,I96535);
not I_5509 (I96596,I2905);
nor I_5510 (I96613,I7813,I7819);
nor I_5511 (I96630,I96613,I7831);
not I_5512 (I96647,I96630);
not I_5513 (I96664,I7828);
nor I_5514 (I96681,I96664,I96613);
not I_5515 (I96698,I96681);
nand I_5516 (I96576,I96647,I96698);
nand I_5517 (I96729,I96630,I7834);
not I_5518 (I96561,I96729);
nor I_5519 (I96585,I96681,I7834);
not I_5520 (I96774,I7810);
nand I_5521 (I96791,I7822,I7804);
nand I_5522 (I96808,I96791,I96774);
nand I_5523 (I96825,I96791,I7810);
not I_5524 (I96842,I96825);
nor I_5525 (I96564,I96842,I96729);
nor I_5526 (I96873,I96842,I7834);
nand I_5527 (I96582,I96647,I96825);
and I_5528 (I96904,I96808,I7816);
nand I_5529 (I96921,I96904,I7813);
not I_5530 (I96938,I96921);
nor I_5531 (I96588,I96938,I96873);
nor I_5532 (I96969,I7810,I7807);
or I_5533 (I96986,I96969,I7807);
nor I_5534 (I97003,I7825,I7804);
nand I_5535 (I97020,I97003,I96986);
not I_5536 (I97037,I97020);
nor I_5537 (I97054,I97037,I96681);
or I_5538 (I97071,I97054,I96921);
nor I_5539 (I96570,I96647,I97071);
nor I_5540 (I97102,I97037,I7834);
DFFARX1 I_5541 (I97102,I2898,I96596,I96573,);
nor I_5542 (I97133,I97037,I96921);
nor I_5543 (I96579,I96842,I97133);
nor I_5544 (I97164,I96921,I97020);
nor I_5545 (I96567,I96698,I97164);
not I_5546 (I97225,I2905);
nor I_5547 (I97242,I137410,I137407);
nor I_5548 (I97259,I97242,I137395);
not I_5549 (I97276,I97259);
not I_5550 (I97293,I137422);
nor I_5551 (I97310,I97293,I97242);
not I_5552 (I97327,I97310);
nand I_5553 (I97205,I97276,I97327);
nand I_5554 (I97358,I97259,I137413);
not I_5555 (I97190,I97358);
nor I_5556 (I97214,I97310,I137413);
not I_5557 (I97403,I137398);
nand I_5558 (I97420,I137416,I137395);
nand I_5559 (I97437,I97420,I97403);
nand I_5560 (I97454,I97420,I137398);
not I_5561 (I97471,I97454);
nor I_5562 (I97193,I97471,I97358);
nor I_5563 (I97502,I97471,I137413);
nand I_5564 (I97211,I97276,I97454);
and I_5565 (I97533,I97437,I137404);
nand I_5566 (I97550,I97533,I137401);
not I_5567 (I97567,I97550);
nor I_5568 (I97217,I97567,I97502);
nor I_5569 (I97598,I137401,I137428);
or I_5570 (I97615,I97598,I137398);
nor I_5571 (I97632,I137419,I137425);
nand I_5572 (I97649,I97632,I97615);
not I_5573 (I97666,I97649);
nor I_5574 (I97683,I97666,I97310);
or I_5575 (I97700,I97683,I97550);
nor I_5576 (I97199,I97276,I97700);
nor I_5577 (I97731,I97666,I137413);
DFFARX1 I_5578 (I97731,I2898,I97225,I97202,);
nor I_5579 (I97762,I97666,I97550);
nor I_5580 (I97208,I97471,I97762);
nor I_5581 (I97793,I97550,I97649);
nor I_5582 (I97196,I97327,I97793);
not I_5583 (I97851,I2905);
or I_5584 (I97868,I223184,I223172);
nor I_5585 (I97885,I223184,I223172);
or I_5586 (I97902,I97885,I223163);
nand I_5587 (I97919,I97868,I223187);
not I_5588 (I97936,I97919);
nor I_5589 (I97953,I97936,I223169);
DFFARX1 I_5590 (I97953,I2898,I97851,I97828,);
not I_5591 (I97984,I223169);
nand I_5592 (I97837,I97902,I97984);
not I_5593 (I98015,I223166);
nand I_5594 (I98032,I223169,I223175);
nand I_5595 (I98049,I98015,I98032);
nand I_5596 (I98066,I223166,I223172);
nor I_5597 (I97819,I98066,I223169);
not I_5598 (I98097,I98066);
nand I_5599 (I98114,I98097,I98049);
nor I_5600 (I97843,I98097,I97919);
nor I_5601 (I98145,I223160,I223178);
or I_5602 (I98162,I98145,I223181);
nor I_5603 (I98179,I223160,I223163);
nand I_5604 (I98196,I98179,I98162);
not I_5605 (I98213,I98196);
nand I_5606 (I98230,I97936,I98213);
nand I_5607 (I98247,I98230,I98114);
not I_5608 (I98264,I98247);
nand I_5609 (I98281,I98097,I98247);
nor I_5610 (I97825,I97902,I98281);
nor I_5611 (I97840,I97936,I98213);
nor I_5612 (I98326,I98196,I97919);
nor I_5613 (I97822,I98264,I98326);
nand I_5614 (I98357,I98196,I98049);
nor I_5615 (I98374,I98066,I98357);
nor I_5616 (I97834,I98374,I223169);
nand I_5617 (I98405,I98196,I97902);
not I_5618 (I97831,I98405);
not I_5619 (I98463,I2905);
or I_5620 (I98480,I221688,I221676);
nor I_5621 (I98497,I221688,I221676);
or I_5622 (I98514,I98497,I221667);
nand I_5623 (I98531,I98480,I221691);
not I_5624 (I98548,I98531);
nor I_5625 (I98565,I98548,I221673);
DFFARX1 I_5626 (I98565,I2898,I98463,I98440,);
not I_5627 (I98596,I221673);
nand I_5628 (I98449,I98514,I98596);
not I_5629 (I98627,I221670);
nand I_5630 (I98644,I221673,I221679);
nand I_5631 (I98661,I98627,I98644);
nand I_5632 (I98678,I221670,I221676);
nor I_5633 (I98431,I98678,I221673);
not I_5634 (I98709,I98678);
nand I_5635 (I98726,I98709,I98661);
nor I_5636 (I98455,I98709,I98531);
nor I_5637 (I98757,I221664,I221682);
or I_5638 (I98774,I98757,I221685);
nor I_5639 (I98791,I221664,I221667);
nand I_5640 (I98808,I98791,I98774);
not I_5641 (I98825,I98808);
nand I_5642 (I98842,I98548,I98825);
nand I_5643 (I98859,I98842,I98726);
not I_5644 (I98876,I98859);
nand I_5645 (I98893,I98709,I98859);
nor I_5646 (I98437,I98514,I98893);
nor I_5647 (I98452,I98548,I98825);
nor I_5648 (I98938,I98808,I98531);
nor I_5649 (I98434,I98876,I98938);
nand I_5650 (I98969,I98808,I98661);
nor I_5651 (I98986,I98678,I98969);
nor I_5652 (I98446,I98986,I221673);
nand I_5653 (I99017,I98808,I98514);
not I_5654 (I98443,I99017);
not I_5655 (I99075,I2905);
or I_5656 (I99092,I214956,I214944);
nor I_5657 (I99109,I214956,I214944);
or I_5658 (I99126,I99109,I214935);
nand I_5659 (I99143,I99092,I214959);
not I_5660 (I99160,I99143);
nor I_5661 (I99177,I99160,I214941);
DFFARX1 I_5662 (I99177,I2898,I99075,I99052,);
not I_5663 (I99208,I214941);
nand I_5664 (I99061,I99126,I99208);
not I_5665 (I99239,I214938);
nand I_5666 (I99256,I214941,I214947);
nand I_5667 (I99273,I99239,I99256);
nand I_5668 (I99290,I214938,I214944);
nor I_5669 (I99043,I99290,I214941);
not I_5670 (I99321,I99290);
nand I_5671 (I99338,I99321,I99273);
nor I_5672 (I99067,I99321,I99143);
nor I_5673 (I99369,I214932,I214950);
or I_5674 (I99386,I99369,I214953);
nor I_5675 (I99403,I214932,I214935);
nand I_5676 (I99420,I99403,I99386);
not I_5677 (I99437,I99420);
nand I_5678 (I99454,I99160,I99437);
nand I_5679 (I99471,I99454,I99338);
not I_5680 (I99488,I99471);
nand I_5681 (I99505,I99321,I99471);
nor I_5682 (I99049,I99126,I99505);
nor I_5683 (I99064,I99160,I99437);
nor I_5684 (I99550,I99420,I99143);
nor I_5685 (I99046,I99488,I99550);
nand I_5686 (I99581,I99420,I99273);
nor I_5687 (I99598,I99290,I99581);
nor I_5688 (I99058,I99598,I214941);
nand I_5689 (I99629,I99420,I99126);
not I_5690 (I99055,I99629);
not I_5691 (I99696,I2905);
or I_5692 (I99713,I182757,I182754);
nand I_5693 (I99730,I182766,I182763);
not I_5694 (I99747,I99730);
and I_5695 (I99764,I99747,I99713);
or I_5696 (I99781,I182751,I182760);
nor I_5697 (I99798,I99781,I182760);
not I_5698 (I99815,I99798);
nor I_5699 (I99832,I99730,I99815);
nand I_5700 (I99849,I99798,I99747);
nor I_5701 (I99866,I99798,I99747);
DFFARX1 I_5702 (I99866,I2898,I99696,I99676,);
nor I_5703 (I99897,I182769,I182751);
or I_5704 (I99914,I99897,I182757);
nor I_5705 (I99931,I182754,I182775);
nand I_5706 (I99948,I99931,I99914);
nand I_5707 (I99965,I99948,I99815);
not I_5708 (I99688,I99965);
nand I_5709 (I99996,I182766,I182772);
nor I_5710 (I99655,I99996,I99764);
not I_5711 (I100027,I99996);
nand I_5712 (I100044,I100027,I99764);
not I_5713 (I99661,I100044);
nor I_5714 (I99664,I99798,I100044);
nor I_5715 (I100089,I99747,I100027);
nor I_5716 (I100106,I99996,I182763);
not I_5717 (I100123,I100106);
nor I_5718 (I99670,I100123,I99832);
nand I_5719 (I99658,I100123,I100044);
nand I_5720 (I100168,I100123,I99849);
nand I_5721 (I100185,I100027,I100168);
nor I_5722 (I99673,I99948,I100185);
nand I_5723 (I99685,I99730,I100123);
nand I_5724 (I99682,I100123,I99948);
nor I_5725 (I100244,I100089,I100106);
nor I_5726 (I99667,I99965,I100244);
and I_5727 (I99679,I99948,I99996);
not I_5728 (I100325,I2905);
or I_5729 (I100342,I438730,I438703);
nand I_5730 (I100359,I438733,I438712);
not I_5731 (I100376,I100359);
and I_5732 (I100393,I100376,I100342);
or I_5733 (I100410,I438721,I438706);
nor I_5734 (I100427,I100410,I438724);
not I_5735 (I100444,I100427);
nor I_5736 (I100461,I100359,I100444);
nand I_5737 (I100478,I100427,I100376);
nor I_5738 (I100495,I100427,I100376);
DFFARX1 I_5739 (I100495,I2898,I100325,I100305,);
nor I_5740 (I100526,I438727,I438706);
or I_5741 (I100543,I100526,I438709);
nor I_5742 (I100560,I438715,I438703);
nand I_5743 (I100577,I100560,I100543);
nand I_5744 (I100594,I100577,I100444);
not I_5745 (I100317,I100594);
nand I_5746 (I100625,I438709,I438718);
nor I_5747 (I100284,I100625,I100393);
not I_5748 (I100656,I100625);
nand I_5749 (I100673,I100656,I100393);
not I_5750 (I100290,I100673);
nor I_5751 (I100293,I100427,I100673);
nor I_5752 (I100718,I100376,I100656);
nor I_5753 (I100735,I100625,I438736);
not I_5754 (I100752,I100735);
nor I_5755 (I100299,I100752,I100461);
nand I_5756 (I100287,I100752,I100673);
nand I_5757 (I100797,I100752,I100478);
nand I_5758 (I100814,I100656,I100797);
nor I_5759 (I100302,I100577,I100814);
nand I_5760 (I100314,I100359,I100752);
nand I_5761 (I100311,I100752,I100577);
nor I_5762 (I100873,I100718,I100735);
nor I_5763 (I100296,I100594,I100873);
and I_5764 (I100308,I100577,I100625);
not I_5765 (I100954,I2905);
or I_5766 (I100971,I71404,I71407);
nand I_5767 (I100988,I71416,I71422);
not I_5768 (I101005,I100988);
and I_5769 (I101022,I101005,I100971);
or I_5770 (I101039,I71428,I71413);
nor I_5771 (I101056,I101039,I71425);
not I_5772 (I101073,I101056);
nor I_5773 (I101090,I100988,I101073);
nand I_5774 (I101107,I101056,I101005);
nor I_5775 (I101124,I101056,I101005);
DFFARX1 I_5776 (I101124,I2898,I100954,I100934,);
nor I_5777 (I101155,I71404,I71419);
or I_5778 (I101172,I101155,I71401);
nor I_5779 (I101189,I71413,I71410);
nand I_5780 (I101206,I101189,I101172);
nand I_5781 (I101223,I101206,I101073);
not I_5782 (I100946,I101223);
nand I_5783 (I101254,I71401,I71410);
nor I_5784 (I100913,I101254,I101022);
not I_5785 (I101285,I101254);
nand I_5786 (I101302,I101285,I101022);
not I_5787 (I100919,I101302);
nor I_5788 (I100922,I101056,I101302);
nor I_5789 (I101347,I101005,I101285);
nor I_5790 (I101364,I101254,I71407);
not I_5791 (I101381,I101364);
nor I_5792 (I100928,I101381,I101090);
nand I_5793 (I100916,I101381,I101302);
nand I_5794 (I101426,I101381,I101107);
nand I_5795 (I101443,I101285,I101426);
nor I_5796 (I100931,I101206,I101443);
nand I_5797 (I100943,I100988,I101381);
nand I_5798 (I100940,I101381,I101206);
nor I_5799 (I101502,I101347,I101364);
nor I_5800 (I100925,I101223,I101502);
and I_5801 (I100937,I101206,I101254);
not I_5802 (I101583,I2905);
or I_5803 (I101600,I38923,I38920);
nand I_5804 (I101617,I38914,I38935);
not I_5805 (I101634,I101617);
and I_5806 (I101651,I101634,I101600);
or I_5807 (I101668,I38929,I38941);
nor I_5808 (I101685,I101668,I38923);
not I_5809 (I101702,I101685);
nor I_5810 (I101719,I101617,I101702);
nand I_5811 (I101736,I101685,I101634);
nor I_5812 (I101753,I101685,I101634);
DFFARX1 I_5813 (I101753,I2898,I101583,I101563,);
nor I_5814 (I101784,I38926,I38926);
or I_5815 (I101801,I101784,I38932);
nor I_5816 (I101818,I38917,I38920);
nand I_5817 (I101835,I101818,I101801);
nand I_5818 (I101852,I101835,I101702);
not I_5819 (I101575,I101852);
nand I_5820 (I101883,I38938,I38914);
nor I_5821 (I101542,I101883,I101651);
not I_5822 (I101914,I101883);
nand I_5823 (I101931,I101914,I101651);
not I_5824 (I101548,I101931);
nor I_5825 (I101551,I101685,I101931);
nor I_5826 (I101976,I101634,I101914);
nor I_5827 (I101993,I101883,I38917);
not I_5828 (I102010,I101993);
nor I_5829 (I101557,I102010,I101719);
nand I_5830 (I101545,I102010,I101931);
nand I_5831 (I102055,I102010,I101736);
nand I_5832 (I102072,I101914,I102055);
nor I_5833 (I101560,I101835,I102072);
nand I_5834 (I101572,I101617,I102010);
nand I_5835 (I101569,I102010,I101835);
nor I_5836 (I102131,I101976,I101993);
nor I_5837 (I101554,I101852,I102131);
and I_5838 (I101566,I101835,I101883);
not I_5839 (I102212,I2905);
or I_5840 (I102229,I422002,I421975);
nand I_5841 (I102246,I422005,I421984);
not I_5842 (I102263,I102246);
and I_5843 (I102280,I102263,I102229);
or I_5844 (I102297,I421993,I421978);
nor I_5845 (I102314,I102297,I421996);
not I_5846 (I102331,I102314);
nor I_5847 (I102348,I102246,I102331);
nand I_5848 (I102365,I102314,I102263);
nor I_5849 (I102382,I102314,I102263);
DFFARX1 I_5850 (I102382,I2898,I102212,I102192,);
nor I_5851 (I102413,I421999,I421978);
or I_5852 (I102430,I102413,I421981);
nor I_5853 (I102447,I421987,I421975);
nand I_5854 (I102464,I102447,I102430);
nand I_5855 (I102481,I102464,I102331);
not I_5856 (I102204,I102481);
nand I_5857 (I102512,I421981,I421990);
nor I_5858 (I102171,I102512,I102280);
not I_5859 (I102543,I102512);
nand I_5860 (I102560,I102543,I102280);
not I_5861 (I102177,I102560);
nor I_5862 (I102180,I102314,I102560);
nor I_5863 (I102605,I102263,I102543);
nor I_5864 (I102622,I102512,I422008);
not I_5865 (I102639,I102622);
nor I_5866 (I102186,I102639,I102348);
nand I_5867 (I102174,I102639,I102560);
nand I_5868 (I102684,I102639,I102365);
nand I_5869 (I102701,I102543,I102684);
nor I_5870 (I102189,I102464,I102701);
nand I_5871 (I102201,I102246,I102639);
nand I_5872 (I102198,I102639,I102464);
nor I_5873 (I102760,I102605,I102622);
nor I_5874 (I102183,I102481,I102760);
and I_5875 (I102195,I102464,I102512);
not I_5876 (I102841,I2905);
or I_5877 (I102858,I64485,I64488);
nand I_5878 (I102875,I64497,I64503);
not I_5879 (I102892,I102875);
and I_5880 (I102909,I102892,I102858);
or I_5881 (I102926,I64509,I64494);
nor I_5882 (I102943,I102926,I64506);
not I_5883 (I102960,I102943);
nor I_5884 (I102977,I102875,I102960);
nand I_5885 (I102994,I102943,I102892);
nor I_5886 (I103011,I102943,I102892);
DFFARX1 I_5887 (I103011,I2898,I102841,I102821,);
nor I_5888 (I103042,I64485,I64500);
or I_5889 (I103059,I103042,I64482);
nor I_5890 (I103076,I64494,I64491);
nand I_5891 (I103093,I103076,I103059);
nand I_5892 (I103110,I103093,I102960);
not I_5893 (I102833,I103110);
nand I_5894 (I103141,I64482,I64491);
nor I_5895 (I102800,I103141,I102909);
not I_5896 (I103172,I103141);
nand I_5897 (I103189,I103172,I102909);
not I_5898 (I102806,I103189);
nor I_5899 (I102809,I102943,I103189);
nor I_5900 (I103234,I102892,I103172);
nor I_5901 (I103251,I103141,I64488);
not I_5902 (I103268,I103251);
nor I_5903 (I102815,I103268,I102977);
nand I_5904 (I102803,I103268,I103189);
nand I_5905 (I103313,I103268,I102994);
nand I_5906 (I103330,I103172,I103313);
nor I_5907 (I102818,I103093,I103330);
nand I_5908 (I102830,I102875,I103268);
nand I_5909 (I102827,I103268,I103093);
nor I_5910 (I103389,I103234,I103251);
nor I_5911 (I102812,I103110,I103389);
and I_5912 (I102824,I103093,I103141);
not I_5913 (I103470,I2905);
or I_5914 (I103487,I62598,I62601);
nand I_5915 (I103504,I62610,I62616);
not I_5916 (I103521,I103504);
and I_5917 (I103538,I103521,I103487);
or I_5918 (I103555,I62622,I62607);
nor I_5919 (I103572,I103555,I62619);
not I_5920 (I103589,I103572);
nor I_5921 (I103606,I103504,I103589);
nand I_5922 (I103623,I103572,I103521);
nor I_5923 (I103640,I103572,I103521);
DFFARX1 I_5924 (I103640,I2898,I103470,I103450,);
nor I_5925 (I103671,I62598,I62613);
or I_5926 (I103688,I103671,I62595);
nor I_5927 (I103705,I62607,I62604);
nand I_5928 (I103722,I103705,I103688);
nand I_5929 (I103739,I103722,I103589);
not I_5930 (I103462,I103739);
nand I_5931 (I103770,I62595,I62604);
nor I_5932 (I103429,I103770,I103538);
not I_5933 (I103801,I103770);
nand I_5934 (I103818,I103801,I103538);
not I_5935 (I103435,I103818);
nor I_5936 (I103438,I103572,I103818);
nor I_5937 (I103863,I103521,I103801);
nor I_5938 (I103880,I103770,I62601);
not I_5939 (I103897,I103880);
nor I_5940 (I103444,I103897,I103606);
nand I_5941 (I103432,I103897,I103818);
nand I_5942 (I103942,I103897,I103623);
nand I_5943 (I103959,I103801,I103942);
nor I_5944 (I103447,I103722,I103959);
nand I_5945 (I103459,I103504,I103897);
nand I_5946 (I103456,I103897,I103722);
nor I_5947 (I104018,I103863,I103880);
nor I_5948 (I103441,I103739,I104018);
and I_5949 (I103453,I103722,I103770);
not I_5950 (I104099,I2905);
or I_5951 (I104116,I368112,I368097);
nand I_5952 (I104133,I368100,I368118);
not I_5953 (I104150,I104133);
and I_5954 (I104167,I104150,I104116);
or I_5955 (I104184,I368091,I368085);
nor I_5956 (I104201,I104184,I368088);
not I_5957 (I104218,I104201);
nor I_5958 (I104235,I104133,I104218);
nand I_5959 (I104252,I104201,I104150);
nor I_5960 (I104269,I104201,I104150);
DFFARX1 I_5961 (I104269,I2898,I104099,I104079,);
nor I_5962 (I104300,I368091,I368109);
or I_5963 (I104317,I104300,I368106);
nor I_5964 (I104334,I368115,I368085);
nand I_5965 (I104351,I104334,I104317);
nand I_5966 (I104368,I104351,I104218);
not I_5967 (I104091,I104368);
nand I_5968 (I104399,I368094,I368103);
nor I_5969 (I104058,I104399,I104167);
not I_5970 (I104430,I104399);
nand I_5971 (I104447,I104430,I104167);
not I_5972 (I104064,I104447);
nor I_5973 (I104067,I104201,I104447);
nor I_5974 (I104492,I104150,I104430);
nor I_5975 (I104509,I104399,I368088);
not I_5976 (I104526,I104509);
nor I_5977 (I104073,I104526,I104235);
nand I_5978 (I104061,I104526,I104447);
nand I_5979 (I104571,I104526,I104252);
nand I_5980 (I104588,I104430,I104571);
nor I_5981 (I104076,I104351,I104588);
nand I_5982 (I104088,I104133,I104526);
nand I_5983 (I104085,I104526,I104351);
nor I_5984 (I104647,I104492,I104509);
nor I_5985 (I104070,I104368,I104647);
and I_5986 (I104082,I104351,I104399);
not I_5987 (I104728,I2905);
or I_5988 (I104745,I215686,I215701);
nand I_5989 (I104762,I215695,I215698);
not I_5990 (I104779,I104762);
and I_5991 (I104796,I104779,I104745);
or I_5992 (I104813,I215683,I215692);
nor I_5993 (I104830,I104813,I215683);
not I_5994 (I104847,I104830);
nor I_5995 (I104864,I104762,I104847);
nand I_5996 (I104881,I104830,I104779);
nor I_5997 (I104898,I104830,I104779);
DFFARX1 I_5998 (I104898,I2898,I104728,I104708,);
nor I_5999 (I104929,I215686,I215680);
or I_6000 (I104946,I104929,I215692);
nor I_6001 (I104963,I215689,I215707);
nand I_6002 (I104980,I104963,I104946);
nand I_6003 (I104997,I104980,I104847);
not I_6004 (I104720,I104997);
nand I_6005 (I105028,I215704,I215689);
nor I_6006 (I104687,I105028,I104796);
not I_6007 (I105059,I105028);
nand I_6008 (I105076,I105059,I104796);
not I_6009 (I104693,I105076);
nor I_6010 (I104696,I104830,I105076);
nor I_6011 (I105121,I104779,I105059);
nor I_6012 (I105138,I105028,I215680);
not I_6013 (I105155,I105138);
nor I_6014 (I104702,I105155,I104864);
nand I_6015 (I104690,I105155,I105076);
nand I_6016 (I105200,I105155,I104881);
nand I_6017 (I105217,I105059,I105200);
nor I_6018 (I104705,I104980,I105217);
nand I_6019 (I104717,I104762,I105155);
nand I_6020 (I104714,I105155,I104980);
nor I_6021 (I105276,I105121,I105138);
nor I_6022 (I104699,I104997,I105276);
and I_6023 (I104711,I104980,I105028);
not I_6024 (I105357,I2905);
or I_6025 (I105374,I419214,I419187);
nand I_6026 (I105391,I419217,I419196);
not I_6027 (I105408,I105391);
and I_6028 (I105425,I105408,I105374);
or I_6029 (I105442,I419205,I419190);
nor I_6030 (I105459,I105442,I419208);
not I_6031 (I105476,I105459);
nor I_6032 (I105493,I105391,I105476);
nand I_6033 (I105510,I105459,I105408);
nor I_6034 (I105527,I105459,I105408);
DFFARX1 I_6035 (I105527,I2898,I105357,I105337,);
nor I_6036 (I105558,I419211,I419190);
or I_6037 (I105575,I105558,I419193);
nor I_6038 (I105592,I419199,I419187);
nand I_6039 (I105609,I105592,I105575);
nand I_6040 (I105626,I105609,I105476);
not I_6041 (I105349,I105626);
nand I_6042 (I105657,I419193,I419202);
nor I_6043 (I105316,I105657,I105425);
not I_6044 (I105688,I105657);
nand I_6045 (I105705,I105688,I105425);
not I_6046 (I105322,I105705);
nor I_6047 (I105325,I105459,I105705);
nor I_6048 (I105750,I105408,I105688);
nor I_6049 (I105767,I105657,I419220);
not I_6050 (I105784,I105767);
nor I_6051 (I105331,I105784,I105493);
nand I_6052 (I105319,I105784,I105705);
nand I_6053 (I105829,I105784,I105510);
nand I_6054 (I105846,I105688,I105829);
nor I_6055 (I105334,I105609,I105846);
nand I_6056 (I105346,I105391,I105784);
nand I_6057 (I105343,I105784,I105609);
nor I_6058 (I105905,I105750,I105767);
nor I_6059 (I105328,I105626,I105905);
and I_6060 (I105340,I105609,I105657);
not I_6061 (I105986,I2905);
or I_6062 (I106003,I9040,I9049);
nand I_6063 (I106020,I9058,I9046);
not I_6064 (I106037,I106020);
and I_6065 (I106054,I106037,I106003);
or I_6066 (I106071,I9043,I9031);
nor I_6067 (I106088,I106071,I9028);
not I_6068 (I106105,I106088);
nor I_6069 (I106122,I106020,I106105);
nand I_6070 (I106139,I106088,I106037);
nor I_6071 (I106156,I106088,I106037);
DFFARX1 I_6072 (I106156,I2898,I105986,I105966,);
nor I_6073 (I106187,I9052,I9031);
or I_6074 (I106204,I106187,I9034);
nor I_6075 (I106221,I9028,I9037);
nand I_6076 (I106238,I106221,I106204);
nand I_6077 (I106255,I106238,I106105);
not I_6078 (I105978,I106255);
nand I_6079 (I106286,I9037,I9034);
nor I_6080 (I105945,I106286,I106054);
not I_6081 (I106317,I106286);
nand I_6082 (I106334,I106317,I106054);
not I_6083 (I105951,I106334);
nor I_6084 (I105954,I106088,I106334);
nor I_6085 (I106379,I106037,I106317);
nor I_6086 (I106396,I106286,I9055);
not I_6087 (I106413,I106396);
nor I_6088 (I105960,I106413,I106122);
nand I_6089 (I105948,I106413,I106334);
nand I_6090 (I106458,I106413,I106139);
nand I_6091 (I106475,I106317,I106458);
nor I_6092 (I105963,I106238,I106475);
nand I_6093 (I105975,I106020,I106413);
nand I_6094 (I105972,I106413,I106238);
nor I_6095 (I106534,I106379,I106396);
nor I_6096 (I105957,I106255,I106534);
and I_6097 (I105969,I106238,I106286);
not I_6098 (I106615,I2905);
or I_6099 (I106632,I225410,I225425);
nand I_6100 (I106649,I225419,I225422);
not I_6101 (I106666,I106649);
and I_6102 (I106683,I106666,I106632);
or I_6103 (I106700,I225407,I225416);
nor I_6104 (I106717,I106700,I225407);
not I_6105 (I106734,I106717);
nor I_6106 (I106751,I106649,I106734);
nand I_6107 (I106768,I106717,I106666);
nor I_6108 (I106785,I106717,I106666);
DFFARX1 I_6109 (I106785,I2898,I106615,I106595,);
nor I_6110 (I106816,I225410,I225404);
or I_6111 (I106833,I106816,I225416);
nor I_6112 (I106850,I225413,I225431);
nand I_6113 (I106867,I106850,I106833);
nand I_6114 (I106884,I106867,I106734);
not I_6115 (I106607,I106884);
nand I_6116 (I106915,I225428,I225413);
nor I_6117 (I106574,I106915,I106683);
not I_6118 (I106946,I106915);
nand I_6119 (I106963,I106946,I106683);
not I_6120 (I106580,I106963);
nor I_6121 (I106583,I106717,I106963);
nor I_6122 (I107008,I106666,I106946);
nor I_6123 (I107025,I106915,I225404);
not I_6124 (I107042,I107025);
nor I_6125 (I106589,I107042,I106751);
nand I_6126 (I106577,I107042,I106963);
nand I_6127 (I107087,I107042,I106768);
nand I_6128 (I107104,I106946,I107087);
nor I_6129 (I106592,I106867,I107104);
nand I_6130 (I106604,I106649,I107042);
nand I_6131 (I106601,I107042,I106867);
nor I_6132 (I107163,I107008,I107025);
nor I_6133 (I106586,I106884,I107163);
and I_6134 (I106598,I106867,I106915);
not I_6135 (I107244,I2905);
or I_6136 (I107261,I185545,I185542);
nand I_6137 (I107278,I185554,I185551);
not I_6138 (I107295,I107278);
and I_6139 (I107312,I107295,I107261);
or I_6140 (I107329,I185539,I185548);
nor I_6141 (I107346,I107329,I185548);
not I_6142 (I107363,I107346);
nor I_6143 (I107380,I107278,I107363);
nand I_6144 (I107397,I107346,I107295);
nor I_6145 (I107414,I107346,I107295);
DFFARX1 I_6146 (I107414,I2898,I107244,I107224,);
nor I_6147 (I107445,I185557,I185539);
or I_6148 (I107462,I107445,I185545);
nor I_6149 (I107479,I185542,I185563);
nand I_6150 (I107496,I107479,I107462);
nand I_6151 (I107513,I107496,I107363);
not I_6152 (I107236,I107513);
nand I_6153 (I107544,I185554,I185560);
nor I_6154 (I107203,I107544,I107312);
not I_6155 (I107575,I107544);
nand I_6156 (I107592,I107575,I107312);
not I_6157 (I107209,I107592);
nor I_6158 (I107212,I107346,I107592);
nor I_6159 (I107637,I107295,I107575);
nor I_6160 (I107654,I107544,I185551);
not I_6161 (I107671,I107654);
nor I_6162 (I107218,I107671,I107380);
nand I_6163 (I107206,I107671,I107592);
nand I_6164 (I107716,I107671,I107397);
nand I_6165 (I107733,I107575,I107716);
nor I_6166 (I107221,I107496,I107733);
nand I_6167 (I107233,I107278,I107671);
nand I_6168 (I107230,I107671,I107496);
nor I_6169 (I107792,I107637,I107654);
nor I_6170 (I107215,I107513,I107792);
and I_6171 (I107227,I107496,I107544);
not I_6172 (I107873,I2905);
or I_6173 (I107890,I280368,I280383);
nand I_6174 (I107907,I280389,I280371);
not I_6175 (I107924,I107907);
and I_6176 (I107941,I107924,I107890);
or I_6177 (I107958,I280374,I280386);
nor I_6178 (I107975,I107958,I280368);
not I_6179 (I107992,I107975);
nor I_6180 (I108009,I107907,I107992);
nand I_6181 (I108026,I107975,I107924);
nor I_6182 (I108043,I107975,I107924);
DFFARX1 I_6183 (I108043,I2898,I107873,I107853,);
nor I_6184 (I108074,I280377,I280365);
or I_6185 (I108091,I108074,I280365);
nor I_6186 (I108108,I280392,I280395);
nand I_6187 (I108125,I108108,I108091);
nand I_6188 (I108142,I108125,I107992);
not I_6189 (I107865,I108142);
nand I_6190 (I108173,I280380,I280371);
nor I_6191 (I107832,I108173,I107941);
not I_6192 (I108204,I108173);
nand I_6193 (I108221,I108204,I107941);
not I_6194 (I107838,I108221);
nor I_6195 (I107841,I107975,I108221);
nor I_6196 (I108266,I107924,I108204);
nor I_6197 (I108283,I108173,I280374);
not I_6198 (I108300,I108283);
nor I_6199 (I107847,I108300,I108009);
nand I_6200 (I107835,I108300,I108221);
nand I_6201 (I108345,I108300,I108026);
nand I_6202 (I108362,I108204,I108345);
nor I_6203 (I107850,I108125,I108362);
nand I_6204 (I107862,I107907,I108300);
nand I_6205 (I107859,I108300,I108125);
nor I_6206 (I108421,I108266,I108283);
nor I_6207 (I107844,I108142,I108421);
and I_6208 (I107856,I108125,I108173);
not I_6209 (I108502,I2905);
or I_6210 (I108519,I75178,I75181);
nand I_6211 (I108536,I75190,I75196);
not I_6212 (I108553,I108536);
and I_6213 (I108570,I108553,I108519);
or I_6214 (I108587,I75202,I75187);
nor I_6215 (I108604,I108587,I75199);
not I_6216 (I108621,I108604);
nor I_6217 (I108638,I108536,I108621);
nand I_6218 (I108655,I108604,I108553);
nor I_6219 (I108672,I108604,I108553);
DFFARX1 I_6220 (I108672,I2898,I108502,I108482,);
nor I_6221 (I108703,I75178,I75193);
or I_6222 (I108720,I108703,I75175);
nor I_6223 (I108737,I75187,I75184);
nand I_6224 (I108754,I108737,I108720);
nand I_6225 (I108771,I108754,I108621);
not I_6226 (I108494,I108771);
nand I_6227 (I108802,I75175,I75184);
nor I_6228 (I108461,I108802,I108570);
not I_6229 (I108833,I108802);
nand I_6230 (I108850,I108833,I108570);
not I_6231 (I108467,I108850);
nor I_6232 (I108470,I108604,I108850);
nor I_6233 (I108895,I108553,I108833);
nor I_6234 (I108912,I108802,I75181);
not I_6235 (I108929,I108912);
nor I_6236 (I108476,I108929,I108638);
nand I_6237 (I108464,I108929,I108850);
nand I_6238 (I108974,I108929,I108655);
nand I_6239 (I108991,I108833,I108974);
nor I_6240 (I108479,I108754,I108991);
nand I_6241 (I108491,I108536,I108929);
nand I_6242 (I108488,I108929,I108754);
nor I_6243 (I109050,I108895,I108912);
nor I_6244 (I108473,I108771,I109050);
and I_6245 (I108485,I108754,I108802);
not I_6246 (I109131,I2905);
or I_6247 (I109148,I417820,I417793);
nand I_6248 (I109165,I417823,I417802);
not I_6249 (I109182,I109165);
and I_6250 (I109199,I109182,I109148);
or I_6251 (I109216,I417811,I417796);
nor I_6252 (I109233,I109216,I417814);
not I_6253 (I109250,I109233);
nor I_6254 (I109267,I109165,I109250);
nand I_6255 (I109284,I109233,I109182);
nor I_6256 (I109301,I109233,I109182);
DFFARX1 I_6257 (I109301,I2898,I109131,I109111,);
nor I_6258 (I109332,I417817,I417796);
or I_6259 (I109349,I109332,I417799);
nor I_6260 (I109366,I417805,I417793);
nand I_6261 (I109383,I109366,I109349);
nand I_6262 (I109400,I109383,I109250);
not I_6263 (I109123,I109400);
nand I_6264 (I109431,I417799,I417808);
nor I_6265 (I109090,I109431,I109199);
not I_6266 (I109462,I109431);
nand I_6267 (I109479,I109462,I109199);
not I_6268 (I109096,I109479);
nor I_6269 (I109099,I109233,I109479);
nor I_6270 (I109524,I109182,I109462);
nor I_6271 (I109541,I109431,I417826);
not I_6272 (I109558,I109541);
nor I_6273 (I109105,I109558,I109267);
nand I_6274 (I109093,I109558,I109479);
nand I_6275 (I109603,I109558,I109284);
nand I_6276 (I109620,I109462,I109603);
nor I_6277 (I109108,I109383,I109620);
nand I_6278 (I109120,I109165,I109558);
nand I_6279 (I109117,I109558,I109383);
nor I_6280 (I109679,I109524,I109541);
nor I_6281 (I109102,I109400,I109679);
and I_6282 (I109114,I109383,I109431);
not I_6283 (I109760,I2905);
or I_6284 (I109777,I63227,I63230);
nand I_6285 (I109794,I63239,I63245);
not I_6286 (I109811,I109794);
and I_6287 (I109828,I109811,I109777);
or I_6288 (I109845,I63251,I63236);
nor I_6289 (I109862,I109845,I63248);
not I_6290 (I109879,I109862);
nor I_6291 (I109896,I109794,I109879);
nand I_6292 (I109913,I109862,I109811);
nor I_6293 (I109930,I109862,I109811);
DFFARX1 I_6294 (I109930,I2898,I109760,I109740,);
nor I_6295 (I109961,I63227,I63242);
or I_6296 (I109978,I109961,I63224);
nor I_6297 (I109995,I63236,I63233);
nand I_6298 (I110012,I109995,I109978);
nand I_6299 (I110029,I110012,I109879);
not I_6300 (I109752,I110029);
nand I_6301 (I110060,I63224,I63233);
nor I_6302 (I109719,I110060,I109828);
not I_6303 (I110091,I110060);
nand I_6304 (I110108,I110091,I109828);
not I_6305 (I109725,I110108);
nor I_6306 (I109728,I109862,I110108);
nor I_6307 (I110153,I109811,I110091);
nor I_6308 (I110170,I110060,I63230);
not I_6309 (I110187,I110170);
nor I_6310 (I109734,I110187,I109896);
nand I_6311 (I109722,I110187,I110108);
nand I_6312 (I110232,I110187,I109913);
nand I_6313 (I110249,I110091,I110232);
nor I_6314 (I109737,I110012,I110249);
nand I_6315 (I109749,I109794,I110187);
nand I_6316 (I109746,I110187,I110012);
nor I_6317 (I110308,I110153,I110170);
nor I_6318 (I109731,I110029,I110308);
and I_6319 (I109743,I110012,I110060);
not I_6320 (I110389,I2905);
or I_6321 (I110406,I397909,I397918);
nand I_6322 (I110423,I397912,I397927);
not I_6323 (I110440,I110423);
and I_6324 (I110457,I110440,I110406);
or I_6325 (I110474,I397924,I397909);
nor I_6326 (I110491,I110474,I397903);
not I_6327 (I110508,I110491);
nor I_6328 (I110525,I110423,I110508);
nand I_6329 (I110542,I110491,I110440);
nor I_6330 (I110559,I110491,I110440);
DFFARX1 I_6331 (I110559,I2898,I110389,I110369,);
nor I_6332 (I110590,I397906,I397918);
or I_6333 (I110607,I110590,I397903);
nor I_6334 (I110624,I397915,I397906);
nand I_6335 (I110641,I110624,I110607);
nand I_6336 (I110658,I110641,I110508);
not I_6337 (I110381,I110658);
nand I_6338 (I110689,I397912,I397921);
nor I_6339 (I110348,I110689,I110457);
not I_6340 (I110720,I110689);
nand I_6341 (I110737,I110720,I110457);
not I_6342 (I110354,I110737);
nor I_6343 (I110357,I110491,I110737);
nor I_6344 (I110782,I110440,I110720);
nor I_6345 (I110799,I110689,I397915);
not I_6346 (I110816,I110799);
nor I_6347 (I110363,I110816,I110525);
nand I_6348 (I110351,I110816,I110737);
nand I_6349 (I110861,I110816,I110542);
nand I_6350 (I110878,I110720,I110861);
nor I_6351 (I110366,I110641,I110878);
nand I_6352 (I110378,I110423,I110816);
nand I_6353 (I110375,I110816,I110641);
nor I_6354 (I110937,I110782,I110799);
nor I_6355 (I110360,I110658,I110937);
and I_6356 (I110372,I110641,I110689);
not I_6357 (I111018,I2905);
or I_6358 (I111035,I2619,I1859);
nand I_6359 (I111052,I1587,I2499);
not I_6360 (I111069,I111052);
and I_6361 (I111086,I111069,I111035);
or I_6362 (I111103,I2099,I2459);
nor I_6363 (I111120,I111103,I2091);
not I_6364 (I111137,I111120);
nor I_6365 (I111154,I111052,I111137);
nand I_6366 (I111171,I111120,I111069);
nor I_6367 (I111188,I111120,I111069);
DFFARX1 I_6368 (I111188,I2898,I111018,I110998,);
nor I_6369 (I111219,I2867,I2507);
or I_6370 (I111236,I111219,I2123);
nor I_6371 (I111253,I2475,I1635);
nand I_6372 (I111270,I111253,I111236);
nand I_6373 (I111287,I111270,I111137);
not I_6374 (I111010,I111287);
nand I_6375 (I111318,I2299,I1995);
nor I_6376 (I110977,I111318,I111086);
not I_6377 (I111349,I111318);
nand I_6378 (I111366,I111349,I111086);
not I_6379 (I110983,I111366);
nor I_6380 (I110986,I111120,I111366);
nor I_6381 (I111411,I111069,I111349);
nor I_6382 (I111428,I111318,I1851);
not I_6383 (I111445,I111428);
nor I_6384 (I110992,I111445,I111154);
nand I_6385 (I110980,I111445,I111366);
nand I_6386 (I111490,I111445,I111171);
nand I_6387 (I111507,I111349,I111490);
nor I_6388 (I110995,I111270,I111507);
nand I_6389 (I111007,I111052,I111445);
nand I_6390 (I111004,I111445,I111270);
nor I_6391 (I111566,I111411,I111428);
nor I_6392 (I110989,I111287,I111566);
and I_6393 (I111001,I111270,I111318);
not I_6394 (I111647,I2905);
or I_6395 (I111664,I4144,I4153);
nand I_6396 (I111681,I4162,I4150);
not I_6397 (I111698,I111681);
and I_6398 (I111715,I111698,I111664);
or I_6399 (I111732,I4147,I4135);
nor I_6400 (I111749,I111732,I4132);
not I_6401 (I111766,I111749);
nor I_6402 (I111783,I111681,I111766);
nand I_6403 (I111800,I111749,I111698);
nor I_6404 (I111817,I111749,I111698);
DFFARX1 I_6405 (I111817,I2898,I111647,I111627,);
nor I_6406 (I111848,I4156,I4135);
or I_6407 (I111865,I111848,I4138);
nor I_6408 (I111882,I4132,I4141);
nand I_6409 (I111899,I111882,I111865);
nand I_6410 (I111916,I111899,I111766);
not I_6411 (I111639,I111916);
nand I_6412 (I111947,I4141,I4138);
nor I_6413 (I111606,I111947,I111715);
not I_6414 (I111978,I111947);
nand I_6415 (I111995,I111978,I111715);
not I_6416 (I111612,I111995);
nor I_6417 (I111615,I111749,I111995);
nor I_6418 (I112040,I111698,I111978);
nor I_6419 (I112057,I111947,I4159);
not I_6420 (I112074,I112057);
nor I_6421 (I111621,I112074,I111783);
nand I_6422 (I111609,I112074,I111995);
nand I_6423 (I112119,I112074,I111800);
nand I_6424 (I112136,I111978,I112119);
nor I_6425 (I111624,I111899,I112136);
nand I_6426 (I111636,I111681,I112074);
nand I_6427 (I111633,I112074,I111899);
nor I_6428 (I112195,I112040,I112057);
nor I_6429 (I111618,I111916,I112195);
and I_6430 (I111630,I111899,I111947);
not I_6431 (I112276,I2905);
or I_6432 (I112293,I7204,I7213);
nand I_6433 (I112310,I7222,I7210);
not I_6434 (I112327,I112310);
and I_6435 (I112344,I112327,I112293);
or I_6436 (I112361,I7207,I7195);
nor I_6437 (I112378,I112361,I7192);
not I_6438 (I112395,I112378);
nor I_6439 (I112412,I112310,I112395);
nand I_6440 (I112429,I112378,I112327);
nor I_6441 (I112446,I112378,I112327);
DFFARX1 I_6442 (I112446,I2898,I112276,I112256,);
nor I_6443 (I112477,I7216,I7195);
or I_6444 (I112494,I112477,I7198);
nor I_6445 (I112511,I7192,I7201);
nand I_6446 (I112528,I112511,I112494);
nand I_6447 (I112545,I112528,I112395);
not I_6448 (I112268,I112545);
nand I_6449 (I112576,I7201,I7198);
nor I_6450 (I112235,I112576,I112344);
not I_6451 (I112607,I112576);
nand I_6452 (I112624,I112607,I112344);
not I_6453 (I112241,I112624);
nor I_6454 (I112244,I112378,I112624);
nor I_6455 (I112669,I112327,I112607);
nor I_6456 (I112686,I112576,I7219);
not I_6457 (I112703,I112686);
nor I_6458 (I112250,I112703,I112412);
nand I_6459 (I112238,I112703,I112624);
nand I_6460 (I112748,I112703,I112429);
nand I_6461 (I112765,I112607,I112748);
nor I_6462 (I112253,I112528,I112765);
nand I_6463 (I112265,I112310,I112703);
nand I_6464 (I112262,I112703,I112528);
nor I_6465 (I112824,I112669,I112686);
nor I_6466 (I112247,I112545,I112824);
and I_6467 (I112259,I112528,I112576);
not I_6468 (I112905,I2905);
or I_6469 (I112922,I405389,I405398);
nand I_6470 (I112939,I405392,I405407);
not I_6471 (I112956,I112939);
and I_6472 (I112973,I112956,I112922);
or I_6473 (I112990,I405404,I405389);
nor I_6474 (I113007,I112990,I405383);
not I_6475 (I113024,I113007);
nor I_6476 (I113041,I112939,I113024);
nand I_6477 (I113058,I113007,I112956);
nor I_6478 (I113075,I113007,I112956);
DFFARX1 I_6479 (I113075,I2898,I112905,I112885,);
nor I_6480 (I113106,I405386,I405398);
or I_6481 (I113123,I113106,I405383);
nor I_6482 (I113140,I405395,I405386);
nand I_6483 (I113157,I113140,I113123);
nand I_6484 (I113174,I113157,I113024);
not I_6485 (I112897,I113174);
nand I_6486 (I113205,I405392,I405401);
nor I_6487 (I112864,I113205,I112973);
not I_6488 (I113236,I113205);
nand I_6489 (I113253,I113236,I112973);
not I_6490 (I112870,I113253);
nor I_6491 (I112873,I113007,I113253);
nor I_6492 (I113298,I112956,I113236);
nor I_6493 (I113315,I113205,I405395);
not I_6494 (I113332,I113315);
nor I_6495 (I112879,I113332,I113041);
nand I_6496 (I112867,I113332,I113253);
nand I_6497 (I113377,I113332,I113058);
nand I_6498 (I113394,I113236,I113377);
nor I_6499 (I112882,I113157,I113394);
nand I_6500 (I112894,I112939,I113332);
nand I_6501 (I112891,I113332,I113157);
nor I_6502 (I113453,I113298,I113315);
nor I_6503 (I112876,I113174,I113453);
and I_6504 (I112888,I113157,I113205);
not I_6505 (I113534,I2905);
or I_6506 (I113551,I276543,I276558);
nand I_6507 (I113568,I276564,I276546);
not I_6508 (I113585,I113568);
and I_6509 (I113602,I113585,I113551);
or I_6510 (I113619,I276549,I276561);
nor I_6511 (I113636,I113619,I276543);
not I_6512 (I113653,I113636);
nor I_6513 (I113670,I113568,I113653);
nand I_6514 (I113687,I113636,I113585);
nor I_6515 (I113704,I113636,I113585);
DFFARX1 I_6516 (I113704,I2898,I113534,I113514,);
nor I_6517 (I113735,I276552,I276540);
or I_6518 (I113752,I113735,I276540);
nor I_6519 (I113769,I276567,I276570);
nand I_6520 (I113786,I113769,I113752);
nand I_6521 (I113803,I113786,I113653);
not I_6522 (I113526,I113803);
nand I_6523 (I113834,I276555,I276546);
nor I_6524 (I113493,I113834,I113602);
not I_6525 (I113865,I113834);
nand I_6526 (I113882,I113865,I113602);
not I_6527 (I113499,I113882);
nor I_6528 (I113502,I113636,I113882);
nor I_6529 (I113927,I113585,I113865);
nor I_6530 (I113944,I113834,I276549);
not I_6531 (I113961,I113944);
nor I_6532 (I113508,I113961,I113670);
nand I_6533 (I113496,I113961,I113882);
nand I_6534 (I114006,I113961,I113687);
nand I_6535 (I114023,I113865,I114006);
nor I_6536 (I113511,I113786,I114023);
nand I_6537 (I113523,I113568,I113961);
nand I_6538 (I113520,I113961,I113786);
nor I_6539 (I114082,I113927,I113944);
nor I_6540 (I113505,I113803,I114082);
and I_6541 (I113517,I113786,I113834);
not I_6542 (I114163,I2905);
or I_6543 (I114180,I186939,I186936);
nand I_6544 (I114197,I186948,I186945);
not I_6545 (I114214,I114197);
and I_6546 (I114231,I114214,I114180);
or I_6547 (I114248,I186933,I186942);
nor I_6548 (I114265,I114248,I186942);
not I_6549 (I114282,I114265);
nor I_6550 (I114299,I114197,I114282);
nand I_6551 (I114316,I114265,I114214);
nor I_6552 (I114333,I114265,I114214);
DFFARX1 I_6553 (I114333,I2898,I114163,I114143,);
nor I_6554 (I114364,I186951,I186933);
or I_6555 (I114381,I114364,I186939);
nor I_6556 (I114398,I186936,I186957);
nand I_6557 (I114415,I114398,I114381);
nand I_6558 (I114432,I114415,I114282);
not I_6559 (I114155,I114432);
nand I_6560 (I114463,I186948,I186954);
nor I_6561 (I114122,I114463,I114231);
not I_6562 (I114494,I114463);
nand I_6563 (I114511,I114494,I114231);
not I_6564 (I114128,I114511);
nor I_6565 (I114131,I114265,I114511);
nor I_6566 (I114556,I114214,I114494);
nor I_6567 (I114573,I114463,I186945);
not I_6568 (I114590,I114573);
nor I_6569 (I114137,I114590,I114299);
nand I_6570 (I114125,I114590,I114511);
nand I_6571 (I114635,I114590,I114316);
nand I_6572 (I114652,I114494,I114635);
nor I_6573 (I114140,I114415,I114652);
nand I_6574 (I114152,I114197,I114590);
nand I_6575 (I114149,I114590,I114415);
nor I_6576 (I114711,I114556,I114573);
nor I_6577 (I114134,I114432,I114711);
and I_6578 (I114146,I114415,I114463);
not I_6579 (I114792,I2905);
or I_6580 (I114809,I1811,I2227);
nand I_6581 (I114826,I1875,I2611);
not I_6582 (I114843,I114826);
and I_6583 (I114860,I114843,I114809);
or I_6584 (I114877,I2115,I1803);
nor I_6585 (I114894,I114877,I2163);
not I_6586 (I114911,I114894);
nor I_6587 (I114928,I114826,I114911);
nand I_6588 (I114945,I114894,I114843);
nor I_6589 (I114962,I114894,I114843);
DFFARX1 I_6590 (I114962,I2898,I114792,I114772,);
nor I_6591 (I114993,I2699,I1659);
or I_6592 (I115010,I114993,I1731);
nor I_6593 (I115027,I2491,I2371);
nand I_6594 (I115044,I115027,I115010);
nand I_6595 (I115061,I115044,I114911);
not I_6596 (I114784,I115061);
nand I_6597 (I115092,I1715,I2219);
nor I_6598 (I114751,I115092,I114860);
not I_6599 (I115123,I115092);
nand I_6600 (I115140,I115123,I114860);
not I_6601 (I114757,I115140);
nor I_6602 (I114760,I114894,I115140);
nor I_6603 (I115185,I114843,I115123);
nor I_6604 (I115202,I115092,I2531);
not I_6605 (I115219,I115202);
nor I_6606 (I114766,I115219,I114928);
nand I_6607 (I114754,I115219,I115140);
nand I_6608 (I115264,I115219,I114945);
nand I_6609 (I115281,I115123,I115264);
nor I_6610 (I114769,I115044,I115281);
nand I_6611 (I114781,I114826,I115219);
nand I_6612 (I114778,I115219,I115044);
nor I_6613 (I115340,I115185,I115202);
nor I_6614 (I114763,I115061,I115340);
and I_6615 (I114775,I115044,I115092);
not I_6616 (I115421,I2905);
or I_6617 (I115438,I170843,I170861);
nand I_6618 (I115455,I170864,I170858);
not I_6619 (I115472,I115455);
and I_6620 (I115489,I115472,I115438);
or I_6621 (I115506,I170852,I170834);
nor I_6622 (I115523,I115506,I170840);
not I_6623 (I115540,I115523);
nor I_6624 (I115557,I115455,I115540);
nand I_6625 (I115574,I115523,I115472);
nor I_6626 (I115591,I115523,I115472);
DFFARX1 I_6627 (I115591,I2898,I115421,I115401,);
nor I_6628 (I115622,I170846,I170867);
or I_6629 (I115639,I115622,I170837);
nor I_6630 (I115656,I170849,I170840);
nand I_6631 (I115673,I115656,I115639);
nand I_6632 (I115690,I115673,I115540);
not I_6633 (I115413,I115690);
nand I_6634 (I115721,I170855,I170837);
nor I_6635 (I115380,I115721,I115489);
not I_6636 (I115752,I115721);
nand I_6637 (I115769,I115752,I115489);
not I_6638 (I115386,I115769);
nor I_6639 (I115389,I115523,I115769);
nor I_6640 (I115814,I115472,I115752);
nor I_6641 (I115831,I115721,I170834);
not I_6642 (I115848,I115831);
nor I_6643 (I115395,I115848,I115557);
nand I_6644 (I115383,I115848,I115769);
nand I_6645 (I115893,I115848,I115574);
nand I_6646 (I115910,I115752,I115893);
nor I_6647 (I115398,I115673,I115910);
nand I_6648 (I115410,I115455,I115848);
nand I_6649 (I115407,I115848,I115673);
nor I_6650 (I115969,I115814,I115831);
nor I_6651 (I115392,I115690,I115969);
and I_6652 (I115404,I115673,I115721);
not I_6653 (I116050,I2905);
or I_6654 (I116067,I173563,I173581);
nand I_6655 (I116084,I173584,I173578);
not I_6656 (I116101,I116084);
and I_6657 (I116118,I116101,I116067);
or I_6658 (I116135,I173572,I173554);
nor I_6659 (I116152,I116135,I173560);
not I_6660 (I116169,I116152);
nor I_6661 (I116186,I116084,I116169);
nand I_6662 (I116203,I116152,I116101);
nor I_6663 (I116220,I116152,I116101);
DFFARX1 I_6664 (I116220,I2898,I116050,I116030,);
nor I_6665 (I116251,I173566,I173587);
or I_6666 (I116268,I116251,I173557);
nor I_6667 (I116285,I173569,I173560);
nand I_6668 (I116302,I116285,I116268);
nand I_6669 (I116319,I116302,I116169);
not I_6670 (I116042,I116319);
nand I_6671 (I116350,I173575,I173557);
nor I_6672 (I116009,I116350,I116118);
not I_6673 (I116381,I116350);
nand I_6674 (I116398,I116381,I116118);
not I_6675 (I116015,I116398);
nor I_6676 (I116018,I116152,I116398);
nor I_6677 (I116443,I116101,I116381);
nor I_6678 (I116460,I116350,I173554);
not I_6679 (I116477,I116460);
nor I_6680 (I116024,I116477,I116186);
nand I_6681 (I116012,I116477,I116398);
nand I_6682 (I116522,I116477,I116203);
nand I_6683 (I116539,I116381,I116522);
nor I_6684 (I116027,I116302,I116539);
nand I_6685 (I116039,I116084,I116477);
nand I_6686 (I116036,I116477,I116302);
nor I_6687 (I116598,I116443,I116460);
nor I_6688 (I116021,I116319,I116598);
and I_6689 (I116033,I116302,I116350);
not I_6690 (I116679,I2905);
or I_6691 (I116696,I279603,I279618);
nand I_6692 (I116713,I279624,I279606);
not I_6693 (I116730,I116713);
and I_6694 (I116747,I116730,I116696);
or I_6695 (I116764,I279609,I279621);
nor I_6696 (I116781,I116764,I279603);
not I_6697 (I116798,I116781);
nor I_6698 (I116815,I116713,I116798);
nand I_6699 (I116832,I116781,I116730);
nor I_6700 (I116849,I116781,I116730);
DFFARX1 I_6701 (I116849,I2898,I116679,I116659,);
nor I_6702 (I116880,I279612,I279600);
or I_6703 (I116897,I116880,I279600);
nor I_6704 (I116914,I279627,I279630);
nand I_6705 (I116931,I116914,I116897);
nand I_6706 (I116948,I116931,I116798);
not I_6707 (I116671,I116948);
nand I_6708 (I116979,I279615,I279606);
nor I_6709 (I116638,I116979,I116747);
not I_6710 (I117010,I116979);
nand I_6711 (I117027,I117010,I116747);
not I_6712 (I116644,I117027);
nor I_6713 (I116647,I116781,I117027);
nor I_6714 (I117072,I116730,I117010);
nor I_6715 (I117089,I116979,I279609);
not I_6716 (I117106,I117089);
nor I_6717 (I116653,I117106,I116815);
nand I_6718 (I116641,I117106,I117027);
nand I_6719 (I117151,I117106,I116832);
nand I_6720 (I117168,I117010,I117151);
nor I_6721 (I116656,I116931,I117168);
nand I_6722 (I116668,I116713,I117106);
nand I_6723 (I116665,I117106,I116931);
nor I_6724 (I117227,I117072,I117089);
nor I_6725 (I116650,I116948,I117227);
and I_6726 (I116662,I116931,I116979);
not I_6727 (I117308,I2905);
or I_6728 (I117325,I90274,I90277);
nand I_6729 (I117342,I90286,I90292);
not I_6730 (I117359,I117342);
and I_6731 (I117376,I117359,I117325);
or I_6732 (I117393,I90298,I90283);
nor I_6733 (I117410,I117393,I90295);
not I_6734 (I117427,I117410);
nor I_6735 (I117444,I117342,I117427);
nand I_6736 (I117461,I117410,I117359);
nor I_6737 (I117478,I117410,I117359);
DFFARX1 I_6738 (I117478,I2898,I117308,I117288,);
nor I_6739 (I117509,I90274,I90289);
or I_6740 (I117526,I117509,I90271);
nor I_6741 (I117543,I90283,I90280);
nand I_6742 (I117560,I117543,I117526);
nand I_6743 (I117577,I117560,I117427);
not I_6744 (I117300,I117577);
nand I_6745 (I117608,I90271,I90280);
nor I_6746 (I117267,I117608,I117376);
not I_6747 (I117639,I117608);
nand I_6748 (I117656,I117639,I117376);
not I_6749 (I117273,I117656);
nor I_6750 (I117276,I117410,I117656);
nor I_6751 (I117701,I117359,I117639);
nor I_6752 (I117718,I117608,I90277);
not I_6753 (I117735,I117718);
nor I_6754 (I117282,I117735,I117444);
nand I_6755 (I117270,I117735,I117656);
nand I_6756 (I117780,I117735,I117461);
nand I_6757 (I117797,I117639,I117780);
nor I_6758 (I117285,I117560,I117797);
nand I_6759 (I117297,I117342,I117735);
nand I_6760 (I117294,I117735,I117560);
nor I_6761 (I117856,I117701,I117718);
nor I_6762 (I117279,I117577,I117856);
and I_6763 (I117291,I117560,I117608);
not I_6764 (I117937,I2905);
or I_6765 (I117954,I2147,I2739);
nand I_6766 (I117971,I2627,I2419);
not I_6767 (I117988,I117971);
and I_6768 (I118005,I117988,I117954);
or I_6769 (I118022,I2643,I2403);
nor I_6770 (I118039,I118022,I2859);
not I_6771 (I118056,I118039);
nor I_6772 (I118073,I117971,I118056);
nand I_6773 (I118090,I118039,I117988);
nor I_6774 (I118107,I118039,I117988);
DFFARX1 I_6775 (I118107,I2898,I117937,I117917,);
nor I_6776 (I118138,I2131,I2547);
or I_6777 (I118155,I118138,I2179);
nor I_6778 (I118172,I2515,I2395);
nand I_6779 (I118189,I118172,I118155);
nand I_6780 (I118206,I118189,I118056);
not I_6781 (I117929,I118206);
nand I_6782 (I118237,I1795,I2715);
nor I_6783 (I117896,I118237,I118005);
not I_6784 (I118268,I118237);
nand I_6785 (I118285,I118268,I118005);
not I_6786 (I117902,I118285);
nor I_6787 (I117905,I118039,I118285);
nor I_6788 (I118330,I117988,I118268);
nor I_6789 (I118347,I118237,I2307);
not I_6790 (I118364,I118347);
nor I_6791 (I117911,I118364,I118073);
nand I_6792 (I117899,I118364,I118285);
nand I_6793 (I118409,I118364,I118090);
nand I_6794 (I118426,I118268,I118409);
nor I_6795 (I117914,I118189,I118426);
nand I_6796 (I117926,I117971,I118364);
nand I_6797 (I117923,I118364,I118189);
nor I_6798 (I118485,I118330,I118347);
nor I_6799 (I117908,I118206,I118485);
and I_6800 (I117920,I118189,I118237);
not I_6801 (I118566,I2905);
or I_6802 (I118583,I433851,I433824);
nand I_6803 (I118600,I433854,I433833);
not I_6804 (I118617,I118600);
and I_6805 (I118634,I118617,I118583);
or I_6806 (I118651,I433842,I433827);
nor I_6807 (I118668,I118651,I433845);
not I_6808 (I118685,I118668);
nor I_6809 (I118702,I118600,I118685);
nand I_6810 (I118719,I118668,I118617);
nor I_6811 (I118736,I118668,I118617);
DFFARX1 I_6812 (I118736,I2898,I118566,I118546,);
nor I_6813 (I118767,I433848,I433827);
or I_6814 (I118784,I118767,I433830);
nor I_6815 (I118801,I433836,I433824);
nand I_6816 (I118818,I118801,I118784);
nand I_6817 (I118835,I118818,I118685);
not I_6818 (I118558,I118835);
nand I_6819 (I118866,I433830,I433839);
nor I_6820 (I118525,I118866,I118634);
not I_6821 (I118897,I118866);
nand I_6822 (I118914,I118897,I118634);
not I_6823 (I118531,I118914);
nor I_6824 (I118534,I118668,I118914);
nor I_6825 (I118959,I118617,I118897);
nor I_6826 (I118976,I118866,I433857);
not I_6827 (I118993,I118976);
nor I_6828 (I118540,I118993,I118702);
nand I_6829 (I118528,I118993,I118914);
nand I_6830 (I119038,I118993,I118719);
nand I_6831 (I119055,I118897,I119038);
nor I_6832 (I118543,I118818,I119055);
nand I_6833 (I118555,I118600,I118993);
nand I_6834 (I118552,I118993,I118818);
nor I_6835 (I119114,I118959,I118976);
nor I_6836 (I118537,I118835,I119114);
and I_6837 (I118549,I118818,I118866);
not I_6838 (I119195,I2905);
or I_6839 (I119212,I73920,I73923);
nand I_6840 (I119229,I73932,I73938);
not I_6841 (I119246,I119229);
and I_6842 (I119263,I119246,I119212);
or I_6843 (I119280,I73944,I73929);
nor I_6844 (I119297,I119280,I73941);
not I_6845 (I119314,I119297);
nor I_6846 (I119331,I119229,I119314);
nand I_6847 (I119348,I119297,I119246);
nor I_6848 (I119365,I119297,I119246);
DFFARX1 I_6849 (I119365,I2898,I119195,I119175,);
nor I_6850 (I119396,I73920,I73935);
or I_6851 (I119413,I119396,I73917);
nor I_6852 (I119430,I73929,I73926);
nand I_6853 (I119447,I119430,I119413);
nand I_6854 (I119464,I119447,I119314);
not I_6855 (I119187,I119464);
nand I_6856 (I119495,I73917,I73926);
nor I_6857 (I119154,I119495,I119263);
not I_6858 (I119526,I119495);
nand I_6859 (I119543,I119526,I119263);
not I_6860 (I119160,I119543);
nor I_6861 (I119163,I119297,I119543);
nor I_6862 (I119588,I119246,I119526);
nor I_6863 (I119605,I119495,I73923);
not I_6864 (I119622,I119605);
nor I_6865 (I119169,I119622,I119331);
nand I_6866 (I119157,I119622,I119543);
nand I_6867 (I119667,I119622,I119348);
nand I_6868 (I119684,I119526,I119667);
nor I_6869 (I119172,I119447,I119684);
nand I_6870 (I119184,I119229,I119622);
nand I_6871 (I119181,I119622,I119447);
nor I_6872 (I119743,I119588,I119605);
nor I_6873 (I119166,I119464,I119743);
and I_6874 (I119178,I119447,I119495);
not I_6875 (I119824,I2905);
or I_6876 (I119841,I74549,I74552);
nand I_6877 (I119858,I74561,I74567);
not I_6878 (I119875,I119858);
and I_6879 (I119892,I119875,I119841);
or I_6880 (I119909,I74573,I74558);
nor I_6881 (I119926,I119909,I74570);
not I_6882 (I119943,I119926);
nor I_6883 (I119960,I119858,I119943);
nand I_6884 (I119977,I119926,I119875);
nor I_6885 (I119994,I119926,I119875);
DFFARX1 I_6886 (I119994,I2898,I119824,I119804,);
nor I_6887 (I120025,I74549,I74564);
or I_6888 (I120042,I120025,I74546);
nor I_6889 (I120059,I74558,I74555);
nand I_6890 (I120076,I120059,I120042);
nand I_6891 (I120093,I120076,I119943);
not I_6892 (I119816,I120093);
nand I_6893 (I120124,I74546,I74555);
nor I_6894 (I119783,I120124,I119892);
not I_6895 (I120155,I120124);
nand I_6896 (I120172,I120155,I119892);
not I_6897 (I119789,I120172);
nor I_6898 (I119792,I119926,I120172);
nor I_6899 (I120217,I119875,I120155);
nor I_6900 (I120234,I120124,I74552);
not I_6901 (I120251,I120234);
nor I_6902 (I119798,I120251,I119960);
nand I_6903 (I119786,I120251,I120172);
nand I_6904 (I120296,I120251,I119977);
nand I_6905 (I120313,I120155,I120296);
nor I_6906 (I119801,I120076,I120313);
nand I_6907 (I119813,I119858,I120251);
nand I_6908 (I119810,I120251,I120076);
nor I_6909 (I120372,I120217,I120234);
nor I_6910 (I119795,I120093,I120372);
and I_6911 (I119807,I120076,I120124);
not I_6912 (I120453,I2905);
or I_6913 (I120470,I87758,I87761);
nand I_6914 (I120487,I87770,I87776);
not I_6915 (I120504,I120487);
and I_6916 (I120521,I120504,I120470);
or I_6917 (I120538,I87782,I87767);
nor I_6918 (I120555,I120538,I87779);
not I_6919 (I120572,I120555);
nor I_6920 (I120589,I120487,I120572);
nand I_6921 (I120606,I120555,I120504);
nor I_6922 (I120623,I120555,I120504);
DFFARX1 I_6923 (I120623,I2898,I120453,I120433,);
nor I_6924 (I120654,I87758,I87773);
or I_6925 (I120671,I120654,I87755);
nor I_6926 (I120688,I87767,I87764);
nand I_6927 (I120705,I120688,I120671);
nand I_6928 (I120722,I120705,I120572);
not I_6929 (I120445,I120722);
nand I_6930 (I120753,I87755,I87764);
nor I_6931 (I120412,I120753,I120521);
not I_6932 (I120784,I120753);
nand I_6933 (I120801,I120784,I120521);
not I_6934 (I120418,I120801);
nor I_6935 (I120421,I120555,I120801);
nor I_6936 (I120846,I120504,I120784);
nor I_6937 (I120863,I120753,I87761);
not I_6938 (I120880,I120863);
nor I_6939 (I120427,I120880,I120589);
nand I_6940 (I120415,I120880,I120801);
nand I_6941 (I120925,I120880,I120606);
nand I_6942 (I120942,I120784,I120925);
nor I_6943 (I120430,I120705,I120942);
nand I_6944 (I120442,I120487,I120880);
nand I_6945 (I120439,I120880,I120705);
nor I_6946 (I121001,I120846,I120863);
nor I_6947 (I120424,I120722,I121001);
and I_6948 (I120436,I120705,I120753);
not I_6949 (I121082,I2905);
or I_6950 (I121099,I249768,I249783);
nand I_6951 (I121116,I249789,I249771);
not I_6952 (I121133,I121116);
and I_6953 (I121150,I121133,I121099);
or I_6954 (I121167,I249774,I249786);
nor I_6955 (I121184,I121167,I249768);
not I_6956 (I121201,I121184);
nor I_6957 (I121218,I121116,I121201);
nand I_6958 (I121235,I121184,I121133);
nor I_6959 (I121252,I121184,I121133);
DFFARX1 I_6960 (I121252,I2898,I121082,I121062,);
nor I_6961 (I121283,I249777,I249765);
or I_6962 (I121300,I121283,I249765);
nor I_6963 (I121317,I249792,I249795);
nand I_6964 (I121334,I121317,I121300);
nand I_6965 (I121351,I121334,I121201);
not I_6966 (I121074,I121351);
nand I_6967 (I121382,I249780,I249771);
nor I_6968 (I121041,I121382,I121150);
not I_6969 (I121413,I121382);
nand I_6970 (I121430,I121413,I121150);
not I_6971 (I121047,I121430);
nor I_6972 (I121050,I121184,I121430);
nor I_6973 (I121475,I121133,I121413);
nor I_6974 (I121492,I121382,I249774);
not I_6975 (I121509,I121492);
nor I_6976 (I121056,I121509,I121218);
nand I_6977 (I121044,I121509,I121430);
nand I_6978 (I121554,I121509,I121235);
nand I_6979 (I121571,I121413,I121554);
nor I_6980 (I121059,I121334,I121571);
nand I_6981 (I121071,I121116,I121509);
nand I_6982 (I121068,I121509,I121334);
nor I_6983 (I121630,I121475,I121492);
nor I_6984 (I121053,I121351,I121630);
and I_6985 (I121065,I121334,I121382);
not I_6986 (I121711,I2905);
or I_6987 (I121728,I235998,I236013);
nand I_6988 (I121745,I236019,I236001);
not I_6989 (I121762,I121745);
and I_6990 (I121779,I121762,I121728);
or I_6991 (I121796,I236004,I236016);
nor I_6992 (I121813,I121796,I235998);
not I_6993 (I121830,I121813);
nor I_6994 (I121847,I121745,I121830);
nand I_6995 (I121864,I121813,I121762);
nor I_6996 (I121881,I121813,I121762);
DFFARX1 I_6997 (I121881,I2898,I121711,I121691,);
nor I_6998 (I121912,I236007,I235995);
or I_6999 (I121929,I121912,I235995);
nor I_7000 (I121946,I236022,I236025);
nand I_7001 (I121963,I121946,I121929);
nand I_7002 (I121980,I121963,I121830);
not I_7003 (I121703,I121980);
nand I_7004 (I122011,I236010,I236001);
nor I_7005 (I121670,I122011,I121779);
not I_7006 (I122042,I122011);
nand I_7007 (I122059,I122042,I121779);
not I_7008 (I121676,I122059);
nor I_7009 (I121679,I121813,I122059);
nor I_7010 (I122104,I121762,I122042);
nor I_7011 (I122121,I122011,I236004);
not I_7012 (I122138,I122121);
nor I_7013 (I121685,I122138,I121847);
nand I_7014 (I121673,I122138,I122059);
nand I_7015 (I122183,I122138,I121864);
nand I_7016 (I122200,I122042,I122183);
nor I_7017 (I121688,I121963,I122200);
nand I_7018 (I121700,I121745,I122138);
nand I_7019 (I121697,I122138,I121963);
nor I_7020 (I122259,I122104,I122121);
nor I_7021 (I121682,I121980,I122259);
and I_7022 (I121694,I121963,I122011);
not I_7023 (I122340,I2905);
or I_7024 (I122357,I231408,I231423);
nand I_7025 (I122374,I231429,I231411);
not I_7026 (I122391,I122374);
and I_7027 (I122408,I122391,I122357);
or I_7028 (I122425,I231414,I231426);
nor I_7029 (I122442,I122425,I231408);
not I_7030 (I122459,I122442);
nor I_7031 (I122476,I122374,I122459);
nand I_7032 (I122493,I122442,I122391);
nor I_7033 (I122510,I122442,I122391);
DFFARX1 I_7034 (I122510,I2898,I122340,I122320,);
nor I_7035 (I122541,I231417,I231405);
or I_7036 (I122558,I122541,I231405);
nor I_7037 (I122575,I231432,I231435);
nand I_7038 (I122592,I122575,I122558);
nand I_7039 (I122609,I122592,I122459);
not I_7040 (I122332,I122609);
nand I_7041 (I122640,I231420,I231411);
nor I_7042 (I122299,I122640,I122408);
not I_7043 (I122671,I122640);
nand I_7044 (I122688,I122671,I122408);
not I_7045 (I122305,I122688);
nor I_7046 (I122308,I122442,I122688);
nor I_7047 (I122733,I122391,I122671);
nor I_7048 (I122750,I122640,I231414);
not I_7049 (I122767,I122750);
nor I_7050 (I122314,I122767,I122476);
nand I_7051 (I122302,I122767,I122688);
nand I_7052 (I122812,I122767,I122493);
nand I_7053 (I122829,I122671,I122812);
nor I_7054 (I122317,I122592,I122829);
nand I_7055 (I122329,I122374,I122767);
nand I_7056 (I122326,I122767,I122592);
nor I_7057 (I122888,I122733,I122750);
nor I_7058 (I122311,I122609,I122888);
and I_7059 (I122323,I122592,I122640);
not I_7060 (I122969,I2905);
or I_7061 (I122986,I189727,I189724);
nand I_7062 (I123003,I189736,I189733);
not I_7063 (I123020,I123003);
and I_7064 (I123037,I123020,I122986);
or I_7065 (I123054,I189721,I189730);
nor I_7066 (I123071,I123054,I189730);
not I_7067 (I123088,I123071);
nor I_7068 (I123105,I123003,I123088);
nand I_7069 (I123122,I123071,I123020);
nor I_7070 (I123139,I123071,I123020);
DFFARX1 I_7071 (I123139,I2898,I122969,I122949,);
nor I_7072 (I123170,I189739,I189721);
or I_7073 (I123187,I123170,I189727);
nor I_7074 (I123204,I189724,I189745);
nand I_7075 (I123221,I123204,I123187);
nand I_7076 (I123238,I123221,I123088);
not I_7077 (I122961,I123238);
nand I_7078 (I123269,I189736,I189742);
nor I_7079 (I122928,I123269,I123037);
not I_7080 (I123300,I123269);
nand I_7081 (I123317,I123300,I123037);
not I_7082 (I122934,I123317);
nor I_7083 (I122937,I123071,I123317);
nor I_7084 (I123362,I123020,I123300);
nor I_7085 (I123379,I123269,I189733);
not I_7086 (I123396,I123379);
nor I_7087 (I122943,I123396,I123105);
nand I_7088 (I122931,I123396,I123317);
nand I_7089 (I123441,I123396,I123122);
nand I_7090 (I123458,I123300,I123441);
nor I_7091 (I122946,I123221,I123458);
nand I_7092 (I122958,I123003,I123396);
nand I_7093 (I122955,I123396,I123221);
nor I_7094 (I123517,I123362,I123379);
nor I_7095 (I122940,I123238,I123517);
and I_7096 (I122952,I123221,I123269);
not I_7097 (I123598,I2905);
or I_7098 (I123615,I46483,I46477);
nand I_7099 (I123632,I46492,I46465);
not I_7100 (I123649,I123632);
and I_7101 (I123666,I123649,I123615);
or I_7102 (I123683,I46474,I46489);
nor I_7103 (I123700,I123683,I46480);
not I_7104 (I123717,I123700);
nor I_7105 (I123734,I123632,I123717);
nand I_7106 (I123751,I123700,I123649);
nor I_7107 (I123768,I123700,I123649);
DFFARX1 I_7108 (I123768,I2898,I123598,I123578,);
nor I_7109 (I123799,I46486,I46471);
or I_7110 (I123816,I123799,I46462);
nor I_7111 (I123833,I46495,I46468);
nand I_7112 (I123850,I123833,I123816);
nand I_7113 (I123867,I123850,I123717);
not I_7114 (I123590,I123867);
nand I_7115 (I123898,I46462,I46498);
nor I_7116 (I123557,I123898,I123666);
not I_7117 (I123929,I123898);
nand I_7118 (I123946,I123929,I123666);
not I_7119 (I123563,I123946);
nor I_7120 (I123566,I123700,I123946);
nor I_7121 (I123991,I123649,I123929);
nor I_7122 (I124008,I123898,I46465);
not I_7123 (I124025,I124008);
nor I_7124 (I123572,I124025,I123734);
nand I_7125 (I123560,I124025,I123946);
nand I_7126 (I124070,I124025,I123751);
nand I_7127 (I124087,I123929,I124070);
nor I_7128 (I123575,I123850,I124087);
nand I_7129 (I123587,I123632,I124025);
nand I_7130 (I123584,I124025,I123850);
nor I_7131 (I124146,I123991,I124008);
nor I_7132 (I123569,I123867,I124146);
and I_7133 (I123581,I123850,I123898);
not I_7134 (I124227,I2905);
or I_7135 (I124244,I271953,I271968);
nand I_7136 (I124261,I271974,I271956);
not I_7137 (I124278,I124261);
and I_7138 (I124295,I124278,I124244);
or I_7139 (I124312,I271959,I271971);
nor I_7140 (I124329,I124312,I271953);
not I_7141 (I124346,I124329);
nor I_7142 (I124363,I124261,I124346);
nand I_7143 (I124380,I124329,I124278);
nor I_7144 (I124397,I124329,I124278);
DFFARX1 I_7145 (I124397,I2898,I124227,I124207,);
nor I_7146 (I124428,I271962,I271950);
or I_7147 (I124445,I124428,I271950);
nor I_7148 (I124462,I271977,I271980);
nand I_7149 (I124479,I124462,I124445);
nand I_7150 (I124496,I124479,I124346);
not I_7151 (I124219,I124496);
nand I_7152 (I124527,I271965,I271956);
nor I_7153 (I124186,I124527,I124295);
not I_7154 (I124558,I124527);
nand I_7155 (I124575,I124558,I124295);
not I_7156 (I124192,I124575);
nor I_7157 (I124195,I124329,I124575);
nor I_7158 (I124620,I124278,I124558);
nor I_7159 (I124637,I124527,I271959);
not I_7160 (I124654,I124637);
nor I_7161 (I124201,I124654,I124363);
nand I_7162 (I124189,I124654,I124575);
nand I_7163 (I124699,I124654,I124380);
nand I_7164 (I124716,I124558,I124699);
nor I_7165 (I124204,I124479,I124716);
nand I_7166 (I124216,I124261,I124654);
nand I_7167 (I124213,I124654,I124479);
nor I_7168 (I124775,I124620,I124637);
nor I_7169 (I124198,I124496,I124775);
and I_7170 (I124210,I124479,I124527);
not I_7171 (I124856,I2905);
or I_7172 (I124873,I75807,I75810);
nand I_7173 (I124890,I75819,I75825);
not I_7174 (I124907,I124890);
and I_7175 (I124924,I124907,I124873);
or I_7176 (I124941,I75831,I75816);
nor I_7177 (I124958,I124941,I75828);
not I_7178 (I124975,I124958);
nor I_7179 (I124992,I124890,I124975);
nand I_7180 (I125009,I124958,I124907);
nor I_7181 (I125026,I124958,I124907);
DFFARX1 I_7182 (I125026,I2898,I124856,I124836,);
nor I_7183 (I125057,I75807,I75822);
or I_7184 (I125074,I125057,I75804);
nor I_7185 (I125091,I75816,I75813);
nand I_7186 (I125108,I125091,I125074);
nand I_7187 (I125125,I125108,I124975);
not I_7188 (I124848,I125125);
nand I_7189 (I125156,I75804,I75813);
nor I_7190 (I124815,I125156,I124924);
not I_7191 (I125187,I125156);
nand I_7192 (I125204,I125187,I124924);
not I_7193 (I124821,I125204);
nor I_7194 (I124824,I124958,I125204);
nor I_7195 (I125249,I124907,I125187);
nor I_7196 (I125266,I125156,I75810);
not I_7197 (I125283,I125266);
nor I_7198 (I124830,I125283,I124992);
nand I_7199 (I124818,I125283,I125204);
nand I_7200 (I125328,I125283,I125009);
nand I_7201 (I125345,I125187,I125328);
nor I_7202 (I124833,I125108,I125345);
nand I_7203 (I124845,I124890,I125283);
nand I_7204 (I124842,I125283,I125108);
nor I_7205 (I125404,I125249,I125266);
nor I_7206 (I124827,I125125,I125404);
and I_7207 (I124839,I125108,I125156);
not I_7208 (I125485,I2905);
or I_7209 (I125502,I164043,I164061);
nand I_7210 (I125519,I164064,I164058);
not I_7211 (I125536,I125519);
and I_7212 (I125553,I125536,I125502);
or I_7213 (I125570,I164052,I164034);
nor I_7214 (I125587,I125570,I164040);
not I_7215 (I125604,I125587);
nor I_7216 (I125621,I125519,I125604);
nand I_7217 (I125638,I125587,I125536);
nor I_7218 (I125655,I125587,I125536);
DFFARX1 I_7219 (I125655,I2898,I125485,I125465,);
nor I_7220 (I125686,I164046,I164067);
or I_7221 (I125703,I125686,I164037);
nor I_7222 (I125720,I164049,I164040);
nand I_7223 (I125737,I125720,I125703);
nand I_7224 (I125754,I125737,I125604);
not I_7225 (I125477,I125754);
nand I_7226 (I125785,I164055,I164037);
nor I_7227 (I125444,I125785,I125553);
not I_7228 (I125816,I125785);
nand I_7229 (I125833,I125816,I125553);
not I_7230 (I125450,I125833);
nor I_7231 (I125453,I125587,I125833);
nor I_7232 (I125878,I125536,I125816);
nor I_7233 (I125895,I125785,I164034);
not I_7234 (I125912,I125895);
nor I_7235 (I125459,I125912,I125621);
nand I_7236 (I125447,I125912,I125833);
nand I_7237 (I125957,I125912,I125638);
nand I_7238 (I125974,I125816,I125957);
nor I_7239 (I125462,I125737,I125974);
nand I_7240 (I125474,I125519,I125912);
nand I_7241 (I125471,I125912,I125737);
nor I_7242 (I126033,I125878,I125895);
nor I_7243 (I125456,I125754,I126033);
and I_7244 (I125468,I125737,I125785);
not I_7245 (I126114,I2905);
or I_7246 (I126131,I168803,I168821);
nand I_7247 (I126148,I168824,I168818);
not I_7248 (I126165,I126148);
and I_7249 (I126182,I126165,I126131);
or I_7250 (I126199,I168812,I168794);
nor I_7251 (I126216,I126199,I168800);
not I_7252 (I126233,I126216);
nor I_7253 (I126250,I126148,I126233);
nand I_7254 (I126267,I126216,I126165);
nor I_7255 (I126284,I126216,I126165);
DFFARX1 I_7256 (I126284,I2898,I126114,I126094,);
nor I_7257 (I126315,I168806,I168827);
or I_7258 (I126332,I126315,I168797);
nor I_7259 (I126349,I168809,I168800);
nand I_7260 (I126366,I126349,I126332);
nand I_7261 (I126383,I126366,I126233);
not I_7262 (I126106,I126383);
nand I_7263 (I126414,I168815,I168797);
nor I_7264 (I126073,I126414,I126182);
not I_7265 (I126445,I126414);
nand I_7266 (I126462,I126445,I126182);
not I_7267 (I126079,I126462);
nor I_7268 (I126082,I126216,I126462);
nor I_7269 (I126507,I126165,I126445);
nor I_7270 (I126524,I126414,I168794);
not I_7271 (I126541,I126524);
nor I_7272 (I126088,I126541,I126250);
nand I_7273 (I126076,I126541,I126462);
nand I_7274 (I126586,I126541,I126267);
nand I_7275 (I126603,I126445,I126586);
nor I_7276 (I126091,I126366,I126603);
nand I_7277 (I126103,I126148,I126541);
nand I_7278 (I126100,I126541,I126366);
nor I_7279 (I126662,I126507,I126524);
nor I_7280 (I126085,I126383,I126662);
and I_7281 (I126097,I126366,I126414);
not I_7282 (I126743,I2905);
or I_7283 (I126760,I61340,I61343);
nand I_7284 (I126777,I61352,I61358);
not I_7285 (I126794,I126777);
and I_7286 (I126811,I126794,I126760);
or I_7287 (I126828,I61364,I61349);
nor I_7288 (I126845,I126828,I61361);
not I_7289 (I126862,I126845);
nor I_7290 (I126879,I126777,I126862);
nand I_7291 (I126896,I126845,I126794);
nor I_7292 (I126913,I126845,I126794);
DFFARX1 I_7293 (I126913,I2898,I126743,I126723,);
nor I_7294 (I126944,I61340,I61355);
or I_7295 (I126961,I126944,I61337);
nor I_7296 (I126978,I61349,I61346);
nand I_7297 (I126995,I126978,I126961);
nand I_7298 (I127012,I126995,I126862);
not I_7299 (I126735,I127012);
nand I_7300 (I127043,I61337,I61346);
nor I_7301 (I126702,I127043,I126811);
not I_7302 (I127074,I127043);
nand I_7303 (I127091,I127074,I126811);
not I_7304 (I126708,I127091);
nor I_7305 (I126711,I126845,I127091);
nor I_7306 (I127136,I126794,I127074);
nor I_7307 (I127153,I127043,I61343);
not I_7308 (I127170,I127153);
nor I_7309 (I126717,I127170,I126879);
nand I_7310 (I126705,I127170,I127091);
nand I_7311 (I127215,I127170,I126896);
nand I_7312 (I127232,I127074,I127215);
nor I_7313 (I126720,I126995,I127232);
nand I_7314 (I126732,I126777,I127170);
nand I_7315 (I126729,I127170,I126995);
nor I_7316 (I127291,I127136,I127153);
nor I_7317 (I126714,I127012,I127291);
and I_7318 (I126726,I126995,I127043);
not I_7319 (I127372,I2905);
or I_7320 (I127389,I159963,I159981);
nand I_7321 (I127406,I159984,I159978);
not I_7322 (I127423,I127406);
and I_7323 (I127440,I127423,I127389);
or I_7324 (I127457,I159972,I159954);
nor I_7325 (I127474,I127457,I159960);
not I_7326 (I127491,I127474);
nor I_7327 (I127508,I127406,I127491);
nand I_7328 (I127525,I127474,I127423);
nor I_7329 (I127542,I127474,I127423);
DFFARX1 I_7330 (I127542,I2898,I127372,I127352,);
nor I_7331 (I127573,I159966,I159987);
or I_7332 (I127590,I127573,I159957);
nor I_7333 (I127607,I159969,I159960);
nand I_7334 (I127624,I127607,I127590);
nand I_7335 (I127641,I127624,I127491);
not I_7336 (I127364,I127641);
nand I_7337 (I127672,I159975,I159957);
nor I_7338 (I127331,I127672,I127440);
not I_7339 (I127703,I127672);
nand I_7340 (I127720,I127703,I127440);
not I_7341 (I127337,I127720);
nor I_7342 (I127340,I127474,I127720);
nor I_7343 (I127765,I127423,I127703);
nor I_7344 (I127782,I127672,I159954);
not I_7345 (I127799,I127782);
nor I_7346 (I127346,I127799,I127508);
nand I_7347 (I127334,I127799,I127720);
nand I_7348 (I127844,I127799,I127525);
nand I_7349 (I127861,I127703,I127844);
nor I_7350 (I127349,I127624,I127861);
nand I_7351 (I127361,I127406,I127799);
nand I_7352 (I127358,I127799,I127624);
nor I_7353 (I127920,I127765,I127782);
nor I_7354 (I127343,I127641,I127920);
and I_7355 (I127355,I127624,I127672);
not I_7356 (I128001,I2905);
or I_7357 (I128018,I232938,I232953);
nand I_7358 (I128035,I232959,I232941);
not I_7359 (I128052,I128035);
and I_7360 (I128069,I128052,I128018);
or I_7361 (I128086,I232944,I232956);
nor I_7362 (I128103,I128086,I232938);
not I_7363 (I128120,I128103);
nor I_7364 (I128137,I128035,I128120);
nand I_7365 (I128154,I128103,I128052);
nor I_7366 (I128171,I128103,I128052);
DFFARX1 I_7367 (I128171,I2898,I128001,I127981,);
nor I_7368 (I128202,I232947,I232935);
or I_7369 (I128219,I128202,I232935);
nor I_7370 (I128236,I232962,I232965);
nand I_7371 (I128253,I128236,I128219);
nand I_7372 (I128270,I128253,I128120);
not I_7373 (I127993,I128270);
nand I_7374 (I128301,I232950,I232941);
nor I_7375 (I127960,I128301,I128069);
not I_7376 (I128332,I128301);
nand I_7377 (I128349,I128332,I128069);
not I_7378 (I127966,I128349);
nor I_7379 (I127969,I128103,I128349);
nor I_7380 (I128394,I128052,I128332);
nor I_7381 (I128411,I128301,I232944);
not I_7382 (I128428,I128411);
nor I_7383 (I127975,I128428,I128137);
nand I_7384 (I127963,I128428,I128349);
nand I_7385 (I128473,I128428,I128154);
nand I_7386 (I128490,I128332,I128473);
nor I_7387 (I127978,I128253,I128490);
nand I_7388 (I127990,I128035,I128428);
nand I_7389 (I127987,I128428,I128253);
nor I_7390 (I128549,I128394,I128411);
nor I_7391 (I127972,I128270,I128549);
and I_7392 (I127984,I128253,I128301);
not I_7393 (I128630,I2905);
or I_7394 (I128647,I43355,I43349);
nand I_7395 (I128664,I43364,I43337);
not I_7396 (I128681,I128664);
and I_7397 (I128698,I128681,I128647);
or I_7398 (I128715,I43346,I43361);
nor I_7399 (I128732,I128715,I43352);
not I_7400 (I128749,I128732);
nor I_7401 (I128766,I128664,I128749);
nand I_7402 (I128783,I128732,I128681);
nor I_7403 (I128800,I128732,I128681);
DFFARX1 I_7404 (I128800,I2898,I128630,I128610,);
nor I_7405 (I128831,I43358,I43343);
or I_7406 (I128848,I128831,I43334);
nor I_7407 (I128865,I43367,I43340);
nand I_7408 (I128882,I128865,I128848);
nand I_7409 (I128899,I128882,I128749);
not I_7410 (I128622,I128899);
nand I_7411 (I128930,I43334,I43370);
nor I_7412 (I128589,I128930,I128698);
not I_7413 (I128961,I128930);
nand I_7414 (I128978,I128961,I128698);
not I_7415 (I128595,I128978);
nor I_7416 (I128598,I128732,I128978);
nor I_7417 (I129023,I128681,I128961);
nor I_7418 (I129040,I128930,I43337);
not I_7419 (I129057,I129040);
nor I_7420 (I128604,I129057,I128766);
nand I_7421 (I128592,I129057,I128978);
nand I_7422 (I129102,I129057,I128783);
nand I_7423 (I129119,I128961,I129102);
nor I_7424 (I128607,I128882,I129119);
nand I_7425 (I128619,I128664,I129057);
nand I_7426 (I128616,I129057,I128882);
nor I_7427 (I129178,I129023,I129040);
nor I_7428 (I128601,I128899,I129178);
and I_7429 (I128613,I128882,I128930);
not I_7430 (I129259,I2905);
or I_7431 (I129276,I52739,I52733);
nand I_7432 (I129293,I52748,I52721);
not I_7433 (I129310,I129293);
and I_7434 (I129327,I129310,I129276);
or I_7435 (I129344,I52730,I52745);
nor I_7436 (I129361,I129344,I52736);
not I_7437 (I129378,I129361);
nor I_7438 (I129395,I129293,I129378);
nand I_7439 (I129412,I129361,I129310);
nor I_7440 (I129429,I129361,I129310);
DFFARX1 I_7441 (I129429,I2898,I129259,I129239,);
nor I_7442 (I129460,I52742,I52727);
or I_7443 (I129477,I129460,I52718);
nor I_7444 (I129494,I52751,I52724);
nand I_7445 (I129511,I129494,I129477);
nand I_7446 (I129528,I129511,I129378);
not I_7447 (I129251,I129528);
nand I_7448 (I129559,I52718,I52754);
nor I_7449 (I129218,I129559,I129327);
not I_7450 (I129590,I129559);
nand I_7451 (I129607,I129590,I129327);
not I_7452 (I129224,I129607);
nor I_7453 (I129227,I129361,I129607);
nor I_7454 (I129652,I129310,I129590);
nor I_7455 (I129669,I129559,I52721);
not I_7456 (I129686,I129669);
nor I_7457 (I129233,I129686,I129395);
nand I_7458 (I129221,I129686,I129607);
nand I_7459 (I129731,I129686,I129412);
nand I_7460 (I129748,I129590,I129731);
nor I_7461 (I129236,I129511,I129748);
nand I_7462 (I129248,I129293,I129686);
nand I_7463 (I129245,I129686,I129511);
nor I_7464 (I129807,I129652,I129669);
nor I_7465 (I129230,I129528,I129807);
and I_7466 (I129242,I129511,I129559);
not I_7467 (I129888,I2905);
or I_7468 (I129905,I35353,I35350);
nand I_7469 (I129922,I35344,I35365);
not I_7470 (I129939,I129922);
and I_7471 (I129956,I129939,I129905);
or I_7472 (I129973,I35359,I35371);
nor I_7473 (I129990,I129973,I35353);
not I_7474 (I130007,I129990);
nor I_7475 (I130024,I129922,I130007);
nand I_7476 (I130041,I129990,I129939);
nor I_7477 (I130058,I129990,I129939);
DFFARX1 I_7478 (I130058,I2898,I129888,I129868,);
nor I_7479 (I130089,I35356,I35356);
or I_7480 (I130106,I130089,I35362);
nor I_7481 (I130123,I35347,I35350);
nand I_7482 (I130140,I130123,I130106);
nand I_7483 (I130157,I130140,I130007);
not I_7484 (I129880,I130157);
nand I_7485 (I130188,I35368,I35344);
nor I_7486 (I129847,I130188,I129956);
not I_7487 (I130219,I130188);
nand I_7488 (I130236,I130219,I129956);
not I_7489 (I129853,I130236);
nor I_7490 (I129856,I129990,I130236);
nor I_7491 (I130281,I129939,I130219);
nor I_7492 (I130298,I130188,I35347);
not I_7493 (I130315,I130298);
nor I_7494 (I129862,I130315,I130024);
nand I_7495 (I129850,I130315,I130236);
nand I_7496 (I130360,I130315,I130041);
nand I_7497 (I130377,I130219,I130360);
nor I_7498 (I129865,I130140,I130377);
nand I_7499 (I129877,I129922,I130315);
nand I_7500 (I129874,I130315,I130140);
nor I_7501 (I130436,I130281,I130298);
nor I_7502 (I129859,I130157,I130436);
and I_7503 (I129871,I130140,I130188);
not I_7504 (I130517,I2905);
or I_7505 (I130534,I247473,I247488);
nand I_7506 (I130551,I247494,I247476);
not I_7507 (I130568,I130551);
and I_7508 (I130585,I130568,I130534);
or I_7509 (I130602,I247479,I247491);
nor I_7510 (I130619,I130602,I247473);
not I_7511 (I130636,I130619);
nor I_7512 (I130653,I130551,I130636);
nand I_7513 (I130670,I130619,I130568);
nor I_7514 (I130687,I130619,I130568);
DFFARX1 I_7515 (I130687,I2898,I130517,I130497,);
nor I_7516 (I130718,I247482,I247470);
or I_7517 (I130735,I130718,I247470);
nor I_7518 (I130752,I247497,I247500);
nand I_7519 (I130769,I130752,I130735);
nand I_7520 (I130786,I130769,I130636);
not I_7521 (I130509,I130786);
nand I_7522 (I130817,I247485,I247476);
nor I_7523 (I130476,I130817,I130585);
not I_7524 (I130848,I130817);
nand I_7525 (I130865,I130848,I130585);
not I_7526 (I130482,I130865);
nor I_7527 (I130485,I130619,I130865);
nor I_7528 (I130910,I130568,I130848);
nor I_7529 (I130927,I130817,I247479);
not I_7530 (I130944,I130927);
nor I_7531 (I130491,I130944,I130653);
nand I_7532 (I130479,I130944,I130865);
nand I_7533 (I130989,I130944,I130670);
nand I_7534 (I131006,I130848,I130989);
nor I_7535 (I130494,I130769,I131006);
nand I_7536 (I130506,I130551,I130944);
nand I_7537 (I130503,I130944,I130769);
nor I_7538 (I131065,I130910,I130927);
nor I_7539 (I130488,I130786,I131065);
and I_7540 (I130500,I130769,I130817);
not I_7541 (I131146,I2905);
or I_7542 (I131163,I410850,I410823);
nand I_7543 (I131180,I410853,I410832);
not I_7544 (I131197,I131180);
and I_7545 (I131214,I131197,I131163);
or I_7546 (I131231,I410841,I410826);
nor I_7547 (I131248,I131231,I410844);
not I_7548 (I131265,I131248);
nor I_7549 (I131282,I131180,I131265);
nand I_7550 (I131299,I131248,I131197);
nor I_7551 (I131316,I131248,I131197);
DFFARX1 I_7552 (I131316,I2898,I131146,I131126,);
nor I_7553 (I131347,I410847,I410826);
or I_7554 (I131364,I131347,I410829);
nor I_7555 (I131381,I410835,I410823);
nand I_7556 (I131398,I131381,I131364);
nand I_7557 (I131415,I131398,I131265);
not I_7558 (I131138,I131415);
nand I_7559 (I131446,I410829,I410838);
nor I_7560 (I131105,I131446,I131214);
not I_7561 (I131477,I131446);
nand I_7562 (I131494,I131477,I131214);
not I_7563 (I131111,I131494);
nor I_7564 (I131114,I131248,I131494);
nor I_7565 (I131539,I131197,I131477);
nor I_7566 (I131556,I131446,I410856);
not I_7567 (I131573,I131556);
nor I_7568 (I131120,I131573,I131282);
nand I_7569 (I131108,I131573,I131494);
nand I_7570 (I131618,I131573,I131299);
nand I_7571 (I131635,I131477,I131618);
nor I_7572 (I131123,I131398,I131635);
nand I_7573 (I131135,I131180,I131573);
nand I_7574 (I131132,I131573,I131398);
nor I_7575 (I131694,I131539,I131556);
nor I_7576 (I131117,I131415,I131694);
and I_7577 (I131129,I131398,I131446);
not I_7578 (I131775,I2905);
or I_7579 (I131792,I95935,I95938);
nand I_7580 (I131809,I95947,I95953);
not I_7581 (I131826,I131809);
and I_7582 (I131843,I131826,I131792);
or I_7583 (I131860,I95959,I95944);
nor I_7584 (I131877,I131860,I95956);
not I_7585 (I131894,I131877);
nor I_7586 (I131911,I131809,I131894);
nand I_7587 (I131928,I131877,I131826);
nor I_7588 (I131945,I131877,I131826);
DFFARX1 I_7589 (I131945,I2898,I131775,I131755,);
nor I_7590 (I131976,I95935,I95950);
or I_7591 (I131993,I131976,I95932);
nor I_7592 (I132010,I95944,I95941);
nand I_7593 (I132027,I132010,I131993);
nand I_7594 (I132044,I132027,I131894);
not I_7595 (I131767,I132044);
nand I_7596 (I132075,I95932,I95941);
nor I_7597 (I131734,I132075,I131843);
not I_7598 (I132106,I132075);
nand I_7599 (I132123,I132106,I131843);
not I_7600 (I131740,I132123);
nor I_7601 (I131743,I131877,I132123);
nor I_7602 (I132168,I131826,I132106);
nor I_7603 (I132185,I132075,I95938);
not I_7604 (I132202,I132185);
nor I_7605 (I131749,I132202,I131911);
nand I_7606 (I131737,I132202,I132123);
nand I_7607 (I132247,I132202,I131928);
nand I_7608 (I132264,I132106,I132247);
nor I_7609 (I131752,I132027,I132264);
nand I_7610 (I131764,I131809,I132202);
nand I_7611 (I131761,I132202,I132027);
nor I_7612 (I132323,I132168,I132185);
nor I_7613 (I131746,I132044,I132323);
and I_7614 (I131758,I132027,I132075);
not I_7615 (I132404,I2905);
or I_7616 (I132421,I80839,I80842);
nand I_7617 (I132438,I80851,I80857);
not I_7618 (I132455,I132438);
and I_7619 (I132472,I132455,I132421);
or I_7620 (I132489,I80863,I80848);
nor I_7621 (I132506,I132489,I80860);
not I_7622 (I132523,I132506);
nor I_7623 (I132540,I132438,I132523);
nand I_7624 (I132557,I132506,I132455);
nor I_7625 (I132574,I132506,I132455);
DFFARX1 I_7626 (I132574,I2898,I132404,I132384,);
nor I_7627 (I132605,I80839,I80854);
or I_7628 (I132622,I132605,I80836);
nor I_7629 (I132639,I80848,I80845);
nand I_7630 (I132656,I132639,I132622);
nand I_7631 (I132673,I132656,I132523);
not I_7632 (I132396,I132673);
nand I_7633 (I132704,I80836,I80845);
nor I_7634 (I132363,I132704,I132472);
not I_7635 (I132735,I132704);
nand I_7636 (I132752,I132735,I132472);
not I_7637 (I132369,I132752);
nor I_7638 (I132372,I132506,I132752);
nor I_7639 (I132797,I132455,I132735);
nor I_7640 (I132814,I132704,I80842);
not I_7641 (I132831,I132814);
nor I_7642 (I132378,I132831,I132540);
nand I_7643 (I132366,I132831,I132752);
nand I_7644 (I132876,I132831,I132557);
nand I_7645 (I132893,I132735,I132876);
nor I_7646 (I132381,I132656,I132893);
nand I_7647 (I132393,I132438,I132831);
nand I_7648 (I132390,I132831,I132656);
nor I_7649 (I132952,I132797,I132814);
nor I_7650 (I132375,I132673,I132952);
and I_7651 (I132387,I132656,I132704);
not I_7652 (I133033,I2905);
or I_7653 (I133050,I157243,I157261);
nand I_7654 (I133067,I157264,I157258);
not I_7655 (I133084,I133067);
and I_7656 (I133101,I133084,I133050);
or I_7657 (I133118,I157252,I157234);
nor I_7658 (I133135,I133118,I157240);
not I_7659 (I133152,I133135);
nor I_7660 (I133169,I133067,I133152);
nand I_7661 (I133186,I133135,I133084);
nor I_7662 (I133203,I133135,I133084);
DFFARX1 I_7663 (I133203,I2898,I133033,I133013,);
nor I_7664 (I133234,I157246,I157267);
or I_7665 (I133251,I133234,I157237);
nor I_7666 (I133268,I157249,I157240);
nand I_7667 (I133285,I133268,I133251);
nand I_7668 (I133302,I133285,I133152);
not I_7669 (I133025,I133302);
nand I_7670 (I133333,I157255,I157237);
nor I_7671 (I132992,I133333,I133101);
not I_7672 (I133364,I133333);
nand I_7673 (I133381,I133364,I133101);
not I_7674 (I132998,I133381);
nor I_7675 (I133001,I133135,I133381);
nor I_7676 (I133426,I133084,I133364);
nor I_7677 (I133443,I133333,I157234);
not I_7678 (I133460,I133443);
nor I_7679 (I133007,I133460,I133169);
nand I_7680 (I132995,I133460,I133381);
nand I_7681 (I133505,I133460,I133186);
nand I_7682 (I133522,I133364,I133505);
nor I_7683 (I133010,I133285,I133522);
nand I_7684 (I133022,I133067,I133460);
nand I_7685 (I133019,I133460,I133285);
nor I_7686 (I133581,I133426,I133443);
nor I_7687 (I133004,I133302,I133581);
and I_7688 (I133016,I133285,I133333);
not I_7689 (I133662,I2905);
or I_7690 (I133679,I246708,I246723);
nand I_7691 (I133696,I246729,I246711);
not I_7692 (I133713,I133696);
and I_7693 (I133730,I133713,I133679);
or I_7694 (I133747,I246714,I246726);
nor I_7695 (I133764,I133747,I246708);
not I_7696 (I133781,I133764);
nor I_7697 (I133798,I133696,I133781);
nand I_7698 (I133815,I133764,I133713);
nor I_7699 (I133832,I133764,I133713);
DFFARX1 I_7700 (I133832,I2898,I133662,I133642,);
nor I_7701 (I133863,I246717,I246705);
or I_7702 (I133880,I133863,I246705);
nor I_7703 (I133897,I246732,I246735);
nand I_7704 (I133914,I133897,I133880);
nand I_7705 (I133931,I133914,I133781);
not I_7706 (I133654,I133931);
nand I_7707 (I133962,I246720,I246711);
nor I_7708 (I133621,I133962,I133730);
not I_7709 (I133993,I133962);
nand I_7710 (I134010,I133993,I133730);
not I_7711 (I133627,I134010);
nor I_7712 (I133630,I133764,I134010);
nor I_7713 (I134055,I133713,I133993);
nor I_7714 (I134072,I133962,I246714);
not I_7715 (I134089,I134072);
nor I_7716 (I133636,I134089,I133798);
nand I_7717 (I133624,I134089,I134010);
nand I_7718 (I134134,I134089,I133815);
nand I_7719 (I134151,I133993,I134134);
nor I_7720 (I133639,I133914,I134151);
nand I_7721 (I133651,I133696,I134089);
nand I_7722 (I133648,I134089,I133914);
nor I_7723 (I134210,I134055,I134072);
nor I_7724 (I133633,I133931,I134210);
and I_7725 (I133645,I133914,I133962);
not I_7726 (I134291,I2905);
or I_7727 (I134308,I409469,I409478);
nand I_7728 (I134325,I409472,I409487);
not I_7729 (I134342,I134325);
and I_7730 (I134359,I134342,I134308);
or I_7731 (I134376,I409484,I409469);
nor I_7732 (I134393,I134376,I409463);
not I_7733 (I134410,I134393);
nor I_7734 (I134427,I134325,I134410);
nand I_7735 (I134444,I134393,I134342);
nor I_7736 (I134461,I134393,I134342);
DFFARX1 I_7737 (I134461,I2898,I134291,I134271,);
nor I_7738 (I134492,I409466,I409478);
or I_7739 (I134509,I134492,I409463);
nor I_7740 (I134526,I409475,I409466);
nand I_7741 (I134543,I134526,I134509);
nand I_7742 (I134560,I134543,I134410);
not I_7743 (I134283,I134560);
nand I_7744 (I134591,I409472,I409481);
nor I_7745 (I134250,I134591,I134359);
not I_7746 (I134622,I134591);
nand I_7747 (I134639,I134622,I134359);
not I_7748 (I134256,I134639);
nor I_7749 (I134259,I134393,I134639);
nor I_7750 (I134684,I134342,I134622);
nor I_7751 (I134701,I134591,I409475);
not I_7752 (I134718,I134701);
nor I_7753 (I134265,I134718,I134427);
nand I_7754 (I134253,I134718,I134639);
nand I_7755 (I134763,I134718,I134444);
nand I_7756 (I134780,I134622,I134763);
nor I_7757 (I134268,I134543,I134780);
nand I_7758 (I134280,I134325,I134718);
nand I_7759 (I134277,I134718,I134543);
nor I_7760 (I134839,I134684,I134701);
nor I_7761 (I134262,I134560,I134839);
and I_7762 (I134274,I134543,I134591);
not I_7763 (I134920,I2905);
or I_7764 (I134937,I283428,I283443);
nand I_7765 (I134954,I283449,I283431);
not I_7766 (I134971,I134954);
and I_7767 (I134988,I134971,I134937);
or I_7768 (I135005,I283434,I283446);
nor I_7769 (I135022,I135005,I283428);
not I_7770 (I135039,I135022);
nor I_7771 (I135056,I134954,I135039);
nand I_7772 (I135073,I135022,I134971);
nor I_7773 (I135090,I135022,I134971);
DFFARX1 I_7774 (I135090,I2898,I134920,I134900,);
nor I_7775 (I135121,I283437,I283425);
or I_7776 (I135138,I135121,I283425);
nor I_7777 (I135155,I283452,I283455);
nand I_7778 (I135172,I135155,I135138);
nand I_7779 (I135189,I135172,I135039);
not I_7780 (I134912,I135189);
nand I_7781 (I135220,I283440,I283431);
nor I_7782 (I134879,I135220,I134988);
not I_7783 (I135251,I135220);
nand I_7784 (I135268,I135251,I134988);
not I_7785 (I134885,I135268);
nor I_7786 (I134888,I135022,I135268);
nor I_7787 (I135313,I134971,I135251);
nor I_7788 (I135330,I135220,I283434);
not I_7789 (I135347,I135330);
nor I_7790 (I134894,I135347,I135056);
nand I_7791 (I134882,I135347,I135268);
nand I_7792 (I135392,I135347,I135073);
nand I_7793 (I135409,I135251,I135392);
nor I_7794 (I134897,I135172,I135409);
nand I_7795 (I134909,I134954,I135347);
nand I_7796 (I134906,I135347,I135172);
nor I_7797 (I135468,I135313,I135330);
nor I_7798 (I134891,I135189,I135468);
and I_7799 (I134903,I135172,I135220);
not I_7800 (I135549,I2905);
or I_7801 (I135566,I72662,I72665);
nand I_7802 (I135583,I72674,I72680);
not I_7803 (I135600,I135583);
and I_7804 (I135617,I135600,I135566);
or I_7805 (I135634,I72686,I72671);
nor I_7806 (I135651,I135634,I72683);
not I_7807 (I135668,I135651);
nor I_7808 (I135685,I135583,I135668);
nand I_7809 (I135702,I135651,I135600);
nor I_7810 (I135719,I135651,I135600);
DFFARX1 I_7811 (I135719,I2898,I135549,I135529,);
nor I_7812 (I135750,I72662,I72677);
or I_7813 (I135767,I135750,I72659);
nor I_7814 (I135784,I72671,I72668);
nand I_7815 (I135801,I135784,I135767);
nand I_7816 (I135818,I135801,I135668);
not I_7817 (I135541,I135818);
nand I_7818 (I135849,I72659,I72668);
nor I_7819 (I135508,I135849,I135617);
not I_7820 (I135880,I135849);
nand I_7821 (I135897,I135880,I135617);
not I_7822 (I135514,I135897);
nor I_7823 (I135517,I135651,I135897);
nor I_7824 (I135942,I135600,I135880);
nor I_7825 (I135959,I135849,I72665);
not I_7826 (I135976,I135959);
nor I_7827 (I135523,I135976,I135685);
nand I_7828 (I135511,I135976,I135897);
nand I_7829 (I136021,I135976,I135702);
nand I_7830 (I136038,I135880,I136021);
nor I_7831 (I135526,I135801,I136038);
nand I_7832 (I135538,I135583,I135976);
nand I_7833 (I135535,I135976,I135801);
nor I_7834 (I136097,I135942,I135959);
nor I_7835 (I135520,I135818,I136097);
and I_7836 (I135532,I135801,I135849);
not I_7837 (I136178,I2905);
or I_7838 (I136195,I237528,I237543);
nand I_7839 (I136212,I237549,I237531);
not I_7840 (I136229,I136212);
and I_7841 (I136246,I136229,I136195);
or I_7842 (I136263,I237534,I237546);
nor I_7843 (I136280,I136263,I237528);
not I_7844 (I136297,I136280);
nor I_7845 (I136314,I136212,I136297);
nand I_7846 (I136331,I136280,I136229);
nor I_7847 (I136348,I136280,I136229);
DFFARX1 I_7848 (I136348,I2898,I136178,I136158,);
nor I_7849 (I136379,I237537,I237525);
or I_7850 (I136396,I136379,I237525);
nor I_7851 (I136413,I237552,I237555);
nand I_7852 (I136430,I136413,I136396);
nand I_7853 (I136447,I136430,I136297);
not I_7854 (I136170,I136447);
nand I_7855 (I136478,I237540,I237531);
nor I_7856 (I136137,I136478,I136246);
not I_7857 (I136509,I136478);
nand I_7858 (I136526,I136509,I136246);
not I_7859 (I136143,I136526);
nor I_7860 (I136146,I136280,I136526);
nor I_7861 (I136571,I136229,I136509);
nor I_7862 (I136588,I136478,I237534);
not I_7863 (I136605,I136588);
nor I_7864 (I136152,I136605,I136314);
nand I_7865 (I136140,I136605,I136526);
nand I_7866 (I136650,I136605,I136331);
nand I_7867 (I136667,I136509,I136650);
nor I_7868 (I136155,I136430,I136667);
nand I_7869 (I136167,I136212,I136605);
nand I_7870 (I136164,I136605,I136430);
nor I_7871 (I136726,I136571,I136588);
nor I_7872 (I136149,I136447,I136726);
and I_7873 (I136161,I136430,I136478);
not I_7874 (I136807,I2905);
or I_7875 (I136824,I36781,I36778);
nand I_7876 (I136841,I36772,I36793);
not I_7877 (I136858,I136841);
and I_7878 (I136875,I136858,I136824);
or I_7879 (I136892,I36787,I36799);
nor I_7880 (I136909,I136892,I36781);
not I_7881 (I136926,I136909);
nor I_7882 (I136943,I136841,I136926);
nand I_7883 (I136960,I136909,I136858);
nor I_7884 (I136977,I136909,I136858);
DFFARX1 I_7885 (I136977,I2898,I136807,I136787,);
nor I_7886 (I137008,I36784,I36784);
or I_7887 (I137025,I137008,I36790);
nor I_7888 (I137042,I36775,I36778);
nand I_7889 (I137059,I137042,I137025);
nand I_7890 (I137076,I137059,I136926);
not I_7891 (I136799,I137076);
nand I_7892 (I137107,I36796,I36772);
nor I_7893 (I136766,I137107,I136875);
not I_7894 (I137138,I137107);
nand I_7895 (I137155,I137138,I136875);
not I_7896 (I136772,I137155);
nor I_7897 (I136775,I136909,I137155);
nor I_7898 (I137200,I136858,I137138);
nor I_7899 (I137217,I137107,I36775);
not I_7900 (I137234,I137217);
nor I_7901 (I136781,I137234,I136943);
nand I_7902 (I136769,I137234,I137155);
nand I_7903 (I137279,I137234,I136960);
nand I_7904 (I137296,I137138,I137279);
nor I_7905 (I136784,I137059,I137296);
nand I_7906 (I136796,I136841,I137234);
nand I_7907 (I136793,I137234,I137059);
nor I_7908 (I137355,I137200,I137217);
nor I_7909 (I136778,I137076,I137355);
and I_7910 (I136790,I137059,I137107);
not I_7911 (I137436,I2905);
or I_7912 (I137453,I18217,I18214);
nand I_7913 (I137470,I18208,I18229);
not I_7914 (I137487,I137470);
and I_7915 (I137504,I137487,I137453);
or I_7916 (I137521,I18223,I18235);
nor I_7917 (I137538,I137521,I18217);
not I_7918 (I137555,I137538);
nor I_7919 (I137572,I137470,I137555);
nand I_7920 (I137589,I137538,I137487);
nor I_7921 (I137606,I137538,I137487);
DFFARX1 I_7922 (I137606,I2898,I137436,I137416,);
nor I_7923 (I137637,I18220,I18220);
or I_7924 (I137654,I137637,I18226);
nor I_7925 (I137671,I18211,I18214);
nand I_7926 (I137688,I137671,I137654);
nand I_7927 (I137705,I137688,I137555);
not I_7928 (I137428,I137705);
nand I_7929 (I137736,I18232,I18208);
nor I_7930 (I137395,I137736,I137504);
not I_7931 (I137767,I137736);
nand I_7932 (I137784,I137767,I137504);
not I_7933 (I137401,I137784);
nor I_7934 (I137404,I137538,I137784);
nor I_7935 (I137829,I137487,I137767);
nor I_7936 (I137846,I137736,I18211);
not I_7937 (I137863,I137846);
nor I_7938 (I137410,I137863,I137572);
nand I_7939 (I137398,I137863,I137784);
nand I_7940 (I137908,I137863,I137589);
nand I_7941 (I137925,I137767,I137908);
nor I_7942 (I137413,I137688,I137925);
nand I_7943 (I137425,I137470,I137863);
nand I_7944 (I137422,I137863,I137688);
nor I_7945 (I137984,I137829,I137846);
nor I_7946 (I137407,I137705,I137984);
and I_7947 (I137419,I137688,I137736);
not I_7948 (I138065,I2905);
or I_7949 (I138082,I211198,I211213);
nand I_7950 (I138099,I211207,I211210);
not I_7951 (I138116,I138099);
and I_7952 (I138133,I138116,I138082);
or I_7953 (I138150,I211195,I211204);
nor I_7954 (I138167,I138150,I211195);
not I_7955 (I138184,I138167);
nor I_7956 (I138201,I138099,I138184);
nand I_7957 (I138218,I138167,I138116);
nor I_7958 (I138235,I138167,I138116);
DFFARX1 I_7959 (I138235,I2898,I138065,I138045,);
nor I_7960 (I138266,I211198,I211192);
or I_7961 (I138283,I138266,I211204);
nor I_7962 (I138300,I211201,I211219);
nand I_7963 (I138317,I138300,I138283);
nand I_7964 (I138334,I138317,I138184);
not I_7965 (I138057,I138334);
nand I_7966 (I138365,I211216,I211201);
nor I_7967 (I138024,I138365,I138133);
not I_7968 (I138396,I138365);
nand I_7969 (I138413,I138396,I138133);
not I_7970 (I138030,I138413);
nor I_7971 (I138033,I138167,I138413);
nor I_7972 (I138458,I138116,I138396);
nor I_7973 (I138475,I138365,I211192);
not I_7974 (I138492,I138475);
nor I_7975 (I138039,I138492,I138201);
nand I_7976 (I138027,I138492,I138413);
nand I_7977 (I138537,I138492,I138218);
nand I_7978 (I138554,I138396,I138537);
nor I_7979 (I138042,I138317,I138554);
nand I_7980 (I138054,I138099,I138492);
nand I_7981 (I138051,I138492,I138317);
nor I_7982 (I138613,I138458,I138475);
nor I_7983 (I138036,I138334,I138613);
and I_7984 (I138048,I138317,I138365);
not I_7985 (I138694,I2905);
or I_7986 (I138711,I84613,I84616);
nand I_7987 (I138728,I84625,I84631);
not I_7988 (I138745,I138728);
and I_7989 (I138762,I138745,I138711);
or I_7990 (I138779,I84637,I84622);
nor I_7991 (I138796,I138779,I84634);
not I_7992 (I138813,I138796);
nor I_7993 (I138830,I138728,I138813);
nand I_7994 (I138847,I138796,I138745);
nor I_7995 (I138864,I138796,I138745);
DFFARX1 I_7996 (I138864,I2898,I138694,I138674,);
nor I_7997 (I138895,I84613,I84628);
or I_7998 (I138912,I138895,I84610);
nor I_7999 (I138929,I84622,I84619);
nand I_8000 (I138946,I138929,I138912);
nand I_8001 (I138963,I138946,I138813);
not I_8002 (I138686,I138963);
nand I_8003 (I138994,I84610,I84619);
nor I_8004 (I138653,I138994,I138762);
not I_8005 (I139025,I138994);
nand I_8006 (I139042,I139025,I138762);
not I_8007 (I138659,I139042);
nor I_8008 (I138662,I138796,I139042);
nor I_8009 (I139087,I138745,I139025);
nor I_8010 (I139104,I138994,I84616);
not I_8011 (I139121,I139104);
nor I_8012 (I138668,I139121,I138830);
nand I_8013 (I138656,I139121,I139042);
nand I_8014 (I139166,I139121,I138847);
nand I_8015 (I139183,I139025,I139166);
nor I_8016 (I138671,I138946,I139183);
nand I_8017 (I138683,I138728,I139121);
nand I_8018 (I138680,I139121,I138946);
nor I_8019 (I139242,I139087,I139104);
nor I_8020 (I138665,I138963,I139242);
and I_8021 (I138677,I138946,I138994);
not I_8022 (I139323,I2905);
or I_8023 (I139340,I259713,I259728);
nand I_8024 (I139357,I259734,I259716);
not I_8025 (I139374,I139357);
and I_8026 (I139391,I139374,I139340);
or I_8027 (I139408,I259719,I259731);
nor I_8028 (I139425,I139408,I259713);
not I_8029 (I139442,I139425);
nor I_8030 (I139459,I139357,I139442);
nand I_8031 (I139476,I139425,I139374);
nor I_8032 (I139493,I139425,I139374);
DFFARX1 I_8033 (I139493,I2898,I139323,I139303,);
nor I_8034 (I139524,I259722,I259710);
or I_8035 (I139541,I139524,I259710);
nor I_8036 (I139558,I259737,I259740);
nand I_8037 (I139575,I139558,I139541);
nand I_8038 (I139592,I139575,I139442);
not I_8039 (I139315,I139592);
nand I_8040 (I139623,I259725,I259716);
nor I_8041 (I139282,I139623,I139391);
not I_8042 (I139654,I139623);
nand I_8043 (I139671,I139654,I139391);
not I_8044 (I139288,I139671);
nor I_8045 (I139291,I139425,I139671);
nor I_8046 (I139716,I139374,I139654);
nor I_8047 (I139733,I139623,I259719);
not I_8048 (I139750,I139733);
nor I_8049 (I139297,I139750,I139459);
nand I_8050 (I139285,I139750,I139671);
nand I_8051 (I139795,I139750,I139476);
nand I_8052 (I139812,I139654,I139795);
nor I_8053 (I139300,I139575,I139812);
nand I_8054 (I139312,I139357,I139750);
nand I_8055 (I139309,I139750,I139575);
nor I_8056 (I139871,I139716,I139733);
nor I_8057 (I139294,I139592,I139871);
and I_8058 (I139306,I139575,I139623);
not I_8059 (I139952,I2905);
or I_8060 (I139969,I242118,I242133);
nand I_8061 (I139986,I242139,I242121);
not I_8062 (I140003,I139986);
and I_8063 (I140020,I140003,I139969);
or I_8064 (I140037,I242124,I242136);
nor I_8065 (I140054,I140037,I242118);
not I_8066 (I140071,I140054);
nor I_8067 (I140088,I139986,I140071);
nand I_8068 (I140105,I140054,I140003);
nor I_8069 (I140122,I140054,I140003);
DFFARX1 I_8070 (I140122,I2898,I139952,I139932,);
nor I_8071 (I140153,I242127,I242115);
or I_8072 (I140170,I140153,I242115);
nor I_8073 (I140187,I242142,I242145);
nand I_8074 (I140204,I140187,I140170);
nand I_8075 (I140221,I140204,I140071);
not I_8076 (I139944,I140221);
nand I_8077 (I140252,I242130,I242121);
nor I_8078 (I139911,I140252,I140020);
not I_8079 (I140283,I140252);
nand I_8080 (I140300,I140283,I140020);
not I_8081 (I139917,I140300);
nor I_8082 (I139920,I140054,I140300);
nor I_8083 (I140345,I140003,I140283);
nor I_8084 (I140362,I140252,I242124);
not I_8085 (I140379,I140362);
nor I_8086 (I139926,I140379,I140088);
nand I_8087 (I139914,I140379,I140300);
nand I_8088 (I140424,I140379,I140105);
nand I_8089 (I140441,I140283,I140424);
nor I_8090 (I139929,I140204,I140441);
nand I_8091 (I139941,I139986,I140379);
nand I_8092 (I139938,I140379,I140204);
nor I_8093 (I140500,I140345,I140362);
nor I_8094 (I139923,I140221,I140500);
and I_8095 (I139935,I140204,I140252);
not I_8096 (I140581,I2905);
or I_8097 (I140598,I4756,I4765);
nand I_8098 (I140615,I4774,I4762);
not I_8099 (I140632,I140615);
and I_8100 (I140649,I140632,I140598);
or I_8101 (I140666,I4759,I4747);
nor I_8102 (I140683,I140666,I4744);
not I_8103 (I140700,I140683);
nor I_8104 (I140717,I140615,I140700);
nand I_8105 (I140734,I140683,I140632);
nor I_8106 (I140751,I140683,I140632);
DFFARX1 I_8107 (I140751,I2898,I140581,I140561,);
nor I_8108 (I140782,I4768,I4747);
or I_8109 (I140799,I140782,I4750);
nor I_8110 (I140816,I4744,I4753);
nand I_8111 (I140833,I140816,I140799);
nand I_8112 (I140850,I140833,I140700);
not I_8113 (I140573,I140850);
nand I_8114 (I140881,I4753,I4750);
nor I_8115 (I140540,I140881,I140649);
not I_8116 (I140912,I140881);
nand I_8117 (I140929,I140912,I140649);
not I_8118 (I140546,I140929);
nor I_8119 (I140549,I140683,I140929);
nor I_8120 (I140974,I140632,I140912);
nor I_8121 (I140991,I140881,I4771);
not I_8122 (I141008,I140991);
nor I_8123 (I140555,I141008,I140717);
nand I_8124 (I140543,I141008,I140929);
nand I_8125 (I141053,I141008,I140734);
nand I_8126 (I141070,I140912,I141053);
nor I_8127 (I140558,I140833,I141070);
nand I_8128 (I140570,I140615,I141008);
nand I_8129 (I140567,I141008,I140833);
nor I_8130 (I141129,I140974,I140991);
nor I_8131 (I140552,I140850,I141129);
and I_8132 (I140564,I140833,I140881);
not I_8133 (I141210,I2905);
or I_8134 (I141227,I89645,I89648);
nand I_8135 (I141244,I89657,I89663);
not I_8136 (I141261,I141244);
and I_8137 (I141278,I141261,I141227);
or I_8138 (I141295,I89669,I89654);
nor I_8139 (I141312,I141295,I89666);
not I_8140 (I141329,I141312);
nor I_8141 (I141346,I141244,I141329);
nand I_8142 (I141363,I141312,I141261);
nor I_8143 (I141380,I141312,I141261);
DFFARX1 I_8144 (I141380,I2898,I141210,I141190,);
nor I_8145 (I141411,I89645,I89660);
or I_8146 (I141428,I141411,I89642);
nor I_8147 (I141445,I89654,I89651);
nand I_8148 (I141462,I141445,I141428);
nand I_8149 (I141479,I141462,I141329);
not I_8150 (I141202,I141479);
nand I_8151 (I141510,I89642,I89651);
nor I_8152 (I141169,I141510,I141278);
not I_8153 (I141541,I141510);
nand I_8154 (I141558,I141541,I141278);
not I_8155 (I141175,I141558);
nor I_8156 (I141178,I141312,I141558);
nor I_8157 (I141603,I141261,I141541);
nor I_8158 (I141620,I141510,I89648);
not I_8159 (I141637,I141620);
nor I_8160 (I141184,I141637,I141346);
nand I_8161 (I141172,I141637,I141558);
nand I_8162 (I141682,I141637,I141363);
nand I_8163 (I141699,I141541,I141682);
nor I_8164 (I141187,I141462,I141699);
nand I_8165 (I141199,I141244,I141637);
nand I_8166 (I141196,I141637,I141462);
nor I_8167 (I141758,I141603,I141620);
nor I_8168 (I141181,I141479,I141758);
and I_8169 (I141193,I141462,I141510);
not I_8170 (I141839,I2905);
or I_8171 (I141856,I406749,I406758);
nand I_8172 (I141873,I406752,I406767);
not I_8173 (I141890,I141873);
and I_8174 (I141907,I141890,I141856);
or I_8175 (I141924,I406764,I406749);
nor I_8176 (I141941,I141924,I406743);
not I_8177 (I141958,I141941);
nor I_8178 (I141975,I141873,I141958);
nand I_8179 (I141992,I141941,I141890);
nor I_8180 (I142009,I141941,I141890);
DFFARX1 I_8181 (I142009,I2898,I141839,I141819,);
nor I_8182 (I142040,I406746,I406758);
or I_8183 (I142057,I142040,I406743);
nor I_8184 (I142074,I406755,I406746);
nand I_8185 (I142091,I142074,I142057);
nand I_8186 (I142108,I142091,I141958);
not I_8187 (I141831,I142108);
nand I_8188 (I142139,I406752,I406761);
nor I_8189 (I141798,I142139,I141907);
not I_8190 (I142170,I142139);
nand I_8191 (I142187,I142170,I141907);
not I_8192 (I141804,I142187);
nor I_8193 (I141807,I141941,I142187);
nor I_8194 (I142232,I141890,I142170);
nor I_8195 (I142249,I142139,I406755);
not I_8196 (I142266,I142249);
nor I_8197 (I141813,I142266,I141975);
nand I_8198 (I141801,I142266,I142187);
nand I_8199 (I142311,I142266,I141992);
nand I_8200 (I142328,I142170,I142311);
nor I_8201 (I141816,I142091,I142328);
nand I_8202 (I141828,I141873,I142266);
nand I_8203 (I141825,I142266,I142091);
nor I_8204 (I142387,I142232,I142249);
nor I_8205 (I141810,I142108,I142387);
and I_8206 (I141822,I142091,I142139);
not I_8207 (I142468,I2905);
or I_8208 (I142485,I428275,I428248);
nand I_8209 (I142502,I428278,I428257);
not I_8210 (I142519,I142502);
and I_8211 (I142536,I142519,I142485);
or I_8212 (I142553,I428266,I428251);
nor I_8213 (I142570,I142553,I428269);
not I_8214 (I142587,I142570);
nor I_8215 (I142604,I142502,I142587);
nand I_8216 (I142621,I142570,I142519);
nor I_8217 (I142638,I142570,I142519);
DFFARX1 I_8218 (I142638,I2898,I142468,I142448,);
nor I_8219 (I142669,I428272,I428251);
or I_8220 (I142686,I142669,I428254);
nor I_8221 (I142703,I428260,I428248);
nand I_8222 (I142720,I142703,I142686);
nand I_8223 (I142737,I142720,I142587);
not I_8224 (I142460,I142737);
nand I_8225 (I142768,I428254,I428263);
nor I_8226 (I142427,I142768,I142536);
not I_8227 (I142799,I142768);
nand I_8228 (I142816,I142799,I142536);
not I_8229 (I142433,I142816);
nor I_8230 (I142436,I142570,I142816);
nor I_8231 (I142861,I142519,I142799);
nor I_8232 (I142878,I142768,I428281);
not I_8233 (I142895,I142878);
nor I_8234 (I142442,I142895,I142604);
nand I_8235 (I142430,I142895,I142816);
nand I_8236 (I142940,I142895,I142621);
nand I_8237 (I142957,I142799,I142940);
nor I_8238 (I142445,I142720,I142957);
nand I_8239 (I142457,I142502,I142895);
nand I_8240 (I142454,I142895,I142720);
nor I_8241 (I143016,I142861,I142878);
nor I_8242 (I142439,I142737,I143016);
and I_8243 (I142451,I142720,I142768);
not I_8244 (I143097,I2905);
or I_8245 (I143114,I24643,I24640);
nand I_8246 (I143131,I24634,I24655);
not I_8247 (I143148,I143131);
and I_8248 (I143165,I143148,I143114);
or I_8249 (I143182,I24649,I24661);
nor I_8250 (I143199,I143182,I24643);
not I_8251 (I143216,I143199);
nor I_8252 (I143233,I143131,I143216);
nand I_8253 (I143250,I143199,I143148);
nor I_8254 (I143267,I143199,I143148);
DFFARX1 I_8255 (I143267,I2898,I143097,I143077,);
nor I_8256 (I143298,I24646,I24646);
or I_8257 (I143315,I143298,I24652);
nor I_8258 (I143332,I24637,I24640);
nand I_8259 (I143349,I143332,I143315);
nand I_8260 (I143366,I143349,I143216);
not I_8261 (I143089,I143366);
nand I_8262 (I143397,I24658,I24634);
nor I_8263 (I143056,I143397,I143165);
not I_8264 (I143428,I143397);
nand I_8265 (I143445,I143428,I143165);
not I_8266 (I143062,I143445);
nor I_8267 (I143065,I143199,I143445);
nor I_8268 (I143490,I143148,I143428);
nor I_8269 (I143507,I143397,I24637);
not I_8270 (I143524,I143507);
nor I_8271 (I143071,I143524,I143233);
nand I_8272 (I143059,I143524,I143445);
nand I_8273 (I143569,I143524,I143250);
nand I_8274 (I143586,I143428,I143569);
nor I_8275 (I143074,I143349,I143586);
nand I_8276 (I143086,I143131,I143524);
nand I_8277 (I143083,I143524,I143349);
nor I_8278 (I143645,I143490,I143507);
nor I_8279 (I143068,I143366,I143645);
and I_8280 (I143080,I143349,I143397);
not I_8281 (I143726,I2905);
or I_8282 (I143743,I385520,I385496);
nand I_8283 (I143760,I385526,I385508);
not I_8284 (I143777,I143760);
and I_8285 (I143794,I143777,I143743);
or I_8286 (I143811,I385514,I385523);
nor I_8287 (I143828,I143811,I385499);
not I_8288 (I143845,I143828);
nor I_8289 (I143862,I143760,I143845);
nand I_8290 (I143879,I143828,I143777);
nor I_8291 (I143896,I143828,I143777);
DFFARX1 I_8292 (I143896,I2898,I143726,I143706,);
nor I_8293 (I143927,I385499,I385505);
or I_8294 (I143944,I143927,I385496);
nor I_8295 (I143961,I385493,I385493);
nand I_8296 (I143978,I143961,I143944);
nand I_8297 (I143995,I143978,I143845);
not I_8298 (I143718,I143995);
nand I_8299 (I144026,I385511,I385517);
nor I_8300 (I143685,I144026,I143794);
not I_8301 (I144057,I144026);
nand I_8302 (I144074,I144057,I143794);
not I_8303 (I143691,I144074);
nor I_8304 (I143694,I143828,I144074);
nor I_8305 (I144119,I143777,I144057);
nor I_8306 (I144136,I144026,I385502);
not I_8307 (I144153,I144136);
nor I_8308 (I143700,I144153,I143862);
nand I_8309 (I143688,I144153,I144074);
nand I_8310 (I144198,I144153,I143879);
nand I_8311 (I144215,I144057,I144198);
nor I_8312 (I143703,I143978,I144215);
nand I_8313 (I143715,I143760,I144153);
nand I_8314 (I143712,I144153,I143978);
nor I_8315 (I144274,I144119,I144136);
nor I_8316 (I143697,I143995,I144274);
and I_8317 (I143709,I143978,I144026);
not I_8318 (I144355,I2905);
or I_8319 (I144372,I323426,I323435);
nor I_8320 (I144389,I323426,I323435);
nor I_8321 (I144406,I144389,I323441);
nand I_8322 (I144423,I144372,I323447);
not I_8323 (I144440,I144423);
not I_8324 (I144457,I323429);
nor I_8325 (I144314,I144406,I144457);
nand I_8326 (I144488,I144406,I323429);
not I_8327 (I144344,I144488);
not I_8328 (I144519,I323438);
nand I_8329 (I144536,I323435,I323444);
nand I_8330 (I144553,I144536,I323438);
not I_8331 (I144570,I144553);
nand I_8332 (I144587,I144406,I144570);
not I_8333 (I144320,I144587);
nor I_8334 (I144332,I144406,I144570);
nor I_8335 (I144632,I144553,I323429);
DFFARX1 I_8336 (I144632,I2898,I144355,I144335,);
nand I_8337 (I144663,I144536,I144519);
and I_8338 (I144680,I144663,I323432);
nand I_8339 (I144697,I144680,I323429);
nor I_8340 (I144714,I144697,I144553);
not I_8341 (I144731,I144697);
nor I_8342 (I144748,I144440,I144731);
nor I_8343 (I144338,I144748,I144457);
nor I_8344 (I144341,I144440,I144697);
nor I_8345 (I144793,I323432,I323450);
or I_8346 (I144810,I144793,I323438);
nor I_8347 (I144827,I323441,I323426);
and I_8348 (I144844,I144827,I144810);
nor I_8349 (I144861,I144844,I144714);
nor I_8350 (I144326,I144861,I144714);
or I_8351 (I144892,I144697,I144861);
nor I_8352 (I144329,I144423,I144892);
nor I_8353 (I144923,I144570,I144844);
nor I_8354 (I144317,I144457,I144923);
nor I_8355 (I144954,I144731,I144844);
nor I_8356 (I144347,I144954,I144488);
nor I_8357 (I144323,I144844,I144587);
not I_8358 (I145035,I2905);
or I_8359 (I145052,I235248,I235251);
nor I_8360 (I145069,I235248,I235251);
nor I_8361 (I145086,I145069,I235233);
nand I_8362 (I145103,I145052,I235260);
not I_8363 (I145120,I145103);
not I_8364 (I145137,I235245);
nor I_8365 (I144994,I145086,I145137);
nand I_8366 (I145168,I145086,I235245);
not I_8367 (I145024,I145168);
not I_8368 (I145199,I235257);
nand I_8369 (I145216,I235236,I235239);
nand I_8370 (I145233,I145216,I235257);
not I_8371 (I145250,I145233);
nand I_8372 (I145267,I145086,I145250);
not I_8373 (I145000,I145267);
nor I_8374 (I145012,I145086,I145250);
nor I_8375 (I145312,I145233,I235245);
DFFARX1 I_8376 (I145312,I2898,I145035,I145015,);
nand I_8377 (I145343,I145216,I145199);
and I_8378 (I145360,I145343,I235233);
nand I_8379 (I145377,I145360,I235242);
nor I_8380 (I145394,I145377,I145233);
not I_8381 (I145411,I145377);
nor I_8382 (I145428,I145120,I145411);
nor I_8383 (I145018,I145428,I145137);
nor I_8384 (I145021,I145120,I145377);
nor I_8385 (I145473,I235230,I235230);
or I_8386 (I145490,I145473,I235254);
nor I_8387 (I145507,I235236,I235239);
and I_8388 (I145524,I145507,I145490);
nor I_8389 (I145541,I145524,I145394);
nor I_8390 (I145006,I145541,I145394);
or I_8391 (I145572,I145377,I145541);
nor I_8392 (I145009,I145103,I145572);
nor I_8393 (I145603,I145250,I145524);
nor I_8394 (I144997,I145137,I145603);
nor I_8395 (I145634,I145411,I145524);
nor I_8396 (I145027,I145634,I145168);
nor I_8397 (I145003,I145524,I145267);
not I_8398 (I145715,I2905);
or I_8399 (I145732,I424066,I424084);
nor I_8400 (I145749,I424066,I424084);
nor I_8401 (I145766,I145749,I424099);
nand I_8402 (I145783,I145732,I424069);
not I_8403 (I145800,I145783);
not I_8404 (I145817,I424072);
nor I_8405 (I145674,I145766,I145817);
nand I_8406 (I145848,I145766,I424072);
not I_8407 (I145704,I145848);
not I_8408 (I145879,I424093);
nand I_8409 (I145896,I424081,I424096);
nand I_8410 (I145913,I145896,I424093);
not I_8411 (I145930,I145913);
nand I_8412 (I145947,I145766,I145930);
not I_8413 (I145680,I145947);
nor I_8414 (I145692,I145766,I145930);
nor I_8415 (I145992,I145913,I424072);
DFFARX1 I_8416 (I145992,I2898,I145715,I145695,);
nand I_8417 (I146023,I145896,I145879);
and I_8418 (I146040,I146023,I424087);
nand I_8419 (I146057,I146040,I424066);
nor I_8420 (I146074,I146057,I145913);
not I_8421 (I146091,I146057);
nor I_8422 (I146108,I145800,I146091);
nor I_8423 (I145698,I146108,I145817);
nor I_8424 (I145701,I145800,I146057);
nor I_8425 (I146153,I424072,I424069);
or I_8426 (I146170,I146153,I424075);
nor I_8427 (I146187,I424090,I424078);
and I_8428 (I146204,I146187,I146170);
nor I_8429 (I146221,I146204,I146074);
nor I_8430 (I145686,I146221,I146074);
or I_8431 (I146252,I146057,I146221);
nor I_8432 (I145689,I145783,I146252);
nor I_8433 (I146283,I145930,I146204);
nor I_8434 (I145677,I145817,I146283);
nor I_8435 (I146314,I146091,I146204);
nor I_8436 (I145707,I146314,I145848);
nor I_8437 (I145683,I146204,I145947);
not I_8438 (I146395,I2905);
or I_8439 (I146412,I141831,I141801);
nor I_8440 (I146429,I141831,I141801);
nor I_8441 (I146446,I146429,I141822);
nand I_8442 (I146463,I146412,I141804);
not I_8443 (I146480,I146463);
not I_8444 (I146497,I141810);
nor I_8445 (I146354,I146446,I146497);
nand I_8446 (I146528,I146446,I141810);
not I_8447 (I146384,I146528);
not I_8448 (I146559,I141816);
nand I_8449 (I146576,I141801,I141813);
nand I_8450 (I146593,I146576,I141816);
not I_8451 (I146610,I146593);
nand I_8452 (I146627,I146446,I146610);
not I_8453 (I146360,I146627);
nor I_8454 (I146372,I146446,I146610);
nor I_8455 (I146672,I146593,I141810);
DFFARX1 I_8456 (I146672,I2898,I146395,I146375,);
nand I_8457 (I146703,I146576,I146559);
and I_8458 (I146720,I146703,I141798);
nand I_8459 (I146737,I146720,I141828);
nor I_8460 (I146754,I146737,I146593);
not I_8461 (I146771,I146737);
nor I_8462 (I146788,I146480,I146771);
nor I_8463 (I146378,I146788,I146497);
nor I_8464 (I146381,I146480,I146737);
nor I_8465 (I146833,I141804,I141825);
or I_8466 (I146850,I146833,I141819);
nor I_8467 (I146867,I141798,I141807);
and I_8468 (I146884,I146867,I146850);
nor I_8469 (I146901,I146884,I146754);
nor I_8470 (I146366,I146901,I146754);
or I_8471 (I146932,I146737,I146901);
nor I_8472 (I146369,I146463,I146932);
nor I_8473 (I146963,I146610,I146884);
nor I_8474 (I146357,I146497,I146963);
nor I_8475 (I146994,I146771,I146884);
nor I_8476 (I146387,I146994,I146528);
nor I_8477 (I146363,I146884,I146627);
not I_8478 (I147075,I2905);
or I_8479 (I147092,I100317,I100287);
nor I_8480 (I147109,I100317,I100287);
nor I_8481 (I147126,I147109,I100308);
nand I_8482 (I147143,I147092,I100290);
not I_8483 (I147160,I147143);
not I_8484 (I147177,I100296);
nor I_8485 (I147034,I147126,I147177);
nand I_8486 (I147208,I147126,I100296);
not I_8487 (I147064,I147208);
not I_8488 (I147239,I100302);
nand I_8489 (I147256,I100287,I100299);
nand I_8490 (I147273,I147256,I100302);
not I_8491 (I147290,I147273);
nand I_8492 (I147307,I147126,I147290);
not I_8493 (I147040,I147307);
nor I_8494 (I147052,I147126,I147290);
nor I_8495 (I147352,I147273,I100296);
DFFARX1 I_8496 (I147352,I2898,I147075,I147055,);
nand I_8497 (I147383,I147256,I147239);
and I_8498 (I147400,I147383,I100284);
nand I_8499 (I147417,I147400,I100314);
nor I_8500 (I147434,I147417,I147273);
not I_8501 (I147451,I147417);
nor I_8502 (I147468,I147160,I147451);
nor I_8503 (I147058,I147468,I147177);
nor I_8504 (I147061,I147160,I147417);
nor I_8505 (I147513,I100290,I100311);
or I_8506 (I147530,I147513,I100305);
nor I_8507 (I147547,I100284,I100293);
and I_8508 (I147564,I147547,I147530);
nor I_8509 (I147581,I147564,I147434);
nor I_8510 (I147046,I147581,I147434);
or I_8511 (I147612,I147417,I147581);
nor I_8512 (I147049,I147143,I147612);
nor I_8513 (I147643,I147290,I147564);
nor I_8514 (I147037,I147177,I147643);
nor I_8515 (I147674,I147451,I147564);
nor I_8516 (I147067,I147674,I147208);
nor I_8517 (I147043,I147564,I147307);
not I_8518 (I147755,I2905);
or I_8519 (I147772,I441491,I441509);
nor I_8520 (I147789,I441491,I441509);
nor I_8521 (I147806,I147789,I441524);
nand I_8522 (I147823,I147772,I441494);
not I_8523 (I147840,I147823);
not I_8524 (I147857,I441497);
nor I_8525 (I147714,I147806,I147857);
nand I_8526 (I147888,I147806,I441497);
not I_8527 (I147744,I147888);
not I_8528 (I147919,I441518);
nand I_8529 (I147936,I441506,I441521);
nand I_8530 (I147953,I147936,I441518);
not I_8531 (I147970,I147953);
nand I_8532 (I147987,I147806,I147970);
not I_8533 (I147720,I147987);
nor I_8534 (I147732,I147806,I147970);
nor I_8535 (I148032,I147953,I441497);
DFFARX1 I_8536 (I148032,I2898,I147755,I147735,);
nand I_8537 (I148063,I147936,I147919);
and I_8538 (I148080,I148063,I441512);
nand I_8539 (I148097,I148080,I441491);
nor I_8540 (I148114,I148097,I147953);
not I_8541 (I148131,I148097);
nor I_8542 (I148148,I147840,I148131);
nor I_8543 (I147738,I148148,I147857);
nor I_8544 (I147741,I147840,I148097);
nor I_8545 (I148193,I441497,I441494);
or I_8546 (I148210,I148193,I441500);
nor I_8547 (I148227,I441515,I441503);
and I_8548 (I148244,I148227,I148210);
nor I_8549 (I148261,I148244,I148114);
nor I_8550 (I147726,I148261,I148114);
or I_8551 (I148292,I148097,I148261);
nor I_8552 (I147729,I147823,I148292);
nor I_8553 (I148323,I147970,I148244);
nor I_8554 (I147717,I147857,I148323);
nor I_8555 (I148354,I148131,I148244);
nor I_8556 (I147747,I148354,I147888);
nor I_8557 (I147723,I148244,I147987);
not I_8558 (I148435,I2905);
or I_8559 (I148452,I229165,I229144);
nor I_8560 (I148469,I229165,I229144);
nor I_8561 (I148486,I148469,I229147);
nand I_8562 (I148503,I148452,I229171);
not I_8563 (I148520,I148503);
not I_8564 (I148537,I229162);
nor I_8565 (I148394,I148486,I148537);
nand I_8566 (I148568,I148486,I229162);
not I_8567 (I148424,I148568);
not I_8568 (I148599,I229159);
nand I_8569 (I148616,I229153,I229144);
nand I_8570 (I148633,I148616,I229159);
not I_8571 (I148650,I148633);
nand I_8572 (I148667,I148486,I148650);
not I_8573 (I148400,I148667);
nor I_8574 (I148412,I148486,I148650);
nor I_8575 (I148712,I148633,I229162);
DFFARX1 I_8576 (I148712,I2898,I148435,I148415,);
nand I_8577 (I148743,I148616,I148599);
and I_8578 (I148760,I148743,I229156);
nand I_8579 (I148777,I148760,I229156);
nor I_8580 (I148794,I148777,I148633);
not I_8581 (I148811,I148777);
nor I_8582 (I148828,I148520,I148811);
nor I_8583 (I148418,I148828,I148537);
nor I_8584 (I148421,I148520,I148777);
nor I_8585 (I148873,I229150,I229153);
or I_8586 (I148890,I148873,I229147);
nor I_8587 (I148907,I229168,I229150);
and I_8588 (I148924,I148907,I148890);
nor I_8589 (I148941,I148924,I148794);
nor I_8590 (I148406,I148941,I148794);
or I_8591 (I148972,I148777,I148941);
nor I_8592 (I148409,I148503,I148972);
nor I_8593 (I149003,I148650,I148924);
nor I_8594 (I148397,I148537,I149003);
nor I_8595 (I149034,I148811,I148924);
nor I_8596 (I148427,I149034,I148568);
nor I_8597 (I148403,I148924,I148667);
not I_8598 (I149115,I2905);
or I_8599 (I149132,I278853,I278856);
nor I_8600 (I149149,I278853,I278856);
nor I_8601 (I149166,I149149,I278838);
nand I_8602 (I149183,I149132,I278865);
not I_8603 (I149200,I149183);
not I_8604 (I149217,I278850);
nor I_8605 (I149074,I149166,I149217);
nand I_8606 (I149248,I149166,I278850);
not I_8607 (I149104,I149248);
not I_8608 (I149279,I278862);
nand I_8609 (I149296,I278841,I278844);
nand I_8610 (I149313,I149296,I278862);
not I_8611 (I149330,I149313);
nand I_8612 (I149347,I149166,I149330);
not I_8613 (I149080,I149347);
nor I_8614 (I149092,I149166,I149330);
nor I_8615 (I149392,I149313,I278850);
DFFARX1 I_8616 (I149392,I2898,I149115,I149095,);
nand I_8617 (I149423,I149296,I149279);
and I_8618 (I149440,I149423,I278838);
nand I_8619 (I149457,I149440,I278847);
nor I_8620 (I149474,I149457,I149313);
not I_8621 (I149491,I149457);
nor I_8622 (I149508,I149200,I149491);
nor I_8623 (I149098,I149508,I149217);
nor I_8624 (I149101,I149200,I149457);
nor I_8625 (I149553,I278835,I278835);
or I_8626 (I149570,I149553,I278859);
nor I_8627 (I149587,I278841,I278844);
and I_8628 (I149604,I149587,I149570);
nor I_8629 (I149621,I149604,I149474);
nor I_8630 (I149086,I149621,I149474);
or I_8631 (I149652,I149457,I149621);
nor I_8632 (I149089,I149183,I149652);
nor I_8633 (I149683,I149330,I149604);
nor I_8634 (I149077,I149217,I149683);
nor I_8635 (I149714,I149491,I149604);
nor I_8636 (I149107,I149714,I149248);
nor I_8637 (I149083,I149604,I149347);
not I_8638 (I149795,I2905);
or I_8639 (I149812,I239838,I239841);
nor I_8640 (I149829,I239838,I239841);
nor I_8641 (I149846,I149829,I239823);
nand I_8642 (I149863,I149812,I239850);
not I_8643 (I149880,I149863);
not I_8644 (I149897,I239835);
nor I_8645 (I149754,I149846,I149897);
nand I_8646 (I149928,I149846,I239835);
not I_8647 (I149784,I149928);
not I_8648 (I149959,I239847);
nand I_8649 (I149976,I239826,I239829);
nand I_8650 (I149993,I149976,I239847);
not I_8651 (I150010,I149993);
nand I_8652 (I150027,I149846,I150010);
not I_8653 (I149760,I150027);
nor I_8654 (I149772,I149846,I150010);
nor I_8655 (I150072,I149993,I239835);
DFFARX1 I_8656 (I150072,I2898,I149795,I149775,);
nand I_8657 (I150103,I149976,I149959);
and I_8658 (I150120,I150103,I239823);
nand I_8659 (I150137,I150120,I239832);
nor I_8660 (I150154,I150137,I149993);
not I_8661 (I150171,I150137);
nor I_8662 (I150188,I149880,I150171);
nor I_8663 (I149778,I150188,I149897);
nor I_8664 (I149781,I149880,I150137);
nor I_8665 (I150233,I239820,I239820);
or I_8666 (I150250,I150233,I239844);
nor I_8667 (I150267,I239826,I239829);
and I_8668 (I150284,I150267,I150250);
nor I_8669 (I150301,I150284,I150154);
nor I_8670 (I149766,I150301,I150154);
or I_8671 (I150332,I150137,I150301);
nor I_8672 (I149769,I149863,I150332);
nor I_8673 (I150363,I150010,I150284);
nor I_8674 (I149757,I149897,I150363);
nor I_8675 (I150394,I150171,I150284);
nor I_8676 (I149787,I150394,I149928);
nor I_8677 (I149763,I150284,I150027);
not I_8678 (I150475,I2905);
or I_8679 (I150492,I268143,I268146);
nor I_8680 (I150509,I268143,I268146);
nor I_8681 (I150526,I150509,I268128);
nand I_8682 (I150543,I150492,I268155);
not I_8683 (I150560,I150543);
not I_8684 (I150577,I268140);
nor I_8685 (I150434,I150526,I150577);
nand I_8686 (I150608,I150526,I268140);
not I_8687 (I150464,I150608);
not I_8688 (I150639,I268152);
nand I_8689 (I150656,I268131,I268134);
nand I_8690 (I150673,I150656,I268152);
not I_8691 (I150690,I150673);
nand I_8692 (I150707,I150526,I150690);
not I_8693 (I150440,I150707);
nor I_8694 (I150452,I150526,I150690);
nor I_8695 (I150752,I150673,I268140);
DFFARX1 I_8696 (I150752,I2898,I150475,I150455,);
nand I_8697 (I150783,I150656,I150639);
and I_8698 (I150800,I150783,I268128);
nand I_8699 (I150817,I150800,I268137);
nor I_8700 (I150834,I150817,I150673);
not I_8701 (I150851,I150817);
nor I_8702 (I150868,I150560,I150851);
nor I_8703 (I150458,I150868,I150577);
nor I_8704 (I150461,I150560,I150817);
nor I_8705 (I150913,I268125,I268125);
or I_8706 (I150930,I150913,I268149);
nor I_8707 (I150947,I268131,I268134);
and I_8708 (I150964,I150947,I150930);
nor I_8709 (I150981,I150964,I150834);
nor I_8710 (I150446,I150981,I150834);
or I_8711 (I151012,I150817,I150981);
nor I_8712 (I150449,I150543,I151012);
nor I_8713 (I151043,I150690,I150964);
nor I_8714 (I150437,I150577,I151043);
nor I_8715 (I151074,I150851,I150964);
nor I_8716 (I150467,I151074,I150608);
nor I_8717 (I150443,I150964,I150707);
not I_8718 (I151155,I2905);
or I_8719 (I151172,I353176,I353185);
nor I_8720 (I151189,I353176,I353185);
nor I_8721 (I151206,I151189,I353191);
nand I_8722 (I151223,I151172,I353197);
not I_8723 (I151240,I151223);
not I_8724 (I151257,I353179);
nor I_8725 (I151114,I151206,I151257);
nand I_8726 (I151288,I151206,I353179);
not I_8727 (I151144,I151288);
not I_8728 (I151319,I353188);
nand I_8729 (I151336,I353185,I353194);
nand I_8730 (I151353,I151336,I353188);
not I_8731 (I151370,I151353);
nand I_8732 (I151387,I151206,I151370);
not I_8733 (I151120,I151387);
nor I_8734 (I151132,I151206,I151370);
nor I_8735 (I151432,I151353,I353179);
DFFARX1 I_8736 (I151432,I2898,I151155,I151135,);
nand I_8737 (I151463,I151336,I151319);
and I_8738 (I151480,I151463,I353182);
nand I_8739 (I151497,I151480,I353179);
nor I_8740 (I151514,I151497,I151353);
not I_8741 (I151531,I151497);
nor I_8742 (I151548,I151240,I151531);
nor I_8743 (I151138,I151548,I151257);
nor I_8744 (I151141,I151240,I151497);
nor I_8745 (I151593,I353182,I353200);
or I_8746 (I151610,I151593,I353188);
nor I_8747 (I151627,I353191,I353176);
and I_8748 (I151644,I151627,I151610);
nor I_8749 (I151661,I151644,I151514);
nor I_8750 (I151126,I151661,I151514);
or I_8751 (I151692,I151497,I151661);
nor I_8752 (I151129,I151223,I151692);
nor I_8753 (I151723,I151370,I151644);
nor I_8754 (I151117,I151257,I151723);
nor I_8755 (I151754,I151531,I151644);
nor I_8756 (I151147,I151754,I151288);
nor I_8757 (I151123,I151644,I151387);
not I_8758 (I151835,I2905);
or I_8759 (I151852,I421278,I421296);
nor I_8760 (I151869,I421278,I421296);
nor I_8761 (I151886,I151869,I421311);
nand I_8762 (I151903,I151852,I421281);
not I_8763 (I151920,I151903);
not I_8764 (I151937,I421284);
nor I_8765 (I151794,I151886,I151937);
nand I_8766 (I151968,I151886,I421284);
not I_8767 (I151824,I151968);
not I_8768 (I151999,I421305);
nand I_8769 (I152016,I421293,I421308);
nand I_8770 (I152033,I152016,I421305);
not I_8771 (I152050,I152033);
nand I_8772 (I152067,I151886,I152050);
not I_8773 (I151800,I152067);
nor I_8774 (I151812,I151886,I152050);
nor I_8775 (I152112,I152033,I421284);
DFFARX1 I_8776 (I152112,I2898,I151835,I151815,);
nand I_8777 (I152143,I152016,I151999);
and I_8778 (I152160,I152143,I421299);
nand I_8779 (I152177,I152160,I421278);
nor I_8780 (I152194,I152177,I152033);
not I_8781 (I152211,I152177);
nor I_8782 (I152228,I151920,I152211);
nor I_8783 (I151818,I152228,I151937);
nor I_8784 (I151821,I151920,I152177);
nor I_8785 (I152273,I421284,I421281);
or I_8786 (I152290,I152273,I421287);
nor I_8787 (I152307,I421302,I421290);
and I_8788 (I152324,I152307,I152290);
nor I_8789 (I152341,I152324,I152194);
nor I_8790 (I151806,I152341,I152194);
or I_8791 (I152372,I152177,I152341);
nor I_8792 (I151809,I151903,I152372);
nor I_8793 (I152403,I152050,I152324);
nor I_8794 (I151797,I151937,I152403);
nor I_8795 (I152434,I152211,I152324);
nor I_8796 (I151827,I152434,I151968);
nor I_8797 (I151803,I152324,I152067);
not I_8798 (I152515,I2905);
or I_8799 (I152532,I362696,I362705);
nor I_8800 (I152549,I362696,I362705);
nor I_8801 (I152566,I152549,I362711);
nand I_8802 (I152583,I152532,I362717);
not I_8803 (I152600,I152583);
not I_8804 (I152617,I362699);
nor I_8805 (I152474,I152566,I152617);
nand I_8806 (I152648,I152566,I362699);
not I_8807 (I152504,I152648);
not I_8808 (I152679,I362708);
nand I_8809 (I152696,I362705,I362714);
nand I_8810 (I152713,I152696,I362708);
not I_8811 (I152730,I152713);
nand I_8812 (I152747,I152566,I152730);
not I_8813 (I152480,I152747);
nor I_8814 (I152492,I152566,I152730);
nor I_8815 (I152792,I152713,I362699);
DFFARX1 I_8816 (I152792,I2898,I152515,I152495,);
nand I_8817 (I152823,I152696,I152679);
and I_8818 (I152840,I152823,I362702);
nand I_8819 (I152857,I152840,I362699);
nor I_8820 (I152874,I152857,I152713);
not I_8821 (I152891,I152857);
nor I_8822 (I152908,I152600,I152891);
nor I_8823 (I152498,I152908,I152617);
nor I_8824 (I152501,I152600,I152857);
nor I_8825 (I152953,I362702,I362720);
or I_8826 (I152970,I152953,I362708);
nor I_8827 (I152987,I362711,I362696);
and I_8828 (I153004,I152987,I152970);
nor I_8829 (I153021,I153004,I152874);
nor I_8830 (I152486,I153021,I152874);
or I_8831 (I153052,I152857,I153021);
nor I_8832 (I152489,I152583,I153052);
nor I_8833 (I153083,I152730,I153004);
nor I_8834 (I152477,I152617,I153083);
nor I_8835 (I153114,I152891,I153004);
nor I_8836 (I152507,I153114,I152648);
nor I_8837 (I152483,I153004,I152747);
not I_8838 (I153195,I2905);
or I_8839 (I153212,I67645,I67642);
nor I_8840 (I153229,I67645,I67642);
nor I_8841 (I153246,I153229,I67627);
nand I_8842 (I153263,I153212,I67651);
not I_8843 (I153280,I153263);
not I_8844 (I153297,I67633);
nor I_8845 (I153154,I153246,I153297);
nand I_8846 (I153328,I153246,I67633);
not I_8847 (I153184,I153328);
not I_8848 (I153359,I67654);
nand I_8849 (I153376,I67630,I67633);
nand I_8850 (I153393,I153376,I67654);
not I_8851 (I153410,I153393);
nand I_8852 (I153427,I153246,I153410);
not I_8853 (I153160,I153427);
nor I_8854 (I153172,I153246,I153410);
nor I_8855 (I153472,I153393,I67633);
DFFARX1 I_8856 (I153472,I2898,I153195,I153175,);
nand I_8857 (I153503,I153376,I153359);
and I_8858 (I153520,I153503,I67639);
nand I_8859 (I153537,I153520,I67639);
nor I_8860 (I153554,I153537,I153393);
not I_8861 (I153571,I153537);
nor I_8862 (I153588,I153280,I153571);
nor I_8863 (I153178,I153588,I153297);
nor I_8864 (I153181,I153280,I153537);
nor I_8865 (I153633,I67648,I67636);
or I_8866 (I153650,I153633,I67636);
nor I_8867 (I153667,I67630,I67627);
and I_8868 (I153684,I153667,I153650);
nor I_8869 (I153701,I153684,I153554);
nor I_8870 (I153166,I153701,I153554);
or I_8871 (I153732,I153537,I153701);
nor I_8872 (I153169,I153263,I153732);
nor I_8873 (I153763,I153410,I153684);
nor I_8874 (I153157,I153297,I153763);
nor I_8875 (I153794,I153571,I153684);
nor I_8876 (I153187,I153794,I153328);
nor I_8877 (I153163,I153684,I153427);
not I_8878 (I153875,I2905);
or I_8879 (I153892,I97825,I97828);
nor I_8880 (I153909,I97825,I97828);
nor I_8881 (I153926,I153909,I97834);
nand I_8882 (I153943,I153892,I97822);
not I_8883 (I153960,I153943);
not I_8884 (I153977,I97819);
nor I_8885 (I153834,I153926,I153977);
nand I_8886 (I154008,I153926,I97819);
not I_8887 (I153864,I154008);
not I_8888 (I154039,I97837);
nand I_8889 (I154056,I97831,I97828);
nand I_8890 (I154073,I154056,I97837);
not I_8891 (I154090,I154073);
nand I_8892 (I154107,I153926,I154090);
not I_8893 (I153840,I154107);
nor I_8894 (I153852,I153926,I154090);
nor I_8895 (I154152,I154073,I97819);
DFFARX1 I_8896 (I154152,I2898,I153875,I153855,);
nand I_8897 (I154183,I154056,I154039);
and I_8898 (I154200,I154183,I97840);
nand I_8899 (I154217,I154200,I97822);
nor I_8900 (I154234,I154217,I154073);
not I_8901 (I154251,I154217);
nor I_8902 (I154268,I153960,I154251);
nor I_8903 (I153858,I154268,I153977);
nor I_8904 (I153861,I153960,I154217);
nor I_8905 (I154313,I97825,I97843);
or I_8906 (I154330,I154313,I97834);
nor I_8907 (I154347,I97831,I97819);
and I_8908 (I154364,I154347,I154330);
nor I_8909 (I154381,I154364,I154234);
nor I_8910 (I153846,I154381,I154234);
or I_8911 (I154412,I154217,I154381);
nor I_8912 (I153849,I153943,I154412);
nor I_8913 (I154443,I154090,I154364);
nor I_8914 (I153837,I153977,I154443);
nor I_8915 (I154474,I154251,I154364);
nor I_8916 (I153867,I154474,I154008);
nor I_8917 (I153843,I154364,I154107);
not I_8918 (I154555,I2905);
or I_8919 (I154572,I67016,I67013);
nor I_8920 (I154589,I67016,I67013);
nor I_8921 (I154606,I154589,I66998);
nand I_8922 (I154623,I154572,I67022);
not I_8923 (I154640,I154623);
not I_8924 (I154657,I67004);
nor I_8925 (I154514,I154606,I154657);
nand I_8926 (I154688,I154606,I67004);
not I_8927 (I154544,I154688);
not I_8928 (I154719,I67025);
nand I_8929 (I154736,I67001,I67004);
nand I_8930 (I154753,I154736,I67025);
not I_8931 (I154770,I154753);
nand I_8932 (I154787,I154606,I154770);
not I_8933 (I154520,I154787);
nor I_8934 (I154532,I154606,I154770);
nor I_8935 (I154832,I154753,I67004);
DFFARX1 I_8936 (I154832,I2898,I154555,I154535,);
nand I_8937 (I154863,I154736,I154719);
and I_8938 (I154880,I154863,I67010);
nand I_8939 (I154897,I154880,I67010);
nor I_8940 (I154914,I154897,I154753);
not I_8941 (I154931,I154897);
nor I_8942 (I154948,I154640,I154931);
nor I_8943 (I154538,I154948,I154657);
nor I_8944 (I154541,I154640,I154897);
nor I_8945 (I154993,I67019,I67007);
or I_8946 (I155010,I154993,I67007);
nor I_8947 (I155027,I67001,I66998);
and I_8948 (I155044,I155027,I155010);
nor I_8949 (I155061,I155044,I154914);
nor I_8950 (I154526,I155061,I154914);
or I_8951 (I155092,I154897,I155061);
nor I_8952 (I154529,I154623,I155092);
nor I_8953 (I155123,I154770,I155044);
nor I_8954 (I154517,I154657,I155123);
nor I_8955 (I155154,I154931,I155044);
nor I_8956 (I154547,I155154,I154688);
nor I_8957 (I154523,I155044,I154787);
not I_8958 (I155235,I2905);
or I_8959 (I155252,I395192,I395192);
nor I_8960 (I155269,I395192,I395192);
nor I_8961 (I155286,I155269,I395204);
nand I_8962 (I155303,I155252,I395183);
not I_8963 (I155320,I155303);
not I_8964 (I155337,I395186);
nor I_8965 (I155194,I155286,I155337);
nand I_8966 (I155368,I155286,I395186);
not I_8967 (I155224,I155368);
not I_8968 (I155399,I395201);
nand I_8969 (I155416,I395195,I395189);
nand I_8970 (I155433,I155416,I395201);
not I_8971 (I155450,I155433);
nand I_8972 (I155467,I155286,I155450);
not I_8973 (I155200,I155467);
nor I_8974 (I155212,I155286,I155450);
nor I_8975 (I155512,I155433,I395186);
DFFARX1 I_8976 (I155512,I2898,I155235,I155215,);
nand I_8977 (I155543,I155416,I155399);
and I_8978 (I155560,I155543,I395195);
nand I_8979 (I155577,I155560,I395189);
nor I_8980 (I155594,I155577,I155433);
not I_8981 (I155611,I155577);
nor I_8982 (I155628,I155320,I155611);
nor I_8983 (I155218,I155628,I155337);
nor I_8984 (I155221,I155320,I155577);
nor I_8985 (I155673,I395186,I395198);
or I_8986 (I155690,I155673,I395198);
nor I_8987 (I155707,I395207,I395183);
and I_8988 (I155724,I155707,I155690);
nor I_8989 (I155741,I155724,I155594);
nor I_8990 (I155206,I155741,I155594);
or I_8991 (I155772,I155577,I155741);
nor I_8992 (I155209,I155303,I155772);
nor I_8993 (I155803,I155450,I155724);
nor I_8994 (I155197,I155337,I155803);
nor I_8995 (I155834,I155611,I155724);
nor I_8996 (I155227,I155834,I155368);
nor I_8997 (I155203,I155724,I155467);
not I_8998 (I155915,I2905);
or I_8999 (I155932,I407432,I407432);
nor I_9000 (I155949,I407432,I407432);
nor I_9001 (I155966,I155949,I407444);
nand I_9002 (I155983,I155932,I407423);
not I_9003 (I156000,I155983);
not I_9004 (I156017,I407426);
nor I_9005 (I155874,I155966,I156017);
nand I_9006 (I156048,I155966,I407426);
not I_9007 (I155904,I156048);
not I_9008 (I156079,I407441);
nand I_9009 (I156096,I407435,I407429);
nand I_9010 (I156113,I156096,I407441);
not I_9011 (I156130,I156113);
nand I_9012 (I156147,I155966,I156130);
not I_9013 (I155880,I156147);
nor I_9014 (I155892,I155966,I156130);
nor I_9015 (I156192,I156113,I407426);
DFFARX1 I_9016 (I156192,I2898,I155915,I155895,);
nand I_9017 (I156223,I156096,I156079);
and I_9018 (I156240,I156223,I407435);
nand I_9019 (I156257,I156240,I407429);
nor I_9020 (I156274,I156257,I156113);
not I_9021 (I156291,I156257);
nor I_9022 (I156308,I156000,I156291);
nor I_9023 (I155898,I156308,I156017);
nor I_9024 (I155901,I156000,I156257);
nor I_9025 (I156353,I407426,I407438);
or I_9026 (I156370,I156353,I407438);
nor I_9027 (I156387,I407447,I407423);
and I_9028 (I156404,I156387,I156370);
nor I_9029 (I156421,I156404,I156274);
nor I_9030 (I155886,I156421,I156274);
or I_9031 (I156452,I156257,I156421);
nor I_9032 (I155889,I155983,I156452);
nor I_9033 (I156483,I156130,I156404);
nor I_9034 (I155877,I156017,I156483);
nor I_9035 (I156514,I156291,I156404);
nor I_9036 (I155907,I156514,I156048);
nor I_9037 (I155883,I156404,I156147);
not I_9038 (I156595,I2905);
or I_9039 (I156612,I55094,I55079);
nor I_9040 (I156629,I55094,I55079);
nor I_9041 (I156646,I156629,I55097);
nand I_9042 (I156663,I156612,I55100);
not I_9043 (I156680,I156663);
not I_9044 (I156697,I55070);
nor I_9045 (I156554,I156646,I156697);
nand I_9046 (I156728,I156646,I55070);
not I_9047 (I156584,I156728);
not I_9048 (I156759,I55064);
nand I_9049 (I156776,I55085,I55064);
nand I_9050 (I156793,I156776,I55064);
not I_9051 (I156810,I156793);
nand I_9052 (I156827,I156646,I156810);
not I_9053 (I156560,I156827);
nor I_9054 (I156572,I156646,I156810);
nor I_9055 (I156872,I156793,I55070);
DFFARX1 I_9056 (I156872,I2898,I156595,I156575,);
nand I_9057 (I156903,I156776,I156759);
and I_9058 (I156920,I156903,I55067);
nand I_9059 (I156937,I156920,I55088);
nor I_9060 (I156954,I156937,I156793);
not I_9061 (I156971,I156937);
nor I_9062 (I156988,I156680,I156971);
nor I_9063 (I156578,I156988,I156697);
nor I_9064 (I156581,I156680,I156937);
nor I_9065 (I157033,I55067,I55073);
or I_9066 (I157050,I157033,I55076);
nor I_9067 (I157067,I55082,I55091);
and I_9068 (I157084,I157067,I157050);
nor I_9069 (I157101,I157084,I156954);
nor I_9070 (I156566,I157101,I156954);
or I_9071 (I157132,I156937,I157101);
nor I_9072 (I156569,I156663,I157132);
nor I_9073 (I157163,I156810,I157084);
nor I_9074 (I156557,I156697,I157163);
nor I_9075 (I157194,I156971,I157084);
nor I_9076 (I156587,I157194,I156728);
nor I_9077 (I156563,I157084,I156827);
not I_9078 (I157275,I2905);
or I_9079 (I157292,I206725,I206704);
nor I_9080 (I157309,I206725,I206704);
nor I_9081 (I157326,I157309,I206707);
nand I_9082 (I157343,I157292,I206731);
not I_9083 (I157360,I157343);
not I_9084 (I157377,I206722);
nor I_9085 (I157234,I157326,I157377);
nand I_9086 (I157408,I157326,I206722);
not I_9087 (I157264,I157408);
not I_9088 (I157439,I206719);
nand I_9089 (I157456,I206713,I206704);
nand I_9090 (I157473,I157456,I206719);
not I_9091 (I157490,I157473);
nand I_9092 (I157507,I157326,I157490);
not I_9093 (I157240,I157507);
nor I_9094 (I157252,I157326,I157490);
nor I_9095 (I157552,I157473,I206722);
DFFARX1 I_9096 (I157552,I2898,I157275,I157255,);
nand I_9097 (I157583,I157456,I157439);
and I_9098 (I157600,I157583,I206716);
nand I_9099 (I157617,I157600,I206716);
nor I_9100 (I157634,I157617,I157473);
not I_9101 (I157651,I157617);
nor I_9102 (I157668,I157360,I157651);
nor I_9103 (I157258,I157668,I157377);
nor I_9104 (I157261,I157360,I157617);
nor I_9105 (I157713,I206710,I206713);
or I_9106 (I157730,I157713,I206707);
nor I_9107 (I157747,I206728,I206710);
and I_9108 (I157764,I157747,I157730);
nor I_9109 (I157781,I157764,I157634);
nor I_9110 (I157246,I157781,I157634);
or I_9111 (I157812,I157617,I157781);
nor I_9112 (I157249,I157343,I157812);
nor I_9113 (I157843,I157490,I157764);
nor I_9114 (I157237,I157377,I157843);
nor I_9115 (I157874,I157651,I157764);
nor I_9116 (I157267,I157874,I157408);
nor I_9117 (I157243,I157764,I157507);
not I_9118 (I157955,I2905);
or I_9119 (I157972,I358531,I358540);
nor I_9120 (I157989,I358531,I358540);
nor I_9121 (I158006,I157989,I358546);
nand I_9122 (I158023,I157972,I358552);
not I_9123 (I158040,I158023);
not I_9124 (I158057,I358534);
nor I_9125 (I157914,I158006,I158057);
nand I_9126 (I158088,I158006,I358534);
not I_9127 (I157944,I158088);
not I_9128 (I158119,I358543);
nand I_9129 (I158136,I358540,I358549);
nand I_9130 (I158153,I158136,I358543);
not I_9131 (I158170,I158153);
nand I_9132 (I158187,I158006,I158170);
not I_9133 (I157920,I158187);
nor I_9134 (I157932,I158006,I158170);
nor I_9135 (I158232,I158153,I358534);
DFFARX1 I_9136 (I158232,I2898,I157955,I157935,);
nand I_9137 (I158263,I158136,I158119);
and I_9138 (I158280,I158263,I358537);
nand I_9139 (I158297,I158280,I358534);
nor I_9140 (I158314,I158297,I158153);
not I_9141 (I158331,I158297);
nor I_9142 (I158348,I158040,I158331);
nor I_9143 (I157938,I158348,I158057);
nor I_9144 (I157941,I158040,I158297);
nor I_9145 (I158393,I358537,I358555);
or I_9146 (I158410,I158393,I358543);
nor I_9147 (I158427,I358546,I358531);
and I_9148 (I158444,I158427,I158410);
nor I_9149 (I158461,I158444,I158314);
nor I_9150 (I157926,I158461,I158314);
or I_9151 (I158492,I158297,I158461);
nor I_9152 (I157929,I158023,I158492);
nor I_9153 (I158523,I158170,I158444);
nor I_9154 (I157917,I158057,I158523);
nor I_9155 (I158554,I158331,I158444);
nor I_9156 (I157947,I158554,I158088);
nor I_9157 (I157923,I158444,I158187);
not I_9158 (I158635,I2905);
or I_9159 (I158652,I351391,I351400);
nor I_9160 (I158669,I351391,I351400);
nor I_9161 (I158686,I158669,I351406);
nand I_9162 (I158703,I158652,I351412);
not I_9163 (I158720,I158703);
not I_9164 (I158737,I351394);
nor I_9165 (I158594,I158686,I158737);
nand I_9166 (I158768,I158686,I351394);
not I_9167 (I158624,I158768);
not I_9168 (I158799,I351403);
nand I_9169 (I158816,I351400,I351409);
nand I_9170 (I158833,I158816,I351403);
not I_9171 (I158850,I158833);
nand I_9172 (I158867,I158686,I158850);
not I_9173 (I158600,I158867);
nor I_9174 (I158612,I158686,I158850);
nor I_9175 (I158912,I158833,I351394);
DFFARX1 I_9176 (I158912,I2898,I158635,I158615,);
nand I_9177 (I158943,I158816,I158799);
and I_9178 (I158960,I158943,I351397);
nand I_9179 (I158977,I158960,I351394);
nor I_9180 (I158994,I158977,I158833);
not I_9181 (I159011,I158977);
nor I_9182 (I159028,I158720,I159011);
nor I_9183 (I158618,I159028,I158737);
nor I_9184 (I158621,I158720,I158977);
nor I_9185 (I159073,I351397,I351415);
or I_9186 (I159090,I159073,I351403);
nor I_9187 (I159107,I351406,I351391);
and I_9188 (I159124,I159107,I159090);
nor I_9189 (I159141,I159124,I158994);
nor I_9190 (I158606,I159141,I158994);
or I_9191 (I159172,I158977,I159141);
nor I_9192 (I158609,I158703,I159172);
nor I_9193 (I159203,I158850,I159124);
nor I_9194 (I158597,I158737,I159203);
nor I_9195 (I159234,I159011,I159124);
nor I_9196 (I158627,I159234,I158768);
nor I_9197 (I158603,I159124,I158867);
not I_9198 (I159315,I2905);
or I_9199 (I159332,I214205,I214184);
nor I_9200 (I159349,I214205,I214184);
nor I_9201 (I159366,I159349,I214187);
nand I_9202 (I159383,I159332,I214211);
not I_9203 (I159400,I159383);
not I_9204 (I159417,I214202);
nor I_9205 (I159274,I159366,I159417);
nand I_9206 (I159448,I159366,I214202);
not I_9207 (I159304,I159448);
not I_9208 (I159479,I214199);
nand I_9209 (I159496,I214193,I214184);
nand I_9210 (I159513,I159496,I214199);
not I_9211 (I159530,I159513);
nand I_9212 (I159547,I159366,I159530);
not I_9213 (I159280,I159547);
nor I_9214 (I159292,I159366,I159530);
nor I_9215 (I159592,I159513,I214202);
DFFARX1 I_9216 (I159592,I2898,I159315,I159295,);
nand I_9217 (I159623,I159496,I159479);
and I_9218 (I159640,I159623,I214196);
nand I_9219 (I159657,I159640,I214196);
nor I_9220 (I159674,I159657,I159513);
not I_9221 (I159691,I159657);
nor I_9222 (I159708,I159400,I159691);
nor I_9223 (I159298,I159708,I159417);
nor I_9224 (I159301,I159400,I159657);
nor I_9225 (I159753,I214190,I214193);
or I_9226 (I159770,I159753,I214187);
nor I_9227 (I159787,I214208,I214190);
and I_9228 (I159804,I159787,I159770);
nor I_9229 (I159821,I159804,I159674);
nor I_9230 (I159286,I159821,I159674);
or I_9231 (I159852,I159657,I159821);
nor I_9232 (I159289,I159383,I159852);
nor I_9233 (I159883,I159530,I159804);
nor I_9234 (I159277,I159417,I159883);
nor I_9235 (I159914,I159691,I159804);
nor I_9236 (I159307,I159914,I159448);
nor I_9237 (I159283,I159804,I159547);
not I_9238 (I159995,I2905);
or I_9239 (I160012,I15376,I15352);
nor I_9240 (I160029,I15376,I15352);
nor I_9241 (I160046,I160029,I15364);
nand I_9242 (I160063,I160012,I15361);
not I_9243 (I160080,I160063);
not I_9244 (I160097,I15352);
nor I_9245 (I159954,I160046,I160097);
nand I_9246 (I160128,I160046,I15352);
not I_9247 (I159984,I160128);
not I_9248 (I160159,I15370);
nand I_9249 (I160176,I15379,I15358);
nand I_9250 (I160193,I160176,I15370);
not I_9251 (I160210,I160193);
nand I_9252 (I160227,I160046,I160210);
not I_9253 (I159960,I160227);
nor I_9254 (I159972,I160046,I160210);
nor I_9255 (I160272,I160193,I15352);
DFFARX1 I_9256 (I160272,I2898,I159995,I159975,);
nand I_9257 (I160303,I160176,I160159);
and I_9258 (I160320,I160303,I15367);
nand I_9259 (I160337,I160320,I15361);
nor I_9260 (I160354,I160337,I160193);
not I_9261 (I160371,I160337);
nor I_9262 (I160388,I160080,I160371);
nor I_9263 (I159978,I160388,I160097);
nor I_9264 (I159981,I160080,I160337);
nor I_9265 (I160433,I15355,I15373);
or I_9266 (I160450,I160433,I15358);
nor I_9267 (I160467,I15355,I15364);
and I_9268 (I160484,I160467,I160450);
nor I_9269 (I160501,I160484,I160354);
nor I_9270 (I159966,I160501,I160354);
or I_9271 (I160532,I160337,I160501);
nor I_9272 (I159969,I160063,I160532);
nor I_9273 (I160563,I160210,I160484);
nor I_9274 (I159957,I160097,I160563);
nor I_9275 (I160594,I160371,I160484);
nor I_9276 (I159987,I160594,I160128);
nor I_9277 (I159963,I160484,I160227);
not I_9278 (I160675,I2905);
or I_9279 (I160692,I86515,I86512);
nor I_9280 (I160709,I86515,I86512);
nor I_9281 (I160726,I160709,I86497);
nand I_9282 (I160743,I160692,I86521);
not I_9283 (I160760,I160743);
not I_9284 (I160777,I86503);
nor I_9285 (I160634,I160726,I160777);
nand I_9286 (I160808,I160726,I86503);
not I_9287 (I160664,I160808);
not I_9288 (I160839,I86524);
nand I_9289 (I160856,I86500,I86503);
nand I_9290 (I160873,I160856,I86524);
not I_9291 (I160890,I160873);
nand I_9292 (I160907,I160726,I160890);
not I_9293 (I160640,I160907);
nor I_9294 (I160652,I160726,I160890);
nor I_9295 (I160952,I160873,I86503);
DFFARX1 I_9296 (I160952,I2898,I160675,I160655,);
nand I_9297 (I160983,I160856,I160839);
and I_9298 (I161000,I160983,I86509);
nand I_9299 (I161017,I161000,I86509);
nor I_9300 (I161034,I161017,I160873);
not I_9301 (I161051,I161017);
nor I_9302 (I161068,I160760,I161051);
nor I_9303 (I160658,I161068,I160777);
nor I_9304 (I160661,I160760,I161017);
nor I_9305 (I161113,I86518,I86506);
or I_9306 (I161130,I161113,I86506);
nor I_9307 (I161147,I86500,I86497);
and I_9308 (I161164,I161147,I161130);
nor I_9309 (I161181,I161164,I161034);
nor I_9310 (I160646,I161181,I161034);
or I_9311 (I161212,I161017,I161181);
nor I_9312 (I160649,I160743,I161212);
nor I_9313 (I161243,I160890,I161164);
nor I_9314 (I160637,I160777,I161243);
nor I_9315 (I161274,I161051,I161164);
nor I_9316 (I160667,I161274,I160808);
nor I_9317 (I160643,I161164,I160907);
not I_9318 (I161355,I2905);
or I_9319 (I161372,I304722,I304698);
nor I_9320 (I161389,I304722,I304698);
nor I_9321 (I161406,I161389,I304698);
nand I_9322 (I161423,I161372,I304716);
not I_9323 (I161440,I161423);
not I_9324 (I161457,I304704);
nor I_9325 (I161314,I161406,I161457);
nand I_9326 (I161488,I161406,I304704);
not I_9327 (I161344,I161488);
not I_9328 (I161519,I304707);
nand I_9329 (I161536,I304701,I304692);
nand I_9330 (I161553,I161536,I304707);
not I_9331 (I161570,I161553);
nand I_9332 (I161587,I161406,I161570);
not I_9333 (I161320,I161587);
nor I_9334 (I161332,I161406,I161570);
nor I_9335 (I161632,I161553,I304704);
DFFARX1 I_9336 (I161632,I2898,I161355,I161335,);
nand I_9337 (I161663,I161536,I161519);
and I_9338 (I161680,I161663,I304719);
nand I_9339 (I161697,I161680,I304713);
nor I_9340 (I161714,I161697,I161553);
not I_9341 (I161731,I161697);
nor I_9342 (I161748,I161440,I161731);
nor I_9343 (I161338,I161748,I161457);
nor I_9344 (I161341,I161440,I161697);
nor I_9345 (I161793,I304710,I304701);
or I_9346 (I161810,I161793,I304692);
nor I_9347 (I161827,I304695,I304695);
and I_9348 (I161844,I161827,I161810);
nor I_9349 (I161861,I161844,I161714);
nor I_9350 (I161326,I161861,I161714);
or I_9351 (I161892,I161697,I161861);
nor I_9352 (I161329,I161423,I161892);
nor I_9353 (I161923,I161570,I161844);
nor I_9354 (I161317,I161457,I161923);
nor I_9355 (I161954,I161731,I161844);
nor I_9356 (I161347,I161954,I161488);
nor I_9357 (I161323,I161844,I161587);
not I_9358 (I162035,I2905);
or I_9359 (I162052,I415005,I415023);
nor I_9360 (I162069,I415005,I415023);
nor I_9361 (I162086,I162069,I415038);
nand I_9362 (I162103,I162052,I415008);
not I_9363 (I162120,I162103);
not I_9364 (I162137,I415011);
nor I_9365 (I161994,I162086,I162137);
nand I_9366 (I162168,I162086,I415011);
not I_9367 (I162024,I162168);
not I_9368 (I162199,I415032);
nand I_9369 (I162216,I415020,I415035);
nand I_9370 (I162233,I162216,I415032);
not I_9371 (I162250,I162233);
nand I_9372 (I162267,I162086,I162250);
not I_9373 (I162000,I162267);
nor I_9374 (I162012,I162086,I162250);
nor I_9375 (I162312,I162233,I415011);
DFFARX1 I_9376 (I162312,I2898,I162035,I162015,);
nand I_9377 (I162343,I162216,I162199);
and I_9378 (I162360,I162343,I415026);
nand I_9379 (I162377,I162360,I415005);
nor I_9380 (I162394,I162377,I162233);
not I_9381 (I162411,I162377);
nor I_9382 (I162428,I162120,I162411);
nor I_9383 (I162018,I162428,I162137);
nor I_9384 (I162021,I162120,I162377);
nor I_9385 (I162473,I415011,I415008);
or I_9386 (I162490,I162473,I415014);
nor I_9387 (I162507,I415029,I415017);
and I_9388 (I162524,I162507,I162490);
nor I_9389 (I162541,I162524,I162394);
nor I_9390 (I162006,I162541,I162394);
or I_9391 (I162572,I162377,I162541);
nor I_9392 (I162009,I162103,I162572);
nor I_9393 (I162603,I162250,I162524);
nor I_9394 (I161997,I162137,I162603);
nor I_9395 (I162634,I162411,I162524);
nor I_9396 (I162027,I162634,I162168);
nor I_9397 (I162003,I162524,I162267);
not I_9398 (I162715,I2905);
or I_9399 (I162732,I217197,I217176);
nor I_9400 (I162749,I217197,I217176);
nor I_9401 (I162766,I162749,I217179);
nand I_9402 (I162783,I162732,I217203);
not I_9403 (I162800,I162783);
not I_9404 (I162817,I217194);
nor I_9405 (I162674,I162766,I162817);
nand I_9406 (I162848,I162766,I217194);
not I_9407 (I162704,I162848);
not I_9408 (I162879,I217191);
nand I_9409 (I162896,I217185,I217176);
nand I_9410 (I162913,I162896,I217191);
not I_9411 (I162930,I162913);
nand I_9412 (I162947,I162766,I162930);
not I_9413 (I162680,I162947);
nor I_9414 (I162692,I162766,I162930);
nor I_9415 (I162992,I162913,I217194);
DFFARX1 I_9416 (I162992,I2898,I162715,I162695,);
nand I_9417 (I163023,I162896,I162879);
and I_9418 (I163040,I163023,I217188);
nand I_9419 (I163057,I163040,I217188);
nor I_9420 (I163074,I163057,I162913);
not I_9421 (I163091,I163057);
nor I_9422 (I163108,I162800,I163091);
nor I_9423 (I162698,I163108,I162817);
nor I_9424 (I162701,I162800,I163057);
nor I_9425 (I163153,I217182,I217185);
or I_9426 (I163170,I163153,I217179);
nor I_9427 (I163187,I217200,I217182);
and I_9428 (I163204,I163187,I163170);
nor I_9429 (I163221,I163204,I163074);
nor I_9430 (I162686,I163221,I163074);
or I_9431 (I163252,I163057,I163221);
nor I_9432 (I162689,I162783,I163252);
nor I_9433 (I163283,I162930,I163204);
nor I_9434 (I162677,I162817,I163283);
nor I_9435 (I163314,I163091,I163204);
nor I_9436 (I162707,I163314,I162848);
nor I_9437 (I162683,I163204,I162947);
not I_9438 (I163395,I2905);
or I_9439 (I163412,I250548,I250551);
nor I_9440 (I163429,I250548,I250551);
nor I_9441 (I163446,I163429,I250533);
nand I_9442 (I163463,I163412,I250560);
not I_9443 (I163480,I163463);
not I_9444 (I163497,I250545);
nor I_9445 (I163354,I163446,I163497);
nand I_9446 (I163528,I163446,I250545);
not I_9447 (I163384,I163528);
not I_9448 (I163559,I250557);
nand I_9449 (I163576,I250536,I250539);
nand I_9450 (I163593,I163576,I250557);
not I_9451 (I163610,I163593);
nand I_9452 (I163627,I163446,I163610);
not I_9453 (I163360,I163627);
nor I_9454 (I163372,I163446,I163610);
nor I_9455 (I163672,I163593,I250545);
DFFARX1 I_9456 (I163672,I2898,I163395,I163375,);
nand I_9457 (I163703,I163576,I163559);
and I_9458 (I163720,I163703,I250533);
nand I_9459 (I163737,I163720,I250542);
nor I_9460 (I163754,I163737,I163593);
not I_9461 (I163771,I163737);
nor I_9462 (I163788,I163480,I163771);
nor I_9463 (I163378,I163788,I163497);
nor I_9464 (I163381,I163480,I163737);
nor I_9465 (I163833,I250530,I250530);
or I_9466 (I163850,I163833,I250554);
nor I_9467 (I163867,I250536,I250539);
and I_9468 (I163884,I163867,I163850);
nor I_9469 (I163901,I163884,I163754);
nor I_9470 (I163366,I163901,I163754);
or I_9471 (I163932,I163737,I163901);
nor I_9472 (I163369,I163463,I163932);
nor I_9473 (I163963,I163610,I163884);
nor I_9474 (I163357,I163497,I163963);
nor I_9475 (I163994,I163771,I163884);
nor I_9476 (I163387,I163994,I163528);
nor I_9477 (I163363,I163884,I163627);
not I_9478 (I164075,I2905);
or I_9479 (I164092,I360316,I360325);
nor I_9480 (I164109,I360316,I360325);
nor I_9481 (I164126,I164109,I360331);
nand I_9482 (I164143,I164092,I360337);
not I_9483 (I164160,I164143);
not I_9484 (I164177,I360319);
nor I_9485 (I164034,I164126,I164177);
nand I_9486 (I164208,I164126,I360319);
not I_9487 (I164064,I164208);
not I_9488 (I164239,I360328);
nand I_9489 (I164256,I360325,I360334);
nand I_9490 (I164273,I164256,I360328);
not I_9491 (I164290,I164273);
nand I_9492 (I164307,I164126,I164290);
not I_9493 (I164040,I164307);
nor I_9494 (I164052,I164126,I164290);
nor I_9495 (I164352,I164273,I360319);
DFFARX1 I_9496 (I164352,I2898,I164075,I164055,);
nand I_9497 (I164383,I164256,I164239);
and I_9498 (I164400,I164383,I360322);
nand I_9499 (I164417,I164400,I360319);
nor I_9500 (I164434,I164417,I164273);
not I_9501 (I164451,I164417);
nor I_9502 (I164468,I164160,I164451);
nor I_9503 (I164058,I164468,I164177);
nor I_9504 (I164061,I164160,I164417);
nor I_9505 (I164513,I360322,I360340);
or I_9506 (I164530,I164513,I360328);
nor I_9507 (I164547,I360331,I360316);
and I_9508 (I164564,I164547,I164530);
nor I_9509 (I164581,I164564,I164434);
nor I_9510 (I164046,I164581,I164434);
or I_9511 (I164612,I164417,I164581);
nor I_9512 (I164049,I164143,I164612);
nor I_9513 (I164643,I164290,I164564);
nor I_9514 (I164037,I164177,I164643);
nor I_9515 (I164674,I164451,I164564);
nor I_9516 (I164067,I164674,I164208);
nor I_9517 (I164043,I164564,I164307);
not I_9518 (I164755,I2905);
or I_9519 (I164772,I36082,I36058);
nor I_9520 (I164789,I36082,I36058);
nor I_9521 (I164806,I164789,I36070);
nand I_9522 (I164823,I164772,I36067);
not I_9523 (I164840,I164823);
not I_9524 (I164857,I36058);
nor I_9525 (I164714,I164806,I164857);
nand I_9526 (I164888,I164806,I36058);
not I_9527 (I164744,I164888);
not I_9528 (I164919,I36076);
nand I_9529 (I164936,I36085,I36064);
nand I_9530 (I164953,I164936,I36076);
not I_9531 (I164970,I164953);
nand I_9532 (I164987,I164806,I164970);
not I_9533 (I164720,I164987);
nor I_9534 (I164732,I164806,I164970);
nor I_9535 (I165032,I164953,I36058);
DFFARX1 I_9536 (I165032,I2898,I164755,I164735,);
nand I_9537 (I165063,I164936,I164919);
and I_9538 (I165080,I165063,I36073);
nand I_9539 (I165097,I165080,I36067);
nor I_9540 (I165114,I165097,I164953);
not I_9541 (I165131,I165097);
nor I_9542 (I165148,I164840,I165131);
nor I_9543 (I164738,I165148,I164857);
nor I_9544 (I164741,I164840,I165097);
nor I_9545 (I165193,I36061,I36079);
or I_9546 (I165210,I165193,I36064);
nor I_9547 (I165227,I36061,I36070);
and I_9548 (I165244,I165227,I165210);
nor I_9549 (I165261,I165244,I165114);
nor I_9550 (I164726,I165261,I165114);
or I_9551 (I165292,I165097,I165261);
nor I_9552 (I164729,I164823,I165292);
nor I_9553 (I165323,I164970,I165244);
nor I_9554 (I164717,I164857,I165323);
nor I_9555 (I165354,I165131,I165244);
nor I_9556 (I164747,I165354,I164888);
nor I_9557 (I164723,I165244,I164987);
not I_9558 (I165435,I2905);
or I_9559 (I165452,I73306,I73303);
nor I_9560 (I165469,I73306,I73303);
nor I_9561 (I165486,I165469,I73288);
nand I_9562 (I165503,I165452,I73312);
not I_9563 (I165520,I165503);
not I_9564 (I165537,I73294);
nor I_9565 (I165394,I165486,I165537);
nand I_9566 (I165568,I165486,I73294);
not I_9567 (I165424,I165568);
not I_9568 (I165599,I73315);
nand I_9569 (I165616,I73291,I73294);
nand I_9570 (I165633,I165616,I73315);
not I_9571 (I165650,I165633);
nand I_9572 (I165667,I165486,I165650);
not I_9573 (I165400,I165667);
nor I_9574 (I165412,I165486,I165650);
nor I_9575 (I165712,I165633,I73294);
DFFARX1 I_9576 (I165712,I2898,I165435,I165415,);
nand I_9577 (I165743,I165616,I165599);
and I_9578 (I165760,I165743,I73300);
nand I_9579 (I165777,I165760,I73300);
nor I_9580 (I165794,I165777,I165633);
not I_9581 (I165811,I165777);
nor I_9582 (I165828,I165520,I165811);
nor I_9583 (I165418,I165828,I165537);
nor I_9584 (I165421,I165520,I165777);
nor I_9585 (I165873,I73309,I73297);
or I_9586 (I165890,I165873,I73297);
nor I_9587 (I165907,I73291,I73288);
and I_9588 (I165924,I165907,I165890);
nor I_9589 (I165941,I165924,I165794);
nor I_9590 (I165406,I165941,I165794);
or I_9591 (I165972,I165777,I165941);
nor I_9592 (I165409,I165503,I165972);
nor I_9593 (I166003,I165650,I165924);
nor I_9594 (I165397,I165537,I166003);
nor I_9595 (I166034,I165811,I165924);
nor I_9596 (I165427,I166034,I165568);
nor I_9597 (I165403,I165924,I165667);
not I_9598 (I166115,I2905);
or I_9599 (I166132,I416399,I416417);
nor I_9600 (I166149,I416399,I416417);
nor I_9601 (I166166,I166149,I416432);
nand I_9602 (I166183,I166132,I416402);
not I_9603 (I166200,I166183);
not I_9604 (I166217,I416405);
nor I_9605 (I166074,I166166,I166217);
nand I_9606 (I166248,I166166,I416405);
not I_9607 (I166104,I166248);
not I_9608 (I166279,I416426);
nand I_9609 (I166296,I416414,I416429);
nand I_9610 (I166313,I166296,I416426);
not I_9611 (I166330,I166313);
nand I_9612 (I166347,I166166,I166330);
not I_9613 (I166080,I166347);
nor I_9614 (I166092,I166166,I166330);
nor I_9615 (I166392,I166313,I416405);
DFFARX1 I_9616 (I166392,I2898,I166115,I166095,);
nand I_9617 (I166423,I166296,I166279);
and I_9618 (I166440,I166423,I416420);
nand I_9619 (I166457,I166440,I416399);
nor I_9620 (I166474,I166457,I166313);
not I_9621 (I166491,I166457);
nor I_9622 (I166508,I166200,I166491);
nor I_9623 (I166098,I166508,I166217);
nor I_9624 (I166101,I166200,I166457);
nor I_9625 (I166553,I416405,I416402);
or I_9626 (I166570,I166553,I416408);
nor I_9627 (I166587,I416423,I416411);
and I_9628 (I166604,I166587,I166570);
nor I_9629 (I166621,I166604,I166474);
nor I_9630 (I166086,I166621,I166474);
or I_9631 (I166652,I166457,I166621);
nor I_9632 (I166089,I166183,I166652);
nor I_9633 (I166683,I166330,I166604);
nor I_9634 (I166077,I166217,I166683);
nor I_9635 (I166714,I166491,I166604);
nor I_9636 (I166107,I166714,I166248);
nor I_9637 (I166083,I166604,I166347);
not I_9638 (I166795,I2905);
or I_9639 (I166812,I83370,I83367);
nor I_9640 (I166829,I83370,I83367);
nor I_9641 (I166846,I166829,I83352);
nand I_9642 (I166863,I166812,I83376);
not I_9643 (I166880,I166863);
not I_9644 (I166897,I83358);
nor I_9645 (I166754,I166846,I166897);
nand I_9646 (I166928,I166846,I83358);
not I_9647 (I166784,I166928);
not I_9648 (I166959,I83379);
nand I_9649 (I166976,I83355,I83358);
nand I_9650 (I166993,I166976,I83379);
not I_9651 (I167010,I166993);
nand I_9652 (I167027,I166846,I167010);
not I_9653 (I166760,I167027);
nor I_9654 (I166772,I166846,I167010);
nor I_9655 (I167072,I166993,I83358);
DFFARX1 I_9656 (I167072,I2898,I166795,I166775,);
nand I_9657 (I167103,I166976,I166959);
and I_9658 (I167120,I167103,I83364);
nand I_9659 (I167137,I167120,I83364);
nor I_9660 (I167154,I167137,I166993);
not I_9661 (I167171,I167137);
nor I_9662 (I167188,I166880,I167171);
nor I_9663 (I166778,I167188,I166897);
nor I_9664 (I166781,I166880,I167137);
nor I_9665 (I167233,I83373,I83361);
or I_9666 (I167250,I167233,I83361);
nor I_9667 (I167267,I83355,I83352);
and I_9668 (I167284,I167267,I167250);
nor I_9669 (I167301,I167284,I167154);
nor I_9670 (I166766,I167301,I167154);
or I_9671 (I167332,I167137,I167301);
nor I_9672 (I166769,I166863,I167332);
nor I_9673 (I167363,I167010,I167284);
nor I_9674 (I166757,I166897,I167363);
nor I_9675 (I167394,I167171,I167284);
nor I_9676 (I166787,I167394,I166928);
nor I_9677 (I166763,I167284,I167027);
not I_9678 (I167475,I2905);
or I_9679 (I167492,I208969,I208948);
nor I_9680 (I167509,I208969,I208948);
nor I_9681 (I167526,I167509,I208951);
nand I_9682 (I167543,I167492,I208975);
not I_9683 (I167560,I167543);
not I_9684 (I167577,I208966);
nor I_9685 (I167434,I167526,I167577);
nand I_9686 (I167608,I167526,I208966);
not I_9687 (I167464,I167608);
not I_9688 (I167639,I208963);
nand I_9689 (I167656,I208957,I208948);
nand I_9690 (I167673,I167656,I208963);
not I_9691 (I167690,I167673);
nand I_9692 (I167707,I167526,I167690);
not I_9693 (I167440,I167707);
nor I_9694 (I167452,I167526,I167690);
nor I_9695 (I167752,I167673,I208966);
DFFARX1 I_9696 (I167752,I2898,I167475,I167455,);
nand I_9697 (I167783,I167656,I167639);
and I_9698 (I167800,I167783,I208960);
nand I_9699 (I167817,I167800,I208960);
nor I_9700 (I167834,I167817,I167673);
not I_9701 (I167851,I167817);
nor I_9702 (I167868,I167560,I167851);
nor I_9703 (I167458,I167868,I167577);
nor I_9704 (I167461,I167560,I167817);
nor I_9705 (I167913,I208954,I208957);
or I_9706 (I167930,I167913,I208951);
nor I_9707 (I167947,I208972,I208954);
and I_9708 (I167964,I167947,I167930);
nor I_9709 (I167981,I167964,I167834);
nor I_9710 (I167446,I167981,I167834);
or I_9711 (I168012,I167817,I167981);
nor I_9712 (I167449,I167543,I168012);
nor I_9713 (I168043,I167690,I167964);
nor I_9714 (I167437,I167577,I168043);
nor I_9715 (I168074,I167851,I167964);
nor I_9716 (I167467,I168074,I167608);
nor I_9717 (I167443,I167964,I167707);
not I_9718 (I168155,I2905);
or I_9719 (I168172,I357341,I357350);
nor I_9720 (I168189,I357341,I357350);
nor I_9721 (I168206,I168189,I357356);
nand I_9722 (I168223,I168172,I357362);
not I_9723 (I168240,I168223);
not I_9724 (I168257,I357344);
nor I_9725 (I168114,I168206,I168257);
nand I_9726 (I168288,I168206,I357344);
not I_9727 (I168144,I168288);
not I_9728 (I168319,I357353);
nand I_9729 (I168336,I357350,I357359);
nand I_9730 (I168353,I168336,I357353);
not I_9731 (I168370,I168353);
nand I_9732 (I168387,I168206,I168370);
not I_9733 (I168120,I168387);
nor I_9734 (I168132,I168206,I168370);
nor I_9735 (I168432,I168353,I357344);
DFFARX1 I_9736 (I168432,I2898,I168155,I168135,);
nand I_9737 (I168463,I168336,I168319);
and I_9738 (I168480,I168463,I357347);
nand I_9739 (I168497,I168480,I357344);
nor I_9740 (I168514,I168497,I168353);
not I_9741 (I168531,I168497);
nor I_9742 (I168548,I168240,I168531);
nor I_9743 (I168138,I168548,I168257);
nor I_9744 (I168141,I168240,I168497);
nor I_9745 (I168593,I357347,I357365);
or I_9746 (I168610,I168593,I357353);
nor I_9747 (I168627,I357356,I357341);
and I_9748 (I168644,I168627,I168610);
nor I_9749 (I168661,I168644,I168514);
nor I_9750 (I168126,I168661,I168514);
or I_9751 (I168692,I168497,I168661);
nor I_9752 (I168129,I168223,I168692);
nor I_9753 (I168723,I168370,I168644);
nor I_9754 (I168117,I168257,I168723);
nor I_9755 (I168754,I168531,I168644);
nor I_9756 (I168147,I168754,I168288);
nor I_9757 (I168123,I168644,I168387);
not I_9758 (I168835,I2905);
or I_9759 (I168852,I388723,I388750);
nor I_9760 (I168869,I388723,I388750);
nor I_9761 (I168886,I168869,I388726);
nand I_9762 (I168903,I168852,I388741);
not I_9763 (I168920,I168903);
not I_9764 (I168937,I388747);
nor I_9765 (I168794,I168886,I168937);
nand I_9766 (I168968,I168886,I388747);
not I_9767 (I168824,I168968);
not I_9768 (I168999,I388738);
nand I_9769 (I169016,I388735,I388729);
nand I_9770 (I169033,I169016,I388738);
not I_9771 (I169050,I169033);
nand I_9772 (I169067,I168886,I169050);
not I_9773 (I168800,I169067);
nor I_9774 (I168812,I168886,I169050);
nor I_9775 (I169112,I169033,I388747);
DFFARX1 I_9776 (I169112,I2898,I168835,I168815,);
nand I_9777 (I169143,I169016,I168999);
and I_9778 (I169160,I169143,I388726);
nand I_9779 (I169177,I169160,I388753);
nor I_9780 (I169194,I169177,I169033);
not I_9781 (I169211,I169177);
nor I_9782 (I169228,I168920,I169211);
nor I_9783 (I168818,I169228,I168937);
nor I_9784 (I168821,I168920,I169177);
nor I_9785 (I169273,I388723,I388729);
or I_9786 (I169290,I169273,I388744);
nor I_9787 (I169307,I388756,I388732);
and I_9788 (I169324,I169307,I169290);
nor I_9789 (I169341,I169324,I169194);
nor I_9790 (I168806,I169341,I169194);
or I_9791 (I169372,I169177,I169341);
nor I_9792 (I168809,I168903,I169372);
nor I_9793 (I169403,I169050,I169324);
nor I_9794 (I168797,I168937,I169403);
nor I_9795 (I169434,I169211,I169324);
nor I_9796 (I168827,I169434,I168968);
nor I_9797 (I168803,I169324,I169067);
not I_9798 (I169515,I2905);
or I_9799 (I169532,I366505,I366499);
nor I_9800 (I169549,I366505,I366499);
nor I_9801 (I169566,I169549,I366511);
nand I_9802 (I169583,I169532,I366514);
not I_9803 (I169600,I169583);
not I_9804 (I169617,I366517);
nor I_9805 (I169474,I169566,I169617);
nand I_9806 (I169648,I169566,I366517);
not I_9807 (I169504,I169648);
not I_9808 (I169679,I366502);
nand I_9809 (I169696,I366493,I366490);
nand I_9810 (I169713,I169696,I366502);
not I_9811 (I169730,I169713);
nand I_9812 (I169747,I169566,I169730);
not I_9813 (I169480,I169747);
nor I_9814 (I169492,I169566,I169730);
nor I_9815 (I169792,I169713,I366517);
DFFARX1 I_9816 (I169792,I2898,I169515,I169495,);
nand I_9817 (I169823,I169696,I169679);
and I_9818 (I169840,I169823,I366487);
nand I_9819 (I169857,I169840,I366496);
nor I_9820 (I169874,I169857,I169713);
not I_9821 (I169891,I169857);
nor I_9822 (I169908,I169600,I169891);
nor I_9823 (I169498,I169908,I169617);
nor I_9824 (I169501,I169600,I169857);
nor I_9825 (I169953,I366490,I366520);
or I_9826 (I169970,I169953,I366487);
nor I_9827 (I169987,I366508,I366493);
and I_9828 (I170004,I169987,I169970);
nor I_9829 (I170021,I170004,I169874);
nor I_9830 (I169486,I170021,I169874);
or I_9831 (I170052,I169857,I170021);
nor I_9832 (I169489,I169583,I170052);
nor I_9833 (I170083,I169730,I170004);
nor I_9834 (I169477,I169617,I170083);
nor I_9835 (I170114,I169891,I170004);
nor I_9836 (I169507,I170114,I169648);
nor I_9837 (I169483,I170004,I169747);
not I_9838 (I170195,I2905);
or I_9839 (I170212,I445673,I445691);
nor I_9840 (I170229,I445673,I445691);
nor I_9841 (I170246,I170229,I445706);
nand I_9842 (I170263,I170212,I445676);
not I_9843 (I170280,I170263);
not I_9844 (I170297,I445679);
nor I_9845 (I170154,I170246,I170297);
nand I_9846 (I170328,I170246,I445679);
not I_9847 (I170184,I170328);
not I_9848 (I170359,I445700);
nand I_9849 (I170376,I445688,I445703);
nand I_9850 (I170393,I170376,I445700);
not I_9851 (I170410,I170393);
nand I_9852 (I170427,I170246,I170410);
not I_9853 (I170160,I170427);
nor I_9854 (I170172,I170246,I170410);
nor I_9855 (I170472,I170393,I445679);
DFFARX1 I_9856 (I170472,I2898,I170195,I170175,);
nand I_9857 (I170503,I170376,I170359);
and I_9858 (I170520,I170503,I445694);
nand I_9859 (I170537,I170520,I445673);
nor I_9860 (I170554,I170537,I170393);
not I_9861 (I170571,I170537);
nor I_9862 (I170588,I170280,I170571);
nor I_9863 (I170178,I170588,I170297);
nor I_9864 (I170181,I170280,I170537);
nor I_9865 (I170633,I445679,I445676);
or I_9866 (I170650,I170633,I445682);
nor I_9867 (I170667,I445697,I445685);
and I_9868 (I170684,I170667,I170650);
nor I_9869 (I170701,I170684,I170554);
nor I_9870 (I170166,I170701,I170554);
or I_9871 (I170732,I170537,I170701);
nor I_9872 (I170169,I170263,I170732);
nor I_9873 (I170763,I170410,I170684);
nor I_9874 (I170157,I170297,I170763);
nor I_9875 (I170794,I170571,I170684);
nor I_9876 (I170187,I170794,I170328);
nor I_9877 (I170163,I170684,I170427);
not I_9878 (I170875,I2905);
or I_9879 (I170892,I260493,I260496);
nor I_9880 (I170909,I260493,I260496);
nor I_9881 (I170926,I170909,I260478);
nand I_9882 (I170943,I170892,I260505);
not I_9883 (I170960,I170943);
not I_9884 (I170977,I260490);
nor I_9885 (I170834,I170926,I170977);
nand I_9886 (I171008,I170926,I260490);
not I_9887 (I170864,I171008);
not I_9888 (I171039,I260502);
nand I_9889 (I171056,I260481,I260484);
nand I_9890 (I171073,I171056,I260502);
not I_9891 (I171090,I171073);
nand I_9892 (I171107,I170926,I171090);
not I_9893 (I170840,I171107);
nor I_9894 (I170852,I170926,I171090);
nor I_9895 (I171152,I171073,I260490);
DFFARX1 I_9896 (I171152,I2898,I170875,I170855,);
nand I_9897 (I171183,I171056,I171039);
and I_9898 (I171200,I171183,I260478);
nand I_9899 (I171217,I171200,I260487);
nor I_9900 (I171234,I171217,I171073);
not I_9901 (I171251,I171217);
nor I_9902 (I171268,I170960,I171251);
nor I_9903 (I170858,I171268,I170977);
nor I_9904 (I170861,I170960,I171217);
nor I_9905 (I171313,I260475,I260475);
or I_9906 (I171330,I171313,I260499);
nor I_9907 (I171347,I260481,I260484);
and I_9908 (I171364,I171347,I171330);
nor I_9909 (I171381,I171364,I171234);
nor I_9910 (I170846,I171381,I171234);
or I_9911 (I171412,I171217,I171381);
nor I_9912 (I170849,I170943,I171412);
nor I_9913 (I171443,I171090,I171364);
nor I_9914 (I170837,I170977,I171443);
nor I_9915 (I171474,I171251,I171364);
nor I_9916 (I170867,I171474,I171008);
nor I_9917 (I170843,I171364,I171107);
not I_9918 (I171555,I2905);
or I_9919 (I171572,I253608,I253611);
nor I_9920 (I171589,I253608,I253611);
nor I_9921 (I171606,I171589,I253593);
nand I_9922 (I171623,I171572,I253620);
not I_9923 (I171640,I171623);
not I_9924 (I171657,I253605);
nor I_9925 (I171514,I171606,I171657);
nand I_9926 (I171688,I171606,I253605);
not I_9927 (I171544,I171688);
not I_9928 (I171719,I253617);
nand I_9929 (I171736,I253596,I253599);
nand I_9930 (I171753,I171736,I253617);
not I_9931 (I171770,I171753);
nand I_9932 (I171787,I171606,I171770);
not I_9933 (I171520,I171787);
nor I_9934 (I171532,I171606,I171770);
nor I_9935 (I171832,I171753,I253605);
DFFARX1 I_9936 (I171832,I2898,I171555,I171535,);
nand I_9937 (I171863,I171736,I171719);
and I_9938 (I171880,I171863,I253593);
nand I_9939 (I171897,I171880,I253602);
nor I_9940 (I171914,I171897,I171753);
not I_9941 (I171931,I171897);
nor I_9942 (I171948,I171640,I171931);
nor I_9943 (I171538,I171948,I171657);
nor I_9944 (I171541,I171640,I171897);
nor I_9945 (I171993,I253590,I253590);
or I_9946 (I172010,I171993,I253614);
nor I_9947 (I172027,I253596,I253599);
and I_9948 (I172044,I172027,I172010);
nor I_9949 (I172061,I172044,I171914);
nor I_9950 (I171526,I172061,I171914);
or I_9951 (I172092,I171897,I172061);
nor I_9952 (I171529,I171623,I172092);
nor I_9953 (I172123,I171770,I172044);
nor I_9954 (I171517,I171657,I172123);
nor I_9955 (I172154,I171931,I172044);
nor I_9956 (I171547,I172154,I171688);
nor I_9957 (I171523,I172044,I171787);
not I_9958 (I172235,I2905);
or I_9959 (I172252,I261258,I261261);
nor I_9960 (I172269,I261258,I261261);
nor I_9961 (I172286,I172269,I261243);
nand I_9962 (I172303,I172252,I261270);
not I_9963 (I172320,I172303);
not I_9964 (I172337,I261255);
nor I_9965 (I172194,I172286,I172337);
nand I_9966 (I172368,I172286,I261255);
not I_9967 (I172224,I172368);
not I_9968 (I172399,I261267);
nand I_9969 (I172416,I261246,I261249);
nand I_9970 (I172433,I172416,I261267);
not I_9971 (I172450,I172433);
nand I_9972 (I172467,I172286,I172450);
not I_9973 (I172200,I172467);
nor I_9974 (I172212,I172286,I172450);
nor I_9975 (I172512,I172433,I261255);
DFFARX1 I_9976 (I172512,I2898,I172235,I172215,);
nand I_9977 (I172543,I172416,I172399);
and I_9978 (I172560,I172543,I261243);
nand I_9979 (I172577,I172560,I261252);
nor I_9980 (I172594,I172577,I172433);
not I_9981 (I172611,I172577);
nor I_9982 (I172628,I172320,I172611);
nor I_9983 (I172218,I172628,I172337);
nor I_9984 (I172221,I172320,I172577);
nor I_9985 (I172673,I261240,I261240);
or I_9986 (I172690,I172673,I261264);
nor I_9987 (I172707,I261246,I261249);
and I_9988 (I172724,I172707,I172690);
nor I_9989 (I172741,I172724,I172594);
nor I_9990 (I172206,I172741,I172594);
or I_9991 (I172772,I172577,I172741);
nor I_9992 (I172209,I172303,I172772);
nor I_9993 (I172803,I172450,I172724);
nor I_9994 (I172197,I172337,I172803);
nor I_9995 (I172834,I172611,I172724);
nor I_9996 (I172227,I172834,I172368);
nor I_9997 (I172203,I172724,I172467);
not I_9998 (I172915,I2905);
or I_9999 (I172932,I138057,I138027);
nor I_10000 (I172949,I138057,I138027);
nor I_10001 (I172966,I172949,I138048);
nand I_10002 (I172983,I172932,I138030);
not I_10003 (I173000,I172983);
not I_10004 (I173017,I138036);
nor I_10005 (I172874,I172966,I173017);
nand I_10006 (I173048,I172966,I138036);
not I_10007 (I172904,I173048);
not I_10008 (I173079,I138042);
nand I_10009 (I173096,I138027,I138039);
nand I_10010 (I173113,I173096,I138042);
not I_10011 (I173130,I173113);
nand I_10012 (I173147,I172966,I173130);
not I_10013 (I172880,I173147);
nor I_10014 (I172892,I172966,I173130);
nor I_10015 (I173192,I173113,I138036);
DFFARX1 I_10016 (I173192,I2898,I172915,I172895,);
nand I_10017 (I173223,I173096,I173079);
and I_10018 (I173240,I173223,I138024);
nand I_10019 (I173257,I173240,I138054);
nor I_10020 (I173274,I173257,I173113);
not I_10021 (I173291,I173257);
nor I_10022 (I173308,I173000,I173291);
nor I_10023 (I172898,I173308,I173017);
nor I_10024 (I172901,I173000,I173257);
nor I_10025 (I173353,I138030,I138051);
or I_10026 (I173370,I173353,I138045);
nor I_10027 (I173387,I138024,I138033);
and I_10028 (I173404,I173387,I173370);
nor I_10029 (I173421,I173404,I173274);
nor I_10030 (I172886,I173421,I173274);
or I_10031 (I173452,I173257,I173421);
nor I_10032 (I172889,I172983,I173452);
nor I_10033 (I173483,I173130,I173404);
nor I_10034 (I172877,I173017,I173483);
nor I_10035 (I173514,I173291,I173404);
nor I_10036 (I172907,I173514,I173048);
nor I_10037 (I172883,I173404,I173147);
not I_10038 (I173595,I2905);
or I_10039 (I173612,I334136,I334145);
nor I_10040 (I173629,I334136,I334145);
nor I_10041 (I173646,I173629,I334151);
nand I_10042 (I173663,I173612,I334157);
not I_10043 (I173680,I173663);
not I_10044 (I173697,I334139);
nor I_10045 (I173554,I173646,I173697);
nand I_10046 (I173728,I173646,I334139);
not I_10047 (I173584,I173728);
not I_10048 (I173759,I334148);
nand I_10049 (I173776,I334145,I334154);
nand I_10050 (I173793,I173776,I334148);
not I_10051 (I173810,I173793);
nand I_10052 (I173827,I173646,I173810);
not I_10053 (I173560,I173827);
nor I_10054 (I173572,I173646,I173810);
nor I_10055 (I173872,I173793,I334139);
DFFARX1 I_10056 (I173872,I2898,I173595,I173575,);
nand I_10057 (I173903,I173776,I173759);
and I_10058 (I173920,I173903,I334142);
nand I_10059 (I173937,I173920,I334139);
nor I_10060 (I173954,I173937,I173793);
not I_10061 (I173971,I173937);
nor I_10062 (I173988,I173680,I173971);
nor I_10063 (I173578,I173988,I173697);
nor I_10064 (I173581,I173680,I173937);
nor I_10065 (I174033,I334142,I334160);
or I_10066 (I174050,I174033,I334148);
nor I_10067 (I174067,I334151,I334136);
and I_10068 (I174084,I174067,I174050);
nor I_10069 (I174101,I174084,I173954);
nor I_10070 (I173566,I174101,I173954);
or I_10071 (I174132,I173937,I174101);
nor I_10072 (I173569,I173663,I174132);
nor I_10073 (I174163,I173810,I174084);
nor I_10074 (I173557,I173697,I174163);
nor I_10075 (I174194,I173971,I174084);
nor I_10076 (I173587,I174194,I173728);
nor I_10077 (I173563,I174084,I173827);
not I_10078 (I174275,I2905);
or I_10079 (I174292,I126106,I126076);
nor I_10080 (I174309,I126106,I126076);
nor I_10081 (I174326,I174309,I126097);
nand I_10082 (I174343,I174292,I126079);
not I_10083 (I174360,I174343);
not I_10084 (I174377,I126085);
nor I_10085 (I174234,I174326,I174377);
nand I_10086 (I174408,I174326,I126085);
not I_10087 (I174264,I174408);
not I_10088 (I174439,I126091);
nand I_10089 (I174456,I126076,I126088);
nand I_10090 (I174473,I174456,I126091);
not I_10091 (I174490,I174473);
nand I_10092 (I174507,I174326,I174490);
not I_10093 (I174240,I174507);
nor I_10094 (I174252,I174326,I174490);
nor I_10095 (I174552,I174473,I126085);
DFFARX1 I_10096 (I174552,I2898,I174275,I174255,);
nand I_10097 (I174583,I174456,I174439);
and I_10098 (I174600,I174583,I126073);
nand I_10099 (I174617,I174600,I126103);
nor I_10100 (I174634,I174617,I174473);
not I_10101 (I174651,I174617);
nor I_10102 (I174668,I174360,I174651);
nor I_10103 (I174258,I174668,I174377);
nor I_10104 (I174261,I174360,I174617);
nor I_10105 (I174713,I126079,I126100);
or I_10106 (I174730,I174713,I126094);
nor I_10107 (I174747,I126073,I126082);
and I_10108 (I174764,I174747,I174730);
nor I_10109 (I174781,I174764,I174634);
nor I_10110 (I174246,I174781,I174634);
or I_10111 (I174812,I174617,I174781);
nor I_10112 (I174249,I174343,I174812);
nor I_10113 (I174843,I174490,I174764);
nor I_10114 (I174237,I174377,I174843);
nor I_10115 (I174874,I174651,I174764);
nor I_10116 (I174267,I174874,I174408);
nor I_10117 (I174243,I174764,I174507);
not I_10118 (I174955,I2905);
or I_10119 (I174972,I392599,I392626);
nor I_10120 (I174989,I392599,I392626);
nor I_10121 (I175006,I174989,I392602);
nand I_10122 (I175023,I174972,I392617);
not I_10123 (I175040,I175023);
not I_10124 (I175057,I392623);
nor I_10125 (I174914,I175006,I175057);
nand I_10126 (I175088,I175006,I392623);
not I_10127 (I174944,I175088);
not I_10128 (I175119,I392614);
nand I_10129 (I175136,I392611,I392605);
nand I_10130 (I175153,I175136,I392614);
not I_10131 (I175170,I175153);
nand I_10132 (I175187,I175006,I175170);
not I_10133 (I174920,I175187);
nor I_10134 (I174932,I175006,I175170);
nor I_10135 (I175232,I175153,I392623);
DFFARX1 I_10136 (I175232,I2898,I174955,I174935,);
nand I_10137 (I175263,I175136,I175119);
and I_10138 (I175280,I175263,I392602);
nand I_10139 (I175297,I175280,I392629);
nor I_10140 (I175314,I175297,I175153);
not I_10141 (I175331,I175297);
nor I_10142 (I175348,I175040,I175331);
nor I_10143 (I174938,I175348,I175057);
nor I_10144 (I174941,I175040,I175297);
nor I_10145 (I175393,I392599,I392605);
or I_10146 (I175410,I175393,I392620);
nor I_10147 (I175427,I392632,I392608);
and I_10148 (I175444,I175427,I175410);
nor I_10149 (I175461,I175444,I175314);
nor I_10150 (I174926,I175461,I175314);
or I_10151 (I175492,I175297,I175461);
nor I_10152 (I174929,I175023,I175492);
nor I_10153 (I175523,I175170,I175444);
nor I_10154 (I174917,I175057,I175523);
nor I_10155 (I175554,I175331,I175444);
nor I_10156 (I174947,I175554,I175088);
nor I_10157 (I174923,I175444,I175187);
not I_10158 (I175635,I2905);
or I_10159 (I175652,I239073,I239076);
nor I_10160 (I175669,I239073,I239076);
nor I_10161 (I175686,I175669,I239058);
nand I_10162 (I175703,I175652,I239085);
not I_10163 (I175720,I175703);
not I_10164 (I175737,I239070);
nor I_10165 (I175594,I175686,I175737);
nand I_10166 (I175768,I175686,I239070);
not I_10167 (I175624,I175768);
not I_10168 (I175799,I239082);
nand I_10169 (I175816,I239061,I239064);
nand I_10170 (I175833,I175816,I239082);
not I_10171 (I175850,I175833);
nand I_10172 (I175867,I175686,I175850);
not I_10173 (I175600,I175867);
nor I_10174 (I175612,I175686,I175850);
nor I_10175 (I175912,I175833,I239070);
DFFARX1 I_10176 (I175912,I2898,I175635,I175615,);
nand I_10177 (I175943,I175816,I175799);
and I_10178 (I175960,I175943,I239058);
nand I_10179 (I175977,I175960,I239067);
nor I_10180 (I175994,I175977,I175833);
not I_10181 (I176011,I175977);
nor I_10182 (I176028,I175720,I176011);
nor I_10183 (I175618,I176028,I175737);
nor I_10184 (I175621,I175720,I175977);
nor I_10185 (I176073,I239055,I239055);
or I_10186 (I176090,I176073,I239079);
nor I_10187 (I176107,I239061,I239064);
and I_10188 (I176124,I176107,I176090);
nor I_10189 (I176141,I176124,I175994);
nor I_10190 (I175606,I176141,I175994);
or I_10191 (I176172,I175977,I176141);
nor I_10192 (I175609,I175703,I176172);
nor I_10193 (I176203,I175850,I176124);
nor I_10194 (I175597,I175737,I176203);
nor I_10195 (I176234,I176011,I176124);
nor I_10196 (I175627,I176234,I175768);
nor I_10197 (I175603,I176124,I175867);
not I_10198 (I176315,I2905);
or I_10199 (I176332,I114784,I114754);
nor I_10200 (I176349,I114784,I114754);
nor I_10201 (I176366,I176349,I114775);
nand I_10202 (I176383,I176332,I114757);
not I_10203 (I176400,I176383);
not I_10204 (I176417,I114763);
nor I_10205 (I176274,I176366,I176417);
nand I_10206 (I176448,I176366,I114763);
not I_10207 (I176304,I176448);
not I_10208 (I176479,I114769);
nand I_10209 (I176496,I114754,I114766);
nand I_10210 (I176513,I176496,I114769);
not I_10211 (I176530,I176513);
nand I_10212 (I176547,I176366,I176530);
not I_10213 (I176280,I176547);
nor I_10214 (I176292,I176366,I176530);
nor I_10215 (I176592,I176513,I114763);
DFFARX1 I_10216 (I176592,I2898,I176315,I176295,);
nand I_10217 (I176623,I176496,I176479);
and I_10218 (I176640,I176623,I114751);
nand I_10219 (I176657,I176640,I114781);
nor I_10220 (I176674,I176657,I176513);
not I_10221 (I176691,I176657);
nor I_10222 (I176708,I176400,I176691);
nor I_10223 (I176298,I176708,I176417);
nor I_10224 (I176301,I176400,I176657);
nor I_10225 (I176753,I114757,I114778);
or I_10226 (I176770,I176753,I114772);
nor I_10227 (I176787,I114751,I114760);
and I_10228 (I176804,I176787,I176770);
nor I_10229 (I176821,I176804,I176674);
nor I_10230 (I176286,I176821,I176674);
or I_10231 (I176852,I176657,I176821);
nor I_10232 (I176289,I176383,I176852);
nor I_10233 (I176883,I176530,I176804);
nor I_10234 (I176277,I176417,I176883);
nor I_10235 (I176914,I176691,I176804);
nor I_10236 (I176307,I176914,I176448);
nor I_10237 (I176283,I176804,I176547);
not I_10238 (I176995,I2905);
or I_10239 (I177012,I245958,I245961);
nor I_10240 (I177029,I245958,I245961);
nor I_10241 (I177046,I177029,I245943);
nand I_10242 (I177063,I177012,I245970);
not I_10243 (I177080,I177063);
not I_10244 (I177097,I245955);
nor I_10245 (I176954,I177046,I177097);
nand I_10246 (I177128,I177046,I245955);
not I_10247 (I176984,I177128);
not I_10248 (I177159,I245967);
nand I_10249 (I177176,I245946,I245949);
nand I_10250 (I177193,I177176,I245967);
not I_10251 (I177210,I177193);
nand I_10252 (I177227,I177046,I177210);
not I_10253 (I176960,I177227);
nor I_10254 (I176972,I177046,I177210);
nor I_10255 (I177272,I177193,I245955);
DFFARX1 I_10256 (I177272,I2898,I176995,I176975,);
nand I_10257 (I177303,I177176,I177159);
and I_10258 (I177320,I177303,I245943);
nand I_10259 (I177337,I177320,I245952);
nor I_10260 (I177354,I177337,I177193);
not I_10261 (I177371,I177337);
nor I_10262 (I177388,I177080,I177371);
nor I_10263 (I176978,I177388,I177097);
nor I_10264 (I176981,I177080,I177337);
nor I_10265 (I177433,I245940,I245940);
or I_10266 (I177450,I177433,I245964);
nor I_10267 (I177467,I245946,I245949);
and I_10268 (I177484,I177467,I177450);
nor I_10269 (I177501,I177484,I177354);
nor I_10270 (I176966,I177501,I177354);
or I_10271 (I177532,I177337,I177501);
nor I_10272 (I176969,I177063,I177532);
nor I_10273 (I177563,I177210,I177484);
nor I_10274 (I176957,I177097,I177563);
nor I_10275 (I177594,I177371,I177484);
nor I_10276 (I176987,I177594,I177128);
nor I_10277 (I176963,I177484,I177227);
not I_10278 (I177672,I2905);
nand I_10279 (I177689,I131764,I131743);
and I_10280 (I177706,I177689,I131734);
DFFARX1 I_10281 (I177706,I2898,I177672,I177732,);
nor I_10282 (I177740,I131749,I131743);
or I_10283 (I177757,I131749,I131743);
not I_10284 (I177774,I131767);
nor I_10285 (I177791,I131761,I131767);
nor I_10286 (I177808,I131746,I131761);
or I_10287 (I177825,I177732,I131746);
nor I_10288 (I177842,I131740,I131737);
not I_10289 (I177859,I177842);
nor I_10290 (I177876,I177842,I177791);
nand I_10291 (I177893,I177876,I177740);
not I_10292 (I177910,I131740);
nand I_10293 (I177927,I177910,I131752);
nand I_10294 (I177944,I177927,I177774);
nand I_10295 (I177961,I177944,I177893);
DFFARX1 I_10296 (I177961,I2898,I177672,I177643,);
and I_10297 (I177992,I177910,I131752);
nor I_10298 (I178009,I177992,I131767);
nor I_10299 (I177655,I177732,I178009);
nor I_10300 (I178040,I131734,I131740);
DFFARX1 I_10301 (I178040,I2898,I177672,I178066,);
nor I_10302 (I177634,I178066,I177859);
not I_10303 (I178088,I178066);
nand I_10304 (I177664,I177808,I178088);
nor I_10305 (I178119,I177825,I131734);
nor I_10306 (I177661,I178066,I178119);
not I_10307 (I178150,I131734);
nand I_10308 (I178167,I131737,I131755);
and I_10309 (I178184,I178167,I177791);
nor I_10310 (I177637,I178184,I177859);
not I_10311 (I178215,I178167);
nor I_10312 (I178232,I177732,I178215);
DFFARX1 I_10313 (I178232,I2898,I177672,I177652,);
or I_10314 (I178263,I178167,I131758);
nand I_10315 (I177640,I177740,I178263);
nor I_10316 (I178294,I178167,I131758);
and I_10317 (I178311,I177808,I178294);
nand I_10318 (I177649,I178311,I177757);
nand I_10319 (I177646,I178311,I178150);
nand I_10320 (I177658,I177808,I178167);
not I_10321 (I178403,I2905);
nand I_10322 (I178420,I267366,I267384);
and I_10323 (I178437,I178420,I267378);
DFFARX1 I_10324 (I178437,I2898,I178403,I178463,);
nor I_10325 (I178471,I267372,I267384);
or I_10326 (I178488,I267372,I267384);
not I_10327 (I178505,I267390);
nor I_10328 (I178522,I267366,I267390);
nor I_10329 (I178539,I267387,I267366);
or I_10330 (I178556,I178463,I267387);
nor I_10331 (I178573,I267360,I267363);
not I_10332 (I178590,I178573);
nor I_10333 (I178607,I178573,I178522);
nand I_10334 (I178624,I178607,I178471);
not I_10335 (I178641,I267360);
nand I_10336 (I178658,I178641,I267369);
nand I_10337 (I178675,I178658,I178505);
nand I_10338 (I178692,I178675,I178624);
DFFARX1 I_10339 (I178692,I2898,I178403,I178374,);
and I_10340 (I178723,I178641,I267369);
nor I_10341 (I178740,I178723,I267390);
nor I_10342 (I178386,I178463,I178740);
nor I_10343 (I178771,I267375,I267369);
DFFARX1 I_10344 (I178771,I2898,I178403,I178797,);
nor I_10345 (I178365,I178797,I178590);
not I_10346 (I178819,I178797);
nand I_10347 (I178395,I178539,I178819);
nor I_10348 (I178850,I178556,I267375);
nor I_10349 (I178392,I178797,I178850);
not I_10350 (I178881,I267375);
nand I_10351 (I178898,I267381,I267360);
and I_10352 (I178915,I178898,I178522);
nor I_10353 (I178368,I178915,I178590);
not I_10354 (I178946,I178898);
nor I_10355 (I178963,I178463,I178946);
DFFARX1 I_10356 (I178963,I2898,I178403,I178383,);
or I_10357 (I178994,I178898,I267363);
nand I_10358 (I178371,I178471,I178994);
nor I_10359 (I179025,I178898,I267363);
and I_10360 (I179042,I178539,I179025);
nand I_10361 (I178380,I179042,I178488);
nand I_10362 (I178377,I179042,I178881);
nand I_10363 (I178389,I178539,I178898);
not I_10364 (I179134,I2905);
nand I_10365 (I179151,I425466,I425478);
and I_10366 (I179168,I179151,I425475);
DFFARX1 I_10367 (I179168,I2898,I179134,I179194,);
nor I_10368 (I179202,I425481,I425478);
or I_10369 (I179219,I425481,I425478);
not I_10370 (I179236,I425493);
nor I_10371 (I179253,I425484,I425493);
nor I_10372 (I179270,I425460,I425484);
or I_10373 (I179287,I179194,I425460);
nor I_10374 (I179304,I425460,I425487);
not I_10375 (I179321,I179304);
nor I_10376 (I179338,I179304,I179253);
nand I_10377 (I179355,I179338,I179202);
not I_10378 (I179372,I425460);
nand I_10379 (I179389,I179372,I425463);
nand I_10380 (I179406,I179389,I179236);
nand I_10381 (I179423,I179406,I179355);
DFFARX1 I_10382 (I179423,I2898,I179134,I179105,);
and I_10383 (I179454,I179372,I425463);
nor I_10384 (I179471,I179454,I425493);
nor I_10385 (I179117,I179194,I179471);
nor I_10386 (I179502,I425469,I425472);
DFFARX1 I_10387 (I179502,I2898,I179134,I179528,);
nor I_10388 (I179096,I179528,I179321);
not I_10389 (I179550,I179528);
nand I_10390 (I179126,I179270,I179550);
nor I_10391 (I179581,I179287,I425469);
nor I_10392 (I179123,I179528,I179581);
not I_10393 (I179612,I425469);
nand I_10394 (I179629,I425490,I425466);
and I_10395 (I179646,I179629,I179253);
nor I_10396 (I179099,I179646,I179321);
not I_10397 (I179677,I179629);
nor I_10398 (I179694,I179194,I179677);
DFFARX1 I_10399 (I179694,I2898,I179134,I179114,);
or I_10400 (I179725,I179629,I425463);
nand I_10401 (I179102,I179202,I179725);
nor I_10402 (I179756,I179629,I425463);
and I_10403 (I179773,I179270,I179756);
nand I_10404 (I179111,I179773,I179219);
nand I_10405 (I179108,I179773,I179612);
nand I_10406 (I179120,I179270,I179629);
not I_10407 (I179865,I2905);
nand I_10408 (I179882,I317128,I317143);
and I_10409 (I179899,I179882,I317119);
DFFARX1 I_10410 (I179899,I2898,I179865,I179925,);
nor I_10411 (I179933,I317125,I317143);
or I_10412 (I179950,I317125,I317143);
not I_10413 (I179967,I317146);
nor I_10414 (I179984,I317122,I317146);
nor I_10415 (I180001,I317149,I317122);
or I_10416 (I180018,I179925,I317149);
nor I_10417 (I180035,I317131,I317134);
not I_10418 (I180052,I180035);
nor I_10419 (I180069,I180035,I179984);
nand I_10420 (I180086,I180069,I179933);
not I_10421 (I180103,I317131);
nand I_10422 (I180120,I180103,I317128);
nand I_10423 (I180137,I180120,I179967);
nand I_10424 (I180154,I180137,I180086);
DFFARX1 I_10425 (I180154,I2898,I179865,I179836,);
and I_10426 (I180185,I180103,I317128);
nor I_10427 (I180202,I180185,I317146);
nor I_10428 (I179848,I179925,I180202);
nor I_10429 (I180233,I317119,I317125);
DFFARX1 I_10430 (I180233,I2898,I179865,I180259,);
nor I_10431 (I179827,I180259,I180052);
not I_10432 (I180281,I180259);
nand I_10433 (I179857,I180001,I180281);
nor I_10434 (I180312,I180018,I317119);
nor I_10435 (I179854,I180259,I180312);
not I_10436 (I180343,I317119);
nand I_10437 (I180360,I317140,I317137);
and I_10438 (I180377,I180360,I179984);
nor I_10439 (I179830,I180377,I180052);
not I_10440 (I180408,I180360);
nor I_10441 (I180425,I179925,I180408);
DFFARX1 I_10442 (I180425,I2898,I179865,I179845,);
or I_10443 (I180456,I180360,I317122);
nand I_10444 (I179833,I179933,I180456);
nor I_10445 (I180487,I180360,I317122);
and I_10446 (I180504,I180001,I180487);
nand I_10447 (I179842,I180504,I179950);
nand I_10448 (I179839,I180504,I180343);
nand I_10449 (I179851,I180001,I180360);
not I_10450 (I180596,I2905);
nand I_10451 (I180613,I32491,I32506);
and I_10452 (I180630,I180613,I32509);
DFFARX1 I_10453 (I180630,I2898,I180596,I180656,);
nor I_10454 (I180664,I32488,I32506);
or I_10455 (I180681,I32488,I32506);
not I_10456 (I180698,I32500);
nor I_10457 (I180715,I32503,I32500);
nor I_10458 (I180732,I32488,I32503);
or I_10459 (I180749,I180656,I32488);
nor I_10460 (I180766,I32515,I32500);
not I_10461 (I180783,I180766);
nor I_10462 (I180800,I180766,I180715);
nand I_10463 (I180817,I180800,I180664);
not I_10464 (I180834,I32515);
nand I_10465 (I180851,I180834,I32497);
nand I_10466 (I180868,I180851,I180698);
nand I_10467 (I180885,I180868,I180817);
DFFARX1 I_10468 (I180885,I2898,I180596,I180567,);
and I_10469 (I180916,I180834,I32497);
nor I_10470 (I180933,I180916,I32500);
nor I_10471 (I180579,I180656,I180933);
nor I_10472 (I180964,I32494,I32491);
DFFARX1 I_10473 (I180964,I2898,I180596,I180990,);
nor I_10474 (I180558,I180990,I180783);
not I_10475 (I181012,I180990);
nand I_10476 (I180588,I180732,I181012);
nor I_10477 (I181043,I180749,I32494);
nor I_10478 (I180585,I180990,I181043);
not I_10479 (I181074,I32494);
nand I_10480 (I181091,I32512,I32497);
and I_10481 (I181108,I181091,I180715);
nor I_10482 (I180561,I181108,I180783);
not I_10483 (I181139,I181091);
nor I_10484 (I181156,I180656,I181139);
DFFARX1 I_10485 (I181156,I2898,I180596,I180576,);
or I_10486 (I181187,I181091,I32494);
nand I_10487 (I180564,I180664,I181187);
nor I_10488 (I181218,I181091,I32494);
and I_10489 (I181235,I180732,I181218);
nand I_10490 (I180573,I181235,I180681);
nand I_10491 (I180570,I181235,I181074);
nand I_10492 (I180582,I180732,I181091);
not I_10493 (I181327,I2905);
nand I_10494 (I181344,I249006,I249024);
and I_10495 (I181361,I181344,I249018);
DFFARX1 I_10496 (I181361,I2898,I181327,I181387,);
nor I_10497 (I181395,I249012,I249024);
or I_10498 (I181412,I249012,I249024);
not I_10499 (I181429,I249030);
nor I_10500 (I181446,I249006,I249030);
nor I_10501 (I181463,I249027,I249006);
or I_10502 (I181480,I181387,I249027);
nor I_10503 (I181497,I249000,I249003);
not I_10504 (I181514,I181497);
nor I_10505 (I181531,I181497,I181446);
nand I_10506 (I181548,I181531,I181395);
not I_10507 (I181565,I249000);
nand I_10508 (I181582,I181565,I249009);
nand I_10509 (I181599,I181582,I181429);
nand I_10510 (I181616,I181599,I181548);
DFFARX1 I_10511 (I181616,I2898,I181327,I181298,);
and I_10512 (I181647,I181565,I249009);
nor I_10513 (I181664,I181647,I249030);
nor I_10514 (I181310,I181387,I181664);
nor I_10515 (I181695,I249015,I249009);
DFFARX1 I_10516 (I181695,I2898,I181327,I181721,);
nor I_10517 (I181289,I181721,I181514);
not I_10518 (I181743,I181721);
nand I_10519 (I181319,I181463,I181743);
nor I_10520 (I181774,I181480,I249015);
nor I_10521 (I181316,I181721,I181774);
not I_10522 (I181805,I249015);
nand I_10523 (I181822,I249021,I249000);
and I_10524 (I181839,I181822,I181446);
nor I_10525 (I181292,I181839,I181514);
not I_10526 (I181870,I181822);
nor I_10527 (I181887,I181387,I181870);
DFFARX1 I_10528 (I181887,I2898,I181327,I181307,);
or I_10529 (I181918,I181822,I249003);
nand I_10530 (I181295,I181395,I181918);
nor I_10531 (I181949,I181822,I249003);
and I_10532 (I181966,I181463,I181949);
nand I_10533 (I181304,I181966,I181412);
nand I_10534 (I181301,I181966,I181805);
nand I_10535 (I181313,I181463,I181822);
not I_10536 (I182058,I2905);
nand I_10537 (I182075,I318590,I318605);
and I_10538 (I182092,I182075,I318581);
DFFARX1 I_10539 (I182092,I2898,I182058,I182118,);
nor I_10540 (I182126,I318587,I318605);
or I_10541 (I182143,I318587,I318605);
not I_10542 (I182160,I318608);
nor I_10543 (I182177,I318584,I318608);
nor I_10544 (I182194,I318611,I318584);
or I_10545 (I182211,I182118,I318611);
nor I_10546 (I182228,I318593,I318596);
not I_10547 (I182245,I182228);
nor I_10548 (I182262,I182228,I182177);
nand I_10549 (I182279,I182262,I182126);
not I_10550 (I182296,I318593);
nand I_10551 (I182313,I182296,I318590);
nand I_10552 (I182330,I182313,I182160);
nand I_10553 (I182347,I182330,I182279);
DFFARX1 I_10554 (I182347,I2898,I182058,I182029,);
and I_10555 (I182378,I182296,I318590);
nor I_10556 (I182395,I182378,I318608);
nor I_10557 (I182041,I182118,I182395);
nor I_10558 (I182426,I318581,I318587);
DFFARX1 I_10559 (I182426,I2898,I182058,I182452,);
nor I_10560 (I182020,I182452,I182245);
not I_10561 (I182474,I182452);
nand I_10562 (I182050,I182194,I182474);
nor I_10563 (I182505,I182211,I318581);
nor I_10564 (I182047,I182452,I182505);
not I_10565 (I182536,I318581);
nand I_10566 (I182553,I318602,I318599);
and I_10567 (I182570,I182553,I182177);
nor I_10568 (I182023,I182570,I182245);
not I_10569 (I182601,I182553);
nor I_10570 (I182618,I182118,I182601);
DFFARX1 I_10571 (I182618,I2898,I182058,I182038,);
or I_10572 (I182649,I182553,I318584);
nand I_10573 (I182026,I182126,I182649);
nor I_10574 (I182680,I182553,I318584);
and I_10575 (I182697,I182194,I182680);
nand I_10576 (I182035,I182697,I182143);
nand I_10577 (I182032,I182697,I182536);
nand I_10578 (I182044,I182194,I182553);
not I_10579 (I182783,I2905);
nand I_10580 (I182800,I294479,I294461);
and I_10581 (I182817,I182800,I294470);
DFFARX1 I_10582 (I182817,I2898,I182783,I182843,);
not I_10583 (I182851,I182843);
nor I_10584 (I182868,I294464,I294461);
not I_10585 (I182885,I182868);
not I_10586 (I182902,I294488);
nand I_10587 (I182919,I294461,I294467);
nand I_10588 (I182936,I182919,I294488);
not I_10589 (I182953,I182936);
nor I_10590 (I182763,I182953,I182843);
nand I_10591 (I182984,I182919,I182902);
and I_10592 (I183001,I182984,I294473);
nand I_10593 (I183018,I183001,I294458);
and I_10594 (I183035,I183018,I182936);
nor I_10595 (I183052,I183018,I182936);
or I_10596 (I183069,I294485,I294467);
nor I_10597 (I183086,I183069,I294464);
not I_10598 (I183103,I183086);
nor I_10599 (I183120,I182885,I183103);
and I_10600 (I182754,I183120,I182851);
nor I_10601 (I183151,I182936,I183103);
nand I_10602 (I183168,I182953,I183086);
nand I_10603 (I183185,I294476,I294482);
nor I_10604 (I182751,I183185,I183086);
nor I_10605 (I183216,I183185,I183103);
not I_10606 (I183233,I183216);
nor I_10607 (I182775,I183035,I183233);
or I_10608 (I183264,I183185,I294458);
nand I_10609 (I183281,I183264,I183168);
not I_10610 (I183298,I183281);
nor I_10611 (I182757,I183298,I183151);
nor I_10612 (I183329,I183264,I183052);
DFFARX1 I_10613 (I183329,I2898,I182783,I182766,);
and I_10614 (I183360,I183018,I183264);
nor I_10615 (I182772,I183360,I182868);
nor I_10616 (I182769,I182851,I183360);
not I_10617 (I183405,I183185);
nand I_10618 (I183422,I183405,I183281);
nor I_10619 (I182760,I182885,I183422);
not I_10620 (I183480,I2905);
nand I_10621 (I183497,I265833,I265830);
and I_10622 (I183514,I183497,I265836);
DFFARX1 I_10623 (I183514,I2898,I183480,I183540,);
not I_10624 (I183548,I183540);
nor I_10625 (I183565,I265842,I265830);
not I_10626 (I183582,I183565);
not I_10627 (I183599,I265833);
nand I_10628 (I183616,I265830,I265839);
nand I_10629 (I183633,I183616,I265833);
not I_10630 (I183650,I183633);
nor I_10631 (I183460,I183650,I183540);
nand I_10632 (I183681,I183616,I183599);
and I_10633 (I183698,I183681,I265860);
nand I_10634 (I183715,I183698,I265848);
and I_10635 (I183732,I183715,I183633);
nor I_10636 (I183749,I183715,I183633);
or I_10637 (I183766,I265839,I265851);
nor I_10638 (I183783,I183766,I265845);
not I_10639 (I183800,I183783);
nor I_10640 (I183817,I183582,I183800);
and I_10641 (I183451,I183817,I183548);
nor I_10642 (I183848,I183633,I183800);
nand I_10643 (I183865,I183650,I183783);
nand I_10644 (I183882,I265854,I265857);
nor I_10645 (I183448,I183882,I183783);
nor I_10646 (I183913,I183882,I183800);
not I_10647 (I183930,I183913);
nor I_10648 (I183472,I183732,I183930);
or I_10649 (I183961,I183882,I265836);
nand I_10650 (I183978,I183961,I183865);
not I_10651 (I183995,I183978);
nor I_10652 (I183454,I183995,I183848);
nor I_10653 (I184026,I183961,I183749);
DFFARX1 I_10654 (I184026,I2898,I183480,I183463,);
and I_10655 (I184057,I183715,I183961);
nor I_10656 (I183469,I184057,I183565);
nor I_10657 (I183466,I183548,I184057);
not I_10658 (I184102,I183882);
nand I_10659 (I184119,I184102,I183978);
nor I_10660 (I183457,I183582,I184119);
not I_10661 (I184177,I2905);
nand I_10662 (I184194,I269658,I269655);
and I_10663 (I184211,I184194,I269661);
DFFARX1 I_10664 (I184211,I2898,I184177,I184237,);
not I_10665 (I184245,I184237);
nor I_10666 (I184262,I269667,I269655);
not I_10667 (I184279,I184262);
not I_10668 (I184296,I269658);
nand I_10669 (I184313,I269655,I269664);
nand I_10670 (I184330,I184313,I269658);
not I_10671 (I184347,I184330);
nor I_10672 (I184157,I184347,I184237);
nand I_10673 (I184378,I184313,I184296);
and I_10674 (I184395,I184378,I269685);
nand I_10675 (I184412,I184395,I269673);
and I_10676 (I184429,I184412,I184330);
nor I_10677 (I184446,I184412,I184330);
or I_10678 (I184463,I269664,I269676);
nor I_10679 (I184480,I184463,I269670);
not I_10680 (I184497,I184480);
nor I_10681 (I184514,I184279,I184497);
and I_10682 (I184148,I184514,I184245);
nor I_10683 (I184545,I184330,I184497);
nand I_10684 (I184562,I184347,I184480);
nand I_10685 (I184579,I269679,I269682);
nor I_10686 (I184145,I184579,I184480);
nor I_10687 (I184610,I184579,I184497);
not I_10688 (I184627,I184610);
nor I_10689 (I184169,I184429,I184627);
or I_10690 (I184658,I184579,I269661);
nand I_10691 (I184675,I184658,I184562);
not I_10692 (I184692,I184675);
nor I_10693 (I184151,I184692,I184545);
nor I_10694 (I184723,I184658,I184446);
DFFARX1 I_10695 (I184723,I2898,I184177,I184160,);
and I_10696 (I184754,I184412,I184658);
nor I_10697 (I184166,I184754,I184262);
nor I_10698 (I184163,I184245,I184754);
not I_10699 (I184799,I184579);
nand I_10700 (I184816,I184799,I184675);
nor I_10701 (I184154,I184279,I184816);
not I_10702 (I184874,I2905);
nand I_10703 (I184891,I428954,I428945);
and I_10704 (I184908,I184891,I428948);
DFFARX1 I_10705 (I184908,I2898,I184874,I184934,);
not I_10706 (I184942,I184934);
nor I_10707 (I184959,I428963,I428945);
not I_10708 (I184976,I184959);
not I_10709 (I184993,I428975);
nand I_10710 (I185010,I428972,I428966);
nand I_10711 (I185027,I185010,I428975);
not I_10712 (I185044,I185027);
nor I_10713 (I184854,I185044,I184934);
nand I_10714 (I185075,I185010,I184993);
and I_10715 (I185092,I185075,I428969);
nand I_10716 (I185109,I185092,I428951);
and I_10717 (I185126,I185109,I185027);
nor I_10718 (I185143,I185109,I185027);
or I_10719 (I185160,I428948,I428960);
nor I_10720 (I185177,I185160,I428957);
not I_10721 (I185194,I185177);
nor I_10722 (I185211,I184976,I185194);
and I_10723 (I184845,I185211,I184942);
nor I_10724 (I185242,I185027,I185194);
nand I_10725 (I185259,I185044,I185177);
nand I_10726 (I185276,I428951,I428978);
nor I_10727 (I184842,I185276,I185177);
nor I_10728 (I185307,I185276,I185194);
not I_10729 (I185324,I185307);
nor I_10730 (I184866,I185126,I185324);
or I_10731 (I185355,I185276,I428945);
nand I_10732 (I185372,I185355,I185259);
not I_10733 (I185389,I185372);
nor I_10734 (I184848,I185389,I185242);
nor I_10735 (I185420,I185355,I185143);
DFFARX1 I_10736 (I185420,I2898,I184874,I184857,);
and I_10737 (I185451,I185109,I185355);
nor I_10738 (I184863,I185451,I184959);
nor I_10739 (I184860,I184942,I185451);
not I_10740 (I185496,I185276);
nand I_10741 (I185513,I185496,I185372);
nor I_10742 (I184851,I184976,I185513);
not I_10743 (I185571,I2905);
nand I_10744 (I185588,I78320,I78338);
and I_10745 (I185605,I185588,I78332);
DFFARX1 I_10746 (I185605,I2898,I185571,I185631,);
not I_10747 (I185639,I185631);
nor I_10748 (I185656,I78326,I78338);
not I_10749 (I185673,I185656);
not I_10750 (I185690,I78344);
nand I_10751 (I185707,I78320,I78341);
nand I_10752 (I185724,I185707,I78344);
not I_10753 (I185741,I185724);
nor I_10754 (I185551,I185741,I185631);
nand I_10755 (I185772,I185707,I185690);
and I_10756 (I185789,I185772,I78329);
nand I_10757 (I185806,I185789,I78329);
and I_10758 (I185823,I185806,I185724);
nor I_10759 (I185840,I185806,I185724);
or I_10760 (I185857,I78323,I78326);
nor I_10761 (I185874,I185857,I78332);
not I_10762 (I185891,I185874);
nor I_10763 (I185908,I185673,I185891);
and I_10764 (I185542,I185908,I185639);
nor I_10765 (I185939,I185724,I185891);
nand I_10766 (I185956,I185741,I185874);
nand I_10767 (I185973,I78335,I78347);
nor I_10768 (I185539,I185973,I185874);
nor I_10769 (I186004,I185973,I185891);
not I_10770 (I186021,I186004);
nor I_10771 (I185563,I185823,I186021);
or I_10772 (I186052,I185973,I78323);
nand I_10773 (I186069,I186052,I185956);
not I_10774 (I186086,I186069);
nor I_10775 (I185545,I186086,I185939);
nor I_10776 (I186117,I186052,I185840);
DFFARX1 I_10777 (I186117,I2898,I185571,I185554,);
and I_10778 (I186148,I185806,I186052);
nor I_10779 (I185560,I186148,I185656);
nor I_10780 (I185557,I185639,I186148);
not I_10781 (I186193,I185973);
nand I_10782 (I186210,I186193,I186069);
nor I_10783 (I185548,I185673,I186210);
not I_10784 (I186268,I2905);
nand I_10785 (I186285,I1907,I2683);
and I_10786 (I186302,I186285,I2851);
DFFARX1 I_10787 (I186302,I2898,I186268,I186328,);
not I_10788 (I186336,I186328);
nor I_10789 (I186353,I2027,I2683);
not I_10790 (I186370,I186353);
not I_10791 (I186387,I2067);
nand I_10792 (I186404,I2555,I1827);
nand I_10793 (I186421,I186404,I2067);
not I_10794 (I186438,I186421);
nor I_10795 (I186248,I186438,I186328);
nand I_10796 (I186469,I186404,I186387);
and I_10797 (I186486,I186469,I2795);
nand I_10798 (I186503,I186486,I2595);
and I_10799 (I186520,I186503,I186421);
nor I_10800 (I186537,I186503,I186421);
or I_10801 (I186554,I2155,I2835);
nor I_10802 (I186571,I186554,I2891);
not I_10803 (I186588,I186571);
nor I_10804 (I186605,I186370,I186588);
and I_10805 (I186239,I186605,I186336);
nor I_10806 (I186636,I186421,I186588);
nand I_10807 (I186653,I186438,I186571);
nand I_10808 (I186670,I2771,I1699);
nor I_10809 (I186236,I186670,I186571);
nor I_10810 (I186701,I186670,I186588);
not I_10811 (I186718,I186701);
nor I_10812 (I186260,I186520,I186718);
or I_10813 (I186749,I186670,I2235);
nand I_10814 (I186766,I186749,I186653);
not I_10815 (I186783,I186766);
nor I_10816 (I186242,I186783,I186636);
nor I_10817 (I186814,I186749,I186537);
DFFARX1 I_10818 (I186814,I2898,I186268,I186251,);
and I_10819 (I186845,I186503,I186749);
nor I_10820 (I186257,I186845,I186353);
nor I_10821 (I186254,I186336,I186845);
not I_10822 (I186890,I186670);
nand I_10823 (I186907,I186890,I186766);
nor I_10824 (I186245,I186370,I186907);
not I_10825 (I186965,I2905);
nand I_10826 (I186982,I255123,I255120);
and I_10827 (I186999,I186982,I255126);
DFFARX1 I_10828 (I186999,I2898,I186965,I187025,);
not I_10829 (I187033,I187025);
nor I_10830 (I187050,I255132,I255120);
not I_10831 (I187067,I187050);
not I_10832 (I187084,I255123);
nand I_10833 (I187101,I255120,I255129);
nand I_10834 (I187118,I187101,I255123);
not I_10835 (I187135,I187118);
nor I_10836 (I186945,I187135,I187025);
nand I_10837 (I187166,I187101,I187084);
and I_10838 (I187183,I187166,I255150);
nand I_10839 (I187200,I187183,I255138);
and I_10840 (I187217,I187200,I187118);
nor I_10841 (I187234,I187200,I187118);
or I_10842 (I187251,I255129,I255141);
nor I_10843 (I187268,I187251,I255135);
not I_10844 (I187285,I187268);
nor I_10845 (I187302,I187067,I187285);
and I_10846 (I186936,I187302,I187033);
nor I_10847 (I187333,I187118,I187285);
nand I_10848 (I187350,I187135,I187268);
nand I_10849 (I187367,I255144,I255147);
nor I_10850 (I186933,I187367,I187268);
nor I_10851 (I187398,I187367,I187285);
not I_10852 (I187415,I187398);
nor I_10853 (I186957,I187217,I187415);
or I_10854 (I187446,I187367,I255126);
nand I_10855 (I187463,I187446,I187350);
not I_10856 (I187480,I187463);
nor I_10857 (I186939,I187480,I187333);
nor I_10858 (I187511,I187446,I187234);
DFFARX1 I_10859 (I187511,I2898,I186965,I186948,);
and I_10860 (I187542,I187200,I187446);
nor I_10861 (I186954,I187542,I187050);
nor I_10862 (I186951,I187033,I187542);
not I_10863 (I187587,I187367);
nand I_10864 (I187604,I187587,I187463);
nor I_10865 (I186942,I187067,I187604);
not I_10866 (I187662,I2905);
nand I_10867 (I187679,I69514,I69532);
and I_10868 (I187696,I187679,I69526);
DFFARX1 I_10869 (I187696,I2898,I187662,I187722,);
not I_10870 (I187730,I187722);
nor I_10871 (I187747,I69520,I69532);
not I_10872 (I187764,I187747);
not I_10873 (I187781,I69538);
nand I_10874 (I187798,I69514,I69535);
nand I_10875 (I187815,I187798,I69538);
not I_10876 (I187832,I187815);
nor I_10877 (I187642,I187832,I187722);
nand I_10878 (I187863,I187798,I187781);
and I_10879 (I187880,I187863,I69523);
nand I_10880 (I187897,I187880,I69523);
and I_10881 (I187914,I187897,I187815);
nor I_10882 (I187931,I187897,I187815);
or I_10883 (I187948,I69517,I69520);
nor I_10884 (I187965,I187948,I69526);
not I_10885 (I187982,I187965);
nor I_10886 (I187999,I187764,I187982);
and I_10887 (I187633,I187999,I187730);
nor I_10888 (I188030,I187815,I187982);
nand I_10889 (I188047,I187832,I187965);
nand I_10890 (I188064,I69529,I69541);
nor I_10891 (I187630,I188064,I187965);
nor I_10892 (I188095,I188064,I187982);
not I_10893 (I188112,I188095);
nor I_10894 (I187654,I187914,I188112);
or I_10895 (I188143,I188064,I69517);
nand I_10896 (I188160,I188143,I188047);
not I_10897 (I188177,I188160);
nor I_10898 (I187636,I188177,I188030);
nor I_10899 (I188208,I188143,I187931);
DFFARX1 I_10900 (I188208,I2898,I187662,I187645,);
and I_10901 (I188239,I187897,I188143);
nor I_10902 (I187651,I188239,I187747);
nor I_10903 (I187648,I187730,I188239);
not I_10904 (I188284,I188064);
nand I_10905 (I188301,I188284,I188160);
nor I_10906 (I187639,I187764,I188301);
not I_10907 (I188359,I2905);
nand I_10908 (I188376,I213463,I213436);
and I_10909 (I188393,I188376,I213448);
DFFARX1 I_10910 (I188393,I2898,I188359,I188419,);
not I_10911 (I188427,I188419);
nor I_10912 (I188444,I213454,I213436);
not I_10913 (I188461,I188444);
not I_10914 (I188478,I213451);
nand I_10915 (I188495,I213445,I213448);
nand I_10916 (I188512,I188495,I213451);
not I_10917 (I188529,I188512);
nor I_10918 (I188339,I188529,I188419);
nand I_10919 (I188560,I188495,I188478);
and I_10920 (I188577,I188560,I213460);
nand I_10921 (I188594,I188577,I213439);
and I_10922 (I188611,I188594,I188512);
nor I_10923 (I188628,I188594,I188512);
or I_10924 (I188645,I213436,I213457);
nor I_10925 (I188662,I188645,I213442);
not I_10926 (I188679,I188662);
nor I_10927 (I188696,I188461,I188679);
and I_10928 (I188330,I188696,I188427);
nor I_10929 (I188727,I188512,I188679);
nand I_10930 (I188744,I188529,I188662);
nand I_10931 (I188761,I213439,I213445);
nor I_10932 (I188327,I188761,I188662);
nor I_10933 (I188792,I188761,I188679);
not I_10934 (I188809,I188792);
nor I_10935 (I188351,I188611,I188809);
or I_10936 (I188840,I188761,I213442);
nand I_10937 (I188857,I188840,I188744);
not I_10938 (I188874,I188857);
nor I_10939 (I188333,I188874,I188727);
nor I_10940 (I188905,I188840,I188628);
DFFARX1 I_10941 (I188905,I2898,I188359,I188342,);
and I_10942 (I188936,I188594,I188840);
nor I_10943 (I188348,I188936,I188444);
nor I_10944 (I188345,I188427,I188936);
not I_10945 (I188981,I188761);
nand I_10946 (I188998,I188981,I188857);
nor I_10947 (I188336,I188461,I188998);
not I_10948 (I189056,I2905);
nand I_10949 (I189073,I275013,I275010);
and I_10950 (I189090,I189073,I275016);
DFFARX1 I_10951 (I189090,I2898,I189056,I189116,);
not I_10952 (I189124,I189116);
nor I_10953 (I189141,I275022,I275010);
not I_10954 (I189158,I189141);
not I_10955 (I189175,I275013);
nand I_10956 (I189192,I275010,I275019);
nand I_10957 (I189209,I189192,I275013);
not I_10958 (I189226,I189209);
nor I_10959 (I189036,I189226,I189116);
nand I_10960 (I189257,I189192,I189175);
and I_10961 (I189274,I189257,I275040);
nand I_10962 (I189291,I189274,I275028);
and I_10963 (I189308,I189291,I189209);
nor I_10964 (I189325,I189291,I189209);
or I_10965 (I189342,I275019,I275031);
nor I_10966 (I189359,I189342,I275025);
not I_10967 (I189376,I189359);
nor I_10968 (I189393,I189158,I189376);
and I_10969 (I189027,I189393,I189124);
nor I_10970 (I189424,I189209,I189376);
nand I_10971 (I189441,I189226,I189359);
nand I_10972 (I189458,I275034,I275037);
nor I_10973 (I189024,I189458,I189359);
nor I_10974 (I189489,I189458,I189376);
not I_10975 (I189506,I189489);
nor I_10976 (I189048,I189308,I189506);
or I_10977 (I189537,I189458,I275016);
nand I_10978 (I189554,I189537,I189441);
not I_10979 (I189571,I189554);
nor I_10980 (I189030,I189571,I189424);
nor I_10981 (I189602,I189537,I189325);
DFFARX1 I_10982 (I189602,I2898,I189056,I189039,);
and I_10983 (I189633,I189291,I189537);
nor I_10984 (I189045,I189633,I189141);
nor I_10985 (I189042,I189124,I189633);
not I_10986 (I189678,I189458);
nand I_10987 (I189695,I189678,I189554);
nor I_10988 (I189033,I189158,I189695);
not I_10989 (I189753,I2905);
nand I_10990 (I189770,I316409,I316391);
and I_10991 (I189787,I189770,I316400);
DFFARX1 I_10992 (I189787,I2898,I189753,I189813,);
not I_10993 (I189821,I189813);
nor I_10994 (I189838,I316394,I316391);
not I_10995 (I189855,I189838);
not I_10996 (I189872,I316418);
nand I_10997 (I189889,I316391,I316397);
nand I_10998 (I189906,I189889,I316418);
not I_10999 (I189923,I189906);
nor I_11000 (I189733,I189923,I189813);
nand I_11001 (I189954,I189889,I189872);
and I_11002 (I189971,I189954,I316403);
nand I_11003 (I189988,I189971,I316388);
and I_11004 (I190005,I189988,I189906);
nor I_11005 (I190022,I189988,I189906);
or I_11006 (I190039,I316415,I316397);
nor I_11007 (I190056,I190039,I316394);
not I_11008 (I190073,I190056);
nor I_11009 (I190090,I189855,I190073);
and I_11010 (I189724,I190090,I189821);
nor I_11011 (I190121,I189906,I190073);
nand I_11012 (I190138,I189923,I190056);
nand I_11013 (I190155,I316406,I316412);
nor I_11014 (I189721,I190155,I190056);
nor I_11015 (I190186,I190155,I190073);
not I_11016 (I190203,I190186);
nor I_11017 (I189745,I190005,I190203);
or I_11018 (I190234,I190155,I316388);
nand I_11019 (I190251,I190234,I190138);
not I_11020 (I190268,I190251);
nor I_11021 (I189727,I190268,I190121);
nor I_11022 (I190299,I190234,I190022);
DFFARX1 I_11023 (I190299,I2898,I189753,I189736,);
and I_11024 (I190330,I189988,I190234);
nor I_11025 (I189742,I190330,I189838);
nor I_11026 (I189739,I189821,I190330);
not I_11027 (I190375,I190155);
nand I_11028 (I190392,I190375,I190251);
nor I_11029 (I189730,I189855,I190392);
not I_11030 (I190450,I2905);
nand I_11031 (I190467,I156554,I156584);
and I_11032 (I190484,I190467,I156560);
DFFARX1 I_11033 (I190484,I2898,I190450,I190510,);
not I_11034 (I190518,I190510);
nor I_11035 (I190535,I156563,I156584);
not I_11036 (I190552,I190535);
not I_11037 (I190569,I156569);
nand I_11038 (I190586,I156575,I156557);
nand I_11039 (I190603,I190586,I156569);
not I_11040 (I190620,I190603);
nor I_11041 (I190430,I190620,I190510);
nand I_11042 (I190651,I190586,I190569);
and I_11043 (I190668,I190651,I156572);
nand I_11044 (I190685,I190668,I156554);
and I_11045 (I190702,I190685,I190603);
nor I_11046 (I190719,I190685,I190603);
or I_11047 (I190736,I156560,I156581);
nor I_11048 (I190753,I190736,I156566);
not I_11049 (I190770,I190753);
nor I_11050 (I190787,I190552,I190770);
and I_11051 (I190421,I190787,I190518);
nor I_11052 (I190818,I190603,I190770);
nand I_11053 (I190835,I190620,I190753);
nand I_11054 (I190852,I156578,I156557);
nor I_11055 (I190418,I190852,I190753);
nor I_11056 (I190883,I190852,I190770);
not I_11057 (I190900,I190883);
nor I_11058 (I190442,I190702,I190900);
or I_11059 (I190931,I190852,I156587);
nand I_11060 (I190948,I190931,I190835);
not I_11061 (I190965,I190948);
nor I_11062 (I190424,I190965,I190818);
nor I_11063 (I190996,I190931,I190719);
DFFARX1 I_11064 (I190996,I2898,I190450,I190433,);
and I_11065 (I191027,I190685,I190931);
nor I_11066 (I190439,I191027,I190535);
nor I_11067 (I190436,I190518,I191027);
not I_11068 (I191072,I190852);
nand I_11069 (I191089,I191072,I190948);
nor I_11070 (I190427,I190552,I191089);
not I_11071 (I191147,I2905);
nand I_11072 (I191164,I233703,I233700);
and I_11073 (I191181,I191164,I233706);
DFFARX1 I_11074 (I191181,I2898,I191147,I191207,);
not I_11075 (I191215,I191207);
nor I_11076 (I191232,I233712,I233700);
not I_11077 (I191249,I191232);
not I_11078 (I191266,I233703);
nand I_11079 (I191283,I233700,I233709);
nand I_11080 (I191300,I191283,I233703);
not I_11081 (I191317,I191300);
nor I_11082 (I191127,I191317,I191207);
nand I_11083 (I191348,I191283,I191266);
and I_11084 (I191365,I191348,I233730);
nand I_11085 (I191382,I191365,I233718);
and I_11086 (I191399,I191382,I191300);
nor I_11087 (I191416,I191382,I191300);
or I_11088 (I191433,I233709,I233721);
nor I_11089 (I191450,I191433,I233715);
not I_11090 (I191467,I191450);
nor I_11091 (I191484,I191249,I191467);
and I_11092 (I191118,I191484,I191215);
nor I_11093 (I191515,I191300,I191467);
nand I_11094 (I191532,I191317,I191450);
nand I_11095 (I191549,I233724,I233727);
nor I_11096 (I191115,I191549,I191450);
nor I_11097 (I191580,I191549,I191467);
not I_11098 (I191597,I191580);
nor I_11099 (I191139,I191399,I191597);
or I_11100 (I191628,I191549,I233706);
nand I_11101 (I191645,I191628,I191532);
not I_11102 (I191662,I191645);
nor I_11103 (I191121,I191662,I191515);
nor I_11104 (I191693,I191628,I191416);
DFFARX1 I_11105 (I191693,I2898,I191147,I191130,);
and I_11106 (I191724,I191382,I191628);
nor I_11107 (I191136,I191724,I191232);
nor I_11108 (I191133,I191215,I191724);
not I_11109 (I191769,I191549);
nand I_11110 (I191786,I191769,I191645);
nor I_11111 (I191124,I191249,I191786);
not I_11112 (I191844,I2905);
nand I_11113 (I191861,I350201,I350213);
and I_11114 (I191878,I191861,I350204);
DFFARX1 I_11115 (I191878,I2898,I191844,I191904,);
not I_11116 (I191912,I191904);
nor I_11117 (I191929,I350216,I350213);
not I_11118 (I191946,I191929);
not I_11119 (I191963,I350222);
nand I_11120 (I191980,I350207,I350210);
nand I_11121 (I191997,I191980,I350222);
not I_11122 (I192014,I191997);
nor I_11123 (I191824,I192014,I191904);
nand I_11124 (I192045,I191980,I191963);
and I_11125 (I192062,I192045,I350219);
nand I_11126 (I192079,I192062,I350207);
and I_11127 (I192096,I192079,I191997);
nor I_11128 (I192113,I192079,I191997);
or I_11129 (I192130,I350225,I350210);
nor I_11130 (I192147,I192130,I350216);
not I_11131 (I192164,I192147);
nor I_11132 (I192181,I191946,I192164);
and I_11133 (I191815,I192181,I191912);
nor I_11134 (I192212,I191997,I192164);
nand I_11135 (I192229,I192014,I192147);
nand I_11136 (I192246,I350201,I350213);
nor I_11137 (I191812,I192246,I192147);
nor I_11138 (I192277,I192246,I192164);
not I_11139 (I192294,I192277);
nor I_11140 (I191836,I192096,I192294);
or I_11141 (I192325,I192246,I350204);
nand I_11142 (I192342,I192325,I192229);
not I_11143 (I192359,I192342);
nor I_11144 (I191818,I192359,I192212);
nor I_11145 (I192390,I192325,I192113);
DFFARX1 I_11146 (I192390,I2898,I191844,I191827,);
and I_11147 (I192421,I192079,I192325);
nor I_11148 (I191833,I192421,I191929);
nor I_11149 (I191830,I191912,I192421);
not I_11150 (I192466,I192246);
nand I_11151 (I192483,I192466,I192342);
nor I_11152 (I191821,I191946,I192483);
not I_11153 (I192541,I2905);
nand I_11154 (I192558,I109743,I109737);
and I_11155 (I192575,I192558,I109728);
DFFARX1 I_11156 (I192575,I2898,I192541,I192601,);
not I_11157 (I192609,I192601);
nor I_11158 (I192626,I109731,I109737);
not I_11159 (I192643,I192626);
not I_11160 (I192660,I109746);
nand I_11161 (I192677,I109722,I109719);
nand I_11162 (I192694,I192677,I109746);
not I_11163 (I192711,I192694);
nor I_11164 (I192521,I192711,I192601);
nand I_11165 (I192742,I192677,I192660);
and I_11166 (I192759,I192742,I109734);
nand I_11167 (I192776,I192759,I109719);
and I_11168 (I192793,I192776,I192694);
nor I_11169 (I192810,I192776,I192694);
or I_11170 (I192827,I109725,I109725);
nor I_11171 (I192844,I192827,I109752);
not I_11172 (I192861,I192844);
nor I_11173 (I192878,I192643,I192861);
and I_11174 (I192512,I192878,I192609);
nor I_11175 (I192909,I192694,I192861);
nand I_11176 (I192926,I192711,I192844);
nand I_11177 (I192943,I109740,I109749);
nor I_11178 (I192509,I192943,I192844);
nor I_11179 (I192974,I192943,I192861);
not I_11180 (I192991,I192974);
nor I_11181 (I192533,I192793,I192991);
or I_11182 (I193022,I192943,I109722);
nand I_11183 (I193039,I193022,I192926);
not I_11184 (I193056,I193039);
nor I_11185 (I192515,I193056,I192909);
nor I_11186 (I193087,I193022,I192810);
DFFARX1 I_11187 (I193087,I2898,I192541,I192524,);
and I_11188 (I193118,I192776,I193022);
nor I_11189 (I192530,I193118,I192626);
nor I_11190 (I192527,I192609,I193118);
not I_11191 (I193163,I192943);
nand I_11192 (I193180,I193163,I193039);
nor I_11193 (I192518,I192643,I193180);
not I_11194 (I193238,I2905);
nand I_11195 (I193255,I220195,I220168);
and I_11196 (I193272,I193255,I220180);
DFFARX1 I_11197 (I193272,I2898,I193238,I193298,);
not I_11198 (I193306,I193298);
nor I_11199 (I193323,I220186,I220168);
not I_11200 (I193340,I193323);
not I_11201 (I193357,I220183);
nand I_11202 (I193374,I220177,I220180);
nand I_11203 (I193391,I193374,I220183);
not I_11204 (I193408,I193391);
nor I_11205 (I193218,I193408,I193298);
nand I_11206 (I193439,I193374,I193357);
and I_11207 (I193456,I193439,I220192);
nand I_11208 (I193473,I193456,I220171);
and I_11209 (I193490,I193473,I193391);
nor I_11210 (I193507,I193473,I193391);
or I_11211 (I193524,I220168,I220189);
nor I_11212 (I193541,I193524,I220174);
not I_11213 (I193558,I193541);
nor I_11214 (I193575,I193340,I193558);
and I_11215 (I193209,I193575,I193306);
nor I_11216 (I193606,I193391,I193558);
nand I_11217 (I193623,I193408,I193541);
nand I_11218 (I193640,I220171,I220177);
nor I_11219 (I193206,I193640,I193541);
nor I_11220 (I193671,I193640,I193558);
not I_11221 (I193688,I193671);
nor I_11222 (I193230,I193490,I193688);
or I_11223 (I193719,I193640,I220174);
nand I_11224 (I193736,I193719,I193623);
not I_11225 (I193753,I193736);
nor I_11226 (I193212,I193753,I193606);
nor I_11227 (I193784,I193719,I193507);
DFFARX1 I_11228 (I193784,I2898,I193238,I193221,);
and I_11229 (I193815,I193473,I193719);
nor I_11230 (I193227,I193815,I193323);
nor I_11231 (I193224,I193306,I193815);
not I_11232 (I193860,I193640);
nand I_11233 (I193877,I193860,I193736);
nor I_11234 (I193215,I193340,I193877);
not I_11235 (I193935,I2905);
nand I_11236 (I193952,I362101,I362113);
and I_11237 (I193969,I193952,I362104);
DFFARX1 I_11238 (I193969,I2898,I193935,I193995,);
not I_11239 (I194003,I193995);
nor I_11240 (I194020,I362116,I362113);
not I_11241 (I194037,I194020);
not I_11242 (I194054,I362122);
nand I_11243 (I194071,I362107,I362110);
nand I_11244 (I194088,I194071,I362122);
not I_11245 (I194105,I194088);
nor I_11246 (I193915,I194105,I193995);
nand I_11247 (I194136,I194071,I194054);
and I_11248 (I194153,I194136,I362119);
nand I_11249 (I194170,I194153,I362107);
and I_11250 (I194187,I194170,I194088);
nor I_11251 (I194204,I194170,I194088);
or I_11252 (I194221,I362125,I362110);
nor I_11253 (I194238,I194221,I362116);
not I_11254 (I194255,I194238);
nor I_11255 (I194272,I194037,I194255);
and I_11256 (I193906,I194272,I194003);
nor I_11257 (I194303,I194088,I194255);
nand I_11258 (I194320,I194105,I194238);
nand I_11259 (I194337,I362101,I362113);
nor I_11260 (I193903,I194337,I194238);
nor I_11261 (I194368,I194337,I194255);
not I_11262 (I194385,I194368);
nor I_11263 (I193927,I194187,I194385);
or I_11264 (I194416,I194337,I362104);
nand I_11265 (I194433,I194416,I194320);
not I_11266 (I194450,I194433);
nor I_11267 (I193909,I194450,I194303);
nor I_11268 (I194481,I194416,I194204);
DFFARX1 I_11269 (I194481,I2898,I193935,I193918,);
and I_11270 (I194512,I194170,I194416);
nor I_11271 (I193924,I194512,I194020);
nor I_11272 (I193921,I194003,I194512);
not I_11273 (I194557,I194337);
nand I_11274 (I194574,I194557,I194433);
nor I_11275 (I193912,I194037,I194574);
not I_11276 (I194632,I2905);
nand I_11277 (I194649,I343061,I343073);
and I_11278 (I194666,I194649,I343064);
DFFARX1 I_11279 (I194666,I2898,I194632,I194692,);
not I_11280 (I194700,I194692);
nor I_11281 (I194717,I343076,I343073);
not I_11282 (I194734,I194717);
not I_11283 (I194751,I343082);
nand I_11284 (I194768,I343067,I343070);
nand I_11285 (I194785,I194768,I343082);
not I_11286 (I194802,I194785);
nor I_11287 (I194612,I194802,I194692);
nand I_11288 (I194833,I194768,I194751);
and I_11289 (I194850,I194833,I343079);
nand I_11290 (I194867,I194850,I343067);
and I_11291 (I194884,I194867,I194785);
nor I_11292 (I194901,I194867,I194785);
or I_11293 (I194918,I343085,I343070);
nor I_11294 (I194935,I194918,I343076);
not I_11295 (I194952,I194935);
nor I_11296 (I194969,I194734,I194952);
and I_11297 (I194603,I194969,I194700);
nor I_11298 (I195000,I194785,I194952);
nand I_11299 (I195017,I194802,I194935);
nand I_11300 (I195034,I343061,I343073);
nor I_11301 (I194600,I195034,I194935);
nor I_11302 (I195065,I195034,I194952);
not I_11303 (I195082,I195065);
nor I_11304 (I194624,I194884,I195082);
or I_11305 (I195113,I195034,I343064);
nand I_11306 (I195130,I195113,I195017);
not I_11307 (I195147,I195130);
nor I_11308 (I194606,I195147,I195000);
nor I_11309 (I195178,I195113,I194901);
DFFARX1 I_11310 (I195178,I2898,I194632,I194615,);
and I_11311 (I195209,I194867,I195113);
nor I_11312 (I194621,I195209,I194717);
nor I_11313 (I194618,I194700,I195209);
not I_11314 (I195254,I195034);
nand I_11315 (I195271,I195254,I195130);
nor I_11316 (I194609,I194734,I195271);
not I_11317 (I195329,I2905);
nand I_11318 (I195346,I284976,I284958);
and I_11319 (I195363,I195346,I284967);
DFFARX1 I_11320 (I195363,I2898,I195329,I195389,);
not I_11321 (I195397,I195389);
nor I_11322 (I195414,I284961,I284958);
not I_11323 (I195431,I195414);
not I_11324 (I195448,I284985);
nand I_11325 (I195465,I284958,I284964);
nand I_11326 (I195482,I195465,I284985);
not I_11327 (I195499,I195482);
nor I_11328 (I195309,I195499,I195389);
nand I_11329 (I195530,I195465,I195448);
and I_11330 (I195547,I195530,I284970);
nand I_11331 (I195564,I195547,I284955);
and I_11332 (I195581,I195564,I195482);
nor I_11333 (I195598,I195564,I195482);
or I_11334 (I195615,I284982,I284964);
nor I_11335 (I195632,I195615,I284961);
not I_11336 (I195649,I195632);
nor I_11337 (I195666,I195431,I195649);
and I_11338 (I195300,I195666,I195397);
nor I_11339 (I195697,I195482,I195649);
nand I_11340 (I195714,I195499,I195632);
nand I_11341 (I195731,I284973,I284979);
nor I_11342 (I195297,I195731,I195632);
nor I_11343 (I195762,I195731,I195649);
not I_11344 (I195779,I195762);
nor I_11345 (I195321,I195581,I195779);
or I_11346 (I195810,I195731,I284955);
nand I_11347 (I195827,I195810,I195714);
not I_11348 (I195844,I195827);
nor I_11349 (I195303,I195844,I195697);
nor I_11350 (I195875,I195810,I195598);
DFFARX1 I_11351 (I195875,I2898,I195329,I195312,);
and I_11352 (I195906,I195564,I195810);
nor I_11353 (I195318,I195906,I195414);
nor I_11354 (I195315,I195397,I195906);
not I_11355 (I195951,I195731);
nand I_11356 (I195968,I195951,I195827);
nor I_11357 (I195306,I195431,I195968);
not I_11358 (I196026,I2905);
nand I_11359 (I196043,I314947,I314929);
and I_11360 (I196060,I196043,I314938);
DFFARX1 I_11361 (I196060,I2898,I196026,I196086,);
not I_11362 (I196094,I196086);
nor I_11363 (I196111,I314932,I314929);
not I_11364 (I196128,I196111);
not I_11365 (I196145,I314956);
nand I_11366 (I196162,I314929,I314935);
nand I_11367 (I196179,I196162,I314956);
not I_11368 (I196196,I196179);
nor I_11369 (I196006,I196196,I196086);
nand I_11370 (I196227,I196162,I196145);
and I_11371 (I196244,I196227,I314941);
nand I_11372 (I196261,I196244,I314926);
and I_11373 (I196278,I196261,I196179);
nor I_11374 (I196295,I196261,I196179);
or I_11375 (I196312,I314953,I314935);
nor I_11376 (I196329,I196312,I314932);
not I_11377 (I196346,I196329);
nor I_11378 (I196363,I196128,I196346);
and I_11379 (I195997,I196363,I196094);
nor I_11380 (I196394,I196179,I196346);
nand I_11381 (I196411,I196196,I196329);
nand I_11382 (I196428,I314944,I314950);
nor I_11383 (I195994,I196428,I196329);
nor I_11384 (I196459,I196428,I196346);
not I_11385 (I196476,I196459);
nor I_11386 (I196018,I196278,I196476);
or I_11387 (I196507,I196428,I314926);
nand I_11388 (I196524,I196507,I196411);
not I_11389 (I196541,I196524);
nor I_11390 (I196000,I196541,I196394);
nor I_11391 (I196572,I196507,I196295);
DFFARX1 I_11392 (I196572,I2898,I196026,I196009,);
and I_11393 (I196603,I196261,I196507);
nor I_11394 (I196015,I196603,I196111);
nor I_11395 (I196012,I196094,I196603);
not I_11396 (I196648,I196428);
nand I_11397 (I196665,I196648,I196524);
nor I_11398 (I196003,I196128,I196665);
not I_11399 (I196723,I2905);
nand I_11400 (I196740,I30352,I30367);
and I_11401 (I196757,I196740,I30361);
DFFARX1 I_11402 (I196757,I2898,I196723,I196783,);
not I_11403 (I196791,I196783);
nor I_11404 (I196808,I30373,I30367);
not I_11405 (I196825,I196808);
not I_11406 (I196842,I30355);
nand I_11407 (I196859,I30364,I30352);
nand I_11408 (I196876,I196859,I30355);
not I_11409 (I196893,I196876);
nor I_11410 (I196703,I196893,I196783);
nand I_11411 (I196924,I196859,I196842);
and I_11412 (I196941,I196924,I30355);
nand I_11413 (I196958,I196941,I30349);
and I_11414 (I196975,I196958,I196876);
nor I_11415 (I196992,I196958,I196876);
or I_11416 (I197009,I30349,I30370);
nor I_11417 (I197026,I197009,I30346);
not I_11418 (I197043,I197026);
nor I_11419 (I197060,I196825,I197043);
and I_11420 (I196694,I197060,I196791);
nor I_11421 (I197091,I196876,I197043);
nand I_11422 (I197108,I196893,I197026);
nand I_11423 (I197125,I30358,I30358);
nor I_11424 (I196691,I197125,I197026);
nor I_11425 (I197156,I197125,I197043);
not I_11426 (I197173,I197156);
nor I_11427 (I196715,I196975,I197173);
or I_11428 (I197204,I197125,I30346);
nand I_11429 (I197221,I197204,I197108);
not I_11430 (I197238,I197221);
nor I_11431 (I196697,I197238,I197091);
nor I_11432 (I197269,I197204,I196992);
DFFARX1 I_11433 (I197269,I2898,I196723,I196706,);
and I_11434 (I197300,I196958,I197204);
nor I_11435 (I196712,I197300,I196808);
nor I_11436 (I196709,I196791,I197300);
not I_11437 (I197345,I197125);
nand I_11438 (I197362,I197345,I197221);
nor I_11439 (I196700,I196825,I197362);
not I_11440 (I197420,I2905);
nand I_11441 (I197437,I55855,I55876);
and I_11442 (I197454,I197437,I55873);
DFFARX1 I_11443 (I197454,I2898,I197420,I197480,);
not I_11444 (I197488,I197480);
nor I_11445 (I197505,I55852,I55876);
not I_11446 (I197522,I197505);
not I_11447 (I197539,I55858);
nand I_11448 (I197556,I55879,I55870);
nand I_11449 (I197573,I197556,I55858);
not I_11450 (I197590,I197573);
nor I_11451 (I197400,I197590,I197480);
nand I_11452 (I197621,I197556,I197539);
and I_11453 (I197638,I197621,I55882);
nand I_11454 (I197655,I197638,I55849);
and I_11455 (I197672,I197655,I197573);
nor I_11456 (I197689,I197655,I197573);
or I_11457 (I197706,I55846,I55861);
nor I_11458 (I197723,I197706,I55846);
not I_11459 (I197740,I197723);
nor I_11460 (I197757,I197522,I197740);
and I_11461 (I197391,I197757,I197488);
nor I_11462 (I197788,I197573,I197740);
nand I_11463 (I197805,I197590,I197723);
nand I_11464 (I197822,I55867,I55864);
nor I_11465 (I197388,I197822,I197723);
nor I_11466 (I197853,I197822,I197740);
not I_11467 (I197870,I197853);
nor I_11468 (I197412,I197672,I197870);
or I_11469 (I197901,I197822,I55849);
nand I_11470 (I197918,I197901,I197805);
not I_11471 (I197935,I197918);
nor I_11472 (I197394,I197935,I197788);
nor I_11473 (I197966,I197901,I197689);
DFFARX1 I_11474 (I197966,I2898,I197420,I197403,);
and I_11475 (I197997,I197655,I197901);
nor I_11476 (I197409,I197997,I197505);
nor I_11477 (I197406,I197488,I197997);
not I_11478 (I198042,I197822);
nand I_11479 (I198059,I198042,I197918);
nor I_11480 (I197397,I197522,I198059);
not I_11481 (I198117,I2905);
nand I_11482 (I198134,I369683,I369695);
and I_11483 (I198151,I198134,I369689);
DFFARX1 I_11484 (I198151,I2898,I198117,I198177,);
not I_11485 (I198185,I198177);
nor I_11486 (I198202,I369683,I369695);
not I_11487 (I198219,I198202);
not I_11488 (I198236,I369704);
nand I_11489 (I198253,I369692,I369713);
nand I_11490 (I198270,I198253,I369704);
not I_11491 (I198287,I198270);
nor I_11492 (I198097,I198287,I198177);
nand I_11493 (I198318,I198253,I198236);
and I_11494 (I198335,I198318,I369698);
nand I_11495 (I198352,I198335,I369707);
and I_11496 (I198369,I198352,I198270);
nor I_11497 (I198386,I198352,I198270);
or I_11498 (I198403,I369716,I369710);
nor I_11499 (I198420,I198403,I369686);
not I_11500 (I198437,I198420);
nor I_11501 (I198454,I198219,I198437);
and I_11502 (I198088,I198454,I198185);
nor I_11503 (I198485,I198270,I198437);
nand I_11504 (I198502,I198287,I198420);
nand I_11505 (I198519,I369689,I369701);
nor I_11506 (I198085,I198519,I198420);
nor I_11507 (I198550,I198519,I198437);
not I_11508 (I198567,I198550);
nor I_11509 (I198109,I198369,I198567);
or I_11510 (I198598,I198519,I369686);
nand I_11511 (I198615,I198598,I198502);
not I_11512 (I198632,I198615);
nor I_11513 (I198091,I198632,I198485);
nor I_11514 (I198663,I198598,I198386);
DFFARX1 I_11515 (I198663,I2898,I198117,I198100,);
and I_11516 (I198694,I198352,I198598);
nor I_11517 (I198106,I198694,I198202);
nor I_11518 (I198103,I198185,I198694);
not I_11519 (I198739,I198519);
nand I_11520 (I198756,I198739,I198615);
nor I_11521 (I198094,I198219,I198756);
not I_11522 (I198814,I2905);
nand I_11523 (I198831,I258948,I258945);
and I_11524 (I198848,I198831,I258951);
DFFARX1 I_11525 (I198848,I2898,I198814,I198874,);
not I_11526 (I198882,I198874);
nor I_11527 (I198899,I258957,I258945);
not I_11528 (I198916,I198899);
not I_11529 (I198933,I258948);
nand I_11530 (I198950,I258945,I258954);
nand I_11531 (I198967,I198950,I258948);
not I_11532 (I198984,I198967);
nor I_11533 (I198794,I198984,I198874);
nand I_11534 (I199015,I198950,I198933);
and I_11535 (I199032,I199015,I258975);
nand I_11536 (I199049,I199032,I258963);
and I_11537 (I199066,I199049,I198967);
nor I_11538 (I199083,I199049,I198967);
or I_11539 (I199100,I258954,I258966);
nor I_11540 (I199117,I199100,I258960);
not I_11541 (I199134,I199117);
nor I_11542 (I199151,I198916,I199134);
and I_11543 (I198785,I199151,I198882);
nor I_11544 (I199182,I198967,I199134);
nand I_11545 (I199199,I198984,I199117);
nand I_11546 (I199216,I258969,I258972);
nor I_11547 (I198782,I199216,I199117);
nor I_11548 (I199247,I199216,I199134);
not I_11549 (I199264,I199247);
nor I_11550 (I198806,I199066,I199264);
or I_11551 (I199295,I199216,I258951);
nand I_11552 (I199312,I199295,I199199);
not I_11553 (I199329,I199312);
nor I_11554 (I198788,I199329,I199182);
nor I_11555 (I199360,I199295,I199083);
DFFARX1 I_11556 (I199360,I2898,I198814,I198797,);
and I_11557 (I199391,I199049,I199295);
nor I_11558 (I198803,I199391,I198899);
nor I_11559 (I198800,I198882,I199391);
not I_11560 (I199436,I199216);
nand I_11561 (I199453,I199436,I199312);
nor I_11562 (I198791,I198916,I199453);
not I_11563 (I199511,I2905);
nand I_11564 (I199528,I431045,I431036);
and I_11565 (I199545,I199528,I431039);
DFFARX1 I_11566 (I199545,I2898,I199511,I199571,);
not I_11567 (I199579,I199571);
nor I_11568 (I199596,I431054,I431036);
not I_11569 (I199613,I199596);
not I_11570 (I199630,I431066);
nand I_11571 (I199647,I431063,I431057);
nand I_11572 (I199664,I199647,I431066);
not I_11573 (I199681,I199664);
nor I_11574 (I199491,I199681,I199571);
nand I_11575 (I199712,I199647,I199630);
and I_11576 (I199729,I199712,I431060);
nand I_11577 (I199746,I199729,I431042);
and I_11578 (I199763,I199746,I199664);
nor I_11579 (I199780,I199746,I199664);
or I_11580 (I199797,I431039,I431051);
nor I_11581 (I199814,I199797,I431048);
not I_11582 (I199831,I199814);
nor I_11583 (I199848,I199613,I199831);
and I_11584 (I199482,I199848,I199579);
nor I_11585 (I199879,I199664,I199831);
nand I_11586 (I199896,I199681,I199814);
nand I_11587 (I199913,I431042,I431069);
nor I_11588 (I199479,I199913,I199814);
nor I_11589 (I199944,I199913,I199831);
not I_11590 (I199961,I199944);
nor I_11591 (I199503,I199763,I199961);
or I_11592 (I199992,I199913,I431036);
nand I_11593 (I200009,I199992,I199896);
not I_11594 (I200026,I200009);
nor I_11595 (I199485,I200026,I199879);
nor I_11596 (I200057,I199992,I199780);
DFFARX1 I_11597 (I200057,I2898,I199511,I199494,);
and I_11598 (I200088,I199746,I199992);
nor I_11599 (I199500,I200088,I199596);
nor I_11600 (I199497,I199579,I200088);
not I_11601 (I200133,I199913);
nand I_11602 (I200150,I200133,I200009);
nor I_11603 (I199488,I199613,I200150);
not I_11604 (I200208,I2905);
nand I_11605 (I200225,I326996,I327008);
and I_11606 (I200242,I200225,I326999);
DFFARX1 I_11607 (I200242,I2898,I200208,I200268,);
not I_11608 (I200276,I200268);
nor I_11609 (I200293,I327011,I327008);
not I_11610 (I200310,I200293);
not I_11611 (I200327,I327017);
nand I_11612 (I200344,I327002,I327005);
nand I_11613 (I200361,I200344,I327017);
not I_11614 (I200378,I200361);
nor I_11615 (I200188,I200378,I200268);
nand I_11616 (I200409,I200344,I200327);
and I_11617 (I200426,I200409,I327014);
nand I_11618 (I200443,I200426,I327002);
and I_11619 (I200460,I200443,I200361);
nor I_11620 (I200477,I200443,I200361);
or I_11621 (I200494,I327020,I327005);
nor I_11622 (I200511,I200494,I327011);
not I_11623 (I200528,I200511);
nor I_11624 (I200545,I200310,I200528);
and I_11625 (I200179,I200545,I200276);
nor I_11626 (I200576,I200361,I200528);
nand I_11627 (I200593,I200378,I200511);
nand I_11628 (I200610,I326996,I327008);
nor I_11629 (I200176,I200610,I200511);
nor I_11630 (I200641,I200610,I200528);
not I_11631 (I200658,I200641);
nor I_11632 (I200200,I200460,I200658);
or I_11633 (I200689,I200610,I326999);
nand I_11634 (I200706,I200689,I200593);
not I_11635 (I200723,I200706);
nor I_11636 (I200182,I200723,I200576);
nor I_11637 (I200754,I200689,I200477);
DFFARX1 I_11638 (I200754,I2898,I200208,I200191,);
and I_11639 (I200785,I200443,I200689);
nor I_11640 (I200197,I200785,I200293);
nor I_11641 (I200194,I200276,I200785);
not I_11642 (I200830,I200610);
nand I_11643 (I200847,I200830,I200706);
nor I_11644 (I200185,I200310,I200847);
not I_11645 (I200905,I2905);
nand I_11646 (I200922,I54291,I54312);
and I_11647 (I200939,I200922,I54309);
DFFARX1 I_11648 (I200939,I2898,I200905,I200965,);
not I_11649 (I200973,I200965);
nor I_11650 (I200990,I54288,I54312);
not I_11651 (I201007,I200990);
not I_11652 (I201024,I54294);
nand I_11653 (I201041,I54315,I54306);
nand I_11654 (I201058,I201041,I54294);
not I_11655 (I201075,I201058);
nor I_11656 (I200885,I201075,I200965);
nand I_11657 (I201106,I201041,I201024);
and I_11658 (I201123,I201106,I54318);
nand I_11659 (I201140,I201123,I54285);
and I_11660 (I201157,I201140,I201058);
nor I_11661 (I201174,I201140,I201058);
or I_11662 (I201191,I54282,I54297);
nor I_11663 (I201208,I201191,I54282);
not I_11664 (I201225,I201208);
nor I_11665 (I201242,I201007,I201225);
and I_11666 (I200876,I201242,I200973);
nor I_11667 (I201273,I201058,I201225);
nand I_11668 (I201290,I201075,I201208);
nand I_11669 (I201307,I54303,I54300);
nor I_11670 (I200873,I201307,I201208);
nor I_11671 (I201338,I201307,I201225);
not I_11672 (I201355,I201338);
nor I_11673 (I200897,I201157,I201355);
or I_11674 (I201386,I201307,I54285);
nand I_11675 (I201403,I201386,I201290);
not I_11676 (I201420,I201403);
nor I_11677 (I200879,I201420,I201273);
nor I_11678 (I201451,I201386,I201174);
DFFARX1 I_11679 (I201451,I2898,I200905,I200888,);
and I_11680 (I201482,I201140,I201386);
nor I_11681 (I200894,I201482,I200990);
nor I_11682 (I200891,I200973,I201482);
not I_11683 (I201527,I201307);
nand I_11684 (I201544,I201527,I201403);
nor I_11685 (I200882,I201007,I201544);
not I_11686 (I201602,I2905);
nand I_11687 (I201619,I256653,I256650);
and I_11688 (I201636,I201619,I256656);
DFFARX1 I_11689 (I201636,I2898,I201602,I201662,);
not I_11690 (I201670,I201662);
nor I_11691 (I201687,I256662,I256650);
not I_11692 (I201704,I201687);
not I_11693 (I201721,I256653);
nand I_11694 (I201738,I256650,I256659);
nand I_11695 (I201755,I201738,I256653);
not I_11696 (I201772,I201755);
nor I_11697 (I201582,I201772,I201662);
nand I_11698 (I201803,I201738,I201721);
and I_11699 (I201820,I201803,I256680);
nand I_11700 (I201837,I201820,I256668);
and I_11701 (I201854,I201837,I201755);
nor I_11702 (I201871,I201837,I201755);
or I_11703 (I201888,I256659,I256671);
nor I_11704 (I201905,I201888,I256665);
not I_11705 (I201922,I201905);
nor I_11706 (I201939,I201704,I201922);
and I_11707 (I201573,I201939,I201670);
nor I_11708 (I201970,I201755,I201922);
nand I_11709 (I201987,I201772,I201905);
nand I_11710 (I202004,I256674,I256677);
nor I_11711 (I201570,I202004,I201905);
nor I_11712 (I202035,I202004,I201922);
not I_11713 (I202052,I202035);
nor I_11714 (I201594,I201854,I202052);
or I_11715 (I202083,I202004,I256656);
nand I_11716 (I202100,I202083,I201987);
not I_11717 (I202117,I202100);
nor I_11718 (I201576,I202117,I201970);
nor I_11719 (I202148,I202083,I201871);
DFFARX1 I_11720 (I202148,I2898,I201602,I201585,);
and I_11721 (I202179,I201837,I202083);
nor I_11722 (I201591,I202179,I201687);
nor I_11723 (I201588,I201670,I202179);
not I_11724 (I202224,I202004);
nand I_11725 (I202241,I202224,I202100);
nor I_11726 (I201579,I201704,I202241);
not I_11727 (I202299,I2905);
nand I_11728 (I202316,I322831,I322843);
and I_11729 (I202333,I202316,I322834);
DFFARX1 I_11730 (I202333,I2898,I202299,I202359,);
not I_11731 (I202367,I202359);
nor I_11732 (I202384,I322846,I322843);
not I_11733 (I202401,I202384);
not I_11734 (I202418,I322852);
nand I_11735 (I202435,I322837,I322840);
nand I_11736 (I202452,I202435,I322852);
not I_11737 (I202469,I202452);
nor I_11738 (I202279,I202469,I202359);
nand I_11739 (I202500,I202435,I202418);
and I_11740 (I202517,I202500,I322849);
nand I_11741 (I202534,I202517,I322837);
and I_11742 (I202551,I202534,I202452);
nor I_11743 (I202568,I202534,I202452);
or I_11744 (I202585,I322855,I322840);
nor I_11745 (I202602,I202585,I322846);
not I_11746 (I202619,I202602);
nor I_11747 (I202636,I202401,I202619);
and I_11748 (I202270,I202636,I202367);
nor I_11749 (I202667,I202452,I202619);
nand I_11750 (I202684,I202469,I202602);
nand I_11751 (I202701,I322831,I322843);
nor I_11752 (I202267,I202701,I202602);
nor I_11753 (I202732,I202701,I202619);
not I_11754 (I202749,I202732);
nor I_11755 (I202291,I202551,I202749);
or I_11756 (I202780,I202701,I322834);
nand I_11757 (I202797,I202780,I202684);
not I_11758 (I202814,I202797);
nor I_11759 (I202273,I202814,I202667);
nor I_11760 (I202845,I202780,I202568);
DFFARX1 I_11761 (I202845,I2898,I202299,I202282,);
and I_11762 (I202876,I202534,I202780);
nor I_11763 (I202288,I202876,I202384);
nor I_11764 (I202285,I202367,I202876);
not I_11765 (I202921,I202701);
nand I_11766 (I202938,I202921,I202797);
nor I_11767 (I202276,I202401,I202938);
not I_11768 (I202999,I2905);
nand I_11769 (I203016,I5989,I5968);
and I_11770 (I203033,I203016,I5983);
DFFARX1 I_11771 (I203033,I2898,I202999,I203059,);
not I_11772 (I203067,I203059);
nor I_11773 (I203084,I5971,I5968);
or I_11774 (I203101,I203059,I203084);
nor I_11775 (I203118,I5986,I5992);
not I_11776 (I203135,I203118);
nor I_11777 (I203152,I203135,I203101);
nor I_11778 (I203169,I5968,I5986);
nor I_11779 (I203186,I203067,I203169);
or I_11780 (I203203,I203169,I5992);
not I_11781 (I203220,I5971);
nor I_11782 (I203237,I203220,I5995);
nor I_11783 (I203254,I203237,I203203);
nor I_11784 (I203271,I203135,I5995);
and I_11785 (I203288,I203271,I5971);
nor I_11786 (I202991,I203288,I203084);
nor I_11787 (I203319,I5995,I5977);
nand I_11788 (I203336,I203319,I203118);
not I_11789 (I203353,I203336);
nor I_11790 (I203370,I203152,I203353);
DFFARX1 I_11791 (I203319,I2898,I202999,I202973,);
nor I_11792 (I203401,I5974,I5968);
nand I_11793 (I203418,I203084,I203401);
not I_11794 (I202967,I203418);
nor I_11795 (I203449,I5974,I5977);
DFFARX1 I_11796 (I203449,I2898,I202999,I203475,);
nor I_11797 (I203483,I203475,I203186);
nor I_11798 (I202970,I203483,I203418);
nor I_11799 (I202964,I203475,I203370);
and I_11800 (I202982,I203169,I5974);
nand I_11801 (I203542,I5980,I5998);
nor I_11802 (I203559,I203542,I5974);
not I_11803 (I203576,I203559);
nor I_11804 (I203593,I203576,I203254);
DFFARX1 I_11805 (I203593,I2898,I202999,I202985,);
nor I_11806 (I203624,I203559,I203118);
nor I_11807 (I202988,I203542,I203288);
nor I_11808 (I203655,I203059,I203542);
nand I_11809 (I202979,I203655,I5974);
not I_11810 (I203686,I203542);
nand I_11811 (I202976,I203624,I203686);
not I_11812 (I203747,I2905);
nand I_11813 (I203764,I281151,I281136);
and I_11814 (I203781,I203764,I281130);
DFFARX1 I_11815 (I203781,I2898,I203747,I203807,);
not I_11816 (I203815,I203807);
nor I_11817 (I203832,I281133,I281136);
or I_11818 (I203849,I203807,I203832);
nor I_11819 (I203866,I281160,I281154);
not I_11820 (I203883,I203866);
nor I_11821 (I203900,I203883,I203849);
nor I_11822 (I203917,I281157,I281160);
nor I_11823 (I203934,I203815,I203917);
or I_11824 (I203951,I203917,I281154);
not I_11825 (I203968,I281145);
nor I_11826 (I203985,I203968,I281136);
nor I_11827 (I204002,I203985,I203951);
nor I_11828 (I204019,I203883,I281136);
and I_11829 (I204036,I204019,I281145);
nor I_11830 (I203739,I204036,I203832);
nor I_11831 (I204067,I281136,I281139);
nand I_11832 (I204084,I204067,I203866);
not I_11833 (I204101,I204084);
nor I_11834 (I204118,I203900,I204101);
DFFARX1 I_11835 (I204067,I2898,I203747,I203721,);
nor I_11836 (I204149,I281142,I281157);
nand I_11837 (I204166,I203832,I204149);
not I_11838 (I203715,I204166);
nor I_11839 (I204197,I281142,I281139);
DFFARX1 I_11840 (I204197,I2898,I203747,I204223,);
nor I_11841 (I204231,I204223,I203934);
nor I_11842 (I203718,I204231,I204166);
nor I_11843 (I203712,I204223,I204118);
and I_11844 (I203730,I203917,I281142);
nand I_11845 (I204290,I281133,I281130);
nor I_11846 (I204307,I204290,I281148);
not I_11847 (I204324,I204307);
nor I_11848 (I204341,I204324,I204002);
DFFARX1 I_11849 (I204341,I2898,I203747,I203733,);
nor I_11850 (I204372,I204307,I203866);
nor I_11851 (I203736,I204290,I204036);
nor I_11852 (I204403,I203807,I204290);
nand I_11853 (I203727,I204403,I281148);
not I_11854 (I204434,I204290);
nand I_11855 (I203724,I204372,I204434);
not I_11856 (I204495,I2905);
nand I_11857 (I204512,I136796,I136799);
and I_11858 (I204529,I204512,I136781);
DFFARX1 I_11859 (I204529,I2898,I204495,I204555,);
not I_11860 (I204563,I204555);
nor I_11861 (I204580,I136766,I136799);
or I_11862 (I204597,I204555,I204580);
nor I_11863 (I204614,I136778,I136775);
not I_11864 (I204631,I204614);
nor I_11865 (I204648,I204631,I204597);
nor I_11866 (I204665,I136784,I136778);
nor I_11867 (I204682,I204563,I204665);
or I_11868 (I204699,I204665,I136775);
not I_11869 (I204716,I136790);
nor I_11870 (I204733,I204716,I136769);
nor I_11871 (I204750,I204733,I204699);
nor I_11872 (I204767,I204631,I136769);
and I_11873 (I204784,I204767,I136790);
nor I_11874 (I204487,I204784,I204580);
nor I_11875 (I204815,I136769,I136769);
nand I_11876 (I204832,I204815,I204614);
not I_11877 (I204849,I204832);
nor I_11878 (I204866,I204648,I204849);
DFFARX1 I_11879 (I204815,I2898,I204495,I204469,);
nor I_11880 (I204897,I136766,I136784);
nand I_11881 (I204914,I204580,I204897);
not I_11882 (I204463,I204914);
nor I_11883 (I204945,I136766,I136772);
DFFARX1 I_11884 (I204945,I2898,I204495,I204971,);
nor I_11885 (I204979,I204971,I204682);
nor I_11886 (I204466,I204979,I204914);
nor I_11887 (I204460,I204971,I204866);
and I_11888 (I204478,I204665,I136766);
nand I_11889 (I205038,I136793,I136787);
nor I_11890 (I205055,I205038,I136772);
not I_11891 (I205072,I205055);
nor I_11892 (I205089,I205072,I204750);
DFFARX1 I_11893 (I205089,I2898,I204495,I204481,);
nor I_11894 (I205120,I205055,I204614);
nor I_11895 (I204484,I205038,I204784);
nor I_11896 (I205151,I204555,I205038);
nand I_11897 (I204475,I205151,I136772);
not I_11898 (I205182,I205038);
nand I_11899 (I204472,I205120,I205182);
not I_11900 (I205243,I2905);
nand I_11901 (I205260,I16093,I16075);
and I_11902 (I205277,I205260,I16066);
DFFARX1 I_11903 (I205277,I2898,I205243,I205303,);
not I_11904 (I205311,I205303);
nor I_11905 (I205328,I16069,I16075);
or I_11906 (I205345,I205303,I205328);
nor I_11907 (I205362,I16084,I16075);
not I_11908 (I205379,I205362);
nor I_11909 (I205396,I205379,I205345);
nor I_11910 (I205413,I16081,I16084);
nor I_11911 (I205430,I205311,I205413);
or I_11912 (I205447,I205413,I16075);
not I_11913 (I205464,I16078);
nor I_11914 (I205481,I205464,I16072);
nor I_11915 (I205498,I205481,I205447);
nor I_11916 (I205515,I205379,I16072);
and I_11917 (I205532,I205515,I16078);
nor I_11918 (I205235,I205532,I205328);
nor I_11919 (I205563,I16072,I16078);
nand I_11920 (I205580,I205563,I205362);
not I_11921 (I205597,I205580);
nor I_11922 (I205614,I205396,I205597);
DFFARX1 I_11923 (I205563,I2898,I205243,I205217,);
nor I_11924 (I205645,I16090,I16081);
nand I_11925 (I205662,I205328,I205645);
not I_11926 (I205211,I205662);
nor I_11927 (I205693,I16090,I16069);
DFFARX1 I_11928 (I205693,I2898,I205243,I205719,);
nor I_11929 (I205727,I205719,I205430);
nor I_11930 (I205214,I205727,I205662);
nor I_11931 (I205208,I205719,I205614);
and I_11932 (I205226,I205413,I16090);
nand I_11933 (I205786,I16087,I16066);
nor I_11934 (I205803,I205786,I16072);
not I_11935 (I205820,I205803);
nor I_11936 (I205837,I205820,I205498);
DFFARX1 I_11937 (I205837,I2898,I205243,I205229,);
nor I_11938 (I205868,I205803,I205362);
nor I_11939 (I205232,I205786,I205532);
nor I_11940 (I205899,I205303,I205786);
nand I_11941 (I205223,I205899,I16072);
not I_11942 (I205930,I205786);
nand I_11943 (I205220,I205868,I205930);
not I_11944 (I205991,I2905);
nand I_11945 (I206008,I381635,I381617);
and I_11946 (I206025,I206008,I381641);
DFFARX1 I_11947 (I206025,I2898,I205991,I206051,);
not I_11948 (I206059,I206051);
nor I_11949 (I206076,I381644,I381617);
or I_11950 (I206093,I206051,I206076);
nor I_11951 (I206110,I381650,I381632);
not I_11952 (I206127,I206110);
nor I_11953 (I206144,I206127,I206093);
nor I_11954 (I206161,I381626,I381650);
nor I_11955 (I206178,I206059,I206161);
or I_11956 (I206195,I206161,I381632);
not I_11957 (I206212,I381623);
nor I_11958 (I206229,I206212,I381638);
nor I_11959 (I206246,I206229,I206195);
nor I_11960 (I206263,I206127,I381638);
and I_11961 (I206280,I206263,I381623);
nor I_11962 (I205983,I206280,I206076);
nor I_11963 (I206311,I381638,I381620);
nand I_11964 (I206328,I206311,I206110);
not I_11965 (I206345,I206328);
nor I_11966 (I206362,I206144,I206345);
DFFARX1 I_11967 (I206311,I2898,I205991,I205965,);
nor I_11968 (I206393,I381623,I381626);
nand I_11969 (I206410,I206076,I206393);
not I_11970 (I205959,I206410);
nor I_11971 (I206441,I381623,I381647);
DFFARX1 I_11972 (I206441,I2898,I205991,I206467,);
nor I_11973 (I206475,I206467,I206178);
nor I_11974 (I205962,I206475,I206410);
nor I_11975 (I205956,I206467,I206362);
and I_11976 (I205974,I206161,I381623);
nand I_11977 (I206534,I381629,I381617);
nor I_11978 (I206551,I206534,I381620);
not I_11979 (I206568,I206551);
nor I_11980 (I206585,I206568,I206246);
DFFARX1 I_11981 (I206585,I2898,I205991,I205977,);
nor I_11982 (I206616,I206551,I206110);
nor I_11983 (I205980,I206534,I206280);
nor I_11984 (I206647,I206051,I206534);
nand I_11985 (I205971,I206647,I381620);
not I_11986 (I206678,I206534);
nand I_11987 (I205968,I206616,I206678);
not I_11988 (I206739,I2905);
nand I_11989 (I206756,I1611,I2107);
and I_11990 (I206773,I206756,I2363);
DFFARX1 I_11991 (I206773,I2898,I206739,I206799,);
not I_11992 (I206807,I206799);
nor I_11993 (I206824,I2043,I2107);
or I_11994 (I206841,I206799,I206824);
nor I_11995 (I206858,I1643,I1835);
not I_11996 (I206875,I206858);
nor I_11997 (I206892,I206875,I206841);
nor I_11998 (I206909,I2723,I1643);
nor I_11999 (I206926,I206807,I206909);
or I_12000 (I206943,I206909,I1835);
not I_12001 (I206960,I2667);
nor I_12002 (I206977,I206960,I2011);
nor I_12003 (I206994,I206977,I206943);
nor I_12004 (I207011,I206875,I2011);
and I_12005 (I207028,I207011,I2667);
nor I_12006 (I206731,I207028,I206824);
nor I_12007 (I207059,I2011,I2819);
nand I_12008 (I207076,I207059,I206858);
not I_12009 (I207093,I207076);
nor I_12010 (I207110,I206892,I207093);
DFFARX1 I_12011 (I207059,I2898,I206739,I206713,);
nor I_12012 (I207141,I1691,I2723);
nand I_12013 (I207158,I206824,I207141);
not I_12014 (I206707,I207158);
nor I_12015 (I207189,I1691,I2083);
DFFARX1 I_12016 (I207189,I2898,I206739,I207215,);
nor I_12017 (I207223,I207215,I206926);
nor I_12018 (I206710,I207223,I207158);
nor I_12019 (I206704,I207215,I207110);
and I_12020 (I206722,I206909,I1691);
nand I_12021 (I207282,I2675,I2243);
nor I_12022 (I207299,I207282,I2075);
not I_12023 (I207316,I207299);
nor I_12024 (I207333,I207316,I206994);
DFFARX1 I_12025 (I207333,I2898,I206739,I206725,);
nor I_12026 (I207364,I207299,I206858);
nor I_12027 (I206728,I207282,I207028);
nor I_12028 (I207395,I206799,I207282);
nand I_12029 (I206719,I207395,I2075);
not I_12030 (I207426,I207282);
nand I_12031 (I206716,I207364,I207426);
not I_12032 (I207487,I2905);
nand I_12033 (I207504,I104717,I104720);
and I_12034 (I207521,I207504,I104702);
DFFARX1 I_12035 (I207521,I2898,I207487,I207547,);
not I_12036 (I207555,I207547);
nor I_12037 (I207572,I104687,I104720);
or I_12038 (I207589,I207547,I207572);
nor I_12039 (I207606,I104699,I104696);
not I_12040 (I207623,I207606);
nor I_12041 (I207640,I207623,I207589);
nor I_12042 (I207657,I104705,I104699);
nor I_12043 (I207674,I207555,I207657);
or I_12044 (I207691,I207657,I104696);
not I_12045 (I207708,I104711);
nor I_12046 (I207725,I207708,I104690);
nor I_12047 (I207742,I207725,I207691);
nor I_12048 (I207759,I207623,I104690);
and I_12049 (I207776,I207759,I104711);
nor I_12050 (I207479,I207776,I207572);
nor I_12051 (I207807,I104690,I104690);
nand I_12052 (I207824,I207807,I207606);
not I_12053 (I207841,I207824);
nor I_12054 (I207858,I207640,I207841);
DFFARX1 I_12055 (I207807,I2898,I207487,I207461,);
nor I_12056 (I207889,I104687,I104705);
nand I_12057 (I207906,I207572,I207889);
not I_12058 (I207455,I207906);
nor I_12059 (I207937,I104687,I104693);
DFFARX1 I_12060 (I207937,I2898,I207487,I207963,);
nor I_12061 (I207971,I207963,I207674);
nor I_12062 (I207458,I207971,I207906);
nor I_12063 (I207452,I207963,I207858);
and I_12064 (I207470,I207657,I104687);
nand I_12065 (I208030,I104714,I104708);
nor I_12066 (I208047,I208030,I104693);
not I_12067 (I208064,I208047);
nor I_12068 (I208081,I208064,I207742);
DFFARX1 I_12069 (I208081,I2898,I207487,I207473,);
nor I_12070 (I208112,I208047,I207606);
nor I_12071 (I207476,I208030,I207776);
nor I_12072 (I208143,I207547,I208030);
nand I_12073 (I207467,I208143,I104693);
not I_12074 (I208174,I208030);
nand I_12075 (I207464,I208112,I208174);
not I_12076 (I208235,I2905);
nand I_12077 (I208252,I390033,I390015);
and I_12078 (I208269,I208252,I390039);
DFFARX1 I_12079 (I208269,I2898,I208235,I208295,);
not I_12080 (I208303,I208295);
nor I_12081 (I208320,I390042,I390015);
or I_12082 (I208337,I208295,I208320);
nor I_12083 (I208354,I390048,I390030);
not I_12084 (I208371,I208354);
nor I_12085 (I208388,I208371,I208337);
nor I_12086 (I208405,I390024,I390048);
nor I_12087 (I208422,I208303,I208405);
or I_12088 (I208439,I208405,I390030);
not I_12089 (I208456,I390021);
nor I_12090 (I208473,I208456,I390036);
nor I_12091 (I208490,I208473,I208439);
nor I_12092 (I208507,I208371,I390036);
and I_12093 (I208524,I208507,I390021);
nor I_12094 (I208227,I208524,I208320);
nor I_12095 (I208555,I390036,I390018);
nand I_12096 (I208572,I208555,I208354);
not I_12097 (I208589,I208572);
nor I_12098 (I208606,I208388,I208589);
DFFARX1 I_12099 (I208555,I2898,I208235,I208209,);
nor I_12100 (I208637,I390021,I390024);
nand I_12101 (I208654,I208320,I208637);
not I_12102 (I208203,I208654);
nor I_12103 (I208685,I390021,I390045);
DFFARX1 I_12104 (I208685,I2898,I208235,I208711,);
nor I_12105 (I208719,I208711,I208422);
nor I_12106 (I208206,I208719,I208654);
nor I_12107 (I208200,I208711,I208606);
and I_12108 (I208218,I208405,I390021);
nand I_12109 (I208778,I390027,I390015);
nor I_12110 (I208795,I208778,I390018);
not I_12111 (I208812,I208795);
nor I_12112 (I208829,I208812,I208490);
DFFARX1 I_12113 (I208829,I2898,I208235,I208221,);
nor I_12114 (I208860,I208795,I208354);
nor I_12115 (I208224,I208778,I208524);
nor I_12116 (I208891,I208295,I208778);
nand I_12117 (I208215,I208891,I390018);
not I_12118 (I208922,I208778);
nand I_12119 (I208212,I208860,I208922);
not I_12120 (I208983,I2905);
nand I_12121 (I209000,I31801,I31783);
and I_12122 (I209017,I209000,I31774);
DFFARX1 I_12123 (I209017,I2898,I208983,I209043,);
not I_12124 (I209051,I209043);
nor I_12125 (I209068,I31777,I31783);
or I_12126 (I209085,I209043,I209068);
nor I_12127 (I209102,I31792,I31783);
not I_12128 (I209119,I209102);
nor I_12129 (I209136,I209119,I209085);
nor I_12130 (I209153,I31789,I31792);
nor I_12131 (I209170,I209051,I209153);
or I_12132 (I209187,I209153,I31783);
not I_12133 (I209204,I31786);
nor I_12134 (I209221,I209204,I31780);
nor I_12135 (I209238,I209221,I209187);
nor I_12136 (I209255,I209119,I31780);
and I_12137 (I209272,I209255,I31786);
nor I_12138 (I208975,I209272,I209068);
nor I_12139 (I209303,I31780,I31786);
nand I_12140 (I209320,I209303,I209102);
not I_12141 (I209337,I209320);
nor I_12142 (I209354,I209136,I209337);
DFFARX1 I_12143 (I209303,I2898,I208983,I208957,);
nor I_12144 (I209385,I31798,I31789);
nand I_12145 (I209402,I209068,I209385);
not I_12146 (I208951,I209402);
nor I_12147 (I209433,I31798,I31777);
DFFARX1 I_12148 (I209433,I2898,I208983,I209459,);
nor I_12149 (I209467,I209459,I209170);
nor I_12150 (I208954,I209467,I209402);
nor I_12151 (I208948,I209459,I209354);
and I_12152 (I208966,I209153,I31798);
nand I_12153 (I209526,I31795,I31774);
nor I_12154 (I209543,I209526,I31780);
not I_12155 (I209560,I209543);
nor I_12156 (I209577,I209560,I209238);
DFFARX1 I_12157 (I209577,I2898,I208983,I208969,);
nor I_12158 (I209608,I209543,I209102);
nor I_12159 (I208972,I209526,I209272);
nor I_12160 (I209639,I209043,I209526);
nand I_12161 (I208963,I209639,I31780);
not I_12162 (I209670,I209526);
nand I_12163 (I208960,I209608,I209670);
not I_12164 (I209731,I2905);
nand I_12165 (I209748,I301774,I301771);
and I_12166 (I209765,I209748,I301768);
DFFARX1 I_12167 (I209765,I2898,I209731,I209791,);
not I_12168 (I209799,I209791);
nor I_12169 (I209816,I301777,I301771);
or I_12170 (I209833,I209791,I209816);
nor I_12171 (I209850,I301795,I301768);
not I_12172 (I209867,I209850);
nor I_12173 (I209884,I209867,I209833);
nor I_12174 (I209901,I301798,I301795);
nor I_12175 (I209918,I209799,I209901);
or I_12176 (I209935,I209901,I301768);
not I_12177 (I209952,I301783);
nor I_12178 (I209969,I209952,I301789);
nor I_12179 (I209986,I209969,I209935);
nor I_12180 (I210003,I209867,I301789);
and I_12181 (I210020,I210003,I301783);
nor I_12182 (I209723,I210020,I209816);
nor I_12183 (I210051,I301789,I301777);
nand I_12184 (I210068,I210051,I209850);
not I_12185 (I210085,I210068);
nor I_12186 (I210102,I209884,I210085);
DFFARX1 I_12187 (I210051,I2898,I209731,I209705,);
nor I_12188 (I210133,I301774,I301798);
nand I_12189 (I210150,I209816,I210133);
not I_12190 (I209699,I210150);
nor I_12191 (I210181,I301774,I301771);
DFFARX1 I_12192 (I210181,I2898,I209731,I210207,);
nor I_12193 (I210215,I210207,I209918);
nor I_12194 (I209702,I210215,I210150);
nor I_12195 (I209696,I210207,I210102);
and I_12196 (I209714,I209901,I301774);
nand I_12197 (I210274,I301780,I301786);
nor I_12198 (I210291,I210274,I301792);
not I_12199 (I210308,I210291);
nor I_12200 (I210325,I210308,I209986);
DFFARX1 I_12201 (I210325,I2898,I209731,I209717,);
nor I_12202 (I210356,I210291,I209850);
nor I_12203 (I209720,I210274,I210020);
nor I_12204 (I210387,I209791,I210274);
nand I_12205 (I209711,I210387,I301792);
not I_12206 (I210418,I210274);
nand I_12207 (I209708,I210356,I210418);
not I_12208 (I210479,I2905);
nand I_12209 (I210496,I172194,I172206);
and I_12210 (I210513,I210496,I172200);
DFFARX1 I_12211 (I210513,I2898,I210479,I210539,);
not I_12212 (I210547,I210539);
nor I_12213 (I210564,I172200,I172206);
or I_12214 (I210581,I210539,I210564);
nor I_12215 (I210598,I172221,I172209);
not I_12216 (I210615,I210598);
nor I_12217 (I210632,I210615,I210581);
nor I_12218 (I210649,I172218,I172221);
nor I_12219 (I210666,I210547,I210649);
or I_12220 (I210683,I210649,I172209);
not I_12221 (I210700,I172212);
nor I_12222 (I210717,I210700,I172194);
nor I_12223 (I210734,I210717,I210683);
nor I_12224 (I210751,I210615,I172194);
and I_12225 (I210768,I210751,I172212);
nor I_12226 (I210471,I210768,I210564);
nor I_12227 (I210799,I172194,I172197);
nand I_12228 (I210816,I210799,I210598);
not I_12229 (I210833,I210816);
nor I_12230 (I210850,I210632,I210833);
DFFARX1 I_12231 (I210799,I2898,I210479,I210453,);
nor I_12232 (I210881,I172224,I172218);
nand I_12233 (I210898,I210564,I210881);
not I_12234 (I210447,I210898);
nor I_12235 (I210929,I172224,I172203);
DFFARX1 I_12236 (I210929,I2898,I210479,I210955,);
nor I_12237 (I210963,I210955,I210666);
nor I_12238 (I210450,I210963,I210898);
nor I_12239 (I210444,I210955,I210850);
and I_12240 (I210462,I210649,I172224);
nand I_12241 (I211022,I172215,I172197);
nor I_12242 (I211039,I211022,I172227);
not I_12243 (I211056,I211039);
nor I_12244 (I211073,I211056,I210734);
DFFARX1 I_12245 (I211073,I2898,I210479,I210465,);
nor I_12246 (I211104,I211039,I210598);
nor I_12247 (I210468,I211022,I210768);
nor I_12248 (I211135,I210539,I211022);
nand I_12249 (I210459,I211135,I172227);
not I_12250 (I211166,I211022);
nand I_12251 (I210456,I211104,I211166);
not I_12252 (I211227,I2905);
nand I_12253 (I211244,I266616,I266601);
and I_12254 (I211261,I211244,I266595);
DFFARX1 I_12255 (I211261,I2898,I211227,I211287,);
not I_12256 (I211295,I211287);
nor I_12257 (I211312,I266598,I266601);
or I_12258 (I211329,I211287,I211312);
nor I_12259 (I211346,I266625,I266619);
not I_12260 (I211363,I211346);
nor I_12261 (I211380,I211363,I211329);
nor I_12262 (I211397,I266622,I266625);
nor I_12263 (I211414,I211295,I211397);
or I_12264 (I211431,I211397,I266619);
not I_12265 (I211448,I266610);
nor I_12266 (I211465,I211448,I266601);
nor I_12267 (I211482,I211465,I211431);
nor I_12268 (I211499,I211363,I266601);
and I_12269 (I211516,I211499,I266610);
nor I_12270 (I211219,I211516,I211312);
nor I_12271 (I211547,I266601,I266604);
nand I_12272 (I211564,I211547,I211346);
not I_12273 (I211581,I211564);
nor I_12274 (I211598,I211380,I211581);
DFFARX1 I_12275 (I211547,I2898,I211227,I211201,);
nor I_12276 (I211629,I266607,I266622);
nand I_12277 (I211646,I211312,I211629);
not I_12278 (I211195,I211646);
nor I_12279 (I211677,I266607,I266604);
DFFARX1 I_12280 (I211677,I2898,I211227,I211703,);
nor I_12281 (I211711,I211703,I211414);
nor I_12282 (I211198,I211711,I211646);
nor I_12283 (I211192,I211703,I211598);
and I_12284 (I211210,I211397,I266607);
nand I_12285 (I211770,I266598,I266595);
nor I_12286 (I211787,I211770,I266613);
not I_12287 (I211804,I211787);
nor I_12288 (I211821,I211804,I211482);
DFFARX1 I_12289 (I211821,I2898,I211227,I211213,);
nor I_12290 (I211852,I211787,I211346);
nor I_12291 (I211216,I211770,I211516);
nor I_12292 (I211883,I211287,I211770);
nand I_12293 (I211207,I211883,I266613);
not I_12294 (I211914,I211770);
nand I_12295 (I211204,I211852,I211914);
not I_12296 (I211975,I2905);
nand I_12297 (I211992,I130506,I130509);
and I_12298 (I212009,I211992,I130491);
DFFARX1 I_12299 (I212009,I2898,I211975,I212035,);
not I_12300 (I212043,I212035);
nor I_12301 (I212060,I130476,I130509);
or I_12302 (I212077,I212035,I212060);
nor I_12303 (I212094,I130488,I130485);
not I_12304 (I212111,I212094);
nor I_12305 (I212128,I212111,I212077);
nor I_12306 (I212145,I130494,I130488);
nor I_12307 (I212162,I212043,I212145);
or I_12308 (I212179,I212145,I130485);
not I_12309 (I212196,I130500);
nor I_12310 (I212213,I212196,I130479);
nor I_12311 (I212230,I212213,I212179);
nor I_12312 (I212247,I212111,I130479);
and I_12313 (I212264,I212247,I130500);
nor I_12314 (I211967,I212264,I212060);
nor I_12315 (I212295,I130479,I130479);
nand I_12316 (I212312,I212295,I212094);
not I_12317 (I212329,I212312);
nor I_12318 (I212346,I212128,I212329);
DFFARX1 I_12319 (I212295,I2898,I211975,I211949,);
nor I_12320 (I212377,I130476,I130494);
nand I_12321 (I212394,I212060,I212377);
not I_12322 (I211943,I212394);
nor I_12323 (I212425,I130476,I130482);
DFFARX1 I_12324 (I212425,I2898,I211975,I212451,);
nor I_12325 (I212459,I212451,I212162);
nor I_12326 (I211946,I212459,I212394);
nor I_12327 (I211940,I212451,I212346);
and I_12328 (I211958,I212145,I130476);
nand I_12329 (I212518,I130503,I130497);
nor I_12330 (I212535,I212518,I130482);
not I_12331 (I212552,I212535);
nor I_12332 (I212569,I212552,I212230);
DFFARX1 I_12333 (I212569,I2898,I211975,I211961,);
nor I_12334 (I212600,I212535,I212094);
nor I_12335 (I211964,I212518,I212264);
nor I_12336 (I212631,I212035,I212518);
nand I_12337 (I211955,I212631,I130482);
not I_12338 (I212662,I212518);
nand I_12339 (I211952,I212600,I212662);
not I_12340 (I212723,I2905);
nand I_12341 (I212740,I128619,I128622);
and I_12342 (I212757,I212740,I128604);
DFFARX1 I_12343 (I212757,I2898,I212723,I212783,);
not I_12344 (I212791,I212783);
nor I_12345 (I212808,I128589,I128622);
or I_12346 (I212825,I212783,I212808);
nor I_12347 (I212842,I128601,I128598);
not I_12348 (I212859,I212842);
nor I_12349 (I212876,I212859,I212825);
nor I_12350 (I212893,I128607,I128601);
nor I_12351 (I212910,I212791,I212893);
or I_12352 (I212927,I212893,I128598);
not I_12353 (I212944,I128613);
nor I_12354 (I212961,I212944,I128592);
nor I_12355 (I212978,I212961,I212927);
nor I_12356 (I212995,I212859,I128592);
and I_12357 (I213012,I212995,I128613);
nor I_12358 (I212715,I213012,I212808);
nor I_12359 (I213043,I128592,I128592);
nand I_12360 (I213060,I213043,I212842);
not I_12361 (I213077,I213060);
nor I_12362 (I213094,I212876,I213077);
DFFARX1 I_12363 (I213043,I2898,I212723,I212697,);
nor I_12364 (I213125,I128589,I128607);
nand I_12365 (I213142,I212808,I213125);
not I_12366 (I212691,I213142);
nor I_12367 (I213173,I128589,I128595);
DFFARX1 I_12368 (I213173,I2898,I212723,I213199,);
nor I_12369 (I213207,I213199,I212910);
nor I_12370 (I212694,I213207,I213142);
nor I_12371 (I212688,I213199,I213094);
and I_12372 (I212706,I212893,I128589);
nand I_12373 (I213266,I128616,I128610);
nor I_12374 (I213283,I213266,I128595);
not I_12375 (I213300,I213283);
nor I_12376 (I213317,I213300,I212978);
DFFARX1 I_12377 (I213317,I2898,I212723,I212709,);
nor I_12378 (I213348,I213283,I212842);
nor I_12379 (I212712,I213266,I213012);
nor I_12380 (I213379,I212783,I213266);
nand I_12381 (I212703,I213379,I128595);
not I_12382 (I213410,I213266);
nand I_12383 (I212700,I213348,I213410);
not I_12384 (I213471,I2905);
nand I_12385 (I213488,I56649,I56631);
and I_12386 (I213505,I213488,I56661);
DFFARX1 I_12387 (I213505,I2898,I213471,I213531,);
not I_12388 (I213539,I213531);
nor I_12389 (I213556,I56631,I56631);
or I_12390 (I213573,I213531,I213556);
nor I_12391 (I213590,I56628,I56640);
not I_12392 (I213607,I213590);
nor I_12393 (I213624,I213607,I213573);
nor I_12394 (I213641,I56655,I56628);
nor I_12395 (I213658,I213539,I213641);
or I_12396 (I213675,I213641,I56640);
not I_12397 (I213692,I56637);
nor I_12398 (I213709,I213692,I56658);
nor I_12399 (I213726,I213709,I213675);
nor I_12400 (I213743,I213607,I56658);
and I_12401 (I213760,I213743,I56637);
nor I_12402 (I213463,I213760,I213556);
nor I_12403 (I213791,I56658,I56634);
nand I_12404 (I213808,I213791,I213590);
not I_12405 (I213825,I213808);
nor I_12406 (I213842,I213624,I213825);
DFFARX1 I_12407 (I213791,I2898,I213471,I213445,);
nor I_12408 (I213873,I56652,I56655);
nand I_12409 (I213890,I213556,I213873);
not I_12410 (I213439,I213890);
nor I_12411 (I213921,I56652,I56646);
DFFARX1 I_12412 (I213921,I2898,I213471,I213947,);
nor I_12413 (I213955,I213947,I213658);
nor I_12414 (I213442,I213955,I213890);
nor I_12415 (I213436,I213947,I213842);
and I_12416 (I213454,I213641,I56652);
nand I_12417 (I214014,I56664,I56628);
nor I_12418 (I214031,I214014,I56643);
not I_12419 (I214048,I214031);
nor I_12420 (I214065,I214048,I213726);
DFFARX1 I_12421 (I214065,I2898,I213471,I213457,);
nor I_12422 (I214096,I214031,I213590);
nor I_12423 (I213460,I214014,I213760);
nor I_12424 (I214127,I213531,I214014);
nand I_12425 (I213451,I214127,I56643);
not I_12426 (I214158,I214014);
nand I_12427 (I213448,I214096,I214158);
not I_12428 (I214219,I2905);
nand I_12429 (I214236,I182047,I182029);
and I_12430 (I214253,I214236,I182020);
DFFARX1 I_12431 (I214253,I2898,I214219,I214279,);
not I_12432 (I214287,I214279);
nor I_12433 (I214304,I182026,I182029);
or I_12434 (I214321,I214279,I214304);
nor I_12435 (I214338,I182023,I182041);
not I_12436 (I214355,I214338);
nor I_12437 (I214372,I214355,I214321);
nor I_12438 (I214389,I182038,I182023);
nor I_12439 (I214406,I214287,I214389);
or I_12440 (I214423,I214389,I182041);
not I_12441 (I214440,I182050);
nor I_12442 (I214457,I214440,I182020);
nor I_12443 (I214474,I214457,I214423);
nor I_12444 (I214491,I214355,I182020);
and I_12445 (I214508,I214491,I182050);
nor I_12446 (I214211,I214508,I214304);
nor I_12447 (I214539,I182020,I182044);
nand I_12448 (I214556,I214539,I214338);
not I_12449 (I214573,I214556);
nor I_12450 (I214590,I214372,I214573);
DFFARX1 I_12451 (I214539,I2898,I214219,I214193,);
nor I_12452 (I214621,I182026,I182038);
nand I_12453 (I214638,I214304,I214621);
not I_12454 (I214187,I214638);
nor I_12455 (I214669,I182026,I182023);
DFFARX1 I_12456 (I214669,I2898,I214219,I214695,);
nor I_12457 (I214703,I214695,I214406);
nor I_12458 (I214190,I214703,I214638);
nor I_12459 (I214184,I214695,I214590);
and I_12460 (I214202,I214389,I182026);
nand I_12461 (I214762,I182035,I182029);
nor I_12462 (I214779,I214762,I182032);
not I_12463 (I214796,I214779);
nor I_12464 (I214813,I214796,I214474);
DFFARX1 I_12465 (I214813,I2898,I214219,I214205,);
nor I_12466 (I214844,I214779,I214338);
nor I_12467 (I214208,I214762,I214508);
nor I_12468 (I214875,I214279,I214762);
nand I_12469 (I214199,I214875,I182032);
not I_12470 (I214906,I214762);
nand I_12471 (I214196,I214844,I214906);
not I_12472 (I214967,I2905);
nand I_12473 (I214984,I6601,I6580);
and I_12474 (I215001,I214984,I6595);
DFFARX1 I_12475 (I215001,I2898,I214967,I215027,);
not I_12476 (I215035,I215027);
nor I_12477 (I215052,I6583,I6580);
or I_12478 (I215069,I215027,I215052);
nor I_12479 (I215086,I6598,I6604);
not I_12480 (I215103,I215086);
nor I_12481 (I215120,I215103,I215069);
nor I_12482 (I215137,I6580,I6598);
nor I_12483 (I215154,I215035,I215137);
or I_12484 (I215171,I215137,I6604);
not I_12485 (I215188,I6583);
nor I_12486 (I215205,I215188,I6607);
nor I_12487 (I215222,I215205,I215171);
nor I_12488 (I215239,I215103,I6607);
and I_12489 (I215256,I215239,I6583);
nor I_12490 (I214959,I215256,I215052);
nor I_12491 (I215287,I6607,I6589);
nand I_12492 (I215304,I215287,I215086);
not I_12493 (I215321,I215304);
nor I_12494 (I215338,I215120,I215321);
DFFARX1 I_12495 (I215287,I2898,I214967,I214941,);
nor I_12496 (I215369,I6586,I6580);
nand I_12497 (I215386,I215052,I215369);
not I_12498 (I214935,I215386);
nor I_12499 (I215417,I6586,I6589);
DFFARX1 I_12500 (I215417,I2898,I214967,I215443,);
nor I_12501 (I215451,I215443,I215154);
nor I_12502 (I214938,I215451,I215386);
nor I_12503 (I214932,I215443,I215338);
and I_12504 (I214950,I215137,I6586);
nand I_12505 (I215510,I6592,I6610);
nor I_12506 (I215527,I215510,I6586);
not I_12507 (I215544,I215527);
nor I_12508 (I215561,I215544,I215222);
DFFARX1 I_12509 (I215561,I2898,I214967,I214953,);
nor I_12510 (I215592,I215527,I215086);
nor I_12511 (I214956,I215510,I215256);
nor I_12512 (I215623,I215027,I215510);
nand I_12513 (I214947,I215623,I6586);
not I_12514 (I215654,I215510);
nand I_12515 (I214944,I215592,I215654);
not I_12516 (I215715,I2905);
nand I_12517 (I215732,I92808,I92799);
and I_12518 (I215749,I215732,I92802);
DFFARX1 I_12519 (I215749,I2898,I215715,I215775,);
not I_12520 (I215783,I215775);
nor I_12521 (I215800,I92796,I92799);
or I_12522 (I215817,I215775,I215800);
nor I_12523 (I215834,I92811,I92796);
not I_12524 (I215851,I215834);
nor I_12525 (I215868,I215851,I215817);
nor I_12526 (I215885,I92814,I92811);
nor I_12527 (I215902,I215783,I215885);
or I_12528 (I215919,I215885,I92796);
not I_12529 (I215936,I92790);
nor I_12530 (I215953,I215936,I92805);
nor I_12531 (I215970,I215953,I215919);
nor I_12532 (I215987,I215851,I92805);
and I_12533 (I216004,I215987,I92790);
nor I_12534 (I215707,I216004,I215800);
nor I_12535 (I216035,I92805,I92793);
nand I_12536 (I216052,I216035,I215834);
not I_12537 (I216069,I216052);
nor I_12538 (I216086,I215868,I216069);
DFFARX1 I_12539 (I216035,I2898,I215715,I215689,);
nor I_12540 (I216117,I92793,I92814);
nand I_12541 (I216134,I215800,I216117);
not I_12542 (I215683,I216134);
nor I_12543 (I216165,I92793,I92787);
DFFARX1 I_12544 (I216165,I2898,I215715,I216191,);
nor I_12545 (I216199,I216191,I215902);
nor I_12546 (I215686,I216199,I216134);
nor I_12547 (I215680,I216191,I216086);
and I_12548 (I215698,I215885,I92793);
nand I_12549 (I216258,I92799,I92790);
nor I_12550 (I216275,I216258,I92787);
not I_12551 (I216292,I216275);
nor I_12552 (I216309,I216292,I215970);
DFFARX1 I_12553 (I216309,I2898,I215715,I215701,);
nor I_12554 (I216340,I216275,I215834);
nor I_12555 (I215704,I216258,I216004);
nor I_12556 (I216371,I215775,I216258);
nand I_12557 (I215695,I216371,I92787);
not I_12558 (I216402,I216258);
nand I_12559 (I215692,I216340,I216402);
not I_12560 (I216463,I2905);
nand I_12561 (I216480,I380989,I380971);
and I_12562 (I216497,I216480,I380995);
DFFARX1 I_12563 (I216497,I2898,I216463,I216523,);
not I_12564 (I216531,I216523);
nor I_12565 (I216548,I380998,I380971);
or I_12566 (I216565,I216523,I216548);
nor I_12567 (I216582,I381004,I380986);
not I_12568 (I216599,I216582);
nor I_12569 (I216616,I216599,I216565);
nor I_12570 (I216633,I380980,I381004);
nor I_12571 (I216650,I216531,I216633);
or I_12572 (I216667,I216633,I380986);
not I_12573 (I216684,I380977);
nor I_12574 (I216701,I216684,I380992);
nor I_12575 (I216718,I216701,I216667);
nor I_12576 (I216735,I216599,I380992);
and I_12577 (I216752,I216735,I380977);
nor I_12578 (I216455,I216752,I216548);
nor I_12579 (I216783,I380992,I380974);
nand I_12580 (I216800,I216783,I216582);
not I_12581 (I216817,I216800);
nor I_12582 (I216834,I216616,I216817);
DFFARX1 I_12583 (I216783,I2898,I216463,I216437,);
nor I_12584 (I216865,I380977,I380980);
nand I_12585 (I216882,I216548,I216865);
not I_12586 (I216431,I216882);
nor I_12587 (I216913,I380977,I381001);
DFFARX1 I_12588 (I216913,I2898,I216463,I216939,);
nor I_12589 (I216947,I216939,I216650);
nor I_12590 (I216434,I216947,I216882);
nor I_12591 (I216428,I216939,I216834);
and I_12592 (I216446,I216633,I380977);
nand I_12593 (I217006,I380983,I380971);
nor I_12594 (I217023,I217006,I380974);
not I_12595 (I217040,I217023);
nor I_12596 (I217057,I217040,I216718);
DFFARX1 I_12597 (I217057,I2898,I216463,I216449,);
nor I_12598 (I217088,I217023,I216582);
nor I_12599 (I216452,I217006,I216752);
nor I_12600 (I217119,I216523,I217006);
nand I_12601 (I216443,I217119,I380974);
not I_12602 (I217150,I217006);
nand I_12603 (I216440,I217088,I217150);
not I_12604 (I217211,I2905);
nand I_12605 (I217228,I25375,I25357);
and I_12606 (I217245,I217228,I25348);
DFFARX1 I_12607 (I217245,I2898,I217211,I217271,);
not I_12608 (I217279,I217271);
nor I_12609 (I217296,I25351,I25357);
or I_12610 (I217313,I217271,I217296);
nor I_12611 (I217330,I25366,I25357);
not I_12612 (I217347,I217330);
nor I_12613 (I217364,I217347,I217313);
nor I_12614 (I217381,I25363,I25366);
nor I_12615 (I217398,I217279,I217381);
or I_12616 (I217415,I217381,I25357);
not I_12617 (I217432,I25360);
nor I_12618 (I217449,I217432,I25354);
nor I_12619 (I217466,I217449,I217415);
nor I_12620 (I217483,I217347,I25354);
and I_12621 (I217500,I217483,I25360);
nor I_12622 (I217203,I217500,I217296);
nor I_12623 (I217531,I25354,I25360);
nand I_12624 (I217548,I217531,I217330);
not I_12625 (I217565,I217548);
nor I_12626 (I217582,I217364,I217565);
DFFARX1 I_12627 (I217531,I2898,I217211,I217185,);
nor I_12628 (I217613,I25372,I25363);
nand I_12629 (I217630,I217296,I217613);
not I_12630 (I217179,I217630);
nor I_12631 (I217661,I25372,I25351);
DFFARX1 I_12632 (I217661,I2898,I217211,I217687,);
nor I_12633 (I217695,I217687,I217398);
nor I_12634 (I217182,I217695,I217630);
nor I_12635 (I217176,I217687,I217582);
and I_12636 (I217194,I217381,I25372);
nand I_12637 (I217754,I25369,I25348);
nor I_12638 (I217771,I217754,I25354);
not I_12639 (I217788,I217771);
nor I_12640 (I217805,I217788,I217466);
DFFARX1 I_12641 (I217805,I2898,I217211,I217197,);
nor I_12642 (I217836,I217771,I217330);
nor I_12643 (I217200,I217754,I217500);
nor I_12644 (I217867,I217271,I217754);
nand I_12645 (I217191,I217867,I25354);
not I_12646 (I217898,I217754);
nand I_12647 (I217188,I217836,I217898);
not I_12648 (I217959,I2905);
nand I_12649 (I217976,I345444,I345441);
and I_12650 (I217993,I217976,I345450);
DFFARX1 I_12651 (I217993,I2898,I217959,I218019,);
not I_12652 (I218027,I218019);
nor I_12653 (I218044,I345447,I345441);
or I_12654 (I218061,I218019,I218044);
nor I_12655 (I218078,I345456,I345450);
not I_12656 (I218095,I218078);
nor I_12657 (I218112,I218095,I218061);
nor I_12658 (I218129,I345444,I345456);
nor I_12659 (I218146,I218027,I218129);
or I_12660 (I218163,I218129,I345450);
not I_12661 (I218180,I345447);
nor I_12662 (I218197,I218180,I345441);
nor I_12663 (I218214,I218197,I218163);
nor I_12664 (I218231,I218095,I345441);
and I_12665 (I218248,I218231,I345447);
nor I_12666 (I217951,I218248,I218044);
nor I_12667 (I218279,I345441,I345459);
nand I_12668 (I218296,I218279,I218078);
not I_12669 (I218313,I218296);
nor I_12670 (I218330,I218112,I218313);
DFFARX1 I_12671 (I218279,I2898,I217959,I217933,);
nor I_12672 (I218361,I345453,I345444);
nand I_12673 (I218378,I218044,I218361);
not I_12674 (I217927,I218378);
nor I_12675 (I218409,I345453,I345465);
DFFARX1 I_12676 (I218409,I2898,I217959,I218435,);
nor I_12677 (I218443,I218435,I218146);
nor I_12678 (I217930,I218443,I218378);
nor I_12679 (I217924,I218435,I218330);
and I_12680 (I217942,I218129,I345453);
nand I_12681 (I218502,I345453,I345462);
nor I_12682 (I218519,I218502,I345456);
not I_12683 (I218536,I218519);
nor I_12684 (I218553,I218536,I218214);
DFFARX1 I_12685 (I218553,I2898,I217959,I217945,);
nor I_12686 (I218584,I218519,I218078);
nor I_12687 (I217948,I218502,I218248);
nor I_12688 (I218615,I218019,I218502);
nand I_12689 (I217939,I218615,I345456);
not I_12690 (I218646,I218502);
nand I_12691 (I217936,I218584,I218646);
not I_12692 (I218707,I2905);
nand I_12693 (I218724,I393263,I393245);
and I_12694 (I218741,I218724,I393269);
DFFARX1 I_12695 (I218741,I2898,I218707,I218767,);
not I_12696 (I218775,I218767);
nor I_12697 (I218792,I393272,I393245);
or I_12698 (I218809,I218767,I218792);
nor I_12699 (I218826,I393278,I393260);
not I_12700 (I218843,I218826);
nor I_12701 (I218860,I218843,I218809);
nor I_12702 (I218877,I393254,I393278);
nor I_12703 (I218894,I218775,I218877);
or I_12704 (I218911,I218877,I393260);
not I_12705 (I218928,I393251);
nor I_12706 (I218945,I218928,I393266);
nor I_12707 (I218962,I218945,I218911);
nor I_12708 (I218979,I218843,I393266);
and I_12709 (I218996,I218979,I393251);
nor I_12710 (I218699,I218996,I218792);
nor I_12711 (I219027,I393266,I393248);
nand I_12712 (I219044,I219027,I218826);
not I_12713 (I219061,I219044);
nor I_12714 (I219078,I218860,I219061);
DFFARX1 I_12715 (I219027,I2898,I218707,I218681,);
nor I_12716 (I219109,I393251,I393254);
nand I_12717 (I219126,I218792,I219109);
not I_12718 (I218675,I219126);
nor I_12719 (I219157,I393251,I393275);
DFFARX1 I_12720 (I219157,I2898,I218707,I219183,);
nor I_12721 (I219191,I219183,I218894);
nor I_12722 (I218678,I219191,I219126);
nor I_12723 (I218672,I219183,I219078);
and I_12724 (I218690,I218877,I393251);
nand I_12725 (I219250,I393257,I393245);
nor I_12726 (I219267,I219250,I393248);
not I_12727 (I219284,I219267);
nor I_12728 (I219301,I219284,I218962);
DFFARX1 I_12729 (I219301,I2898,I218707,I218693,);
nor I_12730 (I219332,I219267,I218826);
nor I_12731 (I218696,I219250,I218996);
nor I_12732 (I219363,I218767,I219250);
nand I_12733 (I218687,I219363,I393248);
not I_12734 (I219394,I219250);
nand I_12735 (I218684,I219332,I219394);
not I_12736 (I219455,I2905);
nand I_12737 (I219472,I89034,I89025);
and I_12738 (I219489,I219472,I89028);
DFFARX1 I_12739 (I219489,I2898,I219455,I219515,);
not I_12740 (I219523,I219515);
nor I_12741 (I219540,I89022,I89025);
or I_12742 (I219557,I219515,I219540);
nor I_12743 (I219574,I89037,I89022);
not I_12744 (I219591,I219574);
nor I_12745 (I219608,I219591,I219557);
nor I_12746 (I219625,I89040,I89037);
nor I_12747 (I219642,I219523,I219625);
or I_12748 (I219659,I219625,I89022);
not I_12749 (I219676,I89016);
nor I_12750 (I219693,I219676,I89031);
nor I_12751 (I219710,I219693,I219659);
nor I_12752 (I219727,I219591,I89031);
and I_12753 (I219744,I219727,I89016);
nor I_12754 (I219447,I219744,I219540);
nor I_12755 (I219775,I89031,I89019);
nand I_12756 (I219792,I219775,I219574);
not I_12757 (I219809,I219792);
nor I_12758 (I219826,I219608,I219809);
DFFARX1 I_12759 (I219775,I2898,I219455,I219429,);
nor I_12760 (I219857,I89019,I89040);
nand I_12761 (I219874,I219540,I219857);
not I_12762 (I219423,I219874);
nor I_12763 (I219905,I89019,I89013);
DFFARX1 I_12764 (I219905,I2898,I219455,I219931,);
nor I_12765 (I219939,I219931,I219642);
nor I_12766 (I219426,I219939,I219874);
nor I_12767 (I219420,I219931,I219826);
and I_12768 (I219438,I219625,I89019);
nand I_12769 (I219998,I89025,I89016);
nor I_12770 (I220015,I219998,I89013);
not I_12771 (I220032,I220015);
nor I_12772 (I220049,I220032,I219710);
DFFARX1 I_12773 (I220049,I2898,I219455,I219441,);
nor I_12774 (I220080,I220015,I219574);
nor I_12775 (I219444,I219998,I219744);
nor I_12776 (I220111,I219515,I219998);
nand I_12777 (I219435,I220111,I89013);
not I_12778 (I220142,I219998);
nand I_12779 (I219432,I220080,I220142);
not I_12780 (I220203,I2905);
nand I_12781 (I220220,I320049,I320046);
and I_12782 (I220237,I220220,I320043);
DFFARX1 I_12783 (I220237,I2898,I220203,I220263,);
not I_12784 (I220271,I220263);
nor I_12785 (I220288,I320052,I320046);
or I_12786 (I220305,I220263,I220288);
nor I_12787 (I220322,I320070,I320043);
not I_12788 (I220339,I220322);
nor I_12789 (I220356,I220339,I220305);
nor I_12790 (I220373,I320073,I320070);
nor I_12791 (I220390,I220271,I220373);
or I_12792 (I220407,I220373,I320043);
not I_12793 (I220424,I320058);
nor I_12794 (I220441,I220424,I320064);
nor I_12795 (I220458,I220441,I220407);
nor I_12796 (I220475,I220339,I320064);
and I_12797 (I220492,I220475,I320058);
nor I_12798 (I220195,I220492,I220288);
nor I_12799 (I220523,I320064,I320052);
nand I_12800 (I220540,I220523,I220322);
not I_12801 (I220557,I220540);
nor I_12802 (I220574,I220356,I220557);
DFFARX1 I_12803 (I220523,I2898,I220203,I220177,);
nor I_12804 (I220605,I320049,I320073);
nand I_12805 (I220622,I220288,I220605);
not I_12806 (I220171,I220622);
nor I_12807 (I220653,I320049,I320046);
DFFARX1 I_12808 (I220653,I2898,I220203,I220679,);
nor I_12809 (I220687,I220679,I220390);
nor I_12810 (I220174,I220687,I220622);
nor I_12811 (I220168,I220679,I220574);
and I_12812 (I220186,I220373,I320049);
nand I_12813 (I220746,I320055,I320061);
nor I_12814 (I220763,I220746,I320067);
not I_12815 (I220780,I220763);
nor I_12816 (I220797,I220780,I220458);
DFFARX1 I_12817 (I220797,I2898,I220203,I220189,);
nor I_12818 (I220828,I220763,I220322);
nor I_12819 (I220192,I220746,I220492);
nor I_12820 (I220859,I220263,I220746);
nand I_12821 (I220183,I220859,I320067);
not I_12822 (I220890,I220746);
nand I_12823 (I220180,I220828,I220890);
not I_12824 (I220951,I2905);
nand I_12825 (I220968,I393909,I393891);
and I_12826 (I220985,I220968,I393915);
DFFARX1 I_12827 (I220985,I2898,I220951,I221011,);
not I_12828 (I221019,I221011);
nor I_12829 (I221036,I393918,I393891);
or I_12830 (I221053,I221011,I221036);
nor I_12831 (I221070,I393924,I393906);
not I_12832 (I221087,I221070);
nor I_12833 (I221104,I221087,I221053);
nor I_12834 (I221121,I393900,I393924);
nor I_12835 (I221138,I221019,I221121);
or I_12836 (I221155,I221121,I393906);
not I_12837 (I221172,I393897);
nor I_12838 (I221189,I221172,I393912);
nor I_12839 (I221206,I221189,I221155);
nor I_12840 (I221223,I221087,I393912);
and I_12841 (I221240,I221223,I393897);
nor I_12842 (I220943,I221240,I221036);
nor I_12843 (I221271,I393912,I393894);
nand I_12844 (I221288,I221271,I221070);
not I_12845 (I221305,I221288);
nor I_12846 (I221322,I221104,I221305);
DFFARX1 I_12847 (I221271,I2898,I220951,I220925,);
nor I_12848 (I221353,I393897,I393900);
nand I_12849 (I221370,I221036,I221353);
not I_12850 (I220919,I221370);
nor I_12851 (I221401,I393897,I393921);
DFFARX1 I_12852 (I221401,I2898,I220951,I221427,);
nor I_12853 (I221435,I221427,I221138);
nor I_12854 (I220922,I221435,I221370);
nor I_12855 (I220916,I221427,I221322);
and I_12856 (I220934,I221121,I393897);
nand I_12857 (I221494,I393903,I393891);
nor I_12858 (I221511,I221494,I393894);
not I_12859 (I221528,I221511);
nor I_12860 (I221545,I221528,I221206);
DFFARX1 I_12861 (I221545,I2898,I220951,I220937,);
nor I_12862 (I221576,I221511,I221070);
nor I_12863 (I220940,I221494,I221240);
nor I_12864 (I221607,I221011,I221494);
nand I_12865 (I220931,I221607,I393894);
not I_12866 (I221638,I221494);
nand I_12867 (I220928,I221576,I221638);
not I_12868 (I221699,I2905);
nand I_12869 (I221716,I28231,I28213);
and I_12870 (I221733,I221716,I28204);
DFFARX1 I_12871 (I221733,I2898,I221699,I221759,);
not I_12872 (I221767,I221759);
nor I_12873 (I221784,I28207,I28213);
or I_12874 (I221801,I221759,I221784);
nor I_12875 (I221818,I28222,I28213);
not I_12876 (I221835,I221818);
nor I_12877 (I221852,I221835,I221801);
nor I_12878 (I221869,I28219,I28222);
nor I_12879 (I221886,I221767,I221869);
or I_12880 (I221903,I221869,I28213);
not I_12881 (I221920,I28216);
nor I_12882 (I221937,I221920,I28210);
nor I_12883 (I221954,I221937,I221903);
nor I_12884 (I221971,I221835,I28210);
and I_12885 (I221988,I221971,I28216);
nor I_12886 (I221691,I221988,I221784);
nor I_12887 (I222019,I28210,I28216);
nand I_12888 (I222036,I222019,I221818);
not I_12889 (I222053,I222036);
nor I_12890 (I222070,I221852,I222053);
DFFARX1 I_12891 (I222019,I2898,I221699,I221673,);
nor I_12892 (I222101,I28228,I28219);
nand I_12893 (I222118,I221784,I222101);
not I_12894 (I221667,I222118);
nor I_12895 (I222149,I28228,I28207);
DFFARX1 I_12896 (I222149,I2898,I221699,I222175,);
nor I_12897 (I222183,I222175,I221886);
nor I_12898 (I221670,I222183,I222118);
nor I_12899 (I221664,I222175,I222070);
and I_12900 (I221682,I221869,I28228);
nand I_12901 (I222242,I28225,I28204);
nor I_12902 (I222259,I222242,I28210);
not I_12903 (I222276,I222259);
nor I_12904 (I222293,I222276,I221954);
DFFARX1 I_12905 (I222293,I2898,I221699,I221685,);
nor I_12906 (I222324,I222259,I221818);
nor I_12907 (I221688,I222242,I221988);
nor I_12908 (I222355,I221759,I222242);
nand I_12909 (I221679,I222355,I28210);
not I_12910 (I222386,I222242);
nand I_12911 (I221676,I222324,I222386);
not I_12912 (I222447,I2905);
nand I_12913 (I222464,I141199,I141202);
and I_12914 (I222481,I222464,I141184);
DFFARX1 I_12915 (I222481,I2898,I222447,I222507,);
not I_12916 (I222515,I222507);
nor I_12917 (I222532,I141169,I141202);
or I_12918 (I222549,I222507,I222532);
nor I_12919 (I222566,I141181,I141178);
not I_12920 (I222583,I222566);
nor I_12921 (I222600,I222583,I222549);
nor I_12922 (I222617,I141187,I141181);
nor I_12923 (I222634,I222515,I222617);
or I_12924 (I222651,I222617,I141178);
not I_12925 (I222668,I141193);
nor I_12926 (I222685,I222668,I141172);
nor I_12927 (I222702,I222685,I222651);
nor I_12928 (I222719,I222583,I141172);
and I_12929 (I222736,I222719,I141193);
nor I_12930 (I222439,I222736,I222532);
nor I_12931 (I222767,I141172,I141172);
nand I_12932 (I222784,I222767,I222566);
not I_12933 (I222801,I222784);
nor I_12934 (I222818,I222600,I222801);
DFFARX1 I_12935 (I222767,I2898,I222447,I222421,);
nor I_12936 (I222849,I141169,I141187);
nand I_12937 (I222866,I222532,I222849);
not I_12938 (I222415,I222866);
nor I_12939 (I222897,I141169,I141175);
DFFARX1 I_12940 (I222897,I2898,I222447,I222923,);
nor I_12941 (I222931,I222923,I222634);
nor I_12942 (I222418,I222931,I222866);
nor I_12943 (I222412,I222923,I222818);
and I_12944 (I222430,I222617,I141169);
nand I_12945 (I222990,I141196,I141190);
nor I_12946 (I223007,I222990,I141175);
not I_12947 (I223024,I223007);
nor I_12948 (I223041,I223024,I222702);
DFFARX1 I_12949 (I223041,I2898,I222447,I222433,);
nor I_12950 (I223072,I223007,I222566);
nor I_12951 (I222436,I222990,I222736);
nor I_12952 (I223103,I222507,I222990);
nand I_12953 (I222427,I223103,I141175);
not I_12954 (I223134,I222990);
nand I_12955 (I222424,I223072,I223134);
not I_12956 (I223195,I2905);
nand I_12957 (I223212,I382281,I382263);
and I_12958 (I223229,I223212,I382287);
DFFARX1 I_12959 (I223229,I2898,I223195,I223255,);
not I_12960 (I223263,I223255);
nor I_12961 (I223280,I382290,I382263);
or I_12962 (I223297,I223255,I223280);
nor I_12963 (I223314,I382296,I382278);
not I_12964 (I223331,I223314);
nor I_12965 (I223348,I223331,I223297);
nor I_12966 (I223365,I382272,I382296);
nor I_12967 (I223382,I223263,I223365);
or I_12968 (I223399,I223365,I382278);
not I_12969 (I223416,I382269);
nor I_12970 (I223433,I223416,I382284);
nor I_12971 (I223450,I223433,I223399);
nor I_12972 (I223467,I223331,I382284);
and I_12973 (I223484,I223467,I382269);
nor I_12974 (I223187,I223484,I223280);
nor I_12975 (I223515,I382284,I382266);
nand I_12976 (I223532,I223515,I223314);
not I_12977 (I223549,I223532);
nor I_12978 (I223566,I223348,I223549);
DFFARX1 I_12979 (I223515,I2898,I223195,I223169,);
nor I_12980 (I223597,I382269,I382272);
nand I_12981 (I223614,I223280,I223597);
not I_12982 (I223163,I223614);
nor I_12983 (I223645,I382269,I382293);
DFFARX1 I_12984 (I223645,I2898,I223195,I223671,);
nor I_12985 (I223679,I223671,I223382);
nor I_12986 (I223166,I223679,I223614);
nor I_12987 (I223160,I223671,I223566);
and I_12988 (I223178,I223365,I382269);
nand I_12989 (I223738,I382275,I382263);
nor I_12990 (I223755,I223738,I382266);
not I_12991 (I223772,I223755);
nor I_12992 (I223789,I223772,I223450);
DFFARX1 I_12993 (I223789,I2898,I223195,I223181,);
nor I_12994 (I223820,I223755,I223314);
nor I_12995 (I223184,I223738,I223484);
nor I_12996 (I223851,I223255,I223738);
nand I_12997 (I223175,I223851,I382266);
not I_12998 (I223882,I223738);
nand I_12999 (I223172,I223820,I223882);
not I_13000 (I223943,I2905);
nand I_13001 (I223960,I23947,I23929);
and I_13002 (I223977,I223960,I23920);
DFFARX1 I_13003 (I223977,I2898,I223943,I224003,);
not I_13004 (I224011,I224003);
nor I_13005 (I224028,I23923,I23929);
or I_13006 (I224045,I224003,I224028);
nor I_13007 (I224062,I23938,I23929);
not I_13008 (I224079,I224062);
nor I_13009 (I224096,I224079,I224045);
nor I_13010 (I224113,I23935,I23938);
nor I_13011 (I224130,I224011,I224113);
or I_13012 (I224147,I224113,I23929);
not I_13013 (I224164,I23932);
nor I_13014 (I224181,I224164,I23926);
nor I_13015 (I224198,I224181,I224147);
nor I_13016 (I224215,I224079,I23926);
and I_13017 (I224232,I224215,I23932);
nor I_13018 (I223935,I224232,I224028);
nor I_13019 (I224263,I23926,I23932);
nand I_13020 (I224280,I224263,I224062);
not I_13021 (I224297,I224280);
nor I_13022 (I224314,I224096,I224297);
DFFARX1 I_13023 (I224263,I2898,I223943,I223917,);
nor I_13024 (I224345,I23944,I23935);
nand I_13025 (I224362,I224028,I224345);
not I_13026 (I223911,I224362);
nor I_13027 (I224393,I23944,I23923);
DFFARX1 I_13028 (I224393,I2898,I223943,I224419,);
nor I_13029 (I224427,I224419,I224130);
nor I_13030 (I223914,I224427,I224362);
nor I_13031 (I223908,I224419,I224314);
and I_13032 (I223926,I224113,I23944);
nand I_13033 (I224486,I23941,I23920);
nor I_13034 (I224503,I224486,I23926);
not I_13035 (I224520,I224503);
nor I_13036 (I224537,I224520,I224198);
DFFARX1 I_13037 (I224537,I2898,I223943,I223929,);
nor I_13038 (I224568,I224503,I224062);
nor I_13039 (I223932,I224486,I224232);
nor I_13040 (I224599,I224003,I224486);
nand I_13041 (I223923,I224599,I23926);
not I_13042 (I224630,I224486);
nand I_13043 (I223920,I224568,I224630);
not I_13044 (I224691,I2905);
nand I_13045 (I224708,I311277,I311274);
and I_13046 (I224725,I224708,I311271);
DFFARX1 I_13047 (I224725,I2898,I224691,I224751,);
not I_13048 (I224759,I224751);
nor I_13049 (I224776,I311280,I311274);
or I_13050 (I224793,I224751,I224776);
nor I_13051 (I224810,I311298,I311271);
not I_13052 (I224827,I224810);
nor I_13053 (I224844,I224827,I224793);
nor I_13054 (I224861,I311301,I311298);
nor I_13055 (I224878,I224759,I224861);
or I_13056 (I224895,I224861,I311271);
not I_13057 (I224912,I311286);
nor I_13058 (I224929,I224912,I311292);
nor I_13059 (I224946,I224929,I224895);
nor I_13060 (I224963,I224827,I311292);
and I_13061 (I224980,I224963,I311286);
nor I_13062 (I224683,I224980,I224776);
nor I_13063 (I225011,I311292,I311280);
nand I_13064 (I225028,I225011,I224810);
not I_13065 (I225045,I225028);
nor I_13066 (I225062,I224844,I225045);
DFFARX1 I_13067 (I225011,I2898,I224691,I224665,);
nor I_13068 (I225093,I311277,I311301);
nand I_13069 (I225110,I224776,I225093);
not I_13070 (I224659,I225110);
nor I_13071 (I225141,I311277,I311274);
DFFARX1 I_13072 (I225141,I2898,I224691,I225167,);
nor I_13073 (I225175,I225167,I224878);
nor I_13074 (I224662,I225175,I225110);
nor I_13075 (I224656,I225167,I225062);
and I_13076 (I224674,I224861,I311277);
nand I_13077 (I225234,I311283,I311289);
nor I_13078 (I225251,I225234,I311295);
not I_13079 (I225268,I225251);
nor I_13080 (I225285,I225268,I224946);
DFFARX1 I_13081 (I225285,I2898,I224691,I224677,);
nor I_13082 (I225316,I225251,I224810);
nor I_13083 (I224680,I225234,I224980);
nor I_13084 (I225347,I224751,I225234);
nand I_13085 (I224671,I225347,I311295);
not I_13086 (I225378,I225234);
nand I_13087 (I224668,I225316,I225378);
not I_13088 (I225439,I2905);
nand I_13089 (I225456,I60100,I60091);
and I_13090 (I225473,I225456,I60094);
DFFARX1 I_13091 (I225473,I2898,I225439,I225499,);
not I_13092 (I225507,I225499);
nor I_13093 (I225524,I60088,I60091);
or I_13094 (I225541,I225499,I225524);
nor I_13095 (I225558,I60103,I60088);
not I_13096 (I225575,I225558);
nor I_13097 (I225592,I225575,I225541);
nor I_13098 (I225609,I60106,I60103);
nor I_13099 (I225626,I225507,I225609);
or I_13100 (I225643,I225609,I60088);
not I_13101 (I225660,I60082);
nor I_13102 (I225677,I225660,I60097);
nor I_13103 (I225694,I225677,I225643);
nor I_13104 (I225711,I225575,I60097);
and I_13105 (I225728,I225711,I60082);
nor I_13106 (I225431,I225728,I225524);
nor I_13107 (I225759,I60097,I60085);
nand I_13108 (I225776,I225759,I225558);
not I_13109 (I225793,I225776);
nor I_13110 (I225810,I225592,I225793);
DFFARX1 I_13111 (I225759,I2898,I225439,I225413,);
nor I_13112 (I225841,I60085,I60106);
nand I_13113 (I225858,I225524,I225841);
not I_13114 (I225407,I225858);
nor I_13115 (I225889,I60085,I60079);
DFFARX1 I_13116 (I225889,I2898,I225439,I225915,);
nor I_13117 (I225923,I225915,I225626);
nor I_13118 (I225410,I225923,I225858);
nor I_13119 (I225404,I225915,I225810);
and I_13120 (I225422,I225609,I60085);
nand I_13121 (I225982,I60091,I60082);
nor I_13122 (I225999,I225982,I60079);
not I_13123 (I226016,I225999);
nor I_13124 (I226033,I226016,I225694);
DFFARX1 I_13125 (I226033,I2898,I225439,I225425,);
nor I_13126 (I226064,I225999,I225558);
nor I_13127 (I225428,I225982,I225728);
nor I_13128 (I226095,I225499,I225982);
nand I_13129 (I225419,I226095,I60079);
not I_13130 (I226126,I225982);
nand I_13131 (I225416,I226064,I226126);
not I_13132 (I226187,I2905);
nand I_13133 (I226204,I329974,I329971);
and I_13134 (I226221,I226204,I329980);
DFFARX1 I_13135 (I226221,I2898,I226187,I226247,);
not I_13136 (I226255,I226247);
nor I_13137 (I226272,I329977,I329971);
or I_13138 (I226289,I226247,I226272);
nor I_13139 (I226306,I329986,I329980);
not I_13140 (I226323,I226306);
nor I_13141 (I226340,I226323,I226289);
nor I_13142 (I226357,I329974,I329986);
nor I_13143 (I226374,I226255,I226357);
or I_13144 (I226391,I226357,I329980);
not I_13145 (I226408,I329977);
nor I_13146 (I226425,I226408,I329971);
nor I_13147 (I226442,I226425,I226391);
nor I_13148 (I226459,I226323,I329971);
and I_13149 (I226476,I226459,I329977);
nor I_13150 (I226179,I226476,I226272);
nor I_13151 (I226507,I329971,I329989);
nand I_13152 (I226524,I226507,I226306);
not I_13153 (I226541,I226524);
nor I_13154 (I226558,I226340,I226541);
DFFARX1 I_13155 (I226507,I2898,I226187,I226161,);
nor I_13156 (I226589,I329983,I329974);
nand I_13157 (I226606,I226272,I226589);
not I_13158 (I226155,I226606);
nor I_13159 (I226637,I329983,I329995);
DFFARX1 I_13160 (I226637,I2898,I226187,I226663,);
nor I_13161 (I226671,I226663,I226374);
nor I_13162 (I226158,I226671,I226606);
nor I_13163 (I226152,I226663,I226558);
and I_13164 (I226170,I226357,I329983);
nand I_13165 (I226730,I329983,I329992);
nor I_13166 (I226747,I226730,I329986);
not I_13167 (I226764,I226747);
nor I_13168 (I226781,I226764,I226442);
DFFARX1 I_13169 (I226781,I2898,I226187,I226173,);
nor I_13170 (I226812,I226747,I226306);
nor I_13171 (I226176,I226730,I226476);
nor I_13172 (I226843,I226247,I226730);
nand I_13173 (I226167,I226843,I329986);
not I_13174 (I226874,I226730);
nand I_13175 (I226164,I226812,I226874);
not I_13176 (I226935,I2905);
nand I_13177 (I226952,I389387,I389369);
and I_13178 (I226969,I226952,I389393);
DFFARX1 I_13179 (I226969,I2898,I226935,I226995,);
not I_13180 (I227003,I226995);
nor I_13181 (I227020,I389396,I389369);
or I_13182 (I227037,I226995,I227020);
nor I_13183 (I227054,I389402,I389384);
not I_13184 (I227071,I227054);
nor I_13185 (I227088,I227071,I227037);
nor I_13186 (I227105,I389378,I389402);
nor I_13187 (I227122,I227003,I227105);
or I_13188 (I227139,I227105,I389384);
not I_13189 (I227156,I389375);
nor I_13190 (I227173,I227156,I389390);
nor I_13191 (I227190,I227173,I227139);
nor I_13192 (I227207,I227071,I389390);
and I_13193 (I227224,I227207,I389375);
nor I_13194 (I226927,I227224,I227020);
nor I_13195 (I227255,I389390,I389372);
nand I_13196 (I227272,I227255,I227054);
not I_13197 (I227289,I227272);
nor I_13198 (I227306,I227088,I227289);
DFFARX1 I_13199 (I227255,I2898,I226935,I226909,);
nor I_13200 (I227337,I389375,I389378);
nand I_13201 (I227354,I227020,I227337);
not I_13202 (I226903,I227354);
nor I_13203 (I227385,I389375,I389399);
DFFARX1 I_13204 (I227385,I2898,I226935,I227411,);
nor I_13205 (I227419,I227411,I227122);
nor I_13206 (I226906,I227419,I227354);
nor I_13207 (I226900,I227411,I227306);
and I_13208 (I226918,I227105,I389375);
nand I_13209 (I227478,I389381,I389369);
nor I_13210 (I227495,I227478,I389372);
not I_13211 (I227512,I227495);
nor I_13212 (I227529,I227512,I227190);
DFFARX1 I_13213 (I227529,I2898,I226935,I226921,);
nor I_13214 (I227560,I227495,I227054);
nor I_13215 (I226924,I227478,I227224);
nor I_13216 (I227591,I226995,I227478);
nand I_13217 (I226915,I227591,I389372);
not I_13218 (I227622,I227478);
nand I_13219 (I226912,I227560,I227622);
not I_13220 (I227683,I2905);
nand I_13221 (I227700,I288616,I288613);
and I_13222 (I227717,I227700,I288610);
DFFARX1 I_13223 (I227717,I2898,I227683,I227743,);
not I_13224 (I227751,I227743);
nor I_13225 (I227768,I288619,I288613);
or I_13226 (I227785,I227743,I227768);
nor I_13227 (I227802,I288637,I288610);
not I_13228 (I227819,I227802);
nor I_13229 (I227836,I227819,I227785);
nor I_13230 (I227853,I288640,I288637);
nor I_13231 (I227870,I227751,I227853);
or I_13232 (I227887,I227853,I288610);
not I_13233 (I227904,I288625);
nor I_13234 (I227921,I227904,I288631);
nor I_13235 (I227938,I227921,I227887);
nor I_13236 (I227955,I227819,I288631);
and I_13237 (I227972,I227955,I288625);
nor I_13238 (I227675,I227972,I227768);
nor I_13239 (I228003,I288631,I288619);
nand I_13240 (I228020,I228003,I227802);
not I_13241 (I228037,I228020);
nor I_13242 (I228054,I227836,I228037);
DFFARX1 I_13243 (I228003,I2898,I227683,I227657,);
nor I_13244 (I228085,I288616,I288640);
nand I_13245 (I228102,I227768,I228085);
not I_13246 (I227651,I228102);
nor I_13247 (I228133,I288616,I288613);
DFFARX1 I_13248 (I228133,I2898,I227683,I228159,);
nor I_13249 (I228167,I228159,I227870);
nor I_13250 (I227654,I228167,I228102);
nor I_13251 (I227648,I228159,I228054);
and I_13252 (I227666,I227853,I288616);
nand I_13253 (I228226,I288622,I288628);
nor I_13254 (I228243,I228226,I288634);
not I_13255 (I228260,I228243);
nor I_13256 (I228277,I228260,I227938);
DFFARX1 I_13257 (I228277,I2898,I227683,I227669,);
nor I_13258 (I228308,I228243,I227802);
nor I_13259 (I227672,I228226,I227972);
nor I_13260 (I228339,I227743,I228226);
nand I_13261 (I227663,I228339,I288634);
not I_13262 (I228370,I228226);
nand I_13263 (I227660,I228308,I228370);
not I_13264 (I228431,I2905);
nand I_13265 (I228448,I312008,I312005);
and I_13266 (I228465,I228448,I312002);
DFFARX1 I_13267 (I228465,I2898,I228431,I228491,);
not I_13268 (I228499,I228491);
nor I_13269 (I228516,I312011,I312005);
or I_13270 (I228533,I228491,I228516);
nor I_13271 (I228550,I312029,I312002);
not I_13272 (I228567,I228550);
nor I_13273 (I228584,I228567,I228533);
nor I_13274 (I228601,I312032,I312029);
nor I_13275 (I228618,I228499,I228601);
or I_13276 (I228635,I228601,I312002);
not I_13277 (I228652,I312017);
nor I_13278 (I228669,I228652,I312023);
nor I_13279 (I228686,I228669,I228635);
nor I_13280 (I228703,I228567,I312023);
and I_13281 (I228720,I228703,I312017);
nor I_13282 (I228423,I228720,I228516);
nor I_13283 (I228751,I312023,I312011);
nand I_13284 (I228768,I228751,I228550);
not I_13285 (I228785,I228768);
nor I_13286 (I228802,I228584,I228785);
DFFARX1 I_13287 (I228751,I2898,I228431,I228405,);
nor I_13288 (I228833,I312008,I312032);
nand I_13289 (I228850,I228516,I228833);
not I_13290 (I228399,I228850);
nor I_13291 (I228881,I312008,I312005);
DFFARX1 I_13292 (I228881,I2898,I228431,I228907,);
nor I_13293 (I228915,I228907,I228618);
nor I_13294 (I228402,I228915,I228850);
nor I_13295 (I228396,I228907,I228802);
and I_13296 (I228414,I228601,I312008);
nand I_13297 (I228974,I312014,I312020);
nor I_13298 (I228991,I228974,I312026);
not I_13299 (I229008,I228991);
nor I_13300 (I229025,I229008,I228686);
DFFARX1 I_13301 (I229025,I2898,I228431,I228417,);
nor I_13302 (I229056,I228991,I228550);
nor I_13303 (I228420,I228974,I228720);
nor I_13304 (I229087,I228491,I228974);
nand I_13305 (I228411,I229087,I312026);
not I_13306 (I229118,I228974);
nand I_13307 (I228408,I229056,I229118);
not I_13308 (I229179,I2905);
nand I_13309 (I229196,I310546,I310543);
and I_13310 (I229213,I229196,I310540);
DFFARX1 I_13311 (I229213,I2898,I229179,I229239,);
not I_13312 (I229247,I229239);
nor I_13313 (I229264,I310549,I310543);
or I_13314 (I229281,I229239,I229264);
nor I_13315 (I229298,I310567,I310540);
not I_13316 (I229315,I229298);
nor I_13317 (I229332,I229315,I229281);
nor I_13318 (I229349,I310570,I310567);
nor I_13319 (I229366,I229247,I229349);
or I_13320 (I229383,I229349,I310540);
not I_13321 (I229400,I310555);
nor I_13322 (I229417,I229400,I310561);
nor I_13323 (I229434,I229417,I229383);
nor I_13324 (I229451,I229315,I310561);
and I_13325 (I229468,I229451,I310555);
nor I_13326 (I229171,I229468,I229264);
nor I_13327 (I229499,I310561,I310549);
nand I_13328 (I229516,I229499,I229298);
not I_13329 (I229533,I229516);
nor I_13330 (I229550,I229332,I229533);
DFFARX1 I_13331 (I229499,I2898,I229179,I229153,);
nor I_13332 (I229581,I310546,I310570);
nand I_13333 (I229598,I229264,I229581);
not I_13334 (I229147,I229598);
nor I_13335 (I229629,I310546,I310543);
DFFARX1 I_13336 (I229629,I2898,I229179,I229655,);
nor I_13337 (I229663,I229655,I229366);
nor I_13338 (I229150,I229663,I229598);
nor I_13339 (I229144,I229655,I229550);
and I_13340 (I229162,I229349,I310546);
nand I_13341 (I229722,I310552,I310558);
nor I_13342 (I229739,I229722,I310564);
not I_13343 (I229756,I229739);
nor I_13344 (I229773,I229756,I229434);
DFFARX1 I_13345 (I229773,I2898,I229179,I229165,);
nor I_13346 (I229804,I229739,I229298);
nor I_13347 (I229168,I229722,I229468);
nor I_13348 (I229835,I229239,I229722);
nand I_13349 (I229159,I229835,I310564);
not I_13350 (I229866,I229722);
nand I_13351 (I229156,I229804,I229866);
not I_13352 (I229927,I2905);
nand I_13353 (I229944,I281916,I281901);
and I_13354 (I229961,I229944,I281895);
DFFARX1 I_13355 (I229961,I2898,I229927,I229987,);
not I_13356 (I229995,I229987);
nor I_13357 (I230012,I281898,I281901);
or I_13358 (I230029,I229987,I230012);
nor I_13359 (I230046,I281925,I281919);
not I_13360 (I230063,I230046);
nor I_13361 (I230080,I230063,I230029);
nor I_13362 (I230097,I281922,I281925);
nor I_13363 (I230114,I229995,I230097);
or I_13364 (I230131,I230097,I281919);
not I_13365 (I230148,I281910);
nor I_13366 (I230165,I230148,I281901);
nor I_13367 (I230182,I230165,I230131);
nor I_13368 (I230199,I230063,I281901);
and I_13369 (I230216,I230199,I281910);
nor I_13370 (I229919,I230216,I230012);
nor I_13371 (I230247,I281901,I281904);
nand I_13372 (I230264,I230247,I230046);
not I_13373 (I230281,I230264);
nor I_13374 (I230298,I230080,I230281);
DFFARX1 I_13375 (I230247,I2898,I229927,I229901,);
nor I_13376 (I230329,I281907,I281922);
nand I_13377 (I230346,I230012,I230329);
not I_13378 (I229895,I230346);
nor I_13379 (I230377,I281907,I281904);
DFFARX1 I_13380 (I230377,I2898,I229927,I230403,);
nor I_13381 (I230411,I230403,I230114);
nor I_13382 (I229898,I230411,I230346);
nor I_13383 (I229892,I230403,I230298);
and I_13384 (I229910,I230097,I281907);
nand I_13385 (I230470,I281898,I281895);
nor I_13386 (I230487,I230470,I281913);
not I_13387 (I230504,I230487);
nor I_13388 (I230521,I230504,I230182);
DFFARX1 I_13389 (I230521,I2898,I229927,I229913,);
nor I_13390 (I230552,I230487,I230046);
nor I_13391 (I229916,I230470,I230216);
nor I_13392 (I230583,I229987,I230470);
nand I_13393 (I229907,I230583,I281913);
not I_13394 (I230614,I230470);
nand I_13395 (I229904,I230552,I230614);
not I_13396 (I230678,I2905);
or I_13397 (I230695,I49614,I49590);
nor I_13398 (I230712,I49614,I49590);
nor I_13399 (I230729,I230712,I49602);
not I_13400 (I230746,I230729);
nand I_13401 (I230763,I230695,I49599);
not I_13402 (I230780,I230763);
not I_13403 (I230797,I49596);
nor I_13404 (I230640,I230797,I230780);
nor I_13405 (I230828,I230797,I230763);
nor I_13406 (I230845,I230729,I49596);
not I_13407 (I230862,I49605);
nand I_13408 (I230879,I49623,I49590);
nand I_13409 (I230896,I230879,I49605);
nor I_13410 (I230913,I230763,I230896);
not I_13411 (I230930,I230913);
nor I_13412 (I230655,I230896,I230828);
not I_13413 (I230961,I230896);
nor I_13414 (I230978,I230961,I230729);
nor I_13415 (I230643,I230797,I230978);
nor I_13416 (I230658,I230896,I230746);
nand I_13417 (I231023,I230879,I230862);
and I_13418 (I231040,I231023,I49626);
nand I_13419 (I231057,I231040,I49617);
not I_13420 (I231074,I231057);
nor I_13421 (I231091,I231074,I49596);
nand I_13422 (I231108,I230845,I231057);
not I_13423 (I230649,I231108);
nor I_13424 (I231139,I49593,I49608);
or I_13425 (I231156,I231139,I49593);
nor I_13426 (I231173,I49611,I49620);
nand I_13427 (I231190,I231173,I231156);
not I_13428 (I231207,I231190);
nor I_13429 (I230670,I231207,I230763);
nand I_13430 (I231238,I231207,I231091);
nand I_13431 (I230646,I231108,I231238);
nor I_13432 (I231269,I231207,I230780);
nor I_13433 (I230667,I231269,I230797);
nor I_13434 (I230661,I231207,I230961);
nor I_13435 (I231314,I231190,I230746);
nor I_13436 (I231331,I231074,I231314);
nor I_13437 (I230652,I231331,I230930);
nor I_13438 (I231362,I230763,I231190);
nor I_13439 (I231379,I231057,I231362);
DFFARX1 I_13440 (I231379,I2898,I230678,I230664,);
not I_13441 (I231443,I2905);
or I_13442 (I231460,I153160,I153175);
nor I_13443 (I231477,I153160,I153175);
nor I_13444 (I231494,I231477,I153166);
not I_13445 (I231511,I231494);
nand I_13446 (I231528,I231460,I153169);
not I_13447 (I231545,I231528);
not I_13448 (I231562,I153154);
nor I_13449 (I231405,I231562,I231545);
nor I_13450 (I231593,I231562,I231528);
nor I_13451 (I231610,I231494,I153154);
not I_13452 (I231627,I153178);
nand I_13453 (I231644,I153157,I153163);
nand I_13454 (I231661,I231644,I153178);
nor I_13455 (I231678,I231528,I231661);
not I_13456 (I231695,I231678);
nor I_13457 (I231420,I231661,I231593);
not I_13458 (I231726,I231661);
nor I_13459 (I231743,I231726,I231494);
nor I_13460 (I231408,I231562,I231743);
nor I_13461 (I231423,I231661,I231511);
nand I_13462 (I231788,I231644,I231627);
and I_13463 (I231805,I231788,I153184);
nand I_13464 (I231822,I231805,I153160);
not I_13465 (I231839,I231822);
nor I_13466 (I231856,I231839,I153154);
nand I_13467 (I231873,I231610,I231822);
not I_13468 (I231414,I231873);
nor I_13469 (I231904,I153187,I153172);
or I_13470 (I231921,I231904,I153157);
nor I_13471 (I231938,I153154,I153181);
nand I_13472 (I231955,I231938,I231921);
not I_13473 (I231972,I231955);
nor I_13474 (I231435,I231972,I231528);
nand I_13475 (I232003,I231972,I231856);
nand I_13476 (I231411,I231873,I232003);
nor I_13477 (I232034,I231972,I231545);
nor I_13478 (I231432,I232034,I231562);
nor I_13479 (I231426,I231972,I231726);
nor I_13480 (I232079,I231955,I231511);
nor I_13481 (I232096,I231839,I232079);
nor I_13482 (I231417,I232096,I231695);
nor I_13483 (I232127,I231528,I231955);
nor I_13484 (I232144,I231822,I232127);
DFFARX1 I_13485 (I232144,I2898,I231443,I231429,);
not I_13486 (I232208,I2905);
or I_13487 (I232225,I326404,I326401);
nor I_13488 (I232242,I326404,I326401);
nor I_13489 (I232259,I232242,I326410);
not I_13490 (I232276,I232259);
nand I_13491 (I232293,I232225,I326422);
not I_13492 (I232310,I232293);
not I_13493 (I232327,I326419);
nor I_13494 (I232170,I232327,I232310);
nor I_13495 (I232358,I232327,I232293);
nor I_13496 (I232375,I232259,I326419);
not I_13497 (I232392,I326425);
nand I_13498 (I232409,I326404,I326413);
nand I_13499 (I232426,I232409,I326425);
nor I_13500 (I232443,I232293,I232426);
not I_13501 (I232460,I232443);
nor I_13502 (I232185,I232426,I232358);
not I_13503 (I232491,I232426);
nor I_13504 (I232508,I232491,I232259);
nor I_13505 (I232173,I232327,I232508);
nor I_13506 (I232188,I232426,I232276);
nand I_13507 (I232553,I232409,I232392);
and I_13508 (I232570,I232553,I326410);
nand I_13509 (I232587,I232570,I326407);
not I_13510 (I232604,I232587);
nor I_13511 (I232621,I232604,I326419);
nand I_13512 (I232638,I232375,I232587);
not I_13513 (I232179,I232638);
nor I_13514 (I232669,I326416,I326401);
or I_13515 (I232686,I232669,I326413);
nor I_13516 (I232703,I326407,I326416);
nand I_13517 (I232720,I232703,I232686);
not I_13518 (I232737,I232720);
nor I_13519 (I232200,I232737,I232293);
nand I_13520 (I232768,I232737,I232621);
nand I_13521 (I232176,I232638,I232768);
nor I_13522 (I232799,I232737,I232310);
nor I_13523 (I232197,I232799,I232327);
nor I_13524 (I232191,I232737,I232491);
nor I_13525 (I232844,I232720,I232276);
nor I_13526 (I232861,I232604,I232844);
nor I_13527 (I232182,I232861,I232460);
nor I_13528 (I232892,I232293,I232720);
nor I_13529 (I232909,I232587,I232892);
DFFARX1 I_13530 (I232909,I2898,I232208,I232194,);
not I_13531 (I232973,I2905);
or I_13532 (I232990,I109114,I109111);
nor I_13533 (I233007,I109114,I109111);
nor I_13534 (I233024,I233007,I109096);
not I_13535 (I233041,I233024);
nand I_13536 (I233058,I232990,I109117);
not I_13537 (I233075,I233058);
not I_13538 (I233092,I109099);
nor I_13539 (I232935,I233092,I233075);
nor I_13540 (I233123,I233092,I233058);
nor I_13541 (I233140,I233024,I109099);
not I_13542 (I233157,I109093);
nand I_13543 (I233174,I109102,I109090);
nand I_13544 (I233191,I233174,I109093);
nor I_13545 (I233208,I233058,I233191);
not I_13546 (I233225,I233208);
nor I_13547 (I232950,I233191,I233123);
not I_13548 (I233256,I233191);
nor I_13549 (I233273,I233256,I233024);
nor I_13550 (I232938,I233092,I233273);
nor I_13551 (I232953,I233191,I233041);
nand I_13552 (I233318,I233174,I233157);
and I_13553 (I233335,I233318,I109123);
nand I_13554 (I233352,I233335,I109120);
not I_13555 (I233369,I233352);
nor I_13556 (I233386,I233369,I109099);
nand I_13557 (I233403,I233140,I233352);
not I_13558 (I232944,I233403);
nor I_13559 (I233434,I109090,I109108);
or I_13560 (I233451,I233434,I109093);
nor I_13561 (I233468,I109105,I109096);
nand I_13562 (I233485,I233468,I233451);
not I_13563 (I233502,I233485);
nor I_13564 (I232965,I233502,I233058);
nand I_13565 (I233533,I233502,I233386);
nand I_13566 (I232941,I233403,I233533);
nor I_13567 (I233564,I233502,I233075);
nor I_13568 (I232962,I233564,I233092);
nor I_13569 (I232956,I233502,I233256);
nor I_13570 (I233609,I233485,I233041);
nor I_13571 (I233626,I233369,I233609);
nor I_13572 (I232947,I233626,I233225);
nor I_13573 (I233657,I233058,I233485);
nor I_13574 (I233674,I233352,I233657);
DFFARX1 I_13575 (I233674,I2898,I232973,I232959,);
not I_13576 (I233738,I2905);
or I_13577 (I233755,I437333,I437330);
nor I_13578 (I233772,I437333,I437330);
nor I_13579 (I233789,I233772,I437318);
not I_13580 (I233806,I233789);
nand I_13581 (I233823,I233755,I437339);
not I_13582 (I233840,I233823);
not I_13583 (I233857,I437309);
nor I_13584 (I233700,I233857,I233840);
nor I_13585 (I233888,I233857,I233823);
nor I_13586 (I233905,I233789,I437309);
not I_13587 (I233922,I437327);
nand I_13588 (I233939,I437342,I437324);
nand I_13589 (I233956,I233939,I437327);
nor I_13590 (I233973,I233823,I233956);
not I_13591 (I233990,I233973);
nor I_13592 (I233715,I233956,I233888);
not I_13593 (I234021,I233956);
nor I_13594 (I234038,I234021,I233789);
nor I_13595 (I233703,I233857,I234038);
nor I_13596 (I233718,I233956,I233806);
nand I_13597 (I234083,I233939,I233922);
and I_13598 (I234100,I234083,I437336);
nand I_13599 (I234117,I234100,I437315);
not I_13600 (I234134,I234117);
nor I_13601 (I234151,I234134,I437309);
nand I_13602 (I234168,I233905,I234117);
not I_13603 (I233709,I234168);
nor I_13604 (I234199,I437321,I437309);
or I_13605 (I234216,I234199,I437312);
nor I_13606 (I234233,I437312,I437315);
nand I_13607 (I234250,I234233,I234216);
not I_13608 (I234267,I234250);
nor I_13609 (I233730,I234267,I233823);
nand I_13610 (I234298,I234267,I234151);
nand I_13611 (I233706,I234168,I234298);
nor I_13612 (I234329,I234267,I233840);
nor I_13613 (I233727,I234329,I233857);
nor I_13614 (I233721,I234267,I234021);
nor I_13615 (I234374,I234250,I233806);
nor I_13616 (I234391,I234134,I234374);
nor I_13617 (I233712,I234391,I233990);
nor I_13618 (I234422,I233823,I234250);
nor I_13619 (I234439,I234117,I234422);
DFFARX1 I_13620 (I234439,I2898,I233738,I233724,);
not I_13621 (I234503,I2905);
or I_13622 (I234520,I228408,I228402);
nor I_13623 (I234537,I228408,I228402);
nor I_13624 (I234554,I234537,I228417);
not I_13625 (I234571,I234554);
nand I_13626 (I234588,I234520,I228420);
not I_13627 (I234605,I234588);
not I_13628 (I234622,I228402);
nor I_13629 (I234465,I234622,I234605);
nor I_13630 (I234653,I234622,I234588);
nor I_13631 (I234670,I234554,I228402);
not I_13632 (I234687,I228405);
nand I_13633 (I234704,I228423,I228396);
nand I_13634 (I234721,I234704,I228405);
nor I_13635 (I234738,I234588,I234721);
not I_13636 (I234755,I234738);
nor I_13637 (I234480,I234721,I234653);
not I_13638 (I234786,I234721);
nor I_13639 (I234803,I234786,I234554);
nor I_13640 (I234468,I234622,I234803);
nor I_13641 (I234483,I234721,I234571);
nand I_13642 (I234848,I234704,I234687);
and I_13643 (I234865,I234848,I228408);
nand I_13644 (I234882,I234865,I228399);
not I_13645 (I234899,I234882);
nor I_13646 (I234916,I234899,I228402);
nand I_13647 (I234933,I234670,I234882);
not I_13648 (I234474,I234933);
nor I_13649 (I234964,I228399,I228405);
or I_13650 (I234981,I234964,I228396);
nor I_13651 (I234998,I228411,I228414);
nand I_13652 (I235015,I234998,I234981);
not I_13653 (I235032,I235015);
nor I_13654 (I234495,I235032,I234588);
nand I_13655 (I235063,I235032,I234916);
nand I_13656 (I234471,I234933,I235063);
nor I_13657 (I235094,I235032,I234605);
nor I_13658 (I234492,I235094,I234622);
nor I_13659 (I234486,I235032,I234786);
nor I_13660 (I235139,I235015,I234571);
nor I_13661 (I235156,I234899,I235139);
nor I_13662 (I234477,I235156,I234755);
nor I_13663 (I235187,I234588,I235015);
nor I_13664 (I235204,I234882,I235187);
DFFARX1 I_13665 (I235204,I2898,I234503,I234489,);
not I_13666 (I235268,I2905);
or I_13667 (I235285,I361509,I361506);
nor I_13668 (I235302,I361509,I361506);
nor I_13669 (I235319,I235302,I361515);
not I_13670 (I235336,I235319);
nand I_13671 (I235353,I235285,I361527);
not I_13672 (I235370,I235353);
not I_13673 (I235387,I361524);
nor I_13674 (I235230,I235387,I235370);
nor I_13675 (I235418,I235387,I235353);
nor I_13676 (I235435,I235319,I361524);
not I_13677 (I235452,I361530);
nand I_13678 (I235469,I361509,I361518);
nand I_13679 (I235486,I235469,I361530);
nor I_13680 (I235503,I235353,I235486);
not I_13681 (I235520,I235503);
nor I_13682 (I235245,I235486,I235418);
not I_13683 (I235551,I235486);
nor I_13684 (I235568,I235551,I235319);
nor I_13685 (I235233,I235387,I235568);
nor I_13686 (I235248,I235486,I235336);
nand I_13687 (I235613,I235469,I235452);
and I_13688 (I235630,I235613,I361515);
nand I_13689 (I235647,I235630,I361512);
not I_13690 (I235664,I235647);
nor I_13691 (I235681,I235664,I361524);
nand I_13692 (I235698,I235435,I235647);
not I_13693 (I235239,I235698);
nor I_13694 (I235729,I361521,I361506);
or I_13695 (I235746,I235729,I361518);
nor I_13696 (I235763,I361512,I361521);
nand I_13697 (I235780,I235763,I235746);
not I_13698 (I235797,I235780);
nor I_13699 (I235260,I235797,I235353);
nand I_13700 (I235828,I235797,I235681);
nand I_13701 (I235236,I235698,I235828);
nor I_13702 (I235859,I235797,I235370);
nor I_13703 (I235257,I235859,I235387);
nor I_13704 (I235251,I235797,I235551);
nor I_13705 (I235904,I235780,I235336);
nor I_13706 (I235921,I235664,I235904);
nor I_13707 (I235242,I235921,I235520);
nor I_13708 (I235952,I235353,I235780);
nor I_13709 (I235969,I235647,I235952);
DFFARX1 I_13710 (I235969,I2898,I235268,I235254,);
not I_13711 (I236033,I2905);
or I_13712 (I236050,I148400,I148415);
nor I_13713 (I236067,I148400,I148415);
nor I_13714 (I236084,I236067,I148406);
not I_13715 (I236101,I236084);
nand I_13716 (I236118,I236050,I148409);
not I_13717 (I236135,I236118);
not I_13718 (I236152,I148394);
nor I_13719 (I235995,I236152,I236135);
nor I_13720 (I236183,I236152,I236118);
nor I_13721 (I236200,I236084,I148394);
not I_13722 (I236217,I148418);
nand I_13723 (I236234,I148397,I148403);
nand I_13724 (I236251,I236234,I148418);
nor I_13725 (I236268,I236118,I236251);
not I_13726 (I236285,I236268);
nor I_13727 (I236010,I236251,I236183);
not I_13728 (I236316,I236251);
nor I_13729 (I236333,I236316,I236084);
nor I_13730 (I235998,I236152,I236333);
nor I_13731 (I236013,I236251,I236101);
nand I_13732 (I236378,I236234,I236217);
and I_13733 (I236395,I236378,I148424);
nand I_13734 (I236412,I236395,I148400);
not I_13735 (I236429,I236412);
nor I_13736 (I236446,I236429,I148394);
nand I_13737 (I236463,I236200,I236412);
not I_13738 (I236004,I236463);
nor I_13739 (I236494,I148427,I148412);
or I_13740 (I236511,I236494,I148397);
nor I_13741 (I236528,I148394,I148421);
nand I_13742 (I236545,I236528,I236511);
not I_13743 (I236562,I236545);
nor I_13744 (I236025,I236562,I236118);
nand I_13745 (I236593,I236562,I236446);
nand I_13746 (I236001,I236463,I236593);
nor I_13747 (I236624,I236562,I236135);
nor I_13748 (I236022,I236624,I236152);
nor I_13749 (I236016,I236562,I236316);
nor I_13750 (I236669,I236545,I236101);
nor I_13751 (I236686,I236429,I236669);
nor I_13752 (I236007,I236686,I236285);
nor I_13753 (I236717,I236118,I236545);
nor I_13754 (I236734,I236412,I236717);
DFFARX1 I_13755 (I236734,I2898,I236033,I236019,);
not I_13756 (I236798,I2905);
or I_13757 (I236815,I335329,I335326);
nor I_13758 (I236832,I335329,I335326);
nor I_13759 (I236849,I236832,I335335);
not I_13760 (I236866,I236849);
nand I_13761 (I236883,I236815,I335347);
not I_13762 (I236900,I236883);
not I_13763 (I236917,I335344);
nor I_13764 (I236760,I236917,I236900);
nor I_13765 (I236948,I236917,I236883);
nor I_13766 (I236965,I236849,I335344);
not I_13767 (I236982,I335350);
nand I_13768 (I236999,I335329,I335338);
nand I_13769 (I237016,I236999,I335350);
nor I_13770 (I237033,I236883,I237016);
not I_13771 (I237050,I237033);
nor I_13772 (I236775,I237016,I236948);
not I_13773 (I237081,I237016);
nor I_13774 (I237098,I237081,I236849);
nor I_13775 (I236763,I236917,I237098);
nor I_13776 (I236778,I237016,I236866);
nand I_13777 (I237143,I236999,I236982);
and I_13778 (I237160,I237143,I335335);
nand I_13779 (I237177,I237160,I335332);
not I_13780 (I237194,I237177);
nor I_13781 (I237211,I237194,I335344);
nand I_13782 (I237228,I236965,I237177);
not I_13783 (I236769,I237228);
nor I_13784 (I237259,I335341,I335326);
or I_13785 (I237276,I237259,I335338);
nor I_13786 (I237293,I335332,I335341);
nand I_13787 (I237310,I237293,I237276);
not I_13788 (I237327,I237310);
nor I_13789 (I236790,I237327,I236883);
nand I_13790 (I237358,I237327,I237211);
nand I_13791 (I236766,I237228,I237358);
nor I_13792 (I237389,I237327,I236900);
nor I_13793 (I236787,I237389,I236917);
nor I_13794 (I236781,I237327,I237081);
nor I_13795 (I237434,I237310,I236866);
nor I_13796 (I237451,I237194,I237434);
nor I_13797 (I236772,I237451,I237050);
nor I_13798 (I237482,I236883,I237310);
nor I_13799 (I237499,I237177,I237482);
DFFARX1 I_13800 (I237499,I2898,I236798,I236784,);
not I_13801 (I237563,I2905);
or I_13802 (I237580,I142451,I142448);
nor I_13803 (I237597,I142451,I142448);
nor I_13804 (I237614,I237597,I142433);
not I_13805 (I237631,I237614);
nand I_13806 (I237648,I237580,I142454);
not I_13807 (I237665,I237648);
not I_13808 (I237682,I142436);
nor I_13809 (I237525,I237682,I237665);
nor I_13810 (I237713,I237682,I237648);
nor I_13811 (I237730,I237614,I142436);
not I_13812 (I237747,I142430);
nand I_13813 (I237764,I142439,I142427);
nand I_13814 (I237781,I237764,I142430);
nor I_13815 (I237798,I237648,I237781);
not I_13816 (I237815,I237798);
nor I_13817 (I237540,I237781,I237713);
not I_13818 (I237846,I237781);
nor I_13819 (I237863,I237846,I237614);
nor I_13820 (I237528,I237682,I237863);
nor I_13821 (I237543,I237781,I237631);
nand I_13822 (I237908,I237764,I237747);
and I_13823 (I237925,I237908,I142460);
nand I_13824 (I237942,I237925,I142457);
not I_13825 (I237959,I237942);
nor I_13826 (I237976,I237959,I142436);
nand I_13827 (I237993,I237730,I237942);
not I_13828 (I237534,I237993);
nor I_13829 (I238024,I142427,I142445);
or I_13830 (I238041,I238024,I142430);
nor I_13831 (I238058,I142442,I142433);
nand I_13832 (I238075,I238058,I238041);
not I_13833 (I238092,I238075);
nor I_13834 (I237555,I238092,I237648);
nand I_13835 (I238123,I238092,I237976);
nand I_13836 (I237531,I237993,I238123);
nor I_13837 (I238154,I238092,I237665);
nor I_13838 (I237552,I238154,I237682);
nor I_13839 (I237546,I238092,I237846);
nor I_13840 (I238199,I238075,I237631);
nor I_13841 (I238216,I237959,I238199);
nor I_13842 (I237537,I238216,I237815);
nor I_13843 (I238247,I237648,I238075);
nor I_13844 (I238264,I237942,I238247);
DFFARX1 I_13845 (I238264,I2898,I237563,I237549,);
not I_13846 (I238328,I2905);
or I_13847 (I238345,I395872,I395884);
nor I_13848 (I238362,I395872,I395884);
nor I_13849 (I238379,I238362,I395866);
not I_13850 (I238396,I238379);
nand I_13851 (I238413,I238345,I395878);
not I_13852 (I238430,I238413);
not I_13853 (I238447,I395872);
nor I_13854 (I238290,I238447,I238430);
nor I_13855 (I238478,I238447,I238413);
nor I_13856 (I238495,I238379,I395872);
not I_13857 (I238512,I395863);
nand I_13858 (I238529,I395881,I395875);
nand I_13859 (I238546,I238529,I395863);
nor I_13860 (I238563,I238413,I238546);
not I_13861 (I238580,I238563);
nor I_13862 (I238305,I238546,I238478);
not I_13863 (I238611,I238546);
nor I_13864 (I238628,I238611,I238379);
nor I_13865 (I238293,I238447,I238628);
nor I_13866 (I238308,I238546,I238396);
nand I_13867 (I238673,I238529,I238512);
and I_13868 (I238690,I238673,I395887);
nand I_13869 (I238707,I238690,I395878);
not I_13870 (I238724,I238707);
nor I_13871 (I238741,I238724,I395872);
nand I_13872 (I238758,I238495,I238707);
not I_13873 (I238299,I238758);
nor I_13874 (I238789,I395875,I395866);
or I_13875 (I238806,I238789,I395863);
nor I_13876 (I238823,I395869,I395869);
nand I_13877 (I238840,I238823,I238806);
not I_13878 (I238857,I238840);
nor I_13879 (I238320,I238857,I238413);
nand I_13880 (I238888,I238857,I238741);
nand I_13881 (I238296,I238758,I238888);
nor I_13882 (I238919,I238857,I238430);
nor I_13883 (I238317,I238919,I238447);
nor I_13884 (I238311,I238857,I238611);
nor I_13885 (I238964,I238840,I238396);
nor I_13886 (I238981,I238724,I238964);
nor I_13887 (I238302,I238981,I238580);
nor I_13888 (I239012,I238413,I238840);
nor I_13889 (I239029,I238707,I239012);
DFFARX1 I_13890 (I239029,I2898,I238328,I238314,);
not I_13891 (I239093,I2905);
or I_13892 (I239110,I367289,I367304);
nor I_13893 (I239127,I367289,I367304);
nor I_13894 (I239144,I239127,I367313);
not I_13895 (I239161,I239144);
nand I_13896 (I239178,I239110,I367301);
not I_13897 (I239195,I239178);
not I_13898 (I239212,I367298);
nor I_13899 (I239055,I239212,I239195);
nor I_13900 (I239243,I239212,I239178);
nor I_13901 (I239260,I239144,I367298);
not I_13902 (I239277,I367292);
nand I_13903 (I239294,I367289,I367310);
nand I_13904 (I239311,I239294,I367292);
nor I_13905 (I239328,I239178,I239311);
not I_13906 (I239345,I239328);
nor I_13907 (I239070,I239311,I239243);
not I_13908 (I239376,I239311);
nor I_13909 (I239393,I239376,I239144);
nor I_13910 (I239058,I239212,I239393);
nor I_13911 (I239073,I239311,I239161);
nand I_13912 (I239438,I239294,I239277);
and I_13913 (I239455,I239438,I367316);
nand I_13914 (I239472,I239455,I367319);
not I_13915 (I239489,I239472);
nor I_13916 (I239506,I239489,I367298);
nand I_13917 (I239523,I239260,I239472);
not I_13918 (I239064,I239523);
nor I_13919 (I239554,I367292,I367286);
or I_13920 (I239571,I239554,I367286);
nor I_13921 (I239588,I367295,I367307);
nand I_13922 (I239605,I239588,I239571);
not I_13923 (I239622,I239605);
nor I_13924 (I239085,I239622,I239178);
nand I_13925 (I239653,I239622,I239506);
nand I_13926 (I239061,I239523,I239653);
nor I_13927 (I239684,I239622,I239195);
nor I_13928 (I239082,I239684,I239212);
nor I_13929 (I239076,I239622,I239376);
nor I_13930 (I239729,I239605,I239161);
nor I_13931 (I239746,I239489,I239729);
nor I_13932 (I239067,I239746,I239345);
nor I_13933 (I239777,I239178,I239605);
nor I_13934 (I239794,I239472,I239777);
DFFARX1 I_13935 (I239794,I2898,I239093,I239079,);
not I_13936 (I239858,I2905);
or I_13937 (I239875,I111001,I110998);
nor I_13938 (I239892,I111001,I110998);
nor I_13939 (I239909,I239892,I110983);
not I_13940 (I239926,I239909);
nand I_13941 (I239943,I239875,I111004);
not I_13942 (I239960,I239943);
not I_13943 (I239977,I110986);
nor I_13944 (I239820,I239977,I239960);
nor I_13945 (I240008,I239977,I239943);
nor I_13946 (I240025,I239909,I110986);
not I_13947 (I240042,I110980);
nand I_13948 (I240059,I110989,I110977);
nand I_13949 (I240076,I240059,I110980);
nor I_13950 (I240093,I239943,I240076);
not I_13951 (I240110,I240093);
nor I_13952 (I239835,I240076,I240008);
not I_13953 (I240141,I240076);
nor I_13954 (I240158,I240141,I239909);
nor I_13955 (I239823,I239977,I240158);
nor I_13956 (I239838,I240076,I239926);
nand I_13957 (I240203,I240059,I240042);
and I_13958 (I240220,I240203,I111010);
nand I_13959 (I240237,I240220,I111007);
not I_13960 (I240254,I240237);
nor I_13961 (I240271,I240254,I110986);
nand I_13962 (I240288,I240025,I240237);
not I_13963 (I239829,I240288);
nor I_13964 (I240319,I110977,I110995);
or I_13965 (I240336,I240319,I110980);
nor I_13966 (I240353,I110992,I110983);
nand I_13967 (I240370,I240353,I240336);
not I_13968 (I240387,I240370);
nor I_13969 (I239850,I240387,I239943);
nand I_13970 (I240418,I240387,I240271);
nand I_13971 (I239826,I240288,I240418);
nor I_13972 (I240449,I240387,I239960);
nor I_13973 (I239847,I240449,I239977);
nor I_13974 (I239841,I240387,I240141);
nor I_13975 (I240494,I240370,I239926);
nor I_13976 (I240511,I240254,I240494);
nor I_13977 (I239832,I240511,I240110);
nor I_13978 (I240542,I239943,I240370);
nor I_13979 (I240559,I240237,I240542);
DFFARX1 I_13980 (I240559,I2898,I239858,I239844,);
not I_13981 (I240623,I2905);
or I_13982 (I240640,I77074,I77086);
nor I_13983 (I240657,I77074,I77086);
nor I_13984 (I240674,I240657,I77083);
not I_13985 (I240691,I240674);
nand I_13986 (I240708,I240640,I77077);
not I_13987 (I240725,I240708);
not I_13988 (I240742,I77071);
nor I_13989 (I240585,I240742,I240725);
nor I_13990 (I240773,I240742,I240708);
nor I_13991 (I240790,I240674,I77071);
not I_13992 (I240807,I77080);
nand I_13993 (I240824,I77068,I77065);
nand I_13994 (I240841,I240824,I77080);
nor I_13995 (I240858,I240708,I240841);
not I_13996 (I240875,I240858);
nor I_13997 (I240600,I240841,I240773);
not I_13998 (I240906,I240841);
nor I_13999 (I240923,I240906,I240674);
nor I_14000 (I240588,I240742,I240923);
nor I_14001 (I240603,I240841,I240691);
nand I_14002 (I240968,I240824,I240807);
and I_14003 (I240985,I240968,I77074);
nand I_14004 (I241002,I240985,I77062);
not I_14005 (I241019,I241002);
nor I_14006 (I241036,I241019,I77071);
nand I_14007 (I241053,I240790,I241002);
not I_14008 (I240594,I241053);
nor I_14009 (I241084,I77068,I77065);
or I_14010 (I241101,I241084,I77071);
nor I_14011 (I241118,I77062,I77089);
nand I_14012 (I241135,I241118,I241101);
not I_14013 (I241152,I241135);
nor I_14014 (I240615,I241152,I240708);
nand I_14015 (I241183,I241152,I241036);
nand I_14016 (I240591,I241053,I241183);
nor I_14017 (I241214,I241152,I240725);
nor I_14018 (I240612,I241214,I240742);
nor I_14019 (I240606,I241152,I240906);
nor I_14020 (I241259,I241135,I240691);
nor I_14021 (I241276,I241019,I241259);
nor I_14022 (I240597,I241276,I240875);
nor I_14023 (I241307,I240708,I241135);
nor I_14024 (I241324,I241002,I241307);
DFFARX1 I_14025 (I241324,I2898,I240623,I240609,);
not I_14026 (I241388,I2905);
or I_14027 (I241405,I346634,I346631);
nor I_14028 (I241422,I346634,I346631);
nor I_14029 (I241439,I241422,I346640);
not I_14030 (I241456,I241439);
nand I_14031 (I241473,I241405,I346652);
not I_14032 (I241490,I241473);
not I_14033 (I241507,I346649);
nor I_14034 (I241350,I241507,I241490);
nor I_14035 (I241538,I241507,I241473);
nor I_14036 (I241555,I241439,I346649);
not I_14037 (I241572,I346655);
nand I_14038 (I241589,I346634,I346643);
nand I_14039 (I241606,I241589,I346655);
nor I_14040 (I241623,I241473,I241606);
not I_14041 (I241640,I241623);
nor I_14042 (I241365,I241606,I241538);
not I_14043 (I241671,I241606);
nor I_14044 (I241688,I241671,I241439);
nor I_14045 (I241353,I241507,I241688);
nor I_14046 (I241368,I241606,I241456);
nand I_14047 (I241733,I241589,I241572);
and I_14048 (I241750,I241733,I346640);
nand I_14049 (I241767,I241750,I346637);
not I_14050 (I241784,I241767);
nor I_14051 (I241801,I241784,I346649);
nand I_14052 (I241818,I241555,I241767);
not I_14053 (I241359,I241818);
nor I_14054 (I241849,I346646,I346631);
or I_14055 (I241866,I241849,I346643);
nor I_14056 (I241883,I346637,I346646);
nand I_14057 (I241900,I241883,I241866);
not I_14058 (I241917,I241900);
nor I_14059 (I241380,I241917,I241473);
nand I_14060 (I241948,I241917,I241801);
nand I_14061 (I241356,I241818,I241948);
nor I_14062 (I241979,I241917,I241490);
nor I_14063 (I241377,I241979,I241507);
nor I_14064 (I241371,I241917,I241671);
nor I_14065 (I242024,I241900,I241456);
nor I_14066 (I242041,I241784,I242024);
nor I_14067 (I241362,I242041,I241640);
nor I_14068 (I242072,I241473,I241900);
nor I_14069 (I242089,I241767,I242072);
DFFARX1 I_14070 (I242089,I2898,I241388,I241374,);
not I_14071 (I242153,I2905);
or I_14072 (I242170,I58204,I58216);
nor I_14073 (I242187,I58204,I58216);
nor I_14074 (I242204,I242187,I58213);
not I_14075 (I242221,I242204);
nand I_14076 (I242238,I242170,I58207);
not I_14077 (I242255,I242238);
not I_14078 (I242272,I58201);
nor I_14079 (I242115,I242272,I242255);
nor I_14080 (I242303,I242272,I242238);
nor I_14081 (I242320,I242204,I58201);
not I_14082 (I242337,I58210);
nand I_14083 (I242354,I58198,I58195);
nand I_14084 (I242371,I242354,I58210);
nor I_14085 (I242388,I242238,I242371);
not I_14086 (I242405,I242388);
nor I_14087 (I242130,I242371,I242303);
not I_14088 (I242436,I242371);
nor I_14089 (I242453,I242436,I242204);
nor I_14090 (I242118,I242272,I242453);
nor I_14091 (I242133,I242371,I242221);
nand I_14092 (I242498,I242354,I242337);
and I_14093 (I242515,I242498,I58204);
nand I_14094 (I242532,I242515,I58192);
not I_14095 (I242549,I242532);
nor I_14096 (I242566,I242549,I58201);
nand I_14097 (I242583,I242320,I242532);
not I_14098 (I242124,I242583);
nor I_14099 (I242614,I58198,I58195);
or I_14100 (I242631,I242614,I58201);
nor I_14101 (I242648,I58192,I58219);
nand I_14102 (I242665,I242648,I242631);
not I_14103 (I242682,I242665);
nor I_14104 (I242145,I242682,I242238);
nand I_14105 (I242713,I242682,I242566);
nand I_14106 (I242121,I242583,I242713);
nor I_14107 (I242744,I242682,I242255);
nor I_14108 (I242142,I242744,I242272);
nor I_14109 (I242136,I242682,I242436);
nor I_14110 (I242789,I242665,I242221);
nor I_14111 (I242806,I242549,I242789);
nor I_14112 (I242127,I242806,I242405);
nor I_14113 (I242837,I242238,I242665);
nor I_14114 (I242854,I242532,I242837);
DFFARX1 I_14115 (I242854,I2898,I242153,I242139,);
not I_14116 (I242918,I2905);
or I_14117 (I242935,I133645,I133642);
nor I_14118 (I242952,I133645,I133642);
nor I_14119 (I242969,I242952,I133627);
not I_14120 (I242986,I242969);
nand I_14121 (I243003,I242935,I133648);
not I_14122 (I243020,I243003);
not I_14123 (I243037,I133630);
nor I_14124 (I242880,I243037,I243020);
nor I_14125 (I243068,I243037,I243003);
nor I_14126 (I243085,I242969,I133630);
not I_14127 (I243102,I133624);
nand I_14128 (I243119,I133633,I133621);
nand I_14129 (I243136,I243119,I133624);
nor I_14130 (I243153,I243003,I243136);
not I_14131 (I243170,I243153);
nor I_14132 (I242895,I243136,I243068);
not I_14133 (I243201,I243136);
nor I_14134 (I243218,I243201,I242969);
nor I_14135 (I242883,I243037,I243218);
nor I_14136 (I242898,I243136,I242986);
nand I_14137 (I243263,I243119,I243102);
and I_14138 (I243280,I243263,I133654);
nand I_14139 (I243297,I243280,I133651);
not I_14140 (I243314,I243297);
nor I_14141 (I243331,I243314,I133630);
nand I_14142 (I243348,I243085,I243297);
not I_14143 (I242889,I243348);
nor I_14144 (I243379,I133621,I133639);
or I_14145 (I243396,I243379,I133624);
nor I_14146 (I243413,I133636,I133627);
nand I_14147 (I243430,I243413,I243396);
not I_14148 (I243447,I243430);
nor I_14149 (I242910,I243447,I243003);
nand I_14150 (I243478,I243447,I243331);
nand I_14151 (I242886,I243348,I243478);
nor I_14152 (I243509,I243447,I243020);
nor I_14153 (I242907,I243509,I243037);
nor I_14154 (I242901,I243447,I243201);
nor I_14155 (I243554,I243430,I242986);
nor I_14156 (I243571,I243314,I243554);
nor I_14157 (I242892,I243571,I243170);
nor I_14158 (I243602,I243003,I243430);
nor I_14159 (I243619,I243297,I243602);
DFFARX1 I_14160 (I243619,I2898,I242918,I242904,);
not I_14161 (I243683,I2905);
or I_14162 (I243700,I402672,I402684);
nor I_14163 (I243717,I402672,I402684);
nor I_14164 (I243734,I243717,I402666);
not I_14165 (I243751,I243734);
nand I_14166 (I243768,I243700,I402678);
not I_14167 (I243785,I243768);
not I_14168 (I243802,I402672);
nor I_14169 (I243645,I243802,I243785);
nor I_14170 (I243833,I243802,I243768);
nor I_14171 (I243850,I243734,I402672);
not I_14172 (I243867,I402663);
nand I_14173 (I243884,I402681,I402675);
nand I_14174 (I243901,I243884,I402663);
nor I_14175 (I243918,I243768,I243901);
not I_14176 (I243935,I243918);
nor I_14177 (I243660,I243901,I243833);
not I_14178 (I243966,I243901);
nor I_14179 (I243983,I243966,I243734);
nor I_14180 (I243648,I243802,I243983);
nor I_14181 (I243663,I243901,I243751);
nand I_14182 (I244028,I243884,I243867);
and I_14183 (I244045,I244028,I402687);
nand I_14184 (I244062,I244045,I402678);
not I_14185 (I244079,I244062);
nor I_14186 (I244096,I244079,I402672);
nand I_14187 (I244113,I243850,I244062);
not I_14188 (I243654,I244113);
nor I_14189 (I244144,I402675,I402666);
or I_14190 (I244161,I244144,I402663);
nor I_14191 (I244178,I402669,I402669);
nand I_14192 (I244195,I244178,I244161);
not I_14193 (I244212,I244195);
nor I_14194 (I243675,I244212,I243768);
nand I_14195 (I244243,I244212,I244096);
nand I_14196 (I243651,I244113,I244243);
nor I_14197 (I244274,I244212,I243785);
nor I_14198 (I243672,I244274,I243802);
nor I_14199 (I243666,I244212,I243966);
nor I_14200 (I244319,I244195,I243751);
nor I_14201 (I244336,I244079,I244319);
nor I_14202 (I243657,I244336,I243935);
nor I_14203 (I244367,I243768,I244195);
nor I_14204 (I244384,I244062,I244367);
DFFARX1 I_14205 (I244384,I2898,I243683,I243669,);
not I_14206 (I244448,I2905);
or I_14207 (I244465,I145000,I145015);
nor I_14208 (I244482,I145000,I145015);
nor I_14209 (I244499,I244482,I145006);
not I_14210 (I244516,I244499);
nand I_14211 (I244533,I244465,I145009);
not I_14212 (I244550,I244533);
not I_14213 (I244567,I144994);
nor I_14214 (I244410,I244567,I244550);
nor I_14215 (I244598,I244567,I244533);
nor I_14216 (I244615,I244499,I144994);
not I_14217 (I244632,I145018);
nand I_14218 (I244649,I144997,I145003);
nand I_14219 (I244666,I244649,I145018);
nor I_14220 (I244683,I244533,I244666);
not I_14221 (I244700,I244683);
nor I_14222 (I244425,I244666,I244598);
not I_14223 (I244731,I244666);
nor I_14224 (I244748,I244731,I244499);
nor I_14225 (I244413,I244567,I244748);
nor I_14226 (I244428,I244666,I244516);
nand I_14227 (I244793,I244649,I244632);
and I_14228 (I244810,I244793,I145024);
nand I_14229 (I244827,I244810,I145000);
not I_14230 (I244844,I244827);
nor I_14231 (I244861,I244844,I144994);
nand I_14232 (I244878,I244615,I244827);
not I_14233 (I244419,I244878);
nor I_14234 (I244909,I145027,I145012);
or I_14235 (I244926,I244909,I144997);
nor I_14236 (I244943,I144994,I145021);
nand I_14237 (I244960,I244943,I244926);
not I_14238 (I244977,I244960);
nor I_14239 (I244440,I244977,I244533);
nand I_14240 (I245008,I244977,I244861);
nand I_14241 (I244416,I244878,I245008);
nor I_14242 (I245039,I244977,I244550);
nor I_14243 (I244437,I245039,I244567);
nor I_14244 (I244431,I244977,I244731);
nor I_14245 (I245084,I244960,I244516);
nor I_14246 (I245101,I244844,I245084);
nor I_14247 (I244422,I245101,I244700);
nor I_14248 (I245132,I244533,I244960);
nor I_14249 (I245149,I244827,I245132);
DFFARX1 I_14250 (I245149,I2898,I244448,I244434,);
not I_14251 (I245213,I2905);
or I_14252 (I245230,I149760,I149775);
nor I_14253 (I245247,I149760,I149775);
nor I_14254 (I245264,I245247,I149766);
not I_14255 (I245281,I245264);
nand I_14256 (I245298,I245230,I149769);
not I_14257 (I245315,I245298);
not I_14258 (I245332,I149754);
nor I_14259 (I245175,I245332,I245315);
nor I_14260 (I245363,I245332,I245298);
nor I_14261 (I245380,I245264,I149754);
not I_14262 (I245397,I149778);
nand I_14263 (I245414,I149757,I149763);
nand I_14264 (I245431,I245414,I149778);
nor I_14265 (I245448,I245298,I245431);
not I_14266 (I245465,I245448);
nor I_14267 (I245190,I245431,I245363);
not I_14268 (I245496,I245431);
nor I_14269 (I245513,I245496,I245264);
nor I_14270 (I245178,I245332,I245513);
nor I_14271 (I245193,I245431,I245281);
nand I_14272 (I245558,I245414,I245397);
and I_14273 (I245575,I245558,I149784);
nand I_14274 (I245592,I245575,I149760);
not I_14275 (I245609,I245592);
nor I_14276 (I245626,I245609,I149754);
nand I_14277 (I245643,I245380,I245592);
not I_14278 (I245184,I245643);
nor I_14279 (I245674,I149787,I149772);
or I_14280 (I245691,I245674,I149757);
nor I_14281 (I245708,I149754,I149781);
nand I_14282 (I245725,I245708,I245691);
not I_14283 (I245742,I245725);
nor I_14284 (I245205,I245742,I245298);
nand I_14285 (I245773,I245742,I245626);
nand I_14286 (I245181,I245643,I245773);
nor I_14287 (I245804,I245742,I245315);
nor I_14288 (I245202,I245804,I245332);
nor I_14289 (I245196,I245742,I245496);
nor I_14290 (I245849,I245725,I245281);
nor I_14291 (I245866,I245609,I245849);
nor I_14292 (I245187,I245866,I245465);
nor I_14293 (I245897,I245298,I245725);
nor I_14294 (I245914,I245592,I245897);
DFFARX1 I_14295 (I245914,I2898,I245213,I245199,);
not I_14296 (I245978,I2905);
or I_14297 (I245995,I13945,I13933);
nor I_14298 (I246012,I13945,I13933);
nor I_14299 (I246029,I246012,I13936);
not I_14300 (I246046,I246029);
nand I_14301 (I246063,I245995,I13924);
not I_14302 (I246080,I246063);
not I_14303 (I246097,I13948);
nor I_14304 (I245940,I246097,I246080);
nor I_14305 (I246128,I246097,I246063);
nor I_14306 (I246145,I246029,I13948);
not I_14307 (I246162,I13924);
nand I_14308 (I246179,I13939,I13930);
nand I_14309 (I246196,I246179,I13924);
nor I_14310 (I246213,I246063,I246196);
not I_14311 (I246230,I246213);
nor I_14312 (I245955,I246196,I246128);
not I_14313 (I246261,I246196);
nor I_14314 (I246278,I246261,I246029);
nor I_14315 (I245943,I246097,I246278);
nor I_14316 (I245958,I246196,I246046);
nand I_14317 (I246323,I246179,I246162);
and I_14318 (I246340,I246323,I13936);
nand I_14319 (I246357,I246340,I13927);
not I_14320 (I246374,I246357);
nor I_14321 (I246391,I246374,I13948);
nand I_14322 (I246408,I246145,I246357);
not I_14323 (I245949,I246408);
nor I_14324 (I246439,I13927,I13951);
or I_14325 (I246456,I246439,I13942);
nor I_14326 (I246473,I13933,I13930);
nand I_14327 (I246490,I246473,I246456);
not I_14328 (I246507,I246490);
nor I_14329 (I245970,I246507,I246063);
nand I_14330 (I246538,I246507,I246391);
nand I_14331 (I245946,I246408,I246538);
nor I_14332 (I246569,I246507,I246080);
nor I_14333 (I245967,I246569,I246097);
nor I_14334 (I245961,I246507,I246261);
nor I_14335 (I246614,I246490,I246046);
nor I_14336 (I246631,I246374,I246614);
nor I_14337 (I245952,I246631,I246230);
nor I_14338 (I246662,I246063,I246490);
nor I_14339 (I246679,I246357,I246662);
DFFARX1 I_14340 (I246679,I2898,I245978,I245964,);
not I_14341 (I246743,I2905);
or I_14342 (I246760,I372576,I372579);
nor I_14343 (I246777,I372576,I372579);
nor I_14344 (I246794,I246777,I372573);
not I_14345 (I246811,I246794);
nand I_14346 (I246828,I246760,I372591);
not I_14347 (I246845,I246828);
not I_14348 (I246862,I372600);
nor I_14349 (I246705,I246862,I246845);
nor I_14350 (I246893,I246862,I246828);
nor I_14351 (I246910,I246794,I372600);
not I_14352 (I246927,I372585);
nand I_14353 (I246944,I372573,I372582);
nand I_14354 (I246961,I246944,I372585);
nor I_14355 (I246978,I246828,I246961);
not I_14356 (I246995,I246978);
nor I_14357 (I246720,I246961,I246893);
not I_14358 (I247026,I246961);
nor I_14359 (I247043,I247026,I246794);
nor I_14360 (I246708,I246862,I247043);
nor I_14361 (I246723,I246961,I246811);
nand I_14362 (I247088,I246944,I246927);
and I_14363 (I247105,I247088,I372576);
nand I_14364 (I247122,I247105,I372579);
not I_14365 (I247139,I247122);
nor I_14366 (I247156,I247139,I372600);
nand I_14367 (I247173,I246910,I247122);
not I_14368 (I246714,I247173);
nor I_14369 (I247204,I372603,I372588);
or I_14370 (I247221,I247204,I372597);
nor I_14371 (I247238,I372606,I372594);
nand I_14372 (I247255,I247238,I247221);
not I_14373 (I247272,I247255);
nor I_14374 (I246735,I247272,I246828);
nand I_14375 (I247303,I247272,I247156);
nand I_14376 (I246711,I247173,I247303);
nor I_14377 (I247334,I247272,I246845);
nor I_14378 (I246732,I247334,I246862);
nor I_14379 (I246726,I247272,I247026);
nor I_14380 (I247379,I247255,I246811);
nor I_14381 (I247396,I247139,I247379);
nor I_14382 (I246717,I247396,I246995);
nor I_14383 (I247427,I246828,I247255);
nor I_14384 (I247444,I247122,I247427);
DFFARX1 I_14385 (I247444,I2898,I246743,I246729,);
not I_14386 (I247508,I2905);
or I_14387 (I247525,I94057,I94069);
nor I_14388 (I247542,I94057,I94069);
nor I_14389 (I247559,I247542,I94066);
not I_14390 (I247576,I247559);
nand I_14391 (I247593,I247525,I94060);
not I_14392 (I247610,I247593);
not I_14393 (I247627,I94054);
nor I_14394 (I247470,I247627,I247610);
nor I_14395 (I247658,I247627,I247593);
nor I_14396 (I247675,I247559,I94054);
not I_14397 (I247692,I94063);
nand I_14398 (I247709,I94051,I94048);
nand I_14399 (I247726,I247709,I94063);
nor I_14400 (I247743,I247593,I247726);
not I_14401 (I247760,I247743);
nor I_14402 (I247485,I247726,I247658);
not I_14403 (I247791,I247726);
nor I_14404 (I247808,I247791,I247559);
nor I_14405 (I247473,I247627,I247808);
nor I_14406 (I247488,I247726,I247576);
nand I_14407 (I247853,I247709,I247692);
and I_14408 (I247870,I247853,I94057);
nand I_14409 (I247887,I247870,I94045);
not I_14410 (I247904,I247887);
nor I_14411 (I247921,I247904,I94054);
nand I_14412 (I247938,I247675,I247887);
not I_14413 (I247479,I247938);
nor I_14414 (I247969,I94051,I94048);
or I_14415 (I247986,I247969,I94054);
nor I_14416 (I248003,I94045,I94072);
nand I_14417 (I248020,I248003,I247986);
not I_14418 (I248037,I248020);
nor I_14419 (I247500,I248037,I247593);
nand I_14420 (I248068,I248037,I247921);
nand I_14421 (I247476,I247938,I248068);
nor I_14422 (I248099,I248037,I247610);
nor I_14423 (I247497,I248099,I247627);
nor I_14424 (I247491,I248037,I247791);
nor I_14425 (I248144,I248020,I247576);
nor I_14426 (I248161,I247904,I248144);
nor I_14427 (I247482,I248161,I247760);
nor I_14428 (I248192,I247593,I248020);
nor I_14429 (I248209,I247887,I248192);
DFFARX1 I_14430 (I248209,I2898,I247508,I247494,);
not I_14431 (I248273,I2905);
or I_14432 (I248290,I160640,I160655);
nor I_14433 (I248307,I160640,I160655);
nor I_14434 (I248324,I248307,I160646);
not I_14435 (I248341,I248324);
nand I_14436 (I248358,I248290,I160649);
not I_14437 (I248375,I248358);
not I_14438 (I248392,I160634);
nor I_14439 (I248235,I248392,I248375);
nor I_14440 (I248423,I248392,I248358);
nor I_14441 (I248440,I248324,I160634);
not I_14442 (I248457,I160658);
nand I_14443 (I248474,I160637,I160643);
nand I_14444 (I248491,I248474,I160658);
nor I_14445 (I248508,I248358,I248491);
not I_14446 (I248525,I248508);
nor I_14447 (I248250,I248491,I248423);
not I_14448 (I248556,I248491);
nor I_14449 (I248573,I248556,I248324);
nor I_14450 (I248238,I248392,I248573);
nor I_14451 (I248253,I248491,I248341);
nand I_14452 (I248618,I248474,I248457);
and I_14453 (I248635,I248618,I160664);
nand I_14454 (I248652,I248635,I160640);
not I_14455 (I248669,I248652);
nor I_14456 (I248686,I248669,I160634);
nand I_14457 (I248703,I248440,I248652);
not I_14458 (I248244,I248703);
nor I_14459 (I248734,I160667,I160652);
or I_14460 (I248751,I248734,I160637);
nor I_14461 (I248768,I160634,I160661);
nand I_14462 (I248785,I248768,I248751);
not I_14463 (I248802,I248785);
nor I_14464 (I248265,I248802,I248358);
nand I_14465 (I248833,I248802,I248686);
nand I_14466 (I248241,I248703,I248833);
nor I_14467 (I248864,I248802,I248375);
nor I_14468 (I248262,I248864,I248392);
nor I_14469 (I248256,I248802,I248556);
nor I_14470 (I248909,I248785,I248341);
nor I_14471 (I248926,I248669,I248909);
nor I_14472 (I248247,I248926,I248525);
nor I_14473 (I248957,I248358,I248785);
nor I_14474 (I248974,I248652,I248957);
DFFARX1 I_14475 (I248974,I2898,I248273,I248259,);
not I_14476 (I249038,I2905);
or I_14477 (I249055,I350799,I350796);
nor I_14478 (I249072,I350799,I350796);
nor I_14479 (I249089,I249072,I350805);
not I_14480 (I249106,I249089);
nand I_14481 (I249123,I249055,I350817);
not I_14482 (I249140,I249123);
not I_14483 (I249157,I350814);
nor I_14484 (I249000,I249157,I249140);
nor I_14485 (I249188,I249157,I249123);
nor I_14486 (I249205,I249089,I350814);
not I_14487 (I249222,I350820);
nand I_14488 (I249239,I350799,I350808);
nand I_14489 (I249256,I249239,I350820);
nor I_14490 (I249273,I249123,I249256);
not I_14491 (I249290,I249273);
nor I_14492 (I249015,I249256,I249188);
not I_14493 (I249321,I249256);
nor I_14494 (I249338,I249321,I249089);
nor I_14495 (I249003,I249157,I249338);
nor I_14496 (I249018,I249256,I249106);
nand I_14497 (I249383,I249239,I249222);
and I_14498 (I249400,I249383,I350805);
nand I_14499 (I249417,I249400,I350802);
not I_14500 (I249434,I249417);
nor I_14501 (I249451,I249434,I350814);
nand I_14502 (I249468,I249205,I249417);
not I_14503 (I249009,I249468);
nor I_14504 (I249499,I350811,I350796);
or I_14505 (I249516,I249499,I350808);
nor I_14506 (I249533,I350802,I350811);
nand I_14507 (I249550,I249533,I249516);
not I_14508 (I249567,I249550);
nor I_14509 (I249030,I249567,I249123);
nand I_14510 (I249598,I249567,I249451);
nand I_14511 (I249006,I249468,I249598);
nor I_14512 (I249629,I249567,I249140);
nor I_14513 (I249027,I249629,I249157);
nor I_14514 (I249021,I249567,I249321);
nor I_14515 (I249674,I249550,I249106);
nor I_14516 (I249691,I249434,I249674);
nor I_14517 (I249012,I249691,I249290);
nor I_14518 (I249722,I249123,I249550);
nor I_14519 (I249739,I249417,I249722);
DFFARX1 I_14520 (I249739,I2898,I249038,I249024,);
not I_14521 (I249803,I2905);
or I_14522 (I249820,I399952,I399964);
nor I_14523 (I249837,I399952,I399964);
nor I_14524 (I249854,I249837,I399946);
not I_14525 (I249871,I249854);
nand I_14526 (I249888,I249820,I399958);
not I_14527 (I249905,I249888);
not I_14528 (I249922,I399952);
nor I_14529 (I249765,I249922,I249905);
nor I_14530 (I249953,I249922,I249888);
nor I_14531 (I249970,I249854,I399952);
not I_14532 (I249987,I399943);
nand I_14533 (I250004,I399961,I399955);
nand I_14534 (I250021,I250004,I399943);
nor I_14535 (I250038,I249888,I250021);
not I_14536 (I250055,I250038);
nor I_14537 (I249780,I250021,I249953);
not I_14538 (I250086,I250021);
nor I_14539 (I250103,I250086,I249854);
nor I_14540 (I249768,I249922,I250103);
nor I_14541 (I249783,I250021,I249871);
nand I_14542 (I250148,I250004,I249987);
and I_14543 (I250165,I250148,I399967);
nand I_14544 (I250182,I250165,I399958);
not I_14545 (I250199,I250182);
nor I_14546 (I250216,I250199,I399952);
nand I_14547 (I250233,I249970,I250182);
not I_14548 (I249774,I250233);
nor I_14549 (I250264,I399955,I399946);
or I_14550 (I250281,I250264,I399943);
nor I_14551 (I250298,I399949,I399949);
nand I_14552 (I250315,I250298,I250281);
not I_14553 (I250332,I250315);
nor I_14554 (I249795,I250332,I249888);
nand I_14555 (I250363,I250332,I250216);
nand I_14556 (I249771,I250233,I250363);
nor I_14557 (I250394,I250332,I249905);
nor I_14558 (I249792,I250394,I249922);
nor I_14559 (I249786,I250332,I250086);
nor I_14560 (I250439,I250315,I249871);
nor I_14561 (I250456,I250199,I250439);
nor I_14562 (I249777,I250456,I250055);
nor I_14563 (I250487,I249888,I250315);
nor I_14564 (I250504,I250182,I250487);
DFFARX1 I_14565 (I250504,I2898,I249803,I249789,);
not I_14566 (I250568,I2905);
or I_14567 (I250585,I180570,I180576);
nor I_14568 (I250602,I180570,I180576);
nor I_14569 (I250619,I250602,I180567);
not I_14570 (I250636,I250619);
nand I_14571 (I250653,I250585,I180558);
not I_14572 (I250670,I250653);
not I_14573 (I250687,I180558);
nor I_14574 (I250530,I250687,I250670);
nor I_14575 (I250718,I250687,I250653);
nor I_14576 (I250735,I250619,I180558);
not I_14577 (I250752,I180564);
nand I_14578 (I250769,I180573,I180585);
nand I_14579 (I250786,I250769,I180564);
nor I_14580 (I250803,I250653,I250786);
not I_14581 (I250820,I250803);
nor I_14582 (I250545,I250786,I250718);
not I_14583 (I250851,I250786);
nor I_14584 (I250868,I250851,I250619);
nor I_14585 (I250533,I250687,I250868);
nor I_14586 (I250548,I250786,I250636);
nand I_14587 (I250913,I250769,I250752);
and I_14588 (I250930,I250913,I180561);
nand I_14589 (I250947,I250930,I180567);
not I_14590 (I250964,I250947);
nor I_14591 (I250981,I250964,I180558);
nand I_14592 (I250998,I250735,I250947);
not I_14593 (I250539,I250998);
nor I_14594 (I251029,I180564,I180582);
or I_14595 (I251046,I251029,I180579);
nor I_14596 (I251063,I180588,I180561);
nand I_14597 (I251080,I251063,I251046);
not I_14598 (I251097,I251080);
nor I_14599 (I250560,I251097,I250653);
nand I_14600 (I251128,I251097,I250981);
nand I_14601 (I250536,I250998,I251128);
nor I_14602 (I251159,I251097,I250670);
nor I_14603 (I250557,I251159,I250687);
nor I_14604 (I250551,I251097,I250851);
nor I_14605 (I251204,I251080,I250636);
nor I_14606 (I251221,I250964,I251204);
nor I_14607 (I250542,I251221,I250820);
nor I_14608 (I251252,I250653,I251080);
nor I_14609 (I251269,I250947,I251252);
DFFARX1 I_14610 (I251269,I2898,I250568,I250554,);
not I_14611 (I251333,I2905);
or I_14612 (I251350,I349609,I349606);
nor I_14613 (I251367,I349609,I349606);
nor I_14614 (I251384,I251367,I349615);
not I_14615 (I251401,I251384);
nand I_14616 (I251418,I251350,I349627);
not I_14617 (I251435,I251418);
not I_14618 (I251452,I349624);
nor I_14619 (I251295,I251452,I251435);
nor I_14620 (I251483,I251452,I251418);
nor I_14621 (I251500,I251384,I349624);
not I_14622 (I251517,I349630);
nand I_14623 (I251534,I349609,I349618);
nand I_14624 (I251551,I251534,I349630);
nor I_14625 (I251568,I251418,I251551);
not I_14626 (I251585,I251568);
nor I_14627 (I251310,I251551,I251483);
not I_14628 (I251616,I251551);
nor I_14629 (I251633,I251616,I251384);
nor I_14630 (I251298,I251452,I251633);
nor I_14631 (I251313,I251551,I251401);
nand I_14632 (I251678,I251534,I251517);
and I_14633 (I251695,I251678,I349615);
nand I_14634 (I251712,I251695,I349612);
not I_14635 (I251729,I251712);
nor I_14636 (I251746,I251729,I349624);
nand I_14637 (I251763,I251500,I251712);
not I_14638 (I251304,I251763);
nor I_14639 (I251794,I349621,I349606);
or I_14640 (I251811,I251794,I349618);
nor I_14641 (I251828,I349612,I349621);
nand I_14642 (I251845,I251828,I251811);
not I_14643 (I251862,I251845);
nor I_14644 (I251325,I251862,I251418);
nand I_14645 (I251893,I251862,I251746);
nand I_14646 (I251301,I251763,I251893);
nor I_14647 (I251924,I251862,I251435);
nor I_14648 (I251322,I251924,I251452);
nor I_14649 (I251316,I251862,I251616);
nor I_14650 (I251969,I251845,I251401);
nor I_14651 (I251986,I251729,I251969);
nor I_14652 (I251307,I251986,I251585);
nor I_14653 (I252017,I251418,I251845);
nor I_14654 (I252034,I251712,I252017);
DFFARX1 I_14655 (I252034,I2898,I251333,I251319,);
not I_14656 (I252098,I2905);
or I_14657 (I252115,I33937,I33925);
nor I_14658 (I252132,I33937,I33925);
nor I_14659 (I252149,I252132,I33928);
not I_14660 (I252166,I252149);
nand I_14661 (I252183,I252115,I33916);
not I_14662 (I252200,I252183);
not I_14663 (I252217,I33940);
nor I_14664 (I252060,I252217,I252200);
nor I_14665 (I252248,I252217,I252183);
nor I_14666 (I252265,I252149,I33940);
not I_14667 (I252282,I33916);
nand I_14668 (I252299,I33931,I33922);
nand I_14669 (I252316,I252299,I33916);
nor I_14670 (I252333,I252183,I252316);
not I_14671 (I252350,I252333);
nor I_14672 (I252075,I252316,I252248);
not I_14673 (I252381,I252316);
nor I_14674 (I252398,I252381,I252149);
nor I_14675 (I252063,I252217,I252398);
nor I_14676 (I252078,I252316,I252166);
nand I_14677 (I252443,I252299,I252282);
and I_14678 (I252460,I252443,I33928);
nand I_14679 (I252477,I252460,I33919);
not I_14680 (I252494,I252477);
nor I_14681 (I252511,I252494,I33940);
nand I_14682 (I252528,I252265,I252477);
not I_14683 (I252069,I252528);
nor I_14684 (I252559,I33919,I33943);
or I_14685 (I252576,I252559,I33934);
nor I_14686 (I252593,I33925,I33922);
nand I_14687 (I252610,I252593,I252576);
not I_14688 (I252627,I252610);
nor I_14689 (I252090,I252627,I252183);
nand I_14690 (I252658,I252627,I252511);
nand I_14691 (I252066,I252528,I252658);
nor I_14692 (I252689,I252627,I252200);
nor I_14693 (I252087,I252689,I252217);
nor I_14694 (I252081,I252627,I252381);
nor I_14695 (I252734,I252610,I252166);
nor I_14696 (I252751,I252494,I252734);
nor I_14697 (I252072,I252751,I252350);
nor I_14698 (I252782,I252183,I252610);
nor I_14699 (I252799,I252477,I252782);
DFFARX1 I_14700 (I252799,I2898,I252098,I252084,);
not I_14701 (I252863,I2905);
or I_14702 (I252880,I306154,I306172);
nor I_14703 (I252897,I306154,I306172);
nor I_14704 (I252914,I252897,I306157);
not I_14705 (I252931,I252914);
nand I_14706 (I252948,I252880,I306166);
not I_14707 (I252965,I252948);
not I_14708 (I252982,I306178);
nor I_14709 (I252825,I252982,I252965);
nor I_14710 (I253013,I252982,I252948);
nor I_14711 (I253030,I252914,I306178);
not I_14712 (I253047,I306175);
nand I_14713 (I253064,I306181,I306154);
nand I_14714 (I253081,I253064,I306175);
nor I_14715 (I253098,I252948,I253081);
not I_14716 (I253115,I253098);
nor I_14717 (I252840,I253081,I253013);
not I_14718 (I253146,I253081);
nor I_14719 (I253163,I253146,I252914);
nor I_14720 (I252828,I252982,I253163);
nor I_14721 (I252843,I253081,I252931);
nand I_14722 (I253208,I253064,I253047);
and I_14723 (I253225,I253208,I306160);
nand I_14724 (I253242,I253225,I306163);
not I_14725 (I253259,I253242);
nor I_14726 (I253276,I253259,I306178);
nand I_14727 (I253293,I253030,I253242);
not I_14728 (I252834,I253293);
nor I_14729 (I253324,I306163,I306184);
or I_14730 (I253341,I253324,I306160);
nor I_14731 (I253358,I306169,I306157);
nand I_14732 (I253375,I253358,I253341);
not I_14733 (I253392,I253375);
nor I_14734 (I252855,I253392,I252948);
nand I_14735 (I253423,I253392,I253276);
nand I_14736 (I252831,I253293,I253423);
nor I_14737 (I253454,I253392,I252965);
nor I_14738 (I252852,I253454,I252982);
nor I_14739 (I252846,I253392,I253146);
nor I_14740 (I253499,I253375,I252931);
nor I_14741 (I253516,I253259,I253499);
nor I_14742 (I252837,I253516,I253115);
nor I_14743 (I253547,I252948,I253375);
nor I_14744 (I253564,I253242,I253547);
DFFARX1 I_14745 (I253564,I2898,I252863,I252849,);
not I_14746 (I253628,I2905);
or I_14747 (I253645,I376452,I376455);
nor I_14748 (I253662,I376452,I376455);
nor I_14749 (I253679,I253662,I376449);
not I_14750 (I253696,I253679);
nand I_14751 (I253713,I253645,I376467);
not I_14752 (I253730,I253713);
not I_14753 (I253747,I376476);
nor I_14754 (I253590,I253747,I253730);
nor I_14755 (I253778,I253747,I253713);
nor I_14756 (I253795,I253679,I376476);
not I_14757 (I253812,I376461);
nand I_14758 (I253829,I376449,I376458);
nand I_14759 (I253846,I253829,I376461);
nor I_14760 (I253863,I253713,I253846);
not I_14761 (I253880,I253863);
nor I_14762 (I253605,I253846,I253778);
not I_14763 (I253911,I253846);
nor I_14764 (I253928,I253911,I253679);
nor I_14765 (I253593,I253747,I253928);
nor I_14766 (I253608,I253846,I253696);
nand I_14767 (I253973,I253829,I253812);
and I_14768 (I253990,I253973,I376452);
nand I_14769 (I254007,I253990,I376455);
not I_14770 (I254024,I254007);
nor I_14771 (I254041,I254024,I376476);
nand I_14772 (I254058,I253795,I254007);
not I_14773 (I253599,I254058);
nor I_14774 (I254089,I376479,I376464);
or I_14775 (I254106,I254089,I376473);
nor I_14776 (I254123,I376482,I376470);
nand I_14777 (I254140,I254123,I254106);
not I_14778 (I254157,I254140);
nor I_14779 (I253620,I254157,I253713);
nand I_14780 (I254188,I254157,I254041);
nand I_14781 (I253596,I254058,I254188);
nor I_14782 (I254219,I254157,I253730);
nor I_14783 (I253617,I254219,I253747);
nor I_14784 (I253611,I254157,I253911);
nor I_14785 (I254264,I254140,I253696);
nor I_14786 (I254281,I254024,I254264);
nor I_14787 (I253602,I254281,I253880);
nor I_14788 (I254312,I253713,I254140);
nor I_14789 (I254329,I254007,I254312);
DFFARX1 I_14790 (I254329,I2898,I253628,I253614,);
not I_14791 (I254393,I2905);
or I_14792 (I254410,I414332,I414329);
nor I_14793 (I254427,I414332,I414329);
nor I_14794 (I254444,I254427,I414317);
not I_14795 (I254461,I254444);
nand I_14796 (I254478,I254410,I414338);
not I_14797 (I254495,I254478);
not I_14798 (I254512,I414308);
nor I_14799 (I254355,I254512,I254495);
nor I_14800 (I254543,I254512,I254478);
nor I_14801 (I254560,I254444,I414308);
not I_14802 (I254577,I414326);
nand I_14803 (I254594,I414341,I414323);
nand I_14804 (I254611,I254594,I414326);
nor I_14805 (I254628,I254478,I254611);
not I_14806 (I254645,I254628);
nor I_14807 (I254370,I254611,I254543);
not I_14808 (I254676,I254611);
nor I_14809 (I254693,I254676,I254444);
nor I_14810 (I254358,I254512,I254693);
nor I_14811 (I254373,I254611,I254461);
nand I_14812 (I254738,I254594,I254577);
and I_14813 (I254755,I254738,I414335);
nand I_14814 (I254772,I254755,I414314);
not I_14815 (I254789,I254772);
nor I_14816 (I254806,I254789,I414308);
nand I_14817 (I254823,I254560,I254772);
not I_14818 (I254364,I254823);
nor I_14819 (I254854,I414320,I414308);
or I_14820 (I254871,I254854,I414311);
nor I_14821 (I254888,I414311,I414314);
nand I_14822 (I254905,I254888,I254871);
not I_14823 (I254922,I254905);
nor I_14824 (I254385,I254922,I254478);
nand I_14825 (I254953,I254922,I254806);
nand I_14826 (I254361,I254823,I254953);
nor I_14827 (I254984,I254922,I254495);
nor I_14828 (I254382,I254984,I254512);
nor I_14829 (I254376,I254922,I254676);
nor I_14830 (I255029,I254905,I254461);
nor I_14831 (I255046,I254789,I255029);
nor I_14832 (I254367,I255046,I254645);
nor I_14833 (I255077,I254478,I254905);
nor I_14834 (I255094,I254772,I255077);
DFFARX1 I_14835 (I255094,I2898,I254393,I254379,);
not I_14836 (I255158,I2905);
or I_14837 (I255175,I193903,I193903);
nor I_14838 (I255192,I193903,I193903);
nor I_14839 (I255209,I255192,I193918);
not I_14840 (I255226,I255209);
nand I_14841 (I255243,I255175,I193915);
not I_14842 (I255260,I255243);
not I_14843 (I255277,I193927);
nor I_14844 (I255120,I255277,I255260);
nor I_14845 (I255308,I255277,I255243);
nor I_14846 (I255325,I255209,I193927);
not I_14847 (I255342,I193906);
nand I_14848 (I255359,I193918,I193909);
nand I_14849 (I255376,I255359,I193906);
nor I_14850 (I255393,I255243,I255376);
not I_14851 (I255410,I255393);
nor I_14852 (I255135,I255376,I255308);
not I_14853 (I255441,I255376);
nor I_14854 (I255458,I255441,I255209);
nor I_14855 (I255123,I255277,I255458);
nor I_14856 (I255138,I255376,I255226);
nand I_14857 (I255503,I255359,I255342);
and I_14858 (I255520,I255503,I193915);
nand I_14859 (I255537,I255520,I193909);
not I_14860 (I255554,I255537);
nor I_14861 (I255571,I255554,I193927);
nand I_14862 (I255588,I255325,I255537);
not I_14863 (I255129,I255588);
nor I_14864 (I255619,I193912,I193912);
or I_14865 (I255636,I255619,I193906);
nor I_14866 (I255653,I193921,I193924);
nand I_14867 (I255670,I255653,I255636);
not I_14868 (I255687,I255670);
nor I_14869 (I255150,I255687,I255243);
nand I_14870 (I255718,I255687,I255571);
nand I_14871 (I255126,I255588,I255718);
nor I_14872 (I255749,I255687,I255260);
nor I_14873 (I255147,I255749,I255277);
nor I_14874 (I255141,I255687,I255441);
nor I_14875 (I255794,I255670,I255226);
nor I_14876 (I255811,I255554,I255794);
nor I_14877 (I255132,I255811,I255410);
nor I_14878 (I255842,I255243,I255670);
nor I_14879 (I255859,I255537,I255842);
DFFARX1 I_14880 (I255859,I2898,I255158,I255144,);
not I_14881 (I255923,I2905);
or I_14882 (I255940,I17515,I17503);
nor I_14883 (I255957,I17515,I17503);
nor I_14884 (I255974,I255957,I17506);
not I_14885 (I255991,I255974);
nand I_14886 (I256008,I255940,I17494);
not I_14887 (I256025,I256008);
not I_14888 (I256042,I17518);
nor I_14889 (I255885,I256042,I256025);
nor I_14890 (I256073,I256042,I256008);
nor I_14891 (I256090,I255974,I17518);
not I_14892 (I256107,I17494);
nand I_14893 (I256124,I17509,I17500);
nand I_14894 (I256141,I256124,I17494);
nor I_14895 (I256158,I256008,I256141);
not I_14896 (I256175,I256158);
nor I_14897 (I255900,I256141,I256073);
not I_14898 (I256206,I256141);
nor I_14899 (I256223,I256206,I255974);
nor I_14900 (I255888,I256042,I256223);
nor I_14901 (I255903,I256141,I255991);
nand I_14902 (I256268,I256124,I256107);
and I_14903 (I256285,I256268,I17506);
nand I_14904 (I256302,I256285,I17497);
not I_14905 (I256319,I256302);
nor I_14906 (I256336,I256319,I17518);
nand I_14907 (I256353,I256090,I256302);
not I_14908 (I255894,I256353);
nor I_14909 (I256384,I17497,I17521);
or I_14910 (I256401,I256384,I17512);
nor I_14911 (I256418,I17503,I17500);
nand I_14912 (I256435,I256418,I256401);
not I_14913 (I256452,I256435);
nor I_14914 (I255915,I256452,I256008);
nand I_14915 (I256483,I256452,I256336);
nand I_14916 (I255891,I256353,I256483);
nor I_14917 (I256514,I256452,I256025);
nor I_14918 (I255912,I256514,I256042);
nor I_14919 (I255906,I256452,I256206);
nor I_14920 (I256559,I256435,I255991);
nor I_14921 (I256576,I256319,I256559);
nor I_14922 (I255897,I256576,I256175);
nor I_14923 (I256607,I256008,I256435);
nor I_14924 (I256624,I256302,I256607);
DFFARX1 I_14925 (I256624,I2898,I255923,I255909,);
not I_14926 (I256688,I2905);
or I_14927 (I256705,I340684,I340681);
nor I_14928 (I256722,I340684,I340681);
nor I_14929 (I256739,I256722,I340690);
not I_14930 (I256756,I256739);
nand I_14931 (I256773,I256705,I340702);
not I_14932 (I256790,I256773);
not I_14933 (I256807,I340699);
nor I_14934 (I256650,I256807,I256790);
nor I_14935 (I256838,I256807,I256773);
nor I_14936 (I256855,I256739,I340699);
not I_14937 (I256872,I340705);
nand I_14938 (I256889,I340684,I340693);
nand I_14939 (I256906,I256889,I340705);
nor I_14940 (I256923,I256773,I256906);
not I_14941 (I256940,I256923);
nor I_14942 (I256665,I256906,I256838);
not I_14943 (I256971,I256906);
nor I_14944 (I256988,I256971,I256739);
nor I_14945 (I256653,I256807,I256988);
nor I_14946 (I256668,I256906,I256756);
nand I_14947 (I257033,I256889,I256872);
and I_14948 (I257050,I257033,I340690);
nand I_14949 (I257067,I257050,I340687);
not I_14950 (I257084,I257067);
nor I_14951 (I257101,I257084,I340699);
nand I_14952 (I257118,I256855,I257067);
not I_14953 (I256659,I257118);
nor I_14954 (I257149,I340696,I340681);
or I_14955 (I257166,I257149,I340693);
nor I_14956 (I257183,I340687,I340696);
nand I_14957 (I257200,I257183,I257166);
not I_14958 (I257217,I257200);
nor I_14959 (I256680,I257217,I256773);
nand I_14960 (I257248,I257217,I257101);
nand I_14961 (I256656,I257118,I257248);
nor I_14962 (I257279,I257217,I256790);
nor I_14963 (I256677,I257279,I256807);
nor I_14964 (I256671,I257217,I256971);
nor I_14965 (I257324,I257200,I256756);
nor I_14966 (I257341,I257084,I257324);
nor I_14967 (I256662,I257341,I256940);
nor I_14968 (I257372,I256773,I257200);
nor I_14969 (I257389,I257067,I257372);
DFFARX1 I_14970 (I257389,I2898,I256688,I256674,);
not I_14971 (I257453,I2905);
or I_14972 (I257470,I435939,I435936);
nor I_14973 (I257487,I435939,I435936);
nor I_14974 (I257504,I257487,I435924);
not I_14975 (I257521,I257504);
nand I_14976 (I257538,I257470,I435945);
not I_14977 (I257555,I257538);
not I_14978 (I257572,I435915);
nor I_14979 (I257415,I257572,I257555);
nor I_14980 (I257603,I257572,I257538);
nor I_14981 (I257620,I257504,I435915);
not I_14982 (I257637,I435933);
nand I_14983 (I257654,I435948,I435930);
nand I_14984 (I257671,I257654,I435933);
nor I_14985 (I257688,I257538,I257671);
not I_14986 (I257705,I257688);
nor I_14987 (I257430,I257671,I257603);
not I_14988 (I257736,I257671);
nor I_14989 (I257753,I257736,I257504);
nor I_14990 (I257418,I257572,I257753);
nor I_14991 (I257433,I257671,I257521);
nand I_14992 (I257798,I257654,I257637);
and I_14993 (I257815,I257798,I435942);
nand I_14994 (I257832,I257815,I435921);
not I_14995 (I257849,I257832);
nor I_14996 (I257866,I257849,I435915);
nand I_14997 (I257883,I257620,I257832);
not I_14998 (I257424,I257883);
nor I_14999 (I257914,I435927,I435915);
or I_15000 (I257931,I257914,I435918);
nor I_15001 (I257948,I435918,I435921);
nand I_15002 (I257965,I257948,I257931);
not I_15003 (I257982,I257965);
nor I_15004 (I257445,I257982,I257538);
nand I_15005 (I258013,I257982,I257866);
nand I_15006 (I257421,I257883,I258013);
nor I_15007 (I258044,I257982,I257555);
nor I_15008 (I257442,I258044,I257572);
nor I_15009 (I257436,I257982,I257736);
nor I_15010 (I258089,I257965,I257521);
nor I_15011 (I258106,I257849,I258089);
nor I_15012 (I257427,I258106,I257705);
nor I_15013 (I258137,I257538,I257965);
nor I_15014 (I258154,I257832,I258137);
DFFARX1 I_15015 (I258154,I2898,I257453,I257439,);
not I_15016 (I258218,I2905);
or I_15017 (I258235,I408792,I408804);
nor I_15018 (I258252,I408792,I408804);
nor I_15019 (I258269,I258252,I408786);
not I_15020 (I258286,I258269);
nand I_15021 (I258303,I258235,I408798);
not I_15022 (I258320,I258303);
not I_15023 (I258337,I408792);
nor I_15024 (I258180,I258337,I258320);
nor I_15025 (I258368,I258337,I258303);
nor I_15026 (I258385,I258269,I408792);
not I_15027 (I258402,I408783);
nand I_15028 (I258419,I408801,I408795);
nand I_15029 (I258436,I258419,I408783);
nor I_15030 (I258453,I258303,I258436);
not I_15031 (I258470,I258453);
nor I_15032 (I258195,I258436,I258368);
not I_15033 (I258501,I258436);
nor I_15034 (I258518,I258501,I258269);
nor I_15035 (I258183,I258337,I258518);
nor I_15036 (I258198,I258436,I258286);
nand I_15037 (I258563,I258419,I258402);
and I_15038 (I258580,I258563,I408807);
nand I_15039 (I258597,I258580,I408798);
not I_15040 (I258614,I258597);
nor I_15041 (I258631,I258614,I408792);
nand I_15042 (I258648,I258385,I258597);
not I_15043 (I258189,I258648);
nor I_15044 (I258679,I408795,I408786);
or I_15045 (I258696,I258679,I408783);
nor I_15046 (I258713,I408789,I408789);
nand I_15047 (I258730,I258713,I258696);
not I_15048 (I258747,I258730);
nor I_15049 (I258210,I258747,I258303);
nand I_15050 (I258778,I258747,I258631);
nand I_15051 (I258186,I258648,I258778);
nor I_15052 (I258809,I258747,I258320);
nor I_15053 (I258207,I258809,I258337);
nor I_15054 (I258201,I258747,I258501);
nor I_15055 (I258854,I258730,I258286);
nor I_15056 (I258871,I258614,I258854);
nor I_15057 (I258192,I258871,I258470);
nor I_15058 (I258902,I258303,I258730);
nor I_15059 (I258919,I258597,I258902);
DFFARX1 I_15060 (I258919,I2898,I258218,I258204,);
not I_15061 (I258983,I2905);
or I_15062 (I259000,I85251,I85263);
nor I_15063 (I259017,I85251,I85263);
nor I_15064 (I259034,I259017,I85260);
not I_15065 (I259051,I259034);
nand I_15066 (I259068,I259000,I85254);
not I_15067 (I259085,I259068);
not I_15068 (I259102,I85248);
nor I_15069 (I258945,I259102,I259085);
nor I_15070 (I259133,I259102,I259068);
nor I_15071 (I259150,I259034,I85248);
not I_15072 (I259167,I85257);
nand I_15073 (I259184,I85245,I85242);
nand I_15074 (I259201,I259184,I85257);
nor I_15075 (I259218,I259068,I259201);
not I_15076 (I259235,I259218);
nor I_15077 (I258960,I259201,I259133);
not I_15078 (I259266,I259201);
nor I_15079 (I259283,I259266,I259034);
nor I_15080 (I258948,I259102,I259283);
nor I_15081 (I258963,I259201,I259051);
nand I_15082 (I259328,I259184,I259167);
and I_15083 (I259345,I259328,I85251);
nand I_15084 (I259362,I259345,I85239);
not I_15085 (I259379,I259362);
nor I_15086 (I259396,I259379,I85248);
nand I_15087 (I259413,I259150,I259362);
not I_15088 (I258954,I259413);
nor I_15089 (I259444,I85245,I85242);
or I_15090 (I259461,I259444,I85248);
nor I_15091 (I259478,I85239,I85266);
nand I_15092 (I259495,I259478,I259461);
not I_15093 (I259512,I259495);
nor I_15094 (I258975,I259512,I259068);
nand I_15095 (I259543,I259512,I259396);
nand I_15096 (I258951,I259413,I259543);
nor I_15097 (I259574,I259512,I259085);
nor I_15098 (I258972,I259574,I259102);
nor I_15099 (I258966,I259512,I259266);
nor I_15100 (I259619,I259495,I259051);
nor I_15101 (I259636,I259379,I259619);
nor I_15102 (I258957,I259636,I259235);
nor I_15103 (I259667,I259068,I259495);
nor I_15104 (I259684,I259362,I259667);
DFFARX1 I_15105 (I259684,I2898,I258983,I258969,);
not I_15106 (I259748,I2905);
or I_15107 (I259765,I291534,I291552);
nor I_15108 (I259782,I291534,I291552);
nor I_15109 (I259799,I259782,I291537);
not I_15110 (I259816,I259799);
nand I_15111 (I259833,I259765,I291546);
not I_15112 (I259850,I259833);
not I_15113 (I259867,I291558);
nor I_15114 (I259710,I259867,I259850);
nor I_15115 (I259898,I259867,I259833);
nor I_15116 (I259915,I259799,I291558);
not I_15117 (I259932,I291555);
nand I_15118 (I259949,I291561,I291534);
nand I_15119 (I259966,I259949,I291555);
nor I_15120 (I259983,I259833,I259966);
not I_15121 (I260000,I259983);
nor I_15122 (I259725,I259966,I259898);
not I_15123 (I260031,I259966);
nor I_15124 (I260048,I260031,I259799);
nor I_15125 (I259713,I259867,I260048);
nor I_15126 (I259728,I259966,I259816);
nand I_15127 (I260093,I259949,I259932);
and I_15128 (I260110,I260093,I291540);
nand I_15129 (I260127,I260110,I291543);
not I_15130 (I260144,I260127);
nor I_15131 (I260161,I260144,I291558);
nand I_15132 (I260178,I259915,I260127);
not I_15133 (I259719,I260178);
nor I_15134 (I260209,I291543,I291564);
or I_15135 (I260226,I260209,I291540);
nor I_15136 (I260243,I291549,I291537);
nand I_15137 (I260260,I260243,I260226);
not I_15138 (I260277,I260260);
nor I_15139 (I259740,I260277,I259833);
nand I_15140 (I260308,I260277,I260161);
nand I_15141 (I259716,I260178,I260308);
nor I_15142 (I260339,I260277,I259850);
nor I_15143 (I259737,I260339,I259867);
nor I_15144 (I259731,I260277,I260031);
nor I_15145 (I260384,I260260,I259816);
nor I_15146 (I260401,I260144,I260384);
nor I_15147 (I259722,I260401,I260000);
nor I_15148 (I260432,I259833,I260260);
nor I_15149 (I260449,I260127,I260432);
DFFARX1 I_15150 (I260449,I2898,I259748,I259734,);
not I_15151 (I260513,I2905);
or I_15152 (I260530,I136161,I136158);
nor I_15153 (I260547,I136161,I136158);
nor I_15154 (I260564,I260547,I136143);
not I_15155 (I260581,I260564);
nand I_15156 (I260598,I260530,I136164);
not I_15157 (I260615,I260598);
not I_15158 (I260632,I136146);
nor I_15159 (I260475,I260632,I260615);
nor I_15160 (I260663,I260632,I260598);
nor I_15161 (I260680,I260564,I136146);
not I_15162 (I260697,I136140);
nand I_15163 (I260714,I136149,I136137);
nand I_15164 (I260731,I260714,I136140);
nor I_15165 (I260748,I260598,I260731);
not I_15166 (I260765,I260748);
nor I_15167 (I260490,I260731,I260663);
not I_15168 (I260796,I260731);
nor I_15169 (I260813,I260796,I260564);
nor I_15170 (I260478,I260632,I260813);
nor I_15171 (I260493,I260731,I260581);
nand I_15172 (I260858,I260714,I260697);
and I_15173 (I260875,I260858,I136170);
nand I_15174 (I260892,I260875,I136167);
not I_15175 (I260909,I260892);
nor I_15176 (I260926,I260909,I136146);
nand I_15177 (I260943,I260680,I260892);
not I_15178 (I260484,I260943);
nor I_15179 (I260974,I136137,I136155);
or I_15180 (I260991,I260974,I136140);
nor I_15181 (I261008,I136152,I136143);
nand I_15182 (I261025,I261008,I260991);
not I_15183 (I261042,I261025);
nor I_15184 (I260505,I261042,I260598);
nand I_15185 (I261073,I261042,I260926);
nand I_15186 (I260481,I260943,I261073);
nor I_15187 (I261104,I261042,I260615);
nor I_15188 (I260502,I261104,I260632);
nor I_15189 (I260496,I261042,I260796);
nor I_15190 (I261149,I261025,I260581);
nor I_15191 (I261166,I260909,I261149);
nor I_15192 (I260487,I261166,I260765);
nor I_15193 (I261197,I260598,I261025);
nor I_15194 (I261214,I260892,I261197);
DFFARX1 I_15195 (I261214,I2898,I260513,I260499,);
not I_15196 (I261278,I2905);
or I_15197 (I261295,I29653,I29641);
nor I_15198 (I261312,I29653,I29641);
nor I_15199 (I261329,I261312,I29644);
not I_15200 (I261346,I261329);
nand I_15201 (I261363,I261295,I29632);
not I_15202 (I261380,I261363);
not I_15203 (I261397,I29656);
nor I_15204 (I261240,I261397,I261380);
nor I_15205 (I261428,I261397,I261363);
nor I_15206 (I261445,I261329,I29656);
not I_15207 (I261462,I29632);
nand I_15208 (I261479,I29647,I29638);
nand I_15209 (I261496,I261479,I29632);
nor I_15210 (I261513,I261363,I261496);
not I_15211 (I261530,I261513);
nor I_15212 (I261255,I261496,I261428);
not I_15213 (I261561,I261496);
nor I_15214 (I261578,I261561,I261329);
nor I_15215 (I261243,I261397,I261578);
nor I_15216 (I261258,I261496,I261346);
nand I_15217 (I261623,I261479,I261462);
and I_15218 (I261640,I261623,I29644);
nand I_15219 (I261657,I261640,I29635);
not I_15220 (I261674,I261657);
nor I_15221 (I261691,I261674,I29656);
nand I_15222 (I261708,I261445,I261657);
not I_15223 (I261249,I261708);
nor I_15224 (I261739,I29635,I29659);
or I_15225 (I261756,I261739,I29650);
nor I_15226 (I261773,I29641,I29638);
nand I_15227 (I261790,I261773,I261756);
not I_15228 (I261807,I261790);
nor I_15229 (I261270,I261807,I261363);
nand I_15230 (I261838,I261807,I261691);
nand I_15231 (I261246,I261708,I261838);
nor I_15232 (I261869,I261807,I261380);
nor I_15233 (I261267,I261869,I261397);
nor I_15234 (I261261,I261807,I261561);
nor I_15235 (I261914,I261790,I261346);
nor I_15236 (I261931,I261674,I261914);
nor I_15237 (I261252,I261931,I261530);
nor I_15238 (I261962,I261363,I261790);
nor I_15239 (I261979,I261657,I261962);
DFFARX1 I_15240 (I261979,I2898,I261278,I261264,);
not I_15241 (I262043,I2905);
or I_15242 (I262060,I39649,I39637);
nor I_15243 (I262077,I39649,I39637);
nor I_15244 (I262094,I262077,I39640);
not I_15245 (I262111,I262094);
nand I_15246 (I262128,I262060,I39628);
not I_15247 (I262145,I262128);
not I_15248 (I262162,I39652);
nor I_15249 (I262005,I262162,I262145);
nor I_15250 (I262193,I262162,I262128);
nor I_15251 (I262210,I262094,I39652);
not I_15252 (I262227,I39628);
nand I_15253 (I262244,I39643,I39634);
nand I_15254 (I262261,I262244,I39628);
nor I_15255 (I262278,I262128,I262261);
not I_15256 (I262295,I262278);
nor I_15257 (I262020,I262261,I262193);
not I_15258 (I262326,I262261);
nor I_15259 (I262343,I262326,I262094);
nor I_15260 (I262008,I262162,I262343);
nor I_15261 (I262023,I262261,I262111);
nand I_15262 (I262388,I262244,I262227);
and I_15263 (I262405,I262388,I39640);
nand I_15264 (I262422,I262405,I39631);
not I_15265 (I262439,I262422);
nor I_15266 (I262456,I262439,I39652);
nand I_15267 (I262473,I262210,I262422);
not I_15268 (I262014,I262473);
nor I_15269 (I262504,I39631,I39655);
or I_15270 (I262521,I262504,I39646);
nor I_15271 (I262538,I39637,I39634);
nand I_15272 (I262555,I262538,I262521);
not I_15273 (I262572,I262555);
nor I_15274 (I262035,I262572,I262128);
nand I_15275 (I262603,I262572,I262456);
nand I_15276 (I262011,I262473,I262603);
nor I_15277 (I262634,I262572,I262145);
nor I_15278 (I262032,I262634,I262162);
nor I_15279 (I262026,I262572,I262326);
nor I_15280 (I262679,I262555,I262111);
nor I_15281 (I262696,I262439,I262679);
nor I_15282 (I262017,I262696,I262295);
nor I_15283 (I262727,I262128,I262555);
nor I_15284 (I262744,I262422,I262727);
DFFARX1 I_15285 (I262744,I2898,I262043,I262029,);
not I_15286 (I262808,I2905);
or I_15287 (I262825,I436636,I436633);
nor I_15288 (I262842,I436636,I436633);
nor I_15289 (I262859,I262842,I436621);
not I_15290 (I262876,I262859);
nand I_15291 (I262893,I262825,I436642);
not I_15292 (I262910,I262893);
not I_15293 (I262927,I436612);
nor I_15294 (I262770,I262927,I262910);
nor I_15295 (I262958,I262927,I262893);
nor I_15296 (I262975,I262859,I436612);
not I_15297 (I262992,I436630);
nand I_15298 (I263009,I436645,I436627);
nand I_15299 (I263026,I263009,I436630);
nor I_15300 (I263043,I262893,I263026);
not I_15301 (I263060,I263043);
nor I_15302 (I262785,I263026,I262958);
not I_15303 (I263091,I263026);
nor I_15304 (I263108,I263091,I262859);
nor I_15305 (I262773,I262927,I263108);
nor I_15306 (I262788,I263026,I262876);
nand I_15307 (I263153,I263009,I262992);
and I_15308 (I263170,I263153,I436639);
nand I_15309 (I263187,I263170,I436618);
not I_15310 (I263204,I263187);
nor I_15311 (I263221,I263204,I436612);
nand I_15312 (I263238,I262975,I263187);
not I_15313 (I262779,I263238);
nor I_15314 (I263269,I436624,I436612);
or I_15315 (I263286,I263269,I436615);
nor I_15316 (I263303,I436615,I436618);
nand I_15317 (I263320,I263303,I263286);
not I_15318 (I263337,I263320);
nor I_15319 (I262800,I263337,I262893);
nand I_15320 (I263368,I263337,I263221);
nand I_15321 (I262776,I263238,I263368);
nor I_15322 (I263399,I263337,I262910);
nor I_15323 (I262797,I263399,I262927);
nor I_15324 (I262791,I263337,I263091);
nor I_15325 (I263444,I263320,I262876);
nor I_15326 (I263461,I263204,I263444);
nor I_15327 (I262782,I263461,I263060);
nor I_15328 (I263492,I262893,I263320);
nor I_15329 (I263509,I263187,I263492);
DFFARX1 I_15330 (I263509,I2898,I262808,I262794,);
not I_15331 (I263573,I2905);
or I_15332 (I263590,I197388,I197388);
nor I_15333 (I263607,I197388,I197388);
nor I_15334 (I263624,I263607,I197403);
not I_15335 (I263641,I263624);
nand I_15336 (I263658,I263590,I197400);
not I_15337 (I263675,I263658);
not I_15338 (I263692,I197412);
nor I_15339 (I263535,I263692,I263675);
nor I_15340 (I263723,I263692,I263658);
nor I_15341 (I263740,I263624,I197412);
not I_15342 (I263757,I197391);
nand I_15343 (I263774,I197403,I197394);
nand I_15344 (I263791,I263774,I197391);
nor I_15345 (I263808,I263658,I263791);
not I_15346 (I263825,I263808);
nor I_15347 (I263550,I263791,I263723);
not I_15348 (I263856,I263791);
nor I_15349 (I263873,I263856,I263624);
nor I_15350 (I263538,I263692,I263873);
nor I_15351 (I263553,I263791,I263641);
nand I_15352 (I263918,I263774,I263757);
and I_15353 (I263935,I263918,I197400);
nand I_15354 (I263952,I263935,I197394);
not I_15355 (I263969,I263952);
nor I_15356 (I263986,I263969,I197412);
nand I_15357 (I264003,I263740,I263952);
not I_15358 (I263544,I264003);
nor I_15359 (I264034,I197397,I197397);
or I_15360 (I264051,I264034,I197391);
nor I_15361 (I264068,I197406,I197409);
nand I_15362 (I264085,I264068,I264051);
not I_15363 (I264102,I264085);
nor I_15364 (I263565,I264102,I263658);
nand I_15365 (I264133,I264102,I263986);
nand I_15366 (I263541,I264003,I264133);
nor I_15367 (I264164,I264102,I263675);
nor I_15368 (I263562,I264164,I263692);
nor I_15369 (I263556,I264102,I263856);
nor I_15370 (I264209,I264085,I263641);
nor I_15371 (I264226,I263969,I264209);
nor I_15372 (I263547,I264226,I263825);
nor I_15373 (I264257,I263658,I264085);
nor I_15374 (I264274,I263952,I264257);
DFFARX1 I_15375 (I264274,I2898,I263573,I263559,);
not I_15376 (I264338,I2905);
or I_15377 (I264355,I50396,I50372);
nor I_15378 (I264372,I50396,I50372);
nor I_15379 (I264389,I264372,I50384);
not I_15380 (I264406,I264389);
nand I_15381 (I264423,I264355,I50381);
not I_15382 (I264440,I264423);
not I_15383 (I264457,I50378);
nor I_15384 (I264300,I264457,I264440);
nor I_15385 (I264488,I264457,I264423);
nor I_15386 (I264505,I264389,I50378);
not I_15387 (I264522,I50387);
nand I_15388 (I264539,I50405,I50372);
nand I_15389 (I264556,I264539,I50387);
nor I_15390 (I264573,I264423,I264556);
not I_15391 (I264590,I264573);
nor I_15392 (I264315,I264556,I264488);
not I_15393 (I264621,I264556);
nor I_15394 (I264638,I264621,I264389);
nor I_15395 (I264303,I264457,I264638);
nor I_15396 (I264318,I264556,I264406);
nand I_15397 (I264683,I264539,I264522);
and I_15398 (I264700,I264683,I50408);
nand I_15399 (I264717,I264700,I50399);
not I_15400 (I264734,I264717);
nor I_15401 (I264751,I264734,I50378);
nand I_15402 (I264768,I264505,I264717);
not I_15403 (I264309,I264768);
nor I_15404 (I264799,I50375,I50390);
or I_15405 (I264816,I264799,I50375);
nor I_15406 (I264833,I50393,I50402);
nand I_15407 (I264850,I264833,I264816);
not I_15408 (I264867,I264850);
nor I_15409 (I264330,I264867,I264423);
nand I_15410 (I264898,I264867,I264751);
nand I_15411 (I264306,I264768,I264898);
nor I_15412 (I264929,I264867,I264440);
nor I_15413 (I264327,I264929,I264457);
nor I_15414 (I264321,I264867,I264621);
nor I_15415 (I264974,I264850,I264406);
nor I_15416 (I264991,I264734,I264974);
nor I_15417 (I264312,I264991,I264590);
nor I_15418 (I265022,I264423,I264850);
nor I_15419 (I265039,I264717,I265022);
DFFARX1 I_15420 (I265039,I2898,I264338,I264324,);
not I_15421 (I265103,I2905);
or I_15422 (I265120,I319312,I319330);
nor I_15423 (I265137,I319312,I319330);
nor I_15424 (I265154,I265137,I319315);
not I_15425 (I265171,I265154);
nand I_15426 (I265188,I265120,I319324);
not I_15427 (I265205,I265188);
not I_15428 (I265222,I319336);
nor I_15429 (I265065,I265222,I265205);
nor I_15430 (I265253,I265222,I265188);
nor I_15431 (I265270,I265154,I319336);
not I_15432 (I265287,I319333);
nand I_15433 (I265304,I319339,I319312);
nand I_15434 (I265321,I265304,I319333);
nor I_15435 (I265338,I265188,I265321);
not I_15436 (I265355,I265338);
nor I_15437 (I265080,I265321,I265253);
not I_15438 (I265386,I265321);
nor I_15439 (I265403,I265386,I265154);
nor I_15440 (I265068,I265222,I265403);
nor I_15441 (I265083,I265321,I265171);
nand I_15442 (I265448,I265304,I265287);
and I_15443 (I265465,I265448,I319318);
nand I_15444 (I265482,I265465,I319321);
not I_15445 (I265499,I265482);
nor I_15446 (I265516,I265499,I319336);
nand I_15447 (I265533,I265270,I265482);
not I_15448 (I265074,I265533);
nor I_15449 (I265564,I319321,I319342);
or I_15450 (I265581,I265564,I319318);
nor I_15451 (I265598,I319327,I319315);
nand I_15452 (I265615,I265598,I265581);
not I_15453 (I265632,I265615);
nor I_15454 (I265095,I265632,I265188);
nand I_15455 (I265663,I265632,I265516);
nand I_15456 (I265071,I265533,I265663);
nor I_15457 (I265694,I265632,I265205);
nor I_15458 (I265092,I265694,I265222);
nor I_15459 (I265086,I265632,I265386);
nor I_15460 (I265739,I265615,I265171);
nor I_15461 (I265756,I265499,I265739);
nor I_15462 (I265077,I265756,I265355);
nor I_15463 (I265787,I265188,I265615);
nor I_15464 (I265804,I265482,I265787);
DFFARX1 I_15465 (I265804,I2898,I265103,I265089,);
not I_15466 (I265868,I2905);
or I_15467 (I265885,I313464,I313482);
nor I_15468 (I265902,I313464,I313482);
nor I_15469 (I265919,I265902,I313467);
not I_15470 (I265936,I265919);
nand I_15471 (I265953,I265885,I313476);
not I_15472 (I265970,I265953);
not I_15473 (I265987,I313488);
nor I_15474 (I265830,I265987,I265970);
nor I_15475 (I266018,I265987,I265953);
nor I_15476 (I266035,I265919,I313488);
not I_15477 (I266052,I313485);
nand I_15478 (I266069,I313491,I313464);
nand I_15479 (I266086,I266069,I313485);
nor I_15480 (I266103,I265953,I266086);
not I_15481 (I266120,I266103);
nor I_15482 (I265845,I266086,I266018);
not I_15483 (I266151,I266086);
nor I_15484 (I266168,I266151,I265919);
nor I_15485 (I265833,I265987,I266168);
nor I_15486 (I265848,I266086,I265936);
nand I_15487 (I266213,I266069,I266052);
and I_15488 (I266230,I266213,I313470);
nand I_15489 (I266247,I266230,I313473);
not I_15490 (I266264,I266247);
nor I_15491 (I266281,I266264,I313488);
nand I_15492 (I266298,I266035,I266247);
not I_15493 (I265839,I266298);
nor I_15494 (I266329,I313473,I313494);
or I_15495 (I266346,I266329,I313470);
nor I_15496 (I266363,I313479,I313467);
nand I_15497 (I266380,I266363,I266346);
not I_15498 (I266397,I266380);
nor I_15499 (I265860,I266397,I265953);
nand I_15500 (I266428,I266397,I266281);
nand I_15501 (I265836,I266298,I266428);
nor I_15502 (I266459,I266397,I265970);
nor I_15503 (I265857,I266459,I265987);
nor I_15504 (I265851,I266397,I266151);
nor I_15505 (I266504,I266380,I265936);
nor I_15506 (I266521,I266264,I266504);
nor I_15507 (I265842,I266521,I266120);
nor I_15508 (I266552,I265953,I266380);
nor I_15509 (I266569,I266247,I266552);
DFFARX1 I_15510 (I266569,I2898,I265868,I265854,);
not I_15511 (I266633,I2905);
or I_15512 (I266650,I338304,I338301);
nor I_15513 (I266667,I338304,I338301);
nor I_15514 (I266684,I266667,I338310);
not I_15515 (I266701,I266684);
nand I_15516 (I266718,I266650,I338322);
not I_15517 (I266735,I266718);
not I_15518 (I266752,I338319);
nor I_15519 (I266595,I266752,I266735);
nor I_15520 (I266783,I266752,I266718);
nor I_15521 (I266800,I266684,I338319);
not I_15522 (I266817,I338325);
nand I_15523 (I266834,I338304,I338313);
nand I_15524 (I266851,I266834,I338325);
nor I_15525 (I266868,I266718,I266851);
not I_15526 (I266885,I266868);
nor I_15527 (I266610,I266851,I266783);
not I_15528 (I266916,I266851);
nor I_15529 (I266933,I266916,I266684);
nor I_15530 (I266598,I266752,I266933);
nor I_15531 (I266613,I266851,I266701);
nand I_15532 (I266978,I266834,I266817);
and I_15533 (I266995,I266978,I338310);
nand I_15534 (I267012,I266995,I338307);
not I_15535 (I267029,I267012);
nor I_15536 (I267046,I267029,I338319);
nand I_15537 (I267063,I266800,I267012);
not I_15538 (I266604,I267063);
nor I_15539 (I267094,I338316,I338301);
or I_15540 (I267111,I267094,I338313);
nor I_15541 (I267128,I338307,I338316);
nand I_15542 (I267145,I267128,I267111);
not I_15543 (I267162,I267145);
nor I_15544 (I266625,I267162,I266718);
nand I_15545 (I267193,I267162,I267046);
nand I_15546 (I266601,I267063,I267193);
nor I_15547 (I267224,I267162,I266735);
nor I_15548 (I266622,I267224,I266752);
nor I_15549 (I266616,I267162,I266916);
nor I_15550 (I267269,I267145,I266701);
nor I_15551 (I267286,I267029,I267269);
nor I_15552 (I266607,I267286,I266885);
nor I_15553 (I267317,I266718,I267145);
nor I_15554 (I267334,I267012,I267317);
DFFARX1 I_15555 (I267334,I2898,I266633,I266619,);
not I_15556 (I267398,I2905);
or I_15557 (I267415,I370485,I370500);
nor I_15558 (I267432,I370485,I370500);
nor I_15559 (I267449,I267432,I370509);
not I_15560 (I267466,I267449);
nand I_15561 (I267483,I267415,I370497);
not I_15562 (I267500,I267483);
not I_15563 (I267517,I370494);
nor I_15564 (I267360,I267517,I267500);
nor I_15565 (I267548,I267517,I267483);
nor I_15566 (I267565,I267449,I370494);
not I_15567 (I267582,I370488);
nand I_15568 (I267599,I370485,I370506);
nand I_15569 (I267616,I267599,I370488);
nor I_15570 (I267633,I267483,I267616);
not I_15571 (I267650,I267633);
nor I_15572 (I267375,I267616,I267548);
not I_15573 (I267681,I267616);
nor I_15574 (I267698,I267681,I267449);
nor I_15575 (I267363,I267517,I267698);
nor I_15576 (I267378,I267616,I267466);
nand I_15577 (I267743,I267599,I267582);
and I_15578 (I267760,I267743,I370512);
nand I_15579 (I267777,I267760,I370515);
not I_15580 (I267794,I267777);
nor I_15581 (I267811,I267794,I370494);
nand I_15582 (I267828,I267565,I267777);
not I_15583 (I267369,I267828);
nor I_15584 (I267859,I370488,I370482);
or I_15585 (I267876,I267859,I370482);
nor I_15586 (I267893,I370491,I370503);
nand I_15587 (I267910,I267893,I267876);
not I_15588 (I267927,I267910);
nor I_15589 (I267390,I267927,I267483);
nand I_15590 (I267958,I267927,I267811);
nand I_15591 (I267366,I267828,I267958);
nor I_15592 (I267989,I267927,I267500);
nor I_15593 (I267387,I267989,I267517);
nor I_15594 (I267381,I267927,I267681);
nor I_15595 (I268034,I267910,I267466);
nor I_15596 (I268051,I267794,I268034);
nor I_15597 (I267372,I268051,I267650);
nor I_15598 (I268082,I267483,I267910);
nor I_15599 (I268099,I267777,I268082);
DFFARX1 I_15600 (I268099,I2898,I267398,I267384,);
not I_15601 (I268163,I2905);
or I_15602 (I268180,I176280,I176295);
nor I_15603 (I268197,I176280,I176295);
nor I_15604 (I268214,I268197,I176286);
not I_15605 (I268231,I268214);
nand I_15606 (I268248,I268180,I176289);
not I_15607 (I268265,I268248);
not I_15608 (I268282,I176274);
nor I_15609 (I268125,I268282,I268265);
nor I_15610 (I268313,I268282,I268248);
nor I_15611 (I268330,I268214,I176274);
not I_15612 (I268347,I176298);
nand I_15613 (I268364,I176277,I176283);
nand I_15614 (I268381,I268364,I176298);
nor I_15615 (I268398,I268248,I268381);
not I_15616 (I268415,I268398);
nor I_15617 (I268140,I268381,I268313);
not I_15618 (I268446,I268381);
nor I_15619 (I268463,I268446,I268214);
nor I_15620 (I268128,I268282,I268463);
nor I_15621 (I268143,I268381,I268231);
nand I_15622 (I268508,I268364,I268347);
and I_15623 (I268525,I268508,I176304);
nand I_15624 (I268542,I268525,I176280);
not I_15625 (I268559,I268542);
nor I_15626 (I268576,I268559,I176274);
nand I_15627 (I268593,I268330,I268542);
not I_15628 (I268134,I268593);
nor I_15629 (I268624,I176307,I176292);
or I_15630 (I268641,I268624,I176277);
nor I_15631 (I268658,I176274,I176301);
nand I_15632 (I268675,I268658,I268641);
not I_15633 (I268692,I268675);
nor I_15634 (I268155,I268692,I268248);
nand I_15635 (I268723,I268692,I268576);
nand I_15636 (I268131,I268593,I268723);
nor I_15637 (I268754,I268692,I268265);
nor I_15638 (I268152,I268754,I268282);
nor I_15639 (I268146,I268692,I268446);
nor I_15640 (I268799,I268675,I268231);
nor I_15641 (I268816,I268559,I268799);
nor I_15642 (I268137,I268816,I268415);
nor I_15643 (I268847,I268248,I268675);
nor I_15644 (I268864,I268542,I268847);
DFFARX1 I_15645 (I268864,I2898,I268163,I268149,);
not I_15646 (I268928,I2905);
or I_15647 (I268945,I410152,I410164);
nor I_15648 (I268962,I410152,I410164);
nor I_15649 (I268979,I268962,I410146);
not I_15650 (I268996,I268979);
nand I_15651 (I269013,I268945,I410158);
not I_15652 (I269030,I269013);
not I_15653 (I269047,I410152);
nor I_15654 (I268890,I269047,I269030);
nor I_15655 (I269078,I269047,I269013);
nor I_15656 (I269095,I268979,I410152);
not I_15657 (I269112,I410143);
nand I_15658 (I269129,I410161,I410155);
nand I_15659 (I269146,I269129,I410143);
nor I_15660 (I269163,I269013,I269146);
not I_15661 (I269180,I269163);
nor I_15662 (I268905,I269146,I269078);
not I_15663 (I269211,I269146);
nor I_15664 (I269228,I269211,I268979);
nor I_15665 (I268893,I269047,I269228);
nor I_15666 (I268908,I269146,I268996);
nand I_15667 (I269273,I269129,I269112);
and I_15668 (I269290,I269273,I410167);
nand I_15669 (I269307,I269290,I410158);
not I_15670 (I269324,I269307);
nor I_15671 (I269341,I269324,I410152);
nand I_15672 (I269358,I269095,I269307);
not I_15673 (I268899,I269358);
nor I_15674 (I269389,I410155,I410146);
or I_15675 (I269406,I269389,I410143);
nor I_15676 (I269423,I410149,I410149);
nand I_15677 (I269440,I269423,I269406);
not I_15678 (I269457,I269440);
nor I_15679 (I268920,I269457,I269013);
nand I_15680 (I269488,I269457,I269341);
nand I_15681 (I268896,I269358,I269488);
nor I_15682 (I269519,I269457,I269030);
nor I_15683 (I268917,I269519,I269047);
nor I_15684 (I268911,I269457,I269211);
nor I_15685 (I269564,I269440,I268996);
nor I_15686 (I269581,I269324,I269564);
nor I_15687 (I268902,I269581,I269180);
nor I_15688 (I269612,I269013,I269440);
nor I_15689 (I269629,I269307,I269612);
DFFARX1 I_15690 (I269629,I2898,I268928,I268914,);
not I_15691 (I269693,I2905);
or I_15692 (I269710,I344849,I344846);
nor I_15693 (I269727,I344849,I344846);
nor I_15694 (I269744,I269727,I344855);
not I_15695 (I269761,I269744);
nand I_15696 (I269778,I269710,I344867);
not I_15697 (I269795,I269778);
not I_15698 (I269812,I344864);
nor I_15699 (I269655,I269812,I269795);
nor I_15700 (I269843,I269812,I269778);
nor I_15701 (I269860,I269744,I344864);
not I_15702 (I269877,I344870);
nand I_15703 (I269894,I344849,I344858);
nand I_15704 (I269911,I269894,I344870);
nor I_15705 (I269928,I269778,I269911);
not I_15706 (I269945,I269928);
nor I_15707 (I269670,I269911,I269843);
not I_15708 (I269976,I269911);
nor I_15709 (I269993,I269976,I269744);
nor I_15710 (I269658,I269812,I269993);
nor I_15711 (I269673,I269911,I269761);
nand I_15712 (I270038,I269894,I269877);
and I_15713 (I270055,I270038,I344855);
nand I_15714 (I270072,I270055,I344852);
not I_15715 (I270089,I270072);
nor I_15716 (I270106,I270089,I344864);
nand I_15717 (I270123,I269860,I270072);
not I_15718 (I269664,I270123);
nor I_15719 (I270154,I344861,I344846);
or I_15720 (I270171,I270154,I344858);
nor I_15721 (I270188,I344852,I344861);
nand I_15722 (I270205,I270188,I270171);
not I_15723 (I270222,I270205);
nor I_15724 (I269685,I270222,I269778);
nand I_15725 (I270253,I270222,I270106);
nand I_15726 (I269661,I270123,I270253);
nor I_15727 (I270284,I270222,I269795);
nor I_15728 (I269682,I270284,I269812);
nor I_15729 (I269676,I270222,I269976);
nor I_15730 (I270329,I270205,I269761);
nor I_15731 (I270346,I270089,I270329);
nor I_15732 (I269667,I270346,I269945);
nor I_15733 (I270377,I269778,I270205);
nor I_15734 (I270394,I270072,I270377);
DFFARX1 I_15735 (I270394,I2898,I269693,I269679,);
not I_15736 (I270458,I2905);
or I_15737 (I270475,I139306,I139303);
nor I_15738 (I270492,I139306,I139303);
nor I_15739 (I270509,I270492,I139288);
not I_15740 (I270526,I270509);
nand I_15741 (I270543,I270475,I139309);
not I_15742 (I270560,I270543);
not I_15743 (I270577,I139291);
nor I_15744 (I270420,I270577,I270560);
nor I_15745 (I270608,I270577,I270543);
nor I_15746 (I270625,I270509,I139291);
not I_15747 (I270642,I139285);
nand I_15748 (I270659,I139294,I139282);
nand I_15749 (I270676,I270659,I139285);
nor I_15750 (I270693,I270543,I270676);
not I_15751 (I270710,I270693);
nor I_15752 (I270435,I270676,I270608);
not I_15753 (I270741,I270676);
nor I_15754 (I270758,I270741,I270509);
nor I_15755 (I270423,I270577,I270758);
nor I_15756 (I270438,I270676,I270526);
nand I_15757 (I270803,I270659,I270642);
and I_15758 (I270820,I270803,I139315);
nand I_15759 (I270837,I270820,I139312);
not I_15760 (I270854,I270837);
nor I_15761 (I270871,I270854,I139291);
nand I_15762 (I270888,I270625,I270837);
not I_15763 (I270429,I270888);
nor I_15764 (I270919,I139282,I139300);
or I_15765 (I270936,I270919,I139285);
nor I_15766 (I270953,I139297,I139288);
nand I_15767 (I270970,I270953,I270936);
not I_15768 (I270987,I270970);
nor I_15769 (I270450,I270987,I270543);
nand I_15770 (I271018,I270987,I270871);
nand I_15771 (I270426,I270888,I271018);
nor I_15772 (I271049,I270987,I270560);
nor I_15773 (I270447,I271049,I270577);
nor I_15774 (I270441,I270987,I270741);
nor I_15775 (I271094,I270970,I270526);
nor I_15776 (I271111,I270854,I271094);
nor I_15777 (I270432,I271111,I270710);
nor I_15778 (I271142,I270543,I270970);
nor I_15779 (I271159,I270837,I271142);
DFFARX1 I_15780 (I271159,I2898,I270458,I270444,);
not I_15781 (I271223,I2905);
or I_15782 (I271240,I222424,I222418);
nor I_15783 (I271257,I222424,I222418);
nor I_15784 (I271274,I271257,I222433);
not I_15785 (I271291,I271274);
nand I_15786 (I271308,I271240,I222436);
not I_15787 (I271325,I271308);
not I_15788 (I271342,I222418);
nor I_15789 (I271185,I271342,I271325);
nor I_15790 (I271373,I271342,I271308);
nor I_15791 (I271390,I271274,I222418);
not I_15792 (I271407,I222421);
nand I_15793 (I271424,I222439,I222412);
nand I_15794 (I271441,I271424,I222421);
nor I_15795 (I271458,I271308,I271441);
not I_15796 (I271475,I271458);
nor I_15797 (I271200,I271441,I271373);
not I_15798 (I271506,I271441);
nor I_15799 (I271523,I271506,I271274);
nor I_15800 (I271188,I271342,I271523);
nor I_15801 (I271203,I271441,I271291);
nand I_15802 (I271568,I271424,I271407);
and I_15803 (I271585,I271568,I222424);
nand I_15804 (I271602,I271585,I222415);
not I_15805 (I271619,I271602);
nor I_15806 (I271636,I271619,I222418);
nand I_15807 (I271653,I271390,I271602);
not I_15808 (I271194,I271653);
nor I_15809 (I271684,I222415,I222421);
or I_15810 (I271701,I271684,I222412);
nor I_15811 (I271718,I222427,I222430);
nand I_15812 (I271735,I271718,I271701);
not I_15813 (I271752,I271735);
nor I_15814 (I271215,I271752,I271308);
nand I_15815 (I271783,I271752,I271636);
nand I_15816 (I271191,I271653,I271783);
nor I_15817 (I271814,I271752,I271325);
nor I_15818 (I271212,I271814,I271342);
nor I_15819 (I271206,I271752,I271506);
nor I_15820 (I271859,I271735,I271291);
nor I_15821 (I271876,I271619,I271859);
nor I_15822 (I271197,I271876,I271475);
nor I_15823 (I271907,I271308,I271735);
nor I_15824 (I271924,I271602,I271907);
DFFARX1 I_15825 (I271924,I2898,I271223,I271209,);
not I_15826 (I271988,I2905);
or I_15827 (I272005,I344254,I344251);
nor I_15828 (I272022,I344254,I344251);
nor I_15829 (I272039,I272022,I344260);
not I_15830 (I272056,I272039);
nand I_15831 (I272073,I272005,I344272);
not I_15832 (I272090,I272073);
not I_15833 (I272107,I344269);
nor I_15834 (I271950,I272107,I272090);
nor I_15835 (I272138,I272107,I272073);
nor I_15836 (I272155,I272039,I344269);
not I_15837 (I272172,I344275);
nand I_15838 (I272189,I344254,I344263);
nand I_15839 (I272206,I272189,I344275);
nor I_15840 (I272223,I272073,I272206);
not I_15841 (I272240,I272223);
nor I_15842 (I271965,I272206,I272138);
not I_15843 (I272271,I272206);
nor I_15844 (I272288,I272271,I272039);
nor I_15845 (I271953,I272107,I272288);
nor I_15846 (I271968,I272206,I272056);
nand I_15847 (I272333,I272189,I272172);
and I_15848 (I272350,I272333,I344260);
nand I_15849 (I272367,I272350,I344257);
not I_15850 (I272384,I272367);
nor I_15851 (I272401,I272384,I344269);
nand I_15852 (I272418,I272155,I272367);
not I_15853 (I271959,I272418);
nor I_15854 (I272449,I344266,I344251);
or I_15855 (I272466,I272449,I344263);
nor I_15856 (I272483,I344257,I344266);
nand I_15857 (I272500,I272483,I272466);
not I_15858 (I272517,I272500);
nor I_15859 (I271980,I272517,I272073);
nand I_15860 (I272548,I272517,I272401);
nand I_15861 (I271956,I272418,I272548);
nor I_15862 (I272579,I272517,I272090);
nor I_15863 (I271977,I272579,I272107);
nor I_15864 (I271971,I272517,I272271);
nor I_15865 (I272624,I272500,I272056);
nor I_15866 (I272641,I272384,I272624);
nor I_15867 (I271962,I272641,I272240);
nor I_15868 (I272672,I272073,I272500);
nor I_15869 (I272689,I272367,I272672);
DFFARX1 I_15870 (I272689,I2898,I271988,I271974,);
not I_15871 (I272753,I2905);
or I_15872 (I272770,I207464,I207458);
nor I_15873 (I272787,I207464,I207458);
nor I_15874 (I272804,I272787,I207473);
not I_15875 (I272821,I272804);
nand I_15876 (I272838,I272770,I207476);
not I_15877 (I272855,I272838);
not I_15878 (I272872,I207458);
nor I_15879 (I272715,I272872,I272855);
nor I_15880 (I272903,I272872,I272838);
nor I_15881 (I272920,I272804,I207458);
not I_15882 (I272937,I207461);
nand I_15883 (I272954,I207479,I207452);
nand I_15884 (I272971,I272954,I207461);
nor I_15885 (I272988,I272838,I272971);
not I_15886 (I273005,I272988);
nor I_15887 (I272730,I272971,I272903);
not I_15888 (I273036,I272971);
nor I_15889 (I273053,I273036,I272804);
nor I_15890 (I272718,I272872,I273053);
nor I_15891 (I272733,I272971,I272821);
nand I_15892 (I273098,I272954,I272937);
and I_15893 (I273115,I273098,I207464);
nand I_15894 (I273132,I273115,I207455);
not I_15895 (I273149,I273132);
nor I_15896 (I273166,I273149,I207458);
nand I_15897 (I273183,I272920,I273132);
not I_15898 (I272724,I273183);
nor I_15899 (I273214,I207455,I207461);
or I_15900 (I273231,I273214,I207452);
nor I_15901 (I273248,I207467,I207470);
nand I_15902 (I273265,I273248,I273231);
not I_15903 (I273282,I273265);
nor I_15904 (I272745,I273282,I272838);
nand I_15905 (I273313,I273282,I273166);
nand I_15906 (I272721,I273183,I273313);
nor I_15907 (I273344,I273282,I272855);
nor I_15908 (I272742,I273344,I272872);
nor I_15909 (I272736,I273282,I273036);
nor I_15910 (I273389,I273265,I272821);
nor I_15911 (I273406,I273149,I273389);
nor I_15912 (I272727,I273406,I273005);
nor I_15913 (I273437,I272838,I273265);
nor I_15914 (I273454,I273132,I273437);
DFFARX1 I_15915 (I273454,I2898,I272753,I272739,);
not I_15916 (I273518,I2905);
or I_15917 (I273535,I420605,I420602);
nor I_15918 (I273552,I420605,I420602);
nor I_15919 (I273569,I273552,I420590);
not I_15920 (I273586,I273569);
nand I_15921 (I273603,I273535,I420611);
not I_15922 (I273620,I273603);
not I_15923 (I273637,I420581);
nor I_15924 (I273480,I273637,I273620);
nor I_15925 (I273668,I273637,I273603);
nor I_15926 (I273685,I273569,I420581);
not I_15927 (I273702,I420599);
nand I_15928 (I273719,I420614,I420596);
nand I_15929 (I273736,I273719,I420599);
nor I_15930 (I273753,I273603,I273736);
not I_15931 (I273770,I273753);
nor I_15932 (I273495,I273736,I273668);
not I_15933 (I273801,I273736);
nor I_15934 (I273818,I273801,I273569);
nor I_15935 (I273483,I273637,I273818);
nor I_15936 (I273498,I273736,I273586);
nand I_15937 (I273863,I273719,I273702);
and I_15938 (I273880,I273863,I420608);
nand I_15939 (I273897,I273880,I420587);
not I_15940 (I273914,I273897);
nor I_15941 (I273931,I273914,I420581);
nand I_15942 (I273948,I273685,I273897);
not I_15943 (I273489,I273948);
nor I_15944 (I273979,I420593,I420581);
or I_15945 (I273996,I273979,I420584);
nor I_15946 (I274013,I420584,I420587);
nand I_15947 (I274030,I274013,I273996);
not I_15948 (I274047,I274030);
nor I_15949 (I273510,I274047,I273603);
nand I_15950 (I274078,I274047,I273931);
nand I_15951 (I273486,I273948,I274078);
nor I_15952 (I274109,I274047,I273620);
nor I_15953 (I273507,I274109,I273637);
nor I_15954 (I273501,I274047,I273801);
nor I_15955 (I274154,I274030,I273586);
nor I_15956 (I274171,I273914,I274154);
nor I_15957 (I273492,I274171,I273770);
nor I_15958 (I274202,I273603,I274030);
nor I_15959 (I274219,I273897,I274202);
DFFARX1 I_15960 (I274219,I2898,I273518,I273504,);
not I_15961 (I274283,I2905);
or I_15962 (I274300,I293727,I293745);
nor I_15963 (I274317,I293727,I293745);
nor I_15964 (I274334,I274317,I293730);
not I_15965 (I274351,I274334);
nand I_15966 (I274368,I274300,I293739);
not I_15967 (I274385,I274368);
not I_15968 (I274402,I293751);
nor I_15969 (I274245,I274402,I274385);
nor I_15970 (I274433,I274402,I274368);
nor I_15971 (I274450,I274334,I293751);
not I_15972 (I274467,I293748);
nand I_15973 (I274484,I293754,I293727);
nand I_15974 (I274501,I274484,I293748);
nor I_15975 (I274518,I274368,I274501);
not I_15976 (I274535,I274518);
nor I_15977 (I274260,I274501,I274433);
not I_15978 (I274566,I274501);
nor I_15979 (I274583,I274566,I274334);
nor I_15980 (I274248,I274402,I274583);
nor I_15981 (I274263,I274501,I274351);
nand I_15982 (I274628,I274484,I274467);
and I_15983 (I274645,I274628,I293733);
nand I_15984 (I274662,I274645,I293736);
not I_15985 (I274679,I274662);
nor I_15986 (I274696,I274679,I293751);
nand I_15987 (I274713,I274450,I274662);
not I_15988 (I274254,I274713);
nor I_15989 (I274744,I293736,I293757);
or I_15990 (I274761,I274744,I293733);
nor I_15991 (I274778,I293742,I293730);
nand I_15992 (I274795,I274778,I274761);
not I_15993 (I274812,I274795);
nor I_15994 (I274275,I274812,I274368);
nand I_15995 (I274843,I274812,I274696);
nand I_15996 (I274251,I274713,I274843);
nor I_15997 (I274874,I274812,I274385);
nor I_15998 (I274272,I274874,I274402);
nor I_15999 (I274266,I274812,I274566);
nor I_16000 (I274919,I274795,I274351);
nor I_16001 (I274936,I274679,I274919);
nor I_16002 (I274257,I274936,I274535);
nor I_16003 (I274967,I274368,I274795);
nor I_16004 (I274984,I274662,I274967);
DFFARX1 I_16005 (I274984,I2898,I274283,I274269,);
not I_16006 (I275048,I2905);
or I_16007 (I275065,I107856,I107853);
nor I_16008 (I275082,I107856,I107853);
nor I_16009 (I275099,I275082,I107838);
not I_16010 (I275116,I275099);
nand I_16011 (I275133,I275065,I107859);
not I_16012 (I275150,I275133);
not I_16013 (I275167,I107841);
nor I_16014 (I275010,I275167,I275150);
nor I_16015 (I275198,I275167,I275133);
nor I_16016 (I275215,I275099,I107841);
not I_16017 (I275232,I107835);
nand I_16018 (I275249,I107844,I107832);
nand I_16019 (I275266,I275249,I107835);
nor I_16020 (I275283,I275133,I275266);
not I_16021 (I275300,I275283);
nor I_16022 (I275025,I275266,I275198);
not I_16023 (I275331,I275266);
nor I_16024 (I275348,I275331,I275099);
nor I_16025 (I275013,I275167,I275348);
nor I_16026 (I275028,I275266,I275116);
nand I_16027 (I275393,I275249,I275232);
and I_16028 (I275410,I275393,I107865);
nand I_16029 (I275427,I275410,I107862);
not I_16030 (I275444,I275427);
nor I_16031 (I275461,I275444,I107841);
nand I_16032 (I275478,I275215,I275427);
not I_16033 (I275019,I275478);
nor I_16034 (I275509,I107832,I107850);
or I_16035 (I275526,I275509,I107835);
nor I_16036 (I275543,I107847,I107838);
nand I_16037 (I275560,I275543,I275526);
not I_16038 (I275577,I275560);
nor I_16039 (I275040,I275577,I275133);
nand I_16040 (I275608,I275577,I275461);
nand I_16041 (I275016,I275478,I275608);
nor I_16042 (I275639,I275577,I275150);
nor I_16043 (I275037,I275639,I275167);
nor I_16044 (I275031,I275577,I275331);
nor I_16045 (I275684,I275560,I275116);
nor I_16046 (I275701,I275444,I275684);
nor I_16047 (I275022,I275701,I275300);
nor I_16048 (I275732,I275133,I275560);
nor I_16049 (I275749,I275427,I275732);
DFFARX1 I_16050 (I275749,I2898,I275048,I275034,);
not I_16051 (I275813,I2905);
or I_16052 (I275830,I82735,I82747);
nor I_16053 (I275847,I82735,I82747);
nor I_16054 (I275864,I275847,I82744);
not I_16055 (I275881,I275864);
nand I_16056 (I275898,I275830,I82738);
not I_16057 (I275915,I275898);
not I_16058 (I275932,I82732);
nor I_16059 (I275775,I275932,I275915);
nor I_16060 (I275963,I275932,I275898);
nor I_16061 (I275980,I275864,I82732);
not I_16062 (I275997,I82741);
nand I_16063 (I276014,I82729,I82726);
nand I_16064 (I276031,I276014,I82741);
nor I_16065 (I276048,I275898,I276031);
not I_16066 (I276065,I276048);
nor I_16067 (I275790,I276031,I275963);
not I_16068 (I276096,I276031);
nor I_16069 (I276113,I276096,I275864);
nor I_16070 (I275778,I275932,I276113);
nor I_16071 (I275793,I276031,I275881);
nand I_16072 (I276158,I276014,I275997);
and I_16073 (I276175,I276158,I82735);
nand I_16074 (I276192,I276175,I82723);
not I_16075 (I276209,I276192);
nor I_16076 (I276226,I276209,I82732);
nand I_16077 (I276243,I275980,I276192);
not I_16078 (I275784,I276243);
nor I_16079 (I276274,I82729,I82726);
or I_16080 (I276291,I276274,I82732);
nor I_16081 (I276308,I82723,I82750);
nand I_16082 (I276325,I276308,I276291);
not I_16083 (I276342,I276325);
nor I_16084 (I275805,I276342,I275898);
nand I_16085 (I276373,I276342,I276226);
nand I_16086 (I275781,I276243,I276373);
nor I_16087 (I276404,I276342,I275915);
nor I_16088 (I275802,I276404,I275932);
nor I_16089 (I275796,I276342,I276096);
nor I_16090 (I276449,I276325,I275881);
nor I_16091 (I276466,I276209,I276449);
nor I_16092 (I275787,I276466,I276065);
nor I_16093 (I276497,I275898,I276325);
nor I_16094 (I276514,I276192,I276497);
DFFARX1 I_16095 (I276514,I2898,I275813,I275799,);
not I_16096 (I276578,I2905);
or I_16097 (I276595,I166080,I166095);
nor I_16098 (I276612,I166080,I166095);
nor I_16099 (I276629,I276612,I166086);
not I_16100 (I276646,I276629);
nand I_16101 (I276663,I276595,I166089);
not I_16102 (I276680,I276663);
not I_16103 (I276697,I166074);
nor I_16104 (I276540,I276697,I276680);
nor I_16105 (I276728,I276697,I276663);
nor I_16106 (I276745,I276629,I166074);
not I_16107 (I276762,I166098);
nand I_16108 (I276779,I166077,I166083);
nand I_16109 (I276796,I276779,I166098);
nor I_16110 (I276813,I276663,I276796);
not I_16111 (I276830,I276813);
nor I_16112 (I276555,I276796,I276728);
not I_16113 (I276861,I276796);
nor I_16114 (I276878,I276861,I276629);
nor I_16115 (I276543,I276697,I276878);
nor I_16116 (I276558,I276796,I276646);
nand I_16117 (I276923,I276779,I276762);
and I_16118 (I276940,I276923,I166104);
nand I_16119 (I276957,I276940,I166080);
not I_16120 (I276974,I276957);
nor I_16121 (I276991,I276974,I166074);
nand I_16122 (I277008,I276745,I276957);
not I_16123 (I276549,I277008);
nor I_16124 (I277039,I166107,I166092);
or I_16125 (I277056,I277039,I166077);
nor I_16126 (I277073,I166074,I166101);
nand I_16127 (I277090,I277073,I277056);
not I_16128 (I277107,I277090);
nor I_16129 (I276570,I277107,I276663);
nand I_16130 (I277138,I277107,I276991);
nand I_16131 (I276546,I277008,I277138);
nor I_16132 (I277169,I277107,I276680);
nor I_16133 (I276567,I277169,I276697);
nor I_16134 (I276561,I277107,I276861);
nor I_16135 (I277214,I277090,I276646);
nor I_16136 (I277231,I276974,I277214);
nor I_16137 (I276552,I277231,I276830);
nor I_16138 (I277262,I276663,I277090);
nor I_16139 (I277279,I276957,I277262);
DFFARX1 I_16140 (I277279,I2898,I276578,I276564,);
not I_16141 (I277343,I2905);
or I_16142 (I277360,I191115,I191115);
nor I_16143 (I277377,I191115,I191115);
nor I_16144 (I277394,I277377,I191130);
not I_16145 (I277411,I277394);
nand I_16146 (I277428,I277360,I191127);
not I_16147 (I277445,I277428);
not I_16148 (I277462,I191139);
nor I_16149 (I277305,I277462,I277445);
nor I_16150 (I277493,I277462,I277428);
nor I_16151 (I277510,I277394,I191139);
not I_16152 (I277527,I191118);
nand I_16153 (I277544,I191130,I191121);
nand I_16154 (I277561,I277544,I191118);
nor I_16155 (I277578,I277428,I277561);
not I_16156 (I277595,I277578);
nor I_16157 (I277320,I277561,I277493);
not I_16158 (I277626,I277561);
nor I_16159 (I277643,I277626,I277394);
nor I_16160 (I277308,I277462,I277643);
nor I_16161 (I277323,I277561,I277411);
nand I_16162 (I277688,I277544,I277527);
and I_16163 (I277705,I277688,I191127);
nand I_16164 (I277722,I277705,I191121);
not I_16165 (I277739,I277722);
nor I_16166 (I277756,I277739,I191139);
nand I_16167 (I277773,I277510,I277722);
not I_16168 (I277314,I277773);
nor I_16169 (I277804,I191124,I191124);
or I_16170 (I277821,I277804,I191118);
nor I_16171 (I277838,I191133,I191136);
nand I_16172 (I277855,I277838,I277821);
not I_16173 (I277872,I277855);
nor I_16174 (I277335,I277872,I277428);
nand I_16175 (I277903,I277872,I277756);
nand I_16176 (I277311,I277773,I277903);
nor I_16177 (I277934,I277872,I277445);
nor I_16178 (I277332,I277934,I277462);
nor I_16179 (I277326,I277872,I277626);
nor I_16180 (I277979,I277855,I277411);
nor I_16181 (I277996,I277739,I277979);
nor I_16182 (I277317,I277996,I277595);
nor I_16183 (I278027,I277428,I277855);
nor I_16184 (I278044,I277722,I278027);
DFFARX1 I_16185 (I278044,I2898,I277343,I277329,);
not I_16186 (I278108,I2905);
or I_16187 (I278125,I80219,I80231);
nor I_16188 (I278142,I80219,I80231);
nor I_16189 (I278159,I278142,I80228);
not I_16190 (I278176,I278159);
nand I_16191 (I278193,I278125,I80222);
not I_16192 (I278210,I278193);
not I_16193 (I278227,I80216);
nor I_16194 (I278070,I278227,I278210);
nor I_16195 (I278258,I278227,I278193);
nor I_16196 (I278275,I278159,I80216);
not I_16197 (I278292,I80225);
nand I_16198 (I278309,I80213,I80210);
nand I_16199 (I278326,I278309,I80225);
nor I_16200 (I278343,I278193,I278326);
not I_16201 (I278360,I278343);
nor I_16202 (I278085,I278326,I278258);
not I_16203 (I278391,I278326);
nor I_16204 (I278408,I278391,I278159);
nor I_16205 (I278073,I278227,I278408);
nor I_16206 (I278088,I278326,I278176);
nand I_16207 (I278453,I278309,I278292);
and I_16208 (I278470,I278453,I80219);
nand I_16209 (I278487,I278470,I80207);
not I_16210 (I278504,I278487);
nor I_16211 (I278521,I278504,I80216);
nand I_16212 (I278538,I278275,I278487);
not I_16213 (I278079,I278538);
nor I_16214 (I278569,I80213,I80210);
or I_16215 (I278586,I278569,I80216);
nor I_16216 (I278603,I80207,I80234);
nand I_16217 (I278620,I278603,I278586);
not I_16218 (I278637,I278620);
nor I_16219 (I278100,I278637,I278193);
nand I_16220 (I278668,I278637,I278521);
nand I_16221 (I278076,I278538,I278668);
nor I_16222 (I278699,I278637,I278210);
nor I_16223 (I278097,I278699,I278227);
nor I_16224 (I278091,I278637,I278391);
nor I_16225 (I278744,I278620,I278176);
nor I_16226 (I278761,I278504,I278744);
nor I_16227 (I278082,I278761,I278360);
nor I_16228 (I278792,I278193,I278620);
nor I_16229 (I278809,I278487,I278792);
DFFARX1 I_16230 (I278809,I2898,I278108,I278094,);
not I_16231 (I278873,I2905);
or I_16232 (I278890,I307616,I307634);
nor I_16233 (I278907,I307616,I307634);
nor I_16234 (I278924,I278907,I307619);
not I_16235 (I278941,I278924);
nand I_16236 (I278958,I278890,I307628);
not I_16237 (I278975,I278958);
not I_16238 (I278992,I307640);
nor I_16239 (I278835,I278992,I278975);
nor I_16240 (I279023,I278992,I278958);
nor I_16241 (I279040,I278924,I307640);
not I_16242 (I279057,I307637);
nand I_16243 (I279074,I307643,I307616);
nand I_16244 (I279091,I279074,I307637);
nor I_16245 (I279108,I278958,I279091);
not I_16246 (I279125,I279108);
nor I_16247 (I278850,I279091,I279023);
not I_16248 (I279156,I279091);
nor I_16249 (I279173,I279156,I278924);
nor I_16250 (I278838,I278992,I279173);
nor I_16251 (I278853,I279091,I278941);
nand I_16252 (I279218,I279074,I279057);
and I_16253 (I279235,I279218,I307622);
nand I_16254 (I279252,I279235,I307625);
not I_16255 (I279269,I279252);
nor I_16256 (I279286,I279269,I307640);
nand I_16257 (I279303,I279040,I279252);
not I_16258 (I278844,I279303);
nor I_16259 (I279334,I307625,I307646);
or I_16260 (I279351,I279334,I307622);
nor I_16261 (I279368,I307631,I307619);
nand I_16262 (I279385,I279368,I279351);
not I_16263 (I279402,I279385);
nor I_16264 (I278865,I279402,I278958);
nand I_16265 (I279433,I279402,I279286);
nand I_16266 (I278841,I279303,I279433);
nor I_16267 (I279464,I279402,I278975);
nor I_16268 (I278862,I279464,I278992);
nor I_16269 (I278856,I279402,I279156);
nor I_16270 (I279509,I279385,I278941);
nor I_16271 (I279526,I279269,I279509);
nor I_16272 (I278847,I279526,I279125);
nor I_16273 (I279557,I278958,I279385);
nor I_16274 (I279574,I279252,I279557);
DFFARX1 I_16275 (I279574,I2898,I278873,I278859,);
not I_16276 (I279638,I2905);
or I_16277 (I279655,I315657,I315675);
nor I_16278 (I279672,I315657,I315675);
nor I_16279 (I279689,I279672,I315660);
not I_16280 (I279706,I279689);
nand I_16281 (I279723,I279655,I315669);
not I_16282 (I279740,I279723);
not I_16283 (I279757,I315681);
nor I_16284 (I279600,I279757,I279740);
nor I_16285 (I279788,I279757,I279723);
nor I_16286 (I279805,I279689,I315681);
not I_16287 (I279822,I315678);
nand I_16288 (I279839,I315684,I315657);
nand I_16289 (I279856,I279839,I315678);
nor I_16290 (I279873,I279723,I279856);
not I_16291 (I279890,I279873);
nor I_16292 (I279615,I279856,I279788);
not I_16293 (I279921,I279856);
nor I_16294 (I279938,I279921,I279689);
nor I_16295 (I279603,I279757,I279938);
nor I_16296 (I279618,I279856,I279706);
nand I_16297 (I279983,I279839,I279822);
and I_16298 (I280000,I279983,I315663);
nand I_16299 (I280017,I280000,I315666);
not I_16300 (I280034,I280017);
nor I_16301 (I280051,I280034,I315681);
nand I_16302 (I280068,I279805,I280017);
not I_16303 (I279609,I280068);
nor I_16304 (I280099,I315666,I315687);
or I_16305 (I280116,I280099,I315663);
nor I_16306 (I280133,I315672,I315660);
nand I_16307 (I280150,I280133,I280116);
not I_16308 (I280167,I280150);
nor I_16309 (I279630,I280167,I279723);
nand I_16310 (I280198,I280167,I280051);
nand I_16311 (I279606,I280068,I280198);
nor I_16312 (I280229,I280167,I279740);
nor I_16313 (I279627,I280229,I279757);
nor I_16314 (I279621,I280167,I279921);
nor I_16315 (I280274,I280150,I279706);
nor I_16316 (I280291,I280034,I280274);
nor I_16317 (I279612,I280291,I279890);
nor I_16318 (I280322,I279723,I280150);
nor I_16319 (I280339,I280017,I280322);
DFFARX1 I_16320 (I280339,I2898,I279638,I279624,);
not I_16321 (I280403,I2905);
or I_16322 (I280420,I349014,I349011);
nor I_16323 (I280437,I349014,I349011);
nor I_16324 (I280454,I280437,I349020);
not I_16325 (I280471,I280454);
nand I_16326 (I280488,I280420,I349032);
not I_16327 (I280505,I280488);
not I_16328 (I280522,I349029);
nor I_16329 (I280365,I280522,I280505);
nor I_16330 (I280553,I280522,I280488);
nor I_16331 (I280570,I280454,I349029);
not I_16332 (I280587,I349035);
nand I_16333 (I280604,I349014,I349023);
nand I_16334 (I280621,I280604,I349035);
nor I_16335 (I280638,I280488,I280621);
not I_16336 (I280655,I280638);
nor I_16337 (I280380,I280621,I280553);
not I_16338 (I280686,I280621);
nor I_16339 (I280703,I280686,I280454);
nor I_16340 (I280368,I280522,I280703);
nor I_16341 (I280383,I280621,I280471);
nand I_16342 (I280748,I280604,I280587);
and I_16343 (I280765,I280748,I349020);
nand I_16344 (I280782,I280765,I349017);
not I_16345 (I280799,I280782);
nor I_16346 (I280816,I280799,I349029);
nand I_16347 (I280833,I280570,I280782);
not I_16348 (I280374,I280833);
nor I_16349 (I280864,I349026,I349011);
or I_16350 (I280881,I280864,I349023);
nor I_16351 (I280898,I349017,I349026);
nand I_16352 (I280915,I280898,I280881);
not I_16353 (I280932,I280915);
nor I_16354 (I280395,I280932,I280488);
nand I_16355 (I280963,I280932,I280816);
nand I_16356 (I280371,I280833,I280963);
nor I_16357 (I280994,I280932,I280505);
nor I_16358 (I280392,I280994,I280522);
nor I_16359 (I280386,I280932,I280686);
nor I_16360 (I281039,I280915,I280471);
nor I_16361 (I281056,I280799,I281039);
nor I_16362 (I280377,I281056,I280655);
nor I_16363 (I281087,I280488,I280915);
nor I_16364 (I281104,I280782,I281087);
DFFARX1 I_16365 (I281104,I2898,I280403,I280389,);
not I_16366 (I281168,I2905);
or I_16367 (I281185,I422696,I422693);
nor I_16368 (I281202,I422696,I422693);
nor I_16369 (I281219,I281202,I422681);
not I_16370 (I281236,I281219);
nand I_16371 (I281253,I281185,I422702);
not I_16372 (I281270,I281253);
not I_16373 (I281287,I422672);
nor I_16374 (I281130,I281287,I281270);
nor I_16375 (I281318,I281287,I281253);
nor I_16376 (I281335,I281219,I422672);
not I_16377 (I281352,I422690);
nand I_16378 (I281369,I422705,I422687);
nand I_16379 (I281386,I281369,I422690);
nor I_16380 (I281403,I281253,I281386);
not I_16381 (I281420,I281403);
nor I_16382 (I281145,I281386,I281318);
not I_16383 (I281451,I281386);
nor I_16384 (I281468,I281451,I281219);
nor I_16385 (I281133,I281287,I281468);
nor I_16386 (I281148,I281386,I281236);
nand I_16387 (I281513,I281369,I281352);
and I_16388 (I281530,I281513,I422699);
nand I_16389 (I281547,I281530,I422678);
not I_16390 (I281564,I281547);
nor I_16391 (I281581,I281564,I422672);
nand I_16392 (I281598,I281335,I281547);
not I_16393 (I281139,I281598);
nor I_16394 (I281629,I422684,I422672);
or I_16395 (I281646,I281629,I422675);
nor I_16396 (I281663,I422675,I422678);
nand I_16397 (I281680,I281663,I281646);
not I_16398 (I281697,I281680);
nor I_16399 (I281160,I281697,I281253);
nand I_16400 (I281728,I281697,I281581);
nand I_16401 (I281136,I281598,I281728);
nor I_16402 (I281759,I281697,I281270);
nor I_16403 (I281157,I281759,I281287);
nor I_16404 (I281151,I281697,I281451);
nor I_16405 (I281804,I281680,I281236);
nor I_16406 (I281821,I281564,I281804);
nor I_16407 (I281142,I281821,I281420);
nor I_16408 (I281852,I281253,I281680);
nor I_16409 (I281869,I281547,I281852);
DFFARX1 I_16410 (I281869,I2898,I281168,I281154,);
not I_16411 (I281933,I2905);
or I_16412 (I281950,I41794,I41770);
nor I_16413 (I281967,I41794,I41770);
nor I_16414 (I281984,I281967,I41782);
not I_16415 (I282001,I281984);
nand I_16416 (I282018,I281950,I41779);
not I_16417 (I282035,I282018);
not I_16418 (I282052,I41776);
nor I_16419 (I281895,I282052,I282035);
nor I_16420 (I282083,I282052,I282018);
nor I_16421 (I282100,I281984,I41776);
not I_16422 (I282117,I41785);
nand I_16423 (I282134,I41803,I41770);
nand I_16424 (I282151,I282134,I41785);
nor I_16425 (I282168,I282018,I282151);
not I_16426 (I282185,I282168);
nor I_16427 (I281910,I282151,I282083);
not I_16428 (I282216,I282151);
nor I_16429 (I282233,I282216,I281984);
nor I_16430 (I281898,I282052,I282233);
nor I_16431 (I281913,I282151,I282001);
nand I_16432 (I282278,I282134,I282117);
and I_16433 (I282295,I282278,I41806);
nand I_16434 (I282312,I282295,I41797);
not I_16435 (I282329,I282312);
nor I_16436 (I282346,I282329,I41776);
nand I_16437 (I282363,I282100,I282312);
not I_16438 (I281904,I282363);
nor I_16439 (I282394,I41773,I41788);
or I_16440 (I282411,I282394,I41773);
nor I_16441 (I282428,I41791,I41800);
nand I_16442 (I282445,I282428,I282411);
not I_16443 (I282462,I282445);
nor I_16444 (I281925,I282462,I282018);
nand I_16445 (I282493,I282462,I282346);
nand I_16446 (I281901,I282363,I282493);
nor I_16447 (I282524,I282462,I282035);
nor I_16448 (I281922,I282524,I282052);
nor I_16449 (I281916,I282462,I282216);
nor I_16450 (I282569,I282445,I282001);
nor I_16451 (I282586,I282329,I282569);
nor I_16452 (I281907,I282586,I282185);
nor I_16453 (I282617,I282018,I282445);
nor I_16454 (I282634,I282312,I282617);
DFFARX1 I_16455 (I282634,I2898,I281933,I281919,);
not I_16456 (I282698,I2905);
or I_16457 (I282715,I34651,I34639);
nor I_16458 (I282732,I34651,I34639);
nor I_16459 (I282749,I282732,I34642);
not I_16460 (I282766,I282749);
nand I_16461 (I282783,I282715,I34630);
not I_16462 (I282800,I282783);
not I_16463 (I282817,I34654);
nor I_16464 (I282660,I282817,I282800);
nor I_16465 (I282848,I282817,I282783);
nor I_16466 (I282865,I282749,I34654);
not I_16467 (I282882,I34630);
nand I_16468 (I282899,I34645,I34636);
nand I_16469 (I282916,I282899,I34630);
nor I_16470 (I282933,I282783,I282916);
not I_16471 (I282950,I282933);
nor I_16472 (I282675,I282916,I282848);
not I_16473 (I282981,I282916);
nor I_16474 (I282998,I282981,I282749);
nor I_16475 (I282663,I282817,I282998);
nor I_16476 (I282678,I282916,I282766);
nand I_16477 (I283043,I282899,I282882);
and I_16478 (I283060,I283043,I34642);
nand I_16479 (I283077,I283060,I34633);
not I_16480 (I283094,I283077);
nor I_16481 (I283111,I283094,I34654);
nand I_16482 (I283128,I282865,I283077);
not I_16483 (I282669,I283128);
nor I_16484 (I283159,I34633,I34657);
or I_16485 (I283176,I283159,I34648);
nor I_16486 (I283193,I34639,I34636);
nand I_16487 (I283210,I283193,I283176);
not I_16488 (I283227,I283210);
nor I_16489 (I282690,I283227,I282783);
nand I_16490 (I283258,I283227,I283111);
nand I_16491 (I282666,I283128,I283258);
nor I_16492 (I283289,I283227,I282800);
nor I_16493 (I282687,I283289,I282817);
nor I_16494 (I282681,I283227,I282981);
nor I_16495 (I283334,I283210,I282766);
nor I_16496 (I283351,I283094,I283334);
nor I_16497 (I282672,I283351,I282950);
nor I_16498 (I283382,I282783,I283210);
nor I_16499 (I283399,I283077,I283382);
DFFARX1 I_16500 (I283399,I2898,I282698,I282684,);
not I_16501 (I283463,I2905);
or I_16502 (I283480,I424787,I424784);
nor I_16503 (I283497,I424787,I424784);
nor I_16504 (I283514,I283497,I424772);
not I_16505 (I283531,I283514);
nand I_16506 (I283548,I283480,I424793);
not I_16507 (I283565,I283548);
not I_16508 (I283582,I424763);
nor I_16509 (I283425,I283582,I283565);
nor I_16510 (I283613,I283582,I283548);
nor I_16511 (I283630,I283514,I424763);
not I_16512 (I283647,I424781);
nand I_16513 (I283664,I424796,I424778);
nand I_16514 (I283681,I283664,I424781);
nor I_16515 (I283698,I283548,I283681);
not I_16516 (I283715,I283698);
nor I_16517 (I283440,I283681,I283613);
not I_16518 (I283746,I283681);
nor I_16519 (I283763,I283746,I283514);
nor I_16520 (I283428,I283582,I283763);
nor I_16521 (I283443,I283681,I283531);
nand I_16522 (I283808,I283664,I283647);
and I_16523 (I283825,I283808,I424790);
nand I_16524 (I283842,I283825,I424769);
not I_16525 (I283859,I283842);
nor I_16526 (I283876,I283859,I424763);
nand I_16527 (I283893,I283630,I283842);
not I_16528 (I283434,I283893);
nor I_16529 (I283924,I424775,I424763);
or I_16530 (I283941,I283924,I424766);
nor I_16531 (I283958,I424766,I424769);
nand I_16532 (I283975,I283958,I283941);
not I_16533 (I283992,I283975);
nor I_16534 (I283455,I283992,I283548);
nand I_16535 (I284023,I283992,I283876);
nand I_16536 (I283431,I283893,I284023);
nor I_16537 (I284054,I283992,I283565);
nor I_16538 (I283452,I284054,I283582);
nor I_16539 (I283446,I283992,I283746);
nor I_16540 (I284099,I283975,I283531);
nor I_16541 (I284116,I283859,I284099);
nor I_16542 (I283437,I284116,I283715);
nor I_16543 (I284147,I283548,I283975);
nor I_16544 (I284164,I283842,I284147);
DFFARX1 I_16545 (I284164,I2898,I283463,I283449,);
not I_16546 (I284228,I2905);
or I_16547 (I284245,I140564,I140561);
nor I_16548 (I284262,I140564,I140561);
nor I_16549 (I284279,I284262,I140546);
not I_16550 (I284296,I284279);
nand I_16551 (I284313,I284245,I140567);
not I_16552 (I284330,I284313);
not I_16553 (I284347,I140549);
nor I_16554 (I284190,I284347,I284330);
nor I_16555 (I284378,I284347,I284313);
nor I_16556 (I284395,I284279,I140549);
not I_16557 (I284412,I140543);
nand I_16558 (I284429,I140552,I140540);
nand I_16559 (I284446,I284429,I140543);
nor I_16560 (I284463,I284313,I284446);
not I_16561 (I284480,I284463);
nor I_16562 (I284205,I284446,I284378);
not I_16563 (I284511,I284446);
nor I_16564 (I284528,I284511,I284279);
nor I_16565 (I284193,I284347,I284528);
nor I_16566 (I284208,I284446,I284296);
nand I_16567 (I284573,I284429,I284412);
and I_16568 (I284590,I284573,I140573);
nand I_16569 (I284607,I284590,I140570);
not I_16570 (I284624,I284607);
nor I_16571 (I284641,I284624,I140549);
nand I_16572 (I284658,I284395,I284607);
not I_16573 (I284199,I284658);
nor I_16574 (I284689,I140540,I140558);
or I_16575 (I284706,I284689,I140543);
nor I_16576 (I284723,I140555,I140546);
nand I_16577 (I284740,I284723,I284706);
not I_16578 (I284757,I284740);
nor I_16579 (I284220,I284757,I284313);
nand I_16580 (I284788,I284757,I284641);
nand I_16581 (I284196,I284658,I284788);
nor I_16582 (I284819,I284757,I284330);
nor I_16583 (I284217,I284819,I284347);
nor I_16584 (I284211,I284757,I284511);
nor I_16585 (I284864,I284740,I284296);
nor I_16586 (I284881,I284624,I284864);
nor I_16587 (I284202,I284881,I284480);
nor I_16588 (I284912,I284313,I284740);
nor I_16589 (I284929,I284607,I284912);
DFFARX1 I_16590 (I284929,I2898,I284228,I284214,);
not I_16591 (I284993,I2905);
nand I_16592 (I285010,I119160,I119181);
and I_16593 (I285027,I119160,I119181);
or I_16594 (I285044,I285027,I119157);
nand I_16595 (I285061,I285044,I285010);
and I_16596 (I285078,I285044,I119187);
and I_16597 (I285095,I285078,I119169);
or I_16598 (I285112,I119172,I119160);
nor I_16599 (I285129,I285112,I119163);
not I_16600 (I285146,I285129);
nand I_16601 (I285163,I285146,I285095);
nand I_16602 (I285180,I119175,I119157);
nor I_16603 (I285197,I285180,I119178);
not I_16604 (I285214,I285197);
nor I_16605 (I285231,I285214,I285061);
not I_16606 (I285248,I285231);
nand I_16607 (I284973,I285146,I285231);
nand I_16608 (I284967,I285095,I285214);
not I_16609 (I285293,I285180);
and I_16610 (I285310,I285293,I285061);
nand I_16611 (I285327,I285180,I285163);
DFFARX1 I_16612 (I285327,I2898,I284993,I284970,);
nor I_16613 (I285358,I119184,I119154);
not I_16614 (I285375,I119166);
nor I_16615 (I285392,I285375,I285358);
nand I_16616 (I285409,I285293,I285392);
not I_16617 (I284955,I285409);
nor I_16618 (I284958,I285129,I285409);
or I_16619 (I285454,I285197,I285392);
nor I_16620 (I284961,I285310,I285454);
nor I_16621 (I285485,I285375,I119154);
and I_16622 (I285502,I285485,I285392);
nor I_16623 (I285519,I285095,I285502);
nor I_16624 (I284979,I285519,I285502);
or I_16625 (I285550,I285146,I285519);
nor I_16626 (I285567,I285485,I285095);
nor I_16627 (I284985,I285567,I285248);
not I_16628 (I285598,I285485);
nor I_16629 (I284982,I285598,I285550);
nand I_16630 (I285629,I285598,I285061);
nor I_16631 (I284964,I285197,I285629);
nor I_16632 (I285660,I285485,I285129);
nand I_16633 (I284976,I285660,I285293);
not I_16634 (I285724,I2905);
nand I_16635 (I285741,I401303,I401318);
and I_16636 (I285758,I401303,I401318);
or I_16637 (I285775,I285758,I401309);
nand I_16638 (I285792,I285775,I285741);
and I_16639 (I285809,I285775,I401309);
and I_16640 (I285826,I285809,I401306);
or I_16641 (I285843,I401303,I401327);
nor I_16642 (I285860,I285843,I401324);
not I_16643 (I285877,I285860);
nand I_16644 (I285894,I285877,I285826);
nand I_16645 (I285911,I401321,I401315);
nor I_16646 (I285928,I285911,I401312);
not I_16647 (I285945,I285928);
nor I_16648 (I285962,I285945,I285792);
not I_16649 (I285979,I285962);
nand I_16650 (I285704,I285877,I285962);
nand I_16651 (I285698,I285826,I285945);
not I_16652 (I286024,I285911);
and I_16653 (I286041,I286024,I285792);
nand I_16654 (I286058,I285911,I285894);
DFFARX1 I_16655 (I286058,I2898,I285724,I285701,);
nor I_16656 (I286089,I401306,I401315);
not I_16657 (I286106,I401312);
nor I_16658 (I286123,I286106,I286089);
nand I_16659 (I286140,I286024,I286123);
not I_16660 (I285686,I286140);
nor I_16661 (I285689,I285860,I286140);
or I_16662 (I286185,I285928,I286123);
nor I_16663 (I285692,I286041,I286185);
nor I_16664 (I286216,I286106,I401318);
and I_16665 (I286233,I286216,I286123);
nor I_16666 (I286250,I285826,I286233);
nor I_16667 (I285710,I286250,I286233);
or I_16668 (I286281,I285877,I286250);
nor I_16669 (I286298,I286216,I285826);
nor I_16670 (I285716,I286298,I285979);
not I_16671 (I286329,I286216);
nor I_16672 (I285713,I286329,I286281);
nand I_16673 (I286360,I286329,I285792);
nor I_16674 (I285695,I285928,I286360);
nor I_16675 (I286391,I286216,I285860);
nand I_16676 (I285707,I286391,I286024);
not I_16677 (I286455,I2905);
nand I_16678 (I286472,I357960,I357945);
and I_16679 (I286489,I357960,I357945);
or I_16680 (I286506,I286489,I357945);
nand I_16681 (I286523,I286506,I286472);
and I_16682 (I286540,I286506,I357939);
and I_16683 (I286557,I286540,I357942);
or I_16684 (I286574,I357936,I357939);
nor I_16685 (I286591,I286574,I357951);
not I_16686 (I286608,I286591);
nand I_16687 (I286625,I286608,I286557);
nand I_16688 (I286642,I357942,I357948);
nor I_16689 (I286659,I286642,I357936);
not I_16690 (I286676,I286659);
nor I_16691 (I286693,I286676,I286523);
not I_16692 (I286710,I286693);
nand I_16693 (I286435,I286608,I286693);
nand I_16694 (I286429,I286557,I286676);
not I_16695 (I286755,I286642);
and I_16696 (I286772,I286755,I286523);
nand I_16697 (I286789,I286642,I286625);
DFFARX1 I_16698 (I286789,I2898,I286455,I286432,);
nor I_16699 (I286820,I357951,I357954);
not I_16700 (I286837,I357957);
nor I_16701 (I286854,I286837,I286820);
nand I_16702 (I286871,I286755,I286854);
not I_16703 (I286417,I286871);
nor I_16704 (I286420,I286591,I286871);
or I_16705 (I286916,I286659,I286854);
nor I_16706 (I286423,I286772,I286916);
nor I_16707 (I286947,I286837,I357948);
and I_16708 (I286964,I286947,I286854);
nor I_16709 (I286981,I286557,I286964);
nor I_16710 (I286441,I286981,I286964);
or I_16711 (I287012,I286608,I286981);
nor I_16712 (I287029,I286947,I286557);
nor I_16713 (I286447,I287029,I286710);
not I_16714 (I287060,I286947);
nor I_16715 (I286444,I287060,I287012);
nand I_16716 (I287091,I287060,I286523);
nor I_16717 (I286426,I286659,I287091);
nor I_16718 (I287122,I286947,I286591);
nand I_16719 (I286438,I287122,I286755);
not I_16720 (I287186,I2905);
nand I_16721 (I287203,I42585,I42552);
and I_16722 (I287220,I42585,I42552);
or I_16723 (I287237,I287220,I42582);
nand I_16724 (I287254,I287237,I287203);
and I_16725 (I287271,I287237,I42552);
and I_16726 (I287288,I287271,I42588);
or I_16727 (I287305,I42579,I42564);
nor I_16728 (I287322,I287305,I42555);
not I_16729 (I287339,I287322);
nand I_16730 (I287356,I287339,I287288);
nand I_16731 (I287373,I42570,I42576);
nor I_16732 (I287390,I287373,I42555);
not I_16733 (I287407,I287390);
nor I_16734 (I287424,I287407,I287254);
not I_16735 (I287441,I287424);
nand I_16736 (I287166,I287339,I287424);
nand I_16737 (I287160,I287288,I287407);
not I_16738 (I287486,I287373);
and I_16739 (I287503,I287486,I287254);
nand I_16740 (I287520,I287373,I287356);
DFFARX1 I_16741 (I287520,I2898,I287186,I287163,);
nor I_16742 (I287551,I42573,I42567);
not I_16743 (I287568,I42558);
nor I_16744 (I287585,I287568,I287551);
nand I_16745 (I287602,I287486,I287585);
not I_16746 (I287148,I287602);
nor I_16747 (I287151,I287322,I287602);
or I_16748 (I287647,I287390,I287585);
nor I_16749 (I287154,I287503,I287647);
nor I_16750 (I287678,I287568,I42561);
and I_16751 (I287695,I287678,I287585);
nor I_16752 (I287712,I287288,I287695);
nor I_16753 (I287172,I287712,I287695);
or I_16754 (I287743,I287339,I287712);
nor I_16755 (I287760,I287678,I287288);
nor I_16756 (I287178,I287760,I287441);
not I_16757 (I287791,I287678);
nor I_16758 (I287175,I287791,I287743);
nand I_16759 (I287822,I287791,I287254);
nor I_16760 (I287157,I287390,I287822);
nor I_16761 (I287853,I287678,I287322);
nand I_16762 (I287169,I287853,I287486);
not I_16763 (I287917,I2905);
nand I_16764 (I287934,I33208,I33208);
and I_16765 (I287951,I33208,I33208);
or I_16766 (I287968,I287951,I33217);
nand I_16767 (I287985,I287968,I287934);
and I_16768 (I288002,I287968,I33202);
and I_16769 (I288019,I288002,I33223);
or I_16770 (I288036,I33202,I33205);
nor I_16771 (I288053,I288036,I33205);
not I_16772 (I288070,I288053);
nand I_16773 (I288087,I288070,I288019);
nand I_16774 (I288104,I33211,I33214);
nor I_16775 (I288121,I288104,I33226);
not I_16776 (I288138,I288121);
nor I_16777 (I288155,I288138,I287985);
not I_16778 (I288172,I288155);
nand I_16779 (I287897,I288070,I288155);
nand I_16780 (I287891,I288019,I288138);
not I_16781 (I288217,I288104);
and I_16782 (I288234,I288217,I287985);
nand I_16783 (I288251,I288104,I288087);
DFFARX1 I_16784 (I288251,I2898,I287917,I287894,);
nor I_16785 (I288282,I33211,I33214);
not I_16786 (I288299,I33220);
nor I_16787 (I288316,I288299,I288282);
nand I_16788 (I288333,I288217,I288316);
not I_16789 (I287879,I288333);
nor I_16790 (I287882,I288053,I288333);
or I_16791 (I288378,I288121,I288316);
nor I_16792 (I287885,I288234,I288378);
nor I_16793 (I288409,I288299,I33229);
and I_16794 (I288426,I288409,I288316);
nor I_16795 (I288443,I288019,I288426);
nor I_16796 (I287903,I288443,I288426);
or I_16797 (I288474,I288070,I288443);
nor I_16798 (I288491,I288409,I288019);
nor I_16799 (I287909,I288491,I288172);
not I_16800 (I288522,I288409);
nor I_16801 (I287906,I288522,I288474);
nand I_16802 (I288553,I288522,I287985);
nor I_16803 (I287888,I288121,I288553);
nor I_16804 (I288584,I288409,I288053);
nand I_16805 (I287900,I288584,I288217);
not I_16806 (I288648,I2905);
nand I_16807 (I288665,I134885,I134906);
and I_16808 (I288682,I134885,I134906);
or I_16809 (I288699,I288682,I134882);
nand I_16810 (I288716,I288699,I288665);
and I_16811 (I288733,I288699,I134912);
and I_16812 (I288750,I288733,I134894);
or I_16813 (I288767,I134897,I134885);
nor I_16814 (I288784,I288767,I134888);
not I_16815 (I288801,I288784);
nand I_16816 (I288818,I288801,I288750);
nand I_16817 (I288835,I134900,I134882);
nor I_16818 (I288852,I288835,I134903);
not I_16819 (I288869,I288852);
nor I_16820 (I288886,I288869,I288716);
not I_16821 (I288903,I288886);
nand I_16822 (I288628,I288801,I288886);
nand I_16823 (I288622,I288750,I288869);
not I_16824 (I288948,I288835);
and I_16825 (I288965,I288948,I288716);
nand I_16826 (I288982,I288835,I288818);
DFFARX1 I_16827 (I288982,I2898,I288648,I288625,);
nor I_16828 (I289013,I134909,I134879);
not I_16829 (I289030,I134891);
nor I_16830 (I289047,I289030,I289013);
nand I_16831 (I289064,I288948,I289047);
not I_16832 (I288610,I289064);
nor I_16833 (I288613,I288784,I289064);
or I_16834 (I289109,I288852,I289047);
nor I_16835 (I288616,I288965,I289109);
nor I_16836 (I289140,I289030,I134879);
and I_16837 (I289157,I289140,I289047);
nor I_16838 (I289174,I288750,I289157);
nor I_16839 (I288634,I289174,I289157);
or I_16840 (I289205,I288801,I289174);
nor I_16841 (I289222,I289140,I288750);
nor I_16842 (I288640,I289222,I288903);
not I_16843 (I289253,I289140);
nor I_16844 (I288637,I289253,I289205);
nand I_16845 (I289284,I289253,I288716);
nor I_16846 (I288619,I288852,I289284);
nor I_16847 (I289315,I289140,I288784);
nand I_16848 (I288631,I289315,I288948);
not I_16849 (I289379,I2905);
nand I_16850 (I289396,I60711,I60735);
and I_16851 (I289413,I60711,I60735);
or I_16852 (I289430,I289413,I60723);
nand I_16853 (I289447,I289430,I289396);
and I_16854 (I289464,I289430,I60717);
and I_16855 (I289481,I289464,I60708);
or I_16856 (I289498,I60720,I60732);
nor I_16857 (I289515,I289498,I60717);
not I_16858 (I289532,I289515);
nand I_16859 (I289549,I289532,I289481);
nand I_16860 (I289566,I60714,I60726);
nor I_16861 (I289583,I289566,I60708);
not I_16862 (I289600,I289583);
nor I_16863 (I289617,I289600,I289447);
not I_16864 (I289634,I289617);
nand I_16865 (I289359,I289532,I289617);
nand I_16866 (I289353,I289481,I289600);
not I_16867 (I289679,I289566);
and I_16868 (I289696,I289679,I289447);
nand I_16869 (I289713,I289566,I289549);
DFFARX1 I_16870 (I289713,I2898,I289379,I289356,);
nor I_16871 (I289744,I60720,I60714);
not I_16872 (I289761,I60729);
nor I_16873 (I289778,I289761,I289744);
nand I_16874 (I289795,I289679,I289778);
not I_16875 (I289341,I289795);
nor I_16876 (I289344,I289515,I289795);
or I_16877 (I289840,I289583,I289778);
nor I_16878 (I289347,I289696,I289840);
nor I_16879 (I289871,I289761,I60711);
and I_16880 (I289888,I289871,I289778);
nor I_16881 (I289905,I289481,I289888);
nor I_16882 (I289365,I289905,I289888);
or I_16883 (I289936,I289532,I289905);
nor I_16884 (I289953,I289871,I289481);
nor I_16885 (I289371,I289953,I289634);
not I_16886 (I289984,I289871);
nor I_16887 (I289368,I289984,I289936);
nand I_16888 (I290015,I289984,I289447);
nor I_16889 (I289350,I289583,I290015);
nor I_16890 (I290046,I289871,I289515);
nand I_16891 (I289362,I290046,I289679);
not I_16892 (I290110,I2905);
nand I_16893 (I290127,I85871,I85895);
and I_16894 (I290144,I85871,I85895);
or I_16895 (I290161,I290144,I85883);
nand I_16896 (I290178,I290161,I290127);
and I_16897 (I290195,I290161,I85877);
and I_16898 (I290212,I290195,I85868);
or I_16899 (I290229,I85880,I85892);
nor I_16900 (I290246,I290229,I85877);
not I_16901 (I290263,I290246);
nand I_16902 (I290280,I290263,I290212);
nand I_16903 (I290297,I85874,I85886);
nor I_16904 (I290314,I290297,I85868);
not I_16905 (I290331,I290314);
nor I_16906 (I290348,I290331,I290178);
not I_16907 (I290365,I290348);
nand I_16908 (I290090,I290263,I290348);
nand I_16909 (I290084,I290212,I290331);
not I_16910 (I290410,I290297);
and I_16911 (I290427,I290410,I290178);
nand I_16912 (I290444,I290297,I290280);
DFFARX1 I_16913 (I290444,I2898,I290110,I290087,);
nor I_16914 (I290475,I85880,I85874);
not I_16915 (I290492,I85889);
nor I_16916 (I290509,I290492,I290475);
nand I_16917 (I290526,I290410,I290509);
not I_16918 (I290072,I290526);
nor I_16919 (I290075,I290246,I290526);
or I_16920 (I290571,I290314,I290509);
nor I_16921 (I290078,I290427,I290571);
nor I_16922 (I290602,I290492,I85871);
and I_16923 (I290619,I290602,I290509);
nor I_16924 (I290636,I290212,I290619);
nor I_16925 (I290096,I290636,I290619);
or I_16926 (I290667,I290263,I290636);
nor I_16927 (I290684,I290602,I290212);
nor I_16928 (I290102,I290684,I290365);
not I_16929 (I290715,I290602);
nor I_16930 (I290099,I290715,I290667);
nand I_16931 (I290746,I290715,I290178);
nor I_16932 (I290081,I290314,I290746);
nor I_16933 (I290777,I290602,I290246);
nand I_16934 (I290093,I290777,I290410);
not I_16935 (I290841,I2905);
nand I_16936 (I290858,I155886,I155880);
and I_16937 (I290875,I155886,I155880);
or I_16938 (I290892,I290875,I155904);
nand I_16939 (I290909,I290892,I290858);
and I_16940 (I290926,I290892,I155901);
and I_16941 (I290943,I290926,I155883);
or I_16942 (I290960,I155889,I155892);
nor I_16943 (I290977,I290960,I155874);
not I_16944 (I290994,I290977);
nand I_16945 (I291011,I290994,I290943);
nand I_16946 (I291028,I155877,I155907);
nor I_16947 (I291045,I291028,I155880);
not I_16948 (I291062,I291045);
nor I_16949 (I291079,I291062,I290909);
not I_16950 (I291096,I291079);
nand I_16951 (I290821,I290994,I291079);
nand I_16952 (I290815,I290943,I291062);
not I_16953 (I291141,I291028);
and I_16954 (I291158,I291141,I290909);
nand I_16955 (I291175,I291028,I291011);
DFFARX1 I_16956 (I291175,I2898,I290841,I290818,);
nor I_16957 (I291206,I155877,I155874);
not I_16958 (I291223,I155898);
nor I_16959 (I291240,I291223,I291206);
nand I_16960 (I291257,I291141,I291240);
not I_16961 (I290803,I291257);
nor I_16962 (I290806,I290977,I291257);
or I_16963 (I291302,I291045,I291240);
nor I_16964 (I290809,I291158,I291302);
nor I_16965 (I291333,I291223,I155895);
and I_16966 (I291350,I291333,I291240);
nor I_16967 (I291367,I290943,I291350);
nor I_16968 (I290827,I291367,I291350);
or I_16969 (I291398,I290994,I291367);
nor I_16970 (I291415,I291333,I290943);
nor I_16971 (I290833,I291415,I291096);
not I_16972 (I291446,I291333);
nor I_16973 (I290830,I291446,I291398);
nand I_16974 (I291477,I291446,I290909);
nor I_16975 (I290812,I291045,I291477);
nor I_16976 (I291508,I291333,I290977);
nand I_16977 (I290824,I291508,I291141);
not I_16978 (I291572,I2905);
nand I_16979 (I291589,I373868,I373874);
and I_16980 (I291606,I373868,I373874);
or I_16981 (I291623,I291606,I373898);
nand I_16982 (I291640,I291623,I291589);
and I_16983 (I291657,I291623,I373865);
and I_16984 (I291674,I291657,I373871);
or I_16985 (I291691,I373868,I373880);
nor I_16986 (I291708,I291691,I373895);
not I_16987 (I291725,I291708);
nand I_16988 (I291742,I291725,I291674);
nand I_16989 (I291759,I373886,I373883);
nor I_16990 (I291776,I291759,I373865);
not I_16991 (I291793,I291776);
nor I_16992 (I291810,I291793,I291640);
not I_16993 (I291827,I291810);
nand I_16994 (I291552,I291725,I291810);
nand I_16995 (I291546,I291674,I291793);
not I_16996 (I291872,I291759);
and I_16997 (I291889,I291872,I291640);
nand I_16998 (I291906,I291759,I291742);
DFFARX1 I_16999 (I291906,I2898,I291572,I291549,);
nor I_17000 (I291937,I373877,I373889);
not I_17001 (I291954,I373871);
nor I_17002 (I291971,I291954,I291937);
nand I_17003 (I291988,I291872,I291971);
not I_17004 (I291534,I291988);
nor I_17005 (I291537,I291708,I291988);
or I_17006 (I292033,I291776,I291971);
nor I_17007 (I291540,I291889,I292033);
nor I_17008 (I292064,I291954,I373892);
and I_17009 (I292081,I292064,I291971);
nor I_17010 (I292098,I291674,I292081);
nor I_17011 (I291558,I292098,I292081);
or I_17012 (I292129,I291725,I292098);
nor I_17013 (I292146,I292064,I291674);
nor I_17014 (I291564,I292146,I291827);
not I_17015 (I292177,I292064);
nor I_17016 (I291561,I292177,I292129);
nand I_17017 (I292208,I292177,I291640);
nor I_17018 (I291543,I291776,I292208);
nor I_17019 (I292239,I292064,I291708);
nand I_17020 (I291555,I292239,I291872);
not I_17021 (I292303,I2905);
nand I_17022 (I292320,I152486,I152480);
and I_17023 (I292337,I152486,I152480);
or I_17024 (I292354,I292337,I152504);
nand I_17025 (I292371,I292354,I292320);
and I_17026 (I292388,I292354,I152501);
and I_17027 (I292405,I292388,I152483);
or I_17028 (I292422,I152489,I152492);
nor I_17029 (I292439,I292422,I152474);
not I_17030 (I292456,I292439);
nand I_17031 (I292473,I292456,I292405);
nand I_17032 (I292490,I152477,I152507);
nor I_17033 (I292507,I292490,I152480);
not I_17034 (I292524,I292507);
nor I_17035 (I292541,I292524,I292371);
not I_17036 (I292558,I292541);
nand I_17037 (I292283,I292456,I292541);
nand I_17038 (I292277,I292405,I292524);
not I_17039 (I292603,I292490);
and I_17040 (I292620,I292603,I292371);
nand I_17041 (I292637,I292490,I292473);
DFFARX1 I_17042 (I292637,I2898,I292303,I292280,);
nor I_17043 (I292668,I152477,I152474);
not I_17044 (I292685,I152498);
nor I_17045 (I292702,I292685,I292668);
nand I_17046 (I292719,I292603,I292702);
not I_17047 (I292265,I292719);
nor I_17048 (I292268,I292439,I292719);
or I_17049 (I292764,I292507,I292702);
nor I_17050 (I292271,I292620,I292764);
nor I_17051 (I292795,I292685,I152495);
and I_17052 (I292812,I292795,I292702);
nor I_17053 (I292829,I292405,I292812);
nor I_17054 (I292289,I292829,I292812);
or I_17055 (I292860,I292456,I292829);
nor I_17056 (I292877,I292795,I292405);
nor I_17057 (I292295,I292877,I292558);
not I_17058 (I292908,I292795);
nor I_17059 (I292292,I292908,I292860);
nand I_17060 (I292939,I292908,I292371);
nor I_17061 (I292274,I292507,I292939);
nor I_17062 (I292970,I292795,I292439);
nand I_17063 (I292286,I292970,I292603);
not I_17064 (I293034,I2905);
nand I_17065 (I293051,I419884,I419890);
and I_17066 (I293068,I419884,I419890);
or I_17067 (I293085,I293068,I419890);
nand I_17068 (I293102,I293085,I293051);
and I_17069 (I293119,I293085,I419905);
and I_17070 (I293136,I293119,I419917);
or I_17071 (I293153,I419887,I419899);
nor I_17072 (I293170,I293153,I419908);
not I_17073 (I293187,I293170);
nand I_17074 (I293204,I293187,I293136);
nand I_17075 (I293221,I419914,I419896);
nor I_17076 (I293238,I293221,I419887);
not I_17077 (I293255,I293238);
nor I_17078 (I293272,I293255,I293102);
not I_17079 (I293289,I293272);
nand I_17080 (I293014,I293187,I293272);
nand I_17081 (I293008,I293136,I293255);
not I_17082 (I293334,I293221);
and I_17083 (I293351,I293334,I293102);
nand I_17084 (I293368,I293221,I293204);
DFFARX1 I_17085 (I293368,I2898,I293034,I293011,);
nor I_17086 (I293399,I419902,I419911);
not I_17087 (I293416,I419893);
nor I_17088 (I293433,I293416,I293399);
nand I_17089 (I293450,I293334,I293433);
not I_17090 (I292996,I293450);
nor I_17091 (I292999,I293170,I293450);
or I_17092 (I293495,I293238,I293433);
nor I_17093 (I293002,I293351,I293495);
nor I_17094 (I293526,I293416,I419884);
and I_17095 (I293543,I293526,I293433);
nor I_17096 (I293560,I293136,I293543);
nor I_17097 (I293020,I293560,I293543);
or I_17098 (I293591,I293187,I293560);
nor I_17099 (I293608,I293526,I293136);
nor I_17100 (I293026,I293608,I293289);
not I_17101 (I293639,I293526);
nor I_17102 (I293023,I293639,I293591);
nand I_17103 (I293670,I293639,I293102);
nor I_17104 (I293005,I293238,I293670);
nor I_17105 (I293701,I293526,I293170);
nand I_17106 (I293017,I293701,I293334);
not I_17107 (I293765,I2905);
nand I_17108 (I293782,I155206,I155200);
and I_17109 (I293799,I155206,I155200);
or I_17110 (I293816,I293799,I155224);
nand I_17111 (I293833,I293816,I293782);
and I_17112 (I293850,I293816,I155221);
and I_17113 (I293867,I293850,I155203);
or I_17114 (I293884,I155209,I155212);
nor I_17115 (I293901,I293884,I155194);
not I_17116 (I293918,I293901);
nand I_17117 (I293935,I293918,I293867);
nand I_17118 (I293952,I155197,I155227);
nor I_17119 (I293969,I293952,I155200);
not I_17120 (I293986,I293969);
nor I_17121 (I294003,I293986,I293833);
not I_17122 (I294020,I294003);
nand I_17123 (I293745,I293918,I294003);
nand I_17124 (I293739,I293867,I293986);
not I_17125 (I294065,I293952);
and I_17126 (I294082,I294065,I293833);
nand I_17127 (I294099,I293952,I293935);
DFFARX1 I_17128 (I294099,I2898,I293765,I293742,);
nor I_17129 (I294130,I155197,I155194);
not I_17130 (I294147,I155218);
nor I_17131 (I294164,I294147,I294130);
nand I_17132 (I294181,I294065,I294164);
not I_17133 (I293727,I294181);
nor I_17134 (I293730,I293901,I294181);
or I_17135 (I294226,I293969,I294164);
nor I_17136 (I293733,I294082,I294226);
nor I_17137 (I294257,I294147,I155215);
and I_17138 (I294274,I294257,I294164);
nor I_17139 (I294291,I293867,I294274);
nor I_17140 (I293751,I294291,I294274);
or I_17141 (I294322,I293918,I294291);
nor I_17142 (I294339,I294257,I293867);
nor I_17143 (I293757,I294339,I294020);
not I_17144 (I294370,I294257);
nor I_17145 (I293754,I294370,I294322);
nand I_17146 (I294401,I294370,I293833);
nor I_17147 (I293736,I293969,I294401);
nor I_17148 (I294432,I294257,I293901);
nand I_17149 (I293748,I294432,I294065);
not I_17150 (I294496,I2905);
nand I_17151 (I294513,I184863,I184860);
and I_17152 (I294530,I184863,I184860);
or I_17153 (I294547,I294530,I184848);
nand I_17154 (I294564,I294547,I294513);
and I_17155 (I294581,I294547,I184848);
and I_17156 (I294598,I294581,I184854);
or I_17157 (I294615,I184845,I184845);
nor I_17158 (I294632,I294615,I184857);
not I_17159 (I294649,I294632);
nand I_17160 (I294666,I294649,I294598);
nand I_17161 (I294683,I184866,I184851);
nor I_17162 (I294700,I294683,I184842);
not I_17163 (I294717,I294700);
nor I_17164 (I294734,I294717,I294564);
not I_17165 (I294751,I294734);
nand I_17166 (I294476,I294649,I294734);
nand I_17167 (I294470,I294598,I294717);
not I_17168 (I294796,I294683);
and I_17169 (I294813,I294796,I294564);
nand I_17170 (I294830,I294683,I294666);
DFFARX1 I_17171 (I294830,I2898,I294496,I294473,);
nor I_17172 (I294861,I184854,I184851);
not I_17173 (I294878,I184857);
nor I_17174 (I294895,I294878,I294861);
nand I_17175 (I294912,I294796,I294895);
not I_17176 (I294458,I294912);
nor I_17177 (I294461,I294632,I294912);
or I_17178 (I294957,I294700,I294895);
nor I_17179 (I294464,I294813,I294957);
nor I_17180 (I294988,I294878,I184842);
and I_17181 (I295005,I294988,I294895);
nor I_17182 (I295022,I294598,I295005);
nor I_17183 (I294482,I295022,I295005);
or I_17184 (I295053,I294649,I295022);
nor I_17185 (I295070,I294988,I294598);
nor I_17186 (I294488,I295070,I294751);
not I_17187 (I295101,I294988);
nor I_17188 (I294485,I295101,I295053);
nand I_17189 (I295132,I295101,I294564);
nor I_17190 (I294467,I294700,I295132);
nor I_17191 (I295163,I294988,I294632);
nand I_17192 (I294479,I295163,I294796);
not I_17193 (I295227,I2905);
nand I_17194 (I295244,I90903,I90927);
and I_17195 (I295261,I90903,I90927);
or I_17196 (I295278,I295261,I90915);
nand I_17197 (I295295,I295278,I295244);
and I_17198 (I295312,I295278,I90909);
and I_17199 (I295329,I295312,I90900);
or I_17200 (I295346,I90912,I90924);
nor I_17201 (I295363,I295346,I90909);
not I_17202 (I295380,I295363);
nand I_17203 (I295397,I295380,I295329);
nand I_17204 (I295414,I90906,I90918);
nor I_17205 (I295431,I295414,I90900);
not I_17206 (I295448,I295431);
nor I_17207 (I295465,I295448,I295295);
not I_17208 (I295482,I295465);
nand I_17209 (I295207,I295380,I295465);
nand I_17210 (I295201,I295329,I295448);
not I_17211 (I295527,I295414);
and I_17212 (I295544,I295527,I295295);
nand I_17213 (I295561,I295414,I295397);
DFFARX1 I_17214 (I295561,I2898,I295227,I295204,);
nor I_17215 (I295592,I90912,I90906);
not I_17216 (I295609,I90921);
nor I_17217 (I295626,I295609,I295592);
nand I_17218 (I295643,I295527,I295626);
not I_17219 (I295189,I295643);
nor I_17220 (I295192,I295363,I295643);
or I_17221 (I295688,I295431,I295626);
nor I_17222 (I295195,I295544,I295688);
nor I_17223 (I295719,I295609,I90903);
and I_17224 (I295736,I295719,I295626);
nor I_17225 (I295753,I295329,I295736);
nor I_17226 (I295213,I295753,I295736);
or I_17227 (I295784,I295380,I295753);
nor I_17228 (I295801,I295719,I295329);
nor I_17229 (I295219,I295801,I295482);
not I_17230 (I295832,I295719);
nor I_17231 (I295216,I295832,I295784);
nand I_17232 (I295863,I295832,I295295);
nor I_17233 (I295198,I295431,I295863);
nor I_17234 (I295894,I295719,I295363);
nand I_17235 (I295210,I295894,I295527);
not I_17236 (I295958,I2905);
nand I_17237 (I295975,I100919,I100940);
and I_17238 (I295992,I100919,I100940);
or I_17239 (I296009,I295992,I100916);
nand I_17240 (I296026,I296009,I295975);
and I_17241 (I296043,I296009,I100946);
and I_17242 (I296060,I296043,I100928);
or I_17243 (I296077,I100931,I100919);
nor I_17244 (I296094,I296077,I100922);
not I_17245 (I296111,I296094);
nand I_17246 (I296128,I296111,I296060);
nand I_17247 (I296145,I100934,I100916);
nor I_17248 (I296162,I296145,I100937);
not I_17249 (I296179,I296162);
nor I_17250 (I296196,I296179,I296026);
not I_17251 (I296213,I296196);
nand I_17252 (I295938,I296111,I296196);
nand I_17253 (I295932,I296060,I296179);
not I_17254 (I296258,I296145);
and I_17255 (I296275,I296258,I296026);
nand I_17256 (I296292,I296145,I296128);
DFFARX1 I_17257 (I296292,I2898,I295958,I295935,);
nor I_17258 (I296323,I100943,I100913);
not I_17259 (I296340,I100925);
nor I_17260 (I296357,I296340,I296323);
nand I_17261 (I296374,I296258,I296357);
not I_17262 (I295920,I296374);
nor I_17263 (I295923,I296094,I296374);
or I_17264 (I296419,I296162,I296357);
nor I_17265 (I295926,I296275,I296419);
nor I_17266 (I296450,I296340,I100913);
and I_17267 (I296467,I296450,I296357);
nor I_17268 (I296484,I296060,I296467);
nor I_17269 (I295944,I296484,I296467);
or I_17270 (I296515,I296111,I296484);
nor I_17271 (I296532,I296450,I296060);
nor I_17272 (I295950,I296532,I296213);
not I_17273 (I296563,I296450);
nor I_17274 (I295947,I296563,I296515);
nand I_17275 (I296594,I296563,I296026);
nor I_17276 (I295929,I296162,I296594);
nor I_17277 (I296625,I296450,I296094);
nand I_17278 (I295941,I296625,I296258);
not I_17279 (I296689,I2905);
nand I_17280 (I296706,I196712,I196709);
and I_17281 (I296723,I196712,I196709);
or I_17282 (I296740,I296723,I196697);
nand I_17283 (I296757,I296740,I296706);
and I_17284 (I296774,I296740,I196697);
and I_17285 (I296791,I296774,I196703);
or I_17286 (I296808,I196694,I196694);
nor I_17287 (I296825,I296808,I196706);
not I_17288 (I296842,I296825);
nand I_17289 (I296859,I296842,I296791);
nand I_17290 (I296876,I196715,I196700);
nor I_17291 (I296893,I296876,I196691);
not I_17292 (I296910,I296893);
nor I_17293 (I296927,I296910,I296757);
not I_17294 (I296944,I296927);
nand I_17295 (I296669,I296842,I296927);
nand I_17296 (I296663,I296791,I296910);
not I_17297 (I296989,I296876);
and I_17298 (I297006,I296989,I296757);
nand I_17299 (I297023,I296876,I296859);
DFFARX1 I_17300 (I297023,I2898,I296689,I296666,);
nor I_17301 (I297054,I196703,I196700);
not I_17302 (I297071,I196706);
nor I_17303 (I297088,I297071,I297054);
nand I_17304 (I297105,I296989,I297088);
not I_17305 (I296651,I297105);
nor I_17306 (I296654,I296825,I297105);
or I_17307 (I297150,I296893,I297088);
nor I_17308 (I296657,I297006,I297150);
nor I_17309 (I297181,I297071,I196691);
and I_17310 (I297198,I297181,I297088);
nor I_17311 (I297215,I296791,I297198);
nor I_17312 (I296675,I297215,I297198);
or I_17313 (I297246,I296842,I297215);
nor I_17314 (I297263,I297181,I296791);
nor I_17315 (I296681,I297263,I296944);
not I_17316 (I297294,I297181);
nor I_17317 (I296678,I297294,I297246);
nand I_17318 (I297325,I297294,I296757);
nor I_17319 (I296660,I296893,I297325);
nor I_17320 (I297356,I297181,I296825);
nand I_17321 (I296672,I297356,I296989);
not I_17322 (I297420,I2905);
nand I_17323 (I297437,I132998,I133019);
and I_17324 (I297454,I132998,I133019);
or I_17325 (I297471,I297454,I132995);
nand I_17326 (I297488,I297471,I297437);
and I_17327 (I297505,I297471,I133025);
and I_17328 (I297522,I297505,I133007);
or I_17329 (I297539,I133010,I132998);
nor I_17330 (I297556,I297539,I133001);
not I_17331 (I297573,I297556);
nand I_17332 (I297590,I297573,I297522);
nand I_17333 (I297607,I133013,I132995);
nor I_17334 (I297624,I297607,I133016);
not I_17335 (I297641,I297624);
nor I_17336 (I297658,I297641,I297488);
not I_17337 (I297675,I297658);
nand I_17338 (I297400,I297573,I297658);
nand I_17339 (I297394,I297522,I297641);
not I_17340 (I297720,I297607);
and I_17341 (I297737,I297720,I297488);
nand I_17342 (I297754,I297607,I297590);
DFFARX1 I_17343 (I297754,I2898,I297420,I297397,);
nor I_17344 (I297785,I133022,I132992);
not I_17345 (I297802,I133004);
nor I_17346 (I297819,I297802,I297785);
nand I_17347 (I297836,I297720,I297819);
not I_17348 (I297382,I297836);
nor I_17349 (I297385,I297556,I297836);
or I_17350 (I297881,I297624,I297819);
nor I_17351 (I297388,I297737,I297881);
nor I_17352 (I297912,I297802,I132992);
and I_17353 (I297929,I297912,I297819);
nor I_17354 (I297946,I297522,I297929);
nor I_17355 (I297406,I297946,I297929);
or I_17356 (I297977,I297573,I297946);
nor I_17357 (I297994,I297912,I297522);
nor I_17358 (I297412,I297994,I297675);
not I_17359 (I298025,I297912);
nor I_17360 (I297409,I298025,I297977);
nand I_17361 (I298056,I298025,I297488);
nor I_17362 (I297391,I297624,I298056);
nor I_17363 (I298087,I297912,I297556);
nand I_17364 (I297403,I298087,I297720);
not I_17365 (I298151,I2905);
nand I_17366 (I298168,I131111,I131132);
and I_17367 (I298185,I131111,I131132);
or I_17368 (I298202,I298185,I131108);
nand I_17369 (I298219,I298202,I298168);
and I_17370 (I298236,I298202,I131138);
and I_17371 (I298253,I298236,I131120);
or I_17372 (I298270,I131123,I131111);
nor I_17373 (I298287,I298270,I131114);
not I_17374 (I298304,I298287);
nand I_17375 (I298321,I298304,I298253);
nand I_17376 (I298338,I131126,I131108);
nor I_17377 (I298355,I298338,I131129);
not I_17378 (I298372,I298355);
nor I_17379 (I298389,I298372,I298219);
not I_17380 (I298406,I298389);
nand I_17381 (I298131,I298304,I298389);
nand I_17382 (I298125,I298253,I298372);
not I_17383 (I298451,I298338);
and I_17384 (I298468,I298451,I298219);
nand I_17385 (I298485,I298338,I298321);
DFFARX1 I_17386 (I298485,I2898,I298151,I298128,);
nor I_17387 (I298516,I131135,I131105);
not I_17388 (I298533,I131117);
nor I_17389 (I298550,I298533,I298516);
nand I_17390 (I298567,I298451,I298550);
not I_17391 (I298113,I298567);
nor I_17392 (I298116,I298287,I298567);
or I_17393 (I298612,I298355,I298550);
nor I_17394 (I298119,I298468,I298612);
nor I_17395 (I298643,I298533,I131105);
and I_17396 (I298660,I298643,I298550);
nor I_17397 (I298677,I298253,I298660);
nor I_17398 (I298137,I298677,I298660);
or I_17399 (I298708,I298304,I298677);
nor I_17400 (I298725,I298643,I298253);
nor I_17401 (I298143,I298725,I298406);
not I_17402 (I298756,I298643);
nor I_17403 (I298140,I298756,I298708);
nand I_17404 (I298787,I298756,I298219);
nor I_17405 (I298122,I298355,I298787);
nor I_17406 (I298818,I298643,I298287);
nand I_17407 (I298134,I298818,I298451);
not I_17408 (I298882,I2905);
nand I_17409 (I298899,I151806,I151800);
and I_17410 (I298916,I151806,I151800);
or I_17411 (I298933,I298916,I151824);
nand I_17412 (I298950,I298933,I298899);
and I_17413 (I298967,I298933,I151821);
and I_17414 (I298984,I298967,I151803);
or I_17415 (I299001,I151809,I151812);
nor I_17416 (I299018,I299001,I151794);
not I_17417 (I299035,I299018);
nand I_17418 (I299052,I299035,I298984);
nand I_17419 (I299069,I151797,I151827);
nor I_17420 (I299086,I299069,I151800);
not I_17421 (I299103,I299086);
nor I_17422 (I299120,I299103,I298950);
not I_17423 (I299137,I299120);
nand I_17424 (I298862,I299035,I299120);
nand I_17425 (I298856,I298984,I299103);
not I_17426 (I299182,I299069);
and I_17427 (I299199,I299182,I298950);
nand I_17428 (I299216,I299069,I299052);
DFFARX1 I_17429 (I299216,I2898,I298882,I298859,);
nor I_17430 (I299247,I151797,I151794);
not I_17431 (I299264,I151818);
nor I_17432 (I299281,I299264,I299247);
nand I_17433 (I299298,I299182,I299281);
not I_17434 (I298844,I299298);
nor I_17435 (I298847,I299018,I299298);
or I_17436 (I299343,I299086,I299281);
nor I_17437 (I298850,I299199,I299343);
nor I_17438 (I299374,I299264,I151815);
and I_17439 (I299391,I299374,I299281);
nor I_17440 (I299408,I298984,I299391);
nor I_17441 (I298868,I299408,I299391);
or I_17442 (I299439,I299035,I299408);
nor I_17443 (I299456,I299374,I298984);
nor I_17444 (I298874,I299456,I299137);
not I_17445 (I299487,I299374);
nor I_17446 (I298871,I299487,I299439);
nand I_17447 (I299518,I299487,I298950);
nor I_17448 (I298853,I299086,I299518);
nor I_17449 (I299549,I299374,I299018);
nand I_17450 (I298865,I299549,I299182);
not I_17451 (I299613,I2905);
nand I_17452 (I299630,I168126,I168120);
and I_17453 (I299647,I168126,I168120);
or I_17454 (I299664,I299647,I168144);
nand I_17455 (I299681,I299664,I299630);
and I_17456 (I299698,I299664,I168141);
and I_17457 (I299715,I299698,I168123);
or I_17458 (I299732,I168129,I168132);
nor I_17459 (I299749,I299732,I168114);
not I_17460 (I299766,I299749);
nand I_17461 (I299783,I299766,I299715);
nand I_17462 (I299800,I168117,I168147);
nor I_17463 (I299817,I299800,I168120);
not I_17464 (I299834,I299817);
nor I_17465 (I299851,I299834,I299681);
not I_17466 (I299868,I299851);
nand I_17467 (I299593,I299766,I299851);
nand I_17468 (I299587,I299715,I299834);
not I_17469 (I299913,I299800);
and I_17470 (I299930,I299913,I299681);
nand I_17471 (I299947,I299800,I299783);
DFFARX1 I_17472 (I299947,I2898,I299613,I299590,);
nor I_17473 (I299978,I168117,I168114);
not I_17474 (I299995,I168138);
nor I_17475 (I300012,I299995,I299978);
nand I_17476 (I300029,I299913,I300012);
not I_17477 (I299575,I300029);
nor I_17478 (I299578,I299749,I300029);
or I_17479 (I300074,I299817,I300012);
nor I_17480 (I299581,I299930,I300074);
nor I_17481 (I300105,I299995,I168135);
and I_17482 (I300122,I300105,I300012);
nor I_17483 (I300139,I299715,I300122);
nor I_17484 (I299599,I300139,I300122);
or I_17485 (I300170,I299766,I300139);
nor I_17486 (I300187,I300105,I299715);
nor I_17487 (I299605,I300187,I299868);
not I_17488 (I300218,I300105);
nor I_17489 (I299602,I300218,I300170);
nand I_17490 (I300249,I300218,I299681);
nor I_17491 (I299584,I299817,I300249);
nor I_17492 (I300280,I300105,I299749);
nand I_17493 (I299596,I300280,I299913);
not I_17494 (I300344,I2905);
nand I_17495 (I300361,I325830,I325815);
and I_17496 (I300378,I325830,I325815);
or I_17497 (I300395,I300378,I325815);
nand I_17498 (I300412,I300395,I300361);
and I_17499 (I300429,I300395,I325809);
and I_17500 (I300446,I300429,I325812);
or I_17501 (I300463,I325806,I325809);
nor I_17502 (I300480,I300463,I325821);
not I_17503 (I300497,I300480);
nand I_17504 (I300514,I300497,I300446);
nand I_17505 (I300531,I325812,I325818);
nor I_17506 (I300548,I300531,I325806);
not I_17507 (I300565,I300548);
nor I_17508 (I300582,I300565,I300412);
not I_17509 (I300599,I300582);
nand I_17510 (I300324,I300497,I300582);
nand I_17511 (I300318,I300446,I300565);
not I_17512 (I300644,I300531);
and I_17513 (I300661,I300644,I300412);
nand I_17514 (I300678,I300531,I300514);
DFFARX1 I_17515 (I300678,I2898,I300344,I300321,);
nor I_17516 (I300709,I325821,I325824);
not I_17517 (I300726,I325827);
nor I_17518 (I300743,I300726,I300709);
nand I_17519 (I300760,I300644,I300743);
not I_17520 (I300306,I300760);
nor I_17521 (I300309,I300480,I300760);
or I_17522 (I300805,I300548,I300743);
nor I_17523 (I300312,I300661,I300805);
nor I_17524 (I300836,I300726,I325818);
and I_17525 (I300853,I300836,I300743);
nor I_17526 (I300870,I300446,I300853);
nor I_17527 (I300330,I300870,I300853);
or I_17528 (I300901,I300497,I300870);
nor I_17529 (I300918,I300836,I300446);
nor I_17530 (I300336,I300918,I300599);
not I_17531 (I300949,I300836);
nor I_17532 (I300333,I300949,I300901);
nand I_17533 (I300980,I300949,I300412);
nor I_17534 (I300315,I300548,I300980);
nor I_17535 (I301011,I300836,I300480);
nand I_17536 (I300327,I301011,I300644);
not I_17537 (I301075,I2905);
nand I_17538 (I301092,I13312,I13315);
and I_17539 (I301109,I13312,I13315);
or I_17540 (I301126,I301109,I13318);
nand I_17541 (I301143,I301126,I301092);
and I_17542 (I301160,I301126,I13342);
and I_17543 (I301177,I301160,I13318);
or I_17544 (I301194,I13339,I13315);
nor I_17545 (I301211,I301194,I13333);
not I_17546 (I301228,I301211);
nand I_17547 (I301245,I301228,I301177);
nand I_17548 (I301262,I13330,I13321);
nor I_17549 (I301279,I301262,I13324);
not I_17550 (I301296,I301279);
nor I_17551 (I301313,I301296,I301143);
not I_17552 (I301330,I301313);
nand I_17553 (I301055,I301228,I301313);
nand I_17554 (I301049,I301177,I301296);
not I_17555 (I301375,I301262);
and I_17556 (I301392,I301375,I301143);
nand I_17557 (I301409,I301262,I301245);
DFFARX1 I_17558 (I301409,I2898,I301075,I301052,);
nor I_17559 (I301440,I13312,I13321);
not I_17560 (I301457,I13336);
nor I_17561 (I301474,I301457,I301440);
nand I_17562 (I301491,I301375,I301474);
not I_17563 (I301037,I301491);
nor I_17564 (I301040,I301211,I301491);
or I_17565 (I301536,I301279,I301474);
nor I_17566 (I301043,I301392,I301536);
nor I_17567 (I301567,I301457,I13327);
and I_17568 (I301584,I301567,I301474);
nor I_17569 (I301601,I301177,I301584);
nor I_17570 (I301061,I301601,I301584);
or I_17571 (I301632,I301228,I301601);
nor I_17572 (I301649,I301567,I301177);
nor I_17573 (I301067,I301649,I301330);
not I_17574 (I301680,I301567);
nor I_17575 (I301064,I301680,I301632);
nand I_17576 (I301711,I301680,I301143);
nor I_17577 (I301046,I301279,I301711);
nor I_17578 (I301742,I301567,I301211);
nand I_17579 (I301058,I301742,I301375);
not I_17580 (I301806,I2905);
nand I_17581 (I301823,I78952,I78976);
and I_17582 (I301840,I78952,I78976);
or I_17583 (I301857,I301840,I78964);
nand I_17584 (I301874,I301857,I301823);
and I_17585 (I301891,I301857,I78958);
and I_17586 (I301908,I301891,I78949);
or I_17587 (I301925,I78961,I78973);
nor I_17588 (I301942,I301925,I78958);
not I_17589 (I301959,I301942);
nand I_17590 (I301976,I301959,I301908);
nand I_17591 (I301993,I78955,I78967);
nor I_17592 (I302010,I301993,I78949);
not I_17593 (I302027,I302010);
nor I_17594 (I302044,I302027,I301874);
not I_17595 (I302061,I302044);
nand I_17596 (I301786,I301959,I302044);
nand I_17597 (I301780,I301908,I302027);
not I_17598 (I302106,I301993);
and I_17599 (I302123,I302106,I301874);
nand I_17600 (I302140,I301993,I301976);
DFFARX1 I_17601 (I302140,I2898,I301806,I301783,);
nor I_17602 (I302171,I78961,I78955);
not I_17603 (I302188,I78970);
nor I_17604 (I302205,I302188,I302171);
nand I_17605 (I302222,I302106,I302205);
not I_17606 (I301768,I302222);
nor I_17607 (I301771,I301942,I302222);
or I_17608 (I302267,I302010,I302205);
nor I_17609 (I301774,I302123,I302267);
nor I_17610 (I302298,I302188,I78952);
and I_17611 (I302315,I302298,I302205);
nor I_17612 (I302332,I301908,I302315);
nor I_17613 (I301792,I302332,I302315);
or I_17614 (I302363,I301959,I302332);
nor I_17615 (I302380,I302298,I301908);
nor I_17616 (I301798,I302380,I302061);
not I_17617 (I302411,I302298);
nor I_17618 (I301795,I302411,I302363);
nand I_17619 (I302442,I302411,I301874);
nor I_17620 (I301777,I302010,I302442);
nor I_17621 (I302473,I302298,I301942);
nand I_17622 (I301789,I302473,I302106);
not I_17623 (I302537,I2905);
nand I_17624 (I302554,I390664,I390670);
and I_17625 (I302571,I390664,I390670);
or I_17626 (I302588,I302571,I390694);
nand I_17627 (I302605,I302588,I302554);
and I_17628 (I302622,I302588,I390661);
and I_17629 (I302639,I302622,I390667);
or I_17630 (I302656,I390664,I390676);
nor I_17631 (I302673,I302656,I390691);
not I_17632 (I302690,I302673);
nand I_17633 (I302707,I302690,I302639);
nand I_17634 (I302724,I390682,I390679);
nor I_17635 (I302741,I302724,I390661);
not I_17636 (I302758,I302741);
nor I_17637 (I302775,I302758,I302605);
not I_17638 (I302792,I302775);
nand I_17639 (I302517,I302690,I302775);
nand I_17640 (I302511,I302639,I302758);
not I_17641 (I302837,I302724);
and I_17642 (I302854,I302837,I302605);
nand I_17643 (I302871,I302724,I302707);
DFFARX1 I_17644 (I302871,I2898,I302537,I302514,);
nor I_17645 (I302902,I390673,I390685);
not I_17646 (I302919,I390667);
nor I_17647 (I302936,I302919,I302902);
nand I_17648 (I302953,I302837,I302936);
not I_17649 (I302499,I302953);
nor I_17650 (I302502,I302673,I302953);
or I_17651 (I302998,I302741,I302936);
nor I_17652 (I302505,I302854,I302998);
nor I_17653 (I303029,I302919,I390688);
and I_17654 (I303046,I303029,I302936);
nor I_17655 (I303063,I302639,I303046);
nor I_17656 (I302523,I303063,I303046);
or I_17657 (I303094,I302690,I303063);
nor I_17658 (I303111,I303029,I302639);
nor I_17659 (I302529,I303111,I302792);
not I_17660 (I303142,I303029);
nor I_17661 (I302526,I303142,I303094);
nand I_17662 (I303173,I303142,I302605);
nor I_17663 (I302508,I302741,I303173);
nor I_17664 (I303204,I303029,I302673);
nand I_17665 (I302520,I303204,I302837);
not I_17666 (I303268,I2905);
nand I_17667 (I303285,I386142,I386148);
and I_17668 (I303302,I386142,I386148);
or I_17669 (I303319,I303302,I386172);
nand I_17670 (I303336,I303319,I303285);
and I_17671 (I303353,I303319,I386139);
and I_17672 (I303370,I303353,I386145);
or I_17673 (I303387,I386142,I386154);
nor I_17674 (I303404,I303387,I386169);
not I_17675 (I303421,I303404);
nand I_17676 (I303438,I303421,I303370);
nand I_17677 (I303455,I386160,I386157);
nor I_17678 (I303472,I303455,I386139);
not I_17679 (I303489,I303472);
nor I_17680 (I303506,I303489,I303336);
not I_17681 (I303523,I303506);
nand I_17682 (I303248,I303421,I303506);
nand I_17683 (I303242,I303370,I303489);
not I_17684 (I303568,I303455);
and I_17685 (I303585,I303568,I303336);
nand I_17686 (I303602,I303455,I303438);
DFFARX1 I_17687 (I303602,I2898,I303268,I303245,);
nor I_17688 (I303633,I386151,I386163);
not I_17689 (I303650,I386145);
nor I_17690 (I303667,I303650,I303633);
nand I_17691 (I303684,I303568,I303667);
not I_17692 (I303230,I303684);
nor I_17693 (I303233,I303404,I303684);
or I_17694 (I303729,I303472,I303667);
nor I_17695 (I303236,I303585,I303729);
nor I_17696 (I303760,I303650,I386166);
and I_17697 (I303777,I303760,I303667);
nor I_17698 (I303794,I303370,I303777);
nor I_17699 (I303254,I303794,I303777);
or I_17700 (I303825,I303421,I303794);
nor I_17701 (I303842,I303760,I303370);
nor I_17702 (I303260,I303842,I303523);
not I_17703 (I303873,I303760);
nor I_17704 (I303257,I303873,I303825);
nand I_17705 (I303904,I303873,I303336);
nor I_17706 (I303239,I303472,I303904);
nor I_17707 (I303935,I303760,I303404);
nand I_17708 (I303251,I303935,I303568);
not I_17709 (I303999,I2905);
nand I_17710 (I304016,I444976,I444982);
and I_17711 (I304033,I444976,I444982);
or I_17712 (I304050,I304033,I444982);
nand I_17713 (I304067,I304050,I304016);
and I_17714 (I304084,I304050,I444997);
and I_17715 (I304101,I304084,I445009);
or I_17716 (I304118,I444979,I444991);
nor I_17717 (I304135,I304118,I445000);
not I_17718 (I304152,I304135);
nand I_17719 (I304169,I304152,I304101);
nand I_17720 (I304186,I445006,I444988);
nor I_17721 (I304203,I304186,I444979);
not I_17722 (I304220,I304203);
nor I_17723 (I304237,I304220,I304067);
not I_17724 (I304254,I304237);
nand I_17725 (I303979,I304152,I304237);
nand I_17726 (I303973,I304101,I304220);
not I_17727 (I304299,I304186);
and I_17728 (I304316,I304299,I304067);
nand I_17729 (I304333,I304186,I304169);
DFFARX1 I_17730 (I304333,I2898,I303999,I303976,);
nor I_17731 (I304364,I444994,I445003);
not I_17732 (I304381,I444985);
nor I_17733 (I304398,I304381,I304364);
nand I_17734 (I304415,I304299,I304398);
not I_17735 (I303961,I304415);
nor I_17736 (I303964,I304135,I304415);
or I_17737 (I304460,I304203,I304398);
nor I_17738 (I303967,I304316,I304460);
nor I_17739 (I304491,I304381,I444976);
and I_17740 (I304508,I304491,I304398);
nor I_17741 (I304525,I304101,I304508);
nor I_17742 (I303985,I304525,I304508);
or I_17743 (I304556,I304152,I304525);
nor I_17744 (I304573,I304491,I304101);
nor I_17745 (I303991,I304573,I304254);
not I_17746 (I304604,I304491);
nor I_17747 (I303988,I304604,I304556);
nand I_17748 (I304635,I304604,I304067);
nor I_17749 (I303970,I304203,I304635);
nor I_17750 (I304666,I304491,I304135);
nand I_17751 (I303982,I304666,I304299);
not I_17752 (I304730,I2905);
nand I_17753 (I304747,I442885,I442891);
and I_17754 (I304764,I442885,I442891);
or I_17755 (I304781,I304764,I442891);
nand I_17756 (I304798,I304781,I304747);
and I_17757 (I304815,I304781,I442906);
and I_17758 (I304832,I304815,I442918);
or I_17759 (I304849,I442888,I442900);
nor I_17760 (I304866,I304849,I442909);
not I_17761 (I304883,I304866);
nand I_17762 (I304900,I304883,I304832);
nand I_17763 (I304917,I442915,I442897);
nor I_17764 (I304934,I304917,I442888);
not I_17765 (I304951,I304934);
nor I_17766 (I304968,I304951,I304798);
not I_17767 (I304985,I304968);
nand I_17768 (I304710,I304883,I304968);
nand I_17769 (I304704,I304832,I304951);
not I_17770 (I305030,I304917);
and I_17771 (I305047,I305030,I304798);
nand I_17772 (I305064,I304917,I304900);
DFFARX1 I_17773 (I305064,I2898,I304730,I304707,);
nor I_17774 (I305095,I442903,I442912);
not I_17775 (I305112,I442894);
nor I_17776 (I305129,I305112,I305095);
nand I_17777 (I305146,I305030,I305129);
not I_17778 (I304692,I305146);
nor I_17779 (I304695,I304866,I305146);
or I_17780 (I305191,I304934,I305129);
nor I_17781 (I304698,I305047,I305191);
nor I_17782 (I305222,I305112,I442885);
and I_17783 (I305239,I305222,I305129);
nor I_17784 (I305256,I304832,I305239);
nor I_17785 (I304716,I305256,I305239);
or I_17786 (I305287,I304883,I305256);
nor I_17787 (I305304,I305222,I304832);
nor I_17788 (I304722,I305304,I304985);
not I_17789 (I305335,I305222);
nor I_17790 (I304719,I305335,I305287);
nand I_17791 (I305366,I305335,I304798);
nor I_17792 (I304701,I304934,I305366);
nor I_17793 (I305397,I305222,I304866);
nand I_17794 (I304713,I305397,I305030);
not I_17795 (I305461,I2905);
nand I_17796 (I305478,I143062,I143083);
and I_17797 (I305495,I143062,I143083);
or I_17798 (I305512,I305495,I143059);
nand I_17799 (I305529,I305512,I305478);
and I_17800 (I305546,I305512,I143089);
and I_17801 (I305563,I305546,I143071);
or I_17802 (I305580,I143074,I143062);
nor I_17803 (I305597,I305580,I143065);
not I_17804 (I305614,I305597);
nand I_17805 (I305631,I305614,I305563);
nand I_17806 (I305648,I143077,I143059);
nor I_17807 (I305665,I305648,I143080);
not I_17808 (I305682,I305665);
nor I_17809 (I305699,I305682,I305529);
not I_17810 (I305716,I305699);
nand I_17811 (I305441,I305614,I305699);
nand I_17812 (I305435,I305563,I305682);
not I_17813 (I305761,I305648);
and I_17814 (I305778,I305761,I305529);
nand I_17815 (I305795,I305648,I305631);
DFFARX1 I_17816 (I305795,I2898,I305461,I305438,);
nor I_17817 (I305826,I143086,I143056);
not I_17818 (I305843,I143068);
nor I_17819 (I305860,I305843,I305826);
nand I_17820 (I305877,I305761,I305860);
not I_17821 (I305423,I305877);
nor I_17822 (I305426,I305597,I305877);
or I_17823 (I305922,I305665,I305860);
nor I_17824 (I305429,I305778,I305922);
nor I_17825 (I305953,I305843,I143056);
and I_17826 (I305970,I305953,I305860);
nor I_17827 (I305987,I305563,I305970);
nor I_17828 (I305447,I305987,I305970);
or I_17829 (I306018,I305614,I305987);
nor I_17830 (I306035,I305953,I305563);
nor I_17831 (I305453,I306035,I305716);
not I_17832 (I306066,I305953);
nor I_17833 (I305450,I306066,I306018);
nand I_17834 (I306097,I306066,I305529);
nor I_17835 (I305432,I305665,I306097);
nor I_17836 (I306128,I305953,I305597);
nand I_17837 (I305444,I306128,I305761);
not I_17838 (I306192,I2905);
nand I_17839 (I306209,I110354,I110375);
and I_17840 (I306226,I110354,I110375);
or I_17841 (I306243,I306226,I110351);
nand I_17842 (I306260,I306243,I306209);
and I_17843 (I306277,I306243,I110381);
and I_17844 (I306294,I306277,I110363);
or I_17845 (I306311,I110366,I110354);
nor I_17846 (I306328,I306311,I110357);
not I_17847 (I306345,I306328);
nand I_17848 (I306362,I306345,I306294);
nand I_17849 (I306379,I110369,I110351);
nor I_17850 (I306396,I306379,I110372);
not I_17851 (I306413,I306396);
nor I_17852 (I306430,I306413,I306260);
not I_17853 (I306447,I306430);
nand I_17854 (I306172,I306345,I306430);
nand I_17855 (I306166,I306294,I306413);
not I_17856 (I306492,I306379);
and I_17857 (I306509,I306492,I306260);
nand I_17858 (I306526,I306379,I306362);
DFFARX1 I_17859 (I306526,I2898,I306192,I306169,);
nor I_17860 (I306557,I110378,I110348);
not I_17861 (I306574,I110360);
nor I_17862 (I306591,I306574,I306557);
nand I_17863 (I306608,I306492,I306591);
not I_17864 (I306154,I306608);
nor I_17865 (I306157,I306328,I306608);
or I_17866 (I306653,I306396,I306591);
nor I_17867 (I306160,I306509,I306653);
nor I_17868 (I306684,I306574,I110348);
and I_17869 (I306701,I306684,I306591);
nor I_17870 (I306718,I306294,I306701);
nor I_17871 (I306178,I306718,I306701);
or I_17872 (I306749,I306345,I306718);
nor I_17873 (I306766,I306684,I306294);
nor I_17874 (I306184,I306766,I306447);
not I_17875 (I306797,I306684);
nor I_17876 (I306181,I306797,I306749);
nand I_17877 (I306828,I306797,I306260);
nor I_17878 (I306163,I306396,I306828);
nor I_17879 (I306859,I306684,I306328);
nand I_17880 (I306175,I306859,I306492);
not I_17881 (I306923,I2905);
nand I_17882 (I306940,I386788,I386794);
and I_17883 (I306957,I386788,I386794);
or I_17884 (I306974,I306957,I386818);
nand I_17885 (I306991,I306974,I306940);
and I_17886 (I307008,I306974,I386785);
and I_17887 (I307025,I307008,I386791);
or I_17888 (I307042,I386788,I386800);
nor I_17889 (I307059,I307042,I386815);
not I_17890 (I307076,I307059);
nand I_17891 (I307093,I307076,I307025);
nand I_17892 (I307110,I386806,I386803);
nor I_17893 (I307127,I307110,I386785);
not I_17894 (I307144,I307127);
nor I_17895 (I307161,I307144,I306991);
not I_17896 (I307178,I307161);
nand I_17897 (I306903,I307076,I307161);
nand I_17898 (I306897,I307025,I307144);
not I_17899 (I307223,I307110);
and I_17900 (I307240,I307223,I306991);
nand I_17901 (I307257,I307110,I307093);
DFFARX1 I_17902 (I307257,I2898,I306923,I306900,);
nor I_17903 (I307288,I386797,I386809);
not I_17904 (I307305,I386791);
nor I_17905 (I307322,I307305,I307288);
nand I_17906 (I307339,I307223,I307322);
not I_17907 (I306885,I307339);
nor I_17908 (I306888,I307059,I307339);
or I_17909 (I307384,I307127,I307322);
nor I_17910 (I306891,I307240,I307384);
nor I_17911 (I307415,I307305,I386812);
and I_17912 (I307432,I307415,I307322);
nor I_17913 (I307449,I307025,I307432);
nor I_17914 (I306909,I307449,I307432);
or I_17915 (I307480,I307076,I307449);
nor I_17916 (I307497,I307415,I307025);
nor I_17917 (I306915,I307497,I307178);
not I_17918 (I307528,I307415);
nor I_17919 (I306912,I307528,I307480);
nand I_17920 (I307559,I307528,I306991);
nor I_17921 (I306894,I307127,I307559);
nor I_17922 (I307590,I307415,I307059);
nand I_17923 (I306906,I307590,I307223);
not I_17924 (I307654,I2905);
nand I_17925 (I307671,I178365,I178371);
and I_17926 (I307688,I178365,I178371);
or I_17927 (I307705,I307688,I178377);
nand I_17928 (I307722,I307705,I307671);
and I_17929 (I307739,I307705,I178386);
and I_17930 (I307756,I307739,I178374);
or I_17931 (I307773,I178374,I178371);
nor I_17932 (I307790,I307773,I178392);
not I_17933 (I307807,I307790);
nand I_17934 (I307824,I307807,I307756);
nand I_17935 (I307841,I178368,I178365);
nor I_17936 (I307858,I307841,I178389);
not I_17937 (I307875,I307858);
nor I_17938 (I307892,I307875,I307722);
not I_17939 (I307909,I307892);
nand I_17940 (I307634,I307807,I307892);
nand I_17941 (I307628,I307756,I307875);
not I_17942 (I307954,I307841);
and I_17943 (I307971,I307954,I307722);
nand I_17944 (I307988,I307841,I307824);
DFFARX1 I_17945 (I307988,I2898,I307654,I307631,);
nor I_17946 (I308019,I178380,I178395);
not I_17947 (I308036,I178368);
nor I_17948 (I308053,I308036,I308019);
nand I_17949 (I308070,I307954,I308053);
not I_17950 (I307616,I308070);
nor I_17951 (I307619,I307790,I308070);
or I_17952 (I308115,I307858,I308053);
nor I_17953 (I307622,I307971,I308115);
nor I_17954 (I308146,I308036,I178383);
and I_17955 (I308163,I308146,I308053);
nor I_17956 (I308180,I307756,I308163);
nor I_17957 (I307640,I308180,I308163);
or I_17958 (I308211,I307807,I308180);
nor I_17959 (I308228,I308146,I307756);
nor I_17960 (I307646,I308228,I307909);
not I_17961 (I308259,I308146);
nor I_17962 (I307643,I308259,I308211);
nand I_17963 (I308290,I308259,I307722);
nor I_17964 (I307625,I307858,I308290);
nor I_17965 (I308321,I308146,I307790);
nand I_17966 (I307637,I308321,I307954);
not I_17967 (I308385,I2905);
nand I_17968 (I308402,I354390,I354375);
and I_17969 (I308419,I354390,I354375);
or I_17970 (I308436,I308419,I354375);
nand I_17971 (I308453,I308436,I308402);
and I_17972 (I308470,I308436,I354369);
and I_17973 (I308487,I308470,I354372);
or I_17974 (I308504,I354366,I354369);
nor I_17975 (I308521,I308504,I354381);
not I_17976 (I308538,I308521);
nand I_17977 (I308555,I308538,I308487);
nand I_17978 (I308572,I354372,I354378);
nor I_17979 (I308589,I308572,I354366);
not I_17980 (I308606,I308589);
nor I_17981 (I308623,I308606,I308453);
not I_17982 (I308640,I308623);
nand I_17983 (I308365,I308538,I308623);
nand I_17984 (I308359,I308487,I308606);
not I_17985 (I308685,I308572);
and I_17986 (I308702,I308685,I308453);
nand I_17987 (I308719,I308572,I308555);
DFFARX1 I_17988 (I308719,I2898,I308385,I308362,);
nor I_17989 (I308750,I354381,I354384);
not I_17990 (I308767,I354387);
nor I_17991 (I308784,I308767,I308750);
nand I_17992 (I308801,I308685,I308784);
not I_17993 (I308347,I308801);
nor I_17994 (I308350,I308521,I308801);
or I_17995 (I308846,I308589,I308784);
nor I_17996 (I308353,I308702,I308846);
nor I_17997 (I308877,I308767,I354378);
and I_17998 (I308894,I308877,I308784);
nor I_17999 (I308911,I308487,I308894);
nor I_18000 (I308371,I308911,I308894);
or I_18001 (I308942,I308538,I308911);
nor I_18002 (I308959,I308877,I308487);
nor I_18003 (I308377,I308959,I308640);
not I_18004 (I308990,I308877);
nor I_18005 (I308374,I308990,I308942);
nand I_18006 (I309021,I308990,I308453);
nor I_18007 (I308356,I308589,I309021);
nor I_18008 (I309052,I308877,I308521);
nand I_18009 (I308368,I309052,I308685);
not I_18010 (I309116,I2905);
nand I_18011 (I309133,I70775,I70799);
and I_18012 (I309150,I70775,I70799);
or I_18013 (I309167,I309150,I70787);
nand I_18014 (I309184,I309167,I309133);
and I_18015 (I309201,I309167,I70781);
and I_18016 (I309218,I309201,I70772);
or I_18017 (I309235,I70784,I70796);
nor I_18018 (I309252,I309235,I70781);
not I_18019 (I309269,I309252);
nand I_18020 (I309286,I309269,I309218);
nand I_18021 (I309303,I70778,I70790);
nor I_18022 (I309320,I309303,I70772);
not I_18023 (I309337,I309320);
nor I_18024 (I309354,I309337,I309184);
not I_18025 (I309371,I309354);
nand I_18026 (I309096,I309269,I309354);
nand I_18027 (I309090,I309218,I309337);
not I_18028 (I309416,I309303);
and I_18029 (I309433,I309416,I309184);
nand I_18030 (I309450,I309303,I309286);
DFFARX1 I_18031 (I309450,I2898,I309116,I309093,);
nor I_18032 (I309481,I70784,I70778);
not I_18033 (I309498,I70793);
nor I_18034 (I309515,I309498,I309481);
nand I_18035 (I309532,I309416,I309515);
not I_18036 (I309078,I309532);
nor I_18037 (I309081,I309252,I309532);
or I_18038 (I309577,I309320,I309515);
nor I_18039 (I309084,I309433,I309577);
nor I_18040 (I309608,I309498,I70775);
and I_18041 (I309625,I309608,I309515);
nor I_18042 (I309642,I309218,I309625);
nor I_18043 (I309102,I309642,I309625);
or I_18044 (I309673,I309269,I309642);
nor I_18045 (I309690,I309608,I309218);
nor I_18046 (I309108,I309690,I309371);
not I_18047 (I309721,I309608);
nor I_18048 (I309105,I309721,I309673);
nand I_18049 (I309752,I309721,I309184);
nor I_18050 (I309087,I309320,I309752);
nor I_18051 (I309783,I309608,I309252);
nand I_18052 (I309099,I309783,I309416);
not I_18053 (I309847,I2905);
nand I_18054 (I309864,I10864,I10867);
and I_18055 (I309881,I10864,I10867);
or I_18056 (I309898,I309881,I10870);
nand I_18057 (I309915,I309898,I309864);
and I_18058 (I309932,I309898,I10894);
and I_18059 (I309949,I309932,I10870);
or I_18060 (I309966,I10891,I10867);
nor I_18061 (I309983,I309966,I10885);
not I_18062 (I310000,I309983);
nand I_18063 (I310017,I310000,I309949);
nand I_18064 (I310034,I10882,I10873);
nor I_18065 (I310051,I310034,I10876);
not I_18066 (I310068,I310051);
nor I_18067 (I310085,I310068,I309915);
not I_18068 (I310102,I310085);
nand I_18069 (I309827,I310000,I310085);
nand I_18070 (I309821,I309949,I310068);
not I_18071 (I310147,I310034);
and I_18072 (I310164,I310147,I309915);
nand I_18073 (I310181,I310034,I310017);
DFFARX1 I_18074 (I310181,I2898,I309847,I309824,);
nor I_18075 (I310212,I10864,I10873);
not I_18076 (I310229,I10888);
nor I_18077 (I310246,I310229,I310212);
nand I_18078 (I310263,I310147,I310246);
not I_18079 (I309809,I310263);
nor I_18080 (I309812,I309983,I310263);
or I_18081 (I310308,I310051,I310246);
nor I_18082 (I309815,I310164,I310308);
nor I_18083 (I310339,I310229,I10879);
and I_18084 (I310356,I310339,I310246);
nor I_18085 (I310373,I309949,I310356);
nor I_18086 (I309833,I310373,I310356);
or I_18087 (I310404,I310000,I310373);
nor I_18088 (I310421,I310339,I309949);
nor I_18089 (I309839,I310421,I310102);
not I_18090 (I310452,I310339);
nor I_18091 (I309836,I310452,I310404);
nand I_18092 (I310483,I310452,I309915);
nor I_18093 (I309818,I310051,I310483);
nor I_18094 (I310514,I310339,I309983);
nand I_18095 (I309830,I310514,I310147);
not I_18096 (I310578,I2905);
nand I_18097 (I310595,I172886,I172880);
and I_18098 (I310612,I172886,I172880);
or I_18099 (I310629,I310612,I172904);
nand I_18100 (I310646,I310629,I310595);
and I_18101 (I310663,I310629,I172901);
and I_18102 (I310680,I310663,I172883);
or I_18103 (I310697,I172889,I172892);
nor I_18104 (I310714,I310697,I172874);
not I_18105 (I310731,I310714);
nand I_18106 (I310748,I310731,I310680);
nand I_18107 (I310765,I172877,I172907);
nor I_18108 (I310782,I310765,I172880);
not I_18109 (I310799,I310782);
nor I_18110 (I310816,I310799,I310646);
not I_18111 (I310833,I310816);
nand I_18112 (I310558,I310731,I310816);
nand I_18113 (I310552,I310680,I310799);
not I_18114 (I310878,I310765);
and I_18115 (I310895,I310878,I310646);
nand I_18116 (I310912,I310765,I310748);
DFFARX1 I_18117 (I310912,I2898,I310578,I310555,);
nor I_18118 (I310943,I172877,I172874);
not I_18119 (I310960,I172898);
nor I_18120 (I310977,I310960,I310943);
nand I_18121 (I310994,I310878,I310977);
not I_18122 (I310540,I310994);
nor I_18123 (I310543,I310714,I310994);
or I_18124 (I311039,I310782,I310977);
nor I_18125 (I310546,I310895,I311039);
nor I_18126 (I311070,I310960,I172895);
and I_18127 (I311087,I311070,I310977);
nor I_18128 (I311104,I310680,I311087);
nor I_18129 (I310564,I311104,I311087);
or I_18130 (I311135,I310731,I311104);
nor I_18131 (I311152,I311070,I310680);
nor I_18132 (I310570,I311152,I310833);
not I_18133 (I311183,I311070);
nor I_18134 (I310567,I311183,I311135);
nand I_18135 (I311214,I311183,I310646);
nor I_18136 (I310549,I310782,I311214);
nor I_18137 (I311245,I311070,I310714);
nand I_18138 (I310561,I311245,I310878);
not I_18139 (I311309,I2905);
nand I_18140 (I311326,I114128,I114149);
and I_18141 (I311343,I114128,I114149);
or I_18142 (I311360,I311343,I114125);
nand I_18143 (I311377,I311360,I311326);
and I_18144 (I311394,I311360,I114155);
and I_18145 (I311411,I311394,I114137);
or I_18146 (I311428,I114140,I114128);
nor I_18147 (I311445,I311428,I114131);
not I_18148 (I311462,I311445);
nand I_18149 (I311479,I311462,I311411);
nand I_18150 (I311496,I114143,I114125);
nor I_18151 (I311513,I311496,I114146);
not I_18152 (I311530,I311513);
nor I_18153 (I311547,I311530,I311377);
not I_18154 (I311564,I311547);
nand I_18155 (I311289,I311462,I311547);
nand I_18156 (I311283,I311411,I311530);
not I_18157 (I311609,I311496);
and I_18158 (I311626,I311609,I311377);
nand I_18159 (I311643,I311496,I311479);
DFFARX1 I_18160 (I311643,I2898,I311309,I311286,);
nor I_18161 (I311674,I114152,I114122);
not I_18162 (I311691,I114134);
nor I_18163 (I311708,I311691,I311674);
nand I_18164 (I311725,I311609,I311708);
not I_18165 (I311271,I311725);
nor I_18166 (I311274,I311445,I311725);
or I_18167 (I311770,I311513,I311708);
nor I_18168 (I311277,I311626,I311770);
nor I_18169 (I311801,I311691,I114122);
and I_18170 (I311818,I311801,I311708);
nor I_18171 (I311835,I311411,I311818);
nor I_18172 (I311295,I311835,I311818);
or I_18173 (I311866,I311462,I311835);
nor I_18174 (I311883,I311801,I311411);
nor I_18175 (I311301,I311883,I311564);
not I_18176 (I311914,I311801);
nor I_18177 (I311298,I311914,I311866);
nand I_18178 (I311945,I311914,I311377);
nor I_18179 (I311280,I311513,I311945);
nor I_18180 (I311976,I311801,I311445);
nand I_18181 (I311292,I311976,I311609);
not I_18182 (I312040,I2905);
nand I_18183 (I312057,I408103,I408118);
and I_18184 (I312074,I408103,I408118);
or I_18185 (I312091,I312074,I408109);
nand I_18186 (I312108,I312091,I312057);
and I_18187 (I312125,I312091,I408109);
and I_18188 (I312142,I312125,I408106);
or I_18189 (I312159,I408103,I408127);
nor I_18190 (I312176,I312159,I408124);
not I_18191 (I312193,I312176);
nand I_18192 (I312210,I312193,I312142);
nand I_18193 (I312227,I408121,I408115);
nor I_18194 (I312244,I312227,I408112);
not I_18195 (I312261,I312244);
nor I_18196 (I312278,I312261,I312108);
not I_18197 (I312295,I312278);
nand I_18198 (I312020,I312193,I312278);
nand I_18199 (I312014,I312142,I312261);
not I_18200 (I312340,I312227);
and I_18201 (I312357,I312340,I312108);
nand I_18202 (I312374,I312227,I312210);
DFFARX1 I_18203 (I312374,I2898,I312040,I312017,);
nor I_18204 (I312405,I408106,I408115);
not I_18205 (I312422,I408112);
nor I_18206 (I312439,I312422,I312405);
nand I_18207 (I312456,I312340,I312439);
not I_18208 (I312002,I312456);
nor I_18209 (I312005,I312176,I312456);
or I_18210 (I312501,I312244,I312439);
nor I_18211 (I312008,I312357,I312501);
nor I_18212 (I312532,I312422,I408118);
and I_18213 (I312549,I312532,I312439);
nor I_18214 (I312566,I312142,I312549);
nor I_18215 (I312026,I312566,I312549);
or I_18216 (I312597,I312193,I312566);
nor I_18217 (I312614,I312532,I312142);
nor I_18218 (I312032,I312614,I312295);
not I_18219 (I312645,I312532);
nor I_18220 (I312029,I312645,I312597);
nand I_18221 (I312676,I312645,I312108);
nor I_18222 (I312011,I312244,I312676);
nor I_18223 (I312707,I312532,I312176);
nand I_18224 (I312023,I312707,I312340);
not I_18225 (I312771,I2905);
nand I_18226 (I312788,I412217,I412223);
and I_18227 (I312805,I412217,I412223);
or I_18228 (I312822,I312805,I412223);
nand I_18229 (I312839,I312822,I312788);
and I_18230 (I312856,I312822,I412238);
and I_18231 (I312873,I312856,I412250);
or I_18232 (I312890,I412220,I412232);
nor I_18233 (I312907,I312890,I412241);
not I_18234 (I312924,I312907);
nand I_18235 (I312941,I312924,I312873);
nand I_18236 (I312958,I412247,I412229);
nor I_18237 (I312975,I312958,I412220);
not I_18238 (I312992,I312975);
nor I_18239 (I313009,I312992,I312839);
not I_18240 (I313026,I313009);
nand I_18241 (I312751,I312924,I313009);
nand I_18242 (I312745,I312873,I312992);
not I_18243 (I313071,I312958);
and I_18244 (I313088,I313071,I312839);
nand I_18245 (I313105,I312958,I312941);
DFFARX1 I_18246 (I313105,I2898,I312771,I312748,);
nor I_18247 (I313136,I412235,I412244);
not I_18248 (I313153,I412226);
nor I_18249 (I313170,I313153,I313136);
nand I_18250 (I313187,I313071,I313170);
not I_18251 (I312733,I313187);
nor I_18252 (I312736,I312907,I313187);
or I_18253 (I313232,I312975,I313170);
nor I_18254 (I312739,I313088,I313232);
nor I_18255 (I313263,I313153,I412217);
and I_18256 (I313280,I313263,I313170);
nor I_18257 (I313297,I312873,I313280);
nor I_18258 (I312757,I313297,I313280);
or I_18259 (I313328,I312924,I313297);
nor I_18260 (I313345,I313263,I312873);
nor I_18261 (I312763,I313345,I313026);
not I_18262 (I313376,I313263);
nor I_18263 (I312760,I313376,I313328);
nand I_18264 (I313407,I313376,I312839);
nor I_18265 (I312742,I312975,I313407);
nor I_18266 (I313438,I313263,I312907);
nand I_18267 (I312754,I313438,I313071);
not I_18268 (I313502,I2905);
nand I_18269 (I313519,I189045,I189042);
and I_18270 (I313536,I189045,I189042);
or I_18271 (I313553,I313536,I189030);
nand I_18272 (I313570,I313553,I313519);
and I_18273 (I313587,I313553,I189030);
and I_18274 (I313604,I313587,I189036);
or I_18275 (I313621,I189027,I189027);
nor I_18276 (I313638,I313621,I189039);
not I_18277 (I313655,I313638);
nand I_18278 (I313672,I313655,I313604);
nand I_18279 (I313689,I189048,I189033);
nor I_18280 (I313706,I313689,I189024);
not I_18281 (I313723,I313706);
nor I_18282 (I313740,I313723,I313570);
not I_18283 (I313757,I313740);
nand I_18284 (I313482,I313655,I313740);
nand I_18285 (I313476,I313604,I313723);
not I_18286 (I313802,I313689);
and I_18287 (I313819,I313802,I313570);
nand I_18288 (I313836,I313689,I313672);
DFFARX1 I_18289 (I313836,I2898,I313502,I313479,);
nor I_18290 (I313867,I189036,I189033);
not I_18291 (I313884,I189039);
nor I_18292 (I313901,I313884,I313867);
nand I_18293 (I313918,I313802,I313901);
not I_18294 (I313464,I313918);
nor I_18295 (I313467,I313638,I313918);
or I_18296 (I313963,I313706,I313901);
nor I_18297 (I313470,I313819,I313963);
nor I_18298 (I313994,I313884,I189024);
and I_18299 (I314011,I313994,I313901);
nor I_18300 (I314028,I313604,I314011);
nor I_18301 (I313488,I314028,I314011);
or I_18302 (I314059,I313655,I314028);
nor I_18303 (I314076,I313994,I313604);
nor I_18304 (I313494,I314076,I313757);
not I_18305 (I314107,I313994);
nor I_18306 (I313491,I314107,I314059);
nand I_18307 (I314138,I314107,I313570);
nor I_18308 (I313473,I313706,I314138);
nor I_18309 (I314169,I313994,I313638);
nand I_18310 (I313485,I314169,I313802);
not I_18311 (I314233,I2905);
nand I_18312 (I314250,I72033,I72057);
and I_18313 (I314267,I72033,I72057);
or I_18314 (I314284,I314267,I72045);
nand I_18315 (I314301,I314284,I314250);
and I_18316 (I314318,I314284,I72039);
and I_18317 (I314335,I314318,I72030);
or I_18318 (I314352,I72042,I72054);
nor I_18319 (I314369,I314352,I72039);
not I_18320 (I314386,I314369);
nand I_18321 (I314403,I314386,I314335);
nand I_18322 (I314420,I72036,I72048);
nor I_18323 (I314437,I314420,I72030);
not I_18324 (I314454,I314437);
nor I_18325 (I314471,I314454,I314301);
not I_18326 (I314488,I314471);
nand I_18327 (I314213,I314386,I314471);
nand I_18328 (I314207,I314335,I314454);
not I_18329 (I314533,I314420);
and I_18330 (I314550,I314533,I314301);
nand I_18331 (I314567,I314420,I314403);
DFFARX1 I_18332 (I314567,I2898,I314233,I314210,);
nor I_18333 (I314598,I72042,I72036);
not I_18334 (I314615,I72051);
nor I_18335 (I314632,I314615,I314598);
nand I_18336 (I314649,I314533,I314632);
not I_18337 (I314195,I314649);
nor I_18338 (I314198,I314369,I314649);
or I_18339 (I314694,I314437,I314632);
nor I_18340 (I314201,I314550,I314694);
nor I_18341 (I314725,I314615,I72033);
and I_18342 (I314742,I314725,I314632);
nor I_18343 (I314759,I314335,I314742);
nor I_18344 (I314219,I314759,I314742);
or I_18345 (I314790,I314386,I314759);
nor I_18346 (I314807,I314725,I314335);
nor I_18347 (I314225,I314807,I314488);
not I_18348 (I314838,I314725);
nor I_18349 (I314222,I314838,I314790);
nand I_18350 (I314869,I314838,I314301);
nor I_18351 (I314204,I314437,I314869);
nor I_18352 (I314900,I314725,I314369);
nand I_18353 (I314216,I314900,I314533);
not I_18354 (I314964,I2905);
nand I_18355 (I314981,I387434,I387440);
and I_18356 (I314998,I387434,I387440);
or I_18357 (I315015,I314998,I387464);
nand I_18358 (I315032,I315015,I314981);
and I_18359 (I315049,I315015,I387431);
and I_18360 (I315066,I315049,I387437);
or I_18361 (I315083,I387434,I387446);
nor I_18362 (I315100,I315083,I387461);
not I_18363 (I315117,I315100);
nand I_18364 (I315134,I315117,I315066);
nand I_18365 (I315151,I387452,I387449);
nor I_18366 (I315168,I315151,I387431);
not I_18367 (I315185,I315168);
nor I_18368 (I315202,I315185,I315032);
not I_18369 (I315219,I315202);
nand I_18370 (I314944,I315117,I315202);
nand I_18371 (I314938,I315066,I315185);
not I_18372 (I315264,I315151);
and I_18373 (I315281,I315264,I315032);
nand I_18374 (I315298,I315151,I315134);
DFFARX1 I_18375 (I315298,I2898,I314964,I314941,);
nor I_18376 (I315329,I387443,I387455);
not I_18377 (I315346,I387437);
nor I_18378 (I315363,I315346,I315329);
nand I_18379 (I315380,I315264,I315363);
not I_18380 (I314926,I315380);
nor I_18381 (I314929,I315100,I315380);
or I_18382 (I315425,I315168,I315363);
nor I_18383 (I314932,I315281,I315425);
nor I_18384 (I315456,I315346,I387458);
and I_18385 (I315473,I315456,I315363);
nor I_18386 (I315490,I315066,I315473);
nor I_18387 (I314950,I315490,I315473);
or I_18388 (I315521,I315117,I315490);
nor I_18389 (I315538,I315456,I315066);
nor I_18390 (I314956,I315538,I315219);
not I_18391 (I315569,I315456);
nor I_18392 (I314953,I315569,I315521);
nand I_18393 (I315600,I315569,I315032);
nor I_18394 (I314935,I315168,I315600);
nor I_18395 (I315631,I315456,I315100);
nand I_18396 (I314947,I315631,I315264);
not I_18397 (I315695,I2905);
nand I_18398 (I315712,I377098,I377104);
and I_18399 (I315729,I377098,I377104);
or I_18400 (I315746,I315729,I377128);
nand I_18401 (I315763,I315746,I315712);
and I_18402 (I315780,I315746,I377095);
and I_18403 (I315797,I315780,I377101);
or I_18404 (I315814,I377098,I377110);
nor I_18405 (I315831,I315814,I377125);
not I_18406 (I315848,I315831);
nand I_18407 (I315865,I315848,I315797);
nand I_18408 (I315882,I377116,I377113);
nor I_18409 (I315899,I315882,I377095);
not I_18410 (I315916,I315899);
nor I_18411 (I315933,I315916,I315763);
not I_18412 (I315950,I315933);
nand I_18413 (I315675,I315848,I315933);
nand I_18414 (I315669,I315797,I315916);
not I_18415 (I315995,I315882);
and I_18416 (I316012,I315995,I315763);
nand I_18417 (I316029,I315882,I315865);
DFFARX1 I_18418 (I316029,I2898,I315695,I315672,);
nor I_18419 (I316060,I377107,I377119);
not I_18420 (I316077,I377101);
nor I_18421 (I316094,I316077,I316060);
nand I_18422 (I316111,I315995,I316094);
not I_18423 (I315657,I316111);
nor I_18424 (I315660,I315831,I316111);
or I_18425 (I316156,I315899,I316094);
nor I_18426 (I315663,I316012,I316156);
nor I_18427 (I316187,I316077,I377122);
and I_18428 (I316204,I316187,I316094);
nor I_18429 (I316221,I315797,I316204);
nor I_18430 (I315681,I316221,I316204);
or I_18431 (I316252,I315848,I316221);
nor I_18432 (I316269,I316187,I315797);
nor I_18433 (I315687,I316269,I315950);
not I_18434 (I316300,I316187);
nor I_18435 (I315684,I316300,I316252);
nand I_18436 (I316331,I316300,I315763);
nor I_18437 (I315666,I315899,I316331);
nor I_18438 (I316362,I316187,I315831);
nand I_18439 (I315678,I316362,I315995);
not I_18440 (I316426,I2905);
nand I_18441 (I316443,I118531,I118552);
and I_18442 (I316460,I118531,I118552);
or I_18443 (I316477,I316460,I118528);
nand I_18444 (I316494,I316477,I316443);
and I_18445 (I316511,I316477,I118558);
and I_18446 (I316528,I316511,I118540);
or I_18447 (I316545,I118543,I118531);
nor I_18448 (I316562,I316545,I118534);
not I_18449 (I316579,I316562);
nand I_18450 (I316596,I316579,I316528);
nand I_18451 (I316613,I118546,I118528);
nor I_18452 (I316630,I316613,I118549);
not I_18453 (I316647,I316630);
nor I_18454 (I316664,I316647,I316494);
not I_18455 (I316681,I316664);
nand I_18456 (I316406,I316579,I316664);
nand I_18457 (I316400,I316528,I316647);
not I_18458 (I316726,I316613);
and I_18459 (I316743,I316726,I316494);
nand I_18460 (I316760,I316613,I316596);
DFFARX1 I_18461 (I316760,I2898,I316426,I316403,);
nor I_18462 (I316791,I118555,I118525);
not I_18463 (I316808,I118537);
nor I_18464 (I316825,I316808,I316791);
nand I_18465 (I316842,I316726,I316825);
not I_18466 (I316388,I316842);
nor I_18467 (I316391,I316562,I316842);
or I_18468 (I316887,I316630,I316825);
nor I_18469 (I316394,I316743,I316887);
nor I_18470 (I316918,I316808,I118525);
and I_18471 (I316935,I316918,I316825);
nor I_18472 (I316952,I316528,I316935);
nor I_18473 (I316412,I316952,I316935);
or I_18474 (I316983,I316579,I316952);
nor I_18475 (I317000,I316918,I316528);
nor I_18476 (I316418,I317000,I316681);
not I_18477 (I317031,I316918);
nor I_18478 (I316415,I317031,I316983);
nand I_18479 (I317062,I317031,I316494);
nor I_18480 (I316397,I316630,I317062);
nor I_18481 (I317093,I316918,I316562);
nand I_18482 (I316409,I317093,I316726);
not I_18483 (I317157,I2905);
nand I_18484 (I317174,I83984,I84008);
and I_18485 (I317191,I83984,I84008);
or I_18486 (I317208,I317191,I83996);
nand I_18487 (I317225,I317208,I317174);
and I_18488 (I317242,I317208,I83990);
and I_18489 (I317259,I317242,I83981);
or I_18490 (I317276,I83993,I84005);
nor I_18491 (I317293,I317276,I83990);
not I_18492 (I317310,I317293);
nand I_18493 (I317327,I317310,I317259);
nand I_18494 (I317344,I83987,I83999);
nor I_18495 (I317361,I317344,I83981);
not I_18496 (I317378,I317361);
nor I_18497 (I317395,I317378,I317225);
not I_18498 (I317412,I317395);
nand I_18499 (I317137,I317310,I317395);
nand I_18500 (I317131,I317259,I317378);
not I_18501 (I317457,I317344);
and I_18502 (I317474,I317457,I317225);
nand I_18503 (I317491,I317344,I317327);
DFFARX1 I_18504 (I317491,I2898,I317157,I317134,);
nor I_18505 (I317522,I83993,I83987);
not I_18506 (I317539,I84002);
nor I_18507 (I317556,I317539,I317522);
nand I_18508 (I317573,I317457,I317556);
not I_18509 (I317119,I317573);
nor I_18510 (I317122,I317293,I317573);
or I_18511 (I317618,I317361,I317556);
nor I_18512 (I317125,I317474,I317618);
nor I_18513 (I317649,I317539,I83984);
and I_18514 (I317666,I317649,I317556);
nor I_18515 (I317683,I317259,I317666);
nor I_18516 (I317143,I317683,I317666);
or I_18517 (I317714,I317310,I317683);
nor I_18518 (I317731,I317649,I317259);
nor I_18519 (I317149,I317731,I317412);
not I_18520 (I317762,I317649);
nor I_18521 (I317146,I317762,I317714);
nand I_18522 (I317793,I317762,I317225);
nor I_18523 (I317128,I317361,I317793);
nor I_18524 (I317824,I317649,I317293);
nand I_18525 (I317140,I317824,I317457);
not I_18526 (I317888,I2905);
nand I_18527 (I317905,I174926,I174920);
and I_18528 (I317922,I174926,I174920);
or I_18529 (I317939,I317922,I174944);
nand I_18530 (I317956,I317939,I317905);
and I_18531 (I317973,I317939,I174941);
and I_18532 (I317990,I317973,I174923);
or I_18533 (I318007,I174929,I174932);
nor I_18534 (I318024,I318007,I174914);
not I_18535 (I318041,I318024);
nand I_18536 (I318058,I318041,I317990);
nand I_18537 (I318075,I174917,I174947);
nor I_18538 (I318092,I318075,I174920);
not I_18539 (I318109,I318092);
nor I_18540 (I318126,I318109,I317956);
not I_18541 (I318143,I318126);
nand I_18542 (I317868,I318041,I318126);
nand I_18543 (I317862,I317990,I318109);
not I_18544 (I318188,I318075);
and I_18545 (I318205,I318188,I317956);
nand I_18546 (I318222,I318075,I318058);
DFFARX1 I_18547 (I318222,I2898,I317888,I317865,);
nor I_18548 (I318253,I174917,I174914);
not I_18549 (I318270,I174938);
nor I_18550 (I318287,I318270,I318253);
nand I_18551 (I318304,I318188,I318287);
not I_18552 (I317850,I318304);
nor I_18553 (I317853,I318024,I318304);
or I_18554 (I318349,I318092,I318287);
nor I_18555 (I317856,I318205,I318349);
nor I_18556 (I318380,I318270,I174935);
and I_18557 (I318397,I318380,I318287);
nor I_18558 (I318414,I317990,I318397);
nor I_18559 (I317874,I318414,I318397);
or I_18560 (I318445,I318041,I318414);
nor I_18561 (I318462,I318380,I317990);
nor I_18562 (I317880,I318462,I318143);
not I_18563 (I318493,I318380);
nor I_18564 (I317877,I318493,I318445);
nand I_18565 (I318524,I318493,I317956);
nor I_18566 (I317859,I318092,I318524);
nor I_18567 (I318555,I318380,I318024);
nand I_18568 (I317871,I318555,I318188);
not I_18569 (I318619,I2905);
nand I_18570 (I318636,I418490,I418496);
and I_18571 (I318653,I418490,I418496);
or I_18572 (I318670,I318653,I418496);
nand I_18573 (I318687,I318670,I318636);
and I_18574 (I318704,I318670,I418511);
and I_18575 (I318721,I318704,I418523);
or I_18576 (I318738,I418493,I418505);
nor I_18577 (I318755,I318738,I418514);
not I_18578 (I318772,I318755);
nand I_18579 (I318789,I318772,I318721);
nand I_18580 (I318806,I418520,I418502);
nor I_18581 (I318823,I318806,I418493);
not I_18582 (I318840,I318823);
nor I_18583 (I318857,I318840,I318687);
not I_18584 (I318874,I318857);
nand I_18585 (I318599,I318772,I318857);
nand I_18586 (I318593,I318721,I318840);
not I_18587 (I318919,I318806);
and I_18588 (I318936,I318919,I318687);
nand I_18589 (I318953,I318806,I318789);
DFFARX1 I_18590 (I318953,I2898,I318619,I318596,);
nor I_18591 (I318984,I418508,I418517);
not I_18592 (I319001,I418499);
nor I_18593 (I319018,I319001,I318984);
nand I_18594 (I319035,I318919,I319018);
not I_18595 (I318581,I319035);
nor I_18596 (I318584,I318755,I319035);
or I_18597 (I319080,I318823,I319018);
nor I_18598 (I318587,I318936,I319080);
nor I_18599 (I319111,I319001,I418490);
and I_18600 (I319128,I319111,I319018);
nor I_18601 (I319145,I318721,I319128);
nor I_18602 (I318605,I319145,I319128);
or I_18603 (I319176,I318772,I319145);
nor I_18604 (I319193,I319111,I318721);
nor I_18605 (I318611,I319193,I318874);
not I_18606 (I319224,I319111);
nor I_18607 (I318608,I319224,I319176);
nand I_18608 (I319255,I319224,I318687);
nor I_18609 (I318590,I318823,I319255);
nor I_18610 (I319286,I319111,I318755);
nand I_18611 (I318602,I319286,I318919);
not I_18612 (I319350,I2905);
nand I_18613 (I319367,I431733,I431739);
and I_18614 (I319384,I431733,I431739);
or I_18615 (I319401,I319384,I431739);
nand I_18616 (I319418,I319401,I319367);
and I_18617 (I319435,I319401,I431754);
and I_18618 (I319452,I319435,I431766);
or I_18619 (I319469,I431736,I431748);
nor I_18620 (I319486,I319469,I431757);
not I_18621 (I319503,I319486);
nand I_18622 (I319520,I319503,I319452);
nand I_18623 (I319537,I431763,I431745);
nor I_18624 (I319554,I319537,I431736);
not I_18625 (I319571,I319554);
nor I_18626 (I319588,I319571,I319418);
not I_18627 (I319605,I319588);
nand I_18628 (I319330,I319503,I319588);
nand I_18629 (I319324,I319452,I319571);
not I_18630 (I319650,I319537);
and I_18631 (I319667,I319650,I319418);
nand I_18632 (I319684,I319537,I319520);
DFFARX1 I_18633 (I319684,I2898,I319350,I319327,);
nor I_18634 (I319715,I431751,I431760);
not I_18635 (I319732,I431742);
nor I_18636 (I319749,I319732,I319715);
nand I_18637 (I319766,I319650,I319749);
not I_18638 (I319312,I319766);
nor I_18639 (I319315,I319486,I319766);
or I_18640 (I319811,I319554,I319749);
nor I_18641 (I319318,I319667,I319811);
nor I_18642 (I319842,I319732,I431733);
and I_18643 (I319859,I319842,I319749);
nor I_18644 (I319876,I319452,I319859);
nor I_18645 (I319336,I319876,I319859);
or I_18646 (I319907,I319503,I319876);
nor I_18647 (I319924,I319842,I319452);
nor I_18648 (I319342,I319924,I319605);
not I_18649 (I319955,I319842);
nor I_18650 (I319339,I319955,I319907);
nand I_18651 (I319986,I319955,I319418);
nor I_18652 (I319321,I319554,I319986);
nor I_18653 (I320017,I319842,I319486);
nand I_18654 (I319333,I320017,I319650);
not I_18655 (I320081,I2905);
nand I_18656 (I320098,I144326,I144320);
and I_18657 (I320115,I144326,I144320);
or I_18658 (I320132,I320115,I144344);
nand I_18659 (I320149,I320132,I320098);
and I_18660 (I320166,I320132,I144341);
and I_18661 (I320183,I320166,I144323);
or I_18662 (I320200,I144329,I144332);
nor I_18663 (I320217,I320200,I144314);
not I_18664 (I320234,I320217);
nand I_18665 (I320251,I320234,I320183);
nand I_18666 (I320268,I144317,I144347);
nor I_18667 (I320285,I320268,I144320);
not I_18668 (I320302,I320285);
nor I_18669 (I320319,I320302,I320149);
not I_18670 (I320336,I320319);
nand I_18671 (I320061,I320234,I320319);
nand I_18672 (I320055,I320183,I320302);
not I_18673 (I320381,I320268);
and I_18674 (I320398,I320381,I320149);
nand I_18675 (I320415,I320268,I320251);
DFFARX1 I_18676 (I320415,I2898,I320081,I320058,);
nor I_18677 (I320446,I144317,I144314);
not I_18678 (I320463,I144338);
nor I_18679 (I320480,I320463,I320446);
nand I_18680 (I320497,I320381,I320480);
not I_18681 (I320043,I320497);
nor I_18682 (I320046,I320217,I320497);
or I_18683 (I320542,I320285,I320480);
nor I_18684 (I320049,I320398,I320542);
nor I_18685 (I320573,I320463,I144335);
and I_18686 (I320590,I320573,I320480);
nor I_18687 (I320607,I320183,I320590);
nor I_18688 (I320067,I320607,I320590);
or I_18689 (I320638,I320234,I320607);
nor I_18690 (I320655,I320573,I320183);
nor I_18691 (I320073,I320655,I320336);
not I_18692 (I320686,I320573);
nor I_18693 (I320070,I320686,I320638);
nand I_18694 (I320717,I320686,I320149);
nor I_18695 (I320052,I320285,I320717);
nor I_18696 (I320748,I320573,I320217);
nand I_18697 (I320064,I320748,I320381);
not I_18698 (I320812,I2905);
nand I_18699 (I320829,I1683,I1923);
and I_18700 (I320846,I1683,I1923);
or I_18701 (I320863,I320846,I1939);
nand I_18702 (I320880,I320863,I320829);
and I_18703 (I320897,I320863,I2803);
and I_18704 (I320914,I320897,I1787);
or I_18705 (I320931,I2539,I1603);
nor I_18706 (I320948,I320931,I2315);
not I_18707 (I320965,I320948);
nand I_18708 (I320982,I320965,I320914);
nand I_18709 (I320999,I2451,I2019);
nor I_18710 (I321016,I320999,I2787);
not I_18711 (I321033,I321016);
nor I_18712 (I321050,I321033,I320880);
not I_18713 (I321067,I321050);
nand I_18714 (I320792,I320965,I321050);
nand I_18715 (I320786,I320914,I321033);
not I_18716 (I321112,I320999);
and I_18717 (I321129,I321112,I320880);
nand I_18718 (I321146,I320999,I320982);
DFFARX1 I_18719 (I321146,I2898,I320812,I320789,);
nor I_18720 (I321177,I1971,I1883);
not I_18721 (I321194,I2355);
nor I_18722 (I321211,I321194,I321177);
nand I_18723 (I321228,I321112,I321211);
not I_18724 (I320774,I321228);
nor I_18725 (I320777,I320948,I321228);
or I_18726 (I321273,I321016,I321211);
nor I_18727 (I320780,I321129,I321273);
nor I_18728 (I321304,I321194,I2387);
and I_18729 (I321321,I321304,I321211);
nor I_18730 (I321338,I320914,I321321);
nor I_18731 (I320798,I321338,I321321);
or I_18732 (I321369,I320965,I321338);
nor I_18733 (I321386,I321304,I320914);
nor I_18734 (I320804,I321386,I321067);
not I_18735 (I321417,I321304);
nor I_18736 (I320801,I321417,I321369);
nand I_18737 (I321448,I321417,I320880);
nor I_18738 (I320783,I321016,I321448);
nor I_18739 (I321479,I321304,I320948);
nand I_18740 (I320795,I321479,I321112);
not I_18741 (I321543,I2905);
nand I_18742 (I321560,I61969,I61993);
and I_18743 (I321577,I61969,I61993);
or I_18744 (I321594,I321577,I61981);
nand I_18745 (I321611,I321594,I321560);
and I_18746 (I321628,I321594,I61975);
and I_18747 (I321645,I321628,I61966);
or I_18748 (I321662,I61978,I61990);
nor I_18749 (I321679,I321662,I61975);
not I_18750 (I321696,I321679);
nand I_18751 (I321713,I321696,I321645);
nand I_18752 (I321730,I61972,I61984);
nor I_18753 (I321747,I321730,I61966);
not I_18754 (I321764,I321747);
nor I_18755 (I321781,I321764,I321611);
not I_18756 (I321798,I321781);
nand I_18757 (I321523,I321696,I321781);
nand I_18758 (I321517,I321645,I321764);
not I_18759 (I321843,I321730);
and I_18760 (I321860,I321843,I321611);
nand I_18761 (I321877,I321730,I321713);
DFFARX1 I_18762 (I321877,I2898,I321543,I321520,);
nor I_18763 (I321908,I61978,I61972);
not I_18764 (I321925,I61987);
nor I_18765 (I321942,I321925,I321908);
nand I_18766 (I321959,I321843,I321942);
not I_18767 (I321505,I321959);
nor I_18768 (I321508,I321679,I321959);
or I_18769 (I322004,I321747,I321942);
nor I_18770 (I321511,I321860,I322004);
nor I_18771 (I322035,I321925,I61969);
and I_18772 (I322052,I322035,I321942);
nor I_18773 (I322069,I321645,I322052);
nor I_18774 (I321529,I322069,I322052);
or I_18775 (I322100,I321696,I322069);
nor I_18776 (I322117,I322035,I321645);
nor I_18777 (I321535,I322117,I321798);
not I_18778 (I322148,I322035);
nor I_18779 (I321532,I322148,I322100);
nand I_18780 (I322179,I322148,I321611);
nor I_18781 (I321514,I321747,I322179);
nor I_18782 (I322210,I322035,I321679);
nand I_18783 (I321526,I322210,I321843);
not I_18784 (I322268,I2905);
or I_18785 (I322285,I135511,I135517);
nand I_18786 (I322302,I135529,I135520);
not I_18787 (I322319,I322302);
nand I_18788 (I322336,I322319,I322285);
or I_18789 (I322353,I135526,I135508);
nor I_18790 (I322370,I322353,I135541);
nand I_18791 (I322387,I322319,I322370);
nor I_18792 (I322404,I322370,I322302);
not I_18793 (I322421,I322404);
not I_18794 (I322438,I322370);
nand I_18795 (I322257,I322336,I322438);
nor I_18796 (I322469,I135511,I135514);
nor I_18797 (I322486,I322469,I135523);
nor I_18798 (I322503,I322486,I322302);
nor I_18799 (I322520,I322438,I322486);
nor I_18800 (I322537,I135532,I135514);
nand I_18801 (I322554,I322537,I322503);
not I_18802 (I322571,I322554);
nor I_18803 (I322242,I322336,I322571);
nand I_18804 (I322239,I322554,I322387);
nand I_18805 (I322616,I322520,I322537);
nand I_18806 (I322260,I322554,I322616);
nand I_18807 (I322647,I135538,I135535);
not I_18808 (I322664,I322647);
nor I_18809 (I322236,I322664,I322302);
nor I_18810 (I322695,I322647,I135508);
not I_18811 (I322712,I322695);
nor I_18812 (I322245,I322336,I322712);
nand I_18813 (I322743,I322438,I322712);
nand I_18814 (I322254,I322421,I322743);
nor I_18815 (I322251,I322319,I322695);
nand I_18816 (I322788,I322647,I322336);
not I_18817 (I322805,I322788);
DFFARX1 I_18818 (I322805,I2898,I322268,I322248,);
not I_18819 (I322863,I2905);
or I_18820 (I322880,I309815,I309827);
nand I_18821 (I322897,I309833,I309830);
not I_18822 (I322914,I322897);
nand I_18823 (I322931,I322914,I322880);
or I_18824 (I322948,I309824,I309809);
nor I_18825 (I322965,I322948,I309839);
nand I_18826 (I322982,I322914,I322965);
nor I_18827 (I322999,I322965,I322897);
not I_18828 (I323016,I322999);
not I_18829 (I323033,I322965);
nand I_18830 (I322852,I322931,I323033);
nor I_18831 (I323064,I309836,I309818);
nor I_18832 (I323081,I323064,I309812);
nor I_18833 (I323098,I323081,I322897);
nor I_18834 (I323115,I323033,I323081);
nor I_18835 (I323132,I309815,I309818);
nand I_18836 (I323149,I323132,I323098);
not I_18837 (I323166,I323149);
nor I_18838 (I322837,I322931,I323166);
nand I_18839 (I322834,I323149,I322982);
nand I_18840 (I323211,I323115,I323132);
nand I_18841 (I322855,I323149,I323211);
nand I_18842 (I323242,I309809,I309821);
not I_18843 (I323259,I323242);
nor I_18844 (I322831,I323259,I322897);
nor I_18845 (I323290,I323242,I309812);
not I_18846 (I323307,I323290);
nor I_18847 (I322840,I322931,I323307);
nand I_18848 (I323338,I323033,I323307);
nand I_18849 (I322849,I323016,I323338);
nor I_18850 (I322846,I322914,I323290);
nand I_18851 (I323383,I323242,I322931);
not I_18852 (I323400,I323383);
DFFARX1 I_18853 (I323400,I2898,I322863,I322843,);
not I_18854 (I323458,I2905);
or I_18855 (I323475,I284217,I284196);
nand I_18856 (I323492,I284193,I284208);
not I_18857 (I323509,I323492);
nand I_18858 (I323526,I323509,I323475);
or I_18859 (I323543,I284205,I284196);
nor I_18860 (I323560,I323543,I284202);
nand I_18861 (I323577,I323509,I323560);
nor I_18862 (I323594,I323560,I323492);
not I_18863 (I323611,I323594);
not I_18864 (I323628,I323560);
nand I_18865 (I323447,I323526,I323628);
nor I_18866 (I323659,I284199,I284199);
nor I_18867 (I323676,I323659,I284220);
nor I_18868 (I323693,I323676,I323492);
nor I_18869 (I323710,I323628,I323676);
nor I_18870 (I323727,I284190,I284211);
nand I_18871 (I323744,I323727,I323693);
not I_18872 (I323761,I323744);
nor I_18873 (I323432,I323526,I323761);
nand I_18874 (I323429,I323744,I323577);
nand I_18875 (I323806,I323710,I323727);
nand I_18876 (I323450,I323744,I323806);
nand I_18877 (I323837,I284193,I284214);
not I_18878 (I323854,I323837);
nor I_18879 (I323426,I323854,I323492);
nor I_18880 (I323885,I323837,I284190);
not I_18881 (I323902,I323885);
nor I_18882 (I323435,I323526,I323902);
nand I_18883 (I323933,I323628,I323902);
nand I_18884 (I323444,I323611,I323933);
nor I_18885 (I323441,I323509,I323885);
nand I_18886 (I323978,I323837,I323526);
not I_18887 (I323995,I323978);
DFFARX1 I_18888 (I323995,I2898,I323458,I323438,);
not I_18889 (I324053,I2905);
or I_18890 (I324070,I170175,I170154);
nand I_18891 (I324087,I170160,I170178);
not I_18892 (I324104,I324087);
nand I_18893 (I324121,I324104,I324070);
or I_18894 (I324138,I170154,I170169);
nor I_18895 (I324155,I324138,I170166);
nand I_18896 (I324172,I324104,I324155);
nor I_18897 (I324189,I324155,I324087);
not I_18898 (I324206,I324189);
not I_18899 (I324223,I324155);
nand I_18900 (I324042,I324121,I324223);
nor I_18901 (I324254,I170172,I170184);
nor I_18902 (I324271,I324254,I170157);
nor I_18903 (I324288,I324271,I324087);
nor I_18904 (I324305,I324223,I324271);
nor I_18905 (I324322,I170163,I170181);
nand I_18906 (I324339,I324322,I324288);
not I_18907 (I324356,I324339);
nor I_18908 (I324027,I324121,I324356);
nand I_18909 (I324024,I324339,I324172);
nand I_18910 (I324401,I324305,I324322);
nand I_18911 (I324045,I324339,I324401);
nand I_18912 (I324432,I170157,I170187);
not I_18913 (I324449,I324432);
nor I_18914 (I324021,I324449,I324087);
nor I_18915 (I324480,I324432,I170160);
not I_18916 (I324497,I324480);
nor I_18917 (I324030,I324121,I324497);
nand I_18918 (I324528,I324223,I324497);
nand I_18919 (I324039,I324206,I324528);
nor I_18920 (I324036,I324104,I324480);
nand I_18921 (I324573,I324432,I324121);
not I_18922 (I324590,I324573);
DFFARX1 I_18923 (I324590,I2898,I324053,I324033,);
not I_18924 (I324648,I2905);
or I_18925 (I324665,I103432,I103438);
nand I_18926 (I324682,I103450,I103441);
not I_18927 (I324699,I324682);
nand I_18928 (I324716,I324699,I324665);
or I_18929 (I324733,I103447,I103429);
nor I_18930 (I324750,I324733,I103462);
nand I_18931 (I324767,I324699,I324750);
nor I_18932 (I324784,I324750,I324682);
not I_18933 (I324801,I324784);
not I_18934 (I324818,I324750);
nand I_18935 (I324637,I324716,I324818);
nor I_18936 (I324849,I103432,I103435);
nor I_18937 (I324866,I324849,I103444);
nor I_18938 (I324883,I324866,I324682);
nor I_18939 (I324900,I324818,I324866);
nor I_18940 (I324917,I103453,I103435);
nand I_18941 (I324934,I324917,I324883);
not I_18942 (I324951,I324934);
nor I_18943 (I324622,I324716,I324951);
nand I_18944 (I324619,I324934,I324767);
nand I_18945 (I324996,I324900,I324917);
nand I_18946 (I324640,I324934,I324996);
nand I_18947 (I325027,I103459,I103456);
not I_18948 (I325044,I325027);
nor I_18949 (I324616,I325044,I324682);
nor I_18950 (I325075,I325027,I103429);
not I_18951 (I325092,I325075);
nor I_18952 (I324625,I324716,I325092);
nand I_18953 (I325123,I324818,I325092);
nand I_18954 (I324634,I324801,I325123);
nor I_18955 (I324631,I324699,I325075);
nand I_18956 (I325168,I325027,I324716);
not I_18957 (I325185,I325168);
DFFARX1 I_18958 (I325185,I2898,I324648,I324628,);
not I_18959 (I325243,I2905);
or I_18960 (I325260,I77718,I77691);
nand I_18961 (I325277,I77703,I77697);
not I_18962 (I325294,I325277);
nand I_18963 (I325311,I325294,I325260);
or I_18964 (I325328,I77700,I77715);
nor I_18965 (I325345,I325328,I77694);
nand I_18966 (I325362,I325294,I325345);
nor I_18967 (I325379,I325345,I325277);
not I_18968 (I325396,I325379);
not I_18969 (I325413,I325345);
nand I_18970 (I325232,I325311,I325413);
nor I_18971 (I325444,I77712,I77694);
nor I_18972 (I325461,I325444,I77700);
nor I_18973 (I325478,I325461,I325277);
nor I_18974 (I325495,I325413,I325461);
nor I_18975 (I325512,I77691,I77709);
nand I_18976 (I325529,I325512,I325478);
not I_18977 (I325546,I325529);
nor I_18978 (I325217,I325311,I325546);
nand I_18979 (I325214,I325529,I325362);
nand I_18980 (I325591,I325495,I325512);
nand I_18981 (I325235,I325529,I325591);
nand I_18982 (I325622,I77697,I77706);
not I_18983 (I325639,I325622);
nor I_18984 (I325211,I325639,I325277);
nor I_18985 (I325670,I325622,I77703);
not I_18986 (I325687,I325670);
nor I_18987 (I325220,I325311,I325687);
nand I_18988 (I325718,I325413,I325687);
nand I_18989 (I325229,I325396,I325718);
nor I_18990 (I325226,I325294,I325670);
nand I_18991 (I325763,I325622,I325311);
not I_18992 (I325780,I325763);
DFFARX1 I_18993 (I325780,I2898,I325243,I325223,);
not I_18994 (I325838,I2905);
or I_18995 (I325855,I171535,I171514);
nand I_18996 (I325872,I171520,I171538);
not I_18997 (I325889,I325872);
nand I_18998 (I325906,I325889,I325855);
or I_18999 (I325923,I171514,I171529);
nor I_19000 (I325940,I325923,I171526);
nand I_19001 (I325957,I325889,I325940);
nor I_19002 (I325974,I325940,I325872);
not I_19003 (I325991,I325974);
not I_19004 (I326008,I325940);
nand I_19005 (I325827,I325906,I326008);
nor I_19006 (I326039,I171532,I171544);
nor I_19007 (I326056,I326039,I171517);
nor I_19008 (I326073,I326056,I325872);
nor I_19009 (I326090,I326008,I326056);
nor I_19010 (I326107,I171523,I171541);
nand I_19011 (I326124,I326107,I326073);
not I_19012 (I326141,I326124);
nor I_19013 (I325812,I325906,I326141);
nand I_19014 (I325809,I326124,I325957);
nand I_19015 (I326186,I326090,I326107);
nand I_19016 (I325830,I326124,I326186);
nand I_19017 (I326217,I171517,I171547);
not I_19018 (I326234,I326217);
nor I_19019 (I325806,I326234,I325872);
nor I_19020 (I326265,I326217,I171520);
not I_19021 (I326282,I326265);
nor I_19022 (I325815,I325906,I326282);
nand I_19023 (I326313,I326008,I326282);
nand I_19024 (I325824,I325991,I326313);
nor I_19025 (I325821,I325889,I326265);
nand I_19026 (I326358,I326217,I325906);
not I_19027 (I326375,I326358);
DFFARX1 I_19028 (I326375,I2898,I325838,I325818,);
not I_19029 (I326433,I2905);
or I_19030 (I326450,I402004,I402001);
nand I_19031 (I326467,I401992,I401989);
not I_19032 (I326484,I326467);
nand I_19033 (I326501,I326484,I326450);
or I_19034 (I326518,I401986,I401998);
nor I_19035 (I326535,I326518,I401989);
nand I_19036 (I326552,I326484,I326535);
nor I_19037 (I326569,I326535,I326467);
not I_19038 (I326586,I326569);
not I_19039 (I326603,I326535);
nand I_19040 (I326422,I326501,I326603);
nor I_19041 (I326634,I401986,I401992);
nor I_19042 (I326651,I326634,I401998);
nor I_19043 (I326668,I326651,I326467);
nor I_19044 (I326685,I326603,I326651);
nor I_19045 (I326702,I401983,I401983);
nand I_19046 (I326719,I326702,I326668);
not I_19047 (I326736,I326719);
nor I_19048 (I326407,I326501,I326736);
nand I_19049 (I326404,I326719,I326552);
nand I_19050 (I326781,I326685,I326702);
nand I_19051 (I326425,I326719,I326781);
nand I_19052 (I326812,I401995,I402007);
not I_19053 (I326829,I326812);
nor I_19054 (I326401,I326829,I326467);
nor I_19055 (I326860,I326812,I401995);
not I_19056 (I326877,I326860);
nor I_19057 (I326410,I326501,I326877);
nand I_19058 (I326908,I326603,I326877);
nand I_19059 (I326419,I326586,I326908);
nor I_19060 (I326416,I326484,I326860);
nand I_19061 (I326953,I326812,I326501);
not I_19062 (I326970,I326953);
DFFARX1 I_19063 (I326970,I2898,I326433,I326413,);
not I_19064 (I327028,I2905);
or I_19065 (I327045,I98434,I98449);
nand I_19066 (I327062,I98446,I98431);
not I_19067 (I327079,I327062);
nand I_19068 (I327096,I327079,I327045);
or I_19069 (I327113,I98440,I98431);
nor I_19070 (I327130,I327113,I98437);
nand I_19071 (I327147,I327079,I327130);
nor I_19072 (I327164,I327130,I327062);
not I_19073 (I327181,I327164);
not I_19074 (I327198,I327130);
nand I_19075 (I327017,I327096,I327198);
nor I_19076 (I327229,I98437,I98443);
nor I_19077 (I327246,I327229,I98455);
nor I_19078 (I327263,I327246,I327062);
nor I_19079 (I327280,I327198,I327246);
nor I_19080 (I327297,I98452,I98434);
nand I_19081 (I327314,I327297,I327263);
not I_19082 (I327331,I327314);
nor I_19083 (I327002,I327096,I327331);
nand I_19084 (I326999,I327314,I327147);
nand I_19085 (I327376,I327280,I327297);
nand I_19086 (I327020,I327314,I327376);
nand I_19087 (I327407,I98443,I98440);
not I_19088 (I327424,I327407);
nor I_19089 (I326996,I327424,I327062);
nor I_19090 (I327455,I327407,I98446);
not I_19091 (I327472,I327455);
nor I_19092 (I327005,I327096,I327472);
nand I_19093 (I327503,I327198,I327472);
nand I_19094 (I327014,I327181,I327503);
nor I_19095 (I327011,I327079,I327455);
nand I_19096 (I327548,I327407,I327096);
not I_19097 (I327565,I327548);
DFFARX1 I_19098 (I327565,I2898,I327028,I327008,);
not I_19099 (I327623,I2905);
or I_19100 (I327640,I248262,I248241);
nand I_19101 (I327657,I248238,I248253);
not I_19102 (I327674,I327657);
nand I_19103 (I327691,I327674,I327640);
or I_19104 (I327708,I248250,I248241);
nor I_19105 (I327725,I327708,I248247);
nand I_19106 (I327742,I327674,I327725);
nor I_19107 (I327759,I327725,I327657);
not I_19108 (I327776,I327759);
not I_19109 (I327793,I327725);
nand I_19110 (I327612,I327691,I327793);
nor I_19111 (I327824,I248244,I248244);
nor I_19112 (I327841,I327824,I248265);
nor I_19113 (I327858,I327841,I327657);
nor I_19114 (I327875,I327793,I327841);
nor I_19115 (I327892,I248235,I248256);
nand I_19116 (I327909,I327892,I327858);
not I_19117 (I327926,I327909);
nor I_19118 (I327597,I327691,I327926);
nand I_19119 (I327594,I327909,I327742);
nand I_19120 (I327971,I327875,I327892);
nand I_19121 (I327615,I327909,I327971);
nand I_19122 (I328002,I248238,I248259);
not I_19123 (I328019,I328002);
nor I_19124 (I327591,I328019,I327657);
nor I_19125 (I328050,I328002,I248235);
not I_19126 (I328067,I328050);
nor I_19127 (I327600,I327691,I328067);
nand I_19128 (I328098,I327793,I328067);
nand I_19129 (I327609,I327776,I328098);
nor I_19130 (I327606,I327674,I328050);
nand I_19131 (I328143,I328002,I327691);
not I_19132 (I328160,I328143);
DFFARX1 I_19133 (I328160,I2898,I327623,I327603,);
not I_19134 (I328218,I2905);
or I_19135 (I328235,I202976,I202979);
nand I_19136 (I328252,I202985,I202976);
not I_19137 (I328269,I328252);
nand I_19138 (I328286,I328269,I328235);
or I_19139 (I328303,I202967,I202967);
nor I_19140 (I328320,I328303,I202964);
nand I_19141 (I328337,I328269,I328320);
nor I_19142 (I328354,I328320,I328252);
not I_19143 (I328371,I328354);
not I_19144 (I328388,I328320);
nand I_19145 (I328207,I328286,I328388);
nor I_19146 (I328419,I202973,I202970);
nor I_19147 (I328436,I328419,I202982);
nor I_19148 (I328453,I328436,I328252);
nor I_19149 (I328470,I328388,I328436);
nor I_19150 (I328487,I202991,I202964);
nand I_19151 (I328504,I328487,I328453);
not I_19152 (I328521,I328504);
nor I_19153 (I328192,I328286,I328521);
nand I_19154 (I328189,I328504,I328337);
nand I_19155 (I328566,I328470,I328487);
nand I_19156 (I328210,I328504,I328566);
nand I_19157 (I328597,I202970,I202973);
not I_19158 (I328614,I328597);
nor I_19159 (I328186,I328614,I328252);
nor I_19160 (I328645,I328597,I202988);
not I_19161 (I328662,I328645);
nor I_19162 (I328195,I328286,I328662);
nand I_19163 (I328693,I328388,I328662);
nand I_19164 (I328204,I328371,I328693);
nor I_19165 (I328201,I328269,I328645);
nand I_19166 (I328738,I328597,I328286);
not I_19167 (I328755,I328738);
DFFARX1 I_19168 (I328755,I2898,I328218,I328198,);
not I_19169 (I328813,I2905);
or I_19170 (I328830,I388107,I388104);
nand I_19171 (I328847,I388089,I388083);
not I_19172 (I328864,I328847);
nand I_19173 (I328881,I328864,I328830);
or I_19174 (I328898,I388110,I388077);
nor I_19175 (I328915,I328898,I388083);
nand I_19176 (I328932,I328864,I328915);
nor I_19177 (I328949,I328915,I328847);
not I_19178 (I328966,I328949);
not I_19179 (I328983,I328915);
nand I_19180 (I328802,I328881,I328983);
nor I_19181 (I329014,I388101,I388092);
nor I_19182 (I329031,I329014,I388095);
nor I_19183 (I329048,I329031,I328847);
nor I_19184 (I329065,I328983,I329031);
nor I_19185 (I329082,I388098,I388080);
nand I_19186 (I329099,I329082,I329048);
not I_19187 (I329116,I329099);
nor I_19188 (I328787,I328881,I329116);
nand I_19189 (I328784,I329099,I328932);
nand I_19190 (I329161,I329065,I329082);
nand I_19191 (I328805,I329099,I329161);
nand I_19192 (I329192,I388077,I388080);
not I_19193 (I329209,I329192);
nor I_19194 (I328781,I329209,I328847);
nor I_19195 (I329240,I329192,I388086);
not I_19196 (I329257,I329240);
nor I_19197 (I328790,I328881,I329257);
nand I_19198 (I329288,I328983,I329257);
nand I_19199 (I328799,I328966,I329288);
nor I_19200 (I328796,I328864,I329240);
nand I_19201 (I329333,I329192,I328881);
not I_19202 (I329350,I329333);
DFFARX1 I_19203 (I329350,I2898,I328813,I328793,);
not I_19204 (I329408,I2905);
or I_19205 (I329425,I429648,I429645);
nand I_19206 (I329442,I429651,I429669);
not I_19207 (I329459,I329442);
nand I_19208 (I329476,I329459,I329425);
or I_19209 (I329493,I429660,I429654);
nor I_19210 (I329510,I329493,I429675);
nand I_19211 (I329527,I329459,I329510);
nor I_19212 (I329544,I329510,I329442);
not I_19213 (I329561,I329544);
not I_19214 (I329578,I329510);
nand I_19215 (I329397,I329476,I329578);
nor I_19216 (I329609,I429642,I429666);
nor I_19217 (I329626,I329609,I429672);
nor I_19218 (I329643,I329626,I329442);
nor I_19219 (I329660,I329578,I329626);
nor I_19220 (I329677,I429642,I429645);
nand I_19221 (I329694,I329677,I329643);
not I_19222 (I329711,I329694);
nor I_19223 (I329382,I329476,I329711);
nand I_19224 (I329379,I329694,I329527);
nand I_19225 (I329756,I329660,I329677);
nand I_19226 (I329400,I329694,I329756);
nand I_19227 (I329787,I429648,I429657);
not I_19228 (I329804,I329787);
nor I_19229 (I329376,I329804,I329442);
nor I_19230 (I329835,I329787,I429663);
not I_19231 (I329852,I329835);
nor I_19232 (I329385,I329476,I329852);
nand I_19233 (I329883,I329578,I329852);
nand I_19234 (I329394,I329561,I329883);
nor I_19235 (I329391,I329459,I329835);
nand I_19236 (I329928,I329787,I329476);
not I_19237 (I329945,I329928);
DFFARX1 I_19238 (I329945,I2898,I329408,I329388,);
not I_19239 (I330003,I2905);
or I_19240 (I330020,I146375,I146354);
nand I_19241 (I330037,I146360,I146378);
not I_19242 (I330054,I330037);
nand I_19243 (I330071,I330054,I330020);
or I_19244 (I330088,I146354,I146369);
nor I_19245 (I330105,I330088,I146366);
nand I_19246 (I330122,I330054,I330105);
nor I_19247 (I330139,I330105,I330037);
not I_19248 (I330156,I330139);
not I_19249 (I330173,I330105);
nand I_19250 (I329992,I330071,I330173);
nor I_19251 (I330204,I146372,I146384);
nor I_19252 (I330221,I330204,I146357);
nor I_19253 (I330238,I330221,I330037);
nor I_19254 (I330255,I330173,I330221);
nor I_19255 (I330272,I146363,I146381);
nand I_19256 (I330289,I330272,I330238);
not I_19257 (I330306,I330289);
nor I_19258 (I329977,I330071,I330306);
nand I_19259 (I329974,I330289,I330122);
nand I_19260 (I330351,I330255,I330272);
nand I_19261 (I329995,I330289,I330351);
nand I_19262 (I330382,I146357,I146387);
not I_19263 (I330399,I330382);
nor I_19264 (I329971,I330399,I330037);
nor I_19265 (I330430,I330382,I146360);
not I_19266 (I330447,I330430);
nor I_19267 (I329980,I330071,I330447);
nand I_19268 (I330478,I330173,I330447);
nand I_19269 (I329989,I330156,I330478);
nor I_19270 (I329986,I330054,I330430);
nand I_19271 (I330523,I330382,I330071);
not I_19272 (I330540,I330523);
DFFARX1 I_19273 (I330540,I2898,I330003,I329983,);
not I_19274 (I330598,I2905);
or I_19275 (I330615,I87153,I87126);
nand I_19276 (I330632,I87138,I87132);
not I_19277 (I330649,I330632);
nand I_19278 (I330666,I330649,I330615);
or I_19279 (I330683,I87135,I87150);
nor I_19280 (I330700,I330683,I87129);
nand I_19281 (I330717,I330649,I330700);
nor I_19282 (I330734,I330700,I330632);
not I_19283 (I330751,I330734);
not I_19284 (I330768,I330700);
nand I_19285 (I330587,I330666,I330768);
nor I_19286 (I330799,I87147,I87129);
nor I_19287 (I330816,I330799,I87135);
nor I_19288 (I330833,I330816,I330632);
nor I_19289 (I330850,I330768,I330816);
nor I_19290 (I330867,I87126,I87144);
nand I_19291 (I330884,I330867,I330833);
not I_19292 (I330901,I330884);
nor I_19293 (I330572,I330666,I330901);
nand I_19294 (I330569,I330884,I330717);
nand I_19295 (I330946,I330850,I330867);
nand I_19296 (I330590,I330884,I330946);
nand I_19297 (I330977,I87132,I87141);
not I_19298 (I330994,I330977);
nor I_19299 (I330566,I330994,I330632);
nor I_19300 (I331025,I330977,I87138);
not I_19301 (I331042,I331025);
nor I_19302 (I330575,I330666,I331042);
nand I_19303 (I331073,I330768,I331042);
nand I_19304 (I330584,I330751,I331073);
nor I_19305 (I330581,I330649,I331025);
nand I_19306 (I331118,I330977,I330666);
not I_19307 (I331135,I331118);
DFFARX1 I_19308 (I331135,I2898,I330598,I330578,);
not I_19309 (I331193,I2905);
or I_19310 (I331210,I14644,I14650);
nand I_19311 (I331227,I14653,I14638);
not I_19312 (I331244,I331227);
nand I_19313 (I331261,I331244,I331210);
or I_19314 (I331278,I14644,I14665);
nor I_19315 (I331295,I331278,I14641);
nand I_19316 (I331312,I331244,I331295);
nor I_19317 (I331329,I331295,I331227);
not I_19318 (I331346,I331329);
not I_19319 (I331363,I331295);
nand I_19320 (I331182,I331261,I331363);
nor I_19321 (I331394,I14647,I14662);
nor I_19322 (I331411,I331394,I14638);
nor I_19323 (I331428,I331411,I331227);
nor I_19324 (I331445,I331363,I331411);
nor I_19325 (I331462,I14650,I14656);
nand I_19326 (I331479,I331462,I331428);
not I_19327 (I331496,I331479);
nor I_19328 (I331167,I331261,I331496);
nand I_19329 (I331164,I331479,I331312);
nand I_19330 (I331541,I331445,I331462);
nand I_19331 (I331185,I331479,I331541);
nand I_19332 (I331572,I14647,I14659);
not I_19333 (I331589,I331572);
nor I_19334 (I331161,I331589,I331227);
nor I_19335 (I331620,I331572,I14641);
not I_19336 (I331637,I331620);
nor I_19337 (I331170,I331261,I331637);
nand I_19338 (I331668,I331363,I331637);
nand I_19339 (I331179,I331346,I331668);
nor I_19340 (I331176,I331244,I331620);
nand I_19341 (I331713,I331572,I331261);
not I_19342 (I331730,I331713);
DFFARX1 I_19343 (I331730,I2898,I331193,I331173,);
not I_19344 (I331788,I2905);
or I_19345 (I331805,I31066,I31072);
nand I_19346 (I331822,I31075,I31060);
not I_19347 (I331839,I331822);
nand I_19348 (I331856,I331839,I331805);
or I_19349 (I331873,I31066,I31087);
nor I_19350 (I331890,I331873,I31063);
nand I_19351 (I331907,I331839,I331890);
nor I_19352 (I331924,I331890,I331822);
not I_19353 (I331941,I331924);
not I_19354 (I331958,I331890);
nand I_19355 (I331777,I331856,I331958);
nor I_19356 (I331989,I31069,I31084);
nor I_19357 (I332006,I331989,I31060);
nor I_19358 (I332023,I332006,I331822);
nor I_19359 (I332040,I331958,I332006);
nor I_19360 (I332057,I31072,I31078);
nand I_19361 (I332074,I332057,I332023);
not I_19362 (I332091,I332074);
nor I_19363 (I331762,I331856,I332091);
nand I_19364 (I331759,I332074,I331907);
nand I_19365 (I332136,I332040,I332057);
nand I_19366 (I331780,I332074,I332136);
nand I_19367 (I332167,I31069,I31081);
not I_19368 (I332184,I332167);
nor I_19369 (I331756,I332184,I331822);
nor I_19370 (I332215,I332167,I31063);
not I_19371 (I332232,I332215);
nor I_19372 (I331765,I331856,I332232);
nand I_19373 (I332263,I331958,I332232);
nand I_19374 (I331774,I331941,I332263);
nor I_19375 (I331771,I331839,I332215);
nand I_19376 (I332308,I332167,I331856);
not I_19377 (I332325,I332308);
DFFARX1 I_19378 (I332325,I2898,I331788,I331768,);
not I_19379 (I332383,I2905);
or I_19380 (I332400,I296657,I296669);
nand I_19381 (I332417,I296675,I296672);
not I_19382 (I332434,I332417);
nand I_19383 (I332451,I332434,I332400);
or I_19384 (I332468,I296666,I296651);
nor I_19385 (I332485,I332468,I296681);
nand I_19386 (I332502,I332434,I332485);
nor I_19387 (I332519,I332485,I332417);
not I_19388 (I332536,I332519);
not I_19389 (I332553,I332485);
nand I_19390 (I332372,I332451,I332553);
nor I_19391 (I332584,I296678,I296660);
nor I_19392 (I332601,I332584,I296654);
nor I_19393 (I332618,I332601,I332417);
nor I_19394 (I332635,I332553,I332601);
nor I_19395 (I332652,I296657,I296660);
nand I_19396 (I332669,I332652,I332618);
not I_19397 (I332686,I332669);
nor I_19398 (I332357,I332451,I332686);
nand I_19399 (I332354,I332669,I332502);
nand I_19400 (I332731,I332635,I332652);
nand I_19401 (I332375,I332669,I332731);
nand I_19402 (I332762,I296651,I296663);
not I_19403 (I332779,I332762);
nor I_19404 (I332351,I332779,I332417);
nor I_19405 (I332810,I332762,I296654);
not I_19406 (I332827,I332810);
nor I_19407 (I332360,I332451,I332827);
nand I_19408 (I332858,I332553,I332827);
nand I_19409 (I332369,I332536,I332858);
nor I_19410 (I332366,I332434,I332810);
nand I_19411 (I332903,I332762,I332451);
not I_19412 (I332920,I332903);
DFFARX1 I_19413 (I332920,I2898,I332383,I332363,);
not I_19414 (I332978,I2905);
or I_19415 (I332995,I230667,I230646);
nand I_19416 (I333012,I230643,I230658);
not I_19417 (I333029,I333012);
nand I_19418 (I333046,I333029,I332995);
or I_19419 (I333063,I230655,I230646);
nor I_19420 (I333080,I333063,I230652);
nand I_19421 (I333097,I333029,I333080);
nor I_19422 (I333114,I333080,I333012);
not I_19423 (I333131,I333114);
not I_19424 (I333148,I333080);
nand I_19425 (I332967,I333046,I333148);
nor I_19426 (I333179,I230649,I230649);
nor I_19427 (I333196,I333179,I230670);
nor I_19428 (I333213,I333196,I333012);
nor I_19429 (I333230,I333148,I333196);
nor I_19430 (I333247,I230640,I230661);
nand I_19431 (I333264,I333247,I333213);
not I_19432 (I333281,I333264);
nor I_19433 (I332952,I333046,I333281);
nand I_19434 (I332949,I333264,I333097);
nand I_19435 (I333326,I333230,I333247);
nand I_19436 (I332970,I333264,I333326);
nand I_19437 (I333357,I230643,I230664);
not I_19438 (I333374,I333357);
nor I_19439 (I332946,I333374,I333012);
nor I_19440 (I333405,I333357,I230640);
not I_19441 (I333422,I333405);
nor I_19442 (I332955,I333046,I333422);
nand I_19443 (I333453,I333148,I333422);
nand I_19444 (I332964,I333131,I333453);
nor I_19445 (I332961,I333029,I333405);
nand I_19446 (I333498,I333357,I333046);
not I_19447 (I333515,I333498);
DFFARX1 I_19448 (I333515,I2898,I332978,I332958,);
not I_19449 (I333573,I2905);
or I_19450 (I333590,I399284,I399281);
nand I_19451 (I333607,I399272,I399269);
not I_19452 (I333624,I333607);
nand I_19453 (I333641,I333624,I333590);
or I_19454 (I333658,I399266,I399278);
nor I_19455 (I333675,I333658,I399269);
nand I_19456 (I333692,I333624,I333675);
nor I_19457 (I333709,I333675,I333607);
not I_19458 (I333726,I333709);
not I_19459 (I333743,I333675);
nand I_19460 (I333562,I333641,I333743);
nor I_19461 (I333774,I399266,I399272);
nor I_19462 (I333791,I333774,I399278);
nor I_19463 (I333808,I333791,I333607);
nor I_19464 (I333825,I333743,I333791);
nor I_19465 (I333842,I399263,I399263);
nand I_19466 (I333859,I333842,I333808);
not I_19467 (I333876,I333859);
nor I_19468 (I333547,I333641,I333876);
nand I_19469 (I333544,I333859,I333692);
nand I_19470 (I333921,I333825,I333842);
nand I_19471 (I333565,I333859,I333921);
nand I_19472 (I333952,I399275,I399287);
not I_19473 (I333969,I333952);
nor I_19474 (I333541,I333969,I333607);
nor I_19475 (I334000,I333952,I399275);
not I_19476 (I334017,I334000);
nor I_19477 (I333550,I333641,I334017);
nand I_19478 (I334048,I333743,I334017);
nand I_19479 (I333559,I333726,I334048);
nor I_19480 (I333556,I333624,I334000);
nand I_19481 (I334093,I333952,I333641);
not I_19482 (I334110,I334093);
DFFARX1 I_19483 (I334110,I2898,I333573,I333553,);
not I_19484 (I334168,I2905);
or I_19485 (I334185,I192524,I192509);
nand I_19486 (I334202,I192518,I192524);
not I_19487 (I334219,I334202);
nand I_19488 (I334236,I334219,I334185);
or I_19489 (I334253,I192527,I192515);
nor I_19490 (I334270,I334253,I192515);
nand I_19491 (I334287,I334219,I334270);
nor I_19492 (I334304,I334270,I334202);
not I_19493 (I334321,I334304);
not I_19494 (I334338,I334270);
nand I_19495 (I334157,I334236,I334338);
nor I_19496 (I334369,I192521,I192521);
nor I_19497 (I334386,I334369,I192530);
nor I_19498 (I334403,I334386,I334202);
nor I_19499 (I334420,I334338,I334386);
nor I_19500 (I334437,I192518,I192533);
nand I_19501 (I334454,I334437,I334403);
not I_19502 (I334471,I334454);
nor I_19503 (I334142,I334236,I334471);
nand I_19504 (I334139,I334454,I334287);
nand I_19505 (I334516,I334420,I334437);
nand I_19506 (I334160,I334454,I334516);
nand I_19507 (I334547,I192512,I192512);
not I_19508 (I334564,I334547);
nor I_19509 (I334136,I334564,I334202);
nor I_19510 (I334595,I334547,I192509);
not I_19511 (I334612,I334595);
nor I_19512 (I334145,I334236,I334612);
nand I_19513 (I334643,I334338,I334612);
nand I_19514 (I334154,I334321,I334643);
nor I_19515 (I334151,I334219,I334595);
nand I_19516 (I334688,I334547,I334236);
not I_19517 (I334705,I334688);
DFFARX1 I_19518 (I334705,I2898,I334168,I334148,);
not I_19519 (I334763,I2905);
or I_19520 (I334780,I365688,I365691);
nand I_19521 (I334797,I365703,I365709);
not I_19522 (I334814,I334797);
nand I_19523 (I334831,I334814,I334780);
or I_19524 (I334848,I365688,I365694);
nor I_19525 (I334865,I334848,I365691);
nand I_19526 (I334882,I334814,I334865);
nor I_19527 (I334899,I334865,I334797);
not I_19528 (I334916,I334899);
not I_19529 (I334933,I334865);
nand I_19530 (I334752,I334831,I334933);
nor I_19531 (I334964,I365712,I365706);
nor I_19532 (I334981,I334964,I365721);
nor I_19533 (I334998,I334981,I334797);
nor I_19534 (I335015,I334933,I334981);
nor I_19535 (I335032,I365715,I365697);
nand I_19536 (I335049,I335032,I334998);
not I_19537 (I335066,I335049);
nor I_19538 (I334737,I334831,I335066);
nand I_19539 (I334734,I335049,I334882);
nand I_19540 (I335111,I335015,I335032);
nand I_19541 (I334755,I335049,I335111);
nand I_19542 (I335142,I365694,I365718);
not I_19543 (I335159,I335142);
nor I_19544 (I334731,I335159,I334797);
nor I_19545 (I335190,I335142,I365700);
not I_19546 (I335207,I335190);
nor I_19547 (I334740,I334831,I335207);
nand I_19548 (I335238,I334933,I335207);
nand I_19549 (I334749,I334916,I335238);
nor I_19550 (I334746,I334814,I335190);
nand I_19551 (I335283,I335142,I334831);
not I_19552 (I335300,I335283);
DFFARX1 I_19553 (I335300,I2898,I334763,I334743,);
not I_19554 (I335358,I2905);
or I_19555 (I335375,I81492,I81465);
nand I_19556 (I335392,I81477,I81471);
not I_19557 (I335409,I335392);
nand I_19558 (I335426,I335409,I335375);
or I_19559 (I335443,I81474,I81489);
nor I_19560 (I335460,I335443,I81468);
nand I_19561 (I335477,I335409,I335460);
nor I_19562 (I335494,I335460,I335392);
not I_19563 (I335511,I335494);
not I_19564 (I335528,I335460);
nand I_19565 (I335347,I335426,I335528);
nor I_19566 (I335559,I81486,I81468);
nor I_19567 (I335576,I335559,I81474);
nor I_19568 (I335593,I335576,I335392);
nor I_19569 (I335610,I335528,I335576);
nor I_19570 (I335627,I81465,I81483);
nand I_19571 (I335644,I335627,I335593);
not I_19572 (I335661,I335644);
nor I_19573 (I335332,I335426,I335661);
nand I_19574 (I335329,I335644,I335477);
nand I_19575 (I335706,I335610,I335627);
nand I_19576 (I335350,I335644,I335706);
nand I_19577 (I335737,I81471,I81480);
not I_19578 (I335754,I335737);
nor I_19579 (I335326,I335754,I335392);
nor I_19580 (I335785,I335737,I81477);
not I_19581 (I335802,I335785);
nor I_19582 (I335335,I335426,I335802);
nand I_19583 (I335833,I335528,I335802);
nand I_19584 (I335344,I335511,I335833);
nor I_19585 (I335341,I335409,I335785);
nand I_19586 (I335878,I335737,I335426);
not I_19587 (I335895,I335878);
DFFARX1 I_19588 (I335895,I2898,I335358,I335338,);
not I_19589 (I335953,I2905);
or I_19590 (I335970,I262797,I262776);
nand I_19591 (I335987,I262773,I262788);
not I_19592 (I336004,I335987);
nand I_19593 (I336021,I336004,I335970);
or I_19594 (I336038,I262785,I262776);
nor I_19595 (I336055,I336038,I262782);
nand I_19596 (I336072,I336004,I336055);
nor I_19597 (I336089,I336055,I335987);
not I_19598 (I336106,I336089);
not I_19599 (I336123,I336055);
nand I_19600 (I335942,I336021,I336123);
nor I_19601 (I336154,I262779,I262779);
nor I_19602 (I336171,I336154,I262800);
nor I_19603 (I336188,I336171,I335987);
nor I_19604 (I336205,I336123,I336171);
nor I_19605 (I336222,I262770,I262791);
nand I_19606 (I336239,I336222,I336188);
not I_19607 (I336256,I336239);
nor I_19608 (I335927,I336021,I336256);
nand I_19609 (I335924,I336239,I336072);
nand I_19610 (I336301,I336205,I336222);
nand I_19611 (I335945,I336239,I336301);
nand I_19612 (I336332,I262773,I262794);
not I_19613 (I336349,I336332);
nor I_19614 (I335921,I336349,I335987);
nor I_19615 (I336380,I336332,I262770);
not I_19616 (I336397,I336380);
nor I_19617 (I335930,I336021,I336397);
nand I_19618 (I336428,I336123,I336397);
nand I_19619 (I335939,I336106,I336428);
nor I_19620 (I335936,I336004,I336380);
nand I_19621 (I336473,I336332,I336021);
not I_19622 (I336490,I336473);
DFFARX1 I_19623 (I336490,I2898,I335953,I335933,);
not I_19624 (I336548,I2905);
or I_19625 (I336565,I290809,I290821);
nand I_19626 (I336582,I290827,I290824);
not I_19627 (I336599,I336582);
nand I_19628 (I336616,I336599,I336565);
or I_19629 (I336633,I290818,I290803);
nor I_19630 (I336650,I336633,I290833);
nand I_19631 (I336667,I336599,I336650);
nor I_19632 (I336684,I336650,I336582);
not I_19633 (I336701,I336684);
not I_19634 (I336718,I336650);
nand I_19635 (I336537,I336616,I336718);
nor I_19636 (I336749,I290830,I290812);
nor I_19637 (I336766,I336749,I290806);
nor I_19638 (I336783,I336766,I336582);
nor I_19639 (I336800,I336718,I336766);
nor I_19640 (I336817,I290809,I290812);
nand I_19641 (I336834,I336817,I336783);
not I_19642 (I336851,I336834);
nor I_19643 (I336522,I336616,I336851);
nand I_19644 (I336519,I336834,I336667);
nand I_19645 (I336896,I336800,I336817);
nand I_19646 (I336540,I336834,I336896);
nand I_19647 (I336927,I290803,I290815);
not I_19648 (I336944,I336927);
nor I_19649 (I336516,I336944,I336582);
nor I_19650 (I336975,I336927,I290806);
not I_19651 (I336992,I336975);
nor I_19652 (I336525,I336616,I336992);
nand I_19653 (I337023,I336718,I336992);
nand I_19654 (I336534,I336701,I337023);
nor I_19655 (I336531,I336599,I336975);
nand I_19656 (I337068,I336927,I336616);
not I_19657 (I337085,I337068);
DFFARX1 I_19658 (I337085,I2898,I336548,I336528,);
not I_19659 (I337143,I2905);
or I_19660 (I337160,I66396,I66369);
nand I_19661 (I337177,I66381,I66375);
not I_19662 (I337194,I337177);
nand I_19663 (I337211,I337194,I337160);
or I_19664 (I337228,I66378,I66393);
nor I_19665 (I337245,I337228,I66372);
nand I_19666 (I337262,I337194,I337245);
nor I_19667 (I337279,I337245,I337177);
not I_19668 (I337296,I337279);
not I_19669 (I337313,I337245);
nand I_19670 (I337132,I337211,I337313);
nor I_19671 (I337344,I66390,I66372);
nor I_19672 (I337361,I337344,I66378);
nor I_19673 (I337378,I337361,I337177);
nor I_19674 (I337395,I337313,I337361);
nor I_19675 (I337412,I66369,I66387);
nand I_19676 (I337429,I337412,I337378);
not I_19677 (I337446,I337429);
nor I_19678 (I337117,I337211,I337446);
nand I_19679 (I337114,I337429,I337262);
nand I_19680 (I337491,I337395,I337412);
nand I_19681 (I337135,I337429,I337491);
nand I_19682 (I337522,I66375,I66384);
not I_19683 (I337539,I337522);
nor I_19684 (I337111,I337539,I337177);
nor I_19685 (I337570,I337522,I66381);
not I_19686 (I337587,I337570);
nor I_19687 (I337120,I337211,I337587);
nand I_19688 (I337618,I337313,I337587);
nand I_19689 (I337129,I337296,I337618);
nor I_19690 (I337126,I337194,I337570);
nand I_19691 (I337663,I337522,I337211);
not I_19692 (I337680,I337663);
DFFARX1 I_19693 (I337680,I2898,I337143,I337123,);
not I_19694 (I337738,I2905);
or I_19695 (I337755,I426163,I426160);
nand I_19696 (I337772,I426166,I426184);
not I_19697 (I337789,I337772);
nand I_19698 (I337806,I337789,I337755);
or I_19699 (I337823,I426175,I426169);
nor I_19700 (I337840,I337823,I426190);
nand I_19701 (I337857,I337789,I337840);
nor I_19702 (I337874,I337840,I337772);
not I_19703 (I337891,I337874);
not I_19704 (I337908,I337840);
nand I_19705 (I337727,I337806,I337908);
nor I_19706 (I337939,I426157,I426181);
nor I_19707 (I337956,I337939,I426187);
nor I_19708 (I337973,I337956,I337772);
nor I_19709 (I337990,I337908,I337956);
nor I_19710 (I338007,I426157,I426160);
nand I_19711 (I338024,I338007,I337973);
not I_19712 (I338041,I338024);
nor I_19713 (I337712,I337806,I338041);
nand I_19714 (I337709,I338024,I337857);
nand I_19715 (I338086,I337990,I338007);
nand I_19716 (I337730,I338024,I338086);
nand I_19717 (I338117,I426163,I426172);
not I_19718 (I338134,I338117);
nor I_19719 (I337706,I338134,I337772);
nor I_19720 (I338165,I338117,I426178);
not I_19721 (I338182,I338165);
nor I_19722 (I337715,I337806,I338182);
nand I_19723 (I338213,I337908,I338182);
nand I_19724 (I337724,I337891,I338213);
nor I_19725 (I337721,I337789,I338165);
nand I_19726 (I338258,I338117,I337806);
not I_19727 (I338275,I338258);
DFFARX1 I_19728 (I338275,I2898,I337738,I337718,);
not I_19729 (I338333,I2905);
or I_19730 (I338350,I439406,I439403);
nand I_19731 (I338367,I439409,I439427);
not I_19732 (I338384,I338367);
nand I_19733 (I338401,I338384,I338350);
or I_19734 (I338418,I439418,I439412);
nor I_19735 (I338435,I338418,I439433);
nand I_19736 (I338452,I338384,I338435);
nor I_19737 (I338469,I338435,I338367);
not I_19738 (I338486,I338469);
not I_19739 (I338503,I338435);
nand I_19740 (I338322,I338401,I338503);
nor I_19741 (I338534,I439400,I439424);
nor I_19742 (I338551,I338534,I439430);
nor I_19743 (I338568,I338551,I338367);
nor I_19744 (I338585,I338503,I338551);
nor I_19745 (I338602,I439400,I439403);
nand I_19746 (I338619,I338602,I338568);
not I_19747 (I338636,I338619);
nor I_19748 (I338307,I338401,I338636);
nand I_19749 (I338304,I338619,I338452);
nand I_19750 (I338681,I338585,I338602);
nand I_19751 (I338325,I338619,I338681);
nand I_19752 (I338712,I439406,I439415);
not I_19753 (I338729,I338712);
nor I_19754 (I338301,I338729,I338367);
nor I_19755 (I338760,I338712,I439421);
not I_19756 (I338777,I338760);
nor I_19757 (I338310,I338401,I338777);
nand I_19758 (I338808,I338503,I338777);
nand I_19759 (I338319,I338486,I338808);
nor I_19760 (I338316,I338384,I338760);
nand I_19761 (I338853,I338712,I338401);
not I_19762 (I338870,I338853);
DFFARX1 I_19763 (I338870,I2898,I338333,I338313,);
not I_19764 (I338928,I2905);
or I_19765 (I338945,I183463,I183448);
nand I_19766 (I338962,I183457,I183463);
not I_19767 (I338979,I338962);
nand I_19768 (I338996,I338979,I338945);
or I_19769 (I339013,I183466,I183454);
nor I_19770 (I339030,I339013,I183454);
nand I_19771 (I339047,I338979,I339030);
nor I_19772 (I339064,I339030,I338962);
not I_19773 (I339081,I339064);
not I_19774 (I339098,I339030);
nand I_19775 (I338917,I338996,I339098);
nor I_19776 (I339129,I183460,I183460);
nor I_19777 (I339146,I339129,I183469);
nor I_19778 (I339163,I339146,I338962);
nor I_19779 (I339180,I339098,I339146);
nor I_19780 (I339197,I183457,I183472);
nand I_19781 (I339214,I339197,I339163);
not I_19782 (I339231,I339214);
nor I_19783 (I338902,I338996,I339231);
nand I_19784 (I338899,I339214,I339047);
nand I_19785 (I339276,I339180,I339197);
nand I_19786 (I338920,I339214,I339276);
nand I_19787 (I339307,I183451,I183451);
not I_19788 (I339324,I339307);
nor I_19789 (I338896,I339324,I338962);
nor I_19790 (I339355,I339307,I183448);
not I_19791 (I339372,I339355);
nor I_19792 (I338905,I338996,I339372);
nand I_19793 (I339403,I339098,I339372);
nand I_19794 (I338914,I339081,I339403);
nor I_19795 (I338911,I338979,I339355);
nand I_19796 (I339448,I339307,I338996);
not I_19797 (I339465,I339448);
DFFARX1 I_19798 (I339465,I2898,I338928,I338908,);
not I_19799 (I339523,I2905);
or I_19800 (I339540,I187645,I187630);
nand I_19801 (I339557,I187639,I187645);
not I_19802 (I339574,I339557);
nand I_19803 (I339591,I339574,I339540);
or I_19804 (I339608,I187648,I187636);
nor I_19805 (I339625,I339608,I187636);
nand I_19806 (I339642,I339574,I339625);
nor I_19807 (I339659,I339625,I339557);
not I_19808 (I339676,I339659);
not I_19809 (I339693,I339625);
nand I_19810 (I339512,I339591,I339693);
nor I_19811 (I339724,I187642,I187642);
nor I_19812 (I339741,I339724,I187651);
nor I_19813 (I339758,I339741,I339557);
nor I_19814 (I339775,I339693,I339741);
nor I_19815 (I339792,I187639,I187654);
nand I_19816 (I339809,I339792,I339758);
not I_19817 (I339826,I339809);
nor I_19818 (I339497,I339591,I339826);
nand I_19819 (I339494,I339809,I339642);
nand I_19820 (I339871,I339775,I339792);
nand I_19821 (I339515,I339809,I339871);
nand I_19822 (I339902,I187633,I187633);
not I_19823 (I339919,I339902);
nor I_19824 (I339491,I339919,I339557);
nor I_19825 (I339950,I339902,I187630);
not I_19826 (I339967,I339950);
nor I_19827 (I339500,I339591,I339967);
nand I_19828 (I339998,I339693,I339967);
nand I_19829 (I339509,I339676,I339998);
nor I_19830 (I339506,I339574,I339950);
nand I_19831 (I340043,I339902,I339591);
not I_19832 (I340060,I340043);
DFFARX1 I_19833 (I340060,I2898,I339523,I339503,);
not I_19834 (I340118,I2905);
or I_19835 (I340135,I440800,I440797);
nand I_19836 (I340152,I440803,I440821);
not I_19837 (I340169,I340152);
nand I_19838 (I340186,I340169,I340135);
or I_19839 (I340203,I440812,I440806);
nor I_19840 (I340220,I340203,I440827);
nand I_19841 (I340237,I340169,I340220);
nor I_19842 (I340254,I340220,I340152);
not I_19843 (I340271,I340254);
not I_19844 (I340288,I340220);
nand I_19845 (I340107,I340186,I340288);
nor I_19846 (I340319,I440794,I440818);
nor I_19847 (I340336,I340319,I440824);
nor I_19848 (I340353,I340336,I340152);
nor I_19849 (I340370,I340288,I340336);
nor I_19850 (I340387,I440794,I440797);
nand I_19851 (I340404,I340387,I340353);
not I_19852 (I340421,I340404);
nor I_19853 (I340092,I340186,I340421);
nand I_19854 (I340089,I340404,I340237);
nand I_19855 (I340466,I340370,I340387);
nand I_19856 (I340110,I340404,I340466);
nand I_19857 (I340497,I440800,I440809);
not I_19858 (I340514,I340497);
nor I_19859 (I340086,I340514,I340152);
nor I_19860 (I340545,I340497,I440815);
not I_19861 (I340562,I340545);
nor I_19862 (I340095,I340186,I340562);
nand I_19863 (I340593,I340288,I340562);
nand I_19864 (I340104,I340271,I340593);
nor I_19865 (I340101,I340169,I340545);
nand I_19866 (I340638,I340497,I340186);
not I_19867 (I340655,I340638);
DFFARX1 I_19868 (I340655,I2898,I340118,I340098,);
not I_19869 (I340713,I2905);
or I_19870 (I340730,I174255,I174234);
nand I_19871 (I340747,I174240,I174258);
not I_19872 (I340764,I340747);
nand I_19873 (I340781,I340764,I340730);
or I_19874 (I340798,I174234,I174249);
nor I_19875 (I340815,I340798,I174246);
nand I_19876 (I340832,I340764,I340815);
nor I_19877 (I340849,I340815,I340747);
not I_19878 (I340866,I340849);
not I_19879 (I340883,I340815);
nand I_19880 (I340702,I340781,I340883);
nor I_19881 (I340914,I174252,I174264);
nor I_19882 (I340931,I340914,I174237);
nor I_19883 (I340948,I340931,I340747);
nor I_19884 (I340965,I340883,I340931);
nor I_19885 (I340982,I174243,I174261);
nand I_19886 (I340999,I340982,I340948);
not I_19887 (I341016,I340999);
nor I_19888 (I340687,I340781,I341016);
nand I_19889 (I340684,I340999,I340832);
nand I_19890 (I341061,I340965,I340982);
nand I_19891 (I340705,I340999,I341061);
nand I_19892 (I341092,I174237,I174267);
not I_19893 (I341109,I341092);
nor I_19894 (I340681,I341109,I340747);
nor I_19895 (I341140,I341092,I174240);
not I_19896 (I341157,I341140);
nor I_19897 (I340690,I340781,I341157);
nand I_19898 (I341188,I340883,I341157);
nand I_19899 (I340699,I340866,I341188);
nor I_19900 (I340696,I340764,I341140);
nand I_19901 (I341233,I341092,I340781);
not I_19902 (I341250,I341233);
DFFARX1 I_19903 (I341250,I2898,I340713,I340693,);
not I_19904 (I341308,I2905);
or I_19905 (I341325,I303236,I303248);
nand I_19906 (I341342,I303254,I303251);
not I_19907 (I341359,I341342);
nand I_19908 (I341376,I341359,I341325);
or I_19909 (I341393,I303245,I303230);
nor I_19910 (I341410,I341393,I303260);
nand I_19911 (I341427,I341359,I341410);
nor I_19912 (I341444,I341410,I341342);
not I_19913 (I341461,I341444);
not I_19914 (I341478,I341410);
nand I_19915 (I341297,I341376,I341478);
nor I_19916 (I341509,I303257,I303239);
nor I_19917 (I341526,I341509,I303233);
nor I_19918 (I341543,I341526,I341342);
nor I_19919 (I341560,I341478,I341526);
nor I_19920 (I341577,I303236,I303239);
nand I_19921 (I341594,I341577,I341543);
not I_19922 (I341611,I341594);
nor I_19923 (I341282,I341376,I341611);
nand I_19924 (I341279,I341594,I341427);
nand I_19925 (I341656,I341560,I341577);
nand I_19926 (I341300,I341594,I341656);
nand I_19927 (I341687,I303230,I303242);
not I_19928 (I341704,I341687);
nor I_19929 (I341276,I341704,I341342);
nor I_19930 (I341735,I341687,I303233);
not I_19931 (I341752,I341735);
nor I_19932 (I341285,I341376,I341752);
nand I_19933 (I341783,I341478,I341752);
nand I_19934 (I341294,I341461,I341783);
nor I_19935 (I341291,I341359,I341735);
nand I_19936 (I341828,I341687,I341376);
not I_19937 (I341845,I341828);
DFFARX1 I_19938 (I341845,I2898,I341308,I341288,);
not I_19939 (I341903,I2905);
or I_19940 (I341920,I106577,I106583);
nand I_19941 (I341937,I106595,I106586);
not I_19942 (I341954,I341937);
nand I_19943 (I341971,I341954,I341920);
or I_19944 (I341988,I106592,I106574);
nor I_19945 (I342005,I341988,I106607);
nand I_19946 (I342022,I341954,I342005);
nor I_19947 (I342039,I342005,I341937);
not I_19948 (I342056,I342039);
not I_19949 (I342073,I342005);
nand I_19950 (I341892,I341971,I342073);
nor I_19951 (I342104,I106577,I106580);
nor I_19952 (I342121,I342104,I106589);
nor I_19953 (I342138,I342121,I341937);
nor I_19954 (I342155,I342073,I342121);
nor I_19955 (I342172,I106598,I106580);
nand I_19956 (I342189,I342172,I342138);
not I_19957 (I342206,I342189);
nor I_19958 (I341877,I341971,I342206);
nand I_19959 (I341874,I342189,I342022);
nand I_19960 (I342251,I342155,I342172);
nand I_19961 (I341895,I342189,I342251);
nand I_19962 (I342282,I106604,I106601);
not I_19963 (I342299,I342282);
nor I_19964 (I341871,I342299,I341937);
nor I_19965 (I342330,I342282,I106574);
not I_19966 (I342347,I342330);
nor I_19967 (I341880,I341971,I342347);
nand I_19968 (I342378,I342073,I342347);
nand I_19969 (I341889,I342056,I342378);
nor I_19970 (I341886,I341954,I342330);
nand I_19971 (I342423,I342282,I341971);
not I_19972 (I342440,I342423);
DFFARX1 I_19973 (I342440,I2898,I341903,I341883,);
not I_19974 (I342498,I2905);
or I_19975 (I342515,I169495,I169474);
nand I_19976 (I342532,I169480,I169498);
not I_19977 (I342549,I342532);
nand I_19978 (I342566,I342549,I342515);
or I_19979 (I342583,I169474,I169489);
nor I_19980 (I342600,I342583,I169486);
nand I_19981 (I342617,I342549,I342600);
nor I_19982 (I342634,I342600,I342532);
not I_19983 (I342651,I342634);
not I_19984 (I342668,I342600);
nand I_19985 (I342487,I342566,I342668);
nor I_19986 (I342699,I169492,I169504);
nor I_19987 (I342716,I342699,I169477);
nor I_19988 (I342733,I342716,I342532);
nor I_19989 (I342750,I342668,I342716);
nor I_19990 (I342767,I169483,I169501);
nand I_19991 (I342784,I342767,I342733);
not I_19992 (I342801,I342784);
nor I_19993 (I342472,I342566,I342801);
nand I_19994 (I342469,I342784,I342617);
nand I_19995 (I342846,I342750,I342767);
nand I_19996 (I342490,I342784,I342846);
nand I_19997 (I342877,I169477,I169507);
not I_19998 (I342894,I342877);
nor I_19999 (I342466,I342894,I342532);
nor I_20000 (I342925,I342877,I169480);
not I_20001 (I342942,I342925);
nor I_20002 (I342475,I342566,I342942);
nand I_20003 (I342973,I342668,I342942);
nand I_20004 (I342484,I342651,I342973);
nor I_20005 (I342481,I342549,I342925);
nand I_20006 (I343018,I342877,I342566);
not I_20007 (I343035,I343018);
DFFARX1 I_20008 (I343035,I2898,I342498,I342478,);
not I_20009 (I343093,I2905);
or I_20010 (I343110,I273507,I273486);
nand I_20011 (I343127,I273483,I273498);
not I_20012 (I343144,I343127);
nand I_20013 (I343161,I343144,I343110);
or I_20014 (I343178,I273495,I273486);
nor I_20015 (I343195,I343178,I273492);
nand I_20016 (I343212,I343144,I343195);
nor I_20017 (I343229,I343195,I343127);
not I_20018 (I343246,I343229);
not I_20019 (I343263,I343195);
nand I_20020 (I343082,I343161,I343263);
nor I_20021 (I343294,I273489,I273489);
nor I_20022 (I343311,I343294,I273510);
nor I_20023 (I343328,I343311,I343127);
nor I_20024 (I343345,I343263,I343311);
nor I_20025 (I343362,I273480,I273501);
nand I_20026 (I343379,I343362,I343328);
not I_20027 (I343396,I343379);
nor I_20028 (I343067,I343161,I343396);
nand I_20029 (I343064,I343379,I343212);
nand I_20030 (I343441,I343345,I343362);
nand I_20031 (I343085,I343379,I343441);
nand I_20032 (I343472,I273483,I273504);
not I_20033 (I343489,I343472);
nor I_20034 (I343061,I343489,I343127);
nor I_20035 (I343520,I343472,I273480);
not I_20036 (I343537,I343520);
nor I_20037 (I343070,I343161,I343537);
nand I_20038 (I343568,I343263,I343537);
nand I_20039 (I343079,I343246,I343568);
nor I_20040 (I343076,I343144,I343520);
nand I_20041 (I343613,I343472,I343161);
not I_20042 (I343630,I343613);
DFFARX1 I_20043 (I343630,I2898,I343093,I343073,);
not I_20044 (I343688,I2905);
or I_20045 (I343705,I122302,I122308);
nand I_20046 (I343722,I122320,I122311);
not I_20047 (I343739,I343722);
nand I_20048 (I343756,I343739,I343705);
or I_20049 (I343773,I122317,I122299);
nor I_20050 (I343790,I343773,I122332);
nand I_20051 (I343807,I343739,I343790);
nor I_20052 (I343824,I343790,I343722);
not I_20053 (I343841,I343824);
not I_20054 (I343858,I343790);
nand I_20055 (I343677,I343756,I343858);
nor I_20056 (I343889,I122302,I122305);
nor I_20057 (I343906,I343889,I122314);
nor I_20058 (I343923,I343906,I343722);
nor I_20059 (I343940,I343858,I343906);
nor I_20060 (I343957,I122323,I122305);
nand I_20061 (I343974,I343957,I343923);
not I_20062 (I343991,I343974);
nor I_20063 (I343662,I343756,I343991);
nand I_20064 (I343659,I343974,I343807);
nand I_20065 (I344036,I343940,I343957);
nand I_20066 (I343680,I343974,I344036);
nand I_20067 (I344067,I122329,I122326);
not I_20068 (I344084,I344067);
nor I_20069 (I343656,I344084,I343722);
nor I_20070 (I344115,I344067,I122299);
not I_20071 (I344132,I344115);
nor I_20072 (I343665,I343756,I344132);
nand I_20073 (I344163,I343858,I344132);
nand I_20074 (I343674,I343841,I344163);
nor I_20075 (I343671,I343739,I344115);
nand I_20076 (I344208,I344067,I343756);
not I_20077 (I344225,I344208);
DFFARX1 I_20078 (I344225,I2898,I343688,I343668,);
not I_20079 (I344283,I2905);
or I_20080 (I344300,I287885,I287897);
nand I_20081 (I344317,I287903,I287900);
not I_20082 (I344334,I344317);
nand I_20083 (I344351,I344334,I344300);
or I_20084 (I344368,I287894,I287879);
nor I_20085 (I344385,I344368,I287909);
nand I_20086 (I344402,I344334,I344385);
nor I_20087 (I344419,I344385,I344317);
not I_20088 (I344436,I344419);
not I_20089 (I344453,I344385);
nand I_20090 (I344272,I344351,I344453);
nor I_20091 (I344484,I287906,I287888);
nor I_20092 (I344501,I344484,I287882);
nor I_20093 (I344518,I344501,I344317);
nor I_20094 (I344535,I344453,I344501);
nor I_20095 (I344552,I287885,I287888);
nand I_20096 (I344569,I344552,I344518);
not I_20097 (I344586,I344569);
nor I_20098 (I344257,I344351,I344586);
nand I_20099 (I344254,I344569,I344402);
nand I_20100 (I344631,I344535,I344552);
nand I_20101 (I344275,I344569,I344631);
nand I_20102 (I344662,I287879,I287891);
not I_20103 (I344679,I344662);
nor I_20104 (I344251,I344679,I344317);
nor I_20105 (I344710,I344662,I287882);
not I_20106 (I344727,I344710);
nor I_20107 (I344260,I344351,I344727);
nand I_20108 (I344758,I344453,I344727);
nand I_20109 (I344269,I344436,I344758);
nor I_20110 (I344266,I344334,I344710);
nand I_20111 (I344803,I344662,I344351);
not I_20112 (I344820,I344803);
DFFARX1 I_20113 (I344820,I2898,I344283,I344263,);
not I_20114 (I344878,I2905);
or I_20115 (I344895,I113496,I113502);
nand I_20116 (I344912,I113514,I113505);
not I_20117 (I344929,I344912);
nand I_20118 (I344946,I344929,I344895);
or I_20119 (I344963,I113511,I113493);
nor I_20120 (I344980,I344963,I113526);
nand I_20121 (I344997,I344929,I344980);
nor I_20122 (I345014,I344980,I344912);
not I_20123 (I345031,I345014);
not I_20124 (I345048,I344980);
nand I_20125 (I344867,I344946,I345048);
nor I_20126 (I345079,I113496,I113499);
nor I_20127 (I345096,I345079,I113508);
nor I_20128 (I345113,I345096,I344912);
nor I_20129 (I345130,I345048,I345096);
nor I_20130 (I345147,I113517,I113499);
nand I_20131 (I345164,I345147,I345113);
not I_20132 (I345181,I345164);
nor I_20133 (I344852,I344946,I345181);
nand I_20134 (I344849,I345164,I344997);
nand I_20135 (I345226,I345130,I345147);
nand I_20136 (I344870,I345164,I345226);
nand I_20137 (I345257,I113523,I113520);
not I_20138 (I345274,I345257);
nor I_20139 (I344846,I345274,I344912);
nor I_20140 (I345305,I345257,I113493);
not I_20141 (I345322,I345305);
nor I_20142 (I344855,I344946,I345322);
nand I_20143 (I345353,I345048,I345322);
nand I_20144 (I344864,I345031,I345353);
nor I_20145 (I344861,I344929,I345305);
nand I_20146 (I345398,I345257,I344946);
not I_20147 (I345415,I345398);
DFFARX1 I_20148 (I345415,I2898,I344878,I344858,);
not I_20149 (I345473,I2905);
or I_20150 (I345490,I124189,I124195);
nand I_20151 (I345507,I124207,I124198);
not I_20152 (I345524,I345507);
nand I_20153 (I345541,I345524,I345490);
or I_20154 (I345558,I124204,I124186);
nor I_20155 (I345575,I345558,I124219);
nand I_20156 (I345592,I345524,I345575);
nor I_20157 (I345609,I345575,I345507);
not I_20158 (I345626,I345609);
not I_20159 (I345643,I345575);
nand I_20160 (I345462,I345541,I345643);
nor I_20161 (I345674,I124189,I124192);
nor I_20162 (I345691,I345674,I124201);
nor I_20163 (I345708,I345691,I345507);
nor I_20164 (I345725,I345643,I345691);
nor I_20165 (I345742,I124210,I124192);
nand I_20166 (I345759,I345742,I345708);
not I_20167 (I345776,I345759);
nor I_20168 (I345447,I345541,I345776);
nand I_20169 (I345444,I345759,I345592);
nand I_20170 (I345821,I345725,I345742);
nand I_20171 (I345465,I345759,I345821);
nand I_20172 (I345852,I124216,I124213);
not I_20173 (I345869,I345852);
nor I_20174 (I345441,I345869,I345507);
nor I_20175 (I345900,I345852,I124186);
not I_20176 (I345917,I345900);
nor I_20177 (I345450,I345541,I345917);
nand I_20178 (I345948,I345643,I345917);
nand I_20179 (I345459,I345626,I345948);
nor I_20180 (I345456,I345524,I345900);
nand I_20181 (I345993,I345852,I345541);
not I_20182 (I346010,I345993);
DFFARX1 I_20183 (I346010,I2898,I345473,I345453,);
not I_20184 (I346068,I2905);
or I_20185 (I346085,I27496,I27502);
nand I_20186 (I346102,I27505,I27490);
not I_20187 (I346119,I346102);
nand I_20188 (I346136,I346119,I346085);
or I_20189 (I346153,I27496,I27517);
nor I_20190 (I346170,I346153,I27493);
nand I_20191 (I346187,I346119,I346170);
nor I_20192 (I346204,I346170,I346102);
not I_20193 (I346221,I346204);
not I_20194 (I346238,I346170);
nand I_20195 (I346057,I346136,I346238);
nor I_20196 (I346269,I27499,I27514);
nor I_20197 (I346286,I346269,I27490);
nor I_20198 (I346303,I346286,I346102);
nor I_20199 (I346320,I346238,I346286);
nor I_20200 (I346337,I27502,I27508);
nand I_20201 (I346354,I346337,I346303);
not I_20202 (I346371,I346354);
nor I_20203 (I346042,I346136,I346371);
nand I_20204 (I346039,I346354,I346187);
nand I_20205 (I346416,I346320,I346337);
nand I_20206 (I346060,I346354,I346416);
nand I_20207 (I346447,I27499,I27511);
not I_20208 (I346464,I346447);
nor I_20209 (I346036,I346464,I346102);
nor I_20210 (I346495,I346447,I27493);
not I_20211 (I346512,I346495);
nor I_20212 (I346045,I346136,I346512);
nand I_20213 (I346543,I346238,I346512);
nand I_20214 (I346054,I346221,I346543);
nor I_20215 (I346051,I346119,I346495);
nand I_20216 (I346588,I346447,I346136);
not I_20217 (I346605,I346588);
DFFARX1 I_20218 (I346605,I2898,I346068,I346048,);
not I_20219 (I346663,I2905);
or I_20220 (I346680,I238317,I238296);
nand I_20221 (I346697,I238293,I238308);
not I_20222 (I346714,I346697);
nand I_20223 (I346731,I346714,I346680);
or I_20224 (I346748,I238305,I238296);
nor I_20225 (I346765,I346748,I238302);
nand I_20226 (I346782,I346714,I346765);
nor I_20227 (I346799,I346765,I346697);
not I_20228 (I346816,I346799);
not I_20229 (I346833,I346765);
nand I_20230 (I346652,I346731,I346833);
nor I_20231 (I346864,I238299,I238299);
nor I_20232 (I346881,I346864,I238320);
nor I_20233 (I346898,I346881,I346697);
nor I_20234 (I346915,I346833,I346881);
nor I_20235 (I346932,I238290,I238311);
nand I_20236 (I346949,I346932,I346898);
not I_20237 (I346966,I346949);
nor I_20238 (I346637,I346731,I346966);
nand I_20239 (I346634,I346949,I346782);
nand I_20240 (I347011,I346915,I346932);
nand I_20241 (I346655,I346949,I347011);
nand I_20242 (I347042,I238293,I238314);
not I_20243 (I347059,I347042);
nor I_20244 (I346631,I347059,I346697);
nor I_20245 (I347090,I347042,I238290);
not I_20246 (I347107,I347090);
nor I_20247 (I346640,I346731,I347107);
nand I_20248 (I347138,I346833,I347107);
nand I_20249 (I346649,I346816,I347138);
nor I_20250 (I346646,I346714,I347090);
nand I_20251 (I347183,I347042,I346731);
not I_20252 (I347200,I347183);
DFFARX1 I_20253 (I347200,I2898,I346663,I346643,);
not I_20254 (I347258,I2905);
or I_20255 (I347275,I265092,I265071);
nand I_20256 (I347292,I265068,I265083);
not I_20257 (I347309,I347292);
nand I_20258 (I347326,I347309,I347275);
or I_20259 (I347343,I265080,I265071);
nor I_20260 (I347360,I347343,I265077);
nand I_20261 (I347377,I347309,I347360);
nor I_20262 (I347394,I347360,I347292);
not I_20263 (I347411,I347394);
not I_20264 (I347428,I347360);
nand I_20265 (I347247,I347326,I347428);
nor I_20266 (I347459,I265074,I265074);
nor I_20267 (I347476,I347459,I265095);
nor I_20268 (I347493,I347476,I347292);
nor I_20269 (I347510,I347428,I347476);
nor I_20270 (I347527,I265065,I265086);
nand I_20271 (I347544,I347527,I347493);
not I_20272 (I347561,I347544);
nor I_20273 (I347232,I347326,I347561);
nand I_20274 (I347229,I347544,I347377);
nand I_20275 (I347606,I347510,I347527);
nand I_20276 (I347250,I347544,I347606);
nand I_20277 (I347637,I265068,I265089);
not I_20278 (I347654,I347637);
nor I_20279 (I347226,I347654,I347292);
nor I_20280 (I347685,I347637,I265065);
not I_20281 (I347702,I347685);
nor I_20282 (I347235,I347326,I347702);
nand I_20283 (I347733,I347428,I347702);
nand I_20284 (I347244,I347411,I347733);
nor I_20285 (I347241,I347309,I347685);
nand I_20286 (I347778,I347637,I347326);
not I_20287 (I347795,I347778);
DFFARX1 I_20288 (I347795,I2898,I347258,I347238,);
not I_20289 (I347853,I2905);
or I_20290 (I347870,I209708,I209711);
nand I_20291 (I347887,I209717,I209708);
not I_20292 (I347904,I347887);
nand I_20293 (I347921,I347904,I347870);
or I_20294 (I347938,I209699,I209699);
nor I_20295 (I347955,I347938,I209696);
nand I_20296 (I347972,I347904,I347955);
nor I_20297 (I347989,I347955,I347887);
not I_20298 (I348006,I347989);
not I_20299 (I348023,I347955);
nand I_20300 (I347842,I347921,I348023);
nor I_20301 (I348054,I209705,I209702);
nor I_20302 (I348071,I348054,I209714);
nor I_20303 (I348088,I348071,I347887);
nor I_20304 (I348105,I348023,I348071);
nor I_20305 (I348122,I209723,I209696);
nand I_20306 (I348139,I348122,I348088);
not I_20307 (I348156,I348139);
nor I_20308 (I347827,I347921,I348156);
nand I_20309 (I347824,I348139,I347972);
nand I_20310 (I348201,I348105,I348122);
nand I_20311 (I347845,I348139,I348201);
nand I_20312 (I348232,I209702,I209705);
not I_20313 (I348249,I348232);
nor I_20314 (I347821,I348249,I347887);
nor I_20315 (I348280,I348232,I209720);
not I_20316 (I348297,I348280);
nor I_20317 (I347830,I347921,I348297);
nand I_20318 (I348328,I348023,I348297);
nand I_20319 (I347839,I348006,I348328);
nor I_20320 (I347836,I347904,I348280);
nand I_20321 (I348373,I348232,I347921);
not I_20322 (I348390,I348373);
DFFARX1 I_20323 (I348390,I2898,I347853,I347833,);
not I_20324 (I348448,I2905);
or I_20325 (I348465,I290078,I290090);
nand I_20326 (I348482,I290096,I290093);
not I_20327 (I348499,I348482);
nand I_20328 (I348516,I348499,I348465);
or I_20329 (I348533,I290087,I290072);
nor I_20330 (I348550,I348533,I290102);
nand I_20331 (I348567,I348499,I348550);
nor I_20332 (I348584,I348550,I348482);
not I_20333 (I348601,I348584);
not I_20334 (I348618,I348550);
nand I_20335 (I348437,I348516,I348618);
nor I_20336 (I348649,I290099,I290081);
nor I_20337 (I348666,I348649,I290075);
nor I_20338 (I348683,I348666,I348482);
nor I_20339 (I348700,I348618,I348666);
nor I_20340 (I348717,I290078,I290081);
nand I_20341 (I348734,I348717,I348683);
not I_20342 (I348751,I348734);
nor I_20343 (I348422,I348516,I348751);
nand I_20344 (I348419,I348734,I348567);
nand I_20345 (I348796,I348700,I348717);
nand I_20346 (I348440,I348734,I348796);
nand I_20347 (I348827,I290072,I290084);
not I_20348 (I348844,I348827);
nor I_20349 (I348416,I348844,I348482);
nor I_20350 (I348875,I348827,I290075);
not I_20351 (I348892,I348875);
nor I_20352 (I348425,I348516,I348892);
nand I_20353 (I348923,I348618,I348892);
nand I_20354 (I348434,I348601,I348923);
nor I_20355 (I348431,I348499,I348875);
nand I_20356 (I348968,I348827,I348516);
not I_20357 (I348985,I348968);
DFFARX1 I_20358 (I348985,I2898,I348448,I348428,);
not I_20359 (I349043,I2905);
or I_20360 (I349060,I198100,I198085);
nand I_20361 (I349077,I198094,I198100);
not I_20362 (I349094,I349077);
nand I_20363 (I349111,I349094,I349060);
or I_20364 (I349128,I198103,I198091);
nor I_20365 (I349145,I349128,I198091);
nand I_20366 (I349162,I349094,I349145);
nor I_20367 (I349179,I349145,I349077);
not I_20368 (I349196,I349179);
not I_20369 (I349213,I349145);
nand I_20370 (I349032,I349111,I349213);
nor I_20371 (I349244,I198097,I198097);
nor I_20372 (I349261,I349244,I198106);
nor I_20373 (I349278,I349261,I349077);
nor I_20374 (I349295,I349213,I349261);
nor I_20375 (I349312,I198094,I198109);
nand I_20376 (I349329,I349312,I349278);
not I_20377 (I349346,I349329);
nor I_20378 (I349017,I349111,I349346);
nand I_20379 (I349014,I349329,I349162);
nand I_20380 (I349391,I349295,I349312);
nand I_20381 (I349035,I349329,I349391);
nand I_20382 (I349422,I198088,I198088);
not I_20383 (I349439,I349422);
nor I_20384 (I349011,I349439,I349077);
nor I_20385 (I349470,I349422,I198085);
not I_20386 (I349487,I349470);
nor I_20387 (I349020,I349111,I349487);
nand I_20388 (I349518,I349213,I349487);
nand I_20389 (I349029,I349196,I349518);
nor I_20390 (I349026,I349094,I349470);
nand I_20391 (I349563,I349422,I349111);
not I_20392 (I349580,I349563);
DFFARX1 I_20393 (I349580,I2898,I349043,I349023,);
not I_20394 (I349638,I2905);
or I_20395 (I349655,I426860,I426857);
nand I_20396 (I349672,I426863,I426881);
not I_20397 (I349689,I349672);
nand I_20398 (I349706,I349689,I349655);
or I_20399 (I349723,I426872,I426866);
nor I_20400 (I349740,I349723,I426887);
nand I_20401 (I349757,I349689,I349740);
nor I_20402 (I349774,I349740,I349672);
not I_20403 (I349791,I349774);
not I_20404 (I349808,I349740);
nand I_20405 (I349627,I349706,I349808);
nor I_20406 (I349839,I426854,I426878);
nor I_20407 (I349856,I349839,I426884);
nor I_20408 (I349873,I349856,I349672);
nor I_20409 (I349890,I349808,I349856);
nor I_20410 (I349907,I426854,I426857);
nand I_20411 (I349924,I349907,I349873);
not I_20412 (I349941,I349924);
nor I_20413 (I349612,I349706,I349941);
nand I_20414 (I349609,I349924,I349757);
nand I_20415 (I349986,I349890,I349907);
nand I_20416 (I349630,I349924,I349986);
nand I_20417 (I350017,I426860,I426869);
not I_20418 (I350034,I350017);
nor I_20419 (I349606,I350034,I349672);
nor I_20420 (I350065,I350017,I426875);
not I_20421 (I350082,I350065);
nor I_20422 (I349615,I349706,I350082);
nand I_20423 (I350113,I349808,I350082);
nand I_20424 (I349624,I349791,I350113);
nor I_20425 (I349621,I349689,I350065);
nand I_20426 (I350158,I350017,I349706);
not I_20427 (I350175,I350158);
DFFARX1 I_20428 (I350175,I2898,I349638,I349618,);
not I_20429 (I350233,I2905);
or I_20430 (I350250,I242907,I242886);
nand I_20431 (I350267,I242883,I242898);
not I_20432 (I350284,I350267);
nand I_20433 (I350301,I350284,I350250);
or I_20434 (I350318,I242895,I242886);
nor I_20435 (I350335,I350318,I242892);
nand I_20436 (I350352,I350284,I350335);
nor I_20437 (I350369,I350335,I350267);
not I_20438 (I350386,I350369);
not I_20439 (I350403,I350335);
nand I_20440 (I350222,I350301,I350403);
nor I_20441 (I350434,I242889,I242889);
nor I_20442 (I350451,I350434,I242910);
nor I_20443 (I350468,I350451,I350267);
nor I_20444 (I350485,I350403,I350451);
nor I_20445 (I350502,I242880,I242901);
nand I_20446 (I350519,I350502,I350468);
not I_20447 (I350536,I350519);
nor I_20448 (I350207,I350301,I350536);
nand I_20449 (I350204,I350519,I350352);
nand I_20450 (I350581,I350485,I350502);
nand I_20451 (I350225,I350519,I350581);
nand I_20452 (I350612,I242883,I242904);
not I_20453 (I350629,I350612);
nor I_20454 (I350201,I350629,I350267);
nor I_20455 (I350660,I350612,I242880);
not I_20456 (I350677,I350660);
nor I_20457 (I350210,I350301,I350677);
nand I_20458 (I350708,I350403,I350677);
nand I_20459 (I350219,I350386,I350708);
nor I_20460 (I350216,I350284,I350660);
nand I_20461 (I350753,I350612,I350301);
not I_20462 (I350770,I350753);
DFFARX1 I_20463 (I350770,I2898,I350233,I350213,);
not I_20464 (I350828,I2905);
or I_20465 (I350845,I2651,I1595);
nand I_20466 (I350862,I1755,I1931);
not I_20467 (I350879,I350862);
nand I_20468 (I350896,I350879,I350845);
or I_20469 (I350913,I2275,I2827);
nor I_20470 (I350930,I350913,I2755);
nand I_20471 (I350947,I350879,I350930);
nor I_20472 (I350964,I350930,I350862);
not I_20473 (I350981,I350964);
not I_20474 (I350998,I350930);
nand I_20475 (I350817,I350896,I350998);
nor I_20476 (I351029,I1779,I2035);
nor I_20477 (I351046,I351029,I2483);
nor I_20478 (I351063,I351046,I350862);
nor I_20479 (I351080,I350998,I351046);
nor I_20480 (I351097,I1843,I1739);
nand I_20481 (I351114,I351097,I351063);
not I_20482 (I351131,I351114);
nor I_20483 (I350802,I350896,I351131);
nand I_20484 (I350799,I351114,I350947);
nand I_20485 (I351176,I351080,I351097);
nand I_20486 (I350820,I351114,I351176);
nand I_20487 (I351207,I2523,I1771);
not I_20488 (I351224,I351207);
nor I_20489 (I350796,I351224,I350862);
nor I_20490 (I351255,I351207,I1747);
not I_20491 (I351272,I351255);
nor I_20492 (I350805,I350896,I351272);
nand I_20493 (I351303,I350998,I351272);
nand I_20494 (I350814,I350981,I351303);
nor I_20495 (I350811,I350879,I351255);
nand I_20496 (I351348,I351207,I350896);
not I_20497 (I351365,I351348);
DFFARX1 I_20498 (I351365,I2898,I350828,I350808,);
not I_20499 (I351423,I2905);
or I_20500 (I351440,I375187,I375184);
nand I_20501 (I351457,I375169,I375163);
not I_20502 (I351474,I351457);
nand I_20503 (I351491,I351474,I351440);
or I_20504 (I351508,I375190,I375157);
nor I_20505 (I351525,I351508,I375163);
nand I_20506 (I351542,I351474,I351525);
nor I_20507 (I351559,I351525,I351457);
not I_20508 (I351576,I351559);
not I_20509 (I351593,I351525);
nand I_20510 (I351412,I351491,I351593);
nor I_20511 (I351624,I375181,I375172);
nor I_20512 (I351641,I351624,I375175);
nor I_20513 (I351658,I351641,I351457);
nor I_20514 (I351675,I351593,I351641);
nor I_20515 (I351692,I375178,I375160);
nand I_20516 (I351709,I351692,I351658);
not I_20517 (I351726,I351709);
nor I_20518 (I351397,I351491,I351726);
nand I_20519 (I351394,I351709,I351542);
nand I_20520 (I351771,I351675,I351692);
nand I_20521 (I351415,I351709,I351771);
nand I_20522 (I351802,I375157,I375160);
not I_20523 (I351819,I351802);
nor I_20524 (I351391,I351819,I351457);
nor I_20525 (I351850,I351802,I375166);
not I_20526 (I351867,I351850);
nor I_20527 (I351400,I351491,I351867);
nand I_20528 (I351898,I351593,I351867);
nand I_20529 (I351409,I351576,I351898);
nor I_20530 (I351406,I351474,I351850);
nand I_20531 (I351943,I351802,I351491);
not I_20532 (I351960,I351943);
DFFARX1 I_20533 (I351960,I2898,I351423,I351403,);
not I_20534 (I352018,I2905);
or I_20535 (I352035,I112867,I112873);
nand I_20536 (I352052,I112885,I112876);
not I_20537 (I352069,I352052);
nand I_20538 (I352086,I352069,I352035);
or I_20539 (I352103,I112882,I112864);
nor I_20540 (I352120,I352103,I112897);
nand I_20541 (I352137,I352069,I352120);
nor I_20542 (I352154,I352120,I352052);
not I_20543 (I352171,I352154);
not I_20544 (I352188,I352120);
nand I_20545 (I352007,I352086,I352188);
nor I_20546 (I352219,I112867,I112870);
nor I_20547 (I352236,I352219,I112879);
nor I_20548 (I352253,I352236,I352052);
nor I_20549 (I352270,I352188,I352236);
nor I_20550 (I352287,I112888,I112870);
nand I_20551 (I352304,I352287,I352253);
not I_20552 (I352321,I352304);
nor I_20553 (I351992,I352086,I352321);
nand I_20554 (I351989,I352304,I352137);
nand I_20555 (I352366,I352270,I352287);
nand I_20556 (I352010,I352304,I352366);
nand I_20557 (I352397,I112894,I112891);
not I_20558 (I352414,I352397);
nor I_20559 (I351986,I352414,I352052);
nor I_20560 (I352445,I352397,I112864);
not I_20561 (I352462,I352445);
nor I_20562 (I351995,I352086,I352462);
nand I_20563 (I352493,I352188,I352462);
nand I_20564 (I352004,I352171,I352493);
nor I_20565 (I352001,I352069,I352445);
nand I_20566 (I352538,I352397,I352086);
not I_20567 (I352555,I352538);
DFFARX1 I_20568 (I352555,I2898,I352018,I351998,);
not I_20569 (I352613,I2905);
or I_20570 (I352630,I94701,I94674);
nand I_20571 (I352647,I94686,I94680);
not I_20572 (I352664,I352647);
nand I_20573 (I352681,I352664,I352630);
or I_20574 (I352698,I94683,I94698);
nor I_20575 (I352715,I352698,I94677);
nand I_20576 (I352732,I352664,I352715);
nor I_20577 (I352749,I352715,I352647);
not I_20578 (I352766,I352749);
not I_20579 (I352783,I352715);
nand I_20580 (I352602,I352681,I352783);
nor I_20581 (I352814,I94695,I94677);
nor I_20582 (I352831,I352814,I94683);
nor I_20583 (I352848,I352831,I352647);
nor I_20584 (I352865,I352783,I352831);
nor I_20585 (I352882,I94674,I94692);
nand I_20586 (I352899,I352882,I352848);
not I_20587 (I352916,I352899);
nor I_20588 (I352587,I352681,I352916);
nand I_20589 (I352584,I352899,I352732);
nand I_20590 (I352961,I352865,I352882);
nand I_20591 (I352605,I352899,I352961);
nand I_20592 (I352992,I94680,I94689);
not I_20593 (I353009,I352992);
nor I_20594 (I352581,I353009,I352647);
nor I_20595 (I353040,I352992,I94686);
not I_20596 (I353057,I353040);
nor I_20597 (I352590,I352681,I353057);
nand I_20598 (I353088,I352783,I353057);
nand I_20599 (I352599,I352766,I353088);
nor I_20600 (I352596,I352664,I353040);
nand I_20601 (I353133,I352992,I352681);
not I_20602 (I353150,I353133);
DFFARX1 I_20603 (I353150,I2898,I352613,I352593,);
not I_20604 (I353208,I2905);
or I_20605 (I353225,I443588,I443585);
nand I_20606 (I353242,I443591,I443609);
not I_20607 (I353259,I353242);
nand I_20608 (I353276,I353259,I353225);
or I_20609 (I353293,I443600,I443594);
nor I_20610 (I353310,I353293,I443615);
nand I_20611 (I353327,I353259,I353310);
nor I_20612 (I353344,I353310,I353242);
not I_20613 (I353361,I353344);
not I_20614 (I353378,I353310);
nand I_20615 (I353197,I353276,I353378);
nor I_20616 (I353409,I443582,I443606);
nor I_20617 (I353426,I353409,I443612);
nor I_20618 (I353443,I353426,I353242);
nor I_20619 (I353460,I353378,I353426);
nor I_20620 (I353477,I443582,I443585);
nand I_20621 (I353494,I353477,I353443);
not I_20622 (I353511,I353494);
nor I_20623 (I353182,I353276,I353511);
nand I_20624 (I353179,I353494,I353327);
nand I_20625 (I353556,I353460,I353477);
nand I_20626 (I353200,I353494,I353556);
nand I_20627 (I353587,I443588,I443597);
not I_20628 (I353604,I353587);
nor I_20629 (I353176,I353604,I353242);
nor I_20630 (I353635,I353587,I443603);
not I_20631 (I353652,I353635);
nor I_20632 (I353185,I353276,I353652);
nand I_20633 (I353683,I353378,I353652);
nand I_20634 (I353194,I353361,I353683);
nor I_20635 (I353191,I353259,I353635);
nand I_20636 (I353728,I353587,I353276);
not I_20637 (I353745,I353728);
DFFARX1 I_20638 (I353745,I2898,I353208,I353188,);
not I_20639 (I353803,I2905);
or I_20640 (I353820,I240612,I240591);
nand I_20641 (I353837,I240588,I240603);
not I_20642 (I353854,I353837);
nand I_20643 (I353871,I353854,I353820);
or I_20644 (I353888,I240600,I240591);
nor I_20645 (I353905,I353888,I240597);
nand I_20646 (I353922,I353854,I353905);
nor I_20647 (I353939,I353905,I353837);
not I_20648 (I353956,I353939);
not I_20649 (I353973,I353905);
nand I_20650 (I353792,I353871,I353973);
nor I_20651 (I354004,I240594,I240594);
nor I_20652 (I354021,I354004,I240615);
nor I_20653 (I354038,I354021,I353837);
nor I_20654 (I354055,I353973,I354021);
nor I_20655 (I354072,I240585,I240606);
nand I_20656 (I354089,I354072,I354038);
not I_20657 (I354106,I354089);
nor I_20658 (I353777,I353871,I354106);
nand I_20659 (I353774,I354089,I353922);
nand I_20660 (I354151,I354055,I354072);
nand I_20661 (I353795,I354089,I354151);
nand I_20662 (I354182,I240588,I240609);
not I_20663 (I354199,I354182);
nor I_20664 (I353771,I354199,I353837);
nor I_20665 (I354230,I354182,I240585);
not I_20666 (I354247,I354230);
nor I_20667 (I353780,I353871,I354247);
nand I_20668 (I354278,I353973,I354247);
nand I_20669 (I353789,I353956,I354278);
nor I_20670 (I353786,I353854,I354230);
nand I_20671 (I354323,I354182,I353871);
not I_20672 (I354340,I354323);
DFFARX1 I_20673 (I354340,I2898,I353803,I353783,);
not I_20674 (I354398,I2905);
or I_20675 (I354415,I122931,I122937);
nand I_20676 (I354432,I122949,I122940);
not I_20677 (I354449,I354432);
nand I_20678 (I354466,I354449,I354415);
or I_20679 (I354483,I122946,I122928);
nor I_20680 (I354500,I354483,I122961);
nand I_20681 (I354517,I354449,I354500);
nor I_20682 (I354534,I354500,I354432);
not I_20683 (I354551,I354534);
not I_20684 (I354568,I354500);
nand I_20685 (I354387,I354466,I354568);
nor I_20686 (I354599,I122931,I122934);
nor I_20687 (I354616,I354599,I122943);
nor I_20688 (I354633,I354616,I354432);
nor I_20689 (I354650,I354568,I354616);
nor I_20690 (I354667,I122952,I122934);
nand I_20691 (I354684,I354667,I354633);
not I_20692 (I354701,I354684);
nor I_20693 (I354372,I354466,I354701);
nand I_20694 (I354369,I354684,I354517);
nand I_20695 (I354746,I354650,I354667);
nand I_20696 (I354390,I354684,I354746);
nand I_20697 (I354777,I122958,I122955);
not I_20698 (I354794,I354777);
nor I_20699 (I354366,I354794,I354432);
nor I_20700 (I354825,I354777,I122928);
not I_20701 (I354842,I354825);
nor I_20702 (I354375,I354466,I354842);
nand I_20703 (I354873,I354568,I354842);
nand I_20704 (I354384,I354551,I354873);
nor I_20705 (I354381,I354449,I354825);
nand I_20706 (I354918,I354777,I354466);
not I_20707 (I354935,I354918);
DFFARX1 I_20708 (I354935,I2898,I354398,I354378,);
not I_20709 (I354993,I2905);
or I_20710 (I355010,I79605,I79578);
nand I_20711 (I355027,I79590,I79584);
not I_20712 (I355044,I355027);
nand I_20713 (I355061,I355044,I355010);
or I_20714 (I355078,I79587,I79602);
nor I_20715 (I355095,I355078,I79581);
nand I_20716 (I355112,I355044,I355095);
nor I_20717 (I355129,I355095,I355027);
not I_20718 (I355146,I355129);
not I_20719 (I355163,I355095);
nand I_20720 (I354982,I355061,I355163);
nor I_20721 (I355194,I79599,I79581);
nor I_20722 (I355211,I355194,I79587);
nor I_20723 (I355228,I355211,I355027);
nor I_20724 (I355245,I355163,I355211);
nor I_20725 (I355262,I79578,I79596);
nand I_20726 (I355279,I355262,I355228);
not I_20727 (I355296,I355279);
nor I_20728 (I354967,I355061,I355296);
nand I_20729 (I354964,I355279,I355112);
nand I_20730 (I355341,I355245,I355262);
nand I_20731 (I354985,I355279,I355341);
nand I_20732 (I355372,I79584,I79593);
not I_20733 (I355389,I355372);
nor I_20734 (I354961,I355389,I355027);
nor I_20735 (I355420,I355372,I79590);
not I_20736 (I355437,I355420);
nor I_20737 (I354970,I355061,I355437);
nand I_20738 (I355468,I355163,I355437);
nand I_20739 (I354979,I355146,I355468);
nor I_20740 (I354976,I355044,I355420);
nand I_20741 (I355513,I355372,I355061);
not I_20742 (I355530,I355513);
DFFARX1 I_20743 (I355530,I2898,I354993,I354973,);
not I_20744 (I355588,I2905);
or I_20745 (I355605,I432436,I432433);
nand I_20746 (I355622,I432439,I432457);
not I_20747 (I355639,I355622);
nand I_20748 (I355656,I355639,I355605);
or I_20749 (I355673,I432448,I432442);
nor I_20750 (I355690,I355673,I432463);
nand I_20751 (I355707,I355639,I355690);
nor I_20752 (I355724,I355690,I355622);
not I_20753 (I355741,I355724);
not I_20754 (I355758,I355690);
nand I_20755 (I355577,I355656,I355758);
nor I_20756 (I355789,I432430,I432454);
nor I_20757 (I355806,I355789,I432460);
nor I_20758 (I355823,I355806,I355622);
nor I_20759 (I355840,I355758,I355806);
nor I_20760 (I355857,I432430,I432433);
nand I_20761 (I355874,I355857,I355823);
not I_20762 (I355891,I355874);
nor I_20763 (I355562,I355656,I355891);
nand I_20764 (I355559,I355874,I355707);
nand I_20765 (I355936,I355840,I355857);
nand I_20766 (I355580,I355874,I355936);
nand I_20767 (I355967,I432436,I432445);
not I_20768 (I355984,I355967);
nor I_20769 (I355556,I355984,I355622);
nor I_20770 (I356015,I355967,I432451);
not I_20771 (I356032,I356015);
nor I_20772 (I355565,I355656,I356032);
nand I_20773 (I356063,I355758,I356032);
nand I_20774 (I355574,I355741,I356063);
nor I_20775 (I355571,I355639,I356015);
nand I_20776 (I356108,I355967,I355656);
not I_20777 (I356125,I356108);
DFFARX1 I_20778 (I356125,I2898,I355588,I355568,);
not I_20779 (I356183,I2905);
or I_20780 (I356200,I163375,I163354);
nand I_20781 (I356217,I163360,I163378);
not I_20782 (I356234,I356217);
nand I_20783 (I356251,I356234,I356200);
or I_20784 (I356268,I163354,I163369);
nor I_20785 (I356285,I356268,I163366);
nand I_20786 (I356302,I356234,I356285);
nor I_20787 (I356319,I356285,I356217);
not I_20788 (I356336,I356319);
not I_20789 (I356353,I356285);
nand I_20790 (I356172,I356251,I356353);
nor I_20791 (I356384,I163372,I163384);
nor I_20792 (I356401,I356384,I163357);
nor I_20793 (I356418,I356401,I356217);
nor I_20794 (I356435,I356353,I356401);
nor I_20795 (I356452,I163363,I163381);
nand I_20796 (I356469,I356452,I356418);
not I_20797 (I356486,I356469);
nor I_20798 (I356157,I356251,I356486);
nand I_20799 (I356154,I356469,I356302);
nand I_20800 (I356531,I356435,I356452);
nand I_20801 (I356175,I356469,I356531);
nand I_20802 (I356562,I163357,I163387);
not I_20803 (I356579,I356562);
nor I_20804 (I356151,I356579,I356217);
nor I_20805 (I356610,I356562,I163360);
not I_20806 (I356627,I356610);
nor I_20807 (I356160,I356251,I356627);
nand I_20808 (I356658,I356353,I356627);
nand I_20809 (I356169,I356336,I356658);
nor I_20810 (I356166,I356234,I356610);
nand I_20811 (I356703,I356562,I356251);
not I_20812 (I356720,I356703);
DFFARX1 I_20813 (I356720,I2898,I356183,I356163,);
not I_20814 (I356778,I2905);
or I_20815 (I356795,I119786,I119792);
nand I_20816 (I356812,I119804,I119795);
not I_20817 (I356829,I356812);
nand I_20818 (I356846,I356829,I356795);
or I_20819 (I356863,I119801,I119783);
nor I_20820 (I356880,I356863,I119816);
nand I_20821 (I356897,I356829,I356880);
nor I_20822 (I356914,I356880,I356812);
not I_20823 (I356931,I356914);
not I_20824 (I356948,I356880);
nand I_20825 (I356767,I356846,I356948);
nor I_20826 (I356979,I119786,I119789);
nor I_20827 (I356996,I356979,I119798);
nor I_20828 (I357013,I356996,I356812);
nor I_20829 (I357030,I356948,I356996);
nor I_20830 (I357047,I119807,I119789);
nand I_20831 (I357064,I357047,I357013);
not I_20832 (I357081,I357064);
nor I_20833 (I356752,I356846,I357081);
nand I_20834 (I356749,I357064,I356897);
nand I_20835 (I357126,I357030,I357047);
nand I_20836 (I356770,I357064,I357126);
nand I_20837 (I357157,I119813,I119810);
not I_20838 (I357174,I357157);
nor I_20839 (I356746,I357174,I356812);
nor I_20840 (I357205,I357157,I119783);
not I_20841 (I357222,I357205);
nor I_20842 (I356755,I356846,I357222);
nand I_20843 (I357253,I356948,I357222);
nand I_20844 (I356764,I356931,I357253);
nor I_20845 (I356761,I356829,I357205);
nand I_20846 (I357298,I357157,I356846);
not I_20847 (I357315,I357298);
DFFARX1 I_20848 (I357315,I2898,I356778,I356758,);
not I_20849 (I357373,I2905);
or I_20850 (I357390,I139914,I139920);
nand I_20851 (I357407,I139932,I139923);
not I_20852 (I357424,I357407);
nand I_20853 (I357441,I357424,I357390);
or I_20854 (I357458,I139929,I139911);
nor I_20855 (I357475,I357458,I139944);
nand I_20856 (I357492,I357424,I357475);
nor I_20857 (I357509,I357475,I357407);
not I_20858 (I357526,I357509);
not I_20859 (I357543,I357475);
nand I_20860 (I357362,I357441,I357543);
nor I_20861 (I357574,I139914,I139917);
nor I_20862 (I357591,I357574,I139926);
nor I_20863 (I357608,I357591,I357407);
nor I_20864 (I357625,I357543,I357591);
nor I_20865 (I357642,I139935,I139917);
nand I_20866 (I357659,I357642,I357608);
not I_20867 (I357676,I357659);
nor I_20868 (I357347,I357441,I357676);
nand I_20869 (I357344,I357659,I357492);
nand I_20870 (I357721,I357625,I357642);
nand I_20871 (I357365,I357659,I357721);
nand I_20872 (I357752,I139941,I139938);
not I_20873 (I357769,I357752);
nor I_20874 (I357341,I357769,I357407);
nor I_20875 (I357800,I357752,I139911);
not I_20876 (I357817,I357800);
nor I_20877 (I357350,I357441,I357817);
nand I_20878 (I357848,I357543,I357817);
nand I_20879 (I357359,I357526,I357848);
nor I_20880 (I357356,I357424,I357800);
nand I_20881 (I357893,I357752,I357441);
not I_20882 (I357910,I357893);
DFFARX1 I_20883 (I357910,I2898,I357373,I357353,);
not I_20884 (I357968,I2905);
or I_20885 (I357985,I104061,I104067);
nand I_20886 (I358002,I104079,I104070);
not I_20887 (I358019,I358002);
nand I_20888 (I358036,I358019,I357985);
or I_20889 (I358053,I104076,I104058);
nor I_20890 (I358070,I358053,I104091);
nand I_20891 (I358087,I358019,I358070);
nor I_20892 (I358104,I358070,I358002);
not I_20893 (I358121,I358104);
not I_20894 (I358138,I358070);
nand I_20895 (I357957,I358036,I358138);
nor I_20896 (I358169,I104061,I104064);
nor I_20897 (I358186,I358169,I104073);
nor I_20898 (I358203,I358186,I358002);
nor I_20899 (I358220,I358138,I358186);
nor I_20900 (I358237,I104082,I104064);
nand I_20901 (I358254,I358237,I358203);
not I_20902 (I358271,I358254);
nor I_20903 (I357942,I358036,I358271);
nand I_20904 (I357939,I358254,I358087);
nand I_20905 (I358316,I358220,I358237);
nand I_20906 (I357960,I358254,I358316);
nand I_20907 (I358347,I104088,I104085);
not I_20908 (I358364,I358347);
nor I_20909 (I357936,I358364,I358002);
nor I_20910 (I358395,I358347,I104058);
not I_20911 (I358412,I358395);
nor I_20912 (I357945,I358036,I358412);
nand I_20913 (I358443,I358138,I358412);
nand I_20914 (I357954,I358121,I358443);
nor I_20915 (I357951,I358019,I358395);
nand I_20916 (I358488,I358347,I358036);
not I_20917 (I358505,I358488);
DFFARX1 I_20918 (I358505,I2898,I357968,I357948,);
not I_20919 (I358563,I2905);
or I_20920 (I358580,I129221,I129227);
nand I_20921 (I358597,I129239,I129230);
not I_20922 (I358614,I358597);
nand I_20923 (I358631,I358614,I358580);
or I_20924 (I358648,I129236,I129218);
nor I_20925 (I358665,I358648,I129251);
nand I_20926 (I358682,I358614,I358665);
nor I_20927 (I358699,I358665,I358597);
not I_20928 (I358716,I358699);
not I_20929 (I358733,I358665);
nand I_20930 (I358552,I358631,I358733);
nor I_20931 (I358764,I129221,I129224);
nor I_20932 (I358781,I358764,I129233);
nor I_20933 (I358798,I358781,I358597);
nor I_20934 (I358815,I358733,I358781);
nor I_20935 (I358832,I129242,I129224);
nand I_20936 (I358849,I358832,I358798);
not I_20937 (I358866,I358849);
nor I_20938 (I358537,I358631,I358866);
nand I_20939 (I358534,I358849,I358682);
nand I_20940 (I358911,I358815,I358832);
nand I_20941 (I358555,I358849,I358911);
nand I_20942 (I358942,I129248,I129245);
not I_20943 (I358959,I358942);
nor I_20944 (I358531,I358959,I358597);
nor I_20945 (I358990,I358942,I129218);
not I_20946 (I359007,I358990);
nor I_20947 (I358540,I358631,I359007);
nand I_20948 (I359038,I358733,I359007);
nand I_20949 (I358549,I358716,I359038);
nor I_20950 (I358546,I358614,I358990);
nand I_20951 (I359083,I358942,I358631);
not I_20952 (I359100,I359083);
DFFARX1 I_20953 (I359100,I2898,I358563,I358543,);
not I_20954 (I359158,I2905);
or I_20955 (I359175,I121673,I121679);
nand I_20956 (I359192,I121691,I121682);
not I_20957 (I359209,I359192);
nand I_20958 (I359226,I359209,I359175);
or I_20959 (I359243,I121688,I121670);
nor I_20960 (I359260,I359243,I121703);
nand I_20961 (I359277,I359209,I359260);
nor I_20962 (I359294,I359260,I359192);
not I_20963 (I359311,I359294);
not I_20964 (I359328,I359260);
nand I_20965 (I359147,I359226,I359328);
nor I_20966 (I359359,I121673,I121676);
nor I_20967 (I359376,I359359,I121685);
nor I_20968 (I359393,I359376,I359192);
nor I_20969 (I359410,I359328,I359376);
nor I_20970 (I359427,I121694,I121676);
nand I_20971 (I359444,I359427,I359393);
not I_20972 (I359461,I359444);
nor I_20973 (I359132,I359226,I359461);
nand I_20974 (I359129,I359444,I359277);
nand I_20975 (I359506,I359410,I359427);
nand I_20976 (I359150,I359444,I359506);
nand I_20977 (I359537,I121700,I121697);
not I_20978 (I359554,I359537);
nor I_20979 (I359126,I359554,I359192);
nor I_20980 (I359585,I359537,I121670);
not I_20981 (I359602,I359585);
nor I_20982 (I359135,I359226,I359602);
nand I_20983 (I359633,I359328,I359602);
nand I_20984 (I359144,I359311,I359633);
nor I_20985 (I359141,I359209,I359585);
nand I_20986 (I359678,I359537,I359226);
not I_20987 (I359695,I359678);
DFFARX1 I_20988 (I359695,I2898,I359158,I359138,);
not I_20989 (I359753,I2905);
or I_20990 (I359770,I123560,I123566);
nand I_20991 (I359787,I123578,I123569);
not I_20992 (I359804,I359787);
nand I_20993 (I359821,I359804,I359770);
or I_20994 (I359838,I123575,I123557);
nor I_20995 (I359855,I359838,I123590);
nand I_20996 (I359872,I359804,I359855);
nor I_20997 (I359889,I359855,I359787);
not I_20998 (I359906,I359889);
not I_20999 (I359923,I359855);
nand I_21000 (I359742,I359821,I359923);
nor I_21001 (I359954,I123560,I123563);
nor I_21002 (I359971,I359954,I123572);
nor I_21003 (I359988,I359971,I359787);
nor I_21004 (I360005,I359923,I359971);
nor I_21005 (I360022,I123581,I123563);
nand I_21006 (I360039,I360022,I359988);
not I_21007 (I360056,I360039);
nor I_21008 (I359727,I359821,I360056);
nand I_21009 (I359724,I360039,I359872);
nand I_21010 (I360101,I360005,I360022);
nand I_21011 (I359745,I360039,I360101);
nand I_21012 (I360132,I123587,I123584);
not I_21013 (I360149,I360132);
nor I_21014 (I359721,I360149,I359787);
nor I_21015 (I360180,I360132,I123557);
not I_21016 (I360197,I360180);
nor I_21017 (I359730,I359821,I360197);
nand I_21018 (I360228,I359923,I360197);
nand I_21019 (I359739,I359906,I360228);
nor I_21020 (I359736,I359804,I360180);
nand I_21021 (I360273,I360132,I359821);
not I_21022 (I360290,I360273);
DFFARX1 I_21023 (I360290,I2898,I359753,I359733,);
not I_21024 (I360348,I2905);
or I_21025 (I360365,I112238,I112244);
nand I_21026 (I360382,I112256,I112247);
not I_21027 (I360399,I360382);
nand I_21028 (I360416,I360399,I360365);
or I_21029 (I360433,I112253,I112235);
nor I_21030 (I360450,I360433,I112268);
nand I_21031 (I360467,I360399,I360450);
nor I_21032 (I360484,I360450,I360382);
not I_21033 (I360501,I360484);
not I_21034 (I360518,I360450);
nand I_21035 (I360337,I360416,I360518);
nor I_21036 (I360549,I112238,I112241);
nor I_21037 (I360566,I360549,I112250);
nor I_21038 (I360583,I360566,I360382);
nor I_21039 (I360600,I360518,I360566);
nor I_21040 (I360617,I112259,I112241);
nand I_21041 (I360634,I360617,I360583);
not I_21042 (I360651,I360634);
nor I_21043 (I360322,I360416,I360651);
nand I_21044 (I360319,I360634,I360467);
nand I_21045 (I360696,I360600,I360617);
nand I_21046 (I360340,I360634,I360696);
nand I_21047 (I360727,I112265,I112262);
not I_21048 (I360744,I360727);
nor I_21049 (I360316,I360744,I360382);
nor I_21050 (I360775,I360727,I112235);
not I_21051 (I360792,I360775);
nor I_21052 (I360325,I360416,I360792);
nand I_21053 (I360823,I360518,I360792);
nand I_21054 (I360334,I360501,I360823);
nor I_21055 (I360331,I360399,I360775);
nand I_21056 (I360868,I360727,I360416);
not I_21057 (I360885,I360868);
DFFARX1 I_21058 (I360885,I2898,I360348,I360328,);
not I_21059 (I360943,I2905);
or I_21060 (I360960,I264327,I264306);
nand I_21061 (I360977,I264303,I264318);
not I_21062 (I360994,I360977);
nand I_21063 (I361011,I360994,I360960);
or I_21064 (I361028,I264315,I264306);
nor I_21065 (I361045,I361028,I264312);
nand I_21066 (I361062,I360994,I361045);
nor I_21067 (I361079,I361045,I360977);
not I_21068 (I361096,I361079);
not I_21069 (I361113,I361045);
nand I_21070 (I360932,I361011,I361113);
nor I_21071 (I361144,I264309,I264309);
nor I_21072 (I361161,I361144,I264330);
nor I_21073 (I361178,I361161,I360977);
nor I_21074 (I361195,I361113,I361161);
nor I_21075 (I361212,I264300,I264321);
nand I_21076 (I361229,I361212,I361178);
not I_21077 (I361246,I361229);
nor I_21078 (I360917,I361011,I361246);
nand I_21079 (I360914,I361229,I361062);
nand I_21080 (I361291,I361195,I361212);
nand I_21081 (I360935,I361229,I361291);
nand I_21082 (I361322,I264303,I264324);
not I_21083 (I361339,I361322);
nor I_21084 (I360911,I361339,I360977);
nor I_21085 (I361370,I361322,I264300);
not I_21086 (I361387,I361370);
nor I_21087 (I360920,I361011,I361387);
nand I_21088 (I361418,I361113,I361387);
nand I_21089 (I360929,I361096,I361418);
nor I_21090 (I360926,I360994,I361370);
nand I_21091 (I361463,I361322,I361011);
not I_21092 (I361480,I361463);
DFFARX1 I_21093 (I361480,I2898,I360943,I360923,);
not I_21094 (I361538,I2905);
or I_21095 (I361555,I302505,I302517);
nand I_21096 (I361572,I302523,I302520);
not I_21097 (I361589,I361572);
nand I_21098 (I361606,I361589,I361555);
or I_21099 (I361623,I302514,I302499);
nor I_21100 (I361640,I361623,I302529);
nand I_21101 (I361657,I361589,I361640);
nor I_21102 (I361674,I361640,I361572);
not I_21103 (I361691,I361674);
not I_21104 (I361708,I361640);
nand I_21105 (I361527,I361606,I361708);
nor I_21106 (I361739,I302526,I302508);
nor I_21107 (I361756,I361739,I302502);
nor I_21108 (I361773,I361756,I361572);
nor I_21109 (I361790,I361708,I361756);
nor I_21110 (I361807,I302505,I302508);
nand I_21111 (I361824,I361807,I361773);
not I_21112 (I361841,I361824);
nor I_21113 (I361512,I361606,I361841);
nand I_21114 (I361509,I361824,I361657);
nand I_21115 (I361886,I361790,I361807);
nand I_21116 (I361530,I361824,I361886);
nand I_21117 (I361917,I302499,I302511);
not I_21118 (I361934,I361917);
nor I_21119 (I361506,I361934,I361572);
nor I_21120 (I361965,I361917,I302502);
not I_21121 (I361982,I361965);
nor I_21122 (I361515,I361606,I361982);
nand I_21123 (I362013,I361708,I361982);
nand I_21124 (I361524,I361691,I362013);
nor I_21125 (I361521,I361589,I361965);
nand I_21126 (I362058,I361917,I361606);
not I_21127 (I362075,I362058);
DFFARX1 I_21128 (I362075,I2898,I361538,I361518,);
not I_21129 (I362133,I2905);
or I_21130 (I362150,I286423,I286435);
nand I_21131 (I362167,I286441,I286438);
not I_21132 (I362184,I362167);
nand I_21133 (I362201,I362184,I362150);
or I_21134 (I362218,I286432,I286417);
nor I_21135 (I362235,I362218,I286447);
nand I_21136 (I362252,I362184,I362235);
nor I_21137 (I362269,I362235,I362167);
not I_21138 (I362286,I362269);
not I_21139 (I362303,I362235);
nand I_21140 (I362122,I362201,I362303);
nor I_21141 (I362334,I286444,I286426);
nor I_21142 (I362351,I362334,I286420);
nor I_21143 (I362368,I362351,I362167);
nor I_21144 (I362385,I362303,I362351);
nor I_21145 (I362402,I286423,I286426);
nand I_21146 (I362419,I362402,I362368);
not I_21147 (I362436,I362419);
nor I_21148 (I362107,I362201,I362436);
nand I_21149 (I362104,I362419,I362252);
nand I_21150 (I362481,I362385,I362402);
nand I_21151 (I362125,I362419,I362481);
nand I_21152 (I362512,I286417,I286429);
not I_21153 (I362529,I362512);
nor I_21154 (I362101,I362529,I362167);
nor I_21155 (I362560,I362512,I286420);
not I_21156 (I362577,I362560);
nor I_21157 (I362110,I362201,I362577);
nand I_21158 (I362608,I362303,I362577);
nand I_21159 (I362119,I362286,I362608);
nor I_21160 (I362116,I362184,I362560);
nand I_21161 (I362653,I362512,I362201);
not I_21162 (I362670,I362653);
DFFARX1 I_21163 (I362670,I2898,I362133,I362113,);
not I_21164 (I362728,I2905);
or I_21165 (I362745,I262032,I262011);
nand I_21166 (I362762,I262008,I262023);
not I_21167 (I362779,I362762);
nand I_21168 (I362796,I362779,I362745);
or I_21169 (I362813,I262020,I262011);
nor I_21170 (I362830,I362813,I262017);
nand I_21171 (I362847,I362779,I362830);
nor I_21172 (I362864,I362830,I362762);
not I_21173 (I362881,I362864);
not I_21174 (I362898,I362830);
nand I_21175 (I362717,I362796,I362898);
nor I_21176 (I362929,I262014,I262014);
nor I_21177 (I362946,I362929,I262035);
nor I_21178 (I362963,I362946,I362762);
nor I_21179 (I362980,I362898,I362946);
nor I_21180 (I362997,I262005,I262026);
nand I_21181 (I363014,I362997,I362963);
not I_21182 (I363031,I363014);
nor I_21183 (I362702,I362796,I363031);
nand I_21184 (I362699,I363014,I362847);
nand I_21185 (I363076,I362980,I362997);
nand I_21186 (I362720,I363014,I363076);
nand I_21187 (I363107,I262008,I262029);
not I_21188 (I363124,I363107);
nor I_21189 (I362696,I363124,I362762);
nor I_21190 (I363155,I363107,I262005);
not I_21191 (I363172,I363155);
nor I_21192 (I362705,I362796,I363172);
nand I_21193 (I363203,I362898,I363172);
nand I_21194 (I362714,I362881,I363203);
nor I_21195 (I362711,I362779,I363155);
nand I_21196 (I363248,I363107,I362796);
not I_21197 (I363265,I363248);
DFFARX1 I_21198 (I363265,I2898,I362728,I362708,);
not I_21199 (I363332,I2905);
or I_21200 (I363349,I157926,I157932);
nand I_21201 (I363366,I157914,I157917);
not I_21202 (I363383,I363366);
nand I_21203 (I363400,I363383,I363349);
not I_21204 (I363417,I363400);
nor I_21205 (I363434,I157941,I157923);
not I_21206 (I363451,I363434);
nor I_21207 (I363468,I363383,I363451);
not I_21208 (I363485,I157938);
nor I_21209 (I363502,I363451,I157920);
nor I_21210 (I363294,I363366,I363502);
nor I_21211 (I363533,I157920,I157941);
not I_21212 (I363550,I157944);
nor I_21213 (I363567,I157914,I157938);
nand I_21214 (I363306,I363468,I363567);
not I_21215 (I363598,I157914);
nand I_21216 (I363615,I363598,I363485);
nor I_21217 (I363632,I363550,I157914);
nor I_21218 (I363649,I363632,I157923);
nor I_21219 (I363312,I363417,I363649);
nor I_21220 (I363680,I363632,I363400);
nand I_21221 (I363303,I363434,I363680);
nor I_21222 (I363711,I157947,I157917);
DFFARX1 I_21223 (I363711,I2898,I363332,I363737,);
not I_21224 (I363745,I363737);
not I_21225 (I363762,I157947);
nor I_21226 (I363779,I157947,I157920);
or I_21227 (I363796,I157947,I157920);
nand I_21228 (I363321,I363615,I363796);
nand I_21229 (I363827,I363745,I157920);
nand I_21230 (I363844,I157935,I157929);
nor I_21231 (I363861,I363844,I157920);
nor I_21232 (I363291,I363366,I363861);
nand I_21233 (I363892,I363745,I363844);
not I_21234 (I363909,I363892);
DFFARX1 I_21235 (I363909,I2898,I363332,I363309,);
nand I_21236 (I363324,I363892,I363827);
nor I_21237 (I363954,I363844,I363417);
not I_21238 (I363297,I363954);
nor I_21239 (I363318,I363954,I363779);
nor I_21240 (I363999,I363844,I363762);
nand I_21241 (I364016,I363737,I363999);
nand I_21242 (I364033,I363533,I364016);
DFFARX1 I_21243 (I364033,I2898,I363332,I363300,);
or I_21244 (I364064,I363844,I157920);
nand I_21245 (I363315,I363615,I364064);
not I_21246 (I364131,I2905);
or I_21247 (I364148,I65120,I65117);
nand I_21248 (I364165,I65138,I65111);
not I_21249 (I364182,I364165);
nand I_21250 (I364199,I364182,I364148);
not I_21251 (I364216,I364199);
nor I_21252 (I364233,I65114,I65120);
not I_21253 (I364250,I364233);
nor I_21254 (I364267,I364182,I364250);
not I_21255 (I364284,I65111);
nor I_21256 (I364301,I364250,I65129);
nor I_21257 (I364093,I364165,I364301);
nor I_21258 (I364332,I65129,I65114);
not I_21259 (I364349,I65132);
nor I_21260 (I364366,I65123,I65111);
nand I_21261 (I364105,I364267,I364366);
not I_21262 (I364397,I65123);
nand I_21263 (I364414,I364397,I364284);
nor I_21264 (I364431,I364349,I65123);
nor I_21265 (I364448,I364431,I65120);
nor I_21266 (I364111,I364216,I364448);
nor I_21267 (I364479,I364431,I364199);
nand I_21268 (I364102,I364233,I364479);
nor I_21269 (I364510,I65117,I65114);
DFFARX1 I_21270 (I364510,I2898,I364131,I364536,);
not I_21271 (I364544,I364536);
not I_21272 (I364561,I65117);
nor I_21273 (I364578,I65117,I65129);
or I_21274 (I364595,I65117,I65129);
nand I_21275 (I364120,I364414,I364595);
nand I_21276 (I364626,I364544,I65135);
nand I_21277 (I364643,I65123,I65126);
nor I_21278 (I364660,I364643,I65135);
nor I_21279 (I364090,I364165,I364660);
nand I_21280 (I364691,I364544,I364643);
not I_21281 (I364708,I364691);
DFFARX1 I_21282 (I364708,I2898,I364131,I364108,);
nand I_21283 (I364123,I364691,I364626);
nor I_21284 (I364753,I364643,I364216);
not I_21285 (I364096,I364753);
nor I_21286 (I364117,I364753,I364578);
nor I_21287 (I364798,I364643,I364561);
nand I_21288 (I364815,I364536,I364798);
nand I_21289 (I364832,I364332,I364815);
DFFARX1 I_21290 (I364832,I2898,I364131,I364099,);
or I_21291 (I364863,I364643,I65135);
nand I_21292 (I364114,I364414,I364863);
not I_21293 (I364930,I2905);
or I_21294 (I364947,I201573,I201585);
nand I_21295 (I364964,I201579,I201582);
not I_21296 (I364981,I364964);
nand I_21297 (I364998,I364981,I364947);
not I_21298 (I365015,I364998);
nor I_21299 (I365032,I201591,I201588);
not I_21300 (I365049,I365032);
nor I_21301 (I365066,I364981,I365049);
not I_21302 (I365083,I201585);
nor I_21303 (I365100,I365049,I201576);
nor I_21304 (I364892,I364964,I365100);
nor I_21305 (I365131,I201576,I201591);
not I_21306 (I365148,I201579);
nor I_21307 (I365165,I201573,I201585);
nand I_21308 (I364904,I365066,I365165);
not I_21309 (I365196,I201573);
nand I_21310 (I365213,I365196,I365083);
nor I_21311 (I365230,I365148,I201573);
nor I_21312 (I365247,I365230,I201588);
nor I_21313 (I364910,I365015,I365247);
nor I_21314 (I365278,I365230,I364998);
nand I_21315 (I364901,I365032,I365278);
nor I_21316 (I365309,I201570,I201594);
DFFARX1 I_21317 (I365309,I2898,I364930,I365335,);
not I_21318 (I365343,I365335);
not I_21319 (I365360,I201570);
nor I_21320 (I365377,I201570,I201576);
or I_21321 (I365394,I201570,I201576);
nand I_21322 (I364919,I365213,I365394);
nand I_21323 (I365425,I365343,I201570);
nand I_21324 (I365442,I201582,I201576);
nor I_21325 (I365459,I365442,I201570);
nor I_21326 (I364889,I364964,I365459);
nand I_21327 (I365490,I365343,I365442);
not I_21328 (I365507,I365490);
DFFARX1 I_21329 (I365507,I2898,I364930,I364907,);
nand I_21330 (I364922,I365490,I365425);
nor I_21331 (I365552,I365442,I365015);
not I_21332 (I364895,I365552);
nor I_21333 (I364916,I365552,I365377);
nor I_21334 (I365597,I365442,I365360);
nand I_21335 (I365614,I365335,I365597);
nand I_21336 (I365631,I365131,I365614);
DFFARX1 I_21337 (I365631,I2898,I364930,I364898,);
or I_21338 (I365662,I365442,I201570);
nand I_21339 (I364913,I365213,I365662);
not I_21340 (I365729,I2905);
or I_21341 (I365746,I337114,I337123);
nand I_21342 (I365763,I337120,I337129);
not I_21343 (I365780,I365763);
nand I_21344 (I365797,I365780,I365746);
not I_21345 (I365814,I365797);
nor I_21346 (I365831,I337135,I337123);
not I_21347 (I365848,I365831);
nor I_21348 (I365865,I365780,I365848);
not I_21349 (I365882,I337111);
nor I_21350 (I365899,I365848,I337132);
nor I_21351 (I365691,I365763,I365899);
nor I_21352 (I365930,I337132,I337135);
not I_21353 (I365947,I337111);
nor I_21354 (I365964,I337114,I337111);
nand I_21355 (I365703,I365865,I365964);
not I_21356 (I365995,I337114);
nand I_21357 (I366012,I365995,I365882);
nor I_21358 (I366029,I365947,I337114);
nor I_21359 (I366046,I366029,I337123);
nor I_21360 (I365709,I365814,I366046);
nor I_21361 (I366077,I366029,I365797);
nand I_21362 (I365700,I365831,I366077);
nor I_21363 (I366108,I337120,I337126);
DFFARX1 I_21364 (I366108,I2898,I365729,I366134,);
not I_21365 (I366142,I366134);
not I_21366 (I366159,I337120);
nor I_21367 (I366176,I337120,I337132);
or I_21368 (I366193,I337120,I337132);
nand I_21369 (I365718,I366012,I366193);
nand I_21370 (I366224,I366142,I337126);
nand I_21371 (I366241,I337117,I337117);
nor I_21372 (I366258,I366241,I337126);
nor I_21373 (I365688,I365763,I366258);
nand I_21374 (I366289,I366142,I366241);
not I_21375 (I366306,I366289);
DFFARX1 I_21376 (I366306,I2898,I365729,I365706,);
nand I_21377 (I365721,I366289,I366224);
nor I_21378 (I366351,I366241,I365814);
not I_21379 (I365694,I366351);
nor I_21380 (I365715,I366351,I366176);
nor I_21381 (I366396,I366241,I366159);
nand I_21382 (I366413,I366134,I366396);
nand I_21383 (I366430,I365930,I366413);
DFFARX1 I_21384 (I366430,I2898,I365729,I365697,);
or I_21385 (I366461,I366241,I337126);
nand I_21386 (I365712,I366012,I366461);
not I_21387 (I366528,I2905);
or I_21388 (I366545,I430369,I430351);
nand I_21389 (I366562,I430366,I430360);
not I_21390 (I366579,I366562);
nand I_21391 (I366596,I366579,I366545);
not I_21392 (I366613,I366596);
nor I_21393 (I366630,I430345,I430372);
not I_21394 (I366647,I366630);
nor I_21395 (I366664,I366579,I366647);
not I_21396 (I366681,I430342);
nor I_21397 (I366698,I366647,I430363);
nor I_21398 (I366490,I366562,I366698);
nor I_21399 (I366729,I430363,I430345);
not I_21400 (I366746,I430354);
nor I_21401 (I366763,I430357,I430342);
nand I_21402 (I366502,I366664,I366763);
not I_21403 (I366794,I430357);
nand I_21404 (I366811,I366794,I366681);
nor I_21405 (I366828,I366746,I430357);
nor I_21406 (I366845,I366828,I430372);
nor I_21407 (I366508,I366613,I366845);
nor I_21408 (I366876,I366828,I366596);
nand I_21409 (I366499,I366630,I366876);
nor I_21410 (I366907,I430345,I430348);
DFFARX1 I_21411 (I366907,I2898,I366528,I366933,);
not I_21412 (I366941,I366933);
not I_21413 (I366958,I430345);
nor I_21414 (I366975,I430345,I430363);
or I_21415 (I366992,I430345,I430363);
nand I_21416 (I366517,I366811,I366992);
nand I_21417 (I367023,I366941,I430342);
nand I_21418 (I367040,I430339,I430339);
nor I_21419 (I367057,I367040,I430342);
nor I_21420 (I366487,I366562,I367057);
nand I_21421 (I367088,I366941,I367040);
not I_21422 (I367105,I367088);
DFFARX1 I_21423 (I367105,I2898,I366528,I366505,);
nand I_21424 (I366520,I367088,I367023);
nor I_21425 (I367150,I367040,I366613);
not I_21426 (I366493,I367150);
nor I_21427 (I366514,I367150,I366975);
nor I_21428 (I367195,I367040,I366958);
nand I_21429 (I367212,I366933,I367195);
nand I_21430 (I367229,I366729,I367212);
DFFARX1 I_21431 (I367229,I2898,I366528,I366496,);
or I_21432 (I367260,I367040,I430342);
nand I_21433 (I366511,I366811,I367260);
not I_21434 (I367327,I2905);
or I_21435 (I367344,I208221,I208203);
nand I_21436 (I367361,I208218,I208227);
not I_21437 (I367378,I367361);
nand I_21438 (I367395,I367378,I367344);
not I_21439 (I367412,I367395);
nor I_21440 (I367429,I208206,I208212);
not I_21441 (I367446,I367429);
nor I_21442 (I367463,I367378,I367446);
not I_21443 (I367480,I208215);
nor I_21444 (I367497,I367446,I208206);
nor I_21445 (I367289,I367361,I367497);
nor I_21446 (I367528,I208206,I208206);
not I_21447 (I367545,I208209);
nor I_21448 (I367562,I208200,I208215);
nand I_21449 (I367301,I367463,I367562);
not I_21450 (I367593,I208200);
nand I_21451 (I367610,I367593,I367480);
nor I_21452 (I367627,I367545,I208200);
nor I_21453 (I367644,I367627,I208212);
nor I_21454 (I367307,I367412,I367644);
nor I_21455 (I367675,I367627,I367395);
nand I_21456 (I367298,I367429,I367675);
nor I_21457 (I367706,I208200,I208212);
DFFARX1 I_21458 (I367706,I2898,I367327,I367732,);
not I_21459 (I367740,I367732);
not I_21460 (I367757,I208200);
nor I_21461 (I367774,I208200,I208206);
or I_21462 (I367791,I208200,I208206);
nand I_21463 (I367316,I367610,I367791);
nand I_21464 (I367822,I367740,I208209);
nand I_21465 (I367839,I208224,I208203);
nor I_21466 (I367856,I367839,I208209);
nor I_21467 (I367286,I367361,I367856);
nand I_21468 (I367887,I367740,I367839);
not I_21469 (I367904,I367887);
DFFARX1 I_21470 (I367904,I2898,I367327,I367304,);
nand I_21471 (I367319,I367887,I367822);
nor I_21472 (I367949,I367839,I367412);
not I_21473 (I367292,I367949);
nor I_21474 (I367313,I367949,I367774);
nor I_21475 (I367994,I367839,I367757);
nand I_21476 (I368011,I367732,I367994);
nand I_21477 (I368028,I367528,I368011);
DFFARX1 I_21478 (I368028,I2898,I367327,I367295,);
or I_21479 (I368059,I367839,I208209);
nand I_21480 (I367310,I367610,I368059);
not I_21481 (I368126,I2905);
or I_21482 (I368143,I10273,I10252);
nand I_21483 (I368160,I10276,I10270);
not I_21484 (I368177,I368160);
nand I_21485 (I368194,I368177,I368143);
not I_21486 (I368211,I368194);
nor I_21487 (I368228,I10255,I10252);
not I_21488 (I368245,I368228);
nor I_21489 (I368262,I368177,I368245);
not I_21490 (I368279,I10261);
nor I_21491 (I368296,I368245,I10267);
nor I_21492 (I368088,I368160,I368296);
nor I_21493 (I368327,I10267,I10255);
not I_21494 (I368344,I10258);
nor I_21495 (I368361,I10264,I10261);
nand I_21496 (I368100,I368262,I368361);
not I_21497 (I368392,I10264);
nand I_21498 (I368409,I368392,I368279);
nor I_21499 (I368426,I368344,I10264);
nor I_21500 (I368443,I368426,I10252);
nor I_21501 (I368106,I368211,I368443);
nor I_21502 (I368474,I368426,I368194);
nand I_21503 (I368097,I368228,I368474);
nor I_21504 (I368505,I10258,I10279);
DFFARX1 I_21505 (I368505,I2898,I368126,I368531,);
not I_21506 (I368539,I368531);
not I_21507 (I368556,I10258);
nor I_21508 (I368573,I10258,I10267);
or I_21509 (I368590,I10258,I10267);
nand I_21510 (I368115,I368409,I368590);
nand I_21511 (I368621,I368539,I10255);
nand I_21512 (I368638,I10261,I10282);
nor I_21513 (I368655,I368638,I10255);
nor I_21514 (I368085,I368160,I368655);
nand I_21515 (I368686,I368539,I368638);
not I_21516 (I368703,I368686);
DFFARX1 I_21517 (I368703,I2898,I368126,I368103,);
nand I_21518 (I368118,I368686,I368621);
nor I_21519 (I368748,I368638,I368211);
not I_21520 (I368091,I368748);
nor I_21521 (I368112,I368748,I368573);
nor I_21522 (I368793,I368638,I368556);
nand I_21523 (I368810,I368531,I368793);
nand I_21524 (I368827,I368327,I368810);
DFFARX1 I_21525 (I368827,I2898,I368126,I368094,);
or I_21526 (I368858,I368638,I10255);
nand I_21527 (I368109,I368409,I368858);
not I_21528 (I368925,I2905);
or I_21529 (I368942,I440127,I440109);
nand I_21530 (I368959,I440124,I440118);
not I_21531 (I368976,I368959);
nand I_21532 (I368993,I368976,I368942);
not I_21533 (I369010,I368993);
nor I_21534 (I369027,I440103,I440130);
not I_21535 (I369044,I369027);
nor I_21536 (I369061,I368976,I369044);
not I_21537 (I369078,I440100);
nor I_21538 (I369095,I369044,I440121);
nor I_21539 (I368887,I368959,I369095);
nor I_21540 (I369126,I440121,I440103);
not I_21541 (I369143,I440112);
nor I_21542 (I369160,I440115,I440100);
nand I_21543 (I368899,I369061,I369160);
not I_21544 (I369191,I440115);
nand I_21545 (I369208,I369191,I369078);
nor I_21546 (I369225,I369143,I440115);
nor I_21547 (I369242,I369225,I440130);
nor I_21548 (I368905,I369010,I369242);
nor I_21549 (I369273,I369225,I368993);
nand I_21550 (I368896,I369027,I369273);
nor I_21551 (I369304,I440103,I440106);
DFFARX1 I_21552 (I369304,I2898,I368925,I369330,);
not I_21553 (I369338,I369330);
not I_21554 (I369355,I440103);
nor I_21555 (I369372,I440103,I440121);
or I_21556 (I369389,I440103,I440121);
nand I_21557 (I368914,I369208,I369389);
nand I_21558 (I369420,I369338,I440100);
nand I_21559 (I369437,I440097,I440097);
nor I_21560 (I369454,I369437,I440100);
nor I_21561 (I368884,I368959,I369454);
nand I_21562 (I369485,I369338,I369437);
not I_21563 (I369502,I369485);
DFFARX1 I_21564 (I369502,I2898,I368925,I368902,);
nand I_21565 (I368917,I369485,I369420);
nor I_21566 (I369547,I369437,I369010);
not I_21567 (I368890,I369547);
nor I_21568 (I368911,I369547,I369372);
nor I_21569 (I369592,I369437,I369355);
nand I_21570 (I369609,I369330,I369592);
nand I_21571 (I369626,I369126,I369609);
DFFARX1 I_21572 (I369626,I2898,I368925,I368893,);
or I_21573 (I369657,I369437,I440100);
nand I_21574 (I368908,I369208,I369657);
not I_21575 (I369724,I2905);
or I_21576 (I369741,I299575,I299578);
nand I_21577 (I369758,I299605,I299587);
not I_21578 (I369775,I369758);
nand I_21579 (I369792,I369775,I369741);
not I_21580 (I369809,I369792);
nor I_21581 (I369826,I299578,I299602);
not I_21582 (I369843,I369826);
nor I_21583 (I369860,I369775,I369843);
not I_21584 (I369877,I299584);
nor I_21585 (I369894,I369843,I299596);
nor I_21586 (I369686,I369758,I369894);
nor I_21587 (I369925,I299596,I299578);
not I_21588 (I369942,I299599);
nor I_21589 (I369959,I299575,I299584);
nand I_21590 (I369698,I369860,I369959);
not I_21591 (I369990,I299575);
nand I_21592 (I370007,I369990,I369877);
nor I_21593 (I370024,I369942,I299575);
nor I_21594 (I370041,I370024,I299602);
nor I_21595 (I369704,I369809,I370041);
nor I_21596 (I370072,I370024,I369792);
nand I_21597 (I369695,I369826,I370072);
nor I_21598 (I370103,I299581,I299581);
DFFARX1 I_21599 (I370103,I2898,I369724,I370129,);
not I_21600 (I370137,I370129);
not I_21601 (I370154,I299581);
nor I_21602 (I370171,I299581,I299596);
or I_21603 (I370188,I299581,I299596);
nand I_21604 (I369713,I370007,I370188);
nand I_21605 (I370219,I370137,I299584);
nand I_21606 (I370236,I299593,I299590);
nor I_21607 (I370253,I370236,I299584);
nor I_21608 (I369683,I369758,I370253);
nand I_21609 (I370284,I370137,I370236);
not I_21610 (I370301,I370284);
DFFARX1 I_21611 (I370301,I2898,I369724,I369701,);
nand I_21612 (I369716,I370284,I370219);
nor I_21613 (I370346,I370236,I369809);
not I_21614 (I369689,I370346);
nor I_21615 (I369710,I370346,I370171);
nor I_21616 (I370391,I370236,I370154);
nand I_21617 (I370408,I370129,I370391);
nand I_21618 (I370425,I369925,I370408);
DFFARX1 I_21619 (I370425,I2898,I369724,I369692,);
or I_21620 (I370456,I370236,I299584);
nand I_21621 (I369707,I370007,I370456);
not I_21622 (I370523,I2905);
or I_21623 (I370540,I99055,I99046);
nand I_21624 (I370557,I99043,I99052);
not I_21625 (I370574,I370557);
nand I_21626 (I370591,I370574,I370540);
not I_21627 (I370608,I370591);
nor I_21628 (I370625,I99049,I99067);
not I_21629 (I370642,I370625);
nor I_21630 (I370659,I370574,I370642);
not I_21631 (I370676,I99049);
nor I_21632 (I370693,I370642,I99058);
nor I_21633 (I370485,I370557,I370693);
nor I_21634 (I370724,I99058,I99049);
not I_21635 (I370741,I99058);
nor I_21636 (I370758,I99055,I99049);
nand I_21637 (I370497,I370659,I370758);
not I_21638 (I370789,I99055);
nand I_21639 (I370806,I370789,I370676);
nor I_21640 (I370823,I370741,I99055);
nor I_21641 (I370840,I370823,I99067);
nor I_21642 (I370503,I370608,I370840);
nor I_21643 (I370871,I370823,I370591);
nand I_21644 (I370494,I370625,I370871);
nor I_21645 (I370902,I99064,I99052);
DFFARX1 I_21646 (I370902,I2898,I370523,I370928,);
not I_21647 (I370936,I370928);
not I_21648 (I370953,I99064);
nor I_21649 (I370970,I99064,I99058);
or I_21650 (I370987,I99064,I99058);
nand I_21651 (I370512,I370806,I370987);
nand I_21652 (I371018,I370936,I99061);
nand I_21653 (I371035,I99046,I99043);
nor I_21654 (I371052,I371035,I99061);
nor I_21655 (I370482,I370557,I371052);
nand I_21656 (I371083,I370936,I371035);
not I_21657 (I371100,I371083);
DFFARX1 I_21658 (I371100,I2898,I370523,I370500,);
nand I_21659 (I370515,I371083,I371018);
nor I_21660 (I371145,I371035,I370608);
not I_21661 (I370488,I371145);
nor I_21662 (I370509,I371145,I370970);
nor I_21663 (I371190,I371035,I370953);
nand I_21664 (I371207,I370928,I371190);
nand I_21665 (I371224,I370724,I371207);
DFFARX1 I_21666 (I371224,I2898,I370523,I370491,);
or I_21667 (I371255,I371035,I99061);
nand I_21668 (I370506,I370806,I371255);
not I_21669 (I371322,I2905);
or I_21670 (I371339,I258198,I258195);
nand I_21671 (I371356,I258180,I258180);
not I_21672 (I371373,I371356);
nand I_21673 (I371390,I371373,I371339);
not I_21674 (I371407,I371390);
nand I_21675 (I371424,I258189,I258207);
and I_21676 (I371441,I371424,I258183);
DFFARX1 I_21677 (I371441,I2898,I371322,I371467,);
nor I_21678 (I371475,I258183,I258207);
not I_21679 (I371492,I371475);
nor I_21680 (I371509,I371467,I371475);
DFFARX1 I_21681 (I371509,I2898,I371322,I371293,);
or I_21682 (I371540,I258186,I258201);
nor I_21683 (I371557,I371540,I258189);
not I_21684 (I371574,I371557);
nor I_21685 (I371281,I371467,I371574);
nand I_21686 (I371305,I371356,I371574);
nor I_21687 (I371619,I258186,I258210);
not I_21688 (I371636,I258204);
nor I_21689 (I371653,I371636,I258192);
not I_21690 (I371670,I371653);
nor I_21691 (I371687,I371670,I371390);
nor I_21692 (I371287,I371492,I371687);
nand I_21693 (I371718,I371670,I371492);
nand I_21694 (I371735,I371407,I371718);
nor I_21695 (I371290,I371574,I371735);
nand I_21696 (I371299,I371356,I371670);
nor I_21697 (I371308,I371467,I371653);
nor I_21698 (I371296,I371653,I371407);
nor I_21699 (I371808,I371619,I371636);
nor I_21700 (I371825,I371373,I371808);
nor I_21701 (I371284,I371574,I371825);
nor I_21702 (I371856,I371467,I371808);
nor I_21703 (I371314,I371653,I371856);
nor I_21704 (I371311,I371856,I371492);
and I_21705 (I371901,I371390,I371808);
nor I_21706 (I371302,I371557,I371901);
not I_21707 (I371968,I2905);
or I_21708 (I371985,I194612,I194603);
nand I_21709 (I372002,I194609,I194615);
not I_21710 (I372019,I372002);
nand I_21711 (I372036,I372019,I371985);
not I_21712 (I372053,I372036);
nand I_21713 (I372070,I194606,I194612);
and I_21714 (I372087,I372070,I194621);
DFFARX1 I_21715 (I372087,I2898,I371968,I372113,);
nor I_21716 (I372121,I194600,I194612);
not I_21717 (I372138,I372121);
nor I_21718 (I372155,I372113,I372121);
DFFARX1 I_21719 (I372155,I2898,I371968,I371939,);
or I_21720 (I372186,I194606,I194609);
nor I_21721 (I372203,I372186,I194618);
not I_21722 (I372220,I372203);
nor I_21723 (I371927,I372113,I372220);
nand I_21724 (I371951,I372002,I372220);
nor I_21725 (I372265,I194615,I194603);
not I_21726 (I372282,I194624);
nor I_21727 (I372299,I372282,I194600);
not I_21728 (I372316,I372299);
nor I_21729 (I372333,I372316,I372036);
nor I_21730 (I371933,I372138,I372333);
nand I_21731 (I372364,I372316,I372138);
nand I_21732 (I372381,I372053,I372364);
nor I_21733 (I371936,I372220,I372381);
nand I_21734 (I371945,I372002,I372316);
nor I_21735 (I371954,I372113,I372299);
nor I_21736 (I371942,I372299,I372053);
nor I_21737 (I372454,I372265,I372282);
nor I_21738 (I372471,I372019,I372454);
nor I_21739 (I371930,I372220,I372471);
nor I_21740 (I372502,I372113,I372454);
nor I_21741 (I371960,I372299,I372502);
nor I_21742 (I371957,I372502,I372138);
and I_21743 (I372547,I372036,I372454);
nor I_21744 (I371948,I372203,I372547);
not I_21745 (I372614,I2905);
or I_21746 (I372631,I340089,I340089);
nand I_21747 (I372648,I340095,I340107);
not I_21748 (I372665,I372648);
nand I_21749 (I372682,I372665,I372631);
not I_21750 (I372699,I372682);
nand I_21751 (I372716,I340095,I340098);
and I_21752 (I372733,I372716,I340101);
DFFARX1 I_21753 (I372733,I2898,I372614,I372759,);
nor I_21754 (I372767,I340086,I340098);
not I_21755 (I372784,I372767);
nor I_21756 (I372801,I372759,I372767);
DFFARX1 I_21757 (I372801,I2898,I372614,I372585,);
or I_21758 (I372832,I340104,I340092);
nor I_21759 (I372849,I372832,I340086);
not I_21760 (I372866,I372849);
nor I_21761 (I372573,I372759,I372866);
nand I_21762 (I372597,I372648,I372866);
nor I_21763 (I372911,I340101,I340092);
not I_21764 (I372928,I340110);
nor I_21765 (I372945,I372928,I340098);
not I_21766 (I372962,I372945);
nor I_21767 (I372979,I372962,I372682);
nor I_21768 (I372579,I372784,I372979);
nand I_21769 (I373010,I372962,I372784);
nand I_21770 (I373027,I372699,I373010);
nor I_21771 (I372582,I372866,I373027);
nand I_21772 (I372591,I372648,I372962);
nor I_21773 (I372600,I372759,I372945);
nor I_21774 (I372588,I372945,I372699);
nor I_21775 (I373100,I372911,I372928);
nor I_21776 (I373117,I372665,I373100);
nor I_21777 (I372576,I372866,I373117);
nor I_21778 (I373148,I372759,I373100);
nor I_21779 (I372606,I372945,I373148);
nor I_21780 (I372603,I373148,I372784);
and I_21781 (I373193,I372682,I373100);
nor I_21782 (I372594,I372849,I373193);
not I_21783 (I373260,I2905);
or I_21784 (I373277,I58821,I58833);
nand I_21785 (I373294,I58833,I58842);
not I_21786 (I373311,I373294);
nand I_21787 (I373328,I373311,I373277);
not I_21788 (I373345,I373328);
nand I_21789 (I373362,I58830,I58824);
and I_21790 (I373379,I373362,I58848);
DFFARX1 I_21791 (I373379,I2898,I373260,I373405,);
nor I_21792 (I373413,I58824,I58824);
not I_21793 (I373430,I373413);
nor I_21794 (I373447,I373405,I373413);
DFFARX1 I_21795 (I373447,I2898,I373260,I373231,);
or I_21796 (I373478,I58836,I58830);
nor I_21797 (I373495,I373478,I58839);
not I_21798 (I373512,I373495);
nor I_21799 (I373219,I373405,I373512);
nand I_21800 (I373243,I373294,I373512);
nor I_21801 (I373557,I58845,I58827);
not I_21802 (I373574,I58827);
nor I_21803 (I373591,I373574,I58821);
not I_21804 (I373608,I373591);
nor I_21805 (I373625,I373608,I373328);
nor I_21806 (I373225,I373430,I373625);
nand I_21807 (I373656,I373608,I373430);
nand I_21808 (I373673,I373345,I373656);
nor I_21809 (I373228,I373512,I373673);
nand I_21810 (I373237,I373294,I373608);
nor I_21811 (I373246,I373405,I373591);
nor I_21812 (I373234,I373591,I373345);
nor I_21813 (I373746,I373557,I373574);
nor I_21814 (I373763,I373311,I373746);
nor I_21815 (I373222,I373512,I373763);
nor I_21816 (I373794,I373405,I373746);
nor I_21817 (I373252,I373591,I373794);
nor I_21818 (I373249,I373794,I373430);
and I_21819 (I373839,I373328,I373746);
nor I_21820 (I373240,I373495,I373839);
not I_21821 (I373906,I2905);
or I_21822 (I373923,I159280,I159301);
nand I_21823 (I373940,I159286,I159277);
not I_21824 (I373957,I373940);
nand I_21825 (I373974,I373957,I373923);
not I_21826 (I373991,I373974);
nand I_21827 (I374008,I159283,I159289);
and I_21828 (I374025,I374008,I159292);
DFFARX1 I_21829 (I374025,I2898,I373906,I374051,);
nor I_21830 (I374059,I159274,I159289);
not I_21831 (I374076,I374059);
nor I_21832 (I374093,I374051,I374059);
DFFARX1 I_21833 (I374093,I2898,I373906,I373877,);
or I_21834 (I374124,I159304,I159298);
nor I_21835 (I374141,I374124,I159277);
not I_21836 (I374158,I374141);
nor I_21837 (I373865,I374051,I374158);
nand I_21838 (I373889,I373940,I374158);
nor I_21839 (I374203,I159280,I159274);
not I_21840 (I374220,I159295);
nor I_21841 (I374237,I374220,I159307);
not I_21842 (I374254,I374237);
nor I_21843 (I374271,I374254,I373974);
nor I_21844 (I373871,I374076,I374271);
nand I_21845 (I374302,I374254,I374076);
nand I_21846 (I374319,I373991,I374302);
nor I_21847 (I373874,I374158,I374319);
nand I_21848 (I373883,I373940,I374254);
nor I_21849 (I373892,I374051,I374237);
nor I_21850 (I373880,I374237,I373991);
nor I_21851 (I374392,I374203,I374220);
nor I_21852 (I374409,I373957,I374392);
nor I_21853 (I373868,I374158,I374409);
nor I_21854 (I374440,I374051,I374392);
nor I_21855 (I373898,I374237,I374440);
nor I_21856 (I373895,I374440,I374076);
and I_21857 (I374485,I373974,I374392);
nor I_21858 (I373886,I374141,I374485);
not I_21859 (I374552,I2905);
or I_21860 (I374569,I95303,I95315);
nand I_21861 (I374586,I95315,I95324);
not I_21862 (I374603,I374586);
nand I_21863 (I374620,I374603,I374569);
not I_21864 (I374637,I374620);
nand I_21865 (I374654,I95312,I95306);
and I_21866 (I374671,I374654,I95330);
DFFARX1 I_21867 (I374671,I2898,I374552,I374697,);
nor I_21868 (I374705,I95306,I95306);
not I_21869 (I374722,I374705);
nor I_21870 (I374739,I374697,I374705);
DFFARX1 I_21871 (I374739,I2898,I374552,I374523,);
or I_21872 (I374770,I95318,I95312);
nor I_21873 (I374787,I374770,I95321);
not I_21874 (I374804,I374787);
nor I_21875 (I374511,I374697,I374804);
nand I_21876 (I374535,I374586,I374804);
nor I_21877 (I374849,I95327,I95309);
not I_21878 (I374866,I95309);
nor I_21879 (I374883,I374866,I95303);
not I_21880 (I374900,I374883);
nor I_21881 (I374917,I374900,I374620);
nor I_21882 (I374517,I374722,I374917);
nand I_21883 (I374948,I374900,I374722);
nand I_21884 (I374965,I374637,I374948);
nor I_21885 (I374520,I374804,I374965);
nand I_21886 (I374529,I374586,I374900);
nor I_21887 (I374538,I374697,I374883);
nor I_21888 (I374526,I374883,I374637);
nor I_21889 (I375038,I374849,I374866);
nor I_21890 (I375055,I374603,I375038);
nor I_21891 (I374514,I374804,I375055);
nor I_21892 (I375086,I374697,I375038);
nor I_21893 (I374544,I374883,I375086);
nor I_21894 (I374541,I375086,I374722);
and I_21895 (I375131,I374620,I375038);
nor I_21896 (I374532,I374787,I375131);
not I_21897 (I375198,I2905);
or I_21898 (I375215,I251313,I251310);
nand I_21899 (I375232,I251295,I251295);
not I_21900 (I375249,I375232);
nand I_21901 (I375266,I375249,I375215);
not I_21902 (I375283,I375266);
nand I_21903 (I375300,I251304,I251322);
and I_21904 (I375317,I375300,I251298);
DFFARX1 I_21905 (I375317,I2898,I375198,I375343,);
nor I_21906 (I375351,I251298,I251322);
not I_21907 (I375368,I375351);
nor I_21908 (I375385,I375343,I375351);
DFFARX1 I_21909 (I375385,I2898,I375198,I375169,);
or I_21910 (I375416,I251301,I251316);
nor I_21911 (I375433,I375416,I251304);
not I_21912 (I375450,I375433);
nor I_21913 (I375157,I375343,I375450);
nand I_21914 (I375181,I375232,I375450);
nor I_21915 (I375495,I251301,I251325);
not I_21916 (I375512,I251319);
nor I_21917 (I375529,I375512,I251307);
not I_21918 (I375546,I375529);
nor I_21919 (I375563,I375546,I375266);
nor I_21920 (I375163,I375368,I375563);
nand I_21921 (I375594,I375546,I375368);
nand I_21922 (I375611,I375283,I375594);
nor I_21923 (I375166,I375450,I375611);
nand I_21924 (I375175,I375232,I375546);
nor I_21925 (I375184,I375343,I375529);
nor I_21926 (I375172,I375529,I375283);
nor I_21927 (I375684,I375495,I375512);
nor I_21928 (I375701,I375249,I375684);
nor I_21929 (I375160,I375450,I375701);
nor I_21930 (I375732,I375343,I375684);
nor I_21931 (I375190,I375529,I375732);
nor I_21932 (I375187,I375732,I375368);
and I_21933 (I375777,I375266,I375684);
nor I_21934 (I375178,I375433,I375777);
not I_21935 (I375844,I2905);
or I_21936 (I375861,I8422,I8437);
nand I_21937 (I375878,I8443,I8440);
not I_21938 (I375895,I375878);
nand I_21939 (I375912,I375895,I375861);
not I_21940 (I375929,I375912);
nand I_21941 (I375946,I8416,I8419);
and I_21942 (I375963,I375946,I8428);
DFFARX1 I_21943 (I375963,I2898,I375844,I375989,);
nor I_21944 (I375997,I8425,I8419);
not I_21945 (I376014,I375997);
nor I_21946 (I376031,I375989,I375997);
DFFARX1 I_21947 (I376031,I2898,I375844,I375815,);
or I_21948 (I376062,I8419,I8422);
nor I_21949 (I376079,I376062,I8425);
not I_21950 (I376096,I376079);
nor I_21951 (I375803,I375989,I376096);
nand I_21952 (I375827,I375878,I376096);
nor I_21953 (I376141,I8431,I8416);
not I_21954 (I376158,I8434);
nor I_21955 (I376175,I376158,I8446);
not I_21956 (I376192,I376175);
nor I_21957 (I376209,I376192,I375912);
nor I_21958 (I375809,I376014,I376209);
nand I_21959 (I376240,I376192,I376014);
nand I_21960 (I376257,I375929,I376240);
nor I_21961 (I375812,I376096,I376257);
nand I_21962 (I375821,I375878,I376192);
nor I_21963 (I375830,I375989,I376175);
nor I_21964 (I375818,I376175,I375929);
nor I_21965 (I376330,I376141,I376158);
nor I_21966 (I376347,I375895,I376330);
nor I_21967 (I375806,I376096,I376347);
nor I_21968 (I376378,I375989,I376330);
nor I_21969 (I375836,I376175,I376378);
nor I_21970 (I375833,I376378,I376014);
and I_21971 (I376423,I375912,I376330);
nor I_21972 (I375824,I376079,I376423);
not I_21973 (I376490,I2905);
or I_21974 (I376507,I153840,I153861);
nand I_21975 (I376524,I153846,I153837);
not I_21976 (I376541,I376524);
nand I_21977 (I376558,I376541,I376507);
not I_21978 (I376575,I376558);
nand I_21979 (I376592,I153843,I153849);
and I_21980 (I376609,I376592,I153852);
DFFARX1 I_21981 (I376609,I2898,I376490,I376635,);
nor I_21982 (I376643,I153834,I153849);
not I_21983 (I376660,I376643);
nor I_21984 (I376677,I376635,I376643);
DFFARX1 I_21985 (I376677,I2898,I376490,I376461,);
or I_21986 (I376708,I153864,I153858);
nor I_21987 (I376725,I376708,I153837);
not I_21988 (I376742,I376725);
nor I_21989 (I376449,I376635,I376742);
nand I_21990 (I376473,I376524,I376742);
nor I_21991 (I376787,I153840,I153834);
not I_21992 (I376804,I153855);
nor I_21993 (I376821,I376804,I153867);
not I_21994 (I376838,I376821);
nor I_21995 (I376855,I376838,I376558);
nor I_21996 (I376455,I376660,I376855);
nand I_21997 (I376886,I376838,I376660);
nand I_21998 (I376903,I376575,I376886);
nor I_21999 (I376458,I376742,I376903);
nand I_22000 (I376467,I376524,I376838);
nor I_22001 (I376476,I376635,I376821);
nor I_22002 (I376464,I376821,I376575);
nor I_22003 (I376976,I376787,I376804);
nor I_22004 (I376993,I376541,I376976);
nor I_22005 (I376452,I376742,I376993);
nor I_22006 (I377024,I376635,I376976);
nor I_22007 (I376482,I376821,I377024);
nor I_22008 (I376479,I377024,I376660);
and I_22009 (I377069,I376558,I376976);
nor I_22010 (I376470,I376725,I377069);
not I_22011 (I377136,I2905);
or I_22012 (I377153,I295195,I295207);
nand I_22013 (I377170,I295195,I295210);
not I_22014 (I377187,I377170);
nand I_22015 (I377204,I377187,I377153);
not I_22016 (I377221,I377204);
nand I_22017 (I377238,I295213,I295189);
and I_22018 (I377255,I377238,I295192);
DFFARX1 I_22019 (I377255,I2898,I377136,I377281,);
nor I_22020 (I377289,I295216,I295189);
not I_22021 (I377306,I377289);
nor I_22022 (I377323,I377281,I377289);
DFFARX1 I_22023 (I377323,I2898,I377136,I377107,);
or I_22024 (I377354,I295198,I295189);
nor I_22025 (I377371,I377354,I295219);
not I_22026 (I377388,I377371);
nor I_22027 (I377095,I377281,I377388);
nand I_22028 (I377119,I377170,I377388);
nor I_22029 (I377433,I295204,I295192);
not I_22030 (I377450,I295201);
nor I_22031 (I377467,I377450,I295198);
not I_22032 (I377484,I377467);
nor I_22033 (I377501,I377484,I377204);
nor I_22034 (I377101,I377306,I377501);
nand I_22035 (I377532,I377484,I377306);
nand I_22036 (I377549,I377221,I377532);
nor I_22037 (I377104,I377388,I377549);
nand I_22038 (I377113,I377170,I377484);
nor I_22039 (I377122,I377281,I377467);
nor I_22040 (I377110,I377467,I377221);
nor I_22041 (I377622,I377433,I377450);
nor I_22042 (I377639,I377187,I377622);
nor I_22043 (I377098,I377388,I377639);
nor I_22044 (I377670,I377281,I377622);
nor I_22045 (I377128,I377467,I377670);
nor I_22046 (I377125,I377670,I377306);
and I_22047 (I377715,I377204,I377622);
nor I_22048 (I377116,I377371,I377715);
not I_22049 (I377782,I2905);
or I_22050 (I377799,I82094,I82106);
nand I_22051 (I377816,I82106,I82115);
not I_22052 (I377833,I377816);
nand I_22053 (I377850,I377833,I377799);
not I_22054 (I377867,I377850);
nand I_22055 (I377884,I82103,I82097);
and I_22056 (I377901,I377884,I82121);
DFFARX1 I_22057 (I377901,I2898,I377782,I377927,);
nor I_22058 (I377935,I82097,I82097);
not I_22059 (I377952,I377935);
nor I_22060 (I377969,I377927,I377935);
DFFARX1 I_22061 (I377969,I2898,I377782,I377753,);
or I_22062 (I378000,I82109,I82103);
nor I_22063 (I378017,I378000,I82112);
not I_22064 (I378034,I378017);
nor I_22065 (I377741,I377927,I378034);
nand I_22066 (I377765,I377816,I378034);
nor I_22067 (I378079,I82118,I82100);
not I_22068 (I378096,I82100);
nor I_22069 (I378113,I378096,I82094);
not I_22070 (I378130,I378113);
nor I_22071 (I378147,I378130,I377850);
nor I_22072 (I377747,I377952,I378147);
nand I_22073 (I378178,I378130,I377952);
nand I_22074 (I378195,I377867,I378178);
nor I_22075 (I377750,I378034,I378195);
nand I_22076 (I377759,I377816,I378130);
nor I_22077 (I377768,I377927,I378113);
nor I_22078 (I377756,I378113,I377867);
nor I_22079 (I378268,I378079,I378096);
nor I_22080 (I378285,I377833,I378268);
nor I_22081 (I377744,I378034,I378285);
nor I_22082 (I378316,I377927,I378268);
nor I_22083 (I377774,I378113,I378316);
nor I_22084 (I377771,I378316,I377952);
and I_22085 (I378361,I377850,I378268);
nor I_22086 (I377762,I378017,I378361);
not I_22087 (I378428,I2905);
or I_22088 (I378445,I415735,I415708);
nand I_22089 (I378462,I415705,I415723);
not I_22090 (I378479,I378462);
nand I_22091 (I378496,I378479,I378445);
not I_22092 (I378513,I378496);
nand I_22093 (I378530,I415726,I415711);
and I_22094 (I378547,I378530,I415729);
DFFARX1 I_22095 (I378547,I2898,I378428,I378573,);
nor I_22096 (I378581,I415702,I415711);
not I_22097 (I378598,I378581);
nor I_22098 (I378615,I378573,I378581);
DFFARX1 I_22099 (I378615,I2898,I378428,I378399,);
or I_22100 (I378646,I415720,I415705);
nor I_22101 (I378663,I378646,I415717);
not I_22102 (I378680,I378663);
nor I_22103 (I378387,I378573,I378680);
nand I_22104 (I378411,I378462,I378680);
nor I_22105 (I378725,I415702,I415714);
not I_22106 (I378742,I415732);
nor I_22107 (I378759,I378742,I415708);
not I_22108 (I378776,I378759);
nor I_22109 (I378793,I378776,I378496);
nor I_22110 (I378393,I378598,I378793);
nand I_22111 (I378824,I378776,I378598);
nand I_22112 (I378841,I378513,I378824);
nor I_22113 (I378396,I378680,I378841);
nand I_22114 (I378405,I378462,I378776);
nor I_22115 (I378414,I378573,I378759);
nor I_22116 (I378402,I378759,I378513);
nor I_22117 (I378914,I378725,I378742);
nor I_22118 (I378931,I378479,I378914);
nor I_22119 (I378390,I378680,I378931);
nor I_22120 (I378962,I378573,I378914);
nor I_22121 (I378420,I378759,I378962);
nor I_22122 (I378417,I378962,I378598);
and I_22123 (I379007,I378496,I378914);
nor I_22124 (I378408,I378663,I379007);
not I_22125 (I379074,I2905);
or I_22126 (I379091,I99688,I99679);
nand I_22127 (I379108,I99661,I99658);
not I_22128 (I379125,I379108);
nand I_22129 (I379142,I379125,I379091);
not I_22130 (I379159,I379142);
nand I_22131 (I379176,I99658,I99673);
and I_22132 (I379193,I379176,I99655);
DFFARX1 I_22133 (I379193,I2898,I379074,I379219,);
nor I_22134 (I379227,I99661,I99673);
not I_22135 (I379244,I379227);
nor I_22136 (I379261,I379219,I379227);
DFFARX1 I_22137 (I379261,I2898,I379074,I379045,);
or I_22138 (I379292,I99670,I99664);
nor I_22139 (I379309,I379292,I99667);
not I_22140 (I379326,I379309);
nor I_22141 (I379033,I379219,I379326);
nand I_22142 (I379057,I379108,I379326);
nor I_22143 (I379371,I99685,I99676);
not I_22144 (I379388,I99682);
nor I_22145 (I379405,I379388,I99655);
not I_22146 (I379422,I379405);
nor I_22147 (I379439,I379422,I379142);
nor I_22148 (I379039,I379244,I379439);
nand I_22149 (I379470,I379422,I379244);
nand I_22150 (I379487,I379159,I379470);
nor I_22151 (I379042,I379326,I379487);
nand I_22152 (I379051,I379108,I379422);
nor I_22153 (I379060,I379219,I379405);
nor I_22154 (I379048,I379405,I379159);
nor I_22155 (I379560,I379371,I379388);
nor I_22156 (I379577,I379125,I379560);
nor I_22157 (I379036,I379326,I379577);
nor I_22158 (I379608,I379219,I379560);
nor I_22159 (I379066,I379405,I379608);
nor I_22160 (I379063,I379608,I379244);
and I_22161 (I379653,I379142,I379560);
nor I_22162 (I379054,I379309,I379653);
not I_22163 (I379720,I2905);
or I_22164 (I379737,I297388,I297400);
nand I_22165 (I379754,I297388,I297403);
not I_22166 (I379771,I379754);
nand I_22167 (I379788,I379771,I379737);
not I_22168 (I379805,I379788);
nand I_22169 (I379822,I297406,I297382);
and I_22170 (I379839,I379822,I297385);
DFFARX1 I_22171 (I379839,I2898,I379720,I379865,);
nor I_22172 (I379873,I297409,I297382);
not I_22173 (I379890,I379873);
nor I_22174 (I379907,I379865,I379873);
DFFARX1 I_22175 (I379907,I2898,I379720,I379691,);
or I_22176 (I379938,I297391,I297382);
nor I_22177 (I379955,I379938,I297412);
not I_22178 (I379972,I379955);
nor I_22179 (I379679,I379865,I379972);
nand I_22180 (I379703,I379754,I379972);
nor I_22181 (I380017,I297397,I297385);
not I_22182 (I380034,I297394);
nor I_22183 (I380051,I380034,I297391);
not I_22184 (I380068,I380051);
nor I_22185 (I380085,I380068,I379788);
nor I_22186 (I379685,I379890,I380085);
nand I_22187 (I380116,I380068,I379890);
nand I_22188 (I380133,I379805,I380116);
nor I_22189 (I379688,I379972,I380133);
nand I_22190 (I379697,I379754,I380068);
nor I_22191 (I379706,I379865,I380051);
nor I_22192 (I379694,I380051,I379805);
nor I_22193 (I380206,I380017,I380034);
nor I_22194 (I380223,I379771,I380206);
nor I_22195 (I379682,I379972,I380223);
nor I_22196 (I380254,I379865,I380206);
nor I_22197 (I379712,I380051,I380254);
nor I_22198 (I379709,I380254,I379890);
and I_22199 (I380299,I379788,I380206);
nor I_22200 (I379700,I379955,I380299);
not I_22201 (I380366,I2905);
or I_22202 (I380383,I404032,I404029);
nand I_22203 (I380400,I404038,I404041);
not I_22204 (I380417,I380400);
nand I_22205 (I380434,I380417,I380383);
not I_22206 (I380451,I380434);
nand I_22207 (I380468,I404029,I404035);
and I_22208 (I380485,I380468,I404026);
DFFARX1 I_22209 (I380485,I2898,I380366,I380511,);
nor I_22210 (I380519,I404023,I404035);
not I_22211 (I380536,I380519);
nor I_22212 (I380553,I380511,I380519);
DFFARX1 I_22213 (I380553,I2898,I380366,I380337,);
or I_22214 (I380584,I404023,I404032);
nor I_22215 (I380601,I380584,I404026);
not I_22216 (I380618,I380601);
nor I_22217 (I380325,I380511,I380618);
nand I_22218 (I380349,I380400,I380618);
nor I_22219 (I380663,I404038,I404044);
not I_22220 (I380680,I404047);
nor I_22221 (I380697,I380680,I404035);
not I_22222 (I380714,I380697);
nor I_22223 (I380731,I380714,I380434);
nor I_22224 (I380331,I380536,I380731);
nand I_22225 (I380762,I380714,I380536);
nand I_22226 (I380779,I380451,I380762);
nor I_22227 (I380334,I380618,I380779);
nand I_22228 (I380343,I380400,I380714);
nor I_22229 (I380352,I380511,I380697);
nor I_22230 (I380340,I380697,I380451);
nor I_22231 (I380852,I380663,I380680);
nor I_22232 (I380869,I380417,I380852);
nor I_22233 (I380328,I380618,I380869);
nor I_22234 (I380900,I380511,I380852);
nor I_22235 (I380358,I380697,I380900);
nor I_22236 (I380355,I380900,I380536);
and I_22237 (I380945,I380434,I380852);
nor I_22238 (I380346,I380601,I380945);
not I_22239 (I381012,I2905);
or I_22240 (I381029,I212691,I212709);
nand I_22241 (I381046,I212700,I212697);
not I_22242 (I381063,I381046);
nand I_22243 (I381080,I381063,I381029);
not I_22244 (I381097,I381080);
nand I_22245 (I381114,I212697,I212691);
and I_22246 (I381131,I381114,I212694);
DFFARX1 I_22247 (I381131,I2898,I381012,I381157,);
nor I_22248 (I381165,I212712,I212691);
not I_22249 (I381182,I381165);
nor I_22250 (I381199,I381157,I381165);
DFFARX1 I_22251 (I381199,I2898,I381012,I380983,);
or I_22252 (I381230,I212706,I212688);
nor I_22253 (I381247,I381230,I212715);
not I_22254 (I381264,I381247);
nor I_22255 (I380971,I381157,I381264);
nand I_22256 (I380995,I381046,I381264);
nor I_22257 (I381309,I212688,I212694);
not I_22258 (I381326,I212703);
nor I_22259 (I381343,I381326,I212700);
not I_22260 (I381360,I381343);
nor I_22261 (I381377,I381360,I381080);
nor I_22262 (I380977,I381182,I381377);
nand I_22263 (I381408,I381360,I381182);
nand I_22264 (I381425,I381097,I381408);
nor I_22265 (I380980,I381264,I381425);
nand I_22266 (I380989,I381046,I381360);
nor I_22267 (I380998,I381157,I381343);
nor I_22268 (I380986,I381343,I381097);
nor I_22269 (I381498,I381309,I381326);
nor I_22270 (I381515,I381063,I381498);
nor I_22271 (I380974,I381264,I381515);
nor I_22272 (I381546,I381157,I381498);
nor I_22273 (I381004,I381343,I381546);
nor I_22274 (I381001,I381546,I381182);
and I_22275 (I381591,I381080,I381498);
nor I_22276 (I380992,I381247,I381591);
not I_22277 (I381658,I2905);
or I_22278 (I381675,I417129,I417102);
nand I_22279 (I381692,I417099,I417117);
not I_22280 (I381709,I381692);
nand I_22281 (I381726,I381709,I381675);
not I_22282 (I381743,I381726);
nand I_22283 (I381760,I417120,I417105);
and I_22284 (I381777,I381760,I417123);
DFFARX1 I_22285 (I381777,I2898,I381658,I381803,);
nor I_22286 (I381811,I417096,I417105);
not I_22287 (I381828,I381811);
nor I_22288 (I381845,I381803,I381811);
DFFARX1 I_22289 (I381845,I2898,I381658,I381629,);
or I_22290 (I381876,I417114,I417099);
nor I_22291 (I381893,I381876,I417111);
not I_22292 (I381910,I381893);
nor I_22293 (I381617,I381803,I381910);
nand I_22294 (I381641,I381692,I381910);
nor I_22295 (I381955,I417096,I417108);
not I_22296 (I381972,I417126);
nor I_22297 (I381989,I381972,I417102);
not I_22298 (I382006,I381989);
nor I_22299 (I382023,I382006,I381726);
nor I_22300 (I381623,I381828,I382023);
nand I_22301 (I382054,I382006,I381828);
nand I_22302 (I382071,I381743,I382054);
nor I_22303 (I381626,I381910,I382071);
nand I_22304 (I381635,I381692,I382006);
nor I_22305 (I381644,I381803,I381989);
nor I_22306 (I381632,I381989,I381743);
nor I_22307 (I382144,I381955,I381972);
nor I_22308 (I382161,I381709,I382144);
nor I_22309 (I381620,I381910,I382161);
nor I_22310 (I382192,I381803,I382144);
nor I_22311 (I381650,I381989,I382192);
nor I_22312 (I381647,I382192,I381828);
and I_22313 (I382237,I381726,I382144);
nor I_22314 (I381638,I381893,I382237);
not I_22315 (I382304,I2905);
or I_22316 (I382321,I102833,I102824);
nand I_22317 (I382338,I102806,I102803);
not I_22318 (I382355,I382338);
nand I_22319 (I382372,I382355,I382321);
not I_22320 (I382389,I382372);
nand I_22321 (I382406,I102803,I102818);
and I_22322 (I382423,I382406,I102800);
DFFARX1 I_22323 (I382423,I2898,I382304,I382449,);
nor I_22324 (I382457,I102806,I102818);
not I_22325 (I382474,I382457);
nor I_22326 (I382491,I382449,I382457);
DFFARX1 I_22327 (I382491,I2898,I382304,I382275,);
or I_22328 (I382522,I102815,I102809);
nor I_22329 (I382539,I382522,I102812);
not I_22330 (I382556,I382539);
nor I_22331 (I382263,I382449,I382556);
nand I_22332 (I382287,I382338,I382556);
nor I_22333 (I382601,I102830,I102821);
not I_22334 (I382618,I102827);
nor I_22335 (I382635,I382618,I102800);
not I_22336 (I382652,I382635);
nor I_22337 (I382669,I382652,I382372);
nor I_22338 (I382269,I382474,I382669);
nand I_22339 (I382700,I382652,I382474);
nand I_22340 (I382717,I382389,I382700);
nor I_22341 (I382272,I382556,I382717);
nand I_22342 (I382281,I382338,I382652);
nor I_22343 (I382290,I382449,I382635);
nor I_22344 (I382278,I382635,I382389);
nor I_22345 (I382790,I382601,I382618);
nor I_22346 (I382807,I382355,I382790);
nor I_22347 (I382266,I382556,I382807);
nor I_22348 (I382838,I382449,I382790);
nor I_22349 (I382296,I382635,I382838);
nor I_22350 (I382293,I382838,I382474);
and I_22351 (I382883,I382372,I382790);
nor I_22352 (I382284,I382539,I382883);
not I_22353 (I382950,I2905);
or I_22354 (I382967,I335924,I335924);
nand I_22355 (I382984,I335930,I335942);
not I_22356 (I383001,I382984);
nand I_22357 (I383018,I383001,I382967);
not I_22358 (I383035,I383018);
nand I_22359 (I383052,I335930,I335933);
and I_22360 (I383069,I383052,I335936);
DFFARX1 I_22361 (I383069,I2898,I382950,I383095,);
nor I_22362 (I383103,I335921,I335933);
not I_22363 (I383120,I383103);
nor I_22364 (I383137,I383095,I383103);
DFFARX1 I_22365 (I383137,I2898,I382950,I382921,);
or I_22366 (I383168,I335939,I335927);
nor I_22367 (I383185,I383168,I335921);
not I_22368 (I383202,I383185);
nor I_22369 (I382909,I383095,I383202);
nand I_22370 (I382933,I382984,I383202);
nor I_22371 (I383247,I335936,I335927);
not I_22372 (I383264,I335945);
nor I_22373 (I383281,I383264,I335933);
not I_22374 (I383298,I383281);
nor I_22375 (I383315,I383298,I383018);
nor I_22376 (I382915,I383120,I383315);
nand I_22377 (I383346,I383298,I383120);
nand I_22378 (I383363,I383035,I383346);
nor I_22379 (I382918,I383202,I383363);
nand I_22380 (I382927,I382984,I383298);
nor I_22381 (I382936,I383095,I383281);
nor I_22382 (I382924,I383281,I383035);
nor I_22383 (I383436,I383247,I383264);
nor I_22384 (I383453,I383001,I383436);
nor I_22385 (I382912,I383202,I383453);
nor I_22386 (I383484,I383095,I383436);
nor I_22387 (I382942,I383281,I383484);
nor I_22388 (I382939,I383484,I383120);
and I_22389 (I383529,I383018,I383436);
nor I_22390 (I382930,I383185,I383529);
not I_22391 (I383596,I2905);
or I_22392 (I383613,I263553,I263550);
nand I_22393 (I383630,I263535,I263535);
not I_22394 (I383647,I383630);
nand I_22395 (I383664,I383647,I383613);
not I_22396 (I383681,I383664);
nand I_22397 (I383698,I263544,I263562);
and I_22398 (I383715,I383698,I263538);
DFFARX1 I_22399 (I383715,I2898,I383596,I383741,);
nor I_22400 (I383749,I263538,I263562);
not I_22401 (I383766,I383749);
nor I_22402 (I383783,I383741,I383749);
DFFARX1 I_22403 (I383783,I2898,I383596,I383567,);
or I_22404 (I383814,I263541,I263556);
nor I_22405 (I383831,I383814,I263544);
not I_22406 (I383848,I383831);
nor I_22407 (I383555,I383741,I383848);
nand I_22408 (I383579,I383630,I383848);
nor I_22409 (I383893,I263541,I263565);
not I_22410 (I383910,I263559);
nor I_22411 (I383927,I383910,I263547);
not I_22412 (I383944,I383927);
nor I_22413 (I383961,I383944,I383664);
nor I_22414 (I383561,I383766,I383961);
nand I_22415 (I383992,I383944,I383766);
nand I_22416 (I384009,I383681,I383992);
nor I_22417 (I383564,I383848,I384009);
nand I_22418 (I383573,I383630,I383944);
nor I_22419 (I383582,I383741,I383927);
nor I_22420 (I383570,I383927,I383681);
nor I_22421 (I384082,I383893,I383910);
nor I_22422 (I384099,I383647,I384082);
nor I_22423 (I383558,I383848,I384099);
nor I_22424 (I384130,I383741,I384082);
nor I_22425 (I383588,I383927,I384130);
nor I_22426 (I383585,I384130,I383766);
and I_22427 (I384175,I383664,I384082);
nor I_22428 (I383576,I383831,I384175);
not I_22429 (I384242,I2905);
or I_22430 (I384259,I92158,I92170);
nand I_22431 (I384276,I92170,I92179);
not I_22432 (I384293,I384276);
nand I_22433 (I384310,I384293,I384259);
not I_22434 (I384327,I384310);
nand I_22435 (I384344,I92167,I92161);
and I_22436 (I384361,I384344,I92185);
DFFARX1 I_22437 (I384361,I2898,I384242,I384387,);
nor I_22438 (I384395,I92161,I92161);
not I_22439 (I384412,I384395);
nor I_22440 (I384429,I384387,I384395);
DFFARX1 I_22441 (I384429,I2898,I384242,I384213,);
or I_22442 (I384460,I92173,I92167);
nor I_22443 (I384477,I384460,I92176);
not I_22444 (I384494,I384477);
nor I_22445 (I384201,I384387,I384494);
nand I_22446 (I384225,I384276,I384494);
nor I_22447 (I384539,I92182,I92164);
not I_22448 (I384556,I92164);
nor I_22449 (I384573,I384556,I92158);
not I_22450 (I384590,I384573);
nor I_22451 (I384607,I384590,I384310);
nor I_22452 (I384207,I384412,I384607);
nand I_22453 (I384638,I384590,I384412);
nand I_22454 (I384655,I384327,I384638);
nor I_22455 (I384210,I384494,I384655);
nand I_22456 (I384219,I384276,I384590);
nor I_22457 (I384228,I384387,I384573);
nor I_22458 (I384216,I384573,I384327);
nor I_22459 (I384728,I384539,I384556);
nor I_22460 (I384745,I384293,I384728);
nor I_22461 (I384204,I384494,I384745);
nor I_22462 (I384776,I384387,I384728);
nor I_22463 (I384234,I384573,I384776);
nor I_22464 (I384231,I384776,I384412);
and I_22465 (I384821,I384310,I384728);
nor I_22466 (I384222,I384477,I384821);
not I_22467 (I384888,I2905);
or I_22468 (I384905,I327594,I327594);
nand I_22469 (I384922,I327600,I327612);
not I_22470 (I384939,I384922);
nand I_22471 (I384956,I384939,I384905);
not I_22472 (I384973,I384956);
nand I_22473 (I384990,I327600,I327603);
and I_22474 (I385007,I384990,I327606);
DFFARX1 I_22475 (I385007,I2898,I384888,I385033,);
nor I_22476 (I385041,I327591,I327603);
not I_22477 (I385058,I385041);
nor I_22478 (I385075,I385033,I385041);
DFFARX1 I_22479 (I385075,I2898,I384888,I384859,);
or I_22480 (I385106,I327609,I327597);
nor I_22481 (I385123,I385106,I327591);
not I_22482 (I385140,I385123);
nor I_22483 (I384847,I385033,I385140);
nand I_22484 (I384871,I384922,I385140);
nor I_22485 (I385185,I327606,I327597);
not I_22486 (I385202,I327615);
nor I_22487 (I385219,I385202,I327603);
not I_22488 (I385236,I385219);
nor I_22489 (I385253,I385236,I384956);
nor I_22490 (I384853,I385058,I385253);
nand I_22491 (I385284,I385236,I385058);
nand I_22492 (I385301,I384973,I385284);
nor I_22493 (I384856,I385140,I385301);
nand I_22494 (I384865,I384922,I385236);
nor I_22495 (I384874,I385033,I385219);
nor I_22496 (I384862,I385219,I384973);
nor I_22497 (I385374,I385185,I385202);
nor I_22498 (I385391,I384939,I385374);
nor I_22499 (I384850,I385140,I385391);
nor I_22500 (I385422,I385033,I385374);
nor I_22501 (I384880,I385219,I385422);
nor I_22502 (I384877,I385422,I385058);
and I_22503 (I385467,I384956,I385374);
nor I_22504 (I384868,I385123,I385467);
not I_22505 (I385534,I2905);
or I_22506 (I385551,I427584,I427557);
nand I_22507 (I385568,I427554,I427572);
not I_22508 (I385585,I385568);
nand I_22509 (I385602,I385585,I385551);
not I_22510 (I385619,I385602);
nand I_22511 (I385636,I427575,I427560);
and I_22512 (I385653,I385636,I427578);
DFFARX1 I_22513 (I385653,I2898,I385534,I385679,);
nor I_22514 (I385687,I427551,I427560);
not I_22515 (I385704,I385687);
nor I_22516 (I385721,I385679,I385687);
DFFARX1 I_22517 (I385721,I2898,I385534,I385505,);
or I_22518 (I385752,I427569,I427554);
nor I_22519 (I385769,I385752,I427566);
not I_22520 (I385786,I385769);
nor I_22521 (I385493,I385679,I385786);
nand I_22522 (I385517,I385568,I385786);
nor I_22523 (I385831,I427551,I427563);
not I_22524 (I385848,I427581);
nor I_22525 (I385865,I385848,I427557);
not I_22526 (I385882,I385865);
nor I_22527 (I385899,I385882,I385602);
nor I_22528 (I385499,I385704,I385899);
nand I_22529 (I385930,I385882,I385704);
nand I_22530 (I385947,I385619,I385930);
nor I_22531 (I385502,I385786,I385947);
nand I_22532 (I385511,I385568,I385882);
nor I_22533 (I385520,I385679,I385865);
nor I_22534 (I385508,I385865,I385619);
nor I_22535 (I386020,I385831,I385848);
nor I_22536 (I386037,I385585,I386020);
nor I_22537 (I385496,I385786,I386037);
nor I_22538 (I386068,I385679,I386020);
nor I_22539 (I385526,I385865,I386068);
nor I_22540 (I385523,I386068,I385704);
and I_22541 (I386113,I385602,I386020);
nor I_22542 (I385514,I385769,I386113);
not I_22543 (I386180,I2905);
or I_22544 (I386197,I217927,I217945);
nand I_22545 (I386214,I217936,I217933);
not I_22546 (I386231,I386214);
nand I_22547 (I386248,I386231,I386197);
not I_22548 (I386265,I386248);
nand I_22549 (I386282,I217933,I217927);
and I_22550 (I386299,I386282,I217930);
DFFARX1 I_22551 (I386299,I2898,I386180,I386325,);
nor I_22552 (I386333,I217948,I217927);
not I_22553 (I386350,I386333);
nor I_22554 (I386367,I386325,I386333);
DFFARX1 I_22555 (I386367,I2898,I386180,I386151,);
or I_22556 (I386398,I217942,I217924);
nor I_22557 (I386415,I386398,I217951);
not I_22558 (I386432,I386415);
nor I_22559 (I386139,I386325,I386432);
nand I_22560 (I386163,I386214,I386432);
nor I_22561 (I386477,I217924,I217930);
not I_22562 (I386494,I217939);
nor I_22563 (I386511,I386494,I217936);
not I_22564 (I386528,I386511);
nor I_22565 (I386545,I386528,I386248);
nor I_22566 (I386145,I386350,I386545);
nand I_22567 (I386576,I386528,I386350);
nand I_22568 (I386593,I386265,I386576);
nor I_22569 (I386148,I386432,I386593);
nand I_22570 (I386157,I386214,I386528);
nor I_22571 (I386166,I386325,I386511);
nor I_22572 (I386154,I386511,I386265);
nor I_22573 (I386666,I386477,I386494);
nor I_22574 (I386683,I386231,I386666);
nor I_22575 (I386142,I386432,I386683);
nor I_22576 (I386714,I386325,I386666);
nor I_22577 (I386172,I386511,I386714);
nor I_22578 (I386169,I386714,I386350);
and I_22579 (I386759,I386248,I386666);
nor I_22580 (I386160,I386415,I386759);
not I_22581 (I386826,I2905);
or I_22582 (I386843,I257433,I257430);
nand I_22583 (I386860,I257415,I257415);
not I_22584 (I386877,I386860);
nand I_22585 (I386894,I386877,I386843);
not I_22586 (I386911,I386894);
nand I_22587 (I386928,I257424,I257442);
and I_22588 (I386945,I386928,I257418);
DFFARX1 I_22589 (I386945,I2898,I386826,I386971,);
nor I_22590 (I386979,I257418,I257442);
not I_22591 (I386996,I386979);
nor I_22592 (I387013,I386971,I386979);
DFFARX1 I_22593 (I387013,I2898,I386826,I386797,);
or I_22594 (I387044,I257421,I257436);
nor I_22595 (I387061,I387044,I257424);
not I_22596 (I387078,I387061);
nor I_22597 (I386785,I386971,I387078);
nand I_22598 (I386809,I386860,I387078);
nor I_22599 (I387123,I257421,I257445);
not I_22600 (I387140,I257439);
nor I_22601 (I387157,I387140,I257427);
not I_22602 (I387174,I387157);
nor I_22603 (I387191,I387174,I386894);
nor I_22604 (I386791,I386996,I387191);
nand I_22605 (I387222,I387174,I386996);
nand I_22606 (I387239,I386911,I387222);
nor I_22607 (I386794,I387078,I387239);
nand I_22608 (I386803,I386860,I387174);
nor I_22609 (I386812,I386971,I387157);
nor I_22610 (I386800,I387157,I386911);
nor I_22611 (I387312,I387123,I387140);
nor I_22612 (I387329,I386877,I387312);
nor I_22613 (I386788,I387078,I387329);
nor I_22614 (I387360,I386971,I387312);
nor I_22615 (I386818,I387157,I387360);
nor I_22616 (I386815,I387360,I386996);
and I_22617 (I387405,I386894,I387312);
nor I_22618 (I386806,I387061,I387405);
not I_22619 (I387472,I2905);
or I_22620 (I387489,I270438,I270435);
nand I_22621 (I387506,I270420,I270420);
not I_22622 (I387523,I387506);
nand I_22623 (I387540,I387523,I387489);
not I_22624 (I387557,I387540);
nand I_22625 (I387574,I270429,I270447);
and I_22626 (I387591,I387574,I270423);
DFFARX1 I_22627 (I387591,I2898,I387472,I387617,);
nor I_22628 (I387625,I270423,I270447);
not I_22629 (I387642,I387625);
nor I_22630 (I387659,I387617,I387625);
DFFARX1 I_22631 (I387659,I2898,I387472,I387443,);
or I_22632 (I387690,I270426,I270441);
nor I_22633 (I387707,I387690,I270429);
not I_22634 (I387724,I387707);
nor I_22635 (I387431,I387617,I387724);
nand I_22636 (I387455,I387506,I387724);
nor I_22637 (I387769,I270426,I270450);
not I_22638 (I387786,I270444);
nor I_22639 (I387803,I387786,I270432);
not I_22640 (I387820,I387803);
nor I_22641 (I387837,I387820,I387540);
nor I_22642 (I387437,I387642,I387837);
nand I_22643 (I387868,I387820,I387642);
nand I_22644 (I387885,I387557,I387868);
nor I_22645 (I387440,I387724,I387885);
nand I_22646 (I387449,I387506,I387820);
nor I_22647 (I387458,I387617,I387803);
nor I_22648 (I387446,I387803,I387557);
nor I_22649 (I387958,I387769,I387786);
nor I_22650 (I387975,I387523,I387958);
nor I_22651 (I387434,I387724,I387975);
nor I_22652 (I388006,I387617,I387958);
nor I_22653 (I387464,I387803,I388006);
nor I_22654 (I387461,I388006,I387642);
and I_22655 (I388051,I387540,I387958);
nor I_22656 (I387452,I387707,I388051);
not I_22657 (I388118,I2905);
or I_22658 (I388135,I41068,I41056);
nand I_22659 (I388152,I41080,I41071);
not I_22660 (I388169,I388152);
nand I_22661 (I388186,I388169,I388135);
not I_22662 (I388203,I388186);
nand I_22663 (I388220,I41059,I41068);
and I_22664 (I388237,I388220,I41077);
DFFARX1 I_22665 (I388237,I2898,I388118,I388263,);
nor I_22666 (I388271,I41062,I41068);
not I_22667 (I388288,I388271);
nor I_22668 (I388305,I388263,I388271);
DFFARX1 I_22669 (I388305,I2898,I388118,I388089,);
or I_22670 (I388336,I41056,I41059);
nor I_22671 (I388353,I388336,I41074);
not I_22672 (I388370,I388353);
nor I_22673 (I388077,I388263,I388370);
nand I_22674 (I388101,I388152,I388370);
nor I_22675 (I388415,I41083,I41065);
not I_22676 (I388432,I41065);
nor I_22677 (I388449,I388432,I41062);
not I_22678 (I388466,I388449);
nor I_22679 (I388483,I388466,I388186);
nor I_22680 (I388083,I388288,I388483);
nand I_22681 (I388514,I388466,I388288);
nand I_22682 (I388531,I388203,I388514);
nor I_22683 (I388086,I388370,I388531);
nand I_22684 (I388095,I388152,I388466);
nor I_22685 (I388104,I388263,I388449);
nor I_22686 (I388092,I388449,I388203);
nor I_22687 (I388604,I388415,I388432);
nor I_22688 (I388621,I388169,I388604);
nor I_22689 (I388080,I388370,I388621);
nor I_22690 (I388652,I388263,I388604);
nor I_22691 (I388110,I388449,I388652);
nor I_22692 (I388107,I388652,I388288);
and I_22693 (I388697,I388186,I388604);
nor I_22694 (I388098,I388353,I388697);
not I_22695 (I388764,I2905);
or I_22696 (I388781,I76433,I76445);
nand I_22697 (I388798,I76445,I76454);
not I_22698 (I388815,I388798);
nand I_22699 (I388832,I388815,I388781);
not I_22700 (I388849,I388832);
nand I_22701 (I388866,I76442,I76436);
and I_22702 (I388883,I388866,I76460);
DFFARX1 I_22703 (I388883,I2898,I388764,I388909,);
nor I_22704 (I388917,I76436,I76436);
not I_22705 (I388934,I388917);
nor I_22706 (I388951,I388909,I388917);
DFFARX1 I_22707 (I388951,I2898,I388764,I388735,);
or I_22708 (I388982,I76448,I76442);
nor I_22709 (I388999,I388982,I76451);
not I_22710 (I389016,I388999);
nor I_22711 (I388723,I388909,I389016);
nand I_22712 (I388747,I388798,I389016);
nor I_22713 (I389061,I76457,I76439);
not I_22714 (I389078,I76439);
nor I_22715 (I389095,I389078,I76433);
not I_22716 (I389112,I389095);
nor I_22717 (I389129,I389112,I388832);
nor I_22718 (I388729,I388934,I389129);
nand I_22719 (I389160,I389112,I388934);
nand I_22720 (I389177,I388849,I389160);
nor I_22721 (I388732,I389016,I389177);
nand I_22722 (I388741,I388798,I389112);
nor I_22723 (I388750,I388909,I389095);
nor I_22724 (I388738,I389095,I388849);
nor I_22725 (I389250,I389061,I389078);
nor I_22726 (I389267,I388815,I389250);
nor I_22727 (I388726,I389016,I389267);
nor I_22728 (I389298,I388909,I389250);
nor I_22729 (I388756,I389095,I389298);
nor I_22730 (I388753,I389298,I388934);
and I_22731 (I389343,I388832,I389250);
nor I_22732 (I388744,I388999,I389343);
not I_22733 (I389410,I2905);
or I_22734 (I389427,I2331,I1667);
nand I_22735 (I389444,I2195,I2347);
not I_22736 (I389461,I389444);
nand I_22737 (I389478,I389461,I389427);
not I_22738 (I389495,I389478);
nand I_22739 (I389512,I1891,I2731);
and I_22740 (I389529,I389512,I2411);
DFFARX1 I_22741 (I389529,I2898,I389410,I389555,);
nor I_22742 (I389563,I2571,I2731);
not I_22743 (I389580,I389563);
nor I_22744 (I389597,I389555,I389563);
DFFARX1 I_22745 (I389597,I2898,I389410,I389381,);
or I_22746 (I389628,I2635,I1979);
nor I_22747 (I389645,I389628,I1651);
not I_22748 (I389662,I389645);
nor I_22749 (I389369,I389555,I389662);
nand I_22750 (I389393,I389444,I389662);
nor I_22751 (I389707,I1579,I2435);
not I_22752 (I389724,I2171);
nor I_22753 (I389741,I389724,I2323);
not I_22754 (I389758,I389741);
nor I_22755 (I389775,I389758,I389478);
nor I_22756 (I389375,I389580,I389775);
nand I_22757 (I389806,I389758,I389580);
nand I_22758 (I389823,I389495,I389806);
nor I_22759 (I389378,I389662,I389823);
nand I_22760 (I389387,I389444,I389758);
nor I_22761 (I389396,I389555,I389741);
nor I_22762 (I389384,I389741,I389495);
nor I_22763 (I389896,I389707,I389724);
nor I_22764 (I389913,I389461,I389896);
nor I_22765 (I389372,I389662,I389913);
nor I_22766 (I389944,I389555,I389896);
nor I_22767 (I389402,I389741,I389944);
nor I_22768 (I389399,I389944,I389580);
and I_22769 (I389989,I389478,I389896);
nor I_22770 (I389390,I389645,I389989);
not I_22771 (I390056,I2905);
or I_22772 (I390073,I116671,I116662);
nand I_22773 (I390090,I116644,I116641);
not I_22774 (I390107,I390090);
nand I_22775 (I390124,I390107,I390073);
not I_22776 (I390141,I390124);
nand I_22777 (I390158,I116641,I116656);
and I_22778 (I390175,I390158,I116638);
DFFARX1 I_22779 (I390175,I2898,I390056,I390201,);
nor I_22780 (I390209,I116644,I116656);
not I_22781 (I390226,I390209);
nor I_22782 (I390243,I390201,I390209);
DFFARX1 I_22783 (I390243,I2898,I390056,I390027,);
or I_22784 (I390274,I116653,I116647);
nor I_22785 (I390291,I390274,I116650);
not I_22786 (I390308,I390291);
nor I_22787 (I390015,I390201,I390308);
nand I_22788 (I390039,I390090,I390308);
nor I_22789 (I390353,I116668,I116659);
not I_22790 (I390370,I116665);
nor I_22791 (I390387,I390370,I116638);
not I_22792 (I390404,I390387);
nor I_22793 (I390421,I390404,I390124);
nor I_22794 (I390021,I390226,I390421);
nand I_22795 (I390452,I390404,I390226);
nand I_22796 (I390469,I390141,I390452);
nor I_22797 (I390024,I390308,I390469);
nand I_22798 (I390033,I390090,I390404);
nor I_22799 (I390042,I390201,I390387);
nor I_22800 (I390030,I390387,I390141);
nor I_22801 (I390542,I390353,I390370);
nor I_22802 (I390559,I390107,I390542);
nor I_22803 (I390018,I390308,I390559);
nor I_22804 (I390590,I390201,I390542);
nor I_22805 (I390048,I390387,I390590);
nor I_22806 (I390045,I390590,I390226);
and I_22807 (I390635,I390124,I390542);
nor I_22808 (I390036,I390291,I390635);
not I_22809 (I390702,I2905);
or I_22810 (I390719,I68256,I68268);
nand I_22811 (I390736,I68268,I68277);
not I_22812 (I390753,I390736);
nand I_22813 (I390770,I390753,I390719);
not I_22814 (I390787,I390770);
nand I_22815 (I390804,I68265,I68259);
and I_22816 (I390821,I390804,I68283);
DFFARX1 I_22817 (I390821,I2898,I390702,I390847,);
nor I_22818 (I390855,I68259,I68259);
not I_22819 (I390872,I390855);
nor I_22820 (I390889,I390847,I390855);
DFFARX1 I_22821 (I390889,I2898,I390702,I390673,);
or I_22822 (I390920,I68271,I68265);
nor I_22823 (I390937,I390920,I68274);
not I_22824 (I390954,I390937);
nor I_22825 (I390661,I390847,I390954);
nand I_22826 (I390685,I390736,I390954);
nor I_22827 (I390999,I68280,I68262);
not I_22828 (I391016,I68262);
nor I_22829 (I391033,I391016,I68256);
not I_22830 (I391050,I391033);
nor I_22831 (I391067,I391050,I390770);
nor I_22832 (I390667,I390872,I391067);
nand I_22833 (I391098,I391050,I390872);
nand I_22834 (I391115,I390787,I391098);
nor I_22835 (I390670,I390954,I391115);
nand I_22836 (I390679,I390736,I391050);
nor I_22837 (I390688,I390847,I391033);
nor I_22838 (I390676,I391033,I390787);
nor I_22839 (I391188,I390999,I391016);
nor I_22840 (I391205,I390753,I391188);
nor I_22841 (I390664,I390954,I391205);
nor I_22842 (I391236,I390847,I391188);
nor I_22843 (I390694,I391033,I391236);
nor I_22844 (I390691,I391236,I390872);
and I_22845 (I391281,I390770,I391188);
nor I_22846 (I390682,I390937,I391281);
not I_22847 (I391348,I2905);
or I_22848 (I391365,I333544,I333544);
nand I_22849 (I391382,I333550,I333562);
not I_22850 (I391399,I391382);
nand I_22851 (I391416,I391399,I391365);
not I_22852 (I391433,I391416);
nand I_22853 (I391450,I333550,I333553);
and I_22854 (I391467,I391450,I333556);
DFFARX1 I_22855 (I391467,I2898,I391348,I391493,);
nor I_22856 (I391501,I333541,I333553);
not I_22857 (I391518,I391501);
nor I_22858 (I391535,I391493,I391501);
DFFARX1 I_22859 (I391535,I2898,I391348,I391319,);
or I_22860 (I391566,I333559,I333547);
nor I_22861 (I391583,I391566,I333541);
not I_22862 (I391600,I391583);
nor I_22863 (I391307,I391493,I391600);
nand I_22864 (I391331,I391382,I391600);
nor I_22865 (I391645,I333556,I333547);
not I_22866 (I391662,I333565);
nor I_22867 (I391679,I391662,I333553);
not I_22868 (I391696,I391679);
nor I_22869 (I391713,I391696,I391416);
nor I_22870 (I391313,I391518,I391713);
nand I_22871 (I391744,I391696,I391518);
nand I_22872 (I391761,I391433,I391744);
nor I_22873 (I391316,I391600,I391761);
nand I_22874 (I391325,I391382,I391696);
nor I_22875 (I391334,I391493,I391679);
nor I_22876 (I391322,I391679,I391433);
nor I_22877 (I391834,I391645,I391662);
nor I_22878 (I391851,I391399,I391834);
nor I_22879 (I391310,I391600,I391851);
nor I_22880 (I391882,I391493,I391834);
nor I_22881 (I391340,I391679,I391882);
nor I_22882 (I391337,I391882,I391518);
and I_22883 (I391927,I391416,I391834);
nor I_22884 (I391328,I391583,I391927);
not I_22885 (I391994,I2905);
or I_22886 (I392011,I121074,I121065);
nand I_22887 (I392028,I121047,I121044);
not I_22888 (I392045,I392028);
nand I_22889 (I392062,I392045,I392011);
not I_22890 (I392079,I392062);
nand I_22891 (I392096,I121044,I121059);
and I_22892 (I392113,I392096,I121041);
DFFARX1 I_22893 (I392113,I2898,I391994,I392139,);
nor I_22894 (I392147,I121047,I121059);
not I_22895 (I392164,I392147);
nor I_22896 (I392181,I392139,I392147);
DFFARX1 I_22897 (I392181,I2898,I391994,I391965,);
or I_22898 (I392212,I121056,I121050);
nor I_22899 (I392229,I392212,I121053);
not I_22900 (I392246,I392229);
nor I_22901 (I391953,I392139,I392246);
nand I_22902 (I391977,I392028,I392246);
nor I_22903 (I392291,I121071,I121062);
not I_22904 (I392308,I121068);
nor I_22905 (I392325,I392308,I121041);
not I_22906 (I392342,I392325);
nor I_22907 (I392359,I392342,I392062);
nor I_22908 (I391959,I392164,I392359);
nand I_22909 (I392390,I392342,I392164);
nand I_22910 (I392407,I392079,I392390);
nor I_22911 (I391962,I392246,I392407);
nand I_22912 (I391971,I392028,I392342);
nor I_22913 (I391980,I392139,I392325);
nor I_22914 (I391968,I392325,I392079);
nor I_22915 (I392480,I392291,I392308);
nor I_22916 (I392497,I392045,I392480);
nor I_22917 (I391956,I392246,I392497);
nor I_22918 (I392528,I392139,I392480);
nor I_22919 (I391986,I392325,I392528);
nor I_22920 (I391983,I392528,I392164);
and I_22921 (I392573,I392062,I392480);
nor I_22922 (I391974,I392229,I392573);
not I_22923 (I392640,I2905);
or I_22924 (I392657,I9646,I9661);
nand I_22925 (I392674,I9667,I9664);
not I_22926 (I392691,I392674);
nand I_22927 (I392708,I392691,I392657);
not I_22928 (I392725,I392708);
nand I_22929 (I392742,I9640,I9643);
and I_22930 (I392759,I392742,I9652);
DFFARX1 I_22931 (I392759,I2898,I392640,I392785,);
nor I_22932 (I392793,I9649,I9643);
not I_22933 (I392810,I392793);
nor I_22934 (I392827,I392785,I392793);
DFFARX1 I_22935 (I392827,I2898,I392640,I392611,);
or I_22936 (I392858,I9643,I9646);
nor I_22937 (I392875,I392858,I9649);
not I_22938 (I392892,I392875);
nor I_22939 (I392599,I392785,I392892);
nand I_22940 (I392623,I392674,I392892);
nor I_22941 (I392937,I9655,I9640);
not I_22942 (I392954,I9658);
nor I_22943 (I392971,I392954,I9670);
not I_22944 (I392988,I392971);
nor I_22945 (I393005,I392988,I392708);
nor I_22946 (I392605,I392810,I393005);
nand I_22947 (I393036,I392988,I392810);
nand I_22948 (I393053,I392725,I393036);
nor I_22949 (I392608,I392892,I393053);
nand I_22950 (I392617,I392674,I392988);
nor I_22951 (I392626,I392785,I392971);
nor I_22952 (I392614,I392971,I392725);
nor I_22953 (I393126,I392937,I392954);
nor I_22954 (I393143,I392691,I393126);
nor I_22955 (I392602,I392892,I393143);
nor I_22956 (I393174,I392785,I393126);
nor I_22957 (I392632,I392971,I393174);
nor I_22958 (I392629,I393174,I392810);
and I_22959 (I393219,I392708,I393126);
nor I_22960 (I392620,I392875,I393219);
not I_22961 (I393286,I2905);
or I_22962 (I393303,I255903,I255900);
nand I_22963 (I393320,I255885,I255885);
not I_22964 (I393337,I393320);
nand I_22965 (I393354,I393337,I393303);
not I_22966 (I393371,I393354);
nand I_22967 (I393388,I255894,I255912);
and I_22968 (I393405,I393388,I255888);
DFFARX1 I_22969 (I393405,I2898,I393286,I393431,);
nor I_22970 (I393439,I255888,I255912);
not I_22971 (I393456,I393439);
nor I_22972 (I393473,I393431,I393439);
DFFARX1 I_22973 (I393473,I2898,I393286,I393257,);
or I_22974 (I393504,I255891,I255906);
nor I_22975 (I393521,I393504,I255894);
not I_22976 (I393538,I393521);
nor I_22977 (I393245,I393431,I393538);
nand I_22978 (I393269,I393320,I393538);
nor I_22979 (I393583,I255891,I255915);
not I_22980 (I393600,I255909);
nor I_22981 (I393617,I393600,I255897);
not I_22982 (I393634,I393617);
nor I_22983 (I393651,I393634,I393354);
nor I_22984 (I393251,I393456,I393651);
nand I_22985 (I393682,I393634,I393456);
nand I_22986 (I393699,I393371,I393682);
nor I_22987 (I393254,I393538,I393699);
nand I_22988 (I393263,I393320,I393634);
nor I_22989 (I393272,I393431,I393617);
nor I_22990 (I393260,I393617,I393371);
nor I_22991 (I393772,I393583,I393600);
nor I_22992 (I393789,I393337,I393772);
nor I_22993 (I393248,I393538,I393789);
nor I_22994 (I393820,I393431,I393772);
nor I_22995 (I393278,I393617,I393820);
nor I_22996 (I393275,I393820,I393456);
and I_22997 (I393865,I393354,I393772);
nor I_22998 (I393266,I393521,I393865);
not I_22999 (I393932,I2905);
or I_23000 (I393949,I47253,I47247);
nand I_23001 (I393966,I47277,I47256);
not I_23002 (I393983,I393966);
nand I_23003 (I394000,I393983,I393949);
not I_23004 (I394017,I394000);
nand I_23005 (I394034,I47262,I47250);
and I_23006 (I394051,I394034,I47244);
DFFARX1 I_23007 (I394051,I2898,I393932,I394077,);
nor I_23008 (I394085,I47274,I47250);
not I_23009 (I394102,I394085);
nor I_23010 (I394119,I394077,I394085);
DFFARX1 I_23011 (I394119,I2898,I393932,I393903,);
or I_23012 (I394150,I47259,I47271);
nor I_23013 (I394167,I394150,I47247);
not I_23014 (I394184,I394167);
nor I_23015 (I393891,I394077,I394184);
nand I_23016 (I393915,I393966,I394184);
nor I_23017 (I394229,I47280,I47244);
not I_23018 (I394246,I47268);
nor I_23019 (I394263,I394246,I47265);
not I_23020 (I394280,I394263);
nor I_23021 (I394297,I394280,I394000);
nor I_23022 (I393897,I394102,I394297);
nand I_23023 (I394328,I394280,I394102);
nand I_23024 (I394345,I394017,I394328);
nor I_23025 (I393900,I394184,I394345);
nand I_23026 (I393909,I393966,I394280);
nor I_23027 (I393918,I394077,I394263);
nor I_23028 (I393906,I394263,I394017);
nor I_23029 (I394418,I394229,I394246);
nor I_23030 (I394435,I393983,I394418);
nor I_23031 (I393894,I394184,I394435);
nor I_23032 (I394466,I394077,I394418);
nor I_23033 (I393924,I394263,I394466);
nor I_23034 (I393921,I394466,I394102);
and I_23035 (I394511,I394000,I394418);
nor I_23036 (I393912,I394167,I394511);
not I_23037 (I394578,I2905);
or I_23038 (I394595,I342469,I342469);
nand I_23039 (I394612,I342475,I342487);
not I_23040 (I394629,I394612);
nand I_23041 (I394646,I394629,I394595);
not I_23042 (I394663,I394646);
nand I_23043 (I394680,I342475,I342478);
and I_23044 (I394697,I394680,I342481);
DFFARX1 I_23045 (I394697,I2898,I394578,I394723,);
nor I_23046 (I394731,I342466,I342478);
not I_23047 (I394748,I394731);
nor I_23048 (I394765,I394723,I394731);
DFFARX1 I_23049 (I394765,I2898,I394578,I394549,);
or I_23050 (I394796,I342484,I342472);
nor I_23051 (I394813,I394796,I342466);
not I_23052 (I394830,I394813);
nor I_23053 (I394537,I394723,I394830);
nand I_23054 (I394561,I394612,I394830);
nor I_23055 (I394875,I342481,I342472);
not I_23056 (I394892,I342490);
nor I_23057 (I394909,I394892,I342478);
not I_23058 (I394926,I394909);
nor I_23059 (I394943,I394926,I394646);
nor I_23060 (I394543,I394748,I394943);
nand I_23061 (I394974,I394926,I394748);
nand I_23062 (I394991,I394663,I394974);
nor I_23063 (I394546,I394830,I394991);
nand I_23064 (I394555,I394612,I394926);
nor I_23065 (I394564,I394723,I394909);
nor I_23066 (I394552,I394909,I394663);
nor I_23067 (I395064,I394875,I394892);
nor I_23068 (I395081,I394629,I395064);
nor I_23069 (I394540,I394830,I395081);
nor I_23070 (I395112,I394723,I395064);
nor I_23071 (I394570,I394909,I395112);
nor I_23072 (I394567,I395112,I394748);
and I_23073 (I395157,I394646,I395064);
nor I_23074 (I394558,I394813,I395157);
not I_23075 (I395215,I2905);
not I_23076 (I395232,I216431);
nand I_23077 (I395249,I216428,I216443);
and I_23078 (I395266,I395249,I216431);
nand I_23079 (I395283,I395249,I395232);
and I_23080 (I395300,I395283,I216440);
nand I_23081 (I395317,I395300,I216440);
or I_23082 (I395334,I216437,I216434);
nor I_23083 (I395351,I395334,I216452);
not I_23084 (I395368,I395351);
and I_23085 (I395385,I395317,I395368);
not I_23086 (I395402,I216434);
nor I_23087 (I395419,I395402,I216449);
nand I_23088 (I395436,I395419,I216437);
not I_23089 (I395453,I395436);
nand I_23090 (I395470,I395453,I395266);
not I_23091 (I395186,I395470);
nor I_23092 (I395189,I395470,I395385);
nand I_23093 (I395192,I395368,I395453);
nand I_23094 (I395529,I395317,I395453);
nand I_23095 (I395546,I395368,I395529);
DFFARX1 I_23096 (I395546,I2898,I395215,I395195,);
nor I_23097 (I395577,I395317,I395402);
and I_23098 (I395594,I395577,I216437);
nor I_23099 (I395204,I395594,I395436);
nand I_23100 (I395625,I395266,I395594);
nand I_23101 (I395207,I395470,I395625);
nand I_23102 (I395656,I216434,I216437);
nor I_23103 (I395673,I216431,I216428);
not I_23104 (I395690,I216446);
nor I_23105 (I395707,I395690,I216455);
nor I_23106 (I395724,I395673,I395690);
not I_23107 (I395741,I395724);
and I_23108 (I395758,I395707,I395741);
nand I_23109 (I395201,I395758,I395656);
nor I_23110 (I395789,I395741,I395436);
not I_23111 (I395806,I395789);
nor I_23112 (I395183,I395707,I395806);
nor I_23113 (I395837,I395724,I395317);
nand I_23114 (I395198,I395837,I395351);
not I_23115 (I395895,I2905);
not I_23116 (I395912,I329388);
nand I_23117 (I395929,I329391,I329379);
and I_23118 (I395946,I395929,I329388);
nand I_23119 (I395963,I395929,I395912);
and I_23120 (I395980,I395963,I329397);
nand I_23121 (I395997,I395980,I329385);
or I_23122 (I396014,I329376,I329391);
nor I_23123 (I396031,I396014,I329379);
not I_23124 (I396048,I396031);
and I_23125 (I396065,I395997,I396048);
not I_23126 (I396082,I329388);
nor I_23127 (I396099,I396082,I329382);
nand I_23128 (I396116,I396099,I329394);
not I_23129 (I396133,I396116);
nand I_23130 (I396150,I396133,I395946);
not I_23131 (I395866,I396150);
nor I_23132 (I395869,I396150,I396065);
nand I_23133 (I395872,I396048,I396133);
nand I_23134 (I396209,I395997,I396133);
nand I_23135 (I396226,I396048,I396209);
DFFARX1 I_23136 (I396226,I2898,I395895,I395875,);
nor I_23137 (I396257,I395997,I396082);
and I_23138 (I396274,I396257,I329394);
nor I_23139 (I395884,I396274,I396116);
nand I_23140 (I396305,I395946,I396274);
nand I_23141 (I395887,I396150,I396305);
nand I_23142 (I396336,I329388,I329394);
nor I_23143 (I396353,I329376,I329385);
not I_23144 (I396370,I329400);
nor I_23145 (I396387,I396370,I329382);
nor I_23146 (I396404,I396353,I396370);
not I_23147 (I396421,I396404);
and I_23148 (I396438,I396387,I396421);
nand I_23149 (I395881,I396438,I396336);
nor I_23150 (I396469,I396421,I396116);
not I_23151 (I396486,I396469);
nor I_23152 (I395863,I396387,I396486);
nor I_23153 (I396517,I396404,I395997);
nand I_23154 (I395878,I396517,I396031);
not I_23155 (I396575,I2905);
not I_23156 (I396592,I338908);
nand I_23157 (I396609,I338911,I338899);
and I_23158 (I396626,I396609,I338908);
nand I_23159 (I396643,I396609,I396592);
and I_23160 (I396660,I396643,I338917);
nand I_23161 (I396677,I396660,I338905);
or I_23162 (I396694,I338896,I338911);
nor I_23163 (I396711,I396694,I338899);
not I_23164 (I396728,I396711);
and I_23165 (I396745,I396677,I396728);
not I_23166 (I396762,I338908);
nor I_23167 (I396779,I396762,I338902);
nand I_23168 (I396796,I396779,I338914);
not I_23169 (I396813,I396796);
nand I_23170 (I396830,I396813,I396626);
not I_23171 (I396546,I396830);
nor I_23172 (I396549,I396830,I396745);
nand I_23173 (I396552,I396728,I396813);
nand I_23174 (I396889,I396677,I396813);
nand I_23175 (I396906,I396728,I396889);
DFFARX1 I_23176 (I396906,I2898,I396575,I396555,);
nor I_23177 (I396937,I396677,I396762);
and I_23178 (I396954,I396937,I338914);
nor I_23179 (I396564,I396954,I396796);
nand I_23180 (I396985,I396626,I396954);
nand I_23181 (I396567,I396830,I396985);
nand I_23182 (I397016,I338908,I338914);
nor I_23183 (I397033,I338896,I338905);
not I_23184 (I397050,I338920);
nor I_23185 (I397067,I397050,I338902);
nor I_23186 (I397084,I397033,I397050);
not I_23187 (I397101,I397084);
and I_23188 (I397118,I397067,I397101);
nand I_23189 (I396561,I397118,I397016);
nor I_23190 (I397149,I397101,I396796);
not I_23191 (I397166,I397149);
nor I_23192 (I396543,I397067,I397166);
nor I_23193 (I397197,I397084,I396677);
nand I_23194 (I396558,I397197,I396711);
not I_23195 (I397255,I2905);
not I_23196 (I397272,I355568);
nand I_23197 (I397289,I355571,I355559);
and I_23198 (I397306,I397289,I355568);
nand I_23199 (I397323,I397289,I397272);
and I_23200 (I397340,I397323,I355577);
nand I_23201 (I397357,I397340,I355565);
or I_23202 (I397374,I355556,I355571);
nor I_23203 (I397391,I397374,I355559);
not I_23204 (I397408,I397391);
and I_23205 (I397425,I397357,I397408);
not I_23206 (I397442,I355568);
nor I_23207 (I397459,I397442,I355562);
nand I_23208 (I397476,I397459,I355574);
not I_23209 (I397493,I397476);
nand I_23210 (I397510,I397493,I397306);
not I_23211 (I397226,I397510);
nor I_23212 (I397229,I397510,I397425);
nand I_23213 (I397232,I397408,I397493);
nand I_23214 (I397569,I397357,I397493);
nand I_23215 (I397586,I397408,I397569);
DFFARX1 I_23216 (I397586,I2898,I397255,I397235,);
nor I_23217 (I397617,I397357,I397442);
and I_23218 (I397634,I397617,I355574);
nor I_23219 (I397244,I397634,I397476);
nand I_23220 (I397665,I397306,I397634);
nand I_23221 (I397247,I397510,I397665);
nand I_23222 (I397696,I355568,I355574);
nor I_23223 (I397713,I355556,I355565);
not I_23224 (I397730,I355580);
nor I_23225 (I397747,I397730,I355562);
nor I_23226 (I397764,I397713,I397730);
not I_23227 (I397781,I397764);
and I_23228 (I397798,I397747,I397781);
nand I_23229 (I397241,I397798,I397696);
nor I_23230 (I397829,I397781,I397476);
not I_23231 (I397846,I397829);
nor I_23232 (I397223,I397747,I397846);
nor I_23233 (I397877,I397764,I397357);
nand I_23234 (I397238,I397877,I397391);
not I_23235 (I397935,I2905);
not I_23236 (I397952,I348428);
nand I_23237 (I397969,I348431,I348419);
and I_23238 (I397986,I397969,I348428);
nand I_23239 (I398003,I397969,I397952);
and I_23240 (I398020,I398003,I348437);
nand I_23241 (I398037,I398020,I348425);
or I_23242 (I398054,I348416,I348431);
nor I_23243 (I398071,I398054,I348419);
not I_23244 (I398088,I398071);
and I_23245 (I398105,I398037,I398088);
not I_23246 (I398122,I348428);
nor I_23247 (I398139,I398122,I348422);
nand I_23248 (I398156,I398139,I348434);
not I_23249 (I398173,I398156);
nand I_23250 (I398190,I398173,I397986);
not I_23251 (I397906,I398190);
nor I_23252 (I397909,I398190,I398105);
nand I_23253 (I397912,I398088,I398173);
nand I_23254 (I398249,I398037,I398173);
nand I_23255 (I398266,I398088,I398249);
DFFARX1 I_23256 (I398266,I2898,I397935,I397915,);
nor I_23257 (I398297,I398037,I398122);
and I_23258 (I398314,I398297,I348434);
nor I_23259 (I397924,I398314,I398156);
nand I_23260 (I398345,I397986,I398314);
nand I_23261 (I397927,I398190,I398345);
nand I_23262 (I398376,I348428,I348434);
nor I_23263 (I398393,I348416,I348425);
not I_23264 (I398410,I348440);
nor I_23265 (I398427,I398410,I348422);
nor I_23266 (I398444,I398393,I398410);
not I_23267 (I398461,I398444);
and I_23268 (I398478,I398427,I398461);
nand I_23269 (I397921,I398478,I398376);
nor I_23270 (I398509,I398461,I398156);
not I_23271 (I398526,I398509);
nor I_23272 (I397903,I398427,I398526);
nor I_23273 (I398557,I398444,I398037);
nand I_23274 (I397918,I398557,I398071);
not I_23275 (I398615,I2905);
not I_23276 (I398632,I195309);
nand I_23277 (I398649,I195318,I195297);
and I_23278 (I398666,I398649,I195309);
nand I_23279 (I398683,I398649,I398632);
and I_23280 (I398700,I398683,I195312);
nand I_23281 (I398717,I398700,I195300);
or I_23282 (I398734,I195315,I195303);
nor I_23283 (I398751,I398734,I195306);
not I_23284 (I398768,I398751);
and I_23285 (I398785,I398717,I398768);
not I_23286 (I398802,I195309);
nor I_23287 (I398819,I398802,I195306);
nand I_23288 (I398836,I398819,I195312);
not I_23289 (I398853,I398836);
nand I_23290 (I398870,I398853,I398666);
not I_23291 (I398586,I398870);
nor I_23292 (I398589,I398870,I398785);
nand I_23293 (I398592,I398768,I398853);
nand I_23294 (I398929,I398717,I398853);
nand I_23295 (I398946,I398768,I398929);
DFFARX1 I_23296 (I398946,I2898,I398615,I398595,);
nor I_23297 (I398977,I398717,I398802);
and I_23298 (I398994,I398977,I195312);
nor I_23299 (I398604,I398994,I398836);
nand I_23300 (I399025,I398666,I398994);
nand I_23301 (I398607,I398870,I399025);
nand I_23302 (I399056,I195309,I195312);
nor I_23303 (I399073,I195300,I195297);
not I_23304 (I399090,I195303);
nor I_23305 (I399107,I399090,I195321);
nor I_23306 (I399124,I399073,I399090);
not I_23307 (I399141,I399124);
and I_23308 (I399158,I399107,I399141);
nand I_23309 (I398601,I399158,I399056);
nor I_23310 (I399189,I399141,I398836);
not I_23311 (I399206,I399189);
nor I_23312 (I398583,I399107,I399206);
nor I_23313 (I399237,I399124,I398717);
nand I_23314 (I398598,I399237,I398751);
not I_23315 (I399295,I2905);
not I_23316 (I399312,I28930);
nand I_23317 (I399329,I28942,I28924);
and I_23318 (I399346,I399329,I28930);
nand I_23319 (I399363,I399329,I399312);
and I_23320 (I399380,I399363,I28939);
nand I_23321 (I399397,I399380,I28918);
or I_23322 (I399414,I28924,I28927);
nor I_23323 (I399431,I399414,I28921);
not I_23324 (I399448,I399431);
and I_23325 (I399465,I399397,I399448);
not I_23326 (I399482,I28930);
nor I_23327 (I399499,I399482,I28921);
nand I_23328 (I399516,I399499,I28933);
not I_23329 (I399533,I399516);
nand I_23330 (I399550,I399533,I399346);
not I_23331 (I399266,I399550);
nor I_23332 (I399269,I399550,I399465);
nand I_23333 (I399272,I399448,I399533);
nand I_23334 (I399609,I399397,I399533);
nand I_23335 (I399626,I399448,I399609);
DFFARX1 I_23336 (I399626,I2898,I399295,I399275,);
nor I_23337 (I399657,I399397,I399482);
and I_23338 (I399674,I399657,I28933);
nor I_23339 (I399284,I399674,I399516);
nand I_23340 (I399705,I399346,I399674);
nand I_23341 (I399287,I399550,I399705);
nand I_23342 (I399736,I28930,I28933);
nor I_23343 (I399753,I28945,I28918);
not I_23344 (I399770,I28936);
nor I_23345 (I399787,I399770,I28927);
nor I_23346 (I399804,I399753,I399770);
not I_23347 (I399821,I399804);
and I_23348 (I399838,I399787,I399821);
nand I_23349 (I399281,I399838,I399736);
nor I_23350 (I399869,I399821,I399516);
not I_23351 (I399886,I399869);
nor I_23352 (I399263,I399787,I399886);
nor I_23353 (I399917,I399804,I399397);
nand I_23354 (I399278,I399917,I399431);
not I_23355 (I399975,I2905);
not I_23356 (I399992,I336528);
nand I_23357 (I400009,I336531,I336519);
and I_23358 (I400026,I400009,I336528);
nand I_23359 (I400043,I400009,I399992);
and I_23360 (I400060,I400043,I336537);
nand I_23361 (I400077,I400060,I336525);
or I_23362 (I400094,I336516,I336531);
nor I_23363 (I400111,I400094,I336519);
not I_23364 (I400128,I400111);
and I_23365 (I400145,I400077,I400128);
not I_23366 (I400162,I336528);
nor I_23367 (I400179,I400162,I336522);
nand I_23368 (I400196,I400179,I336534);
not I_23369 (I400213,I400196);
nand I_23370 (I400230,I400213,I400026);
not I_23371 (I399946,I400230);
nor I_23372 (I399949,I400230,I400145);
nand I_23373 (I399952,I400128,I400213);
nand I_23374 (I400289,I400077,I400213);
nand I_23375 (I400306,I400128,I400289);
DFFARX1 I_23376 (I400306,I2898,I399975,I399955,);
nor I_23377 (I400337,I400077,I400162);
and I_23378 (I400354,I400337,I336534);
nor I_23379 (I399964,I400354,I400196);
nand I_23380 (I400385,I400026,I400354);
nand I_23381 (I399967,I400230,I400385);
nand I_23382 (I400416,I336528,I336534);
nor I_23383 (I400433,I336516,I336525);
not I_23384 (I400450,I336540);
nor I_23385 (I400467,I400450,I336522);
nor I_23386 (I400484,I400433,I400450);
not I_23387 (I400501,I400484);
and I_23388 (I400518,I400467,I400501);
nand I_23389 (I399961,I400518,I400416);
nor I_23390 (I400549,I400501,I400196);
not I_23391 (I400566,I400549);
nor I_23392 (I399943,I400467,I400566);
nor I_23393 (I400597,I400484,I400077);
nand I_23394 (I399958,I400597,I400111);
not I_23395 (I400655,I2905);
not I_23396 (I400672,I205211);
nand I_23397 (I400689,I205208,I205223);
and I_23398 (I400706,I400689,I205211);
nand I_23399 (I400723,I400689,I400672);
and I_23400 (I400740,I400723,I205220);
nand I_23401 (I400757,I400740,I205220);
or I_23402 (I400774,I205217,I205214);
nor I_23403 (I400791,I400774,I205232);
not I_23404 (I400808,I400791);
and I_23405 (I400825,I400757,I400808);
not I_23406 (I400842,I205214);
nor I_23407 (I400859,I400842,I205229);
nand I_23408 (I400876,I400859,I205217);
not I_23409 (I400893,I400876);
nand I_23410 (I400910,I400893,I400706);
not I_23411 (I400626,I400910);
nor I_23412 (I400629,I400910,I400825);
nand I_23413 (I400632,I400808,I400893);
nand I_23414 (I400969,I400757,I400893);
nand I_23415 (I400986,I400808,I400969);
DFFARX1 I_23416 (I400986,I2898,I400655,I400635,);
nor I_23417 (I401017,I400757,I400842);
and I_23418 (I401034,I401017,I205217);
nor I_23419 (I400644,I401034,I400876);
nand I_23420 (I401065,I400706,I401034);
nand I_23421 (I400647,I400910,I401065);
nand I_23422 (I401096,I205214,I205217);
nor I_23423 (I401113,I205211,I205208);
not I_23424 (I401130,I205226);
nor I_23425 (I401147,I401130,I205235);
nor I_23426 (I401164,I401113,I401130);
not I_23427 (I401181,I401164);
and I_23428 (I401198,I401147,I401181);
nand I_23429 (I400641,I401198,I401096);
nor I_23430 (I401229,I401181,I400876);
not I_23431 (I401246,I401229);
nor I_23432 (I400623,I401147,I401246);
nor I_23433 (I401277,I401164,I400757);
nand I_23434 (I400638,I401277,I400791);
not I_23435 (I401335,I2905);
not I_23436 (I401352,I377765);
nand I_23437 (I401369,I377768,I377762);
and I_23438 (I401386,I401369,I377765);
nand I_23439 (I401403,I401369,I401352);
and I_23440 (I401420,I401403,I377747);
nand I_23441 (I401437,I401420,I377759);
or I_23442 (I401454,I377771,I377774);
nor I_23443 (I401471,I401454,I377753);
not I_23444 (I401488,I401471);
and I_23445 (I401505,I401437,I401488);
not I_23446 (I401522,I377744);
nor I_23447 (I401539,I401522,I377741);
nand I_23448 (I401556,I401539,I377744);
not I_23449 (I401573,I401556);
nand I_23450 (I401590,I401573,I401386);
not I_23451 (I401306,I401590);
nor I_23452 (I401309,I401590,I401505);
nand I_23453 (I401312,I401488,I401573);
nand I_23454 (I401649,I401437,I401573);
nand I_23455 (I401666,I401488,I401649);
DFFARX1 I_23456 (I401666,I2898,I401335,I401315,);
nor I_23457 (I401697,I401437,I401522);
and I_23458 (I401714,I401697,I377744);
nor I_23459 (I401324,I401714,I401556);
nand I_23460 (I401745,I401386,I401714);
nand I_23461 (I401327,I401590,I401745);
nand I_23462 (I401776,I377744,I377744);
nor I_23463 (I401793,I377756,I377747);
not I_23464 (I401810,I377741);
nor I_23465 (I401827,I401810,I377750);
nor I_23466 (I401844,I401793,I401810);
not I_23467 (I401861,I401844);
and I_23468 (I401878,I401827,I401861);
nand I_23469 (I401321,I401878,I401776);
nor I_23470 (I401909,I401861,I401556);
not I_23471 (I401926,I401909);
nor I_23472 (I401303,I401827,I401926);
nor I_23473 (I401957,I401844,I401437);
nand I_23474 (I401318,I401957,I401471);
not I_23475 (I402015,I2905);
not I_23476 (I402032,I351998);
nand I_23477 (I402049,I352001,I351989);
and I_23478 (I402066,I402049,I351998);
nand I_23479 (I402083,I402049,I402032);
and I_23480 (I402100,I402083,I352007);
nand I_23481 (I402117,I402100,I351995);
or I_23482 (I402134,I351986,I352001);
nor I_23483 (I402151,I402134,I351989);
not I_23484 (I402168,I402151);
and I_23485 (I402185,I402117,I402168);
not I_23486 (I402202,I351998);
nor I_23487 (I402219,I402202,I351992);
nand I_23488 (I402236,I402219,I352004);
not I_23489 (I402253,I402236);
nand I_23490 (I402270,I402253,I402066);
not I_23491 (I401986,I402270);
nor I_23492 (I401989,I402270,I402185);
nand I_23493 (I401992,I402168,I402253);
nand I_23494 (I402329,I402117,I402253);
nand I_23495 (I402346,I402168,I402329);
DFFARX1 I_23496 (I402346,I2898,I402015,I401995,);
nor I_23497 (I402377,I402117,I402202);
and I_23498 (I402394,I402377,I352004);
nor I_23499 (I402004,I402394,I402236);
nand I_23500 (I402425,I402066,I402394);
nand I_23501 (I402007,I402270,I402425);
nand I_23502 (I402456,I351998,I352004);
nor I_23503 (I402473,I351986,I351995);
not I_23504 (I402490,I352010);
nor I_23505 (I402507,I402490,I351992);
nor I_23506 (I402524,I402473,I402490);
not I_23507 (I402541,I402524);
and I_23508 (I402558,I402507,I402541);
nand I_23509 (I402001,I402558,I402456);
nor I_23510 (I402589,I402541,I402236);
not I_23511 (I402606,I402589);
nor I_23512 (I401983,I402507,I402606);
nor I_23513 (I402637,I402524,I402117);
nand I_23514 (I401998,I402637,I402151);
not I_23515 (I402695,I2905);
not I_23516 (I402712,I364102);
nand I_23517 (I402729,I364090,I364096);
and I_23518 (I402746,I402729,I364102);
nand I_23519 (I402763,I402729,I402712);
and I_23520 (I402780,I402763,I364090);
nand I_23521 (I402797,I402780,I364120);
or I_23522 (I402814,I364096,I364123);
nor I_23523 (I402831,I402814,I364093);
not I_23524 (I402848,I402831);
and I_23525 (I402865,I402797,I402848);
not I_23526 (I402882,I364114);
nor I_23527 (I402899,I402882,I364111);
nand I_23528 (I402916,I402899,I364105);
not I_23529 (I402933,I402916);
nand I_23530 (I402950,I402933,I402746);
not I_23531 (I402666,I402950);
nor I_23532 (I402669,I402950,I402865);
nand I_23533 (I402672,I402848,I402933);
nand I_23534 (I403009,I402797,I402933);
nand I_23535 (I403026,I402848,I403009);
DFFARX1 I_23536 (I403026,I2898,I402695,I402675,);
nor I_23537 (I403057,I402797,I402882);
and I_23538 (I403074,I403057,I364105);
nor I_23539 (I402684,I403074,I402916);
nand I_23540 (I403105,I402746,I403074);
nand I_23541 (I402687,I402950,I403105);
nand I_23542 (I403136,I364114,I364105);
nor I_23543 (I403153,I364108,I364117);
not I_23544 (I403170,I364099);
nor I_23545 (I403187,I403170,I364093);
nor I_23546 (I403204,I403153,I403170);
not I_23547 (I403221,I403204);
and I_23548 (I403238,I403187,I403221);
nand I_23549 (I402681,I403238,I403136);
nor I_23550 (I403269,I403221,I402916);
not I_23551 (I403286,I403269);
nor I_23552 (I402663,I403187,I403286);
nor I_23553 (I403317,I403204,I402797);
nand I_23554 (I402678,I403317,I402831);
not I_23555 (I403375,I2905);
not I_23556 (I403392,I223911);
nand I_23557 (I403409,I223908,I223923);
and I_23558 (I403426,I403409,I223911);
nand I_23559 (I403443,I403409,I403392);
and I_23560 (I403460,I403443,I223920);
nand I_23561 (I403477,I403460,I223920);
or I_23562 (I403494,I223917,I223914);
nor I_23563 (I403511,I403494,I223932);
not I_23564 (I403528,I403511);
and I_23565 (I403545,I403477,I403528);
not I_23566 (I403562,I223914);
nor I_23567 (I403579,I403562,I223929);
nand I_23568 (I403596,I403579,I223917);
not I_23569 (I403613,I403596);
nand I_23570 (I403630,I403613,I403426);
not I_23571 (I403346,I403630);
nor I_23572 (I403349,I403630,I403545);
nand I_23573 (I403352,I403528,I403613);
nand I_23574 (I403689,I403477,I403613);
nand I_23575 (I403706,I403528,I403689);
DFFARX1 I_23576 (I403706,I2898,I403375,I403355,);
nor I_23577 (I403737,I403477,I403562);
and I_23578 (I403754,I403737,I223917);
nor I_23579 (I403364,I403754,I403596);
nand I_23580 (I403785,I403426,I403754);
nand I_23581 (I403367,I403630,I403785);
nand I_23582 (I403816,I223914,I223917);
nor I_23583 (I403833,I223911,I223908);
not I_23584 (I403850,I223926);
nor I_23585 (I403867,I403850,I223935);
nor I_23586 (I403884,I403833,I403850);
not I_23587 (I403901,I403884);
and I_23588 (I403918,I403867,I403901);
nand I_23589 (I403361,I403918,I403816);
nor I_23590 (I403949,I403901,I403596);
not I_23591 (I403966,I403949);
nor I_23592 (I403343,I403867,I403966);
nor I_23593 (I403997,I403884,I403477);
nand I_23594 (I403358,I403997,I403511);
not I_23595 (I404055,I2905);
not I_23596 (I404072,I2883);
nand I_23597 (I404089,I2443,I1819);
and I_23598 (I404106,I404089,I2883);
nand I_23599 (I404123,I404089,I404072);
and I_23600 (I404140,I404123,I1675);
nand I_23601 (I404157,I404140,I1763);
or I_23602 (I404174,I1963,I1707);
nor I_23603 (I404191,I404174,I1619);
not I_23604 (I404208,I404191);
and I_23605 (I404225,I404157,I404208);
not I_23606 (I404242,I2379);
nor I_23607 (I404259,I404242,I2003);
nand I_23608 (I404276,I404259,I2779);
not I_23609 (I404293,I404276);
nand I_23610 (I404310,I404293,I404106);
not I_23611 (I404026,I404310);
nor I_23612 (I404029,I404310,I404225);
nand I_23613 (I404032,I404208,I404293);
nand I_23614 (I404369,I404157,I404293);
nand I_23615 (I404386,I404208,I404369);
DFFARX1 I_23616 (I404386,I2898,I404055,I404035,);
nor I_23617 (I404417,I404157,I404242);
and I_23618 (I404434,I404417,I2779);
nor I_23619 (I404044,I404434,I404276);
nand I_23620 (I404465,I404106,I404434);
nand I_23621 (I404047,I404310,I404465);
nand I_23622 (I404496,I2379,I2779);
nor I_23623 (I404513,I1627,I2659);
not I_23624 (I404530,I2187);
nor I_23625 (I404547,I404530,I2139);
nor I_23626 (I404564,I404513,I404530);
not I_23627 (I404581,I404564);
and I_23628 (I404598,I404547,I404581);
nand I_23629 (I404041,I404598,I404496);
nor I_23630 (I404629,I404581,I404276);
not I_23631 (I404646,I404629);
nor I_23632 (I404023,I404547,I404646);
nor I_23633 (I404677,I404564,I404157);
nand I_23634 (I404038,I404677,I404191);
not I_23635 (I404735,I2905);
not I_23636 (I404752,I356758);
nand I_23637 (I404769,I356761,I356749);
and I_23638 (I404786,I404769,I356758);
nand I_23639 (I404803,I404769,I404752);
and I_23640 (I404820,I404803,I356767);
nand I_23641 (I404837,I404820,I356755);
or I_23642 (I404854,I356746,I356761);
nor I_23643 (I404871,I404854,I356749);
not I_23644 (I404888,I404871);
and I_23645 (I404905,I404837,I404888);
not I_23646 (I404922,I356758);
nor I_23647 (I404939,I404922,I356752);
nand I_23648 (I404956,I404939,I356764);
not I_23649 (I404973,I404956);
nand I_23650 (I404990,I404973,I404786);
not I_23651 (I404706,I404990);
nor I_23652 (I404709,I404990,I404905);
nand I_23653 (I404712,I404888,I404973);
nand I_23654 (I405049,I404837,I404973);
nand I_23655 (I405066,I404888,I405049);
DFFARX1 I_23656 (I405066,I2898,I404735,I404715,);
nor I_23657 (I405097,I404837,I404922);
and I_23658 (I405114,I405097,I356764);
nor I_23659 (I404724,I405114,I404956);
nand I_23660 (I405145,I404786,I405114);
nand I_23661 (I404727,I404990,I405145);
nand I_23662 (I405176,I356758,I356764);
nor I_23663 (I405193,I356746,I356755);
not I_23664 (I405210,I356770);
nor I_23665 (I405227,I405210,I356752);
nor I_23666 (I405244,I405193,I405210);
not I_23667 (I405261,I405244);
and I_23668 (I405278,I405227,I405261);
nand I_23669 (I404721,I405278,I405176);
nor I_23670 (I405309,I405261,I404956);
not I_23671 (I405326,I405309);
nor I_23672 (I404703,I405227,I405326);
nor I_23673 (I405357,I405244,I404837);
nand I_23674 (I404718,I405357,I404871);
not I_23675 (I405415,I2905);
not I_23676 (I405432,I181310);
nand I_23677 (I405449,I181301,I181304);
and I_23678 (I405466,I405449,I181310);
nand I_23679 (I405483,I405449,I405432);
and I_23680 (I405500,I405483,I181298);
nand I_23681 (I405517,I405500,I181298);
or I_23682 (I405534,I181316,I181292);
nor I_23683 (I405551,I405534,I181289);
not I_23684 (I405568,I405551);
and I_23685 (I405585,I405517,I405568);
not I_23686 (I405602,I181289);
nor I_23687 (I405619,I405602,I181307);
nand I_23688 (I405636,I405619,I181313);
not I_23689 (I405653,I405636);
nand I_23690 (I405670,I405653,I405466);
not I_23691 (I405386,I405670);
nor I_23692 (I405389,I405670,I405585);
nand I_23693 (I405392,I405568,I405653);
nand I_23694 (I405729,I405517,I405653);
nand I_23695 (I405746,I405568,I405729);
DFFARX1 I_23696 (I405746,I2898,I405415,I405395,);
nor I_23697 (I405777,I405517,I405602);
and I_23698 (I405794,I405777,I181313);
nor I_23699 (I405404,I405794,I405636);
nand I_23700 (I405825,I405466,I405794);
nand I_23701 (I405407,I405670,I405825);
nand I_23702 (I405856,I181289,I181313);
nor I_23703 (I405873,I181295,I181292);
not I_23704 (I405890,I181319);
nor I_23705 (I405907,I405890,I181295);
nor I_23706 (I405924,I405873,I405890);
not I_23707 (I405941,I405924);
and I_23708 (I405958,I405907,I405941);
nand I_23709 (I405401,I405958,I405856);
nor I_23710 (I405989,I405941,I405636);
not I_23711 (I406006,I405989);
nor I_23712 (I405383,I405907,I406006);
nor I_23713 (I406037,I405924,I405517);
nand I_23714 (I405398,I406037,I405551);
not I_23715 (I406095,I2905);
not I_23716 (I406112,I391977);
nand I_23717 (I406129,I391980,I391974);
and I_23718 (I406146,I406129,I391977);
nand I_23719 (I406163,I406129,I406112);
and I_23720 (I406180,I406163,I391959);
nand I_23721 (I406197,I406180,I391971);
or I_23722 (I406214,I391983,I391986);
nor I_23723 (I406231,I406214,I391965);
not I_23724 (I406248,I406231);
and I_23725 (I406265,I406197,I406248);
not I_23726 (I406282,I391956);
nor I_23727 (I406299,I406282,I391953);
nand I_23728 (I406316,I406299,I391956);
not I_23729 (I406333,I406316);
nand I_23730 (I406350,I406333,I406146);
not I_23731 (I406066,I406350);
nor I_23732 (I406069,I406350,I406265);
nand I_23733 (I406072,I406248,I406333);
nand I_23734 (I406409,I406197,I406333);
nand I_23735 (I406426,I406248,I406409);
DFFARX1 I_23736 (I406426,I2898,I406095,I406075,);
nor I_23737 (I406457,I406197,I406282);
and I_23738 (I406474,I406457,I391956);
nor I_23739 (I406084,I406474,I406316);
nand I_23740 (I406505,I406146,I406474);
nand I_23741 (I406087,I406350,I406505);
nand I_23742 (I406536,I391956,I391956);
nor I_23743 (I406553,I391968,I391959);
not I_23744 (I406570,I391953);
nor I_23745 (I406587,I406570,I391962);
nor I_23746 (I406604,I406553,I406570);
not I_23747 (I406621,I406604);
and I_23748 (I406638,I406587,I406621);
nand I_23749 (I406081,I406638,I406536);
nor I_23750 (I406669,I406621,I406316);
not I_23751 (I406686,I406669);
nor I_23752 (I406063,I406587,I406686);
nor I_23753 (I406717,I406604,I406197);
nand I_23754 (I406078,I406717,I406231);
not I_23755 (I406775,I2905);
not I_23756 (I406792,I371305);
nand I_23757 (I406809,I371308,I371302);
and I_23758 (I406826,I406809,I371305);
nand I_23759 (I406843,I406809,I406792);
and I_23760 (I406860,I406843,I371287);
nand I_23761 (I406877,I406860,I371299);
or I_23762 (I406894,I371311,I371314);
nor I_23763 (I406911,I406894,I371293);
not I_23764 (I406928,I406911);
and I_23765 (I406945,I406877,I406928);
not I_23766 (I406962,I371284);
nor I_23767 (I406979,I406962,I371281);
nand I_23768 (I406996,I406979,I371284);
not I_23769 (I407013,I406996);
nand I_23770 (I407030,I407013,I406826);
not I_23771 (I406746,I407030);
nor I_23772 (I406749,I407030,I406945);
nand I_23773 (I406752,I406928,I407013);
nand I_23774 (I407089,I406877,I407013);
nand I_23775 (I407106,I406928,I407089);
DFFARX1 I_23776 (I407106,I2898,I406775,I406755,);
nor I_23777 (I407137,I406877,I406962);
and I_23778 (I407154,I407137,I371284);
nor I_23779 (I406764,I407154,I406996);
nand I_23780 (I407185,I406826,I407154);
nand I_23781 (I406767,I407030,I407185);
nand I_23782 (I407216,I371284,I371284);
nor I_23783 (I407233,I371296,I371287);
not I_23784 (I407250,I371281);
nor I_23785 (I407267,I407250,I371290);
nor I_23786 (I407284,I407233,I407250);
not I_23787 (I407301,I407284);
and I_23788 (I407318,I407267,I407301);
nand I_23789 (I406761,I407318,I407216);
nor I_23790 (I407349,I407301,I406996);
not I_23791 (I407366,I407349);
nor I_23792 (I406743,I407267,I407366);
nor I_23793 (I407397,I407284,I406877);
nand I_23794 (I406758,I407397,I406911);
not I_23795 (I407455,I2905);
not I_23796 (I407472,I384225);
nand I_23797 (I407489,I384228,I384222);
and I_23798 (I407506,I407489,I384225);
nand I_23799 (I407523,I407489,I407472);
and I_23800 (I407540,I407523,I384207);
nand I_23801 (I407557,I407540,I384219);
or I_23802 (I407574,I384231,I384234);
nor I_23803 (I407591,I407574,I384213);
not I_23804 (I407608,I407591);
and I_23805 (I407625,I407557,I407608);
not I_23806 (I407642,I384204);
nor I_23807 (I407659,I407642,I384201);
nand I_23808 (I407676,I407659,I384204);
not I_23809 (I407693,I407676);
nand I_23810 (I407710,I407693,I407506);
not I_23811 (I407426,I407710);
nor I_23812 (I407429,I407710,I407625);
nand I_23813 (I407432,I407608,I407693);
nand I_23814 (I407769,I407557,I407693);
nand I_23815 (I407786,I407608,I407769);
DFFARX1 I_23816 (I407786,I2898,I407455,I407435,);
nor I_23817 (I407817,I407557,I407642);
and I_23818 (I407834,I407817,I384204);
nor I_23819 (I407444,I407834,I407676);
nand I_23820 (I407865,I407506,I407834);
nand I_23821 (I407447,I407710,I407865);
nand I_23822 (I407896,I384204,I384204);
nor I_23823 (I407913,I384216,I384207);
not I_23824 (I407930,I384201);
nor I_23825 (I407947,I407930,I384210);
nor I_23826 (I407964,I407913,I407930);
not I_23827 (I407981,I407964);
and I_23828 (I407998,I407947,I407981);
nand I_23829 (I407441,I407998,I407896);
nor I_23830 (I408029,I407981,I407676);
not I_23831 (I408046,I408029);
nor I_23832 (I407423,I407947,I408046);
nor I_23833 (I408077,I407964,I407557);
nand I_23834 (I407438,I408077,I407591);
not I_23835 (I408135,I2905);
not I_23836 (I408152,I352593);
nand I_23837 (I408169,I352596,I352584);
and I_23838 (I408186,I408169,I352593);
nand I_23839 (I408203,I408169,I408152);
and I_23840 (I408220,I408203,I352602);
nand I_23841 (I408237,I408220,I352590);
or I_23842 (I408254,I352581,I352596);
nor I_23843 (I408271,I408254,I352584);
not I_23844 (I408288,I408271);
and I_23845 (I408305,I408237,I408288);
not I_23846 (I408322,I352593);
nor I_23847 (I408339,I408322,I352587);
nand I_23848 (I408356,I408339,I352599);
not I_23849 (I408373,I408356);
nand I_23850 (I408390,I408373,I408186);
not I_23851 (I408106,I408390);
nor I_23852 (I408109,I408390,I408305);
nand I_23853 (I408112,I408288,I408373);
nand I_23854 (I408449,I408237,I408373);
nand I_23855 (I408466,I408288,I408449);
DFFARX1 I_23856 (I408466,I2898,I408135,I408115,);
nor I_23857 (I408497,I408237,I408322);
and I_23858 (I408514,I408497,I352599);
nor I_23859 (I408124,I408514,I408356);
nand I_23860 (I408545,I408186,I408514);
nand I_23861 (I408127,I408390,I408545);
nand I_23862 (I408576,I352593,I352599);
nor I_23863 (I408593,I352581,I352590);
not I_23864 (I408610,I352605);
nor I_23865 (I408627,I408610,I352587);
nor I_23866 (I408644,I408593,I408610);
not I_23867 (I408661,I408644);
and I_23868 (I408678,I408627,I408661);
nand I_23869 (I408121,I408678,I408576);
nor I_23870 (I408709,I408661,I408356);
not I_23871 (I408726,I408709);
nor I_23872 (I408103,I408627,I408726);
nor I_23873 (I408757,I408644,I408237);
nand I_23874 (I408118,I408757,I408271);
not I_23875 (I408815,I2905);
not I_23876 (I408832,I204463);
nand I_23877 (I408849,I204460,I204475);
and I_23878 (I408866,I408849,I204463);
nand I_23879 (I408883,I408849,I408832);
and I_23880 (I408900,I408883,I204472);
nand I_23881 (I408917,I408900,I204472);
or I_23882 (I408934,I204469,I204466);
nor I_23883 (I408951,I408934,I204484);
not I_23884 (I408968,I408951);
and I_23885 (I408985,I408917,I408968);
not I_23886 (I409002,I204466);
nor I_23887 (I409019,I409002,I204481);
nand I_23888 (I409036,I409019,I204469);
not I_23889 (I409053,I409036);
nand I_23890 (I409070,I409053,I408866);
not I_23891 (I408786,I409070);
nor I_23892 (I408789,I409070,I408985);
nand I_23893 (I408792,I408968,I409053);
nand I_23894 (I409129,I408917,I409053);
nand I_23895 (I409146,I408968,I409129);
DFFARX1 I_23896 (I409146,I2898,I408815,I408795,);
nor I_23897 (I409177,I408917,I409002);
and I_23898 (I409194,I409177,I204469);
nor I_23899 (I408804,I409194,I409036);
nand I_23900 (I409225,I408866,I409194);
nand I_23901 (I408807,I409070,I409225);
nand I_23902 (I409256,I204466,I204469);
nor I_23903 (I409273,I204463,I204460);
not I_23904 (I409290,I204478);
nor I_23905 (I409307,I409290,I204487);
nor I_23906 (I409324,I409273,I409290);
not I_23907 (I409341,I409324);
and I_23908 (I409358,I409307,I409341);
nand I_23909 (I408801,I409358,I409256);
nor I_23910 (I409389,I409341,I409036);
not I_23911 (I409406,I409389);
nor I_23912 (I408783,I409307,I409406);
nor I_23913 (I409437,I409324,I408917);
nand I_23914 (I408798,I409437,I408951);
not I_23915 (I409495,I2905);
not I_23916 (I409512,I21076);
nand I_23917 (I409529,I21088,I21070);
and I_23918 (I409546,I409529,I21076);
nand I_23919 (I409563,I409529,I409512);
and I_23920 (I409580,I409563,I21085);
nand I_23921 (I409597,I409580,I21064);
or I_23922 (I409614,I21070,I21073);
nor I_23923 (I409631,I409614,I21067);
not I_23924 (I409648,I409631);
and I_23925 (I409665,I409597,I409648);
not I_23926 (I409682,I21076);
nor I_23927 (I409699,I409682,I21067);
nand I_23928 (I409716,I409699,I21079);
not I_23929 (I409733,I409716);
nand I_23930 (I409750,I409733,I409546);
not I_23931 (I409466,I409750);
nor I_23932 (I409469,I409750,I409665);
nand I_23933 (I409472,I409648,I409733);
nand I_23934 (I409809,I409597,I409733);
nand I_23935 (I409826,I409648,I409809);
DFFARX1 I_23936 (I409826,I2898,I409495,I409475,);
nor I_23937 (I409857,I409597,I409682);
and I_23938 (I409874,I409857,I21079);
nor I_23939 (I409484,I409874,I409716);
nand I_23940 (I409905,I409546,I409874);
nand I_23941 (I409487,I409750,I409905);
nand I_23942 (I409936,I21076,I21079);
nor I_23943 (I409953,I21091,I21064);
not I_23944 (I409970,I21082);
nor I_23945 (I409987,I409970,I21073);
nor I_23946 (I410004,I409953,I409970);
not I_23947 (I410021,I410004);
and I_23948 (I410038,I409987,I410021);
nand I_23949 (I409481,I410038,I409936);
nor I_23950 (I410069,I410021,I409716);
not I_23951 (I410086,I410069);
nor I_23952 (I409463,I409987,I410086);
nor I_23953 (I410117,I410004,I409597);
nand I_23954 (I409478,I410117,I409631);
not I_23955 (I410175,I2905);
not I_23956 (I410192,I334743);
nand I_23957 (I410209,I334746,I334734);
and I_23958 (I410226,I410209,I334743);
nand I_23959 (I410243,I410209,I410192);
and I_23960 (I410260,I410243,I334752);
nand I_23961 (I410277,I410260,I334740);
or I_23962 (I410294,I334731,I334746);
nor I_23963 (I410311,I410294,I334734);
not I_23964 (I410328,I410311);
and I_23965 (I410345,I410277,I410328);
not I_23966 (I410362,I334743);
nor I_23967 (I410379,I410362,I334737);
nand I_23968 (I410396,I410379,I334749);
not I_23969 (I410413,I410396);
nand I_23970 (I410430,I410413,I410226);
not I_23971 (I410146,I410430);
nor I_23972 (I410149,I410430,I410345);
nand I_23973 (I410152,I410328,I410413);
nand I_23974 (I410489,I410277,I410413);
nand I_23975 (I410506,I410328,I410489);
DFFARX1 I_23976 (I410506,I2898,I410175,I410155,);
nor I_23977 (I410537,I410277,I410362);
and I_23978 (I410554,I410537,I334749);
nor I_23979 (I410164,I410554,I410396);
nand I_23980 (I410585,I410226,I410554);
nand I_23981 (I410167,I410430,I410585);
nand I_23982 (I410616,I334743,I334749);
nor I_23983 (I410633,I334731,I334740);
not I_23984 (I410650,I334755);
nor I_23985 (I410667,I410650,I334737);
nor I_23986 (I410684,I410633,I410650);
not I_23987 (I410701,I410684);
and I_23988 (I410718,I410667,I410701);
nand I_23989 (I410161,I410718,I410616);
nor I_23990 (I410749,I410701,I410396);
not I_23991 (I410766,I410749);
nor I_23992 (I410143,I410667,I410766);
nor I_23993 (I410797,I410684,I410277);
nand I_23994 (I410158,I410797,I410311);
not I_23995 (I410864,I2905);
nand I_23996 (I410881,I341883,I341877);
and I_23997 (I410898,I410881,I341895);
DFFARX1 I_23998 (I410898,I2898,I410864,I410924,);
not I_23999 (I410932,I410924);
nor I_24000 (I410949,I341880,I341877);
not I_24001 (I410966,I341892);
nand I_24002 (I410983,I341886,I341874);
nand I_24003 (I411000,I410983,I410966);
nand I_24004 (I411017,I410983,I341892);
not I_24005 (I411034,I411017);
and I_24006 (I411051,I411000,I341871);
and I_24007 (I411068,I411051,I341889);
or I_24008 (I411085,I341880,I341877);
nor I_24009 (I411102,I411085,I341886);
nor I_24010 (I411119,I411034,I411102);
not I_24011 (I411136,I411102);
nor I_24012 (I411153,I411136,I410949);
nor I_24013 (I410856,I411102,I411068);
nand I_24014 (I411184,I341871,I341874);
nor I_24015 (I411201,I411184,I341883);
not I_24016 (I411218,I411201);
nor I_24017 (I410823,I411068,I411218);
nor I_24018 (I410826,I411218,I411119);
nand I_24019 (I411263,I410932,I411218);
nor I_24020 (I410835,I411153,I411263);
nor I_24021 (I410847,I411201,I411034);
not I_24022 (I411308,I411184);
nand I_24023 (I411325,I411308,I410949);
not I_24024 (I410829,I411325);
nor I_24025 (I410832,I410924,I411325);
and I_24026 (I411370,I411068,I411308);
nor I_24027 (I411387,I411201,I411370);
nor I_24028 (I410838,I411387,I411370);
not I_24029 (I411418,I411387);
nand I_24030 (I411435,I411068,I411418);
nor I_24031 (I410841,I410932,I411435);
nor I_24032 (I411466,I411068,I411308);
DFFARX1 I_24033 (I411466,I2898,I410864,I410844,);
nand I_24034 (I410853,I411017,I411184);
nand I_24035 (I410850,I411184,I411136);
not I_24036 (I411561,I2905);
nand I_24037 (I411578,I198794,I198800);
and I_24038 (I411595,I411578,I198788);
DFFARX1 I_24039 (I411595,I2898,I411561,I411621,);
not I_24040 (I411629,I411621);
nor I_24041 (I411646,I198788,I198800);
not I_24042 (I411663,I198782);
nand I_24043 (I411680,I198791,I198785);
nand I_24044 (I411697,I411680,I411663);
nand I_24045 (I411714,I411680,I198782);
not I_24046 (I411731,I411714);
and I_24047 (I411748,I411697,I198794);
and I_24048 (I411765,I411748,I198797);
or I_24049 (I411782,I198797,I198782);
nor I_24050 (I411799,I411782,I198803);
nor I_24051 (I411816,I411731,I411799);
not I_24052 (I411833,I411799);
nor I_24053 (I411850,I411833,I411646);
nor I_24054 (I411553,I411799,I411765);
nand I_24055 (I411881,I198806,I198791);
nor I_24056 (I411898,I411881,I198785);
not I_24057 (I411915,I411898);
nor I_24058 (I411520,I411765,I411915);
nor I_24059 (I411523,I411915,I411816);
nand I_24060 (I411960,I411629,I411915);
nor I_24061 (I411532,I411850,I411960);
nor I_24062 (I411544,I411898,I411731);
not I_24063 (I412005,I411881);
nand I_24064 (I412022,I412005,I411646);
not I_24065 (I411526,I412022);
nor I_24066 (I411529,I411621,I412022);
and I_24067 (I412067,I411765,I412005);
nor I_24068 (I412084,I411898,I412067);
nor I_24069 (I411535,I412084,I412067);
not I_24070 (I412115,I412084);
nand I_24071 (I412132,I411765,I412115);
nor I_24072 (I411538,I411629,I412132);
nor I_24073 (I412163,I411765,I412005);
DFFARX1 I_24074 (I412163,I2898,I411561,I411541,);
nand I_24075 (I411550,I411714,I411881);
nand I_24076 (I411547,I411881,I411833);
not I_24077 (I412258,I2905);
nand I_24078 (I412275,I57440,I57425);
and I_24079 (I412292,I412275,I57419);
DFFARX1 I_24080 (I412292,I2898,I412258,I412318,);
not I_24081 (I412326,I412318);
nor I_24082 (I412343,I57422,I57425);
not I_24083 (I412360,I57410);
nand I_24084 (I412377,I57410,I57431);
nand I_24085 (I412394,I412377,I412360);
nand I_24086 (I412411,I412377,I57410);
not I_24087 (I412428,I412411);
and I_24088 (I412445,I412394,I57413);
and I_24089 (I412462,I412445,I57434);
or I_24090 (I412479,I57413,I57428);
nor I_24091 (I412496,I412479,I57446);
nor I_24092 (I412513,I412428,I412496);
not I_24093 (I412530,I412496);
nor I_24094 (I412547,I412530,I412343);
nor I_24095 (I412250,I412496,I412462);
nand I_24096 (I412578,I57437,I57443);
nor I_24097 (I412595,I412578,I57416);
not I_24098 (I412612,I412595);
nor I_24099 (I412217,I412462,I412612);
nor I_24100 (I412220,I412612,I412513);
nand I_24101 (I412657,I412326,I412612);
nor I_24102 (I412229,I412547,I412657);
nor I_24103 (I412241,I412595,I412428);
not I_24104 (I412702,I412578);
nand I_24105 (I412719,I412702,I412343);
not I_24106 (I412223,I412719);
nor I_24107 (I412226,I412318,I412719);
and I_24108 (I412764,I412462,I412702);
nor I_24109 (I412781,I412595,I412764);
nor I_24110 (I412232,I412781,I412764);
not I_24111 (I412812,I412781);
nand I_24112 (I412829,I412462,I412812);
nor I_24113 (I412235,I412326,I412829);
nor I_24114 (I412860,I412462,I412702);
DFFARX1 I_24115 (I412860,I2898,I412258,I412238,);
nand I_24116 (I412247,I412411,I412578);
nand I_24117 (I412244,I412578,I412530);
not I_24118 (I412955,I2905);
nand I_24119 (I412972,I320789,I320801);
and I_24120 (I412989,I412972,I320798);
DFFARX1 I_24121 (I412989,I2898,I412955,I413015,);
not I_24122 (I413023,I413015);
nor I_24123 (I413040,I320780,I320801);
not I_24124 (I413057,I320780);
nand I_24125 (I413074,I320774,I320777);
nand I_24126 (I413091,I413074,I413057);
nand I_24127 (I413108,I413074,I320780);
not I_24128 (I413125,I413108);
and I_24129 (I413142,I413091,I320783);
and I_24130 (I413159,I413142,I320792);
or I_24131 (I413176,I320774,I320804);
nor I_24132 (I413193,I413176,I320777);
nor I_24133 (I413210,I413125,I413193);
not I_24134 (I413227,I413193);
nor I_24135 (I413244,I413227,I413040);
nor I_24136 (I412947,I413193,I413159);
nand I_24137 (I413275,I320795,I320786);
nor I_24138 (I413292,I413275,I320783);
not I_24139 (I413309,I413292);
nor I_24140 (I412914,I413159,I413309);
nor I_24141 (I412917,I413309,I413210);
nand I_24142 (I413354,I413023,I413309);
nor I_24143 (I412926,I413244,I413354);
nor I_24144 (I412938,I413292,I413125);
not I_24145 (I413399,I413275);
nand I_24146 (I413416,I413399,I413040);
not I_24147 (I412920,I413416);
nor I_24148 (I412923,I413015,I413416);
and I_24149 (I413461,I413159,I413399);
nor I_24150 (I413478,I413292,I413461);
nor I_24151 (I412929,I413478,I413461);
not I_24152 (I413509,I413478);
nand I_24153 (I413526,I413159,I413509);
nor I_24154 (I412932,I413023,I413526);
nor I_24155 (I413557,I413159,I413399);
DFFARX1 I_24156 (I413557,I2898,I412955,I412935,);
nand I_24157 (I412944,I413108,I413275);
nand I_24158 (I412941,I413275,I413227);
not I_24159 (I413652,I2905);
nand I_24160 (I413669,I293011,I293023);
and I_24161 (I413686,I413669,I293020);
DFFARX1 I_24162 (I413686,I2898,I413652,I413712,);
not I_24163 (I413720,I413712);
nor I_24164 (I413737,I293002,I293023);
not I_24165 (I413754,I293002);
nand I_24166 (I413771,I292996,I292999);
nand I_24167 (I413788,I413771,I413754);
nand I_24168 (I413805,I413771,I293002);
not I_24169 (I413822,I413805);
and I_24170 (I413839,I413788,I293005);
and I_24171 (I413856,I413839,I293014);
or I_24172 (I413873,I292996,I293026);
nor I_24173 (I413890,I413873,I292999);
nor I_24174 (I413907,I413822,I413890);
not I_24175 (I413924,I413890);
nor I_24176 (I413941,I413924,I413737);
nor I_24177 (I413644,I413890,I413856);
nand I_24178 (I413972,I293017,I293008);
nor I_24179 (I413989,I413972,I293005);
not I_24180 (I414006,I413989);
nor I_24181 (I413611,I413856,I414006);
nor I_24182 (I413614,I414006,I413907);
nand I_24183 (I414051,I413720,I414006);
nor I_24184 (I413623,I413941,I414051);
nor I_24185 (I413635,I413989,I413822);
not I_24186 (I414096,I413972);
nand I_24187 (I414113,I414096,I413737);
not I_24188 (I413617,I414113);
nor I_24189 (I413620,I413712,I414113);
and I_24190 (I414158,I413856,I414096);
nor I_24191 (I414175,I413989,I414158);
nor I_24192 (I413626,I414175,I414158);
not I_24193 (I414206,I414175);
nand I_24194 (I414223,I413856,I414206);
nor I_24195 (I413629,I413720,I414223);
nor I_24196 (I414254,I413856,I414096);
DFFARX1 I_24197 (I414254,I2898,I413652,I413632,);
nand I_24198 (I413641,I413805,I413972);
nand I_24199 (I413638,I413972,I413924);
not I_24200 (I414349,I2905);
nand I_24201 (I414366,I312748,I312760);
and I_24202 (I414383,I414366,I312757);
DFFARX1 I_24203 (I414383,I2898,I414349,I414409,);
not I_24204 (I414417,I414409);
nor I_24205 (I414434,I312739,I312760);
not I_24206 (I414451,I312739);
nand I_24207 (I414468,I312733,I312736);
nand I_24208 (I414485,I414468,I414451);
nand I_24209 (I414502,I414468,I312739);
not I_24210 (I414519,I414502);
and I_24211 (I414536,I414485,I312742);
and I_24212 (I414553,I414536,I312751);
or I_24213 (I414570,I312733,I312763);
nor I_24214 (I414587,I414570,I312736);
nor I_24215 (I414604,I414519,I414587);
not I_24216 (I414621,I414587);
nor I_24217 (I414638,I414621,I414434);
nor I_24218 (I414341,I414587,I414553);
nand I_24219 (I414669,I312754,I312745);
nor I_24220 (I414686,I414669,I312742);
not I_24221 (I414703,I414686);
nor I_24222 (I414308,I414553,I414703);
nor I_24223 (I414311,I414703,I414604);
nand I_24224 (I414748,I414417,I414703);
nor I_24225 (I414320,I414638,I414748);
nor I_24226 (I414332,I414686,I414519);
not I_24227 (I414793,I414669);
nand I_24228 (I414810,I414793,I414434);
not I_24229 (I414314,I414810);
nor I_24230 (I414317,I414409,I414810);
and I_24231 (I414855,I414553,I414793);
nor I_24232 (I414872,I414686,I414855);
nor I_24233 (I414323,I414872,I414855);
not I_24234 (I414903,I414872);
nand I_24235 (I414920,I414553,I414903);
nor I_24236 (I414326,I414417,I414920);
nor I_24237 (I414951,I414553,I414793);
DFFARX1 I_24238 (I414951,I2898,I414349,I414329,);
nand I_24239 (I414338,I414502,I414669);
nand I_24240 (I414335,I414669,I414621);
not I_24241 (I415046,I2905);
nand I_24242 (I415063,I200188,I200194);
and I_24243 (I415080,I415063,I200182);
DFFARX1 I_24244 (I415080,I2898,I415046,I415106,);
not I_24245 (I415114,I415106);
nor I_24246 (I415131,I200182,I200194);
not I_24247 (I415148,I200176);
nand I_24248 (I415165,I200185,I200179);
nand I_24249 (I415182,I415165,I415148);
nand I_24250 (I415199,I415165,I200176);
not I_24251 (I415216,I415199);
and I_24252 (I415233,I415182,I200188);
and I_24253 (I415250,I415233,I200191);
or I_24254 (I415267,I200191,I200176);
nor I_24255 (I415284,I415267,I200197);
nor I_24256 (I415301,I415216,I415284);
not I_24257 (I415318,I415284);
nor I_24258 (I415335,I415318,I415131);
nor I_24259 (I415038,I415284,I415250);
nand I_24260 (I415366,I200200,I200185);
nor I_24261 (I415383,I415366,I200179);
not I_24262 (I415400,I415383);
nor I_24263 (I415005,I415250,I415400);
nor I_24264 (I415008,I415400,I415301);
nand I_24265 (I415445,I415114,I415400);
nor I_24266 (I415017,I415335,I415445);
nor I_24267 (I415029,I415383,I415216);
not I_24268 (I415490,I415366);
nand I_24269 (I415507,I415490,I415131);
not I_24270 (I415011,I415507);
nor I_24271 (I415014,I415106,I415507);
and I_24272 (I415552,I415250,I415490);
nor I_24273 (I415569,I415383,I415552);
nor I_24274 (I415020,I415569,I415552);
not I_24275 (I415600,I415569);
nand I_24276 (I415617,I415250,I415600);
nor I_24277 (I415023,I415114,I415617);
nor I_24278 (I415648,I415250,I415490);
DFFARX1 I_24279 (I415648,I2898,I415046,I415026,);
nand I_24280 (I415035,I415199,I415366);
nand I_24281 (I415032,I415366,I415318);
not I_24282 (I415743,I2905);
nand I_24283 (I415760,I347833,I347827);
and I_24284 (I415777,I415760,I347845);
DFFARX1 I_24285 (I415777,I2898,I415743,I415803,);
not I_24286 (I415811,I415803);
nor I_24287 (I415828,I347830,I347827);
not I_24288 (I415845,I347842);
nand I_24289 (I415862,I347836,I347824);
nand I_24290 (I415879,I415862,I415845);
nand I_24291 (I415896,I415862,I347842);
not I_24292 (I415913,I415896);
and I_24293 (I415930,I415879,I347821);
and I_24294 (I415947,I415930,I347839);
or I_24295 (I415964,I347830,I347827);
nor I_24296 (I415981,I415964,I347836);
nor I_24297 (I415998,I415913,I415981);
not I_24298 (I416015,I415981);
nor I_24299 (I416032,I416015,I415828);
nor I_24300 (I415735,I415981,I415947);
nand I_24301 (I416063,I347821,I347824);
nor I_24302 (I416080,I416063,I347833);
not I_24303 (I416097,I416080);
nor I_24304 (I415702,I415947,I416097);
nor I_24305 (I415705,I416097,I415998);
nand I_24306 (I416142,I415811,I416097);
nor I_24307 (I415714,I416032,I416142);
nor I_24308 (I415726,I416080,I415913);
not I_24309 (I416187,I416063);
nand I_24310 (I416204,I416187,I415828);
not I_24311 (I415708,I416204);
nor I_24312 (I415711,I415803,I416204);
and I_24313 (I416249,I415947,I416187);
nor I_24314 (I416266,I416080,I416249);
nor I_24315 (I415717,I416266,I416249);
not I_24316 (I416297,I416266);
nand I_24317 (I416314,I415947,I416297);
nor I_24318 (I415720,I415811,I416314);
nor I_24319 (I416345,I415947,I416187);
DFFARX1 I_24320 (I416345,I2898,I415743,I415723,);
nand I_24321 (I415732,I415896,I416063);
nand I_24322 (I415729,I416063,I416015);
not I_24323 (I416440,I2905);
nand I_24324 (I416457,I346048,I346042);
and I_24325 (I416474,I416457,I346060);
DFFARX1 I_24326 (I416474,I2898,I416440,I416500,);
not I_24327 (I416508,I416500);
nor I_24328 (I416525,I346045,I346042);
not I_24329 (I416542,I346057);
nand I_24330 (I416559,I346051,I346039);
nand I_24331 (I416576,I416559,I416542);
nand I_24332 (I416593,I416559,I346057);
not I_24333 (I416610,I416593);
and I_24334 (I416627,I416576,I346036);
and I_24335 (I416644,I416627,I346054);
or I_24336 (I416661,I346045,I346042);
nor I_24337 (I416678,I416661,I346051);
nor I_24338 (I416695,I416610,I416678);
not I_24339 (I416712,I416678);
nor I_24340 (I416729,I416712,I416525);
nor I_24341 (I416432,I416678,I416644);
nand I_24342 (I416760,I346036,I346039);
nor I_24343 (I416777,I416760,I346048);
not I_24344 (I416794,I416777);
nor I_24345 (I416399,I416644,I416794);
nor I_24346 (I416402,I416794,I416695);
nand I_24347 (I416839,I416508,I416794);
nor I_24348 (I416411,I416729,I416839);
nor I_24349 (I416423,I416777,I416610);
not I_24350 (I416884,I416760);
nand I_24351 (I416901,I416884,I416525);
not I_24352 (I416405,I416901);
nor I_24353 (I416408,I416500,I416901);
and I_24354 (I416946,I416644,I416884);
nor I_24355 (I416963,I416777,I416946);
nor I_24356 (I416414,I416963,I416946);
not I_24357 (I416994,I416963);
nand I_24358 (I417011,I416644,I416994);
nor I_24359 (I416417,I416508,I417011);
nor I_24360 (I417042,I416644,I416884);
DFFARX1 I_24361 (I417042,I2898,I416440,I416420,);
nand I_24362 (I416429,I416593,I416760);
nand I_24363 (I416426,I416760,I416712);
not I_24364 (I417137,I2905);
nand I_24365 (I417154,I48056,I48041);
and I_24366 (I417171,I417154,I48035);
DFFARX1 I_24367 (I417171,I2898,I417137,I417197,);
not I_24368 (I417205,I417197);
nor I_24369 (I417222,I48038,I48041);
not I_24370 (I417239,I48026);
nand I_24371 (I417256,I48026,I48047);
nand I_24372 (I417273,I417256,I417239);
nand I_24373 (I417290,I417256,I48026);
not I_24374 (I417307,I417290);
and I_24375 (I417324,I417273,I48029);
and I_24376 (I417341,I417324,I48050);
or I_24377 (I417358,I48029,I48044);
nor I_24378 (I417375,I417358,I48062);
nor I_24379 (I417392,I417307,I417375);
not I_24380 (I417409,I417375);
nor I_24381 (I417426,I417409,I417222);
nor I_24382 (I417129,I417375,I417341);
nand I_24383 (I417457,I48053,I48059);
nor I_24384 (I417474,I417457,I48032);
not I_24385 (I417491,I417474);
nor I_24386 (I417096,I417341,I417491);
nor I_24387 (I417099,I417491,I417392);
nand I_24388 (I417536,I417205,I417491);
nor I_24389 (I417108,I417426,I417536);
nor I_24390 (I417120,I417474,I417307);
not I_24391 (I417581,I417457);
nand I_24392 (I417598,I417581,I417222);
not I_24393 (I417102,I417598);
nor I_24394 (I417105,I417197,I417598);
and I_24395 (I417643,I417341,I417581);
nor I_24396 (I417660,I417474,I417643);
nor I_24397 (I417111,I417660,I417643);
not I_24398 (I417691,I417660);
nand I_24399 (I417708,I417341,I417691);
nor I_24400 (I417114,I417205,I417708);
nor I_24401 (I417739,I417341,I417581);
DFFARX1 I_24402 (I417739,I2898,I417137,I417117,);
nand I_24403 (I417126,I417290,I417457);
nand I_24404 (I417123,I417457,I417409);
not I_24405 (I417834,I2905);
nand I_24406 (I417851,I2920,I2929);
and I_24407 (I417868,I417851,I2917);
DFFARX1 I_24408 (I417868,I2898,I417834,I417894,);
not I_24409 (I417902,I417894);
nor I_24410 (I417919,I2926,I2929);
not I_24411 (I417936,I2917);
nand I_24412 (I417953,I2908,I2914);
nand I_24413 (I417970,I417953,I417936);
nand I_24414 (I417987,I417953,I2917);
not I_24415 (I418004,I417987);
and I_24416 (I418021,I417970,I2911);
and I_24417 (I418038,I418021,I2908);
or I_24418 (I418055,I2911,I2932);
nor I_24419 (I418072,I418055,I2938);
nor I_24420 (I418089,I418004,I418072);
not I_24421 (I418106,I418072);
nor I_24422 (I418123,I418106,I417919);
nor I_24423 (I417826,I418072,I418038);
nand I_24424 (I418154,I2923,I2914);
nor I_24425 (I418171,I418154,I2935);
not I_24426 (I418188,I418171);
nor I_24427 (I417793,I418038,I418188);
nor I_24428 (I417796,I418188,I418089);
nand I_24429 (I418233,I417902,I418188);
nor I_24430 (I417805,I418123,I418233);
nor I_24431 (I417817,I418171,I418004);
not I_24432 (I418278,I418154);
nand I_24433 (I418295,I418278,I417919);
not I_24434 (I417799,I418295);
nor I_24435 (I417802,I417894,I418295);
and I_24436 (I418340,I418038,I418278);
nor I_24437 (I418357,I418171,I418340);
nor I_24438 (I417808,I418357,I418340);
not I_24439 (I418388,I418357);
nand I_24440 (I418405,I418038,I418388);
nor I_24441 (I417811,I417902,I418405);
nor I_24442 (I418436,I418038,I418278);
DFFARX1 I_24443 (I418436,I2898,I417834,I417814,);
nand I_24444 (I417823,I417987,I418154);
nand I_24445 (I417820,I418154,I418106);
not I_24446 (I418531,I2905);
nand I_24447 (I418548,I305438,I305450);
and I_24448 (I418565,I418548,I305447);
DFFARX1 I_24449 (I418565,I2898,I418531,I418591,);
not I_24450 (I418599,I418591);
nor I_24451 (I418616,I305429,I305450);
not I_24452 (I418633,I305429);
nand I_24453 (I418650,I305423,I305426);
nand I_24454 (I418667,I418650,I418633);
nand I_24455 (I418684,I418650,I305429);
not I_24456 (I418701,I418684);
and I_24457 (I418718,I418667,I305432);
and I_24458 (I418735,I418718,I305441);
or I_24459 (I418752,I305423,I305453);
nor I_24460 (I418769,I418752,I305426);
nor I_24461 (I418786,I418701,I418769);
not I_24462 (I418803,I418769);
nor I_24463 (I418820,I418803,I418616);
nor I_24464 (I418523,I418769,I418735);
nand I_24465 (I418851,I305444,I305435);
nor I_24466 (I418868,I418851,I305432);
not I_24467 (I418885,I418868);
nor I_24468 (I418490,I418735,I418885);
nor I_24469 (I418493,I418885,I418786);
nand I_24470 (I418930,I418599,I418885);
nor I_24471 (I418502,I418820,I418930);
nor I_24472 (I418514,I418868,I418701);
not I_24473 (I418975,I418851);
nand I_24474 (I418992,I418975,I418616);
not I_24475 (I418496,I418992);
nor I_24476 (I418499,I418591,I418992);
and I_24477 (I419037,I418735,I418975);
nor I_24478 (I419054,I418868,I419037);
nor I_24479 (I418505,I419054,I419037);
not I_24480 (I419085,I419054);
nand I_24481 (I419102,I418735,I419085);
nor I_24482 (I418508,I418599,I419102);
nor I_24483 (I419133,I418735,I418975);
DFFARX1 I_24484 (I419133,I2898,I418531,I418511,);
nand I_24485 (I418520,I418684,I418851);
nand I_24486 (I418517,I418851,I418803);
not I_24487 (I419228,I2905);
nand I_24488 (I419245,I105954,I105951);
and I_24489 (I419262,I419245,I105957);
DFFARX1 I_24490 (I419262,I2898,I419228,I419288,);
not I_24491 (I419296,I419288);
nor I_24492 (I419313,I105951,I105951);
not I_24493 (I419330,I105963);
nand I_24494 (I419347,I105975,I105960);
nand I_24495 (I419364,I419347,I419330);
nand I_24496 (I419381,I419347,I105963);
not I_24497 (I419398,I419381);
and I_24498 (I419415,I419364,I105948);
and I_24499 (I419432,I419415,I105945);
or I_24500 (I419449,I105948,I105972);
nor I_24501 (I419466,I419449,I105969);
nor I_24502 (I419483,I419398,I419466);
not I_24503 (I419500,I419466);
nor I_24504 (I419517,I419500,I419313);
nor I_24505 (I419220,I419466,I419432);
nand I_24506 (I419548,I105978,I105945);
nor I_24507 (I419565,I419548,I105966);
not I_24508 (I419582,I419565);
nor I_24509 (I419187,I419432,I419582);
nor I_24510 (I419190,I419582,I419483);
nand I_24511 (I419627,I419296,I419582);
nor I_24512 (I419199,I419517,I419627);
nor I_24513 (I419211,I419565,I419398);
not I_24514 (I419672,I419548);
nand I_24515 (I419689,I419672,I419313);
not I_24516 (I419193,I419689);
nor I_24517 (I419196,I419288,I419689);
and I_24518 (I419734,I419432,I419672);
nor I_24519 (I419751,I419565,I419734);
nor I_24520 (I419202,I419751,I419734);
not I_24521 (I419782,I419751);
nand I_24522 (I419799,I419432,I419782);
nor I_24523 (I419205,I419296,I419799);
nor I_24524 (I419830,I419432,I419672);
DFFARX1 I_24525 (I419830,I2898,I419228,I419208,);
nand I_24526 (I419217,I419381,I419548);
nand I_24527 (I419214,I419548,I419500);
not I_24528 (I419925,I2905);
nand I_24529 (I419942,I303976,I303988);
and I_24530 (I419959,I419942,I303985);
DFFARX1 I_24531 (I419959,I2898,I419925,I419985,);
not I_24532 (I419993,I419985);
nor I_24533 (I420010,I303967,I303988);
not I_24534 (I420027,I303967);
nand I_24535 (I420044,I303961,I303964);
nand I_24536 (I420061,I420044,I420027);
nand I_24537 (I420078,I420044,I303967);
not I_24538 (I420095,I420078);
and I_24539 (I420112,I420061,I303970);
and I_24540 (I420129,I420112,I303979);
or I_24541 (I420146,I303961,I303991);
nor I_24542 (I420163,I420146,I303964);
nor I_24543 (I420180,I420095,I420163);
not I_24544 (I420197,I420163);
nor I_24545 (I420214,I420197,I420010);
nor I_24546 (I419917,I420163,I420129);
nand I_24547 (I420245,I303982,I303973);
nor I_24548 (I420262,I420245,I303970);
not I_24549 (I420279,I420262);
nor I_24550 (I419884,I420129,I420279);
nor I_24551 (I419887,I420279,I420180);
nand I_24552 (I420324,I419993,I420279);
nor I_24553 (I419896,I420214,I420324);
nor I_24554 (I419908,I420262,I420095);
not I_24555 (I420369,I420245);
nand I_24556 (I420386,I420369,I420010);
not I_24557 (I419890,I420386);
nor I_24558 (I419893,I419985,I420386);
and I_24559 (I420431,I420129,I420369);
nor I_24560 (I420448,I420262,I420431);
nor I_24561 (I419899,I420448,I420431);
not I_24562 (I420479,I420448);
nand I_24563 (I420496,I420129,I420479);
nor I_24564 (I419902,I419993,I420496);
nor I_24565 (I420527,I420129,I420369);
DFFARX1 I_24566 (I420527,I2898,I419925,I419905,);
nand I_24567 (I419914,I420078,I420245);
nand I_24568 (I419911,I420245,I420197);
not I_24569 (I420622,I2905);
nand I_24570 (I420639,I175600,I175627);
and I_24571 (I420656,I420639,I175594);
DFFARX1 I_24572 (I420656,I2898,I420622,I420682,);
not I_24573 (I420690,I420682);
nor I_24574 (I420707,I175609,I175627);
not I_24575 (I420724,I175615);
nand I_24576 (I420741,I175597,I175624);
nand I_24577 (I420758,I420741,I420724);
nand I_24578 (I420775,I420741,I175615);
not I_24579 (I420792,I420775);
and I_24580 (I420809,I420758,I175612);
and I_24581 (I420826,I420809,I175606);
or I_24582 (I420843,I175597,I175603);
nor I_24583 (I420860,I420843,I175600);
nor I_24584 (I420877,I420792,I420860);
not I_24585 (I420894,I420860);
nor I_24586 (I420911,I420894,I420707);
nor I_24587 (I420614,I420860,I420826);
nand I_24588 (I420942,I175621,I175618);
nor I_24589 (I420959,I420942,I175594);
not I_24590 (I420976,I420959);
nor I_24591 (I420581,I420826,I420976);
nor I_24592 (I420584,I420976,I420877);
nand I_24593 (I421021,I420690,I420976);
nor I_24594 (I420593,I420911,I421021);
nor I_24595 (I420605,I420959,I420792);
not I_24596 (I421066,I420942);
nand I_24597 (I421083,I421066,I420707);
not I_24598 (I420587,I421083);
nor I_24599 (I420590,I420682,I421083);
and I_24600 (I421128,I420826,I421066);
nor I_24601 (I421145,I420959,I421128);
nor I_24602 (I420596,I421145,I421128);
not I_24603 (I421176,I421145);
nand I_24604 (I421193,I420826,I421176);
nor I_24605 (I420599,I420690,I421193);
nor I_24606 (I421224,I420826,I421066);
DFFARX1 I_24607 (I421224,I2898,I420622,I420602,);
nand I_24608 (I420611,I420775,I420942);
nand I_24609 (I420608,I420942,I420894);
not I_24610 (I421319,I2905);
nand I_24611 (I421336,I384868,I384853);
and I_24612 (I421353,I421336,I384859);
DFFARX1 I_24613 (I421353,I2898,I421319,I421379,);
not I_24614 (I421387,I421379);
nor I_24615 (I421404,I384850,I384853);
not I_24616 (I421421,I384880);
nand I_24617 (I421438,I384853,I384877);
nand I_24618 (I421455,I421438,I421421);
nand I_24619 (I421472,I421438,I384880);
not I_24620 (I421489,I421472);
and I_24621 (I421506,I421455,I384850);
and I_24622 (I421523,I421506,I384847);
or I_24623 (I421540,I384862,I384847);
nor I_24624 (I421557,I421540,I384874);
nor I_24625 (I421574,I421489,I421557);
not I_24626 (I421591,I421557);
nor I_24627 (I421608,I421591,I421404);
nor I_24628 (I421311,I421557,I421523);
nand I_24629 (I421639,I384871,I384865);
nor I_24630 (I421656,I421639,I384856);
not I_24631 (I421673,I421656);
nor I_24632 (I421278,I421523,I421673);
nor I_24633 (I421281,I421673,I421574);
nand I_24634 (I421718,I421387,I421673);
nor I_24635 (I421290,I421608,I421718);
nor I_24636 (I421302,I421656,I421489);
not I_24637 (I421763,I421639);
nand I_24638 (I421780,I421763,I421404);
not I_24639 (I421284,I421780);
nor I_24640 (I421287,I421379,I421780);
and I_24641 (I421825,I421523,I421763);
nor I_24642 (I421842,I421656,I421825);
nor I_24643 (I421293,I421842,I421825);
not I_24644 (I421873,I421842);
nand I_24645 (I421890,I421523,I421873);
nor I_24646 (I421296,I421387,I421890);
nor I_24647 (I421921,I421523,I421763);
DFFARX1 I_24648 (I421921,I2898,I421319,I421299,);
nand I_24649 (I421308,I421472,I421639);
nand I_24650 (I421305,I421639,I421591);
not I_24651 (I422016,I2905);
nand I_24652 (I422033,I12100,I12109);
and I_24653 (I422050,I422033,I12097);
DFFARX1 I_24654 (I422050,I2898,I422016,I422076,);
not I_24655 (I422084,I422076);
nor I_24656 (I422101,I12106,I12109);
not I_24657 (I422118,I12097);
nand I_24658 (I422135,I12088,I12094);
nand I_24659 (I422152,I422135,I422118);
nand I_24660 (I422169,I422135,I12097);
not I_24661 (I422186,I422169);
and I_24662 (I422203,I422152,I12091);
and I_24663 (I422220,I422203,I12088);
or I_24664 (I422237,I12091,I12112);
nor I_24665 (I422254,I422237,I12118);
nor I_24666 (I422271,I422186,I422254);
not I_24667 (I422288,I422254);
nor I_24668 (I422305,I422288,I422101);
nor I_24669 (I422008,I422254,I422220);
nand I_24670 (I422336,I12103,I12094);
nor I_24671 (I422353,I422336,I12115);
not I_24672 (I422370,I422353);
nor I_24673 (I421975,I422220,I422370);
nor I_24674 (I421978,I422370,I422271);
nand I_24675 (I422415,I422084,I422370);
nor I_24676 (I421987,I422305,I422415);
nor I_24677 (I421999,I422353,I422186);
not I_24678 (I422460,I422336);
nand I_24679 (I422477,I422460,I422101);
not I_24680 (I421981,I422477);
nor I_24681 (I421984,I422076,I422477);
and I_24682 (I422522,I422220,I422460);
nor I_24683 (I422539,I422353,I422522);
nor I_24684 (I421990,I422539,I422522);
not I_24685 (I422570,I422539);
nand I_24686 (I422587,I422220,I422570);
nor I_24687 (I421993,I422084,I422587);
nor I_24688 (I422618,I422220,I422460);
DFFARX1 I_24689 (I422618,I2898,I422016,I421996,);
nand I_24690 (I422005,I422169,I422336);
nand I_24691 (I422002,I422336,I422288);
not I_24692 (I422713,I2905);
nand I_24693 (I422730,I379054,I379039);
and I_24694 (I422747,I422730,I379045);
DFFARX1 I_24695 (I422747,I2898,I422713,I422773,);
not I_24696 (I422781,I422773);
nor I_24697 (I422798,I379036,I379039);
not I_24698 (I422815,I379066);
nand I_24699 (I422832,I379039,I379063);
nand I_24700 (I422849,I422832,I422815);
nand I_24701 (I422866,I422832,I379066);
not I_24702 (I422883,I422866);
and I_24703 (I422900,I422849,I379036);
and I_24704 (I422917,I422900,I379033);
or I_24705 (I422934,I379048,I379033);
nor I_24706 (I422951,I422934,I379060);
nor I_24707 (I422968,I422883,I422951);
not I_24708 (I422985,I422951);
nor I_24709 (I423002,I422985,I422798);
nor I_24710 (I422705,I422951,I422917);
nand I_24711 (I423033,I379057,I379051);
nor I_24712 (I423050,I423033,I379042);
not I_24713 (I423067,I423050);
nor I_24714 (I422672,I422917,I423067);
nor I_24715 (I422675,I423067,I422968);
nand I_24716 (I423112,I422781,I423067);
nor I_24717 (I422684,I423002,I423112);
nor I_24718 (I422696,I423050,I422883);
not I_24719 (I423157,I423033);
nand I_24720 (I423174,I423157,I422798);
not I_24721 (I422678,I423174);
nor I_24722 (I422681,I422773,I423174);
and I_24723 (I423219,I422917,I423157);
nor I_24724 (I423236,I423050,I423219);
nor I_24725 (I422687,I423236,I423219);
not I_24726 (I423267,I423236);
nand I_24727 (I423284,I422917,I423267);
nor I_24728 (I422690,I422781,I423284);
nor I_24729 (I423315,I422917,I423157);
DFFARX1 I_24730 (I423315,I2898,I422713,I422693,);
nand I_24731 (I422702,I422866,I423033);
nand I_24732 (I422699,I423033,I422985);
not I_24733 (I423410,I2905);
nand I_24734 (I423427,I205956,I205974);
and I_24735 (I423444,I423427,I205965);
DFFARX1 I_24736 (I423444,I2898,I423410,I423470,);
not I_24737 (I423478,I423470);
nor I_24738 (I423495,I205968,I205974);
not I_24739 (I423512,I205965);
nand I_24740 (I423529,I205959,I205983);
nand I_24741 (I423546,I423529,I423512);
nand I_24742 (I423563,I423529,I205965);
not I_24743 (I423580,I423563);
and I_24744 (I423597,I423546,I205968);
and I_24745 (I423614,I423597,I205962);
or I_24746 (I423631,I205962,I205956);
nor I_24747 (I423648,I423631,I205977);
nor I_24748 (I423665,I423580,I423648);
not I_24749 (I423682,I423648);
nor I_24750 (I423699,I423682,I423495);
nor I_24751 (I423402,I423648,I423614);
nand I_24752 (I423730,I205980,I205971);
nor I_24753 (I423747,I423730,I205959);
not I_24754 (I423764,I423747);
nor I_24755 (I423369,I423614,I423764);
nor I_24756 (I423372,I423764,I423665);
nand I_24757 (I423809,I423478,I423764);
nor I_24758 (I423381,I423699,I423809);
nor I_24759 (I423393,I423747,I423580);
not I_24760 (I423854,I423730);
nand I_24761 (I423871,I423854,I423495);
not I_24762 (I423375,I423871);
nor I_24763 (I423378,I423470,I423871);
and I_24764 (I423916,I423614,I423854);
nor I_24765 (I423933,I423747,I423916);
nor I_24766 (I423384,I423933,I423916);
not I_24767 (I423964,I423933);
nand I_24768 (I423981,I423614,I423964);
nor I_24769 (I423387,I423478,I423981);
nor I_24770 (I424012,I423614,I423854);
DFFARX1 I_24771 (I424012,I2898,I423410,I423390,);
nand I_24772 (I423399,I423563,I423730);
nand I_24773 (I423396,I423730,I423682);
not I_24774 (I424107,I2905);
nand I_24775 (I424124,I374532,I374517);
and I_24776 (I424141,I424124,I374523);
DFFARX1 I_24777 (I424141,I2898,I424107,I424167,);
not I_24778 (I424175,I424167);
nor I_24779 (I424192,I374514,I374517);
not I_24780 (I424209,I374544);
nand I_24781 (I424226,I374517,I374541);
nand I_24782 (I424243,I424226,I424209);
nand I_24783 (I424260,I424226,I374544);
not I_24784 (I424277,I424260);
and I_24785 (I424294,I424243,I374514);
and I_24786 (I424311,I424294,I374511);
or I_24787 (I424328,I374526,I374511);
nor I_24788 (I424345,I424328,I374538);
nor I_24789 (I424362,I424277,I424345);
not I_24790 (I424379,I424345);
nor I_24791 (I424396,I424379,I424192);
nor I_24792 (I424099,I424345,I424311);
nand I_24793 (I424427,I374535,I374529);
nor I_24794 (I424444,I424427,I374520);
not I_24795 (I424461,I424444);
nor I_24796 (I424066,I424311,I424461);
nor I_24797 (I424069,I424461,I424362);
nand I_24798 (I424506,I424175,I424461);
nor I_24799 (I424078,I424396,I424506);
nor I_24800 (I424090,I424444,I424277);
not I_24801 (I424551,I424427);
nand I_24802 (I424568,I424551,I424192);
not I_24803 (I424072,I424568);
nor I_24804 (I424075,I424167,I424568);
and I_24805 (I424613,I424311,I424551);
nor I_24806 (I424630,I424444,I424613);
nor I_24807 (I424081,I424630,I424613);
not I_24808 (I424661,I424630);
nand I_24809 (I424678,I424311,I424661);
nor I_24810 (I424084,I424175,I424678);
nor I_24811 (I424709,I424311,I424551);
DFFARX1 I_24812 (I424709,I2898,I424107,I424087,);
nand I_24813 (I424096,I424260,I424427);
nand I_24814 (I424093,I424427,I424379);
not I_24815 (I424804,I2905);
nand I_24816 (I424821,I394558,I394543);
and I_24817 (I424838,I424821,I394549);
DFFARX1 I_24818 (I424838,I2898,I424804,I424864,);
not I_24819 (I424872,I424864);
nor I_24820 (I424889,I394540,I394543);
not I_24821 (I424906,I394570);
nand I_24822 (I424923,I394543,I394567);
nand I_24823 (I424940,I424923,I424906);
nand I_24824 (I424957,I424923,I394570);
not I_24825 (I424974,I424957);
and I_24826 (I424991,I424940,I394540);
and I_24827 (I425008,I424991,I394537);
or I_24828 (I425025,I394552,I394537);
nor I_24829 (I425042,I425025,I394564);
nor I_24830 (I425059,I424974,I425042);
not I_24831 (I425076,I425042);
nor I_24832 (I425093,I425076,I424889);
nor I_24833 (I424796,I425042,I425008);
nand I_24834 (I425124,I394561,I394555);
nor I_24835 (I425141,I425124,I394546);
not I_24836 (I425158,I425141);
nor I_24837 (I424763,I425008,I425158);
nor I_24838 (I424766,I425158,I425059);
nand I_24839 (I425203,I424872,I425158);
nor I_24840 (I424775,I425093,I425203);
nor I_24841 (I424787,I425141,I424974);
not I_24842 (I425248,I425124);
nand I_24843 (I425265,I425248,I424889);
not I_24844 (I424769,I425265);
nor I_24845 (I424772,I424864,I425265);
and I_24846 (I425310,I425008,I425248);
nor I_24847 (I425327,I425141,I425310);
nor I_24848 (I424778,I425327,I425310);
not I_24849 (I425358,I425327);
nand I_24850 (I425375,I425008,I425358);
nor I_24851 (I424781,I424872,I425375);
nor I_24852 (I425406,I425008,I425248);
DFFARX1 I_24853 (I425406,I2898,I424804,I424784,);
nand I_24854 (I424793,I424957,I425124);
nand I_24855 (I424790,I425124,I425076);
not I_24856 (I425501,I2905);
nand I_24857 (I425518,I371948,I371933);
and I_24858 (I425535,I425518,I371939);
DFFARX1 I_24859 (I425535,I2898,I425501,I425561,);
not I_24860 (I425569,I425561);
nor I_24861 (I425586,I371930,I371933);
not I_24862 (I425603,I371960);
nand I_24863 (I425620,I371933,I371957);
nand I_24864 (I425637,I425620,I425603);
nand I_24865 (I425654,I425620,I371960);
not I_24866 (I425671,I425654);
and I_24867 (I425688,I425637,I371930);
and I_24868 (I425705,I425688,I371927);
or I_24869 (I425722,I371942,I371927);
nor I_24870 (I425739,I425722,I371954);
nor I_24871 (I425756,I425671,I425739);
not I_24872 (I425773,I425739);
nor I_24873 (I425790,I425773,I425586);
nor I_24874 (I425493,I425739,I425705);
nand I_24875 (I425821,I371951,I371945);
nor I_24876 (I425838,I425821,I371936);
not I_24877 (I425855,I425838);
nor I_24878 (I425460,I425705,I425855);
nor I_24879 (I425463,I425855,I425756);
nand I_24880 (I425900,I425569,I425855);
nor I_24881 (I425472,I425790,I425900);
nor I_24882 (I425484,I425838,I425671);
not I_24883 (I425945,I425821);
nand I_24884 (I425962,I425945,I425586);
not I_24885 (I425466,I425962);
nor I_24886 (I425469,I425561,I425962);
and I_24887 (I426007,I425705,I425945);
nor I_24888 (I426024,I425838,I426007);
nor I_24889 (I425475,I426024,I426007);
not I_24890 (I426055,I426024);
nand I_24891 (I426072,I425705,I426055);
nor I_24892 (I425478,I425569,I426072);
nor I_24893 (I426103,I425705,I425945);
DFFARX1 I_24894 (I426103,I2898,I425501,I425481,);
nand I_24895 (I425490,I425654,I425821);
nand I_24896 (I425487,I425821,I425773);
not I_24897 (I426198,I2905);
nand I_24898 (I426215,I117905,I117902);
and I_24899 (I426232,I426215,I117908);
DFFARX1 I_24900 (I426232,I2898,I426198,I426258,);
not I_24901 (I426266,I426258);
nor I_24902 (I426283,I117902,I117902);
not I_24903 (I426300,I117914);
nand I_24904 (I426317,I117926,I117911);
nand I_24905 (I426334,I426317,I426300);
nand I_24906 (I426351,I426317,I117914);
not I_24907 (I426368,I426351);
and I_24908 (I426385,I426334,I117899);
and I_24909 (I426402,I426385,I117896);
or I_24910 (I426419,I117899,I117923);
nor I_24911 (I426436,I426419,I117920);
nor I_24912 (I426453,I426368,I426436);
not I_24913 (I426470,I426436);
nor I_24914 (I426487,I426470,I426283);
nor I_24915 (I426190,I426436,I426402);
nand I_24916 (I426518,I117929,I117896);
nor I_24917 (I426535,I426518,I117917);
not I_24918 (I426552,I426535);
nor I_24919 (I426157,I426402,I426552);
nor I_24920 (I426160,I426552,I426453);
nand I_24921 (I426597,I426266,I426552);
nor I_24922 (I426169,I426487,I426597);
nor I_24923 (I426181,I426535,I426368);
not I_24924 (I426642,I426518);
nand I_24925 (I426659,I426642,I426283);
not I_24926 (I426163,I426659);
nor I_24927 (I426166,I426258,I426659);
and I_24928 (I426704,I426402,I426642);
nor I_24929 (I426721,I426535,I426704);
nor I_24930 (I426172,I426721,I426704);
not I_24931 (I426752,I426721);
nand I_24932 (I426769,I426402,I426752);
nor I_24933 (I426175,I426266,I426769);
nor I_24934 (I426800,I426402,I426642);
DFFARX1 I_24935 (I426800,I2898,I426198,I426178,);
nand I_24936 (I426187,I426351,I426518);
nand I_24937 (I426184,I426518,I426470);
not I_24938 (I426895,I2905);
nand I_24939 (I426912,I3532,I3541);
and I_24940 (I426929,I426912,I3529);
DFFARX1 I_24941 (I426929,I2898,I426895,I426955,);
not I_24942 (I426963,I426955);
nor I_24943 (I426980,I3538,I3541);
not I_24944 (I426997,I3529);
nand I_24945 (I427014,I3520,I3526);
nand I_24946 (I427031,I427014,I426997);
nand I_24947 (I427048,I427014,I3529);
not I_24948 (I427065,I427048);
and I_24949 (I427082,I427031,I3523);
and I_24950 (I427099,I427082,I3520);
or I_24951 (I427116,I3523,I3544);
nor I_24952 (I427133,I427116,I3550);
nor I_24953 (I427150,I427065,I427133);
not I_24954 (I427167,I427133);
nor I_24955 (I427184,I427167,I426980);
nor I_24956 (I426887,I427133,I427099);
nand I_24957 (I427215,I3535,I3526);
nor I_24958 (I427232,I427215,I3547);
not I_24959 (I427249,I427232);
nor I_24960 (I426854,I427099,I427249);
nor I_24961 (I426857,I427249,I427150);
nand I_24962 (I427294,I426963,I427249);
nor I_24963 (I426866,I427184,I427294);
nor I_24964 (I426878,I427232,I427065);
not I_24965 (I427339,I427215);
nand I_24966 (I427356,I427339,I426980);
not I_24967 (I426860,I427356);
nor I_24968 (I426863,I426955,I427356);
and I_24969 (I427401,I427099,I427339);
nor I_24970 (I427418,I427232,I427401);
nor I_24971 (I426869,I427418,I427401);
not I_24972 (I427449,I427418);
nand I_24973 (I427466,I427099,I427449);
nor I_24974 (I426872,I426963,I427466);
nor I_24975 (I427497,I427099,I427339);
DFFARX1 I_24976 (I427497,I2898,I426895,I426875,);
nand I_24977 (I426884,I427048,I427215);
nand I_24978 (I426881,I427215,I427167);
not I_24979 (I427592,I2905);
nand I_24980 (I427609,I364904,I364916);
and I_24981 (I427626,I427609,I364922);
DFFARX1 I_24982 (I427626,I2898,I427592,I427652,);
not I_24983 (I427660,I427652);
nor I_24984 (I427677,I364898,I364916);
not I_24985 (I427694,I364907);
nand I_24986 (I427711,I364913,I364889);
nand I_24987 (I427728,I427711,I427694);
nand I_24988 (I427745,I427711,I364907);
not I_24989 (I427762,I427745);
and I_24990 (I427779,I427728,I364910);
and I_24991 (I427796,I427779,I364892);
or I_24992 (I427813,I364892,I364919);
nor I_24993 (I427830,I427813,I364895);
nor I_24994 (I427847,I427762,I427830);
not I_24995 (I427864,I427830);
nor I_24996 (I427881,I427864,I427677);
nor I_24997 (I427584,I427830,I427796);
nand I_24998 (I427912,I364895,I364889);
nor I_24999 (I427929,I427912,I364901);
not I_25000 (I427946,I427929);
nor I_25001 (I427551,I427796,I427946);
nor I_25002 (I427554,I427946,I427847);
nand I_25003 (I427991,I427660,I427946);
nor I_25004 (I427563,I427881,I427991);
nor I_25005 (I427575,I427929,I427762);
not I_25006 (I428036,I427912);
nand I_25007 (I428053,I428036,I427677);
not I_25008 (I427557,I428053);
nor I_25009 (I427560,I427652,I428053);
and I_25010 (I428098,I427796,I428036);
nor I_25011 (I428115,I427929,I428098);
nor I_25012 (I427566,I428115,I428098);
not I_25013 (I428146,I428115);
nand I_25014 (I428163,I427796,I428146);
nor I_25015 (I427569,I427660,I428163);
nor I_25016 (I428194,I427796,I428036);
DFFARX1 I_25017 (I428194,I2898,I427592,I427572,);
nand I_25018 (I427581,I427745,I427912);
nand I_25019 (I427578,I427912,I427864);
not I_25020 (I428289,I2905);
nand I_25021 (I428306,I224656,I224674);
and I_25022 (I428323,I428306,I224665);
DFFARX1 I_25023 (I428323,I2898,I428289,I428349,);
not I_25024 (I428357,I428349);
nor I_25025 (I428374,I224668,I224674);
not I_25026 (I428391,I224665);
nand I_25027 (I428408,I224659,I224683);
nand I_25028 (I428425,I428408,I428391);
nand I_25029 (I428442,I428408,I224665);
not I_25030 (I428459,I428442);
and I_25031 (I428476,I428425,I224668);
and I_25032 (I428493,I428476,I224662);
or I_25033 (I428510,I224662,I224656);
nor I_25034 (I428527,I428510,I224677);
nor I_25035 (I428544,I428459,I428527);
not I_25036 (I428561,I428527);
nor I_25037 (I428578,I428561,I428374);
nor I_25038 (I428281,I428527,I428493);
nand I_25039 (I428609,I224680,I224671);
nor I_25040 (I428626,I428609,I224659);
not I_25041 (I428643,I428626);
nor I_25042 (I428248,I428493,I428643);
nor I_25043 (I428251,I428643,I428544);
nand I_25044 (I428688,I428357,I428643);
nor I_25045 (I428260,I428578,I428688);
nor I_25046 (I428272,I428626,I428459);
not I_25047 (I428733,I428609);
nand I_25048 (I428750,I428733,I428374);
not I_25049 (I428254,I428750);
nor I_25050 (I428257,I428349,I428750);
and I_25051 (I428795,I428493,I428733);
nor I_25052 (I428812,I428626,I428795);
nor I_25053 (I428263,I428812,I428795);
not I_25054 (I428843,I428812);
nand I_25055 (I428860,I428493,I428843);
nor I_25056 (I428266,I428357,I428860);
nor I_25057 (I428891,I428493,I428733);
DFFARX1 I_25058 (I428891,I2898,I428289,I428269,);
nand I_25059 (I428278,I428442,I428609);
nand I_25060 (I428275,I428609,I428561);
not I_25061 (I428986,I2905);
nand I_25062 (I429003,I166760,I166787);
and I_25063 (I429020,I429003,I166754);
DFFARX1 I_25064 (I429020,I2898,I428986,I429046,);
not I_25065 (I429054,I429046);
nor I_25066 (I429071,I166769,I166787);
not I_25067 (I429088,I166775);
nand I_25068 (I429105,I166757,I166784);
nand I_25069 (I429122,I429105,I429088);
nand I_25070 (I429139,I429105,I166775);
not I_25071 (I429156,I429139);
and I_25072 (I429173,I429122,I166772);
and I_25073 (I429190,I429173,I166766);
or I_25074 (I429207,I166757,I166763);
nor I_25075 (I429224,I429207,I166760);
nor I_25076 (I429241,I429156,I429224);
not I_25077 (I429258,I429224);
nor I_25078 (I429275,I429258,I429071);
nor I_25079 (I428978,I429224,I429190);
nand I_25080 (I429306,I166781,I166778);
nor I_25081 (I429323,I429306,I166754);
not I_25082 (I429340,I429323);
nor I_25083 (I428945,I429190,I429340);
nor I_25084 (I428948,I429340,I429241);
nand I_25085 (I429385,I429054,I429340);
nor I_25086 (I428957,I429275,I429385);
nor I_25087 (I428969,I429323,I429156);
not I_25088 (I429430,I429306);
nand I_25089 (I429447,I429430,I429071);
not I_25090 (I428951,I429447);
nor I_25091 (I428954,I429046,I429447);
and I_25092 (I429492,I429190,I429430);
nor I_25093 (I429509,I429323,I429492);
nor I_25094 (I428960,I429509,I429492);
not I_25095 (I429540,I429509);
nand I_25096 (I429557,I429190,I429540);
nor I_25097 (I428963,I429054,I429557);
nor I_25098 (I429588,I429190,I429430);
DFFARX1 I_25099 (I429588,I2898,I428986,I428966,);
nand I_25100 (I428975,I429139,I429306);
nand I_25101 (I428972,I429306,I429258);
not I_25102 (I429683,I2905);
nand I_25103 (I429700,I186248,I186254);
and I_25104 (I429717,I429700,I186242);
DFFARX1 I_25105 (I429717,I2898,I429683,I429743,);
not I_25106 (I429751,I429743);
nor I_25107 (I429768,I186242,I186254);
not I_25108 (I429785,I186236);
nand I_25109 (I429802,I186245,I186239);
nand I_25110 (I429819,I429802,I429785);
nand I_25111 (I429836,I429802,I186236);
not I_25112 (I429853,I429836);
and I_25113 (I429870,I429819,I186248);
and I_25114 (I429887,I429870,I186251);
or I_25115 (I429904,I186251,I186236);
nor I_25116 (I429921,I429904,I186257);
nor I_25117 (I429938,I429853,I429921);
not I_25118 (I429955,I429921);
nor I_25119 (I429972,I429955,I429768);
nor I_25120 (I429675,I429921,I429887);
nand I_25121 (I430003,I186260,I186245);
nor I_25122 (I430020,I430003,I186239);
not I_25123 (I430037,I430020);
nor I_25124 (I429642,I429887,I430037);
nor I_25125 (I429645,I430037,I429938);
nand I_25126 (I430082,I429751,I430037);
nor I_25127 (I429654,I429972,I430082);
nor I_25128 (I429666,I430020,I429853);
not I_25129 (I430127,I430003);
nand I_25130 (I430144,I430127,I429768);
not I_25131 (I429648,I430144);
nor I_25132 (I429651,I429743,I430144);
and I_25133 (I430189,I429887,I430127);
nor I_25134 (I430206,I430020,I430189);
nor I_25135 (I429657,I430206,I430189);
not I_25136 (I430237,I430206);
nand I_25137 (I430254,I429887,I430237);
nor I_25138 (I429660,I429751,I430254);
nor I_25139 (I430285,I429887,I430127);
DFFARX1 I_25140 (I430285,I2898,I429683,I429663,);
nand I_25141 (I429672,I429836,I430003);
nand I_25142 (I429669,I430003,I429955);
not I_25143 (I430380,I2905);
nand I_25144 (I430397,I134259,I134256);
and I_25145 (I430414,I430397,I134262);
DFFARX1 I_25146 (I430414,I2898,I430380,I430440,);
not I_25147 (I430448,I430440);
nor I_25148 (I430465,I134256,I134256);
not I_25149 (I430482,I134268);
nand I_25150 (I430499,I134280,I134265);
nand I_25151 (I430516,I430499,I430482);
nand I_25152 (I430533,I430499,I134268);
not I_25153 (I430550,I430533);
and I_25154 (I430567,I430516,I134253);
and I_25155 (I430584,I430567,I134250);
or I_25156 (I430601,I134253,I134277);
nor I_25157 (I430618,I430601,I134274);
nor I_25158 (I430635,I430550,I430618);
not I_25159 (I430652,I430618);
nor I_25160 (I430669,I430652,I430465);
nor I_25161 (I430372,I430618,I430584);
nand I_25162 (I430700,I134283,I134250);
nor I_25163 (I430717,I430700,I134271);
not I_25164 (I430734,I430717);
nor I_25165 (I430339,I430584,I430734);
nor I_25166 (I430342,I430734,I430635);
nand I_25167 (I430779,I430448,I430734);
nor I_25168 (I430351,I430669,I430779);
nor I_25169 (I430363,I430717,I430550);
not I_25170 (I430824,I430700);
nand I_25171 (I430841,I430824,I430465);
not I_25172 (I430345,I430841);
nor I_25173 (I430348,I430440,I430841);
and I_25174 (I430886,I430584,I430824);
nor I_25175 (I430903,I430717,I430886);
nor I_25176 (I430354,I430903,I430886);
not I_25177 (I430934,I430903);
nand I_25178 (I430951,I430584,I430934);
nor I_25179 (I430357,I430448,I430951);
nor I_25180 (I430982,I430584,I430824);
DFFARX1 I_25181 (I430982,I2898,I430380,I430360,);
nand I_25182 (I430369,I430533,I430700);
nand I_25183 (I430366,I430700,I430652);
not I_25184 (I431077,I2905);
nand I_25185 (I431094,I117276,I117273);
and I_25186 (I431111,I431094,I117279);
DFFARX1 I_25187 (I431111,I2898,I431077,I431137,);
not I_25188 (I431145,I431137);
nor I_25189 (I431162,I117273,I117273);
not I_25190 (I431179,I117285);
nand I_25191 (I431196,I117297,I117282);
nand I_25192 (I431213,I431196,I431179);
nand I_25193 (I431230,I431196,I117285);
not I_25194 (I431247,I431230);
and I_25195 (I431264,I431213,I117270);
and I_25196 (I431281,I431264,I117267);
or I_25197 (I431298,I117270,I117294);
nor I_25198 (I431315,I431298,I117291);
nor I_25199 (I431332,I431247,I431315);
not I_25200 (I431349,I431315);
nor I_25201 (I431366,I431349,I431162);
nor I_25202 (I431069,I431315,I431281);
nand I_25203 (I431397,I117300,I117267);
nor I_25204 (I431414,I431397,I117288);
not I_25205 (I431431,I431414);
nor I_25206 (I431036,I431281,I431431);
nor I_25207 (I431039,I431431,I431332);
nand I_25208 (I431476,I431145,I431431);
nor I_25209 (I431048,I431366,I431476);
nor I_25210 (I431060,I431414,I431247);
not I_25211 (I431521,I431397);
nand I_25212 (I431538,I431521,I431162);
not I_25213 (I431042,I431538);
nor I_25214 (I431045,I431137,I431538);
and I_25215 (I431583,I431281,I431521);
nor I_25216 (I431600,I431414,I431583);
nor I_25217 (I431051,I431600,I431583);
not I_25218 (I431631,I431600);
nand I_25219 (I431648,I431281,I431631);
nor I_25220 (I431054,I431145,I431648);
nor I_25221 (I431679,I431281,I431521);
DFFARX1 I_25222 (I431679,I2898,I431077,I431057,);
nand I_25223 (I431066,I431230,I431397);
nand I_25224 (I431063,I431397,I431349);
not I_25225 (I431774,I2905);
nand I_25226 (I431791,I138662,I138659);
and I_25227 (I431808,I431791,I138665);
DFFARX1 I_25228 (I431808,I2898,I431774,I431834,);
not I_25229 (I431842,I431834);
nor I_25230 (I431859,I138659,I138659);
not I_25231 (I431876,I138671);
nand I_25232 (I431893,I138683,I138668);
nand I_25233 (I431910,I431893,I431876);
nand I_25234 (I431927,I431893,I138671);
not I_25235 (I431944,I431927);
and I_25236 (I431961,I431910,I138656);
and I_25237 (I431978,I431961,I138653);
or I_25238 (I431995,I138656,I138680);
nor I_25239 (I432012,I431995,I138677);
nor I_25240 (I432029,I431944,I432012);
not I_25241 (I432046,I432012);
nor I_25242 (I432063,I432046,I431859);
nor I_25243 (I431766,I432012,I431978);
nand I_25244 (I432094,I138686,I138653);
nor I_25245 (I432111,I432094,I138674);
not I_25246 (I432128,I432111);
nor I_25247 (I431733,I431978,I432128);
nor I_25248 (I431736,I432128,I432029);
nand I_25249 (I432173,I431842,I432128);
nor I_25250 (I431745,I432063,I432173);
nor I_25251 (I431757,I432111,I431944);
not I_25252 (I432218,I432094);
nand I_25253 (I432235,I432218,I431859);
not I_25254 (I431739,I432235);
nor I_25255 (I431742,I431834,I432235);
and I_25256 (I432280,I431978,I432218);
nor I_25257 (I432297,I432111,I432280);
nor I_25258 (I431748,I432297,I432280);
not I_25259 (I432328,I432297);
nand I_25260 (I432345,I431978,I432328);
nor I_25261 (I431751,I431842,I432345);
nor I_25262 (I432376,I431978,I432218);
DFFARX1 I_25263 (I432376,I2898,I431774,I431754,);
nand I_25264 (I431763,I431927,I432094);
nand I_25265 (I431760,I432094,I432046);
not I_25266 (I432471,I2905);
nand I_25267 (I432488,I331768,I331762);
and I_25268 (I432505,I432488,I331780);
DFFARX1 I_25269 (I432505,I2898,I432471,I432531,);
not I_25270 (I432539,I432531);
nor I_25271 (I432556,I331765,I331762);
not I_25272 (I432573,I331777);
nand I_25273 (I432590,I331771,I331759);
nand I_25274 (I432607,I432590,I432573);
nand I_25275 (I432624,I432590,I331777);
not I_25276 (I432641,I432624);
and I_25277 (I432658,I432607,I331756);
and I_25278 (I432675,I432658,I331774);
or I_25279 (I432692,I331765,I331762);
nor I_25280 (I432709,I432692,I331771);
nor I_25281 (I432726,I432641,I432709);
not I_25282 (I432743,I432709);
nor I_25283 (I432760,I432743,I432556);
nor I_25284 (I432463,I432709,I432675);
nand I_25285 (I432791,I331756,I331759);
nor I_25286 (I432808,I432791,I331768);
not I_25287 (I432825,I432808);
nor I_25288 (I432430,I432675,I432825);
nor I_25289 (I432433,I432825,I432726);
nand I_25290 (I432870,I432539,I432825);
nor I_25291 (I432442,I432760,I432870);
nor I_25292 (I432454,I432808,I432641);
not I_25293 (I432915,I432791);
nand I_25294 (I432932,I432915,I432556);
not I_25295 (I432436,I432932);
nor I_25296 (I432439,I432531,I432932);
and I_25297 (I432977,I432675,I432915);
nor I_25298 (I432994,I432808,I432977);
nor I_25299 (I432445,I432994,I432977);
not I_25300 (I433025,I432994);
nand I_25301 (I433042,I432675,I433025);
nor I_25302 (I432448,I432539,I433042);
nor I_25303 (I433073,I432675,I432915);
DFFARX1 I_25304 (I433073,I2898,I432471,I432451,);
nand I_25305 (I432460,I432624,I432791);
nand I_25306 (I432457,I432791,I432743);
not I_25307 (I433168,I2905);
nand I_25308 (I433185,I219420,I219438);
and I_25309 (I433202,I433185,I219429);
DFFARX1 I_25310 (I433202,I2898,I433168,I433228,);
not I_25311 (I433236,I433228);
nor I_25312 (I433253,I219432,I219438);
not I_25313 (I433270,I219429);
nand I_25314 (I433287,I219423,I219447);
nand I_25315 (I433304,I433287,I433270);
nand I_25316 (I433321,I433287,I219429);
not I_25317 (I433338,I433321);
and I_25318 (I433355,I433304,I219432);
and I_25319 (I433372,I433355,I219426);
or I_25320 (I433389,I219426,I219420);
nor I_25321 (I433406,I433389,I219441);
nor I_25322 (I433423,I433338,I433406);
not I_25323 (I433440,I433406);
nor I_25324 (I433457,I433440,I433253);
nor I_25325 (I433160,I433406,I433372);
nand I_25326 (I433488,I219444,I219435);
nor I_25327 (I433505,I433488,I219423);
not I_25328 (I433522,I433505);
nor I_25329 (I433127,I433372,I433522);
nor I_25330 (I433130,I433522,I433423);
nand I_25331 (I433567,I433236,I433522);
nor I_25332 (I433139,I433457,I433567);
nor I_25333 (I433151,I433505,I433338);
not I_25334 (I433612,I433488);
nand I_25335 (I433629,I433612,I433253);
not I_25336 (I433133,I433629);
nor I_25337 (I433136,I433228,I433629);
and I_25338 (I433674,I433372,I433612);
nor I_25339 (I433691,I433505,I433674);
nor I_25340 (I433142,I433691,I433674);
not I_25341 (I433722,I433691);
nand I_25342 (I433739,I433372,I433722);
nor I_25343 (I433145,I433236,I433739);
nor I_25344 (I433770,I433372,I433612);
DFFARX1 I_25345 (I433770,I2898,I433168,I433148,);
nand I_25346 (I433157,I433321,I433488);
nand I_25347 (I433154,I433488,I433440);
not I_25348 (I433865,I2905);
nand I_25349 (I433882,I124824,I124821);
and I_25350 (I433899,I433882,I124827);
DFFARX1 I_25351 (I433899,I2898,I433865,I433925,);
not I_25352 (I433933,I433925);
nor I_25353 (I433950,I124821,I124821);
not I_25354 (I433967,I124833);
nand I_25355 (I433984,I124845,I124830);
nand I_25356 (I434001,I433984,I433967);
nand I_25357 (I434018,I433984,I124833);
not I_25358 (I434035,I434018);
and I_25359 (I434052,I434001,I124818);
and I_25360 (I434069,I434052,I124815);
or I_25361 (I434086,I124818,I124842);
nor I_25362 (I434103,I434086,I124839);
nor I_25363 (I434120,I434035,I434103);
not I_25364 (I434137,I434103);
nor I_25365 (I434154,I434137,I433950);
nor I_25366 (I433857,I434103,I434069);
nand I_25367 (I434185,I124848,I124815);
nor I_25368 (I434202,I434185,I124836);
not I_25369 (I434219,I434202);
nor I_25370 (I433824,I434069,I434219);
nor I_25371 (I433827,I434219,I434120);
nand I_25372 (I434264,I433933,I434219);
nor I_25373 (I433836,I434154,I434264);
nor I_25374 (I433848,I434202,I434035);
not I_25375 (I434309,I434185);
nand I_25376 (I434326,I434309,I433950);
not I_25377 (I433830,I434326);
nor I_25378 (I433833,I433925,I434326);
and I_25379 (I434371,I434069,I434309);
nor I_25380 (I434388,I434202,I434371);
nor I_25381 (I433839,I434388,I434371);
not I_25382 (I434419,I434388);
nand I_25383 (I434436,I434069,I434419);
nor I_25384 (I433842,I433933,I434436);
nor I_25385 (I434467,I434069,I434309);
DFFARX1 I_25386 (I434467,I2898,I433865,I433845,);
nand I_25387 (I433854,I434018,I434185);
nand I_25388 (I433851,I434185,I434137);
not I_25389 (I434562,I2905);
nand I_25390 (I434579,I12712,I12721);
and I_25391 (I434596,I434579,I12709);
DFFARX1 I_25392 (I434596,I2898,I434562,I434622,);
not I_25393 (I434630,I434622);
nor I_25394 (I434647,I12718,I12721);
not I_25395 (I434664,I12709);
nand I_25396 (I434681,I12700,I12706);
nand I_25397 (I434698,I434681,I434664);
nand I_25398 (I434715,I434681,I12709);
not I_25399 (I434732,I434715);
and I_25400 (I434749,I434698,I12703);
and I_25401 (I434766,I434749,I12700);
or I_25402 (I434783,I12703,I12724);
nor I_25403 (I434800,I434783,I12730);
nor I_25404 (I434817,I434732,I434800);
not I_25405 (I434834,I434800);
nor I_25406 (I434851,I434834,I434647);
nor I_25407 (I434554,I434800,I434766);
nand I_25408 (I434882,I12715,I12706);
nor I_25409 (I434899,I434882,I12727);
not I_25410 (I434916,I434899);
nor I_25411 (I434521,I434766,I434916);
nor I_25412 (I434524,I434916,I434817);
nand I_25413 (I434961,I434630,I434916);
nor I_25414 (I434533,I434851,I434961);
nor I_25415 (I434545,I434899,I434732);
not I_25416 (I435006,I434882);
nand I_25417 (I435023,I435006,I434647);
not I_25418 (I434527,I435023);
nor I_25419 (I434530,I434622,I435023);
and I_25420 (I435068,I434766,I435006);
nor I_25421 (I435085,I434899,I435068);
nor I_25422 (I434536,I435085,I435068);
not I_25423 (I435116,I435085);
nand I_25424 (I435133,I434766,I435116);
nor I_25425 (I434539,I434630,I435133);
nor I_25426 (I435164,I434766,I435006);
DFFARX1 I_25427 (I435164,I2898,I434562,I434542,);
nand I_25428 (I434551,I434715,I434882);
nand I_25429 (I434548,I434882,I434834);
not I_25430 (I435259,I2905);
nand I_25431 (I435276,I126711,I126708);
and I_25432 (I435293,I435276,I126714);
DFFARX1 I_25433 (I435293,I2898,I435259,I435319,);
not I_25434 (I435327,I435319);
nor I_25435 (I435344,I126708,I126708);
not I_25436 (I435361,I126720);
nand I_25437 (I435378,I126732,I126717);
nand I_25438 (I435395,I435378,I435361);
nand I_25439 (I435412,I435378,I126720);
not I_25440 (I435429,I435412);
and I_25441 (I435446,I435395,I126705);
and I_25442 (I435463,I435446,I126702);
or I_25443 (I435480,I126705,I126729);
nor I_25444 (I435497,I435480,I126726);
nor I_25445 (I435514,I435429,I435497);
not I_25446 (I435531,I435497);
nor I_25447 (I435548,I435531,I435344);
nor I_25448 (I435251,I435497,I435463);
nand I_25449 (I435579,I126735,I126702);
nor I_25450 (I435596,I435579,I126723);
not I_25451 (I435613,I435596);
nor I_25452 (I435218,I435463,I435613);
nor I_25453 (I435221,I435613,I435514);
nand I_25454 (I435658,I435327,I435613);
nor I_25455 (I435230,I435548,I435658);
nor I_25456 (I435242,I435596,I435429);
not I_25457 (I435703,I435579);
nand I_25458 (I435720,I435703,I435344);
not I_25459 (I435224,I435720);
nor I_25460 (I435227,I435319,I435720);
and I_25461 (I435765,I435463,I435703);
nor I_25462 (I435782,I435596,I435765);
nor I_25463 (I435233,I435782,I435765);
not I_25464 (I435813,I435782);
nand I_25465 (I435830,I435463,I435813);
nor I_25466 (I435236,I435327,I435830);
nor I_25467 (I435861,I435463,I435703);
DFFARX1 I_25468 (I435861,I2898,I435259,I435239,);
nand I_25469 (I435248,I435412,I435579);
nand I_25470 (I435245,I435579,I435531);
not I_25471 (I435956,I2905);
nand I_25472 (I435973,I63865,I63877);
and I_25473 (I435990,I435973,I63853);
DFFARX1 I_25474 (I435990,I2898,I435956,I436016,);
not I_25475 (I436024,I436016);
nor I_25476 (I436041,I63862,I63877);
not I_25477 (I436058,I63862);
nand I_25478 (I436075,I63874,I63880);
nand I_25479 (I436092,I436075,I436058);
nand I_25480 (I436109,I436075,I63862);
not I_25481 (I436126,I436109);
and I_25482 (I436143,I436092,I63853);
and I_25483 (I436160,I436143,I63859);
or I_25484 (I436177,I63859,I63856);
nor I_25485 (I436194,I436177,I63865);
nor I_25486 (I436211,I436126,I436194);
not I_25487 (I436228,I436194);
nor I_25488 (I436245,I436228,I436041);
nor I_25489 (I435948,I436194,I436160);
nand I_25490 (I436276,I63871,I63868);
nor I_25491 (I436293,I436276,I63856);
not I_25492 (I436310,I436293);
nor I_25493 (I435915,I436160,I436310);
nor I_25494 (I435918,I436310,I436211);
nand I_25495 (I436355,I436024,I436310);
nor I_25496 (I435927,I436245,I436355);
nor I_25497 (I435939,I436293,I436126);
not I_25498 (I436400,I436276);
nand I_25499 (I436417,I436400,I436041);
not I_25500 (I435921,I436417);
nor I_25501 (I435924,I436016,I436417);
and I_25502 (I436462,I436160,I436400);
nor I_25503 (I436479,I436293,I436462);
nor I_25504 (I435930,I436479,I436462);
not I_25505 (I436510,I436479);
nand I_25506 (I436527,I436160,I436510);
nor I_25507 (I435933,I436024,I436527);
nor I_25508 (I436558,I436160,I436400);
DFFARX1 I_25509 (I436558,I2898,I435956,I435936,);
nand I_25510 (I435945,I436109,I436276);
nand I_25511 (I435942,I436276,I436228);
not I_25512 (I436653,I2905);
nand I_25513 (I436670,I337718,I337712);
and I_25514 (I436687,I436670,I337730);
DFFARX1 I_25515 (I436687,I2898,I436653,I436713,);
not I_25516 (I436721,I436713);
nor I_25517 (I436738,I337715,I337712);
not I_25518 (I436755,I337727);
nand I_25519 (I436772,I337721,I337709);
nand I_25520 (I436789,I436772,I436755);
nand I_25521 (I436806,I436772,I337727);
not I_25522 (I436823,I436806);
and I_25523 (I436840,I436789,I337706);
and I_25524 (I436857,I436840,I337724);
or I_25525 (I436874,I337715,I337712);
nor I_25526 (I436891,I436874,I337721);
nor I_25527 (I436908,I436823,I436891);
not I_25528 (I436925,I436891);
nor I_25529 (I436942,I436925,I436738);
nor I_25530 (I436645,I436891,I436857);
nand I_25531 (I436973,I337706,I337709);
nor I_25532 (I436990,I436973,I337718);
not I_25533 (I437007,I436990);
nor I_25534 (I436612,I436857,I437007);
nor I_25535 (I436615,I437007,I436908);
nand I_25536 (I437052,I436721,I437007);
nor I_25537 (I436624,I436942,I437052);
nor I_25538 (I436636,I436990,I436823);
not I_25539 (I437097,I436973);
nand I_25540 (I437114,I437097,I436738);
not I_25541 (I436618,I437114);
nor I_25542 (I436621,I436713,I437114);
and I_25543 (I437159,I436857,I437097);
nor I_25544 (I437176,I436990,I437159);
nor I_25545 (I436627,I437176,I437159);
not I_25546 (I437207,I437176);
nand I_25547 (I437224,I436857,I437207);
nor I_25548 (I436630,I436721,I437224);
nor I_25549 (I437255,I436857,I437097);
DFFARX1 I_25550 (I437255,I2898,I436653,I436633,);
nand I_25551 (I436642,I436806,I436973);
nand I_25552 (I436639,I436973,I436925);
not I_25553 (I437350,I2905);
nand I_25554 (I437367,I96573,I96585);
and I_25555 (I437384,I437367,I96561);
DFFARX1 I_25556 (I437384,I2898,I437350,I437410,);
not I_25557 (I437418,I437410);
nor I_25558 (I437435,I96570,I96585);
not I_25559 (I437452,I96570);
nand I_25560 (I437469,I96582,I96588);
nand I_25561 (I437486,I437469,I437452);
nand I_25562 (I437503,I437469,I96570);
not I_25563 (I437520,I437503);
and I_25564 (I437537,I437486,I96561);
and I_25565 (I437554,I437537,I96567);
or I_25566 (I437571,I96567,I96564);
nor I_25567 (I437588,I437571,I96573);
nor I_25568 (I437605,I437520,I437588);
not I_25569 (I437622,I437588);
nor I_25570 (I437639,I437622,I437435);
nor I_25571 (I437342,I437588,I437554);
nand I_25572 (I437670,I96579,I96576);
nor I_25573 (I437687,I437670,I96564);
not I_25574 (I437704,I437687);
nor I_25575 (I437309,I437554,I437704);
nor I_25576 (I437312,I437704,I437605);
nand I_25577 (I437749,I437418,I437704);
nor I_25578 (I437321,I437639,I437749);
nor I_25579 (I437333,I437687,I437520);
not I_25580 (I437794,I437670);
nand I_25581 (I437811,I437794,I437435);
not I_25582 (I437315,I437811);
nor I_25583 (I437318,I437410,I437811);
and I_25584 (I437856,I437554,I437794);
nor I_25585 (I437873,I437687,I437856);
nor I_25586 (I437324,I437873,I437856);
not I_25587 (I437904,I437873);
nand I_25588 (I437921,I437554,I437904);
nor I_25589 (I437327,I437418,I437921);
nor I_25590 (I437952,I437554,I437794);
DFFARX1 I_25591 (I437952,I2898,I437350,I437330,);
nand I_25592 (I437339,I437503,I437670);
nand I_25593 (I437336,I437670,I437622);
not I_25594 (I438047,I2905);
nand I_25595 (I438064,I161320,I161347);
and I_25596 (I438081,I438064,I161314);
DFFARX1 I_25597 (I438081,I2898,I438047,I438107,);
not I_25598 (I438115,I438107);
nor I_25599 (I438132,I161329,I161347);
not I_25600 (I438149,I161335);
nand I_25601 (I438166,I161317,I161344);
nand I_25602 (I438183,I438166,I438149);
nand I_25603 (I438200,I438166,I161335);
not I_25604 (I438217,I438200);
and I_25605 (I438234,I438183,I161332);
and I_25606 (I438251,I438234,I161326);
or I_25607 (I438268,I161317,I161323);
nor I_25608 (I438285,I438268,I161320);
nor I_25609 (I438302,I438217,I438285);
not I_25610 (I438319,I438285);
nor I_25611 (I438336,I438319,I438132);
nor I_25612 (I438039,I438285,I438251);
nand I_25613 (I438367,I161341,I161338);
nor I_25614 (I438384,I438367,I161314);
not I_25615 (I438401,I438384);
nor I_25616 (I438006,I438251,I438401);
nor I_25617 (I438009,I438401,I438302);
nand I_25618 (I438446,I438115,I438401);
nor I_25619 (I438018,I438336,I438446);
nor I_25620 (I438030,I438384,I438217);
not I_25621 (I438491,I438367);
nand I_25622 (I438508,I438491,I438132);
not I_25623 (I438012,I438508);
nor I_25624 (I438015,I438107,I438508);
and I_25625 (I438553,I438251,I438491);
nor I_25626 (I438570,I438384,I438553);
nor I_25627 (I438021,I438570,I438553);
not I_25628 (I438601,I438570);
nand I_25629 (I438618,I438251,I438601);
nor I_25630 (I438024,I438115,I438618);
nor I_25631 (I438649,I438251,I438491);
DFFARX1 I_25632 (I438649,I2898,I438047,I438027,);
nand I_25633 (I438036,I438200,I438367);
nand I_25634 (I438033,I438367,I438319);
not I_25635 (I438744,I2905);
nand I_25636 (I438761,I19636,I19645);
and I_25637 (I438778,I438761,I19639);
DFFARX1 I_25638 (I438778,I2898,I438744,I438804,);
not I_25639 (I438812,I438804);
nor I_25640 (I438829,I19642,I19645);
not I_25641 (I438846,I19636);
nand I_25642 (I438863,I19663,I19648);
nand I_25643 (I438880,I438863,I438846);
nand I_25644 (I438897,I438863,I19636);
not I_25645 (I438914,I438897);
and I_25646 (I438931,I438880,I19651);
and I_25647 (I438948,I438931,I19645);
or I_25648 (I438965,I19642,I19648);
nor I_25649 (I438982,I438965,I19654);
nor I_25650 (I438999,I438914,I438982);
not I_25651 (I439016,I438982);
nor I_25652 (I439033,I439016,I438829);
nor I_25653 (I438736,I438982,I438948);
nand I_25654 (I439064,I19657,I19660);
nor I_25655 (I439081,I439064,I19639);
not I_25656 (I439098,I439081);
nor I_25657 (I438703,I438948,I439098);
nor I_25658 (I438706,I439098,I438999);
nand I_25659 (I439143,I438812,I439098);
nor I_25660 (I438715,I439033,I439143);
nor I_25661 (I438727,I439081,I438914);
not I_25662 (I439188,I439064);
nand I_25663 (I439205,I439188,I438829);
not I_25664 (I438709,I439205);
nor I_25665 (I438712,I438804,I439205);
and I_25666 (I439250,I438948,I439188);
nor I_25667 (I439267,I439081,I439250);
nor I_25668 (I438718,I439267,I439250);
not I_25669 (I439298,I439267);
nand I_25670 (I439315,I438948,I439298);
nor I_25671 (I438721,I438812,I439315);
nor I_25672 (I439346,I438948,I439188);
DFFARX1 I_25673 (I439346,I2898,I438744,I438724,);
nand I_25674 (I438733,I438897,I439064);
nand I_25675 (I438730,I439064,I439016);
not I_25676 (I439441,I2905);
nand I_25677 (I439458,I2427,I1947);
and I_25678 (I439475,I439458,I1915);
DFFARX1 I_25679 (I439475,I2898,I439441,I439501,);
not I_25680 (I439509,I439501);
nor I_25681 (I439526,I2467,I1947);
not I_25682 (I439543,I2875);
nand I_25683 (I439560,I2763,I2579);
nand I_25684 (I439577,I439560,I439543);
nand I_25685 (I439594,I439560,I2875);
not I_25686 (I439611,I439594);
and I_25687 (I439628,I439577,I2587);
and I_25688 (I439645,I439628,I1723);
or I_25689 (I439662,I1867,I1987);
nor I_25690 (I439679,I439662,I2707);
nor I_25691 (I439696,I439611,I439679);
not I_25692 (I439713,I439679);
nor I_25693 (I439730,I439713,I439526);
nor I_25694 (I439433,I439679,I439645);
nand I_25695 (I439761,I2811,I2603);
nor I_25696 (I439778,I439761,I2563);
not I_25697 (I439795,I439778);
nor I_25698 (I439400,I439645,I439795);
nor I_25699 (I439403,I439795,I439696);
nand I_25700 (I439840,I439509,I439795);
nor I_25701 (I439412,I439730,I439840);
nor I_25702 (I439424,I439778,I439611);
not I_25703 (I439885,I439761);
nand I_25704 (I439902,I439885,I439526);
not I_25705 (I439406,I439902);
nor I_25706 (I439409,I439501,I439902);
and I_25707 (I439947,I439645,I439885);
nor I_25708 (I439964,I439778,I439947);
nor I_25709 (I439415,I439964,I439947);
not I_25710 (I439995,I439964);
nand I_25711 (I440012,I439645,I439995);
nor I_25712 (I439418,I439509,I440012);
nor I_25713 (I440043,I439645,I439885);
DFFARX1 I_25714 (I440043,I2898,I439441,I439421,);
nand I_25715 (I439430,I439594,I439761);
nand I_25716 (I439427,I439761,I439713);
not I_25717 (I440138,I2905);
nand I_25718 (I440155,I359733,I359727);
and I_25719 (I440172,I440155,I359745);
DFFARX1 I_25720 (I440172,I2898,I440138,I440198,);
not I_25721 (I440206,I440198);
nor I_25722 (I440223,I359730,I359727);
not I_25723 (I440240,I359742);
nand I_25724 (I440257,I359736,I359724);
nand I_25725 (I440274,I440257,I440240);
nand I_25726 (I440291,I440257,I359742);
not I_25727 (I440308,I440291);
and I_25728 (I440325,I440274,I359721);
and I_25729 (I440342,I440325,I359739);
or I_25730 (I440359,I359730,I359727);
nor I_25731 (I440376,I440359,I359736);
nor I_25732 (I440393,I440308,I440376);
not I_25733 (I440410,I440376);
nor I_25734 (I440427,I440410,I440223);
nor I_25735 (I440130,I440376,I440342);
nand I_25736 (I440458,I359721,I359724);
nor I_25737 (I440475,I440458,I359733);
not I_25738 (I440492,I440475);
nor I_25739 (I440097,I440342,I440492);
nor I_25740 (I440100,I440492,I440393);
nand I_25741 (I440537,I440206,I440492);
nor I_25742 (I440109,I440427,I440537);
nor I_25743 (I440121,I440475,I440308);
not I_25744 (I440582,I440458);
nand I_25745 (I440599,I440582,I440223);
not I_25746 (I440103,I440599);
nor I_25747 (I440106,I440198,I440599);
and I_25748 (I440644,I440342,I440582);
nor I_25749 (I440661,I440475,I440644);
nor I_25750 (I440112,I440661,I440644);
not I_25751 (I440692,I440661);
nand I_25752 (I440709,I440342,I440692);
nor I_25753 (I440115,I440206,I440709);
nor I_25754 (I440740,I440342,I440582);
DFFARX1 I_25755 (I440740,I2898,I440138,I440118,);
nand I_25756 (I440127,I440291,I440458);
nand I_25757 (I440124,I440458,I440410);
not I_25758 (I440835,I2905);
nand I_25759 (I440852,I93428,I93440);
and I_25760 (I440869,I440852,I93416);
DFFARX1 I_25761 (I440869,I2898,I440835,I440895,);
not I_25762 (I440903,I440895);
nor I_25763 (I440920,I93425,I93440);
not I_25764 (I440937,I93425);
nand I_25765 (I440954,I93437,I93443);
nand I_25766 (I440971,I440954,I440937);
nand I_25767 (I440988,I440954,I93425);
not I_25768 (I441005,I440988);
and I_25769 (I441022,I440971,I93416);
and I_25770 (I441039,I441022,I93422);
or I_25771 (I441056,I93422,I93419);
nor I_25772 (I441073,I441056,I93428);
nor I_25773 (I441090,I441005,I441073);
not I_25774 (I441107,I441073);
nor I_25775 (I441124,I441107,I440920);
nor I_25776 (I440827,I441073,I441039);
nand I_25777 (I441155,I93434,I93431);
nor I_25778 (I441172,I441155,I93419);
not I_25779 (I441189,I441172);
nor I_25780 (I440794,I441039,I441189);
nor I_25781 (I440797,I441189,I441090);
nand I_25782 (I441234,I440903,I441189);
nor I_25783 (I440806,I441124,I441234);
nor I_25784 (I440818,I441172,I441005);
not I_25785 (I441279,I441155);
nand I_25786 (I441296,I441279,I440920);
not I_25787 (I440800,I441296);
nor I_25788 (I440803,I440895,I441296);
and I_25789 (I441341,I441039,I441279);
nor I_25790 (I441358,I441172,I441341);
nor I_25791 (I440809,I441358,I441341);
not I_25792 (I441389,I441358);
nand I_25793 (I441406,I441039,I441389);
nor I_25794 (I440812,I440903,I441406);
nor I_25795 (I441437,I441039,I441279);
DFFARX1 I_25796 (I441437,I2898,I440835,I440815,);
nand I_25797 (I440824,I440988,I441155);
nand I_25798 (I440821,I441155,I441107);
not I_25799 (I441532,I2905);
nand I_25800 (I441549,I292280,I292292);
and I_25801 (I441566,I441549,I292289);
DFFARX1 I_25802 (I441566,I2898,I441532,I441592,);
not I_25803 (I441600,I441592);
nor I_25804 (I441617,I292271,I292292);
not I_25805 (I441634,I292271);
nand I_25806 (I441651,I292265,I292268);
nand I_25807 (I441668,I441651,I441634);
nand I_25808 (I441685,I441651,I292271);
not I_25809 (I441702,I441685);
and I_25810 (I441719,I441668,I292274);
and I_25811 (I441736,I441719,I292283);
or I_25812 (I441753,I292265,I292295);
nor I_25813 (I441770,I441753,I292268);
nor I_25814 (I441787,I441702,I441770);
not I_25815 (I441804,I441770);
nor I_25816 (I441821,I441804,I441617);
nor I_25817 (I441524,I441770,I441736);
nand I_25818 (I441852,I292286,I292277);
nor I_25819 (I441869,I441852,I292274);
not I_25820 (I441886,I441869);
nor I_25821 (I441491,I441736,I441886);
nor I_25822 (I441494,I441886,I441787);
nand I_25823 (I441931,I441600,I441886);
nor I_25824 (I441503,I441821,I441931);
nor I_25825 (I441515,I441869,I441702);
not I_25826 (I441976,I441852);
nand I_25827 (I441993,I441976,I441617);
not I_25828 (I441497,I441993);
nor I_25829 (I441500,I441592,I441993);
and I_25830 (I442038,I441736,I441976);
nor I_25831 (I442055,I441869,I442038);
nor I_25832 (I441506,I442055,I442038);
not I_25833 (I442086,I442055);
nand I_25834 (I442103,I441736,I442086);
nor I_25835 (I441509,I441600,I442103);
nor I_25836 (I442134,I441736,I441976);
DFFARX1 I_25837 (I442134,I2898,I441532,I441512,);
nand I_25838 (I441521,I441685,I441852);
nand I_25839 (I441518,I441852,I441804);
not I_25840 (I442229,I2905);
nand I_25841 (I442246,I37486,I37495);
and I_25842 (I442263,I442246,I37489);
DFFARX1 I_25843 (I442263,I2898,I442229,I442289,);
not I_25844 (I442297,I442289);
nor I_25845 (I442314,I37492,I37495);
not I_25846 (I442331,I37486);
nand I_25847 (I442348,I37513,I37498);
nand I_25848 (I442365,I442348,I442331);
nand I_25849 (I442382,I442348,I37486);
not I_25850 (I442399,I442382);
and I_25851 (I442416,I442365,I37501);
and I_25852 (I442433,I442416,I37495);
or I_25853 (I442450,I37492,I37498);
nor I_25854 (I442467,I442450,I37504);
nor I_25855 (I442484,I442399,I442467);
not I_25856 (I442501,I442467);
nor I_25857 (I442518,I442501,I442314);
nor I_25858 (I442221,I442467,I442433);
nand I_25859 (I442549,I37507,I37510);
nor I_25860 (I442566,I442549,I37489);
not I_25861 (I442583,I442566);
nor I_25862 (I442188,I442433,I442583);
nor I_25863 (I442191,I442583,I442484);
nand I_25864 (I442628,I442297,I442583);
nor I_25865 (I442200,I442518,I442628);
nor I_25866 (I442212,I442566,I442399);
not I_25867 (I442673,I442549);
nand I_25868 (I442690,I442673,I442314);
not I_25869 (I442194,I442690);
nor I_25870 (I442197,I442289,I442690);
and I_25871 (I442735,I442433,I442673);
nor I_25872 (I442752,I442566,I442735);
nor I_25873 (I442203,I442752,I442735);
not I_25874 (I442783,I442752);
nand I_25875 (I442800,I442433,I442783);
nor I_25876 (I442206,I442297,I442800);
nor I_25877 (I442831,I442433,I442673);
DFFARX1 I_25878 (I442831,I2898,I442229,I442209,);
nand I_25879 (I442218,I442382,I442549);
nand I_25880 (I442215,I442549,I442501);
not I_25881 (I442926,I2905);
nand I_25882 (I442943,I59462,I59474);
and I_25883 (I442960,I442943,I59450);
DFFARX1 I_25884 (I442960,I2898,I442926,I442986,);
not I_25885 (I442994,I442986);
nor I_25886 (I443011,I59459,I59474);
not I_25887 (I443028,I59459);
nand I_25888 (I443045,I59471,I59477);
nand I_25889 (I443062,I443045,I443028);
nand I_25890 (I443079,I443045,I59459);
not I_25891 (I443096,I443079);
and I_25892 (I443113,I443062,I59450);
and I_25893 (I443130,I443113,I59456);
or I_25894 (I443147,I59456,I59453);
nor I_25895 (I443164,I443147,I59462);
nor I_25896 (I443181,I443096,I443164);
not I_25897 (I443198,I443164);
nor I_25898 (I443215,I443198,I443011);
nor I_25899 (I442918,I443164,I443130);
nand I_25900 (I443246,I59468,I59465);
nor I_25901 (I443263,I443246,I59453);
not I_25902 (I443280,I443263);
nor I_25903 (I442885,I443130,I443280);
nor I_25904 (I442888,I443280,I443181);
nand I_25905 (I443325,I442994,I443280);
nor I_25906 (I442897,I443215,I443325);
nor I_25907 (I442909,I443263,I443096);
not I_25908 (I443370,I443246);
nand I_25909 (I443387,I443370,I443011);
not I_25910 (I442891,I443387);
nor I_25911 (I442894,I442986,I443387);
and I_25912 (I443432,I443130,I443370);
nor I_25913 (I443449,I443263,I443432);
nor I_25914 (I442900,I443449,I443432);
not I_25915 (I443480,I443449);
nand I_25916 (I443497,I443130,I443480);
nor I_25917 (I442903,I442994,I443497);
nor I_25918 (I443528,I443130,I443370);
DFFARX1 I_25919 (I443528,I2898,I442926,I442906,);
nand I_25920 (I442915,I443079,I443246);
nand I_25921 (I442912,I443246,I443198);
not I_25922 (I443623,I2905);
nand I_25923 (I443640,I325223,I325217);
and I_25924 (I443657,I443640,I325235);
DFFARX1 I_25925 (I443657,I2898,I443623,I443683,);
not I_25926 (I443691,I443683);
nor I_25927 (I443708,I325220,I325217);
not I_25928 (I443725,I325232);
nand I_25929 (I443742,I325226,I325214);
nand I_25930 (I443759,I443742,I443725);
nand I_25931 (I443776,I443742,I325232);
not I_25932 (I443793,I443776);
and I_25933 (I443810,I443759,I325211);
and I_25934 (I443827,I443810,I325229);
or I_25935 (I443844,I325220,I325217);
nor I_25936 (I443861,I443844,I325226);
nor I_25937 (I443878,I443793,I443861);
not I_25938 (I443895,I443861);
nor I_25939 (I443912,I443895,I443708);
nor I_25940 (I443615,I443861,I443827);
nand I_25941 (I443943,I325211,I325214);
nor I_25942 (I443960,I443943,I325223);
not I_25943 (I443977,I443960);
nor I_25944 (I443582,I443827,I443977);
nor I_25945 (I443585,I443977,I443878);
nand I_25946 (I444022,I443691,I443977);
nor I_25947 (I443594,I443912,I444022);
nor I_25948 (I443606,I443960,I443793);
not I_25949 (I444067,I443943);
nand I_25950 (I444084,I444067,I443708);
not I_25951 (I443588,I444084);
nor I_25952 (I443591,I443683,I444084);
and I_25953 (I444129,I443827,I444067);
nor I_25954 (I444146,I443960,I444129);
nor I_25955 (I443597,I444146,I444129);
not I_25956 (I444177,I444146);
nand I_25957 (I444194,I443827,I444177);
nor I_25958 (I443600,I443691,I444194);
nor I_25959 (I444225,I443827,I444067);
DFFARX1 I_25960 (I444225,I2898,I443623,I443603,);
nand I_25961 (I443612,I443776,I443943);
nand I_25962 (I443609,I443943,I443895);
not I_25963 (I444320,I2905);
nand I_25964 (I444337,I176960,I176987);
and I_25965 (I444354,I444337,I176954);
DFFARX1 I_25966 (I444354,I2898,I444320,I444380,);
not I_25967 (I444388,I444380);
nor I_25968 (I444405,I176969,I176987);
not I_25969 (I444422,I176975);
nand I_25970 (I444439,I176957,I176984);
nand I_25971 (I444456,I444439,I444422);
nand I_25972 (I444473,I444439,I176975);
not I_25973 (I444490,I444473);
and I_25974 (I444507,I444456,I176972);
and I_25975 (I444524,I444507,I176966);
or I_25976 (I444541,I176957,I176963);
nor I_25977 (I444558,I444541,I176960);
nor I_25978 (I444575,I444490,I444558);
not I_25979 (I444592,I444558);
nor I_25980 (I444609,I444592,I444405);
nor I_25981 (I444312,I444558,I444524);
nand I_25982 (I444640,I176981,I176978);
nor I_25983 (I444657,I444640,I176954);
not I_25984 (I444674,I444657);
nor I_25985 (I444279,I444524,I444674);
nor I_25986 (I444282,I444674,I444575);
nand I_25987 (I444719,I444388,I444674);
nor I_25988 (I444291,I444609,I444719);
nor I_25989 (I444303,I444657,I444490);
not I_25990 (I444764,I444640);
nand I_25991 (I444781,I444764,I444405);
not I_25992 (I444285,I444781);
nor I_25993 (I444288,I444380,I444781);
and I_25994 (I444826,I444524,I444764);
nor I_25995 (I444843,I444657,I444826);
nor I_25996 (I444294,I444843,I444826);
not I_25997 (I444874,I444843);
nand I_25998 (I444891,I444524,I444874);
nor I_25999 (I444297,I444388,I444891);
nor I_26000 (I444922,I444524,I444764);
DFFARX1 I_26001 (I444922,I2898,I444320,I444300,);
nand I_26002 (I444309,I444473,I444640);
nand I_26003 (I444306,I444640,I444592);
not I_26004 (I445017,I2905);
nand I_26005 (I445034,I301052,I301064);
and I_26006 (I445051,I445034,I301061);
DFFARX1 I_26007 (I445051,I2898,I445017,I445077,);
not I_26008 (I445085,I445077);
nor I_26009 (I445102,I301043,I301064);
not I_26010 (I445119,I301043);
nand I_26011 (I445136,I301037,I301040);
nand I_26012 (I445153,I445136,I445119);
nand I_26013 (I445170,I445136,I301043);
not I_26014 (I445187,I445170);
and I_26015 (I445204,I445153,I301046);
and I_26016 (I445221,I445204,I301055);
or I_26017 (I445238,I301037,I301067);
nor I_26018 (I445255,I445238,I301040);
nor I_26019 (I445272,I445187,I445255);
not I_26020 (I445289,I445255);
nor I_26021 (I445306,I445289,I445102);
nor I_26022 (I445009,I445255,I445221);
nand I_26023 (I445337,I301058,I301049);
nor I_26024 (I445354,I445337,I301046);
not I_26025 (I445371,I445354);
nor I_26026 (I444976,I445221,I445371);
nor I_26027 (I444979,I445371,I445272);
nand I_26028 (I445416,I445085,I445371);
nor I_26029 (I444988,I445306,I445416);
nor I_26030 (I445000,I445354,I445187);
not I_26031 (I445461,I445337);
nand I_26032 (I445478,I445461,I445102);
not I_26033 (I444982,I445478);
nor I_26034 (I444985,I445077,I445478);
and I_26035 (I445523,I445221,I445461);
nor I_26036 (I445540,I445354,I445523);
nor I_26037 (I444991,I445540,I445523);
not I_26038 (I445571,I445540);
nand I_26039 (I445588,I445221,I445571);
nor I_26040 (I444994,I445085,I445588);
nor I_26041 (I445619,I445221,I445461);
DFFARX1 I_26042 (I445619,I2898,I445017,I444997,);
nand I_26043 (I445006,I445170,I445337);
nand I_26044 (I445003,I445337,I445289);
not I_26045 (I445714,I2905);
nand I_26046 (I445731,I391328,I391313);
and I_26047 (I445748,I445731,I391319);
DFFARX1 I_26048 (I445748,I2898,I445714,I445774,);
not I_26049 (I445782,I445774);
nor I_26050 (I445799,I391310,I391313);
not I_26051 (I445816,I391340);
nand I_26052 (I445833,I391313,I391337);
nand I_26053 (I445850,I445833,I445816);
nand I_26054 (I445867,I445833,I391340);
not I_26055 (I445884,I445867);
and I_26056 (I445901,I445850,I391310);
and I_26057 (I445918,I445901,I391307);
or I_26058 (I445935,I391322,I391307);
nor I_26059 (I445952,I445935,I391334);
nor I_26060 (I445969,I445884,I445952);
not I_26061 (I445986,I445952);
nor I_26062 (I446003,I445986,I445799);
nor I_26063 (I445706,I445952,I445918);
nand I_26064 (I446034,I391331,I391325);
nor I_26065 (I446051,I446034,I391316);
not I_26066 (I446068,I446051);
nor I_26067 (I445673,I445918,I446068);
nor I_26068 (I445676,I446068,I445969);
nand I_26069 (I446113,I445782,I446068);
nor I_26070 (I445685,I446003,I446113);
nor I_26071 (I445697,I446051,I445884);
not I_26072 (I446158,I446034);
nand I_26073 (I446175,I446158,I445799);
not I_26074 (I445679,I446175);
nor I_26075 (I445682,I445774,I446175);
and I_26076 (I446220,I445918,I446158);
nor I_26077 (I446237,I446051,I446220);
nor I_26078 (I445688,I446237,I446220);
not I_26079 (I446268,I446237);
nand I_26080 (I446285,I445918,I446268);
nor I_26081 (I445691,I445782,I446285);
nor I_26082 (I446316,I445918,I446158);
DFFARX1 I_26083 (I446316,I2898,I445714,I445694,);
nand I_26084 (I445703,I445867,I446034);
nand I_26085 (I445700,I446034,I445986);
endmodule


