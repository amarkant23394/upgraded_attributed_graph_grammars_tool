module test_final(G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4,n_431_0_l_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n4_1_r_4,blif_clk_net_1_r_9,n5_9,G42_1_r_4,);
nor I_1(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_2(n_573_1_r_4,G2_0_l_4,n16_4);
nor I_3(n_549_1_r_4,n22_4,n23_4);
nand I_4(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_5(n19_4,blif_clk_net_1_r_9,n5_9,ACVQN2_3_r_4,);
nor I_6(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_7(n19_4,blif_clk_net_1_r_9,n5_9,ACVQN1_5_r_4,);
not I_8(P6_5_r_4,P6_5_r_internal_4);
or I_9(n_431_0_l_4,IN_8_0_l_4,n26_4);
DFFARX1 I_10(n_431_0_l_4,blif_clk_net_1_r_9,n5_9,G78_0_l_4,);
DFFARX1 I_11(IN_2_5_l_4,blif_clk_net_1_r_9,n5_9,ACVQN1_5_l_4,);
not I_12(n16_4,ACVQN1_5_l_4);
DFFARX1 I_13(IN_1_5_l_4,blif_clk_net_1_r_9,n5_9,n17_internal_4,);
not I_14(n17_4,n17_internal_4);
nor I_15(n4_1_r_4,n30_4,n31_4);
nand I_16(n19_4,G1_0_l_4,n33_4);
DFFARX1 I_17(G78_0_l_4,blif_clk_net_1_r_9,n5_9,n15_internal_4,);
not I_18(n15_4,n15_internal_4);
DFFARX1 I_19(ACVQN1_5_l_4,blif_clk_net_1_r_9,n5_9,P6_5_r_internal_4,);
and I_20(n20_4,IN_11_0_l_4,n16_4);
nor I_21(n21_4,G2_0_l_4,IN_10_0_l_4);
nand I_22(n22_4,G78_0_l_4,n25_4);
nand I_23(n23_4,IN_11_0_l_4,n24_4);
not I_24(n24_4,G2_0_l_4);
not I_25(n25_4,IN_10_0_l_4);
and I_26(n26_4,IN_2_0_l_4,n27_4);
nor I_27(n27_4,IN_4_0_l_4,n28_4);
not I_28(n28_4,G1_0_l_4);
not I_29(n29_4,n30_4);
nand I_30(n30_4,IN_7_0_l_4,n32_4);
nand I_31(n31_4,IN_11_0_l_4,n25_4);
nor I_32(n32_4,G2_0_l_4,n33_4);
not I_33(n33_4,IN_5_0_l_4);
DFFARX1 I_34(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_35(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_36(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_37(n_549_1_r_9,n17_9,n18_9);
or I_38(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_39(n_452_1_r_9,n26_9,n25_9);
nor I_40(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_41(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_42(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_43(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_44(N3_2_l_9,n22_9,n_573_1_r_4);
not I_45(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_46(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_47(n16_9,n27_9);
DFFARX1 I_48(n_569_1_r_4,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_49(n15_9,n26_9);
DFFARX1 I_50(n_573_1_r_4,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_51(n29_9,n29_internal_9);
and I_52(N1_4_l_9,n24_9,n_572_1_r_4);
DFFARX1 I_53(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_54(ACVQN1_5_r_4,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_55(n28_9,n28_internal_9);
nor I_56(n4_1_r_9,n27_9,n26_9);
nor I_57(N3_2_r_9,n15_9,n21_9);
nor I_58(N1_4_r_9,n16_9,n21_9);
nor I_59(n_42_2_l_9,G42_1_r_4,n_572_1_r_4);
not I_60(n17_9,n_452_1_r_9);
nand I_61(n18_9,n27_9,n15_9);
nor I_62(n19_9,n29_9,n20_9);
not I_63(n20_9,P6_5_r_4);
and I_64(n21_9,n23_9,P6_5_r_4);
nand I_65(n22_9,ACVQN2_3_r_4,n_572_1_r_4);
nor I_66(n23_9,n29_9,n28_9);
nand I_67(n24_9,n_549_1_r_4,n_266_and_0_3_r_4);
endmodule


