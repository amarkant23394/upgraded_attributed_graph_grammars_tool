module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_5_r_13,n9_13,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
nor I_34(N1371_0_r_13,n59_13,n61_13);
nor I_35(N1508_0_r_13,n59_13,n60_13);
not I_36(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_37(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_38(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_39(n_102_5_r_13,N1508_0_r_12,N1507_6_r_12);
nand I_40(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_41(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_42(n_572_7_r_13,n40_13,n41_13);
nand I_43(n_573_7_r_13,n37_13,n38_13);
nor I_44(n_549_7_r_13,n46_13,n47_13);
nand I_45(n_569_7_r_13,n37_13,n43_13);
nand I_46(n_452_7_r_13,n52_13,n53_13);
nor I_47(n4_7_l_13,N1371_0_r_12,N1508_6_r_12);
not I_48(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_49(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_50(n33_13,n62_13);
nand I_51(n_431_5_r_13,n54_13,n55_13);
not I_52(n1_13,n52_13);
nor I_53(n34_13,n35_13,n36_13);
nor I_54(n35_13,n42_13,N1371_0_r_12);
nand I_55(n36_13,n50_13,n58_13);
nand I_56(n37_13,n44_13,n45_13);
or I_57(n38_13,n39_13,N1508_6_r_12);
nand I_58(n39_13,N1507_6_r_12,N6147_9_r_12);
not I_59(n40_13,n36_13);
nor I_60(n41_13,n35_13,N1508_0_r_12);
not I_61(n42_13,n_569_7_r_12);
or I_62(n43_13,N1371_0_r_12,N6147_9_r_12);
not I_63(n44_13,N1371_0_r_12);
not I_64(n45_13,n_572_7_r_12);
nor I_65(n46_13,n39_13,n40_13);
nor I_66(n47_13,N1371_0_r_12,N6147_9_r_12);
nor I_67(n48_13,n50_13,n51_13);
nor I_68(n49_13,n_572_7_r_12,N1371_0_r_12);
not I_69(n50_13,n59_13);
not I_70(n51_13,n_102_5_r_13);
nand I_71(n52_13,n33_13,n39_13);
nand I_72(n53_13,n33_13,N1508_6_r_12);
nor I_73(n54_13,N1508_0_r_12,N6147_9_r_12);
nand I_74(n55_13,n62_13,n56_13);
nor I_75(n56_13,n39_13,n57_13);
not I_76(n57_13,N1371_0_r_12);
or I_77(n58_13,n_549_7_r_12,n_569_7_r_12);
nand I_78(n59_13,G42_7_r_12,n_572_7_r_12);
nor I_79(n60_13,n51_13,N6147_9_r_12);
nor I_80(n61_13,n39_13,N1508_6_r_12);
endmodule


