module test_I10038(I8107,I1477,I7621,I6321,I7714,I10069,I1470,I10038);
input I8107,I1477,I7621,I6321,I7714,I10069,I1470;
output I10038;
wire I7850,I10538,I10103,I7731,I10490,I10052,I7977,I10349,I10332,I7556,I7550,I10086,I7570,I7544,I7532;
nor I_0(I7850,I7731);
nor I_1(I10538,I10490,I10103);
DFFARX1 I_2(I10086,I1470,I10052,,,I10103,);
not I_3(I7731,I7714);
DFFARX1 I_4(I7556,I1470,I10052,,,I10490,);
not I_5(I10052,I1477);
DFFARX1 I_6(I6321,I1470,I7570,,,I7977,);
and I_7(I10349,I10332,I7550);
nand I_8(I10038,I10349,I10538);
DFFARX1 I_9(I7532,I1470,I10052,,,I10332,);
nand I_10(I7556,I7621,I7850);
nand I_11(I7550,I7977,I7731);
and I_12(I10086,I10069,I7544);
not I_13(I7570,I1477);
DFFARX1 I_14(I7621,I1470,I7570,,,I7544,);
DFFARX1 I_15(I8107,I1470,I7570,,,I7532,);
endmodule


