module test_I11201(I10647,I1470,I11201);
input I10647,I1470;
output I11201;
wire I10961,I9720,I10664,I9474,I9737,I9471,I10715,I9542,I9638,I11184,I11167,I9816,I9771,I9459,I8178,I11150,I10732,I9477,I9754,I9465,I9621,I9689;
nand I_0(I10961,I10664,I9459);
not I_1(I9720,I9689);
not I_2(I10664,I9471);
or I_3(I9474,I9542);
nor I_4(I9737,I9621,I9720);
nor I_5(I9471,I9689,I9542);
nor I_6(I10715,I10664,I9477);
DFFARX1 I_7(I1470,,,I9542,);
nor I_8(I9638,I9621);
nand I_9(I11184,I11167,I10732);
not I_10(I11167,I11150);
DFFARX1 I_11(I1470,,,I9816,);
and I_12(I9771,I9754,I8178);
nand I_13(I9459,I9771,I9737);
DFFARX1 I_14(I1470,,,I8178,);
DFFARX1 I_15(I9474,I1470,I10647,,,I11150,);
nand I_16(I10732,I10715,I9465);
nor I_17(I9477,I9771);
DFFARX1 I_18(I1470,,,I9754,);
nand I_19(I9465,I9816,I9638);
and I_20(I11201,I10961,I11184);
DFFARX1 I_21(I1470,,,I9621,);
DFFARX1 I_22(I1470,,,I9689,);
endmodule


