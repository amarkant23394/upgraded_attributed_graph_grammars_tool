module test_I16852(I12605,I15047,I1477,I1470,I15194,I15423,I16852);
input I12605,I15047,I1477,I1470,I15194,I15423;
output I16852;
wire I14948,I15502,I15211,I15064,I14936,I16835,I12587,I15519,I14965,I15228,I15485,I14957;
DFFARX1 I_0(I15519,I1470,I14965,,,I14948,);
not I_1(I15502,I15485);
DFFARX1 I_2(I15194,I1470,I14965,,,I15211,);
nand I_3(I15064,I15047,I12587);
DFFARX1 I_4(I15064,I1470,I14965,,,I14936,);
nand I_5(I16835,I14936,I14948);
and I_6(I16852,I16835,I14957);
DFFARX1 I_7(I1470,,,I12587,);
or I_8(I15519,I15502,I15423);
not I_9(I14965,I1477);
nor I_10(I15228,I15211,I15064);
DFFARX1 I_11(I12605,I1470,I14965,,,I15485,);
nand I_12(I14957,I15502,I15228);
endmodule


