module test_I4527(I1477,I2311,I1239,I1303,I1470,I4527);
input I1477,I2311,I1239,I1303,I1470;
output I4527;
wire I2167,I4629,I4595,I4544,I2328,I2633,I2540,I4561,I2458,I2152,I4578,I2161,I2345,I2173,I2181,I2509,I2557,I2232;
nand I_0(I2167,I2633,I2328);
nor I_1(I4629,I2167,I2173);
DFFARX1 I_2(I4578,I1470,I4544,,,I4595,);
not I_3(I4544,I1477);
nor I_4(I2328,I2232,I2311);
or I_5(I4527,I4629,I4595);
DFFARX1 I_6(I1239,I1470,I2181,,,I2633,);
DFFARX1 I_7(I1470,I2181,,,I2540,);
nand I_8(I4561,I2152,I2173);
DFFARX1 I_9(I1470,I2181,,,I2458,);
DFFARX1 I_10(I2458,I1470,I2181,,,I2152,);
and I_11(I4578,I4561,I2161);
nand I_12(I2161,I2345,I2311);
DFFARX1 I_13(I1470,I2181,,,I2345,);
nand I_14(I2173,I2557,I2509);
not I_15(I2181,I1477);
nor I_16(I2509,I2458,I2232);
and I_17(I2557,I2540,I1303);
DFFARX1 I_18(I1470,I2181,,,I2232,);
endmodule


