module test_I16452(I13177,I1477,I13186,I13162,I1470,I16452);
input I13177,I1477,I13186,I13162,I1470;
output I16452;
wire I14362,I14667,I14455,I14421,I16435,I14715,I14684,I14350,I14650,I14808,I14537,I14359,I14370,I14825,I13159,I14438,I13189,I14732;
DFFARX1 I_0(I14825,I1470,I14370,,,I14362,);
and I_1(I14667,I14650,I13189);
DFFARX1 I_2(I13177,I1470,I14370,,,I14455,);
DFFARX1 I_3(I1470,I14370,,,I14421,);
nand I_4(I16435,I14359,I14350);
not I_5(I14715,I14667);
nand I_6(I14684,I14667,I14537);
nand I_7(I14350,I14455,I14732);
and I_8(I16452,I16435,I14362);
DFFARX1 I_9(I1470,I14370,,,I14650,);
DFFARX1 I_10(I13162,I1470,I14370,,,I14808,);
DFFARX1 I_11(I1470,I14370,,,I14537,);
nor I_12(I14359,I14667,I14438);
not I_13(I14370,I1477);
and I_14(I14825,I14808,I14684);
DFFARX1 I_15(I1470,,,I13159,);
nor I_16(I14438,I13159,I13186);
DFFARX1 I_17(I1470,,,I13189,);
nor I_18(I14732,I14421,I14715);
endmodule


