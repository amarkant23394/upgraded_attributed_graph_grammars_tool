module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_5_r_7,n6_7,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
nor I_34(N1371_0_r_7,n53_7,n52_7);
nor I_35(N1508_0_r_7,n51_7,n52_7);
nand I_36(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_37(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_38(n_576_5_r_7,n31_7,n32_7);
nor I_39(n_102_5_r_7,N1508_0_r_12,N1507_6_r_12);
nand I_40(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_41(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_42(n_572_7_r_7,n54_7,n33_7);
nand I_43(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_44(n_549_7_r_7,n53_7,n36_7);
nand I_45(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_46(n_452_7_r_7,n_572_7_r_12,n_549_7_r_12);
nor I_47(n4_7_l_7,G42_7_r_12,n_572_7_r_12);
not I_48(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_49(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_50(n30_7,n53_7);
and I_51(N3_8_l_7,n50_7,N6147_9_r_12);
DFFARX1 I_52(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_53(n_431_5_r_7,n40_7,n41_7);
nor I_54(n4_7_r_7,n54_7,n49_7);
and I_55(n31_7,n_102_5_r_7,n39_7);
not I_56(n32_7,G42_7_r_12);
nor I_57(n33_7,n34_7,N1508_6_r_12);
and I_58(n34_7,n35_7,N1371_0_r_12);
not I_59(n35_7,N1371_0_r_12);
nor I_60(n36_7,n37_7,G42_7_r_12);
or I_61(n37_7,n54_7,N1508_0_r_12);
or I_62(n38_7,N1508_6_r_12,N1507_6_r_12);
nor I_63(n39_7,n_452_7_r_7,N1508_0_r_12);
nand I_64(n40_7,n46_7,n47_7);
nand I_65(n41_7,n42_7,n43_7);
nor I_66(n42_7,n44_7,n45_7);
nor I_67(n43_7,N1508_6_r_12,N1507_6_r_12);
nor I_68(n44_7,n_569_7_r_12,N1371_0_r_12);
nor I_69(n45_7,N1507_6_r_12,N1508_6_r_12);
nand I_70(n46_7,n35_7,N1371_0_r_12);
not I_71(n47_7,N1508_6_r_12);
or I_72(n48_7,n_452_7_r_7,N1508_0_r_12);
not I_73(n49_7,n_452_7_r_7);
nand I_74(n50_7,N1508_6_r_12,n_549_7_r_12);
and I_75(n51_7,n_452_7_r_7,n45_7);
not I_76(n52_7,n44_7);
endmodule


