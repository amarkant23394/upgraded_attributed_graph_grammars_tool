module test_I10349(I6657,I6843,I6309,I6705,I1470_clk,I1477_rst,I10349);
input I6657,I6843,I6309,I6705,I1470_clk,I1477_rst;
output I10349;
wire I8107,I7731,I8090,I7977,I7532,I10052_rst,I10332,I7570_rst,I7550,I6321,I6329_rst,I6297,I7714;
not I_0(I8107,I8090);
not I_1(I7731,I7714);
DFFARX1 I_2 (I6309,I1470_clk,I7570_rst,I8090);
DFFARX1 I_3 (I6321,I1470_clk,I7570_rst,I7977);
DFFARX1 I_4 (I8107,I1470_clk,I7570_rst,I7532);
not I_5(I10052_rst,I1477_rst);
DFFARX1 I_6 (I7532,I1470_clk,I10052_rst,I10332);
not I_7(I7570_rst,I1477_rst);
nand I_8(I7550,I7977,I7731);
and I_9(I10349,I10332,I7550);
nand I_10(I6321,I6705,I6657);
not I_11(I6329_rst,I1477_rst);
DFFARX1 I_12 (I6843,I1470_clk,I6329_rst,I6297);
not I_13(I7714,I6297);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule