module test_final(G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3,n4_1_l_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n4_1_r_3,blif_clk_net_1_r_8,n8_8,G42_1_r_3,);
nor I_1(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_2(n_573_1_r_3,n26_3,n27_3);
nor I_3(n_549_1_r_3,n40_3,n32_3);
nand I_4(n_569_1_r_3,n27_3,n31_3);
and I_5(n_452_1_r_3,G18_1_l_3,n26_3);
nor I_6(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_7(N3_2_r_3,blif_clk_net_1_r_8,n8_8,G199_2_r_3,);
DFFARX1 I_8(n_572_1_l_3,blif_clk_net_1_r_8,n8_8,ACVQN2_3_r_3,);
nor I_9(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_10(n4_1_l_3,G18_1_l_3,IN_1_1_l_3);
DFFARX1 I_11(n4_1_l_3,blif_clk_net_1_r_8,n8_8,G42_1_l_3,);
not I_12(n22_3,G42_1_l_3);
DFFARX1 I_13(IN_1_3_l_3,blif_clk_net_1_r_8,n8_8,n40_3,);
DFFARX1 I_14(IN_2_3_l_3,blif_clk_net_1_r_8,n8_8,n25_internal_3,);
not I_15(n25_3,n25_internal_3);
nor I_16(n4_1_r_3,n40_3,n36_3);
nor I_17(N3_2_r_3,n26_3,n37_3);
nor I_18(n_572_1_l_3,G15_1_l_3,IN_7_1_l_3);
DFFARX1 I_19(G42_1_l_3,blif_clk_net_1_r_8,n8_8,ACVQN1_3_r_3,);
nor I_20(n26_3,IN_5_1_l_3,IN_9_1_l_3);
not I_21(n27_3,IN_10_1_l_3);
nor I_22(n28_3,IN_10_1_l_3,n29_3);
nor I_23(n29_3,G15_1_l_3,n30_3);
not I_24(n30_3,IN_4_1_l_3);
nor I_25(n31_3,IN_9_1_l_3,n40_3);
nor I_26(n32_3,n25_3,n33_3);
nand I_27(n33_3,IN_4_3_l_3,n22_3);
or I_28(n34_3,IN_9_1_l_3,IN_10_1_l_3);
nand I_29(n35_3,IN_4_3_l_3,ACVQN1_3_r_3);
nor I_30(n36_3,G18_1_l_3,IN_5_1_l_3);
nor I_31(n37_3,n38_3,n39_3);
not I_32(n38_3,n_572_1_l_3);
nand I_33(n39_3,n27_3,n30_3);
DFFARX1 I_34(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_35(n_572_1_r_8,n39_8,n23_8);
and I_36(n_549_1_r_8,n38_8,n23_8);
nand I_37(n_569_1_r_8,n38_8,n24_8);
nor I_38(n_452_1_r_8,n25_8,n26_8);
nor I_39(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_40(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_41(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_42(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_43(n_431_0_l_8,n29_8,n_572_1_r_3);
not I_44(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_45(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_46(n19_8,G78_0_l_8);
DFFARX1 I_47(n_573_1_r_3,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_48(n22_8,n39_8);
DFFARX1 I_49(ACVQN2_3_r_3,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_50(n4_1_r_8,G78_0_l_8,n33_8);
nor I_51(N3_2_r_8,n22_8,n35_8);
nor I_52(N1_4_r_8,n27_8,n37_8);
nand I_53(n23_8,n32_8,n_266_and_0_3_r_3);
not I_54(n24_8,n23_8);
nand I_55(n25_8,n36_8,G42_1_r_3);
nand I_56(n26_8,n27_8,n28_8);
nor I_57(n27_8,n31_8,n_569_1_r_3);
not I_58(n28_8,n_42_2_r_3);
and I_59(n29_8,n30_8,G42_1_r_3);
nor I_60(n30_8,n31_8,G199_2_r_3);
not I_61(n31_8,n_549_1_r_3);
and I_62(n32_8,n28_8,n_569_1_r_3);
nand I_63(n33_8,n28_8,n34_8);
not I_64(n34_8,n25_8);
nor I_65(n35_8,n34_8,n_42_2_r_3);
not I_66(n36_8,n_452_1_r_3);
nor I_67(n37_8,n19_8,n38_8);
endmodule


