module test_I3637(I1637,I1383,I1477,I1423,I1586,I1470,I3637);
input I1637,I1383,I1477,I1423,I1586,I1470;
output I3637;
wire I1518,I3388,I1668,I3620,I1880,I1603,I1492,I1483;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
not I_2(I1668,I1637);
nor I_3(I3620,I1492,I1483);
DFFARX1 I_4(I3620,I1470,I3388,,,I3637,);
DFFARX1 I_5(I1383,I1470,I1518,,,I1880,);
nand I_6(I1603,I1586,I1423);
nand I_7(I1492,I1603,I1668);
DFFARX1 I_8(I1880,I1470,I1518,,,I1483,);
endmodule


