module test_I4181(I1415,I2776,I3217,I2946,I1477,I1470,I4181);
input I1415,I2776,I3217,I2946,I1477,I1470;
output I4181;
wire I2759,I3234,I4147,I2963,I4164,I2739,I2980,I2748,I2736,I3983;
not I_0(I2759,I1477);
nor I_1(I3234,I3217);
nand I_2(I4147,I2739,I2736);
DFFARX1 I_3(I2946,I1470,I2759,,,I2963,);
and I_4(I4164,I4147,I2748);
nor I_5(I2739,I3217,I2980);
DFFARX1 I_6(I4164,I1470,I3983,,,I4181,);
nand I_7(I2980,I2776,I1415);
or I_8(I2748,I2980,I2963);
DFFARX1 I_9(I3234,I1470,I2759,,,I2736,);
not I_10(I3983,I1477);
endmodule


