module test_I13313(I9320,I1477,I1470,I9210,I13313);
input I9320,I1477,I1470,I9210;
output I13313;
wire I11672,I8836,I13197,I11293,I11310;
DFFARX1 I_0(I11293,I1470,I13197,,,I13313,);
DFFARX1 I_1(I8836,I1470,I11310,,,I11672,);
nand I_2(I8836,I9320,I9210);
not I_3(I13197,I1477);
not I_4(I11293,I11672);
not I_5(I11310,I1477);
endmodule


