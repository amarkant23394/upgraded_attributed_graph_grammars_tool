module test_I17304(I15016,I1477,I1470,I15245,I17304);
input I15016,I1477,I1470,I15245;
output I17304;
wire I14927,I14948,I15485,I14951,I17287,I17205,I16818,I17270,I15519,I14965,I16886,I15502;
DFFARX1 I_0(I15502,I1470,I14965,,,I14927,);
DFFARX1 I_1(I15519,I1470,I14965,,,I14948,);
DFFARX1 I_2(I1470,I14965,,,I15485,);
nand I_3(I14951,I15016,I15245);
and I_4(I17304,I17205,I17287);
nor I_5(I17287,I16886,I17270);
DFFARX1 I_6(I14927,I1470,I16818,,,I17205,);
not I_7(I16818,I1477);
not I_8(I17270,I17205);
or I_9(I15519,I15502);
not I_10(I14965,I1477);
nor I_11(I16886,I14951,I14948);
not I_12(I15502,I15485);
endmodule


