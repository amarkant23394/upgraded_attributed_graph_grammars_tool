module test_I13618(I8836,I1477,I1470,I8848,I8851,I13618);
input I8836,I1477,I1470,I8848,I8851;
output I13618;
wire I13313,I11672,I11378,I13601,I11429,I13197,I11299,I11293,I11395,I11310;
DFFARX1 I_0(I11293,I1470,I13197,,,I13313,);
DFFARX1 I_1(I8836,I1470,I11310,,,I11672,);
nor I_2(I11378,I8848);
DFFARX1 I_3(I11299,I1470,I13197,,,I13601,);
not I_4(I11429,I8848);
not I_5(I13197,I1477);
nor I_6(I11299,I11395,I11429);
not I_7(I11293,I11672);
nand I_8(I11395,I11378,I8851);
not I_9(I11310,I1477);
nand I_10(I13618,I13601,I13313);
endmodule


