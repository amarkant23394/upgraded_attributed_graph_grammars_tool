module test_I8233(I5994,I1477,I1470,I8233);
input I5994,I1477,I1470;
output I8233;
wire I5751,I6028,I6011,I4521,I5722;
not I_0(I8233,I5722);
not I_1(I5751,I1477);
DFFARX1 I_2(I6011,I1470,I5751,,,I6028,);
and I_3(I6011,I5994,I4521);
DFFARX1 I_4(I1470,,,I4521,);
DFFARX1 I_5(I6028,I1470,I5751,,,I5722,);
endmodule


