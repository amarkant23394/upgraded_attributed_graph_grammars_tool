module test_I17464(I1477,I15662,I13749,I15781,I16069,I15696,I15628,I1470,I17464);
input I1477,I15662,I13749,I15781,I16069,I15696,I15628,I1470;
output I17464;
wire I13746,I14083,I15832,I15815,I15611,I15928,I15597,I15588,I16145,I16162,I17447,I16086,I13767,I15594,I15798;
not I_0(I13746,I14083);
DFFARX1 I_1(I1470,,,I14083,);
nand I_2(I15832,I15628,I13749);
DFFARX1 I_3(I15798,I1470,I15611,,,I15815,);
not I_4(I15611,I1477);
DFFARX1 I_5(I13746,I1470,I15611,,,I15928,);
nor I_6(I15597,I15832,I16162);
DFFARX1 I_7(I16086,I1470,I15611,,,I15588,);
not I_8(I16145,I16069);
and I_9(I16162,I15696,I16145);
nor I_10(I17447,I15597,I15588);
nor I_11(I16086,I16069,I15662);
DFFARX1 I_12(I1470,,,I13767,);
or I_13(I15594,I15928,I15815);
nand I_14(I17464,I17447,I15594);
or I_15(I15798,I15781,I13767);
endmodule


