module test_I12814(I1477,I10664,I9638,I9477,I10913,I1470,I12814);
input I1477,I10664,I9638,I9477,I10913,I1470;
output I12814;
wire I10647,I10978,I10961,I10715,I10797,I11167,I9816,I10766,I11150,I10732,I10621,I11232,I10624,I9465;
not I_0(I10647,I1477);
and I_1(I10978,I10961,I10913);
nand I_2(I10961,I10664);
nand I_3(I12814,I10624,I10621);
nor I_4(I10715,I10664,I9477);
not I_5(I10797,I10766);
not I_6(I11167,I11150);
DFFARX1 I_7(I1470,,,I9816,);
not I_8(I10766,I9477);
DFFARX1 I_9(I1470,I10647,,,I11150,);
nand I_10(I10732,I10715,I9465);
nand I_11(I10621,I10732,I10797);
or I_12(I11232,I11167,I10978);
DFFARX1 I_13(I11232,I1470,I10647,,,I10624,);
nand I_14(I9465,I9816,I9638);
endmodule


