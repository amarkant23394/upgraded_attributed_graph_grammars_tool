module test_I1684(I1263,I1207,I1684);
input I1263,I1207;
output I1684;
wire I1359;
not I_0(I1359,I1263);
nand I_1(I1684,I1359,I1207);
endmodule


