module test_I6028(I1477,I1470,I4824,I4773,I6028);
input I1477,I1470,I4824,I4773;
output I6028;
wire I4917,I5994,I5751,I6011,I4521,I4512,I4506,I4544,I4869,I4674,I4790;
nor I_0(I4917,I4869,I4674);
nand I_1(I5994,I4512,I4506);
not I_2(I5751,I1477);
DFFARX1 I_3(I6011,I1470,I5751,,,I6028,);
and I_4(I6011,I5994,I4521);
DFFARX1 I_5(I4917,I1470,I4544,,,I4521,);
nand I_6(I4512,I4824,I4790);
nand I_7(I4506,I4869,I4773);
not I_8(I4544,I1477);
DFFARX1 I_9(I1470,I4544,,,I4869,);
DFFARX1 I_10(I1470,I4544,,,I4674,);
nor I_11(I4790,I4674,I4773);
endmodule


