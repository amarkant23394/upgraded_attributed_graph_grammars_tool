module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_5_r_11,n9_11,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
not I_36(N1372_1_r_11,n53_11);
nor I_37(N1508_1_r_11,n39_11,n53_11);
nor I_38(N6147_2_r_11,n48_11,n49_11);
nor I_39(N6147_3_r_11,n44_11,n45_11);
nand I_40(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_41(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_42(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_43(n_102_5_r_11,n39_11);
nand I_44(n_547_5_r_11,n36_11,n37_11);
nor I_45(N1507_6_r_11,n52_11,n57_11);
nor I_46(N1508_6_r_11,n46_11,n51_11);
nor I_47(N1372_10_r_11,n43_11,n47_11);
nor I_48(N1508_10_r_11,n55_11,n56_11);
nand I_49(n_431_5_r_11,n40_11,n41_11);
not I_50(n9_11,blif_reset_net_5_r_11);
nor I_51(n36_11,n38_11,n39_11);
not I_52(n37_11,n40_11);
nor I_53(n38_11,n60_11,N1371_0_r_5);
nor I_54(n39_11,n54_11,N1508_1_r_5);
nand I_55(n40_11,G42_7_r_5,N1508_0_r_5);
nand I_56(n41_11,n_102_5_r_11,n42_11);
and I_57(n42_11,n58_11,N1507_6_r_5);
not I_58(n43_11,n44_11);
nor I_59(n44_11,n40_11,n_572_7_r_5);
nand I_60(n45_11,n46_11,n47_11);
not I_61(n46_11,n38_11);
nand I_62(n47_11,n59_11,n62_11);
and I_63(n48_11,n37_11,n47_11);
or I_64(n49_11,n44_11,n50_11);
nor I_65(n50_11,n60_11,n61_11);
or I_66(n51_11,n_102_5_r_11,n52_11);
nor I_67(n52_11,n42_11,n57_11);
nand I_68(n53_11,n37_11,n50_11);
or I_69(n54_11,N1372_1_r_5,N1508_6_r_5);
nor I_70(n55_11,n38_11,n42_11);
not I_71(n56_11,N1372_10_r_11);
and I_72(n57_11,n38_11,n50_11);
and I_73(n58_11,n59_11,n_452_7_r_5);
or I_74(n59_11,n63_11,N1508_0_r_5);
not I_75(n60_11,N6147_2_r_5);
nor I_76(n61_11,N1371_0_r_5,n_569_7_r_5);
nand I_77(n62_11,n_573_7_r_5,N1372_1_r_5);
and I_78(n63_11,n_573_7_r_5,N1372_1_r_5);
endmodule


