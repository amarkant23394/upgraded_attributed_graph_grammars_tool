module test_I2963(I1391,I2895,I1311,I1263,I1470_clk,I1477_rst,I2963);
input I1391,I2895,I1311,I1263,I1470_clk,I1477_rst;
output I2963;
wire I2929,I2946,I2759_rst,I2912;
and I_0(I2929,I2912,I1391);
DFFARX1 I_1 (I2946,I1470_clk,I2759_rst,I2963);
or I_2(I2946,I2929,I1263);
not I_3(I2759_rst,I1477_rst);
nor I_4(I2912,I2895,I1311);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule