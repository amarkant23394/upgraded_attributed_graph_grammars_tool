module test_I2748(I1415,I1391,I1263,I1477,I1470,I2912,I1407,I2748);
input I1415,I1391,I1263,I1477,I1470,I2912,I1407;
output I2748;
wire I2759,I2946,I2929,I2963,I2980,I2776;
not I_0(I2759,I1477);
or I_1(I2946,I2929,I1263);
and I_2(I2929,I2912,I1391);
DFFARX1 I_3(I2946,I1470,I2759,,,I2963,);
or I_4(I2748,I2980,I2963);
nand I_5(I2980,I2776,I1415);
not I_6(I2776,I1407);
endmodule


