module Benchmark_testing100(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I3114,I3117,I3093,I3105,I3120,I3108,I3102,I3096,I3099,I3111);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458;
output I3114,I3117,I3093,I3105,I3120,I3108,I3102,I3096,I3099,I3111;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I1493,I2575,I1519,I1527,I1544,I2572,I2587,I1561,I2569,I1587,I2566,I1604,I1612,I1629,I1461,I1660,I1677,I1473,I1717,I1482,I1739,I2581,I1756,I2584,I1782,I1799,I1485,I1821,I1470,I1852,I2578,I1869,I1886,I1903,I1479,I1934,I1467,I1476,I1464,I2020,I2046,I2054,I2071,I2088,I2114,I2122,I2148,I2156,I2173,I2190,I2207,I2003,I2247,I2255,I2272,I2289,I2306,I2006,I2337,I2354,I2380,I2388,I1988,I2419,I1997,I2450,I2467,I2009,I2498,I2000,I1991,I1994,I2012,I2595,I2621,I2629,I2646,I2663,I2689,I2720,I2728,I2745,I2771,I2779,I2819,I2855,I2872,I2898,I2906,I2923,I2954,I2971,I2988,I3019,I3050,I3067,I3128,I3154,I3171,I3179,I3196,I3213,I3230,I3247,I3264,I3295,I3312,I3343,I3360,I3377,I3408,I3448,I3456,I3473,I3490,I3507,I3538,I3555,I3572,I3598,I3620,I3637,I3668,I3713;
not I_0 (I1493,I1458);
DFFARX1 I_1 (I2575,I1451,I1493,I1519,);
not I_2 (I1527,I1519);
nand I_3 (I1544,I2572,I2587);
and I_4 (I1561,I1544,I2569);
DFFARX1 I_5 (I1561,I1451,I1493,I1587,);
DFFARX1 I_6 (I2566,I1451,I1493,I1604,);
and I_7 (I1612,I1604,I2566);
nor I_8 (I1629,I1587,I1612);
DFFARX1 I_9 (I1629,I1451,I1493,I1461,);
nand I_10 (I1660,I1604,I2566);
nand I_11 (I1677,I1527,I1660);
not I_12 (I1473,I1677);
DFFARX1 I_13 (I2569,I1451,I1493,I1717,);
DFFARX1 I_14 (I1717,I1451,I1493,I1482,);
nand I_15 (I1739,I2581,I2572);
and I_16 (I1756,I1739,I2584);
DFFARX1 I_17 (I1756,I1451,I1493,I1782,);
DFFARX1 I_18 (I1782,I1451,I1493,I1799,);
not I_19 (I1485,I1799);
not I_20 (I1821,I1782);
nand I_21 (I1470,I1821,I1660);
nor I_22 (I1852,I2578,I2572);
not I_23 (I1869,I1852);
nor I_24 (I1886,I1821,I1869);
nor I_25 (I1903,I1527,I1886);
DFFARX1 I_26 (I1903,I1451,I1493,I1479,);
nor I_27 (I1934,I1587,I1869);
nor I_28 (I1467,I1782,I1934);
nor I_29 (I1476,I1717,I1852);
nor I_30 (I1464,I1587,I1852);
not I_31 (I2020,I1458);
DFFARX1 I_32 (I1464,I1451,I2020,I2046,);
not I_33 (I2054,I2046);
nand I_34 (I2071,I1473,I1482);
and I_35 (I2088,I2071,I1461);
DFFARX1 I_36 (I2088,I1451,I2020,I2114,);
not I_37 (I2122,I1464);
DFFARX1 I_38 (I1479,I1451,I2020,I2148,);
not I_39 (I2156,I2148);
nor I_40 (I2173,I2156,I2054);
and I_41 (I2190,I2173,I1464);
nor I_42 (I2207,I2156,I2122);
nor I_43 (I2003,I2114,I2207);
DFFARX1 I_44 (I1470,I1451,I2020,I2247,);
nor I_45 (I2255,I2247,I2114);
not I_46 (I2272,I2255);
not I_47 (I2289,I2247);
nor I_48 (I2306,I2289,I2190);
DFFARX1 I_49 (I2306,I1451,I2020,I2006,);
nand I_50 (I2337,I1485,I1461);
and I_51 (I2354,I2337,I1467);
DFFARX1 I_52 (I2354,I1451,I2020,I2380,);
nor I_53 (I2388,I2380,I2247);
DFFARX1 I_54 (I2388,I1451,I2020,I1988,);
nand I_55 (I2419,I2380,I2289);
nand I_56 (I1997,I2272,I2419);
not I_57 (I2450,I2380);
nor I_58 (I2467,I2450,I2190);
DFFARX1 I_59 (I2467,I1451,I2020,I2009,);
nor I_60 (I2498,I1476,I1461);
or I_61 (I2000,I2247,I2498);
nor I_62 (I1991,I2380,I2498);
or I_63 (I1994,I2114,I2498);
DFFARX1 I_64 (I2498,I1451,I2020,I2012,);
not I_65 (I2595,I1458);
DFFARX1 I_66 (I1380,I1451,I2595,I2621,);
not I_67 (I2629,I2621);
nand I_68 (I2646,I1372,I1396);
and I_69 (I2663,I2646,I1420);
DFFARX1 I_70 (I2663,I1451,I2595,I2689,);
DFFARX1 I_71 (I2689,I1451,I2595,I2584,);
DFFARX1 I_72 (I1428,I1451,I2595,I2720,);
nand I_73 (I2728,I2720,I1444);
not I_74 (I2745,I2728);
DFFARX1 I_75 (I2745,I1451,I2595,I2771,);
not I_76 (I2779,I2771);
nor I_77 (I2587,I2629,I2779);
DFFARX1 I_78 (I1412,I1451,I2595,I2819,);
nor I_79 (I2578,I2819,I2689);
nor I_80 (I2569,I2819,I2745);
nand I_81 (I2855,I1388,I1436);
and I_82 (I2872,I2855,I1404);
DFFARX1 I_83 (I2872,I1451,I2595,I2898,);
not I_84 (I2906,I2898);
nand I_85 (I2923,I2906,I2819);
nand I_86 (I2572,I2906,I2728);
nor I_87 (I2954,I1364,I1436);
and I_88 (I2971,I2819,I2954);
nor I_89 (I2988,I2906,I2971);
DFFARX1 I_90 (I2988,I1451,I2595,I2581,);
nor I_91 (I3019,I2621,I2954);
DFFARX1 I_92 (I3019,I1451,I2595,I2566,);
nor I_93 (I3050,I2898,I2954);
not I_94 (I3067,I3050);
nand I_95 (I2575,I3067,I2923);
not I_96 (I3128,I1458);
DFFARX1 I_97 (I1994,I1451,I3128,I3154,);
DFFARX1 I_98 (I1988,I1451,I3128,I3171,);
not I_99 (I3179,I3171);
not I_100 (I3196,I2003);
nor I_101 (I3213,I3196,I1988);
not I_102 (I3230,I1997);
nor I_103 (I3247,I3213,I2006);
nor I_104 (I3264,I3171,I3247);
DFFARX1 I_105 (I3264,I1451,I3128,I3114,);
nor I_106 (I3295,I2006,I1988);
nand I_107 (I3312,I3295,I2003);
DFFARX1 I_108 (I3312,I1451,I3128,I3117,);
nor I_109 (I3343,I3230,I2006);
nand I_110 (I3360,I3343,I1991);
nor I_111 (I3377,I3154,I3360);
DFFARX1 I_112 (I3377,I1451,I3128,I3093,);
not I_113 (I3408,I3360);
nand I_114 (I3105,I3171,I3408);
DFFARX1 I_115 (I3360,I1451,I3128,I3448,);
not I_116 (I3456,I3448);
not I_117 (I3473,I2006);
not I_118 (I3490,I2000);
nor I_119 (I3507,I3490,I1997);
nor I_120 (I3120,I3456,I3507);
nor I_121 (I3538,I3490,I2009);
and I_122 (I3555,I3538,I2012);
or I_123 (I3572,I3555,I1991);
DFFARX1 I_124 (I3572,I1451,I3128,I3598,);
nor I_125 (I3108,I3598,I3154);
not I_126 (I3620,I3598);
and I_127 (I3637,I3620,I3154);
nor I_128 (I3102,I3179,I3637);
nand I_129 (I3668,I3620,I3230);
nor I_130 (I3096,I3490,I3668);
nand I_131 (I3099,I3620,I3408);
nand I_132 (I3713,I3230,I2000);
nor I_133 (I3111,I3473,I3713);
endmodule


