module test_final(IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_10,blif_reset_net_1_r_10,G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10);
input IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_10,blif_reset_net_1_r_10;
output G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10;
wire G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5,N3_2_l_5,G199_2_l_5,ACVQN2_3_l_5,n13_5,ACVQN1_3_l_5,N1_4_l_5,n21_5,n15_5,n22_5,n4_1_r_5,n11_internal_5,n11_5,n_42_2_l_5,n1_5,P6_5_r_internal_5,n16_5,n17_5,n18_5,n19_5,n20_5,n_452_1_r_10,N3_2_l_10,n4_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10;
DFFARX1 I_0(n4_1_r_5,blif_clk_net_1_r_10,n4_10,G42_1_r_5,);
nor I_1(n_572_1_r_5,n21_5,n22_5);
nand I_2(n_573_1_r_5,n13_5,n16_5);
nor I_3(n_549_1_r_5,n21_5,n17_5);
nand I_4(n_569_1_r_5,n13_5,n15_5);
nor I_5(n_452_1_r_5,n22_5,n_42_2_l_5);
DFFARX1 I_6(G199_2_l_5,blif_clk_net_1_r_10,n4_10,ACVQN2_3_r_5,);
nor I_7(n_266_and_0_3_r_5,n11_5,n16_5);
DFFARX1 I_8(n_42_2_l_5,blif_clk_net_1_r_10,n4_10,ACVQN1_5_r_5,);
not I_9(P6_5_r_5,P6_5_r_internal_5);
and I_10(N3_2_l_5,IN_6_2_l_5,n19_5);
DFFARX1 I_11(N3_2_l_5,blif_clk_net_1_r_10,n4_10,G199_2_l_5,);
DFFARX1 I_12(IN_1_3_l_5,blif_clk_net_1_r_10,n4_10,ACVQN2_3_l_5,);
not I_13(n13_5,ACVQN2_3_l_5);
DFFARX1 I_14(IN_2_3_l_5,blif_clk_net_1_r_10,n4_10,ACVQN1_3_l_5,);
and I_15(N1_4_l_5,IN_6_4_l_5,n20_5);
DFFARX1 I_16(N1_4_l_5,blif_clk_net_1_r_10,n4_10,n21_5,);
not I_17(n15_5,n21_5);
DFFARX1 I_18(IN_3_4_l_5,blif_clk_net_1_r_10,n4_10,n22_5,);
nor I_19(n4_1_r_5,G199_2_l_5,n22_5);
DFFARX1 I_20(ACVQN2_3_l_5,blif_clk_net_1_r_10,n4_10,n11_internal_5,);
not I_21(n11_5,n11_internal_5);
nor I_22(n_42_2_l_5,IN_1_2_l_5,IN_3_2_l_5);
not I_23(n1_5,n18_5);
DFFARX1 I_24(n1_5,blif_clk_net_1_r_10,n4_10,P6_5_r_internal_5,);
not I_25(n16_5,n_42_2_l_5);
nor I_26(n17_5,n22_5,n18_5);
nand I_27(n18_5,IN_4_3_l_5,ACVQN1_3_l_5);
nand I_28(n19_5,IN_2_2_l_5,IN_3_2_l_5);
nand I_29(n20_5,IN_1_4_l_5,IN_2_4_l_5);
DFFARX1 I_30(n4_1_r_10,blif_clk_net_1_r_10,n4_10,G42_1_r_10,);
nor I_31(n_572_1_r_10,n26_10,n3_10);
nand I_32(n_573_1_r_10,n16_10,n18_10);
nand I_33(n_549_1_r_10,n19_10,n20_10);
nor I_34(n_452_1_r_10,n25_10,n21_10);
nor I_35(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_36(N3_2_r_10,blif_clk_net_1_r_10,n4_10,G199_2_r_10,);
DFFARX1 I_37(G199_4_l_10,blif_clk_net_1_r_10,n4_10,ACVQN2_3_r_10,);
nor I_38(n_266_and_0_3_r_10,n17_10,n13_10);
and I_39(N3_2_l_10,n23_10,n_569_1_r_5);
not I_40(n4_10,blif_reset_net_1_r_10);
DFFARX1 I_41(N3_2_l_10,blif_clk_net_1_r_10,n4_10,n25_10,);
not I_42(n16_10,n25_10);
DFFARX1 I_43(n_452_1_r_5,blif_clk_net_1_r_10,n4_10,n26_10,);
DFFARX1 I_44(n_266_and_0_3_r_5,blif_clk_net_1_r_10,n4_10,ACVQN1_3_l_10,);
and I_45(N1_4_l_10,n24_10,ACVQN2_3_r_5);
DFFARX1 I_46(N1_4_l_10,blif_clk_net_1_r_10,n4_10,G199_4_l_10,);
DFFARX1 I_47(n_549_1_r_5,blif_clk_net_1_r_10,n4_10,n27_10,);
not I_48(n17_10,n27_10);
nor I_49(n4_1_r_10,n27_10,n21_10);
nor I_50(N3_2_r_10,n16_10,n22_10);
not I_51(n3_10,n18_10);
DFFARX1 I_52(n3_10,blif_clk_net_1_r_10,n4_10,n13_internal_10,);
not I_53(n13_10,n13_internal_10);
nand I_54(n18_10,ACVQN1_3_l_10,n_572_1_r_5);
not I_55(n19_10,n_452_1_r_10);
nand I_56(n20_10,n16_10,n26_10);
nor I_57(n21_10,n_573_1_r_5,ACVQN1_5_r_5);
and I_58(n22_10,n26_10,n21_10);
nand I_59(n23_10,n_573_1_r_5,P6_5_r_5);
nand I_60(n24_10,G42_1_r_5,n_572_1_r_5);
endmodule


