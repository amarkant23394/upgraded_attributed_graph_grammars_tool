module test_I16903(I1477,I15423,I14999,I1470,I15126,I15502,I16903);
input I1477,I15423,I14999,I1470,I15126,I15502;
output I16903;
wire I14948,I14951,I14965,I12581,I16835,I16852,I14957,I16818,I15211,I15228,I15016,I14936,I16869,I15519,I15245,I16886;
DFFARX1 I_0(I15519,I1470,I14965,,,I14948,);
nand I_1(I14951,I15016,I15245);
not I_2(I14965,I1477);
nor I_3(I16903,I16886,I16869);
DFFARX1 I_4(I1470,,,I12581,);
nand I_5(I16835,I14936,I14948);
and I_6(I16852,I16835,I14957);
nand I_7(I14957,I15502,I15228);
not I_8(I16818,I1477);
DFFARX1 I_9(I1470,I14965,,,I15211,);
nor I_10(I15228,I15211);
nand I_11(I15016,I14999,I12581);
DFFARX1 I_12(I1470,I14965,,,I14936,);
DFFARX1 I_13(I16852,I1470,I16818,,,I16869,);
or I_14(I15519,I15502,I15423);
nor I_15(I15245,I15211,I15126);
nor I_16(I16886,I14951,I14948);
endmodule


