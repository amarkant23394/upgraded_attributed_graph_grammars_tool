module test_I6688(I2733,I4418,I1477,I1470,I4068,I6688);
input I2733,I4418,I1477,I1470,I4068;
output I6688;
wire I4246,I3948,I6329,I4452,I4263,I4435,I3983;
DFFARX1 I_0(I1470,I3983,,,I4246,);
DFFARX1 I_1(I4452,I1470,I3983,,,I3948,);
not I_2(I6329,I1477);
DFFARX1 I_3(I3948,I1470,I6329,,,I6688,);
or I_4(I4452,I4263,I4435);
and I_5(I4263,I4246,I2733);
and I_6(I4435,I4068,I4418);
not I_7(I3983,I1477);
endmodule


