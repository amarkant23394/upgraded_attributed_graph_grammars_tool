module test_I3960(I2810,I3217,I1477,I1470,I3960);
input I2810,I3217,I1477,I1470;
output I3960;
wire I3124,I2727,I4113,I3076,I4308,I4356,I2751,I3983;
DFFARX1 I_0(I4356,I1470,I3983,,,I3960,);
nor I_1(I3124,I3076);
nand I_2(I2727,I2810,I3124);
DFFARX1 I_3(I2751,I1470,I3983,,,I4113,);
DFFARX1 I_4(I1470,,,I3076,);
DFFARX1 I_5(I2727,I1470,I3983,,,I4308,);
nor I_6(I4356,I4308,I4113);
nor I_7(I2751,I3076,I3217);
not I_8(I3983,I1477);
endmodule


