module test_I3246_rst(I1301_rst,I3246_rst);
,I3246_rst);
input I1301_rst;
output I3246_rst;
wire ;
not I_0(I3246_rst,I1301_rst);
endmodule


