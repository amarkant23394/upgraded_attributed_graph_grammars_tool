module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_7_r_3,n10_3,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
not I_39(N1372_1_r_3,n40_3);
nor I_40(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_41(N1507_6_r_3,n31_3,n42_3);
nor I_42(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_43(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_44(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_45(n_573_7_r_3,n30_3,n31_3);
nor I_46(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_47(n_569_7_r_3,n30_3,n32_3);
nor I_48(n_452_7_r_3,n35_3,N1508_4_r_15);
not I_49(N6147_9_r_3,n32_3);
nor I_50(N6134_9_r_3,n36_3,n37_3);
not I_51(I_BUFF_1_9_r_3,n45_3);
nor I_52(n4_7_r_3,I_BUFF_1_9_r_3,N1508_4_r_15);
not I_53(n10_3,blif_reset_net_7_r_3);
not I_54(n30_3,n39_3);
not I_55(n31_3,n35_3);
nand I_56(n32_3,n41_3,n_576_5_r_15);
nor I_57(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_58(n34_3,n46_3,N1508_6_r_15);
nor I_59(n35_3,n43_3,n44_3);
not I_60(n36_3,n34_3);
nor I_61(n37_3,N6147_9_r_3,N1508_4_r_15);
or I_62(n38_3,n_572_7_r_3,n34_3);
nor I_63(n39_3,n44_3,n_429_or_0_5_r_15);
nand I_64(n40_3,n39_3,N1508_4_r_15);
nand I_65(n41_3,N1508_1_r_15,N1372_4_r_15);
nor I_66(n42_3,n34_3,n45_3);
not I_67(n43_3,N1508_1_r_15);
nor I_68(n44_3,N1508_4_r_15,n_576_5_r_15);
nand I_69(n45_3,n49_3,n50_3);
and I_70(n46_3,n47_3,n_429_or_0_5_r_15);
nand I_71(n47_3,n41_3,n48_3);
not I_72(n48_3,n_576_5_r_15);
nor I_73(n49_3,G78_5_r_15,n_547_5_r_15);
or I_74(n50_3,n51_3,G78_5_r_15);
nor I_75(n51_3,N1372_4_r_15,N1507_6_r_15);
endmodule


