module test_I4561(I1303,I1477,I1247,I1470,I2424,I1327,I2215,I4561);
input I1303,I1477,I1247,I1470,I2424,I1327,I2215;
output I4561;
wire I2540,I2441,I2173,I2181,I2509,I2557,I2458,I2232,I2152;
DFFARX1 I_0(I1247,I1470,I2181,,,I2540,);
and I_1(I2441,I2424,I1327);
nand I_2(I2173,I2557,I2509);
not I_3(I2181,I1477);
nor I_4(I2509,I2458,I2232);
nand I_5(I4561,I2152,I2173);
and I_6(I2557,I2540,I1303);
DFFARX1 I_7(I2441,I1470,I2181,,,I2458,);
DFFARX1 I_8(I2215,I1470,I2181,,,I2232,);
DFFARX1 I_9(I2458,I1470,I2181,,,I2152,);
endmodule


