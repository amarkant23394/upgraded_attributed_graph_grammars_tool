module test_I2736(I1351,I1319,I1431,I1477,I1470,I1335,I2736);
input I1351,I1319,I1431,I1477,I1470,I1335;
output I2736;
wire I3217,I2759,I2810,I3234,I3200,I2793;
not I_0(I3217,I3200);
not I_1(I2759,I1477);
nand I_2(I2810,I2793,I1335);
nor I_3(I3234,I3217,I2810);
DFFARX1 I_4(I1431,I1470,I2759,,,I3200,);
nor I_5(I2793,I1351,I1319);
DFFARX1 I_6(I3234,I1470,I2759,,,I2736,);
endmodule


