module test_I14083(I12270,I10041,I1470_clk,I1477_rst,I14083);
input I12270,I10041,I1470_clk,I1477_rst;
output I14083;
wire I13775_rst,I11962,I11956,I14066,I14049,I11973_rst,I12349;
not I_0(I13775_rst,I1477_rst);
nor I_1(I11962,I12349,I12270);
DFFARX1 I_2 (I14066,I1470_clk,I13775_rst,I14083);
not I_3(I11956,I12349);
and I_4(I14066,I14049,I11956);
DFFARX1 I_5 (I11962,I1470_clk,I13775_rst,I14049);
not I_6(I11973_rst,I1477_rst);
DFFARX1 I_7 (I10041,I1470_clk,I11973_rst,I12349);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule