module test_I4130(I1447,I2946,I3045,I1477,I1470,I4130);
input I1447,I2946,I3045,I1477,I1470;
output I4130;
wire I3217,I2742,I2759,I3155,I3200,I4113,I3076,I2963,I4068,I2724,I2751,I3983;
not I_0(I3217,I3200);
or I_1(I2742,I3076,I2963);
not I_2(I2759,I1477);
or I_3(I3155,I3076,I3045);
DFFARX1 I_4(I1470,I2759,,,I3200,);
DFFARX1 I_5(I2751,I1470,I3983,,,I4113,);
DFFARX1 I_6(I1447,I1470,I2759,,,I3076,);
DFFARX1 I_7(I2946,I1470,I2759,,,I2963,);
nor I_8(I4068,I2742,I2724);
nor I_9(I4130,I4113,I4068);
DFFARX1 I_10(I3155,I1470,I2759,,,I2724,);
nor I_11(I2751,I3076,I3217);
not I_12(I3983,I1477);
endmodule


