module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_7_r_1,n9_1,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
and I_42(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_43(N1508_0_r_1,n40_1,n44_1);
nor I_44(N1507_6_r_1,n43_1,n49_1);
nor I_45(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_46(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_47(n_572_7_r_1,n29_1,n30_1);
not I_48(n_573_7_r_1,n_452_7_r_1);
nor I_49(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_50(n_569_7_r_1,n30_1,n31_1);
nor I_51(n_452_7_r_1,n30_1,n32_1);
nor I_52(N6147_9_r_1,n35_1,n36_1);
nand I_53(N6134_9_r_1,n38_1,n39_1);
not I_54(I_BUFF_1_9_r_1,n40_1);
nor I_55(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_56(n9_1,blif_reset_net_7_r_1);
nor I_57(n29_1,n34_1,N6147_2_r_11);
nor I_58(n30_1,n33_1,n34_1);
nor I_59(n31_1,n54_1,N6147_2_r_11);
not I_60(n32_1,n48_1);
nor I_61(n33_1,N6147_3_r_11,n_547_5_r_11);
not I_62(n34_1,n_576_5_r_11);
nor I_63(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_64(n36_1,n29_1);
not I_65(n37_1,n41_1);
nand I_66(n38_1,I_BUFF_1_9_r_1,N6147_3_r_11);
nand I_67(n39_1,n37_1,n40_1);
nand I_68(n40_1,N1508_1_r_11,N1372_1_r_11);
nand I_69(n41_1,n52_1,G78_5_r_11);
or I_70(n42_1,n36_1,n43_1);
nor I_71(n43_1,n32_1,n49_1);
nand I_72(n44_1,n45_1,n46_1);
nand I_73(n45_1,n47_1,n48_1);
not I_74(n46_1,N6147_3_r_11);
not I_75(n47_1,n31_1);
nand I_76(n48_1,n50_1,N1508_1_r_11);
nor I_77(n49_1,n41_1,n47_1);
and I_78(n50_1,n51_1,n_429_or_0_5_r_11);
nand I_79(n51_1,n52_1,n53_1);
nand I_80(n52_1,N1372_1_r_11,N1508_10_r_11);
not I_81(n53_1,G78_5_r_11);
or I_82(n54_1,N1507_6_r_11,N1508_6_r_11);
nor I_83(n55_1,n29_1,N6147_3_r_11);
endmodule


