module test_final(IN_1_0_l_0,IN_2_0_l_0,IN_4_0_l_0,IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_6_1_l_0,IN_1_5_l_0,IN_2_5_l_0,IN_3_5_l_0,IN_6_5_l_0,blif_reset_net_0_r_6,blif_clk_net_0_r_6,ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6);
input IN_1_0_l_0,IN_2_0_l_0,IN_4_0_l_0,IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_6_1_l_0,IN_1_5_l_0,IN_2_5_l_0,IN_3_5_l_0,IN_6_5_l_0,blif_reset_net_0_r_6,blif_clk_net_0_r_6;
output ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6;
wire n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0,n1_0_r_6,ACVQN1_2_l_6,P6_2_l_6,P6_internal_2_l_6,n_429_or_0_3_l_6,n12_3_l_6,n_431_3_l_6,G78_3_l_6,n_576_3_l_6,n11_3_l_6,n_102_3_l_6,n_547_3_l_6,n13_3_l_6,n14_3_l_6,n15_3_l_6,n16_3_l_6,ACVQN1_0_r_6,P6_internal_2_r_6,n12_3_r_6,n_431_3_r_6,n11_3_r_6,n13_3_r_6,n14_3_r_6,n15_3_r_6,n16_3_r_6,N3_5_r_6,n3_5_r_6;
nand I_0(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_1(n_431_3_r_0,blif_clk_net_0_r_6,n1_0_r_6,G78_3_r_0,);
nand I_2(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_3(n_102_3_r_0,n_42_5_l_0);
nand I_4(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_5(n4_4_r_0,blif_clk_net_0_r_6,n1_0_r_6,G42_4_r_0,);
nor I_6(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_7(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_8(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_9(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_10(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
DFFARX1 I_11(IN_1_0_l_0,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_l_0,);
and I_12(n_266_and_0_0_l_0,IN_4_0_l_0,ACVQN1_0_l_0);
DFFARX1 I_13(IN_2_0_l_0,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_l_0,);
and I_14(N1_1_l_0,IN_6_1_l_0,n3_1_l_0);
DFFARX1 I_15(N1_1_l_0,blif_clk_net_0_r_6,n1_0_r_6,G199_1_l_0,);
DFFARX1 I_16(IN_3_1_l_0,blif_clk_net_0_r_6,n1_0_r_6,G214_1_l_0,);
nand I_17(n3_1_l_0,IN_1_1_l_0,IN_2_1_l_0);
nor I_18(n_42_5_l_0,IN_1_5_l_0,IN_3_5_l_0);
and I_19(N3_5_l_0,IN_6_5_l_0,n3_5_l_0);
DFFARX1 I_20(N3_5_l_0,blif_clk_net_0_r_6,n1_0_r_6,G199_5_l_0,);
nand I_21(n3_5_l_0,IN_2_5_l_0,IN_3_5_l_0);
not I_22(n12_3_r_0,G199_1_l_0);
or I_23(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_24(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_25(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_26(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_27(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_28(n16_3_r_0,ACVQN2_0_l_0);
nor I_29(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_30(n_87_4_r_0,G199_5_l_0);
and I_31(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
DFFARX1 I_32(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_r_6,);
and I_33(n_266_and_0_0_r_6,n_429_or_0_3_l_6,ACVQN1_0_r_6);
DFFARX1 I_34(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_r_6,);
not I_35(P6_2_r_6,P6_internal_2_r_6);
nand I_36(n_429_or_0_3_r_6,n_102_3_l_6,n12_3_r_6);
DFFARX1 I_37(n_431_3_r_6,blif_clk_net_0_r_6,n1_0_r_6,G78_3_r_6,);
nand I_38(n_576_3_r_6,P6_2_l_6,n11_3_r_6);
not I_39(n_102_3_r_6,ACVQN1_2_l_6);
nand I_40(n_547_3_r_6,n_576_3_l_6,n13_3_r_6);
nor I_41(n_42_5_r_6,ACVQN1_2_l_6,n_429_or_0_3_l_6);
DFFARX1 I_42(N3_5_r_6,blif_clk_net_0_r_6,n1_0_r_6,G199_5_r_6,);
not I_43(n1_0_r_6,blif_reset_net_0_r_6);
DFFARX1 I_44(n_547_3_r_0,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_l_6,);
not I_45(P6_2_l_6,P6_internal_2_l_6);
DFFARX1 I_46(n_576_3_r_0,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_l_6,);
nand I_47(n_429_or_0_3_l_6,n12_3_l_6,n_429_or_0_3_r_0);
not I_48(n12_3_l_6,n_102_3_r_0);
or I_49(n_431_3_l_6,n14_3_l_6,n_452_4_r_0);
DFFARX1 I_50(n_431_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,G78_3_l_6,);
nand I_51(n_576_3_l_6,n11_3_l_6,G78_3_r_0);
nor I_52(n11_3_l_6,n12_3_l_6,n_549_4_r_0);
not I_53(n_102_3_l_6,n_549_4_r_0);
nand I_54(n_547_3_l_6,n13_3_l_6,n_569_4_r_0);
nor I_55(n13_3_l_6,n_572_4_r_0,n_549_4_r_0);
and I_56(n14_3_l_6,n15_3_l_6,n_573_4_r_0);
nor I_57(n15_3_l_6,n16_3_l_6,G42_4_r_0);
not I_58(n16_3_l_6,n_429_or_0_3_r_0);
DFFARX1 I_59(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_r_6,);
DFFARX1 I_60(n_576_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_r_6,);
not I_61(n12_3_r_6,P6_2_l_6);
or I_62(n_431_3_r_6,n_429_or_0_3_l_6,n14_3_r_6);
nor I_63(n11_3_r_6,ACVQN1_2_l_6,n12_3_r_6);
nor I_64(n13_3_r_6,ACVQN1_2_l_6,n_547_3_l_6);
and I_65(n14_3_r_6,ACVQN1_2_l_6,n15_3_r_6);
nor I_66(n15_3_r_6,P6_2_l_6,n16_3_r_6);
not I_67(n16_3_r_6,n_102_3_l_6);
and I_68(N3_5_r_6,n_102_3_l_6,n3_5_r_6);
nand I_69(n3_5_r_6,n_429_or_0_3_l_6,n_547_3_l_6);
endmodule


