module test_I5722(I4917,I1477,I4512,I4506,I1470,I5722);
input I4917,I1477,I4512,I4506,I1470;
output I5722;
wire I5994,I5751,I6028,I6011,I4521,I4544;
nand I_0(I5994,I4512,I4506);
not I_1(I5751,I1477);
DFFARX1 I_2(I6011,I1470,I5751,,,I6028,);
and I_3(I6011,I5994,I4521);
DFFARX1 I_4(I4917,I1470,I4544,,,I4521,);
not I_5(I4544,I1477);
DFFARX1 I_6(I6028,I1470,I5751,,,I5722,);
endmodule


