module test_I14244(I1477,I12024,I12041,I10026,I12270,I12106,I1470,I14244);
input I1477,I12024,I12041,I10026,I12270,I12106,I1470;
output I14244;
wire I12058,I12380,I13775,I13843,I11965,I12287,I12239,I12349,I11938,I12304,I14227,I14162,I11973,I11959;
nor I_0(I14244,I13843,I14227);
nand I_1(I12058,I12041,I10026);
nor I_2(I12380,I12349,I12024);
not I_3(I13775,I1477);
nor I_4(I13843,I11959,I11965);
DFFARX1 I_5(I12304,I1470,I11973,,,I11965,);
nand I_6(I12287,I12270,I12024);
DFFARX1 I_7(I1470,I11973,,,I12239,);
DFFARX1 I_8(I1470,I11973,,,I12349,);
and I_9(I11938,I12270,I12239);
and I_10(I12304,I12106,I12287);
not I_11(I14227,I14162);
DFFARX1 I_12(I11938,I1470,I13775,,,I14162,);
not I_13(I11973,I1477);
nand I_14(I11959,I12058,I12380);
endmodule


