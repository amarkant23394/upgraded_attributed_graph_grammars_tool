module test_I1543(I1231,I1279,I1475,I1294,I1301,I1287,I1239,I1543);
input I1231,I1279,I1475,I1294,I1301,I1287,I1239;
output I1543;
wire I1376,I1526,I1342,I1509,I1359,I1393,I1492;
nor I_0(I1543,I1393,I1526);
and I_1(I1376,I1359,I1231);
not I_2(I1526,I1509);
not I_3(I1342,I1301);
DFFARX1 I_4(I1492,I1294,I1342,,,I1509,);
nand I_5(I1359,I1287,I1239);
DFFARX1 I_6(I1376,I1294,I1342,,,I1393,);
and I_7(I1492,I1475,I1279);
endmodule


