module test_I2263(I1343,I1231,I1477,I1470,I1271,I2263);
input I1343,I1231,I1477,I1470,I1271;
output I2263;
wire I2181,I2232,I2198,I2215;
not I_0(I2181,I1477);
DFFARX1 I_1(I2215,I1470,I2181,,,I2232,);
nand I_2(I2198,I1343,I1231);
DFFARX1 I_3(I2232,I1470,I2181,,,I2263,);
and I_4(I2215,I2198,I1271);
endmodule


