module test_I8181(I1477,I6248,I6127,I1470,I8181);
input I1477,I6248,I6127,I1470;
output I8181;
wire I8527,I6265,I8233,I8360,I8216,I5751,I5713,I8592,I5915,I5719,I5722;
nand I_0(I8527,I8233,I5713);
and I_1(I6265,I5915,I6248);
not I_2(I8233,I5722);
and I_3(I8181,I8360,I8592);
not I_4(I8360,I5719);
not I_5(I8216,I1477);
not I_6(I5751,I1477);
DFFARX1 I_7(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_8(I8527,I1470,I8216,,,I8592,);
DFFARX1 I_9(I1470,I5751,,,I5915,);
DFFARX1 I_10(I6265,I1470,I5751,,,I5719,);
DFFARX1 I_11(I1470,I5751,,,I5722,);
endmodule


