module test_I3653(I1908,I1294,I1301,I3653);
input I1908,I1294,I1301;
output I3653;
wire I2668,I2733,I3168,I1914,I2583,I3280,I2945,I2572,I2563,I2548,I3297,I2560,I2651,I2993,I3246,I2702,I3622,I3086,I3103;
nand I_0(I2668,I2651,I1914);
not I_1(I2733,I2702);
or I_2(I3168,I3103);
DFFARX1 I_3(I1294,,,I1914,);
not I_4(I2583,I1301);
nor I_5(I3280,I2548,I2560);
DFFARX1 I_6(I1294,I2583,,,I2945,);
nor I_7(I2572,I2668,I2702);
nand I_8(I2563,I3103,I2993);
DFFARX1 I_9(I2945,I1294,I2583,,,I2548,);
nor I_10(I3653,I3622,I3297);
nand I_11(I3297,I3280,I2563);
DFFARX1 I_12(I3168,I1294,I2583,,,I2560,);
nor I_13(I2651,I1908);
nor I_14(I2993,I2945,I2733);
not I_15(I3246,I1301);
not I_16(I2702,I1908);
DFFARX1 I_17(I2572,I1294,I3246,,,I3622,);
DFFARX1 I_18(I1294,I2583,,,I3086,);
not I_19(I3103,I3086);
endmodule


