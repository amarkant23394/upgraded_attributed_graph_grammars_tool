module test_final(G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_0,blif_reset_net_1_r_0,G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0);
input G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_0,blif_reset_net_1_r_0;
output G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0;
wire G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8,n_431_0_l_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n_569_1_r_0,n4_1_l_0,n6_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0;
DFFARX1 I_0(n4_1_r_8,blif_clk_net_1_r_0,n6_0,G42_1_r_8,);
nor I_1(n_572_1_r_8,n39_8,n23_8);
and I_2(n_549_1_r_8,n38_8,n23_8);
nand I_3(n_569_1_r_8,n38_8,n24_8);
nor I_4(n_452_1_r_8,n25_8,n26_8);
nor I_5(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_6(N3_2_r_8,blif_clk_net_1_r_0,n6_0,G199_2_r_8,);
DFFARX1 I_7(N1_4_r_8,blif_clk_net_1_r_0,n6_0,G199_4_r_8,);
DFFARX1 I_8(G78_0_l_8,blif_clk_net_1_r_0,n6_0,G214_4_r_8,);
or I_9(n_431_0_l_8,IN_8_0_l_8,n29_8);
DFFARX1 I_10(n_431_0_l_8,blif_clk_net_1_r_0,n6_0,G78_0_l_8,);
not I_11(n19_8,G78_0_l_8);
DFFARX1 I_12(IN_2_5_l_8,blif_clk_net_1_r_0,n6_0,n39_8,);
not I_13(n22_8,n39_8);
DFFARX1 I_14(IN_1_5_l_8,blif_clk_net_1_r_0,n6_0,n38_8,);
nor I_15(n4_1_r_8,G78_0_l_8,n33_8);
nor I_16(N3_2_r_8,n22_8,n35_8);
nor I_17(N1_4_r_8,n27_8,n37_8);
nand I_18(n23_8,IN_7_0_l_8,n32_8);
not I_19(n24_8,n23_8);
nand I_20(n25_8,IN_11_0_l_8,n36_8);
nand I_21(n26_8,n27_8,n28_8);
nor I_22(n27_8,IN_5_0_l_8,n31_8);
not I_23(n28_8,G2_0_l_8);
and I_24(n29_8,IN_2_0_l_8,n30_8);
nor I_25(n30_8,IN_4_0_l_8,n31_8);
not I_26(n31_8,G1_0_l_8);
and I_27(n32_8,IN_5_0_l_8,n28_8);
nand I_28(n33_8,n28_8,n34_8);
not I_29(n34_8,n25_8);
nor I_30(n35_8,G2_0_l_8,n34_8);
not I_31(n36_8,IN_10_0_l_8);
nor I_32(n37_8,n19_8,n38_8);
DFFARX1 I_33(n4_1_r_0,blif_clk_net_1_r_0,n6_0,G42_1_r_0,);
nor I_34(n_572_1_r_0,n23_0,G214_4_r_8);
nand I_35(n_573_1_r_0,n21_0,n22_0);
nand I_36(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_37(n_569_1_r_0,n21_0,n26_0);
nor I_38(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_39(N3_2_r_0,blif_clk_net_1_r_0,n6_0,G199_2_r_0,);
DFFARX1 I_40(N1_4_r_0,blif_clk_net_1_r_0,n6_0,G199_4_r_0,);
DFFARX1 I_41(n2_0,blif_clk_net_1_r_0,n6_0,G214_4_r_0,);
nor I_42(n4_1_l_0,n_569_1_r_8,G42_1_r_8);
not I_43(n6_0,blif_reset_net_1_r_0);
DFFARX1 I_44(n4_1_l_0,blif_clk_net_1_r_0,n6_0,n37_0,);
DFFARX1 I_45(n_549_1_r_8,blif_clk_net_1_r_0,n6_0,n38_0,);
not I_46(n20_0,n38_0);
DFFARX1 I_47(n_572_1_r_8,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_0,);
nor I_48(n4_1_r_0,n23_0,n_572_1_r_8);
nor I_49(N3_2_r_0,n31_0,n32_0);
nor I_50(N1_4_r_0,n29_0,n32_0);
not I_51(n2_0,n31_0);
nor I_52(n21_0,n37_0,G199_2_r_8);
not I_53(n22_0,G214_4_r_8);
nand I_54(n23_0,n20_0,n30_0);
nand I_55(n24_0,n38_0,n25_0);
nor I_56(n25_0,n_572_1_r_8,G199_2_r_8);
not I_57(n26_0,n_572_1_r_8);
not I_58(n27_0,n29_0);
nor I_59(n28_0,n_452_1_r_8,G199_4_r_8);
nand I_60(n29_0,n26_0,n33_0);
not I_61(n30_0,G199_2_r_8);
nand I_62(n31_0,ACVQN1_3_l_0,n_42_2_r_8);
and I_63(n32_0,n35_0,n36_0);
nand I_64(n33_0,n34_0,G42_1_r_8);
not I_65(n34_0,G199_4_r_8);
nor I_66(n35_0,n_569_1_r_8,G199_4_r_8);
nor I_67(n36_0,n_452_1_r_8,G214_4_r_8);
endmodule


