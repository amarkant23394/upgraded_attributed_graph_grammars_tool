module test_I9943(I8527,I1477,I9655,I8193,I5737,I8208,I1470,I9943);
input I8527,I1477,I9655,I8193,I5737,I8208,I1470;
output I9943;
wire I8202,I8496,I8216,I9816,I9909,I5719,I8377,I8250,I9491,I9672,I8181,I8360,I8592,I8462,I9926,I9576,I8267,I9689;
nand I_0(I8202,I8267,I8496);
nor I_1(I8496,I8462,I8377);
not I_2(I8216,I1477);
DFFARX1 I_3(I8193,I1470,I9491,,,I9816,);
not I_4(I9909,I9816);
DFFARX1 I_5(I1470,,,I5719,);
not I_6(I8377,I8360);
nor I_7(I8250,I5719);
not I_8(I9491,I1477);
and I_9(I9672,I9655,I8208);
and I_10(I8181,I8360,I8592);
not I_11(I8360,I5719);
DFFARX1 I_12(I8527,I1470,I8216,,,I8592,);
and I_13(I9943,I9576,I9926);
DFFARX1 I_14(I1470,I8216,,,I8462,);
nor I_15(I9926,I9689,I9909);
nor I_16(I9576,I8181,I8202);
nand I_17(I8267,I8250,I5737);
DFFARX1 I_18(I9672,I1470,I9491,,,I9689,);
endmodule


