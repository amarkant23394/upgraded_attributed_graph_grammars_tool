module test_I16202(I14667,I1477,I14520,I1470,I16202);
input I14667,I1477,I14520,I1470;
output I16202;
wire I14901,I14537,I14344,I14808,I16534,I16240,I14370,I16551,I14335,I14715;
DFFARX1 I_0(I14808,I1470,I14370,,,I14901,);
DFFARX1 I_1(I16551,I1470,I16240,,,I16202,);
DFFARX1 I_2(I14520,I1470,I14370,,,I14537,);
nand I_3(I14344,I14537,I14715);
DFFARX1 I_4(I1470,I14370,,,I14808,);
DFFARX1 I_5(I14335,I1470,I16240,,,I16534,);
not I_6(I16240,I1477);
not I_7(I14370,I1477);
and I_8(I16551,I16534,I14344);
and I_9(I14335,I14808,I14901);
not I_10(I14715,I14667);
endmodule


