module test_final(IN_1_1_l,IN_2_1_l,IN_3_1_l,G18_7_l,G15_7_l,IN_1_7_l,IN_4_7_l,IN_5_7_l,IN_7_7_l,IN_9_7_l,IN_10_7_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_5_r,blif_reset_net_5_r,N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N1372_4_r,N1508_4_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,N1507_6_r,N1508_6_r);
input IN_1_1_l,IN_2_1_l,IN_3_1_l,G18_7_l,G15_7_l,IN_1_7_l,IN_4_7_l,IN_5_7_l,IN_7_7_l,IN_9_7_l,IN_10_7_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_5_r,blif_reset_net_5_r;
output N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N1372_4_r,N1508_4_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,N1507_6_r,N1508_6_r;
wire N1372_1_l,N1508_1_l,n4_1_l,G42_7_l,n_87_7_l,n_572_7_l,n_573_7_l,n_549_7_l,n_569_7_l,n_452_7_l,n4_7_l,n7_7_l,N1372_10_l,N1508_10_l,n5_10_l,n6_10_l,n3_0_r,n4_0_r,n4_1_r,n6_4_r,n7_4_r,n8_4_r,n_431_5_r,n2_5_r,n11_5_r,n12_5_r,n13_5_r,n14_5_r,n15_5_r,n16_5_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r;
not I_0(N1372_1_l,n4_1_l);
nor I_1(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_2(n4_1_l,IN_1_1_l,IN_2_1_l);
DFFARX1 I_3(n4_7_l,blif_clk_net_5_r,n2_5_r,G42_7_l,);
not I_4(n_87_7_l,G15_7_l);
nor I_5(n_572_7_l,G15_7_l,IN_7_7_l);
or I_6(n_573_7_l,IN_5_7_l,IN_9_7_l);
nor I_7(n_549_7_l,IN_10_7_l,n7_7_l);
or I_8(n_569_7_l,IN_9_7_l,IN_10_7_l);
nor I_9(n_452_7_l,G18_7_l,IN_5_7_l);
nor I_10(n4_7_l,G18_7_l,IN_1_7_l);
and I_11(n7_7_l,IN_4_7_l,n_87_7_l);
not I_12(N1372_10_l,n6_10_l);
nor I_13(N1508_10_l,n5_10_l,n6_10_l);
nor I_14(n5_10_l,IN_3_10_l,IN_4_10_l);
nand I_15(n6_10_l,IN_1_10_l,IN_2_10_l);
nor I_16(N1371_0_r,n4_0_r,n_573_7_l);
nor I_17(N1508_0_r,n3_0_r,n4_0_r);
nor I_18(n3_0_r,N1508_1_l,N1508_10_l);
not I_19(n4_0_r,G42_7_l);
not I_20(N1372_1_r,n4_1_r);
nor I_21(N1508_1_r,n4_1_r,n_572_7_l);
nand I_22(n4_1_r,n_573_7_l,n_452_7_l);
not I_23(N1372_4_r,n7_4_r);
nor I_24(N1508_4_r,n6_4_r,n7_4_r);
nor I_25(n6_4_r,n8_4_r,n_569_7_l);
nand I_26(n7_4_r,N1508_1_l,n_572_7_l);
and I_27(n8_4_r,N1372_1_l,n_549_7_l);
nand I_28(n_429_or_0_5_r,n12_5_r,N1508_1_l);
DFFARX1 I_29(n_431_5_r,blif_clk_net_5_r,n2_5_r,G78_5_r,);
nand I_30(n_576_5_r,n11_5_r,n_569_7_l);
not I_31(n_102_5_r,n_452_7_l);
nand I_32(n_547_5_r,n13_5_r,n_549_7_l);
or I_33(n_431_5_r,n14_5_r,n_572_7_l);
not I_34(n2_5_r,blif_reset_net_5_r);
nor I_35(n11_5_r,n12_5_r,n_452_7_l);
not I_36(n12_5_r,N1372_10_l);
nor I_37(n13_5_r,N1372_1_l,n_452_7_l);
and I_38(n14_5_r,n15_5_r,n_573_7_l);
nor I_39(n15_5_r,n16_5_r,N1372_10_l);
not I_40(n16_5_r,N1508_1_l);
nor I_41(N1507_6_r,n8_6_r,n9_6_r);
and I_42(N1508_6_r,n6_6_r,N1508_10_l);
nor I_43(n6_6_r,n7_6_r,n8_6_r);
not I_44(n7_6_r,G42_7_l);
nor I_45(n8_6_r,n9_6_r,N1372_1_l);
and I_46(n9_6_r,G42_7_l,n_549_7_l);
endmodule


