module test_I14571(I1477,I14503,I1470,I13525,I13171,I14571);
input I1477,I14503,I1470,I13525,I13171;
output I14571;
wire I14554,I13601,I13183,I14520,I14404,I13186,I14421,I13174,I14537,I14387,I14370;
not I_0(I14554,I14537);
DFFARX1 I_1(I1470,,,I13601,);
nand I_2(I13183,I13601,I13525);
nor I_3(I14571,I14421,I14554);
and I_4(I14520,I14503,I13174);
and I_5(I14404,I14387,I13183);
nor I_6(I13186,I13601);
DFFARX1 I_7(I14404,I1470,I14370,,,I14421,);
DFFARX1 I_8(I1470,,,I13174,);
DFFARX1 I_9(I14520,I1470,I14370,,,I14537,);
nand I_10(I14387,I13171,I13186);
not I_11(I14370,I1477);
endmodule


