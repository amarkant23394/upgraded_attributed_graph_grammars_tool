module test_I17270(I1477,I1470,I17270);
input I1477,I1470;
output I17270;
wire I14927,I17205,I16818,I14965,I15485,I15502;
DFFARX1 I_0(I15502,I1470,I14965,,,I14927,);
DFFARX1 I_1(I14927,I1470,I16818,,,I17205,);
not I_2(I16818,I1477);
not I_3(I17270,I17205);
not I_4(I14965,I1477);
DFFARX1 I_5(I1470,I14965,,,I15485,);
not I_6(I15502,I15485);
endmodule


