module test_I17287(I14999,I15502,I1477,I1470,I15423,I15126,I17287);
input I14999,I15502,I1477,I1470,I15423,I15126;
output I17287;
wire I14927,I14948,I15016,I15211,I14951,I17205,I16818,I17270,I15519,I14965,I15245,I12581,I16886;
DFFARX1 I_0(I15502,I1470,I14965,,,I14927,);
DFFARX1 I_1(I15519,I1470,I14965,,,I14948,);
nand I_2(I15016,I14999,I12581);
DFFARX1 I_3(I1470,I14965,,,I15211,);
nand I_4(I14951,I15016,I15245);
nor I_5(I17287,I16886,I17270);
DFFARX1 I_6(I14927,I1470,I16818,,,I17205,);
not I_7(I16818,I1477);
not I_8(I17270,I17205);
or I_9(I15519,I15502,I15423);
not I_10(I14965,I1477);
nor I_11(I15245,I15211,I15126);
DFFARX1 I_12(I1470,,,I12581,);
nor I_13(I16886,I14951,I14948);
endmodule


