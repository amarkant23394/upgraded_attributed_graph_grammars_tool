module test_I2458(I1327,I1223,I1255,I1477,I1470,I2458);
input I1327,I1223,I1255,I1477,I1470;
output I2458;
wire I2441,I2181,I2424;
and I_0(I2441,I2424,I1327);
not I_1(I2181,I1477);
DFFARX1 I_2(I2441,I1470,I2181,,,I2458,);
nand I_3(I2424,I1223,I1255);
endmodule


