module test_I15585(I13761,I1477,I15628,I1470,I13843,I14278,I15585);
input I13761,I1477,I15628,I1470,I13843,I14278;
output I15585;
wire I14083,I13752,I15696,I13746,I16052,I13775,I15611,I15959,I13758,I15679,I15928,I16069;
DFFARX1 I_0(I1470,I13775,,,I14083,);
DFFARX1 I_1(I14278,I1470,I13775,,,I13752,);
nand I_2(I15696,I15679,I13758);
not I_3(I13746,I14083);
DFFARX1 I_4(I13752,I1470,I15611,,,I16052,);
not I_5(I13775,I1477);
nand I_6(I15585,I16069,I15959);
not I_7(I15611,I1477);
nor I_8(I15959,I15928,I15696);
not I_9(I13758,I13843);
nor I_10(I15679,I15628,I13761);
DFFARX1 I_11(I13746,I1470,I15611,,,I15928,);
not I_12(I16069,I16052);
endmodule


