module test_I10978(I1477,I10862,I9462,I9465,I1470,I10978);
input I1477,I10862,I9462,I9465,I1470;
output I10978;
wire I10879,I10647,I10961,I10664,I9720,I9737,I9471,I10715,I9542,I9771,I9459,I10896,I10749,I8178,I10732,I9754,I10913,I9621,I9689;
or I_0(I10879,I10862,I9462);
not I_1(I10647,I1477);
and I_2(I10978,I10961,I10913);
nand I_3(I10961,I10664,I9459);
not I_4(I10664,I9471);
not I_5(I9720,I9689);
nor I_6(I9737,I9621,I9720);
nor I_7(I9471,I9689,I9542);
nor I_8(I10715,I10664);
DFFARX1 I_9(I1470,,,I9542,);
and I_10(I9771,I9754,I8178);
nand I_11(I9459,I9771,I9737);
DFFARX1 I_12(I10879,I1470,I10647,,,I10896,);
not I_13(I10749,I10732);
DFFARX1 I_14(I1470,,,I8178,);
nand I_15(I10732,I10715,I9465);
DFFARX1 I_16(I1470,,,I9754,);
nor I_17(I10913,I10896,I10749);
DFFARX1 I_18(I1470,,,I9621,);
DFFARX1 I_19(I1470,,,I9689,);
endmodule


