module test_I7731(I6826,I1477,I1470,I7731);
input I6826,I1477,I1470;
output I7731;
wire I6297,I7714,I6329,I6493,I6843;
DFFARX1 I_0(I6843,I1470,I6329,,,I6297,);
not I_1(I7714,I6297);
not I_2(I6329,I1477);
DFFARX1 I_3(I1470,I6329,,,I6493,);
and I_4(I6843,I6493,I6826);
not I_5(I7731,I7714);
endmodule


