module test_final(IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_11,blif_reset_net_1_r_11,G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11);
input IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_11,blif_reset_net_1_r_11;
output G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11;
wire G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1,N3_2_l_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1,n_431_0_l_11,n9_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11;
DFFARX1 I_0(n4_1_r_1,blif_clk_net_1_r_11,n9_11,G42_1_r_1,);
nor I_1(n_572_1_r_1,n26_1,n19_1);
nand I_2(n_573_1_r_1,n16_1,n18_1);
nor I_3(n_549_1_r_1,n20_1,n21_1);
nor I_4(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_5(G199_4_l_1,blif_clk_net_1_r_11,n9_11,ACVQN2_3_r_1,);
nor I_6(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_7(N1_4_r_1,blif_clk_net_1_r_11,n9_11,G199_4_r_1,);
DFFARX1 I_8(G199_4_l_1,blif_clk_net_1_r_11,n9_11,G214_4_r_1,);
and I_9(N3_2_l_1,IN_6_2_l_1,n23_1);
DFFARX1 I_10(N3_2_l_1,blif_clk_net_1_r_11,n9_11,n26_1,);
not I_11(n17_1,n26_1);
DFFARX1 I_12(IN_1_3_l_1,blif_clk_net_1_r_11,n9_11,n16_internal_1,);
not I_13(n16_1,n16_internal_1);
DFFARX1 I_14(IN_2_3_l_1,blif_clk_net_1_r_11,n9_11,ACVQN1_3_l_1,);
and I_15(N1_4_l_1,IN_6_4_l_1,n25_1);
DFFARX1 I_16(N1_4_l_1,blif_clk_net_1_r_11,n9_11,G199_4_l_1,);
DFFARX1 I_17(IN_3_4_l_1,blif_clk_net_1_r_11,n9_11,G214_4_l_1,);
nor I_18(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_19(G214_4_l_1,blif_clk_net_1_r_11,n9_11,n14_internal_1,);
not I_20(n14_1,n14_internal_1);
nor I_21(N1_4_r_1,n17_1,n24_1);
nand I_22(n18_1,IN_4_3_l_1,ACVQN1_3_l_1);
nor I_23(n19_1,IN_1_2_l_1,IN_3_2_l_1);
not I_24(n20_1,n18_1);
nor I_25(n21_1,n26_1,n22_1);
not I_26(n22_1,n19_1);
nand I_27(n23_1,IN_2_2_l_1,IN_3_2_l_1);
nor I_28(n24_1,n18_1,n22_1);
nand I_29(n25_1,IN_1_4_l_1,IN_2_4_l_1);
DFFARX1 I_30(n4_1_r_11,blif_clk_net_1_r_11,n9_11,G42_1_r_11,);
nor I_31(n_572_1_r_11,n29_11,n30_11);
nand I_32(n_573_1_r_11,n26_11,n28_11);
nor I_33(n_549_1_r_11,n27_11,n32_11);
nand I_34(n_569_1_r_11,n45_11,n28_11);
nor I_35(n_452_1_r_11,n43_11,n44_11);
nor I_36(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_37(N3_2_r_11,blif_clk_net_1_r_11,n9_11,G199_2_r_11,);
DFFARX1 I_38(n24_11,blif_clk_net_1_r_11,n9_11,ACVQN2_3_r_11,);
nor I_39(n_266_and_0_3_r_11,n20_11,n37_11);
or I_40(n_431_0_l_11,n33_11,G199_4_r_1);
not I_41(n9_11,blif_reset_net_1_r_11);
DFFARX1 I_42(n_431_0_l_11,blif_clk_net_1_r_11,n9_11,n43_11,);
not I_43(n26_11,n43_11);
DFFARX1 I_44(G42_1_r_1,blif_clk_net_1_r_11,n9_11,n44_11,);
DFFARX1 I_45(n_452_1_r_1,blif_clk_net_1_r_11,n9_11,n45_11,);
not I_46(n27_11,n45_11);
nor I_47(n4_1_r_11,n44_11,n25_11);
nor I_48(N3_2_r_11,n45_11,n40_11);
nand I_49(n24_11,n39_11,ACVQN2_3_r_1);
nand I_50(n25_11,n38_11,G42_1_r_1);
DFFARX1 I_51(n25_11,blif_clk_net_1_r_11,n9_11,n20_internal_11,);
not I_52(n20_11,n20_internal_11);
not I_53(n28_11,n25_11);
not I_54(n29_11,n_266_and_0_3_r_1);
nand I_55(n30_11,n26_11,n31_11);
not I_56(n31_11,n_549_1_r_1);
and I_57(n32_11,n26_11,n44_11);
and I_58(n33_11,n34_11,G214_4_r_1);
nor I_59(n34_11,n29_11,n_572_1_r_1);
not I_60(n35_11,n_573_1_r_1);
nand I_61(n36_11,n31_11,n_266_and_0_3_r_1);
nor I_62(n37_11,n29_11,n_549_1_r_1);
nor I_63(n38_11,n31_11,n_573_1_r_1);
nor I_64(n39_11,n_572_1_r_1,n_573_1_r_1);
nor I_65(n40_11,n41_11,n_573_1_r_1);
nor I_66(n41_11,n42_11,n_572_1_r_1);
not I_67(n42_11,ACVQN2_3_r_1);
endmodule


