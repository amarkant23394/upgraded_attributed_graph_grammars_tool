module test_I1784(I1439,I1477,I1215,I1423,I1279,I1470,I1716,I1535,I1784);
input I1439,I1477,I1215,I1423,I1279,I1470,I1716,I1535;
output I1784;
wire I1518,I1750,I1733,I1586,I1603,I1620,I1767;
not I_0(I1518,I1477);
or I_1(I1750,I1733,I1279);
and I_2(I1733,I1716,I1439);
nor I_3(I1784,I1767,I1620);
nor I_4(I1586,I1535,I1215);
nand I_5(I1603,I1586,I1423);
not I_6(I1620,I1603);
DFFARX1 I_7(I1750,I1470,I1518,,,I1767,);
endmodule


