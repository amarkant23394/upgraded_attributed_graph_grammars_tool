module test_I1526(I1271,I1231,I1207,I1526);
input I1271,I1231,I1207;
output I1526;
wire I1492,I1509;
not I_0(I1492,I1207);
and I_1(I1526,I1509,I1271);
nor I_2(I1509,I1492,I1231);
endmodule


