module test_I5105_rst(I1477_rst,I5105_rst);
,I5105_rst);
input I1477_rst;
output I5105_rst;
wire ;
not I_0(I5105_rst,I1477_rst);
endmodule


