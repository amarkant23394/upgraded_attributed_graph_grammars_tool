module test_I1475(I1215,I1475);
input I1215;
output I1475;
wire ;
not I_0(I1475,I1215);
endmodule


