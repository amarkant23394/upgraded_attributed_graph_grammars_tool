module test_I12157(I7621,I1477,I7850,I1470,I10202,I12157);
input I7621,I1477,I7850,I1470,I10202;
output I12157;
wire I7556,I12140,I10219,I10014,I10490,I10052,I10035;
nand I_0(I7556,I7621,I7850);
not I_1(I12140,I10014);
DFFARX1 I_2(I10202,I1470,I10052,,,I10219,);
DFFARX1 I_3(I10219,I1470,I10052,,,I10014,);
nor I_4(I12157,I12140,I10035);
DFFARX1 I_5(I7556,I1470,I10052,,,I10490,);
not I_6(I10052,I1477);
not I_7(I10035,I10490);
endmodule


