module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_16,blif_reset_net_1_r_16,G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_16,blif_reset_net_1_r_16;
output G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n4_1_l_16,n7_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_16,n7_16,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_16,n7_16,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_16,n7_16,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_16,n7_16,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_16,n7_16,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_16,n7_16,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_16,n7_16,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_16,n7_16,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_16,n7_16,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_16,blif_clk_net_1_r_16,n7_16,G42_1_r_16,);
nor I_34(n_572_1_r_16,n20_16,n21_16);
nand I_35(n_573_1_r_16,n18_16,n19_16);
nor I_36(n_549_1_r_16,n23_16,n24_16);
nand I_37(n_569_1_r_16,n18_16,n22_16);
nor I_38(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_39(N1_4_r_16,blif_clk_net_1_r_16,n7_16,G199_4_r_16,);
DFFARX1 I_40(n6_16,blif_clk_net_1_r_16,n7_16,G214_4_r_16,);
DFFARX1 I_41(n_573_1_l_16,blif_clk_net_1_r_16,n7_16,ACVQN1_5_r_16,);
not I_42(P6_5_r_16,P6_5_r_internal_16);
nor I_43(n4_1_l_16,n_573_1_r_9,G214_4_r_9);
not I_44(n7_16,blif_reset_net_1_r_16);
DFFARX1 I_45(n4_1_l_16,blif_clk_net_1_r_16,n7_16,n29_16,);
DFFARX1 I_46(G199_4_r_9,blif_clk_net_1_r_16,n7_16,n16_internal_16,);
not I_47(n16_16,n16_internal_16);
DFFARX1 I_48(G199_2_r_9,blif_clk_net_1_r_16,n7_16,ACVQN1_3_l_16,);
nor I_49(n4_1_r_16,n29_16,n21_16);
nor I_50(N1_4_r_16,n27_16,n28_16);
not I_51(n6_16,n19_16);
or I_52(n_573_1_l_16,n_569_1_r_9,G42_1_r_9);
nor I_53(n_452_1_l_16,n_573_1_r_9,n_569_1_r_9);
DFFARX1 I_54(n_452_1_l_16,blif_clk_net_1_r_16,n7_16,P6_5_r_internal_16,);
not I_55(n18_16,n20_16);
nor I_56(n19_16,n_42_2_r_9,G42_1_r_9);
nor I_57(n20_16,n_549_1_r_9,n_572_1_r_9);
nor I_58(n21_16,n25_16,n_42_2_r_9);
nand I_59(n22_16,ACVQN1_3_l_16,n_572_1_r_9);
not I_60(n23_16,n22_16);
nor I_61(n24_16,n16_16,n20_16);
nor I_62(n25_16,n26_16,n_549_1_r_9);
not I_63(n26_16,G42_1_r_9);
and I_64(n27_16,n29_16,G42_1_r_9);
not I_65(n28_16,n_452_1_l_16);
endmodule


