module test_I11559(I11491,I1477,I9083,I8981,I1470,I6896,I11559);
input I11491,I1477,I9083,I8981,I1470,I6896;
output I11559;
wire I8824,I11542,I11508,I8842,I11525,I8833,I9179,I8862,I11310;
nand I_0(I8824,I9083,I8981);
or I_1(I11542,I11525,I8833);
nor I_2(I11508,I11491,I8842);
nor I_3(I8842,I9083);
and I_4(I11525,I11508,I8824);
not I_5(I8833,I9179);
DFFARX1 I_6(I6896,I1470,I8862,,,I9179,);
not I_7(I8862,I1477);
DFFARX1 I_8(I11542,I1470,I11310,,,I11559,);
not I_9(I11310,I1477);
endmodule


