module Benchmark_testing45000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2507,I2514,I56747,I56759,I56768,I56771,I56756,I56765,I56753,I56762,I56750,I78881,I78893,I78902,I78905,I78890,I78899,I78887,I78896,I78884,I123513,I123489,I123501,I123495,I123510,I123504,I123498,I123492,I123507,I124703,I124679,I124691,I124685,I124700,I124694,I124688,I124682,I124697,I173234,I173258,I173240,I173243,I173231,I173249,I173252,I173237,I173246,I173255,I242771,I242750,I242744,I242759,I242747,I242762,I242753,I242756,I242768,I242765,I307957,I307954,I307945,I307948,I307942,I307951,I307939,I307963,I307960,I371534,I371537,I371519,I371528,I371540,I371531,I371522,I371525,I371543,I471344,I471347,I471338,I471329,I471332,I471341,I471326,I471335,I549224,I549206,I549209,I549218,I549221,I549215,I549203,I549212,I639293,I639272,I639275,I639290,I639287,I639284,I639281,I639269,I639278,I678087,I678066,I678072,I678081,I678084,I678063,I678078,I678075,I678069,I718611,I718626,I718608,I718620,I718635,I718632,I718629,I718623,I718617,I718614);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2507,I2514;
output I56747,I56759,I56768,I56771,I56756,I56765,I56753,I56762,I56750,I78881,I78893,I78902,I78905,I78890,I78899,I78887,I78896,I78884,I123513,I123489,I123501,I123495,I123510,I123504,I123498,I123492,I123507,I124703,I124679,I124691,I124685,I124700,I124694,I124688,I124682,I124697,I173234,I173258,I173240,I173243,I173231,I173249,I173252,I173237,I173246,I173255,I242771,I242750,I242744,I242759,I242747,I242762,I242753,I242756,I242768,I242765,I307957,I307954,I307945,I307948,I307942,I307951,I307939,I307963,I307960,I371534,I371537,I371519,I371528,I371540,I371531,I371522,I371525,I371543,I471344,I471347,I471338,I471329,I471332,I471341,I471326,I471335,I549224,I549206,I549209,I549218,I549221,I549215,I549203,I549212,I639293,I639272,I639275,I639290,I639287,I639284,I639281,I639269,I639278,I678087,I678066,I678072,I678081,I678084,I678063,I678078,I678075,I678069,I718611,I718626,I718608,I718620,I718635,I718632,I718629,I718623,I718617,I718614;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2507,I2514,I2546,I399865,I2572,I2580,I399844,I2597,I2538,I399853,I2637,I2645,I2662,I399859,I2679,I399856,I2696,I2713,I2517,I2744,I2761,I2778,I399847,I399841,I2520,I2809,I2826,I399862,I2843,I2860,I2877,I2894,I2529,I2925,I399850,I2942,I2959,I2535,I2990,I2532,I3021,I3047,I3055,I3072,I2526,I2523,I3141,I567722,I3167,I3175,I567734,I3192,I3133,I567719,I3232,I3240,I3257,I3274,I567716,I3291,I3308,I3112,I3339,I3356,I3373,I567725,I3115,I3404,I3421,I567731,I3438,I3455,I3472,I3489,I3124,I3520,I567728,I3537,I3554,I3130,I3585,I3127,I3616,I567737,I3642,I3650,I3667,I3121,I3118,I3736,I628902,I3762,I3770,I3787,I3728,I628917,I3827,I3835,I3852,I628914,I3869,I628923,I3886,I3903,I3707,I3934,I3951,I3968,I628911,I628920,I3710,I3999,I4016,I628908,I4033,I628899,I4050,I4067,I4084,I3719,I4115,I628905,I4132,I4149,I3725,I4180,I3722,I4211,I4237,I4245,I4262,I3716,I3713,I4331,I577460,I4357,I4365,I4382,I4323,I577475,I4422,I4430,I4447,I577472,I4464,I577481,I4481,I4498,I4302,I4529,I4546,I4563,I577469,I577478,I4305,I4594,I4611,I577466,I4628,I577457,I4645,I4662,I4679,I4314,I4710,I577463,I4727,I4744,I4320,I4775,I4317,I4806,I4832,I4840,I4857,I4311,I4308,I4926,I457633,I4952,I4960,I457624,I4977,I4918,I457630,I5017,I5025,I5042,I5059,I457636,I5076,I5093,I4897,I5124,I5141,I5158,I457645,I457642,I4900,I5189,I5206,I5223,I457627,I5240,I5257,I5274,I4909,I5305,I5322,I5339,I4915,I5370,I4912,I5401,I457639,I5427,I5435,I5452,I4906,I4903,I5521,I456052,I5547,I5555,I456043,I5572,I5513,I456049,I5612,I5620,I5637,I5654,I456055,I5671,I5688,I5492,I5719,I5736,I5753,I456064,I456061,I5495,I5784,I5801,I5818,I456046,I5835,I5852,I5869,I5504,I5900,I5917,I5934,I5510,I5965,I5507,I5996,I456058,I6022,I6030,I6047,I5501,I5498,I6116,I489299,I6142,I6150,I489290,I6167,I6108,I489293,I6207,I6215,I6232,I489305,I6249,I489284,I6266,I6283,I6087,I6314,I6331,I6348,I489296,I489302,I6090,I6379,I6396,I489287,I6413,I489278,I6430,I6447,I6464,I6099,I6495,I6512,I6529,I6105,I6560,I6102,I6591,I489281,I6617,I6625,I6642,I6096,I6093,I6714,I501576,I6740,I6757,I6765,I6782,I501552,I501579,I6799,I501564,I6825,I6706,I6697,I501570,I6870,I6878,I501555,I6895,I6694,I501573,I6935,I6943,I6700,I6688,I6988,I501558,I501561,I7005,I7031,I7039,I6682,I7070,I7087,I501567,I7104,I7121,I7138,I6703,I7169,I6691,I6685,I7241,I591931,I7267,I7284,I7292,I7309,I591919,I591910,I7326,I591907,I7352,I7233,I7224,I591913,I7397,I7405,I591925,I7422,I7221,I591922,I7462,I7470,I7227,I7215,I7515,I591916,I7532,I591928,I7558,I7566,I7209,I7597,I7614,I7631,I7648,I7665,I7230,I7696,I7218,I7212,I7768,I517080,I7794,I7811,I7819,I7836,I517056,I517083,I7853,I517068,I7879,I7760,I7751,I517074,I7924,I7932,I517059,I7949,I7748,I517077,I7989,I7997,I7754,I7742,I8042,I517062,I517065,I8059,I8085,I8093,I7736,I8124,I8141,I517071,I8158,I8175,I8192,I7757,I8223,I7745,I7739,I8295,I225431,I8321,I8338,I8346,I8363,I225428,I225422,I8380,I225416,I8406,I8287,I8278,I225404,I8451,I8459,I225413,I8476,I8275,I225410,I8516,I8524,I8281,I8269,I8569,I225407,I225425,I8586,I8612,I8620,I8263,I8651,I8668,I225419,I8685,I8702,I8719,I8284,I8750,I8272,I8266,I8822,I667096,I8848,I8865,I8873,I8890,I667099,I667093,I8907,I667102,I8933,I8814,I8805,I667090,I8978,I8986,I667105,I9003,I8802,I667081,I9043,I9051,I8808,I8796,I9096,I667084,I9113,I9139,I9147,I8790,I9178,I9195,I667087,I9212,I9229,I9246,I8811,I9277,I8799,I8793,I9349,I646885,I9375,I9392,I9400,I9417,I646903,I646897,I9434,I646906,I9460,I9341,I9332,I646891,I9505,I9513,I646900,I9530,I9329,I646888,I9570,I9578,I9335,I9323,I9623,I646909,I646894,I9640,I9666,I9674,I9317,I9705,I9722,I9739,I9756,I9773,I9338,I9804,I9326,I9320,I9876,I140155,I9902,I9919,I9927,I9944,I140173,I140158,I9961,I140161,I9987,I9868,I9859,I140149,I10032,I10040,I140152,I10057,I9856,I140164,I10097,I10105,I9862,I9850,I10150,I140170,I140167,I10167,I10193,I10201,I9844,I10232,I10249,I10266,I10283,I10300,I9865,I10331,I9853,I9847,I10403,I722773,I10429,I10446,I10454,I10471,I722776,I722782,I10488,I722791,I10514,I10395,I10386,I722794,I10559,I10567,I722785,I10584,I10383,I10624,I10632,I10389,I10377,I10677,I722800,I722779,I10694,I722788,I10720,I10728,I10371,I10759,I10776,I722797,I10793,I10810,I10827,I10392,I10858,I10380,I10374,I10930,I589041,I10956,I10973,I10981,I10998,I589029,I589020,I11015,I589017,I11041,I10922,I10913,I589023,I11086,I11094,I589035,I11111,I10910,I589032,I11151,I11159,I10916,I10904,I11204,I589026,I11221,I589038,I11247,I11255,I10898,I11286,I11303,I11320,I11337,I11354,I10919,I11385,I10907,I10901,I11457,I11483,I11500,I11508,I11525,I11542,I11568,I11449,I11440,I11613,I11621,I11638,I11437,I11678,I11686,I11443,I11431,I11731,I11748,I11774,I11782,I11425,I11813,I11830,I11847,I11864,I11881,I11446,I11912,I11434,I11428,I11984,I266136,I12010,I12027,I12035,I12052,I266139,I12069,I266160,I12095,I11976,I11967,I266148,I12140,I12148,I266151,I12165,I11964,I266157,I12205,I12213,I11970,I11958,I12258,I266154,I266142,I12275,I266145,I12301,I12309,I11952,I12340,I12357,I266163,I12374,I12391,I12408,I11973,I12439,I11961,I11955,I12511,I585573,I12537,I12554,I12562,I12579,I585561,I585552,I12596,I585549,I12622,I12503,I12494,I585555,I12667,I12675,I585567,I12692,I12491,I585564,I12732,I12740,I12497,I12485,I12785,I585558,I12802,I585570,I12828,I12836,I12479,I12867,I12884,I12901,I12918,I12935,I12500,I12966,I12488,I12482,I13038,I641445,I13064,I13081,I13089,I13106,I641463,I641457,I13123,I641466,I13149,I13030,I13021,I641451,I13194,I13202,I641460,I13219,I13018,I641448,I13259,I13267,I13024,I13012,I13312,I641469,I641454,I13329,I13355,I13363,I13006,I13394,I13411,I13428,I13445,I13462,I13027,I13493,I13015,I13009,I13565,I261240,I13591,I13608,I13616,I13633,I261243,I13650,I261264,I13676,I13557,I13548,I261252,I13721,I13729,I261255,I13746,I13545,I261261,I13786,I13794,I13551,I13539,I13839,I261258,I261246,I13856,I261249,I13882,I13890,I13533,I13921,I13938,I261267,I13955,I13972,I13989,I13554,I14020,I13542,I13536,I14092,I711468,I14118,I14135,I14143,I14160,I711471,I711477,I14177,I711486,I14203,I14084,I14075,I711489,I14248,I14256,I711480,I14273,I14072,I14313,I14321,I14078,I14066,I14366,I711495,I711474,I14383,I711483,I14409,I14417,I14060,I14448,I14465,I711492,I14482,I14499,I14516,I14081,I14547,I14069,I14063,I14619,I220688,I14645,I14662,I14670,I14687,I220685,I220679,I14704,I220673,I14730,I14611,I14602,I220661,I14775,I14783,I220670,I14800,I14599,I220667,I14840,I14848,I14605,I14593,I14893,I220664,I220682,I14910,I14936,I14944,I14587,I14975,I14992,I220676,I15009,I15026,I15043,I14608,I15074,I14596,I14590,I15146,I195392,I15172,I15189,I15197,I15214,I195389,I195383,I15231,I195377,I15257,I15138,I15129,I195365,I15302,I15310,I195374,I15327,I15126,I195371,I15367,I15375,I15132,I15120,I15420,I195368,I195386,I15437,I15463,I15471,I15114,I15502,I15519,I195380,I15536,I15553,I15570,I15135,I15601,I15123,I15117,I15673,I594243,I15699,I15716,I15724,I15741,I594231,I594222,I15758,I594219,I15784,I15665,I15656,I594225,I15829,I15837,I594237,I15854,I15653,I594234,I15894,I15902,I15659,I15647,I15947,I594228,I15964,I594240,I15990,I15998,I15641,I16029,I16046,I16063,I16080,I16097,I15662,I16128,I15650,I15644,I16200,I44102,I16226,I16243,I16251,I16268,I44117,I16285,I44120,I16311,I16192,I16183,I44114,I16356,I16364,I44123,I16381,I16180,I44099,I16421,I16429,I16186,I16174,I16474,I44105,I16491,I44108,I16517,I16525,I16168,I16556,I16573,I44111,I16590,I16607,I16624,I16189,I16655,I16177,I16171,I16727,I364011,I16753,I16770,I16778,I16795,I364026,I364029,I16812,I364008,I16838,I16719,I16710,I364014,I16883,I16891,I364020,I16908,I16707,I16948,I16956,I16713,I16701,I17001,I364023,I364005,I17018,I364017,I17044,I17052,I16695,I17083,I17100,I17117,I17134,I17151,I16716,I17182,I16704,I16698,I17254,I580949,I17280,I17297,I17305,I17322,I580937,I580928,I17339,I580925,I17365,I17246,I17237,I580931,I17410,I17418,I580943,I17435,I17234,I580940,I17475,I17483,I17240,I17228,I17528,I580934,I17545,I580946,I17571,I17579,I17222,I17610,I17627,I17644,I17661,I17678,I17243,I17709,I17231,I17225,I17781,I679812,I17807,I17824,I17832,I17849,I679815,I679809,I17866,I679818,I17892,I17773,I17764,I679806,I17937,I17945,I679821,I17962,I17761,I679797,I18002,I18010,I17767,I17755,I18055,I679800,I18072,I18098,I18106,I17749,I18137,I18154,I679803,I18171,I18188,I18205,I17770,I18236,I17758,I17752,I18308,I704923,I18334,I18351,I18359,I18376,I704926,I704932,I18393,I704941,I18419,I18300,I18291,I704944,I18464,I18472,I704935,I18489,I18288,I18529,I18537,I18294,I18282,I18582,I704950,I704929,I18599,I704938,I18625,I18633,I18276,I18664,I18681,I704947,I18698,I18715,I18732,I18297,I18763,I18285,I18279,I18835,I287922,I18861,I18878,I18886,I18903,I287928,I287916,I18920,I287913,I18946,I18827,I18818,I287925,I18991,I18999,I287919,I19016,I18815,I287937,I19056,I19064,I18821,I18809,I19109,I287931,I287934,I19126,I19152,I19160,I18803,I19191,I19208,I19225,I19242,I19259,I18824,I19290,I18812,I18806,I19362,I38305,I19388,I19405,I19413,I19430,I38320,I19447,I38323,I19473,I19354,I19345,I38317,I19518,I19526,I38326,I19543,I19342,I38302,I19583,I19591,I19348,I19336,I19636,I38308,I19653,I38311,I19679,I19687,I19330,I19718,I19735,I38314,I19752,I19769,I19786,I19351,I19817,I19339,I19333,I19889,I588463,I19915,I19932,I19940,I19957,I588451,I588442,I19974,I588439,I20000,I19881,I19872,I588445,I20045,I20053,I588457,I20070,I19869,I588454,I20110,I20118,I19875,I19863,I20163,I588448,I20180,I588460,I20206,I20214,I19857,I20245,I20262,I20279,I20296,I20313,I19878,I20344,I19866,I19860,I20416,I48318,I20442,I20459,I20467,I20484,I48333,I20501,I48336,I20527,I20408,I20399,I48330,I20572,I20580,I48339,I20597,I20396,I48315,I20637,I20645,I20402,I20390,I20690,I48321,I20707,I48324,I20733,I20741,I20384,I20772,I20789,I48327,I20806,I20823,I20840,I20405,I20871,I20393,I20387,I20943,I243832,I20969,I20986,I20994,I21011,I243835,I21028,I243856,I21054,I20935,I20926,I243844,I21099,I21107,I243847,I21124,I20923,I243853,I21164,I21172,I20929,I20917,I21217,I243850,I243838,I21234,I243841,I21260,I21268,I20911,I21299,I21316,I243859,I21333,I21350,I21367,I20932,I21398,I20920,I20914,I21470,I403893,I21496,I21513,I21521,I21538,I403908,I403911,I21555,I403890,I21581,I21462,I21453,I403896,I21626,I21634,I403902,I21651,I21450,I21691,I21699,I21456,I21444,I21744,I403905,I403887,I21761,I403899,I21787,I21795,I21438,I21826,I21843,I21860,I21877,I21894,I21459,I21925,I21447,I21441,I21997,I540233,I22023,I22040,I22048,I22065,I540227,I540248,I22082,I22108,I21989,I21980,I540230,I22153,I22161,I540239,I22178,I21977,I22218,I22226,I21983,I21971,I22271,I540245,I22288,I540236,I22314,I22322,I21965,I22353,I22370,I540242,I22387,I22404,I22421,I21986,I22452,I21974,I21968,I22524,I605803,I22550,I22567,I22575,I22592,I605791,I605782,I22609,I605779,I22635,I22516,I22507,I605785,I22680,I22688,I605797,I22705,I22504,I605794,I22745,I22753,I22510,I22498,I22798,I605788,I22815,I605800,I22841,I22849,I22492,I22880,I22897,I22914,I22931,I22948,I22513,I22979,I22501,I22495,I23051,I182744,I23077,I23094,I23102,I23119,I182741,I182735,I23136,I182729,I23162,I23043,I23034,I182717,I23207,I23215,I182726,I23232,I23031,I182723,I23272,I23280,I23037,I23025,I23325,I182720,I182738,I23342,I23368,I23376,I23019,I23407,I23424,I182732,I23441,I23458,I23475,I23040,I23506,I23028,I23022,I23578,I332230,I23604,I23621,I23629,I23646,I332215,I332233,I23663,I332227,I23689,I23570,I23561,I332224,I23734,I23742,I23759,I23558,I332218,I23799,I23807,I23564,I23552,I23852,I332239,I332221,I23869,I332236,I23895,I23903,I23546,I23934,I23951,I23968,I23985,I24002,I23567,I24033,I23555,I23549,I24105,I58858,I24131,I24148,I24156,I24173,I58873,I24190,I58876,I24216,I24097,I24088,I58870,I24261,I24269,I58879,I24286,I24085,I58855,I24326,I24334,I24091,I24079,I24379,I58861,I24396,I58864,I24422,I24430,I24073,I24461,I24478,I58867,I24495,I24512,I24529,I24094,I24560,I24082,I24076,I24632,I612739,I24658,I24675,I24683,I24700,I612727,I612718,I24717,I612715,I24743,I24624,I24615,I612721,I24788,I24796,I612733,I24813,I24612,I612730,I24853,I24861,I24618,I24606,I24906,I612724,I24923,I612736,I24949,I24957,I24600,I24988,I25005,I25022,I25039,I25056,I24621,I25087,I24609,I24603,I25159,I531292,I25185,I25202,I25210,I25227,I531268,I531295,I25244,I531280,I25270,I25151,I25142,I531286,I25315,I25323,I531271,I25340,I25139,I531289,I25380,I25388,I25145,I25133,I25433,I531274,I531277,I25450,I25476,I25484,I25127,I25515,I25532,I531283,I25549,I25566,I25583,I25148,I25614,I25136,I25130,I25686,I568844,I25712,I25729,I25737,I25754,I568838,I568859,I25771,I25797,I25678,I25669,I568841,I25842,I25850,I568850,I25867,I25666,I25907,I25915,I25672,I25660,I25960,I568856,I25977,I568847,I26003,I26011,I25654,I26042,I26059,I568853,I26076,I26093,I26110,I25675,I26141,I25663,I25657,I26213,I26239,I26256,I26264,I26281,I26298,I26324,I26205,I26196,I26369,I26377,I26394,I26193,I26434,I26442,I26199,I26187,I26487,I26504,I26530,I26538,I26181,I26569,I26586,I26603,I26620,I26637,I26202,I26668,I26190,I26184,I26740,I443404,I26766,I26783,I26791,I26808,I443395,I443416,I26825,I443398,I26851,I26732,I26723,I26896,I26904,I443413,I26921,I26720,I443407,I26961,I26969,I26726,I26714,I27014,I443401,I443410,I27031,I27057,I27065,I26708,I27096,I27113,I27130,I27147,I27164,I26729,I27195,I26717,I26711,I27267,I209621,I27293,I27310,I27318,I27335,I209618,I209612,I27352,I209606,I27378,I27259,I27250,I209594,I27423,I27431,I209603,I27448,I27247,I209600,I27488,I27496,I27253,I27241,I27541,I209597,I209615,I27558,I27584,I27592,I27235,I27623,I27640,I209609,I27657,I27674,I27691,I27256,I27722,I27244,I27238,I27794,I652325,I27820,I27837,I27845,I27862,I652343,I652337,I27879,I652346,I27905,I27786,I27777,I652331,I27950,I27958,I652340,I27975,I27774,I652328,I28015,I28023,I27780,I27768,I28068,I652349,I652334,I28085,I28111,I28119,I27762,I28150,I28167,I28184,I28201,I28218,I27783,I28249,I27771,I27765,I28321,I94340,I28347,I28364,I28372,I28389,I94358,I94343,I28406,I94346,I28432,I28313,I28304,I94334,I28477,I28485,I94337,I28502,I28301,I94349,I28542,I28550,I28307,I28295,I28595,I94355,I94352,I28612,I28638,I28646,I28289,I28677,I28694,I28711,I28728,I28745,I28310,I28776,I28298,I28292,I28848,I299227,I28874,I28891,I28899,I28916,I299233,I299221,I28933,I299218,I28959,I28840,I28831,I299230,I29004,I29012,I299224,I29029,I28828,I299242,I29069,I29077,I28834,I28822,I29122,I299236,I299239,I29139,I29165,I29173,I28816,I29204,I29221,I29238,I29255,I29272,I28837,I29303,I28825,I28819,I29375,I155030,I29401,I29418,I29426,I29443,I155048,I155033,I29460,I155036,I29486,I29367,I29358,I155024,I29531,I29539,I155027,I29556,I29355,I155039,I29596,I29604,I29361,I29349,I29649,I155045,I155042,I29666,I29692,I29700,I29343,I29731,I29748,I29765,I29782,I29799,I29364,I29830,I29352,I29346,I29902,I317202,I29928,I29945,I29953,I29970,I317187,I317205,I29987,I317199,I30013,I29894,I29885,I317196,I30058,I30066,I30083,I29882,I317190,I30123,I30131,I29888,I29876,I30176,I317211,I317193,I30193,I317208,I30219,I30227,I29870,I30258,I30275,I30292,I30309,I30326,I29891,I30357,I29879,I29873,I30429,I528708,I30455,I30472,I30480,I30497,I528684,I528711,I30514,I528696,I30540,I30421,I30412,I528702,I30585,I30593,I528687,I30610,I30409,I528705,I30650,I30658,I30415,I30403,I30703,I528690,I528693,I30720,I30746,I30754,I30397,I30785,I30802,I528699,I30819,I30836,I30853,I30418,I30884,I30406,I30400,I30956,I497700,I30982,I30999,I31007,I31024,I497676,I497703,I31041,I497688,I31067,I30948,I30939,I497694,I31112,I31120,I497679,I31137,I30936,I497697,I31177,I31185,I30942,I30930,I31230,I497682,I497685,I31247,I31273,I31281,I30924,I31312,I31329,I497691,I31346,I31363,I31380,I30945,I31411,I30933,I30927,I31483,I621409,I31509,I31526,I31534,I31551,I621397,I621388,I31568,I621385,I31594,I31475,I31466,I621391,I31639,I31647,I621403,I31664,I31463,I621400,I31704,I31712,I31469,I31457,I31757,I621394,I31774,I621406,I31800,I31808,I31451,I31839,I31856,I31873,I31890,I31907,I31472,I31938,I31460,I31454,I32010,I684428,I32036,I32053,I32061,I32078,I684419,I684425,I32095,I684404,I32121,I32002,I31993,I684422,I32166,I32174,I32191,I31990,I684416,I32231,I32239,I31996,I31984,I32284,I684410,I684431,I32301,I684413,I32327,I32335,I31978,I32366,I32383,I684407,I32400,I32417,I32434,I31999,I32465,I31987,I31981,I32537,I700758,I32563,I32580,I32588,I32605,I700761,I700767,I32622,I700776,I32648,I32529,I32520,I700779,I32693,I32701,I700770,I32718,I32517,I32758,I32766,I32523,I32511,I32811,I700785,I700764,I32828,I700773,I32854,I32862,I32505,I32893,I32910,I700782,I32927,I32944,I32961,I32526,I32992,I32514,I32508,I33064,I512558,I33090,I33107,I33115,I33132,I512534,I512561,I33149,I512546,I33175,I33056,I33047,I512552,I33220,I33228,I512537,I33245,I33044,I512555,I33285,I33293,I33050,I33038,I33338,I512540,I512543,I33355,I33381,I33389,I33032,I33420,I33437,I512549,I33454,I33471,I33488,I33053,I33519,I33041,I33035,I33591,I686087,I33617,I33625,I33642,I686093,I686111,I33659,I686108,I33685,I686105,I33702,I33710,I686099,I33727,I33559,I33758,I33775,I33571,I33815,I33580,I33837,I686102,I686090,I33854,I686114,I33880,I33897,I33583,I33919,I33568,I33950,I686096,I33967,I33984,I34001,I33577,I34032,I33565,I33574,I33562,I34118,I633529,I34144,I34152,I34169,I633544,I633523,I34186,I633526,I34212,I633547,I34229,I34237,I34254,I34086,I34285,I34302,I34098,I34342,I34107,I34364,I633535,I633532,I34381,I633538,I34407,I34424,I34110,I34446,I34095,I34477,I633541,I34494,I34511,I34528,I34104,I34559,I34092,I34101,I34089,I34645,I221742,I34671,I34679,I34696,I221724,I221739,I34713,I221715,I34739,I221718,I34756,I34764,I221733,I34781,I34613,I34812,I34829,I34625,I221736,I34869,I34634,I34891,I221727,I34908,I221721,I34934,I34951,I34637,I34973,I34622,I35004,I221730,I35021,I35038,I35055,I34631,I35086,I34619,I34628,I34616,I35172,I35198,I35206,I35223,I35240,I35266,I35283,I35291,I35308,I35140,I35339,I35356,I35152,I35396,I35161,I35418,I35435,I35461,I35478,I35164,I35500,I35149,I35531,I35548,I35565,I35582,I35158,I35613,I35146,I35155,I35143,I35699,I658859,I35725,I35733,I35750,I658853,I658874,I35767,I658865,I35793,I658856,I35810,I35818,I658868,I35835,I35667,I35866,I35883,I35679,I35923,I35688,I35945,I658877,I658862,I35962,I35988,I36005,I35691,I36027,I35676,I36058,I658871,I36075,I36092,I36109,I35685,I36140,I35673,I35682,I35670,I36226,I36252,I36260,I36277,I36294,I36320,I36337,I36345,I36362,I36194,I36393,I36410,I36206,I36450,I36215,I36472,I36489,I36515,I36532,I36218,I36554,I36203,I36585,I36602,I36619,I36636,I36212,I36667,I36200,I36209,I36197,I36753,I154441,I36779,I36787,I36804,I154435,I154429,I36821,I154450,I36847,I154447,I36864,I36872,I154444,I36889,I36721,I36920,I36937,I36733,I36977,I36742,I36999,I154432,I37016,I154453,I37042,I37059,I36745,I37081,I36730,I37112,I154438,I37129,I37146,I37163,I36739,I37194,I36727,I36736,I36724,I37280,I158606,I37306,I37314,I37331,I158600,I158594,I37348,I158615,I37374,I158612,I37391,I37399,I158609,I37416,I37248,I37447,I37464,I37260,I37504,I37269,I37526,I158597,I37543,I158618,I37569,I37586,I37272,I37608,I37257,I37639,I158603,I37656,I37673,I37690,I37266,I37721,I37254,I37263,I37251,I37807,I224377,I37833,I37841,I37858,I224359,I224374,I37875,I224350,I37901,I224353,I37918,I37926,I224368,I37943,I37775,I37974,I37991,I37787,I224371,I38031,I37796,I38053,I224362,I38070,I224356,I38096,I38113,I37799,I38135,I37784,I38166,I224365,I38183,I38200,I38217,I37793,I38248,I37781,I37790,I37778,I38334,I314884,I38360,I38368,I38385,I314896,I314881,I38402,I314875,I38428,I314890,I38445,I38453,I314878,I38470,I38501,I38518,I314887,I38558,I38580,I314893,I314899,I38597,I38623,I38640,I38662,I38693,I38710,I38727,I38744,I38775,I38861,I337426,I38887,I38895,I38912,I337438,I337423,I38929,I337417,I38955,I337432,I38972,I38980,I337420,I38997,I38829,I39028,I39045,I38841,I337429,I39085,I38850,I39107,I337435,I337441,I39124,I39150,I39167,I38853,I39189,I38838,I39220,I39237,I39254,I39271,I38847,I39302,I38835,I38844,I38832,I39388,I478305,I39414,I39422,I39439,I478323,I478317,I39456,I478296,I39482,I478314,I39499,I39507,I478299,I39524,I39356,I39555,I39572,I39368,I478311,I39612,I39377,I39634,I478320,I478308,I39651,I478302,I39677,I39694,I39380,I39716,I39365,I39747,I39764,I39781,I39798,I39374,I39829,I39362,I39371,I39359,I39915,I102676,I39941,I39949,I39966,I102670,I102664,I39983,I102685,I40009,I102682,I40026,I40034,I102679,I40051,I39883,I40082,I40099,I39895,I40139,I39904,I40161,I102667,I40178,I102688,I40204,I40221,I39907,I40243,I39892,I40274,I102673,I40291,I40308,I40325,I39901,I40356,I39889,I39898,I39886,I40442,I105056,I40468,I40476,I40493,I105050,I105044,I40510,I105065,I40536,I105062,I40553,I40561,I105059,I40578,I40410,I40609,I40626,I40422,I40666,I40431,I40688,I105047,I40705,I105068,I40731,I40748,I40434,I40770,I40419,I40801,I105053,I40818,I40835,I40852,I40428,I40883,I40416,I40425,I40413,I40969,I366907,I40995,I41003,I41020,I366898,I366916,I41037,I366895,I41063,I41080,I41088,I366901,I41105,I40937,I41136,I41153,I40949,I41193,I40958,I41215,I366913,I366904,I41232,I366919,I41258,I41275,I40961,I41297,I40946,I41328,I366910,I41345,I41362,I41379,I40955,I41410,I40943,I40952,I40940,I41496,I112791,I41522,I41530,I41547,I112785,I112779,I41564,I112800,I41590,I112797,I41607,I41615,I112794,I41632,I41464,I41663,I41680,I41476,I41720,I41485,I41742,I112782,I41759,I112803,I41785,I41802,I41488,I41824,I41473,I41855,I112788,I41872,I41889,I41906,I41482,I41937,I41470,I41479,I41467,I42023,I199081,I42049,I42057,I42074,I199063,I199078,I42091,I199054,I42117,I199057,I42134,I42142,I199072,I42159,I41991,I42190,I42207,I42003,I199075,I42247,I42012,I42269,I199066,I42286,I199060,I42312,I42329,I42015,I42351,I42000,I42382,I199069,I42399,I42416,I42433,I42009,I42464,I41997,I42006,I41994,I42550,I189595,I42576,I42584,I42601,I189577,I189592,I42618,I189568,I42644,I189571,I42661,I42669,I189586,I42686,I42518,I42717,I42734,I42530,I189589,I42774,I42539,I42796,I189580,I42813,I189574,I42839,I42856,I42542,I42878,I42527,I42909,I189583,I42926,I42943,I42960,I42536,I42991,I42524,I42533,I42521,I43077,I587867,I43103,I43111,I43128,I587882,I587861,I43145,I587864,I43171,I587885,I43188,I43196,I43213,I43045,I43244,I43261,I43057,I43301,I43066,I43323,I587873,I587870,I43340,I587876,I43366,I43383,I43069,I43405,I43054,I43436,I587879,I43453,I43470,I43487,I43063,I43518,I43051,I43060,I43048,I43604,I342050,I43630,I43638,I43655,I342062,I342047,I43672,I342041,I43698,I342056,I43715,I43723,I342044,I43740,I43572,I43771,I43788,I43584,I342053,I43828,I43593,I43850,I342059,I342065,I43867,I43893,I43910,I43596,I43932,I43581,I43963,I43980,I43997,I44014,I43590,I44045,I43578,I43587,I43575,I44131,I365173,I44157,I44165,I44182,I365164,I365182,I44199,I365161,I44225,I44242,I44250,I365167,I44267,I44298,I44315,I44355,I44377,I365179,I365170,I44394,I365185,I44420,I44437,I44459,I44490,I365176,I44507,I44524,I44541,I44572,I44658,I44684,I44692,I44709,I44726,I44752,I44769,I44777,I44794,I44626,I44825,I44842,I44638,I44882,I44647,I44904,I44921,I44947,I44964,I44650,I44986,I44635,I45017,I45034,I45051,I45068,I44644,I45099,I44632,I44641,I44629,I45185,I429175,I45211,I45219,I45236,I429172,I429187,I45253,I429169,I45279,I429166,I45296,I45304,I45321,I45153,I45352,I45369,I45165,I45409,I45174,I45431,I429181,I45448,I429184,I45474,I45491,I45177,I45513,I45162,I45544,I429178,I45561,I45578,I45595,I45171,I45626,I45159,I45168,I45156,I45712,I642539,I45738,I45746,I45763,I642533,I642554,I45780,I642545,I45806,I642536,I45823,I45831,I642548,I45848,I45680,I45879,I45896,I45692,I45936,I45701,I45958,I642557,I642542,I45975,I46001,I46018,I45704,I46040,I45689,I46071,I642551,I46088,I46105,I46122,I45698,I46153,I45686,I45695,I45683,I46239,I214891,I46265,I46273,I46290,I214873,I214888,I46307,I214864,I46333,I214867,I46350,I46358,I214882,I46375,I46207,I46406,I46423,I46219,I214885,I46463,I46228,I46485,I214876,I46502,I214870,I46528,I46545,I46231,I46567,I46216,I46598,I214879,I46615,I46632,I46649,I46225,I46680,I46213,I46222,I46210,I46766,I46792,I46800,I46817,I46834,I46860,I46877,I46885,I46902,I46734,I46933,I46950,I46746,I46990,I46755,I47012,I47029,I47055,I47072,I46758,I47094,I46743,I47125,I47142,I47159,I47176,I46752,I47207,I46740,I46749,I46737,I47293,I139566,I47319,I47327,I47344,I139560,I139554,I47361,I139575,I47387,I139572,I47404,I47412,I139569,I47429,I47261,I47460,I47477,I47273,I47517,I47282,I47539,I139557,I47556,I139578,I47582,I47599,I47285,I47621,I47270,I47652,I139563,I47669,I47686,I47703,I47279,I47734,I47267,I47276,I47264,I47820,I173785,I47846,I47854,I47871,I173767,I173782,I47888,I173758,I47914,I173761,I47931,I47939,I173776,I47956,I47788,I47987,I48004,I47800,I173779,I48044,I47809,I48066,I173770,I48083,I173764,I48109,I48126,I47812,I48148,I47797,I48179,I173773,I48196,I48213,I48230,I47806,I48261,I47794,I47803,I47791,I48347,I372109,I48373,I48381,I48398,I372100,I372118,I48415,I372097,I48441,I48458,I48466,I372103,I48483,I48514,I48531,I48571,I48593,I372115,I372106,I48610,I372121,I48636,I48653,I48675,I48706,I372112,I48723,I48740,I48757,I48788,I48874,I48900,I48908,I48925,I48942,I48968,I48985,I48993,I49010,I48842,I49041,I49058,I48854,I49098,I48863,I49120,I49137,I49163,I49180,I48866,I49202,I48851,I49233,I49250,I49267,I49284,I48860,I49315,I48848,I48857,I48845,I49401,I260170,I49427,I49435,I49452,I260164,I260155,I49469,I260176,I49495,I260158,I49512,I49520,I260152,I49537,I49369,I49568,I49585,I49381,I49625,I49390,I49647,I260179,I260161,I49664,I260167,I49690,I49707,I49393,I49729,I49378,I49760,I260173,I49777,I49794,I49811,I49387,I49842,I49375,I49384,I49372,I49928,I666524,I49954,I49962,I49979,I666527,I666521,I49996,I666518,I50022,I666503,I50039,I50047,I666512,I50064,I49896,I50095,I50112,I49908,I50152,I49917,I50174,I666506,I666509,I50191,I666515,I50217,I50234,I49920,I50256,I49905,I50287,I50304,I50321,I50338,I49914,I50369,I49902,I49911,I49899,I50455,I597693,I50481,I50489,I50506,I597708,I597687,I50523,I597690,I50549,I597711,I50566,I50574,I50591,I50423,I50622,I50639,I50435,I50679,I50444,I50701,I597699,I597696,I50718,I597702,I50744,I50761,I50447,I50783,I50432,I50814,I597705,I50831,I50848,I50865,I50441,I50896,I50429,I50438,I50426,I50982,I111601,I51008,I51016,I51033,I111595,I111589,I51050,I111610,I51076,I111607,I51093,I51101,I111604,I51118,I50950,I51149,I51166,I50962,I51206,I50971,I51228,I111592,I51245,I111613,I51271,I51288,I50974,I51310,I50959,I51341,I111598,I51358,I51375,I51392,I50968,I51423,I50956,I50965,I50953,I51509,I97916,I51535,I51543,I51560,I97910,I97904,I51577,I97925,I51603,I97922,I51620,I51628,I97919,I51645,I51477,I51676,I51693,I51489,I51733,I51498,I51755,I97907,I51772,I97928,I51798,I51815,I51501,I51837,I51486,I51868,I97913,I51885,I51902,I51919,I51495,I51950,I51483,I51492,I51480,I52036,I52062,I52070,I52087,I52104,I52130,I52147,I52155,I52172,I52004,I52203,I52220,I52016,I52260,I52025,I52282,I52299,I52325,I52342,I52028,I52364,I52013,I52395,I52412,I52429,I52446,I52022,I52477,I52010,I52019,I52007,I52563,I112196,I52589,I52597,I52614,I112190,I112184,I52631,I112205,I52657,I112202,I52674,I52682,I112199,I52699,I52531,I52730,I52747,I52543,I52787,I52552,I52809,I112187,I52826,I112208,I52852,I52869,I52555,I52891,I52540,I52922,I112193,I52939,I52956,I52973,I52549,I53004,I52537,I52546,I52534,I53090,I127666,I53116,I53124,I53141,I127660,I127654,I53158,I127675,I53184,I127672,I53201,I53209,I127669,I53226,I53058,I53257,I53274,I53070,I53314,I53079,I53336,I127657,I53353,I127678,I53379,I53396,I53082,I53418,I53067,I53449,I127663,I53466,I53483,I53500,I53076,I53531,I53064,I53073,I53061,I53617,I236234,I53643,I53651,I53668,I236228,I236219,I53685,I236240,I53711,I236222,I53728,I53736,I236216,I53753,I53585,I53784,I53801,I53597,I53841,I53606,I53863,I236243,I236225,I53880,I236231,I53906,I53923,I53609,I53945,I53594,I53976,I236237,I53993,I54010,I54027,I53603,I54058,I53591,I53600,I53588,I54144,I181163,I54170,I54178,I54195,I181145,I181160,I54212,I181136,I54238,I181139,I54255,I54263,I181154,I54280,I54112,I54311,I54328,I54124,I181157,I54368,I54133,I54390,I181148,I54407,I181142,I54433,I54450,I54136,I54472,I54121,I54503,I181151,I54520,I54537,I54554,I54130,I54585,I54118,I54127,I54115,I54671,I312572,I54697,I54705,I54722,I312584,I312569,I54739,I312563,I54765,I312578,I54782,I54790,I312566,I54807,I54639,I54838,I54855,I54651,I312575,I54895,I54660,I54917,I312581,I312587,I54934,I54960,I54977,I54663,I54999,I54648,I55030,I55047,I55064,I55081,I54657,I55112,I54645,I54654,I54642,I55198,I689465,I55224,I55232,I55249,I689459,I689480,I55266,I689456,I55292,I689477,I55309,I55317,I689474,I55334,I55166,I55365,I55382,I55178,I689462,I55422,I55187,I55444,I689471,I689468,I55461,I689453,I55487,I55504,I55190,I55526,I55175,I55557,I55574,I55591,I55608,I55184,I55639,I55172,I55181,I55169,I55725,I451836,I55751,I55759,I55776,I451833,I451848,I55793,I451830,I55819,I451827,I55836,I55844,I55861,I55693,I55892,I55909,I55705,I55949,I55714,I55971,I451842,I55988,I451845,I56014,I56031,I55717,I56053,I55702,I56084,I451839,I56101,I56118,I56135,I55711,I56166,I55699,I55708,I55696,I56252,I442877,I56278,I56286,I56303,I442874,I442889,I56320,I442871,I56346,I442868,I56363,I56371,I56388,I56220,I56419,I56436,I56232,I56476,I56241,I56498,I442883,I56515,I442886,I56541,I56558,I56244,I56580,I56229,I56611,I442880,I56628,I56645,I56662,I56238,I56693,I56226,I56235,I56223,I56779,I191703,I56805,I56813,I56830,I191685,I191700,I56847,I191676,I56873,I191679,I56890,I56898,I191694,I56915,I56946,I56963,I191697,I57003,I57025,I191688,I57042,I191682,I57068,I57085,I57107,I57138,I191691,I57155,I57172,I57189,I57220,I57306,I402165,I57332,I57340,I57357,I402156,I402174,I57374,I402153,I57400,I57417,I57425,I402159,I57442,I57274,I57473,I57490,I57286,I57530,I57295,I57552,I402171,I402162,I57569,I402177,I57595,I57612,I57298,I57634,I57283,I57665,I402168,I57682,I57699,I57716,I57292,I57747,I57280,I57289,I57277,I57833,I210675,I57859,I57867,I57884,I210657,I210672,I57901,I210648,I57927,I210651,I57944,I57952,I210666,I57969,I57801,I58000,I58017,I57813,I210669,I58057,I57822,I58079,I210660,I58096,I210654,I58122,I58139,I57825,I58161,I57810,I58192,I210663,I58209,I58226,I58243,I57819,I58274,I57807,I57816,I57804,I58360,I436553,I58386,I58394,I58411,I436550,I436565,I58428,I436547,I58454,I436544,I58471,I58479,I58496,I58328,I58527,I58544,I58340,I58584,I58349,I58606,I436559,I58623,I436562,I58649,I58666,I58352,I58688,I58337,I58719,I436556,I58736,I58753,I58770,I58346,I58801,I58334,I58343,I58331,I58887,I598849,I58913,I58921,I58938,I598864,I598843,I58955,I598846,I58981,I598867,I58998,I59006,I59023,I59054,I59071,I59111,I59133,I598855,I598852,I59150,I598858,I59176,I59193,I59215,I59246,I598861,I59263,I59280,I59297,I59328,I59414,I108626,I59440,I59448,I59465,I108620,I108614,I59482,I108635,I59508,I108632,I59525,I59533,I108629,I59550,I59382,I59581,I59598,I59394,I59638,I59403,I59660,I108617,I59677,I108638,I59703,I59720,I59406,I59742,I59391,I59773,I108623,I59790,I59807,I59824,I59400,I59855,I59388,I59397,I59385,I59941,I93751,I59967,I59975,I59992,I93745,I93739,I60009,I93760,I60035,I93757,I60052,I60060,I93754,I60077,I59909,I60108,I60125,I59921,I60165,I59930,I60187,I93742,I60204,I93763,I60230,I60247,I59933,I60269,I59918,I60300,I93748,I60317,I60334,I60351,I59927,I60382,I59915,I59924,I59912,I60468,I84835,I60494,I60502,I60519,I84832,I84814,I60536,I84820,I60562,I84829,I60579,I60587,I84823,I60604,I60436,I60635,I60652,I60448,I84838,I60692,I60457,I60714,I84826,I84817,I60731,I60757,I60774,I60460,I60796,I60445,I60827,I84841,I60844,I60861,I60878,I60454,I60909,I60442,I60451,I60439,I60995,I61021,I61029,I61046,I61063,I61089,I61106,I61114,I61131,I60963,I61162,I61179,I60975,I61219,I60984,I61241,I61258,I61284,I61301,I60987,I61323,I60972,I61354,I61371,I61388,I61405,I60981,I61436,I60969,I60978,I60966,I61522,I61548,I61556,I61573,I61590,I61616,I61633,I61641,I61658,I61490,I61689,I61706,I61502,I61746,I61511,I61768,I61785,I61811,I61828,I61514,I61850,I61499,I61881,I61898,I61915,I61932,I61508,I61963,I61496,I61505,I61493,I62049,I602317,I62075,I62083,I62100,I602332,I602311,I62117,I602314,I62143,I602335,I62160,I62168,I62185,I62017,I62216,I62233,I62029,I62273,I62038,I62295,I602323,I602320,I62312,I602326,I62338,I62355,I62041,I62377,I62026,I62408,I602329,I62425,I62442,I62459,I62035,I62490,I62023,I62032,I62020,I62576,I405055,I62602,I62610,I62627,I405046,I405064,I62644,I405043,I62670,I62687,I62695,I405049,I62712,I62544,I62743,I62760,I62556,I62800,I62565,I62822,I405061,I405052,I62839,I405067,I62865,I62882,I62568,I62904,I62553,I62935,I405058,I62952,I62969,I62986,I62562,I63017,I62550,I62559,I62547,I63103,I605207,I63129,I63137,I63154,I605222,I605201,I63171,I605204,I63197,I605225,I63214,I63222,I63239,I63071,I63270,I63287,I63083,I63327,I63092,I63349,I605213,I605210,I63366,I605216,I63392,I63409,I63095,I63431,I63080,I63462,I605219,I63479,I63496,I63513,I63089,I63544,I63077,I63086,I63074,I63630,I226485,I63656,I63664,I63681,I226467,I226482,I63698,I226458,I63724,I226461,I63741,I63749,I226476,I63766,I63598,I63797,I63814,I63610,I226479,I63854,I63619,I63876,I226470,I63893,I226464,I63919,I63936,I63622,I63958,I63607,I63989,I226473,I64006,I64023,I64040,I63616,I64071,I63604,I63613,I63601,I64157,I611565,I64183,I64191,I64208,I611580,I611559,I64225,I611562,I64251,I611583,I64268,I64276,I64293,I64125,I64324,I64341,I64137,I64381,I64146,I64403,I611571,I611568,I64420,I611574,I64446,I64463,I64149,I64485,I64134,I64516,I611577,I64533,I64550,I64567,I64143,I64598,I64131,I64140,I64128,I64684,I241674,I64710,I64718,I64735,I241668,I241659,I64752,I241680,I64778,I241662,I64795,I64803,I241656,I64820,I64652,I64851,I64868,I64664,I64908,I64673,I64930,I241683,I241665,I64947,I241671,I64973,I64990,I64676,I65012,I64661,I65043,I241677,I65060,I65077,I65094,I64670,I65125,I64658,I64667,I64655,I65211,I280842,I65237,I65245,I65262,I280836,I280827,I65279,I280848,I65305,I280830,I65322,I65330,I280824,I65347,I65179,I65378,I65395,I65191,I65435,I65200,I65457,I280851,I280833,I65474,I280839,I65500,I65517,I65203,I65539,I65188,I65570,I280845,I65587,I65604,I65621,I65197,I65652,I65185,I65194,I65182,I65738,I645259,I65764,I65772,I65789,I645253,I645274,I65806,I645265,I65832,I645256,I65849,I65857,I645268,I65874,I65706,I65905,I65922,I65718,I65962,I65727,I65984,I645277,I645262,I66001,I66027,I66044,I65730,I66066,I65715,I66097,I645271,I66114,I66131,I66148,I65724,I66179,I65712,I65721,I65709,I66265,I209094,I66291,I66299,I66316,I209076,I209091,I66333,I209067,I66359,I209070,I66376,I66384,I209085,I66401,I66233,I66432,I66449,I66245,I209088,I66489,I66254,I66511,I209079,I66528,I209073,I66554,I66571,I66257,I66593,I66242,I66624,I209082,I66641,I66658,I66675,I66251,I66706,I66239,I66248,I66236,I66792,I662667,I66818,I66826,I66843,I662661,I662682,I66860,I662673,I66886,I662664,I66903,I66911,I662676,I66928,I66760,I66959,I66976,I66772,I67016,I66781,I67038,I662685,I662670,I67055,I67081,I67098,I66784,I67120,I66769,I67151,I662679,I67168,I67185,I67202,I66778,I67233,I66766,I66775,I66763,I67319,I296246,I67345,I67353,I67370,I296267,I296261,I67387,I296243,I67413,I67430,I67438,I296255,I67455,I67287,I67486,I67503,I67299,I296252,I67543,I67308,I67565,I296258,I296249,I67582,I67608,I67625,I67311,I67647,I67296,I67678,I296264,I67695,I67712,I67729,I67305,I67760,I67293,I67302,I67290,I67846,I645803,I67872,I67880,I67897,I645797,I645818,I67914,I645809,I67940,I645800,I67957,I67965,I645812,I67982,I67814,I68013,I68030,I67826,I68070,I67835,I68092,I645821,I645806,I68109,I68135,I68152,I67838,I68174,I67823,I68205,I645815,I68222,I68239,I68256,I67832,I68287,I67820,I67829,I67817,I68373,I480889,I68399,I68407,I68424,I480907,I480901,I68441,I480880,I68467,I480898,I68484,I68492,I480883,I68509,I68341,I68540,I68557,I68353,I480895,I68597,I68362,I68619,I480904,I480892,I68636,I480886,I68662,I68679,I68365,I68701,I68350,I68732,I68749,I68766,I68783,I68359,I68814,I68347,I68356,I68344,I68900,I90181,I68926,I68934,I68951,I90175,I90169,I68968,I90190,I68994,I90187,I69011,I69019,I90184,I69036,I68868,I69067,I69084,I68880,I69124,I68889,I69146,I90172,I69163,I90193,I69189,I69206,I68892,I69228,I68877,I69259,I90178,I69276,I69293,I69310,I68886,I69341,I68874,I68883,I68871,I69427,I698390,I69453,I69461,I69478,I698384,I698405,I69495,I698381,I69521,I698402,I69538,I69546,I698399,I69563,I69395,I69594,I69611,I69407,I698387,I69651,I69416,I69673,I698396,I698393,I69690,I698378,I69716,I69733,I69419,I69755,I69404,I69786,I69803,I69820,I69837,I69413,I69868,I69401,I69410,I69398,I69954,I401009,I69980,I69988,I70005,I401000,I401018,I70022,I400997,I70048,I70065,I70073,I401003,I70090,I69922,I70121,I70138,I69934,I70178,I69943,I70200,I401015,I401006,I70217,I401021,I70243,I70260,I69946,I70282,I69931,I70313,I401012,I70330,I70347,I70364,I69940,I70395,I69928,I69937,I69925,I70481,I170096,I70507,I70515,I70532,I170078,I170093,I70549,I170069,I70575,I170072,I70592,I70600,I170087,I70617,I70449,I70648,I70665,I70461,I170090,I70705,I70470,I70727,I170081,I70744,I170075,I70770,I70787,I70473,I70809,I70458,I70840,I170084,I70857,I70874,I70891,I70467,I70922,I70455,I70464,I70452,I71008,I703745,I71034,I71042,I71059,I703739,I703760,I71076,I703736,I71102,I703757,I71119,I71127,I703754,I71144,I70976,I71175,I71192,I70988,I703742,I71232,I70997,I71254,I703751,I703748,I71271,I703733,I71297,I71314,I71000,I71336,I70985,I71367,I71384,I71401,I71418,I70994,I71449,I70982,I70991,I70979,I71535,I407367,I71561,I71569,I71586,I407358,I407376,I71603,I407355,I71629,I71646,I71654,I407361,I71671,I71503,I71702,I71719,I71515,I71759,I71524,I71781,I407373,I407364,I71798,I407379,I71824,I71841,I71527,I71863,I71512,I71894,I407370,I71911,I71928,I71945,I71521,I71976,I71509,I71518,I71506,I72062,I152656,I72088,I72096,I72113,I152650,I152644,I72130,I152665,I72156,I152662,I72173,I72181,I152659,I72198,I72030,I72229,I72246,I72042,I72286,I72051,I72308,I152647,I72325,I152668,I72351,I72368,I72054,I72390,I72039,I72421,I152653,I72438,I72455,I72472,I72048,I72503,I72036,I72045,I72033,I72589,I141946,I72615,I72623,I72640,I141940,I141934,I72657,I141955,I72683,I141952,I72700,I72708,I141949,I72725,I72557,I72756,I72773,I72569,I72813,I72578,I72835,I141937,I72852,I141958,I72878,I72895,I72581,I72917,I72566,I72948,I141943,I72965,I72982,I72999,I72575,I73030,I72563,I72572,I72560,I73116,I661579,I73142,I73150,I73167,I661573,I661594,I73184,I661585,I73210,I661576,I73227,I73235,I661588,I73252,I73084,I73283,I73300,I73096,I73340,I73105,I73362,I661597,I661582,I73379,I73405,I73422,I73108,I73444,I73093,I73475,I661591,I73492,I73509,I73526,I73102,I73557,I73090,I73099,I73087,I73643,I73669,I73677,I73694,I73711,I73737,I73754,I73762,I73779,I73611,I73810,I73827,I73623,I73867,I73632,I73889,I73906,I73932,I73949,I73635,I73971,I73620,I74002,I74019,I74036,I74053,I73629,I74084,I73617,I73626,I73614,I74170,I358237,I74196,I74204,I74221,I358228,I358246,I74238,I358225,I74264,I74281,I74289,I358231,I74306,I74138,I74337,I74354,I74150,I74394,I74159,I74416,I358243,I358234,I74433,I358249,I74459,I74476,I74162,I74498,I74147,I74529,I358240,I74546,I74563,I74580,I74156,I74611,I74144,I74153,I74141,I74697,I493163,I74723,I74731,I74748,I493181,I493175,I74765,I493154,I74791,I493172,I74808,I74816,I493157,I74833,I74665,I74864,I74881,I74677,I493169,I74921,I74686,I74943,I493178,I493166,I74960,I493160,I74986,I75003,I74689,I75025,I74674,I75056,I75073,I75090,I75107,I74683,I75138,I74671,I74680,I74668,I75224,I265066,I75250,I75258,I75275,I265060,I265051,I75292,I265072,I75318,I265054,I75335,I75343,I265048,I75360,I75192,I75391,I75408,I75204,I75448,I75213,I75470,I265075,I265057,I75487,I265063,I75513,I75530,I75216,I75552,I75201,I75583,I265069,I75600,I75617,I75634,I75210,I75665,I75198,I75207,I75195,I75751,I386559,I75777,I75785,I75802,I386550,I386568,I75819,I386547,I75845,I75862,I75870,I386553,I75887,I75719,I75918,I75935,I75731,I75975,I75740,I75997,I386565,I386556,I76014,I386571,I76040,I76057,I75743,I76079,I75728,I76110,I386562,I76127,I76144,I76161,I75737,I76192,I75725,I75734,I75722,I76278,I701365,I76304,I76312,I76329,I701359,I701380,I76346,I701356,I76372,I701377,I76389,I76397,I701374,I76414,I76246,I76445,I76462,I76258,I701362,I76502,I76267,I76524,I701371,I701368,I76541,I701353,I76567,I76584,I76270,I76606,I76255,I76637,I76654,I76671,I76688,I76264,I76719,I76252,I76261,I76249,I76805,I125881,I76831,I76839,I76856,I125875,I125869,I76873,I125890,I76899,I125887,I76916,I76924,I125884,I76941,I76773,I76972,I76989,I76785,I77029,I76794,I77051,I125872,I77068,I125893,I77094,I77111,I76797,I77133,I76782,I77164,I125878,I77181,I77198,I77215,I76791,I77246,I76779,I76788,I76776,I77332,I388871,I77358,I77366,I77383,I388862,I388880,I77400,I388859,I77426,I77443,I77451,I388865,I77468,I77300,I77499,I77516,I77312,I77556,I77321,I77578,I388877,I388868,I77595,I388883,I77621,I77638,I77324,I77660,I77309,I77691,I388874,I77708,I77725,I77742,I77318,I77773,I77306,I77315,I77303,I77859,I172204,I77885,I77893,I77910,I172186,I172201,I77927,I172177,I77953,I172180,I77970,I77978,I172195,I77995,I77827,I78026,I78043,I77839,I172198,I78083,I77848,I78105,I172189,I78122,I172183,I78148,I78165,I77851,I78187,I77836,I78218,I172192,I78235,I78252,I78269,I77845,I78300,I77833,I77842,I77830,I78386,I216999,I78412,I78420,I78437,I216981,I216996,I78454,I216972,I78480,I216975,I78497,I78505,I216990,I78522,I78354,I78553,I78570,I78366,I216993,I78610,I78375,I78632,I216984,I78649,I216978,I78675,I78692,I78378,I78714,I78363,I78745,I216987,I78762,I78779,I78796,I78372,I78827,I78360,I78369,I78357,I78913,I661035,I78939,I78947,I78964,I661029,I661050,I78981,I661041,I79007,I661032,I79024,I79032,I661044,I79049,I79080,I79097,I79137,I79159,I661053,I661038,I79176,I79202,I79219,I79241,I79272,I661047,I79289,I79306,I79323,I79354,I79440,I616767,I79466,I79474,I79491,I616782,I616761,I79508,I616764,I79534,I616785,I79551,I79559,I79576,I79408,I79607,I79624,I79420,I79664,I79429,I79686,I616773,I616770,I79703,I616776,I79729,I79746,I79432,I79768,I79417,I79799,I616779,I79816,I79833,I79850,I79426,I79881,I79414,I79423,I79411,I79967,I79993,I80001,I80018,I80035,I80061,I80078,I80086,I80103,I79935,I80134,I80151,I79947,I80191,I79956,I80213,I80230,I80256,I80273,I79959,I80295,I79944,I80326,I80343,I80360,I80377,I79953,I80408,I79941,I79950,I79938,I80494,I582665,I80520,I80528,I80545,I582680,I582659,I80562,I582662,I80588,I582683,I80605,I80613,I80630,I80462,I80661,I80678,I80474,I80718,I80483,I80740,I582671,I582668,I80757,I582674,I80783,I80800,I80486,I80822,I80471,I80853,I582677,I80870,I80887,I80904,I80480,I80935,I80468,I80477,I80465,I81021,I183271,I81047,I81055,I81072,I183253,I183268,I81089,I183244,I81115,I183247,I81132,I81140,I183262,I81157,I80989,I81188,I81205,I81001,I183265,I81245,I81010,I81267,I183256,I81284,I183250,I81310,I81327,I81013,I81349,I80998,I81380,I183259,I81397,I81414,I81431,I81007,I81462,I80995,I81004,I80992,I81548,I470808,I81574,I81582,I81599,I470805,I470820,I81616,I470802,I81642,I470799,I81659,I81667,I81684,I81516,I81715,I81732,I81528,I81772,I81537,I81794,I470814,I81811,I470817,I81837,I81854,I81540,I81876,I81525,I81907,I470811,I81924,I81941,I81958,I81534,I81989,I81522,I81531,I81519,I82075,I457106,I82101,I82109,I82126,I457103,I457118,I82143,I457100,I82169,I457097,I82186,I82194,I82211,I82043,I82242,I82259,I82055,I82299,I82064,I82321,I457112,I82338,I457115,I82364,I82381,I82067,I82403,I82052,I82434,I457109,I82451,I82468,I82485,I82061,I82516,I82049,I82058,I82046,I82602,I506729,I82628,I82636,I82653,I506747,I506741,I82670,I506720,I82696,I506738,I82713,I82721,I506723,I82738,I82570,I82769,I82786,I82582,I506735,I82826,I82591,I82848,I506744,I506732,I82865,I506726,I82891,I82908,I82594,I82930,I82579,I82961,I82978,I82995,I83012,I82588,I83043,I82576,I82585,I82573,I83129,I342628,I83155,I83163,I83180,I342640,I342625,I83197,I342619,I83223,I342634,I83240,I83248,I342622,I83265,I83097,I83296,I83313,I83109,I342631,I83353,I83118,I83375,I342637,I342643,I83392,I83418,I83435,I83121,I83457,I83106,I83488,I83505,I83522,I83539,I83115,I83570,I83103,I83112,I83100,I83659,I458157,I83685,I83693,I83719,I83727,I458154,I83744,I458166,I83761,I83636,I83792,I458160,I83630,I83823,I458172,I83840,I83857,I458163,I458151,I83874,I83891,I83908,I83645,I83642,I83648,I83967,I83984,I84001,I84027,I83627,I84058,I84066,I458169,I83651,I84097,I84114,I84131,I83633,I84162,I84179,I83624,I83639,I84254,I196428,I84280,I84288,I196425,I84314,I84322,I196422,I84339,I196434,I84356,I84231,I84387,I196443,I84225,I84418,I196440,I84435,I84452,I196419,I84469,I84486,I84503,I84240,I84237,I84243,I84562,I84579,I84596,I196431,I196446,I84622,I84222,I84653,I84661,I196437,I84246,I84692,I84709,I84726,I84228,I84757,I84774,I84219,I84234,I84849,I674020,I84875,I84883,I674017,I84909,I84917,I674035,I84934,I674029,I84951,I84982,I674023,I85013,I85030,I85047,I674026,I674032,I85064,I85081,I85098,I85157,I85174,I85191,I674038,I85217,I85248,I85256,I674041,I85287,I85304,I85321,I85352,I85369,I85444,I228080,I85470,I85478,I228074,I85504,I85512,I228071,I85529,I228062,I85546,I85421,I85577,I228065,I85415,I85608,I228068,I85625,I85642,I228056,I228083,I85659,I85676,I85693,I85430,I85427,I85433,I85752,I85769,I85786,I228059,I85812,I85412,I85843,I85851,I228077,I85436,I85882,I85899,I85916,I85418,I85947,I85964,I85409,I85424,I86039,I201171,I86065,I86073,I201168,I86099,I86107,I201165,I86124,I201177,I86141,I86016,I86172,I201186,I86010,I86203,I201183,I86220,I86237,I201162,I86254,I86271,I86288,I86025,I86022,I86028,I86347,I86364,I86381,I201174,I201189,I86407,I86007,I86438,I86446,I201180,I86031,I86477,I86494,I86511,I86013,I86542,I86559,I86004,I86019,I86634,I471859,I86660,I86668,I86694,I86702,I471856,I86719,I471868,I86736,I86611,I86767,I471862,I86605,I86798,I471874,I86815,I86832,I471865,I471853,I86849,I86866,I86883,I86620,I86617,I86623,I86942,I86959,I86976,I87002,I86602,I87033,I87041,I471871,I86626,I87072,I87089,I87106,I86608,I87137,I87154,I86599,I86614,I87229,I87255,I87263,I87289,I87297,I87314,I87331,I87206,I87362,I87200,I87393,I87410,I87427,I87444,I87461,I87478,I87215,I87212,I87218,I87537,I87554,I87571,I87597,I87197,I87628,I87636,I87221,I87667,I87684,I87701,I87203,I87732,I87749,I87194,I87209,I87824,I617920,I87850,I87858,I617917,I87884,I87892,I617926,I87909,I87926,I87801,I87957,I617929,I87795,I87988,I617923,I88005,I88022,I617938,I88039,I88056,I88073,I87810,I87807,I87813,I88132,I88149,I88166,I617941,I617935,I88192,I87792,I88223,I88231,I617932,I87816,I88262,I88279,I88296,I87798,I88327,I88344,I87789,I87804,I88416,I603467,I88442,I88459,I88408,I88481,I88507,I88515,I88532,I603470,I88549,I603482,I88566,I88583,I603488,I88600,I603479,I88617,I603485,I88634,I88384,I88665,I88682,I88699,I88716,I88396,I88390,I88761,I603476,I88405,I88399,I88806,I88823,I603473,I88840,I603491,I88857,I88883,I88891,I88393,I88387,I88945,I88953,I88402,I89011,I554255,I89037,I89054,I89003,I89076,I554264,I89102,I89110,I89127,I554258,I89144,I554252,I89161,I89178,I554267,I89195,I89212,I554261,I89229,I88979,I89260,I89277,I89294,I89311,I88991,I88985,I89356,I89000,I88994,I89401,I89418,I554273,I89435,I554270,I89452,I89478,I89486,I88988,I88982,I89540,I89548,I88997,I89606,I367485,I89632,I89649,I89598,I89671,I367482,I89697,I89705,I89722,I367488,I89739,I367473,I89756,I89773,I367476,I89790,I367497,I89807,I367494,I89824,I89574,I89855,I89872,I89889,I89906,I89586,I89580,I89951,I89595,I89589,I89996,I90013,I367479,I90030,I367491,I90047,I90073,I90081,I89583,I89577,I90135,I90143,I89592,I90201,I594797,I90227,I90244,I90266,I90292,I90300,I90317,I594800,I90334,I594812,I90351,I90368,I594818,I90385,I594809,I90402,I594815,I90419,I90450,I90467,I90484,I90501,I90546,I594806,I90591,I90608,I594803,I90625,I594821,I90642,I90668,I90676,I90730,I90738,I90796,I531929,I90822,I90839,I90788,I90861,I531938,I90887,I90895,I90912,I531926,I90929,I531917,I90946,I90963,I531923,I90980,I531941,I90997,I531914,I91014,I90764,I91045,I91062,I91079,I91096,I90776,I90770,I91141,I531920,I90785,I90779,I91186,I91203,I531932,I91220,I91237,I531935,I91263,I91271,I90773,I90767,I91325,I91333,I90782,I91391,I91417,I91434,I91383,I91456,I91482,I91490,I91507,I91524,I91541,I91558,I91575,I91592,I91609,I91359,I91640,I91657,I91674,I91691,I91371,I91365,I91736,I91380,I91374,I91781,I91798,I91815,I91832,I91858,I91866,I91368,I91362,I91920,I91928,I91377,I91986,I615605,I92012,I92029,I91978,I92051,I92077,I92085,I92102,I615608,I92119,I615620,I92136,I92153,I615626,I92170,I615617,I92187,I615623,I92204,I91954,I92235,I92252,I92269,I92286,I91966,I91960,I92331,I615614,I91975,I91969,I92376,I92393,I615611,I92410,I615629,I92427,I92453,I92461,I91963,I91957,I92515,I92523,I91972,I92581,I340322,I92607,I92624,I92573,I92646,I340313,I92672,I92680,I92697,I340331,I92714,I340328,I92731,I92748,I340307,I92765,I340310,I92782,I340319,I92799,I92549,I92830,I92847,I92864,I92881,I92561,I92555,I92926,I340325,I92570,I92564,I92971,I92988,I93005,I340316,I93022,I93048,I93056,I92558,I92552,I93110,I93118,I92567,I93176,I665928,I93202,I93219,I93168,I93241,I665940,I93267,I93275,I93292,I665934,I93309,I665946,I93326,I93343,I665931,I93360,I665943,I93377,I665925,I93394,I93144,I93425,I93442,I93459,I93476,I93156,I93150,I93521,I665937,I93165,I93159,I93566,I93583,I93600,I93617,I665949,I93643,I93651,I93153,I93147,I93705,I93713,I93162,I93771,I719224,I93797,I93814,I93836,I719215,I93862,I93870,I93887,I719209,I93904,I719203,I93921,I93938,I719230,I93955,I93972,I719227,I93989,I94020,I94037,I94054,I94071,I94116,I719212,I94161,I94178,I719218,I94195,I719221,I94212,I719206,I94238,I94246,I94300,I94308,I94366,I94392,I94409,I94431,I94457,I94465,I94482,I94499,I94516,I94533,I94550,I94567,I94584,I94615,I94632,I94649,I94666,I94711,I94756,I94773,I94790,I94807,I94833,I94841,I94895,I94903,I94961,I510611,I94987,I95004,I94953,I95026,I510620,I95052,I95060,I95077,I510608,I95094,I510599,I95111,I95128,I510605,I95145,I510623,I95162,I510596,I95179,I94929,I95210,I95227,I95244,I95261,I94941,I94935,I95306,I510602,I94950,I94944,I95351,I95368,I510614,I95385,I95402,I510617,I95428,I95436,I94938,I94932,I95490,I95498,I94947,I95556,I355347,I95582,I95599,I95548,I95621,I355344,I95647,I95655,I95672,I355350,I95689,I355335,I95706,I95723,I355338,I95740,I355359,I95757,I355356,I95774,I95524,I95805,I95822,I95839,I95856,I95536,I95530,I95901,I95545,I95539,I95946,I95963,I355341,I95980,I355353,I95997,I96023,I96031,I95533,I95527,I96085,I96093,I95542,I96151,I223823,I96177,I96194,I96143,I96216,I223838,I96242,I96250,I96267,I223835,I96284,I96301,I96318,I223832,I96335,I223847,I96352,I223844,I96369,I96119,I96400,I96417,I96434,I96451,I96131,I96125,I96496,I223841,I96140,I96134,I96541,I96558,I223829,I96575,I223850,I96592,I223826,I96618,I96626,I96128,I96122,I96680,I96688,I96137,I96746,I231344,I96772,I96789,I96738,I96811,I231332,I96837,I96845,I96862,I231341,I96879,I231338,I96896,I96913,I231329,I96930,I231335,I96947,I231320,I96964,I96714,I96995,I97012,I97029,I97046,I96726,I96720,I97091,I96735,I96729,I97136,I97153,I231326,I97170,I231323,I97187,I231347,I97213,I97221,I96723,I96717,I97275,I97283,I96732,I97341,I221188,I97367,I97384,I97333,I97406,I221203,I97432,I97440,I97457,I221200,I97474,I97491,I97508,I221197,I97525,I221212,I97542,I221209,I97559,I97309,I97590,I97607,I97624,I97641,I97321,I97315,I97686,I221206,I97330,I97324,I97731,I97748,I221194,I97765,I221215,I97782,I221191,I97808,I97816,I97318,I97312,I97870,I97878,I97327,I97936,I682112,I97962,I97979,I98001,I682124,I98027,I98035,I98052,I682118,I98069,I682130,I98086,I98103,I682115,I98120,I682127,I98137,I682109,I98154,I98185,I98202,I98219,I98236,I98281,I682121,I98326,I98343,I98360,I98377,I682133,I98403,I98411,I98465,I98473,I98531,I472913,I98557,I98574,I98523,I98596,I472907,I98622,I98630,I98647,I472925,I98664,I98681,I98698,I98715,I472919,I98732,I472910,I98749,I98499,I98780,I98797,I98814,I98831,I98511,I98505,I98876,I472922,I98520,I98514,I98921,I98938,I472928,I98955,I98972,I472916,I98998,I99006,I98508,I98502,I99060,I99068,I98517,I99126,I618495,I99152,I99169,I99118,I99191,I99217,I99225,I99242,I618498,I99259,I618510,I99276,I99293,I618516,I99310,I618507,I99327,I618513,I99344,I99094,I99375,I99392,I99409,I99426,I99106,I99100,I99471,I618504,I99115,I99109,I99516,I99533,I618501,I99550,I618519,I99567,I99593,I99601,I99103,I99097,I99655,I99663,I99112,I99721,I562670,I99747,I99764,I99713,I99786,I562679,I99812,I99820,I99837,I562673,I99854,I562667,I99871,I99888,I562682,I99905,I99922,I562676,I99939,I99689,I99970,I99987,I100004,I100021,I99701,I99695,I100066,I99710,I99704,I100111,I100128,I562688,I100145,I562685,I100162,I100188,I100196,I99698,I99692,I100250,I100258,I99707,I100316,I622541,I100342,I100359,I100308,I100381,I100407,I100415,I100432,I622544,I100449,I622556,I100466,I100483,I622562,I100500,I622553,I100517,I622559,I100534,I100284,I100565,I100582,I100599,I100616,I100296,I100290,I100661,I622550,I100305,I100299,I100706,I100723,I622547,I100740,I622565,I100757,I100783,I100791,I100293,I100287,I100845,I100853,I100302,I100911,I444455,I100937,I100954,I100903,I100976,I444449,I101002,I101010,I101027,I444467,I101044,I101061,I101078,I101095,I444461,I101112,I444452,I101129,I100879,I101160,I101177,I101194,I101211,I100891,I100885,I101256,I444464,I100900,I100894,I101301,I101318,I444470,I101335,I101352,I444458,I101378,I101386,I100888,I100882,I101440,I101448,I100897,I101506,I572255,I101532,I101549,I101498,I101571,I101597,I101605,I101622,I572258,I101639,I572270,I101656,I101673,I572276,I101690,I572267,I101707,I572273,I101724,I101474,I101755,I101772,I101789,I101806,I101486,I101480,I101851,I572264,I101495,I101489,I101896,I101913,I572261,I101930,I572279,I101947,I101973,I101981,I101483,I101477,I102035,I102043,I101492,I102101,I720414,I102127,I102144,I102093,I102166,I720405,I102192,I102200,I102217,I720399,I102234,I720393,I102251,I102268,I720420,I102285,I102302,I720417,I102319,I102069,I102350,I102367,I102384,I102401,I102081,I102075,I102446,I720402,I102090,I102084,I102491,I102508,I720408,I102525,I720411,I102542,I720396,I102568,I102576,I102078,I102072,I102630,I102638,I102087,I102696,I102722,I102739,I102761,I102787,I102795,I102812,I102829,I102846,I102863,I102880,I102897,I102914,I102945,I102962,I102979,I102996,I103041,I103086,I103103,I103120,I103137,I103163,I103171,I103225,I103233,I103291,I494461,I103317,I103334,I103283,I103356,I494470,I103382,I103390,I103407,I494458,I103424,I494449,I103441,I103458,I494455,I103475,I494473,I103492,I494446,I103509,I103259,I103540,I103557,I103574,I103591,I103271,I103265,I103636,I494452,I103280,I103274,I103681,I103698,I494464,I103715,I103732,I494467,I103758,I103766,I103268,I103262,I103820,I103828,I103277,I103886,I479603,I103912,I103929,I103878,I103951,I479612,I103977,I103985,I104002,I479600,I104019,I479591,I104036,I104053,I479597,I104070,I479615,I104087,I479588,I104104,I103854,I104135,I104152,I104169,I104186,I103866,I103860,I104231,I479594,I103875,I103869,I104276,I104293,I479606,I104310,I104327,I479609,I104353,I104361,I103863,I103857,I104415,I104423,I103872,I104481,I218553,I104507,I104524,I104473,I104546,I218568,I104572,I104580,I104597,I218565,I104614,I104631,I104648,I218562,I104665,I218577,I104682,I218574,I104699,I104449,I104730,I104747,I104764,I104781,I104461,I104455,I104826,I218571,I104470,I104464,I104871,I104888,I218559,I104905,I218580,I104922,I218556,I104948,I104956,I104458,I104452,I105010,I105018,I104467,I105076,I295065,I105102,I105119,I105141,I295059,I105167,I105175,I105192,I295074,I105209,I295071,I105226,I105243,I295062,I105260,I295053,I105277,I295056,I105294,I105325,I105342,I105359,I105376,I105421,I295077,I105466,I105483,I295068,I105500,I105517,I105543,I105551,I105605,I105613,I105671,I233520,I105697,I105714,I105663,I105736,I233508,I105762,I105770,I105787,I233517,I105804,I233514,I105821,I105838,I233505,I105855,I233511,I105872,I233496,I105889,I105639,I105920,I105937,I105954,I105971,I105651,I105645,I106016,I105660,I105654,I106061,I106078,I233502,I106095,I233499,I106112,I233523,I106138,I106146,I105648,I105642,I106200,I106208,I105657,I106266,I438658,I106292,I106309,I106258,I106331,I438652,I106357,I106365,I106382,I438670,I106399,I106416,I106433,I106450,I438664,I106467,I438655,I106484,I106234,I106515,I106532,I106549,I106566,I106246,I106240,I106611,I438667,I106255,I106249,I106656,I106673,I438673,I106690,I106707,I438661,I106733,I106741,I106243,I106237,I106795,I106803,I106252,I106861,I355925,I106887,I106904,I106853,I106926,I355922,I106952,I106960,I106977,I355928,I106994,I355913,I107011,I107028,I355916,I107045,I355937,I107062,I355934,I107079,I106829,I107110,I107127,I107144,I107161,I106841,I106835,I107206,I106850,I106844,I107251,I107268,I355919,I107285,I355931,I107302,I107328,I107336,I106838,I106832,I107390,I107398,I106847,I107456,I530637,I107482,I107499,I107448,I107521,I530646,I107547,I107555,I107572,I530634,I107589,I530625,I107606,I107623,I530631,I107640,I530649,I107657,I530622,I107674,I107424,I107705,I107722,I107739,I107756,I107436,I107430,I107801,I530628,I107445,I107439,I107846,I107863,I530640,I107880,I107897,I530643,I107923,I107931,I107433,I107427,I107985,I107993,I107442,I108051,I652887,I108077,I108094,I108043,I108116,I652872,I108142,I108150,I108167,I652890,I108184,I108201,I108218,I652893,I108235,I652884,I108252,I652881,I108269,I108019,I108300,I108317,I108334,I108351,I108031,I108025,I108396,I652878,I108040,I108034,I108441,I108458,I652869,I108475,I652875,I108492,I108518,I108526,I108028,I108022,I108580,I108588,I108037,I108646,I578613,I108672,I108689,I108711,I108737,I108745,I108762,I578616,I108779,I578628,I108796,I108813,I578634,I108830,I578625,I108847,I578631,I108864,I108895,I108912,I108929,I108946,I108991,I578622,I109036,I109053,I578619,I109070,I578637,I109087,I109113,I109121,I109175,I109183,I109241,I514487,I109267,I109284,I109233,I109306,I514496,I109332,I109340,I109357,I514484,I109374,I514475,I109391,I109408,I514481,I109425,I514499,I109442,I514472,I109459,I109209,I109490,I109507,I109524,I109541,I109221,I109215,I109586,I514478,I109230,I109224,I109631,I109648,I514490,I109665,I109682,I514493,I109708,I109716,I109218,I109212,I109770,I109778,I109227,I109836,I712084,I109862,I109879,I109828,I109901,I712075,I109927,I109935,I109952,I712069,I109969,I712063,I109986,I110003,I712090,I110020,I110037,I712087,I110054,I109804,I110085,I110102,I110119,I110136,I109816,I109810,I110181,I712072,I109825,I109819,I110226,I110243,I712078,I110260,I712081,I110277,I712066,I110303,I110311,I109813,I109807,I110365,I110373,I109822,I110431,I599421,I110457,I110474,I110423,I110496,I110522,I110530,I110547,I599424,I110564,I599436,I110581,I110598,I599442,I110615,I599433,I110632,I599439,I110649,I110399,I110680,I110697,I110714,I110731,I110411,I110405,I110776,I599430,I110420,I110414,I110821,I110838,I599427,I110855,I599445,I110872,I110898,I110906,I110408,I110402,I110960,I110968,I110417,I111026,I217499,I111052,I111069,I111018,I111091,I217514,I111117,I111125,I111142,I217511,I111159,I111176,I111193,I217508,I111210,I217523,I111227,I217520,I111244,I110994,I111275,I111292,I111309,I111326,I111006,I111000,I111371,I217517,I111015,I111009,I111416,I111433,I217505,I111450,I217526,I111467,I217502,I111493,I111501,I111003,I110997,I111555,I111563,I111012,I111621,I111647,I111664,I111686,I111712,I111720,I111737,I111754,I111771,I111788,I111805,I111822,I111839,I111870,I111887,I111904,I111921,I111966,I112011,I112028,I112045,I112062,I112088,I112096,I112150,I112158,I112216,I277040,I112242,I112259,I112281,I277028,I112307,I112315,I112332,I277037,I112349,I277034,I112366,I112383,I277025,I112400,I277031,I112417,I277016,I112434,I112465,I112482,I112499,I112516,I112561,I112606,I112623,I277022,I112640,I277019,I112657,I277043,I112683,I112691,I112745,I112753,I112811,I630633,I112837,I112854,I112876,I112902,I112910,I112927,I630636,I112944,I630648,I112961,I112978,I630654,I112995,I630645,I113012,I630651,I113029,I113060,I113077,I113094,I113111,I113156,I630642,I113201,I113218,I630639,I113235,I630657,I113252,I113278,I113286,I113340,I113348,I113406,I469751,I113432,I113449,I113398,I113471,I469745,I113497,I113505,I113522,I469763,I113539,I113556,I113573,I113590,I469757,I113607,I469748,I113624,I113374,I113655,I113672,I113689,I113706,I113386,I113380,I113751,I469760,I113395,I113389,I113796,I113813,I469766,I113830,I113847,I469754,I113873,I113881,I113383,I113377,I113935,I113943,I113392,I114001,I684992,I114027,I114044,I113993,I114066,I684965,I114092,I114100,I114117,I684989,I114134,I684986,I114151,I114168,I114185,I684983,I114202,I684971,I114219,I113969,I114250,I114267,I114284,I114301,I113981,I113975,I114346,I684977,I113990,I113984,I114391,I114408,I684980,I114425,I684968,I114442,I684974,I114468,I114476,I113978,I113972,I114530,I114538,I113987,I114596,I347255,I114622,I114639,I114588,I114661,I347252,I114687,I114695,I114712,I347258,I114729,I347243,I114746,I114763,I347246,I114780,I347267,I114797,I347264,I114814,I114564,I114845,I114862,I114879,I114896,I114576,I114570,I114941,I114585,I114579,I114986,I115003,I347249,I115020,I347261,I115037,I115063,I115071,I114573,I114567,I115125,I115133,I114582,I115191,I300420,I115217,I115234,I115183,I115256,I300414,I115282,I115290,I115307,I300429,I115324,I300426,I115341,I115358,I300417,I115375,I300408,I115392,I300411,I115409,I115159,I115440,I115457,I115474,I115491,I115171,I115165,I115536,I300432,I115180,I115174,I115581,I115598,I300423,I115615,I115632,I115658,I115666,I115168,I115162,I115720,I115728,I115177,I115786,I369219,I115812,I115829,I115778,I115851,I369216,I115877,I115885,I115902,I369222,I115919,I369207,I115936,I115953,I369210,I115970,I369231,I115987,I369228,I116004,I115754,I116035,I116052,I116069,I116086,I115766,I115760,I116131,I115775,I115769,I116176,I116193,I369213,I116210,I369225,I116227,I116253,I116261,I115763,I115757,I116315,I116323,I115772,I116381,I675754,I116407,I116424,I116373,I116446,I675766,I116472,I116480,I116497,I675760,I116514,I675772,I116531,I116548,I675757,I116565,I675769,I116582,I675751,I116599,I116349,I116630,I116647,I116664,I116681,I116361,I116355,I116726,I675763,I116370,I116364,I116771,I116788,I116805,I116822,I675775,I116848,I116856,I116358,I116352,I116910,I116918,I116367,I116976,I576879,I117002,I117019,I116968,I117041,I117067,I117075,I117092,I576882,I117109,I576894,I117126,I117143,I576900,I117160,I576891,I117177,I576897,I117194,I116944,I117225,I117242,I117259,I117276,I116956,I116950,I117321,I576888,I116965,I116959,I117366,I117383,I576885,I117400,I576903,I117417,I117443,I117451,I116953,I116947,I117505,I117513,I116962,I117571,I353613,I117597,I117614,I117563,I117636,I353610,I117662,I117670,I117687,I353616,I117704,I353601,I117721,I117738,I353604,I117755,I353625,I117772,I353622,I117789,I117539,I117820,I117837,I117854,I117871,I117551,I117545,I117916,I117560,I117554,I117961,I117978,I353607,I117995,I353619,I118012,I118038,I118046,I117548,I117542,I118100,I118108,I117557,I118166,I118192,I118209,I118158,I118231,I118257,I118265,I118282,I118299,I118316,I118333,I118350,I118367,I118384,I118134,I118415,I118432,I118449,I118466,I118146,I118140,I118511,I118155,I118149,I118556,I118573,I118590,I118607,I118633,I118641,I118143,I118137,I118695,I118703,I118152,I118761,I548645,I118787,I118804,I118753,I118826,I548654,I118852,I118860,I118877,I548648,I118894,I548642,I118911,I118928,I548657,I118945,I118962,I548651,I118979,I118729,I119010,I119027,I119044,I119061,I118741,I118735,I119106,I118750,I118744,I119151,I119168,I548663,I119185,I548660,I119202,I119228,I119236,I118738,I118732,I119290,I119298,I118747,I119356,I119382,I119399,I119348,I119421,I119447,I119455,I119472,I119489,I119506,I119523,I119540,I119557,I119574,I119324,I119605,I119622,I119639,I119656,I119336,I119330,I119701,I119345,I119339,I119746,I119763,I119780,I119797,I119823,I119831,I119333,I119327,I119885,I119893,I119342,I119951,I252016,I119977,I119994,I119943,I120016,I252004,I120042,I120050,I120067,I252013,I120084,I252010,I120101,I120118,I252001,I120135,I252007,I120152,I251992,I120169,I119919,I120200,I120217,I120234,I120251,I119931,I119925,I120296,I119940,I119934,I120341,I120358,I251998,I120375,I251995,I120392,I252019,I120418,I120426,I119928,I119922,I120480,I120488,I119937,I120546,I638147,I120572,I120589,I120538,I120611,I120637,I120645,I120662,I638150,I120679,I638162,I120696,I120713,I638168,I120730,I638159,I120747,I638165,I120764,I120514,I120795,I120812,I120829,I120846,I120526,I120520,I120891,I638156,I120535,I120529,I120936,I120953,I638153,I120970,I638171,I120987,I121013,I121021,I120523,I120517,I121075,I121083,I120532,I121141,I595375,I121167,I121184,I121133,I121206,I121232,I121240,I121257,I595378,I121274,I595390,I121291,I121308,I595396,I121325,I595387,I121342,I595393,I121359,I121109,I121390,I121407,I121424,I121441,I121121,I121115,I121486,I595384,I121130,I121124,I121531,I121548,I595381,I121565,I595399,I121582,I121608,I121616,I121118,I121112,I121670,I121678,I121127,I121736,I631789,I121762,I121779,I121728,I121801,I121827,I121835,I121852,I631792,I121869,I631804,I121886,I121903,I631810,I121920,I631801,I121937,I631807,I121954,I121704,I121985,I122002,I122019,I122036,I121716,I121710,I122081,I631798,I121725,I121719,I122126,I122143,I631795,I122160,I631813,I122177,I122203,I122211,I121713,I121707,I122265,I122273,I121722,I122331,I476602,I122357,I122374,I122323,I122396,I476596,I122422,I122430,I122447,I476614,I122464,I122481,I122498,I122515,I476608,I122532,I476599,I122549,I122299,I122580,I122597,I122614,I122631,I122311,I122305,I122676,I476611,I122320,I122314,I122721,I122738,I476617,I122755,I122772,I476605,I122798,I122806,I122308,I122302,I122860,I122868,I122317,I122926,I634101,I122952,I122969,I122918,I122991,I123017,I123025,I123042,I634104,I123059,I634116,I123076,I123093,I634122,I123110,I634113,I123127,I634119,I123144,I122894,I123175,I123192,I123209,I123226,I122906,I122900,I123271,I634110,I122915,I122909,I123316,I123333,I634107,I123350,I634125,I123367,I123393,I123401,I122903,I122897,I123455,I123463,I122912,I123521,I440766,I123547,I123564,I123586,I440760,I123612,I123620,I123637,I440778,I123654,I123671,I123688,I123705,I440772,I123722,I440763,I123739,I123770,I123787,I123804,I123821,I123866,I440775,I123911,I123928,I440781,I123945,I123962,I440769,I123988,I123996,I124050,I124058,I124116,I620807,I124142,I124159,I124108,I124181,I124207,I124215,I124232,I620810,I124249,I620822,I124266,I124283,I620828,I124300,I620819,I124317,I620825,I124334,I124084,I124365,I124382,I124399,I124416,I124096,I124090,I124461,I620816,I124105,I124099,I124506,I124523,I620813,I124540,I620831,I124557,I124583,I124591,I124093,I124087,I124645,I124653,I124102,I124711,I124737,I124754,I124776,I124802,I124810,I124827,I124844,I124861,I124878,I124895,I124912,I124929,I124960,I124977,I124994,I125011,I125056,I125101,I125118,I125135,I125152,I125178,I125186,I125240,I125248,I125306,I515779,I125332,I125349,I125298,I125371,I515788,I125397,I125405,I125422,I515776,I125439,I515767,I125456,I125473,I515773,I125490,I515791,I125507,I515764,I125524,I125274,I125555,I125572,I125589,I125606,I125286,I125280,I125651,I515770,I125295,I125289,I125696,I125713,I515782,I125730,I125747,I515785,I125773,I125781,I125283,I125277,I125835,I125843,I125292,I125901,I125927,I125944,I125966,I125992,I126000,I126017,I126034,I126051,I126068,I126085,I126102,I126119,I126150,I126167,I126184,I126201,I126246,I126291,I126308,I126325,I126342,I126368,I126376,I126430,I126438,I126496,I595953,I126522,I126539,I126488,I126561,I126587,I126595,I126612,I595956,I126629,I595968,I126646,I126663,I595974,I126680,I595965,I126697,I595971,I126714,I126464,I126745,I126762,I126779,I126796,I126476,I126470,I126841,I595962,I126485,I126479,I126886,I126903,I595959,I126920,I595977,I126937,I126963,I126971,I126473,I126467,I127025,I127033,I126482,I127091,I127117,I127134,I127083,I127156,I127182,I127190,I127207,I127224,I127241,I127258,I127275,I127292,I127309,I127059,I127340,I127357,I127374,I127391,I127071,I127065,I127436,I127080,I127074,I127481,I127498,I127515,I127532,I127558,I127566,I127068,I127062,I127620,I127628,I127077,I127686,I593641,I127712,I127729,I127751,I127777,I127785,I127802,I593644,I127819,I593656,I127836,I127853,I593662,I127870,I593653,I127887,I593659,I127904,I127935,I127952,I127969,I127986,I128031,I593650,I128076,I128093,I593647,I128110,I593665,I128127,I128153,I128161,I128215,I128223,I128281,I597109,I128307,I128324,I128273,I128346,I128372,I128380,I128397,I597112,I128414,I597124,I128431,I128448,I597130,I128465,I597121,I128482,I597127,I128499,I128249,I128530,I128547,I128564,I128581,I128261,I128255,I128626,I597118,I128270,I128264,I128671,I128688,I597115,I128705,I597133,I128722,I128748,I128756,I128258,I128252,I128810,I128818,I128267,I128876,I305642,I128902,I128919,I128868,I128941,I305633,I128967,I128975,I128992,I305651,I129009,I305648,I129026,I129043,I305627,I129060,I305630,I129077,I305639,I129094,I128844,I129125,I129142,I129159,I129176,I128856,I128850,I129221,I305645,I128865,I128859,I129266,I129283,I129300,I305636,I129317,I129343,I129351,I128853,I128847,I129405,I129413,I128862,I129471,I411413,I129497,I129514,I129463,I129536,I411410,I129562,I129570,I129587,I411416,I129604,I411401,I129621,I129638,I411404,I129655,I411425,I129672,I411422,I129689,I129439,I129720,I129737,I129754,I129771,I129451,I129445,I129816,I129460,I129454,I129861,I129878,I411407,I129895,I411419,I129912,I129938,I129946,I129448,I129442,I130000,I130008,I129457,I130066,I130092,I130109,I130058,I130131,I130157,I130165,I130182,I130199,I130216,I130233,I130250,I130267,I130284,I130034,I130315,I130332,I130349,I130366,I130046,I130040,I130411,I130055,I130049,I130456,I130473,I130490,I130507,I130533,I130541,I130043,I130037,I130595,I130603,I130052,I130661,I309110,I130687,I130704,I130653,I130726,I309101,I130752,I130760,I130777,I309119,I130794,I309116,I130811,I130828,I309095,I130845,I309098,I130862,I309107,I130879,I130629,I130910,I130927,I130944,I130961,I130641,I130635,I131006,I309113,I130650,I130644,I131051,I131068,I131085,I309104,I131102,I131128,I131136,I130638,I130632,I131190,I131198,I130647,I131256,I468697,I131282,I131299,I131248,I131321,I468691,I131347,I131355,I131372,I468709,I131389,I131406,I131423,I131440,I468703,I131457,I468694,I131474,I131224,I131505,I131522,I131539,I131556,I131236,I131230,I131601,I468706,I131245,I131239,I131646,I131663,I468712,I131680,I131697,I468700,I131723,I131731,I131233,I131227,I131785,I131793,I131242,I131851,I524823,I131877,I131894,I131843,I131916,I524832,I131942,I131950,I131967,I524820,I131984,I524811,I132001,I132018,I524817,I132035,I524835,I132052,I524808,I132069,I131819,I132100,I132117,I132134,I132151,I131831,I131825,I132196,I524814,I131840,I131834,I132241,I132258,I524826,I132275,I132292,I524829,I132318,I132326,I131828,I131822,I132380,I132388,I131837,I132446,I418927,I132472,I132489,I132438,I132511,I418924,I132537,I132545,I132562,I418930,I132579,I418915,I132596,I132613,I418918,I132630,I418939,I132647,I418936,I132664,I132414,I132695,I132712,I132729,I132746,I132426,I132420,I132791,I132435,I132429,I132836,I132853,I418921,I132870,I418933,I132887,I132913,I132921,I132423,I132417,I132975,I132983,I132432,I133041,I504797,I133067,I133084,I133033,I133106,I504806,I133132,I133140,I133157,I504794,I133174,I504785,I133191,I133208,I504791,I133225,I504809,I133242,I504782,I133259,I133009,I133290,I133307,I133324,I133341,I133021,I133015,I133386,I504788,I133030,I133024,I133431,I133448,I504800,I133465,I133482,I504803,I133508,I133516,I133018,I133012,I133570,I133578,I133027,I133636,I451306,I133662,I133679,I133628,I133701,I451300,I133727,I133735,I133752,I451318,I133769,I133786,I133803,I133820,I451312,I133837,I451303,I133854,I133604,I133885,I133902,I133919,I133936,I133616,I133610,I133981,I451315,I133625,I133619,I134026,I134043,I451321,I134060,I134077,I451309,I134103,I134111,I133613,I133607,I134165,I134173,I133622,I134231,I673442,I134257,I134274,I134223,I134296,I673454,I134322,I134330,I134347,I673448,I134364,I673460,I134381,I134398,I673445,I134415,I673457,I134432,I673439,I134449,I134199,I134480,I134497,I134514,I134531,I134211,I134205,I134576,I673451,I134220,I134214,I134621,I134638,I134655,I134672,I673463,I134698,I134706,I134208,I134202,I134760,I134768,I134217,I134826,I643095,I134852,I134869,I134818,I134891,I643080,I134917,I134925,I134942,I643098,I134959,I134976,I134993,I643101,I135010,I643092,I135027,I643089,I135044,I134794,I135075,I135092,I135109,I135126,I134806,I134800,I135171,I643086,I134815,I134809,I135216,I135233,I643077,I135250,I643083,I135267,I135293,I135301,I134803,I134797,I135355,I135363,I134812,I135421,I293875,I135447,I135464,I135413,I135486,I293869,I135512,I135520,I135537,I293884,I135554,I293881,I135571,I135588,I293872,I135605,I293863,I135622,I293866,I135639,I135389,I135670,I135687,I135704,I135721,I135401,I135395,I135766,I293887,I135410,I135404,I135811,I135828,I293878,I135845,I135862,I135888,I135896,I135398,I135392,I135950,I135958,I135407,I136016,I166380,I136042,I136059,I136008,I136081,I166395,I136107,I136115,I136132,I166392,I136149,I136166,I136183,I166389,I136200,I166404,I136217,I166401,I136234,I135984,I136265,I136282,I136299,I136316,I135996,I135990,I136361,I166398,I136005,I135999,I136406,I136423,I166386,I136440,I166407,I136457,I166383,I136483,I136491,I135993,I135987,I136545,I136553,I136002,I136611,I626009,I136637,I136654,I136603,I136676,I136702,I136710,I136727,I626012,I136744,I626024,I136761,I136778,I626030,I136795,I626021,I136812,I626027,I136829,I136579,I136860,I136877,I136894,I136911,I136591,I136585,I136956,I626018,I136600,I136594,I137001,I137018,I626015,I137035,I626033,I137052,I137078,I137086,I136588,I136582,I137140,I137148,I136597,I137206,I486709,I137232,I137249,I137198,I137271,I486718,I137297,I137305,I137322,I486706,I137339,I486697,I137356,I137373,I486703,I137390,I486721,I137407,I486694,I137424,I137174,I137455,I137472,I137489,I137506,I137186,I137180,I137551,I486700,I137195,I137189,I137596,I137613,I486712,I137630,I137647,I486715,I137673,I137681,I137183,I137177,I137735,I137743,I137192,I137801,I370375,I137827,I137844,I137793,I137866,I370372,I137892,I137900,I137917,I370378,I137934,I370363,I137951,I137968,I370366,I137985,I370387,I138002,I370384,I138019,I137769,I138050,I138067,I138084,I138101,I137781,I137775,I138146,I137790,I137784,I138191,I138208,I370369,I138225,I370381,I138242,I138268,I138276,I137778,I137772,I138330,I138338,I137787,I138396,I527407,I138422,I138439,I138388,I138461,I527416,I138487,I138495,I138512,I527404,I138529,I527395,I138546,I138563,I527401,I138580,I527419,I138597,I527392,I138614,I138364,I138645,I138662,I138679,I138696,I138376,I138370,I138741,I527398,I138385,I138379,I138786,I138803,I527410,I138820,I138837,I527413,I138863,I138871,I138373,I138367,I138925,I138933,I138382,I138991,I139017,I139034,I138983,I139056,I139082,I139090,I139107,I139124,I139141,I139158,I139175,I139192,I139209,I138959,I139240,I139257,I139274,I139291,I138971,I138965,I139336,I138980,I138974,I139381,I139398,I139415,I139432,I139458,I139466,I138968,I138962,I139520,I139528,I138977,I139586,I321826,I139612,I139629,I139651,I321817,I139677,I139685,I139702,I321835,I139719,I321832,I139736,I139753,I321811,I139770,I321814,I139787,I321823,I139804,I139835,I139852,I139869,I139886,I139931,I321829,I139976,I139993,I140010,I321820,I140027,I140053,I140061,I140115,I140123,I140181,I680378,I140207,I140224,I140246,I680390,I140272,I140280,I140297,I680384,I140314,I680396,I140331,I140348,I680381,I140365,I680393,I140382,I680375,I140399,I140430,I140447,I140464,I140481,I140526,I680387,I140571,I140588,I140605,I140622,I680399,I140648,I140656,I140710,I140718,I140776,I227536,I140802,I140819,I140768,I140841,I227524,I140867,I140875,I140892,I227533,I140909,I227530,I140926,I140943,I227521,I140960,I227527,I140977,I227512,I140994,I140744,I141025,I141042,I141059,I141076,I140756,I140750,I141121,I140765,I140759,I141166,I141183,I227518,I141200,I227515,I141217,I227539,I141243,I141251,I140753,I140747,I141305,I141313,I140762,I141371,I685553,I141397,I141414,I141363,I141436,I685526,I141462,I141470,I141487,I685550,I141504,I685547,I141521,I141538,I141555,I685544,I141572,I685532,I141589,I141339,I141620,I141637,I141654,I141671,I141351,I141345,I141716,I685538,I141360,I141354,I141761,I141778,I685541,I141795,I685529,I141812,I685535,I141838,I141846,I141348,I141342,I141900,I141908,I141357,I141966,I631211,I141992,I142009,I142031,I142057,I142065,I142082,I631214,I142099,I631226,I142116,I142133,I631232,I142150,I631223,I142167,I631229,I142184,I142215,I142232,I142249,I142266,I142311,I631220,I142356,I142373,I631217,I142390,I631235,I142407,I142433,I142441,I142495,I142503,I142561,I516425,I142587,I142604,I142553,I142626,I516434,I142652,I142660,I142677,I516422,I142694,I516413,I142711,I142728,I516419,I142745,I516437,I142762,I516410,I142779,I142529,I142810,I142827,I142844,I142861,I142541,I142535,I142906,I516416,I142550,I142544,I142951,I142968,I516428,I142985,I143002,I516431,I143028,I143036,I142538,I142532,I143090,I143098,I142547,I143156,I279760,I143182,I143199,I143148,I143221,I279748,I143247,I143255,I143272,I279757,I143289,I279754,I143306,I143323,I279745,I143340,I279751,I143357,I279736,I143374,I143124,I143405,I143422,I143439,I143456,I143136,I143130,I143501,I143145,I143139,I143546,I143563,I279742,I143580,I279739,I143597,I279763,I143623,I143631,I143133,I143127,I143685,I143693,I143142,I143751,I482833,I143777,I143794,I143743,I143816,I482842,I143842,I143850,I143867,I482830,I143884,I482821,I143901,I143918,I482827,I143935,I482845,I143952,I482818,I143969,I143719,I144000,I144017,I144034,I144051,I143731,I143725,I144096,I482824,I143740,I143734,I144141,I144158,I482836,I144175,I144192,I482839,I144218,I144226,I143728,I143722,I144280,I144288,I143737,I144346,I365751,I144372,I144389,I144338,I144411,I365748,I144437,I144445,I144462,I365754,I144479,I365739,I144496,I144513,I365742,I144530,I365763,I144547,I365760,I144564,I144314,I144595,I144612,I144629,I144646,I144326,I144320,I144691,I144335,I144329,I144736,I144753,I365745,I144770,I365757,I144787,I144813,I144821,I144323,I144317,I144875,I144883,I144332,I144941,I169015,I144967,I144984,I144933,I145006,I169030,I145032,I145040,I145057,I169027,I145074,I145091,I145108,I169024,I145125,I169039,I145142,I169036,I145159,I144909,I145190,I145207,I145224,I145241,I144921,I144915,I145286,I169033,I144930,I144924,I145331,I145348,I169021,I145365,I169042,I145382,I169018,I145408,I145416,I144918,I144912,I145470,I145478,I144927,I145536,I581503,I145562,I145579,I145528,I145601,I145627,I145635,I145652,I581506,I145669,I581518,I145686,I145703,I581524,I145720,I581515,I145737,I581521,I145754,I145504,I145785,I145802,I145819,I145836,I145516,I145510,I145881,I581512,I145525,I145519,I145926,I145943,I581509,I145960,I581527,I145977,I146003,I146011,I145513,I145507,I146065,I146073,I145522,I146131,I348411,I146157,I146174,I146123,I146196,I348408,I146222,I146230,I146247,I348414,I146264,I348399,I146281,I146298,I348402,I146315,I348423,I146332,I348420,I146349,I146099,I146380,I146397,I146414,I146431,I146111,I146105,I146476,I146120,I146114,I146521,I146538,I348405,I146555,I348417,I146572,I146598,I146606,I146108,I146102,I146660,I146668,I146117,I146726,I259088,I146752,I146769,I146718,I146791,I259076,I146817,I146825,I146842,I259085,I146859,I259082,I146876,I146893,I259073,I146910,I259079,I146927,I259064,I146944,I146694,I146975,I146992,I147009,I147026,I146706,I146700,I147071,I146715,I146709,I147116,I147133,I259070,I147150,I259067,I147167,I259091,I147193,I147201,I146703,I146697,I147255,I147263,I146712,I147321,I260720,I147347,I147364,I147313,I147386,I260708,I147412,I147420,I147437,I260717,I147454,I260714,I147471,I147488,I260705,I147505,I260711,I147522,I260696,I147539,I147289,I147570,I147587,I147604,I147621,I147301,I147295,I147666,I147310,I147304,I147711,I147728,I260702,I147745,I260699,I147762,I260723,I147788,I147796,I147298,I147292,I147850,I147858,I147307,I147916,I352457,I147942,I147959,I147908,I147981,I352454,I148007,I148015,I148032,I352460,I148049,I352445,I148066,I148083,I352448,I148100,I352469,I148117,I352466,I148134,I147884,I148165,I148182,I148199,I148216,I147896,I147890,I148261,I147905,I147899,I148306,I148323,I352451,I148340,I352463,I148357,I148383,I148391,I147893,I147887,I148445,I148453,I147902,I148511,I198527,I148537,I148554,I148503,I148576,I198542,I148602,I148610,I148627,I198539,I148644,I148661,I148678,I198536,I148695,I198551,I148712,I198548,I148729,I148479,I148760,I148777,I148794,I148811,I148491,I148485,I148856,I198545,I148500,I148494,I148901,I148918,I198533,I148935,I198554,I148952,I198530,I148978,I148986,I148488,I148482,I149040,I149048,I148497,I149106,I149132,I149149,I149098,I149171,I149197,I149205,I149222,I149239,I149256,I149273,I149290,I149307,I149324,I149074,I149355,I149372,I149389,I149406,I149086,I149080,I149451,I149095,I149089,I149496,I149513,I149530,I149547,I149573,I149581,I149083,I149077,I149635,I149643,I149092,I149701,I713869,I149727,I149744,I149693,I149766,I713860,I149792,I149800,I149817,I713854,I149834,I713848,I149851,I149868,I713875,I149885,I149902,I713872,I149919,I149669,I149950,I149967,I149984,I150001,I149681,I149675,I150046,I713857,I149690,I149684,I150091,I150108,I713863,I150125,I713866,I150142,I713851,I150168,I150176,I149678,I149672,I150230,I150238,I149687,I150296,I590751,I150322,I150339,I150288,I150361,I150387,I150395,I150412,I590754,I150429,I590766,I150446,I150463,I590772,I150480,I590763,I150497,I590769,I150514,I150264,I150545,I150562,I150579,I150596,I150276,I150270,I150641,I590760,I150285,I150279,I150686,I150703,I590757,I150720,I590775,I150737,I150763,I150771,I150273,I150267,I150825,I150833,I150282,I150891,I540791,I150917,I150934,I150883,I150956,I540800,I150982,I150990,I151007,I540794,I151024,I540788,I151041,I151058,I540803,I151075,I151092,I540797,I151109,I150859,I151140,I151157,I151174,I151191,I150871,I150865,I151236,I150880,I150874,I151281,I151298,I540809,I151315,I540806,I151332,I151358,I151366,I150868,I150862,I151420,I151428,I150877,I151486,I151512,I151529,I151478,I151551,I151577,I151585,I151602,I151619,I151636,I151653,I151670,I151687,I151704,I151454,I151735,I151752,I151769,I151786,I151466,I151460,I151831,I151475,I151469,I151876,I151893,I151910,I151927,I151953,I151961,I151463,I151457,I152015,I152023,I151472,I152081,I327606,I152107,I152124,I152073,I152146,I327597,I152172,I152180,I152197,I327615,I152214,I327612,I152231,I152248,I327591,I152265,I327594,I152282,I327603,I152299,I152049,I152330,I152347,I152364,I152381,I152061,I152055,I152426,I327609,I152070,I152064,I152471,I152488,I152505,I327600,I152522,I152548,I152556,I152058,I152052,I152610,I152618,I152067,I152676,I283760,I152702,I152719,I152741,I283754,I152767,I152775,I152792,I283769,I152809,I283766,I152826,I152843,I283757,I152860,I283748,I152877,I283751,I152894,I152925,I152942,I152959,I152976,I153021,I283772,I153066,I153083,I283763,I153100,I153117,I153143,I153151,I153205,I153213,I153271,I398697,I153297,I153314,I153263,I153336,I398694,I153362,I153370,I153387,I398700,I153404,I398685,I153421,I153438,I398688,I153455,I398709,I153472,I398706,I153489,I153239,I153520,I153537,I153554,I153571,I153251,I153245,I153616,I153260,I153254,I153661,I153678,I398691,I153695,I398703,I153712,I153738,I153746,I153248,I153242,I153800,I153808,I153257,I153866,I636413,I153892,I153909,I153858,I153931,I153957,I153965,I153982,I636416,I153999,I636428,I154016,I154033,I636434,I154050,I636425,I154067,I636431,I154084,I153834,I154115,I154132,I154149,I154166,I153846,I153840,I154211,I636422,I153855,I153849,I154256,I154273,I636419,I154290,I636437,I154307,I154333,I154341,I153843,I153837,I154395,I154403,I153852,I154461,I350145,I154487,I154504,I154526,I350142,I154552,I154560,I154577,I350148,I154594,I350133,I154611,I154628,I350136,I154645,I350157,I154662,I350154,I154679,I154710,I154727,I154744,I154761,I154806,I154851,I154868,I350139,I154885,I350151,I154902,I154928,I154936,I154990,I154998,I155056,I269968,I155082,I155099,I155121,I269956,I155147,I155155,I155172,I269965,I155189,I269962,I155206,I155223,I269953,I155240,I269959,I155257,I269944,I155274,I155305,I155322,I155339,I155356,I155401,I155446,I155463,I269950,I155480,I269947,I155497,I269971,I155523,I155531,I155585,I155593,I155651,I587283,I155677,I155694,I155643,I155716,I155742,I155750,I155767,I587286,I155784,I587298,I155801,I155818,I587304,I155835,I587295,I155852,I587301,I155869,I155619,I155900,I155917,I155934,I155951,I155631,I155625,I155996,I587292,I155640,I155634,I156041,I156058,I587289,I156075,I587307,I156092,I156118,I156126,I155628,I155622,I156180,I156188,I155637,I156246,I156272,I156289,I156238,I156311,I156337,I156345,I156362,I156379,I156396,I156413,I156430,I156447,I156464,I156214,I156495,I156512,I156529,I156546,I156226,I156220,I156591,I156235,I156229,I156636,I156653,I156670,I156687,I156713,I156721,I156223,I156217,I156775,I156783,I156232,I156841,I235152,I156867,I156884,I156833,I156906,I235140,I156932,I156940,I156957,I235149,I156974,I235146,I156991,I157008,I235137,I157025,I235143,I157042,I235128,I157059,I156809,I157090,I157107,I157124,I157141,I156821,I156815,I157186,I156830,I156824,I157231,I157248,I235134,I157265,I235131,I157282,I235155,I157308,I157316,I156818,I156812,I157370,I157378,I156827,I157436,I201689,I157462,I157479,I157428,I157501,I201704,I157527,I157535,I157552,I201701,I157569,I157586,I157603,I201698,I157620,I201713,I157637,I201710,I157654,I157404,I157685,I157702,I157719,I157736,I157416,I157410,I157781,I201707,I157425,I157419,I157826,I157843,I201695,I157860,I201716,I157877,I201692,I157903,I157911,I157413,I157407,I157965,I157973,I157422,I158031,I169542,I158057,I158074,I158023,I158096,I169557,I158122,I158130,I158147,I169554,I158164,I158181,I158198,I169551,I158215,I169566,I158232,I169563,I158249,I157999,I158280,I158297,I158314,I158331,I158011,I158005,I158376,I169560,I158020,I158014,I158421,I158438,I169548,I158455,I169569,I158472,I169545,I158498,I158506,I158008,I158002,I158560,I158568,I158017,I158626,I158652,I158669,I158691,I158717,I158725,I158742,I158759,I158776,I158793,I158810,I158827,I158844,I158875,I158892,I158909,I158926,I158971,I159016,I159033,I159050,I159067,I159093,I159101,I159155,I159163,I159221,I447090,I159247,I159264,I159213,I159286,I447084,I159312,I159320,I159337,I447102,I159354,I159371,I159388,I159405,I447096,I159422,I447087,I159439,I159189,I159470,I159487,I159504,I159521,I159201,I159195,I159566,I447099,I159210,I159204,I159611,I159628,I447105,I159645,I159662,I447093,I159688,I159696,I159198,I159192,I159750,I159758,I159207,I159816,I159842,I159859,I159808,I159881,I159907,I159915,I159932,I159949,I159966,I159983,I160000,I160017,I160034,I159784,I160065,I160082,I160099,I160116,I159796,I159790,I160161,I159805,I159799,I160206,I160223,I160240,I160257,I160283,I160291,I159793,I159787,I160345,I160353,I159802,I160411,I351879,I160437,I160454,I160403,I160476,I351876,I160502,I160510,I160527,I351882,I160544,I351867,I160561,I160578,I351870,I160595,I351891,I160612,I351888,I160629,I160379,I160660,I160677,I160694,I160711,I160391,I160385,I160756,I160400,I160394,I160801,I160818,I351873,I160835,I351885,I160852,I160878,I160886,I160388,I160382,I160940,I160948,I160397,I161006,I161032,I161049,I160998,I161071,I161097,I161105,I161122,I161139,I161156,I161173,I161190,I161207,I161224,I160974,I161255,I161272,I161289,I161306,I160986,I160980,I161351,I160995,I160989,I161396,I161413,I161430,I161447,I161473,I161481,I160983,I160977,I161535,I161543,I160992,I161601,I706729,I161627,I161644,I161593,I161666,I706720,I161692,I161700,I161717,I706714,I161734,I706708,I161751,I161768,I706735,I161785,I161802,I706732,I161819,I161569,I161850,I161867,I161884,I161901,I161581,I161575,I161946,I706717,I161590,I161584,I161991,I162008,I706723,I162025,I706726,I162042,I706711,I162068,I162076,I161578,I161572,I162130,I162138,I161587,I162199,I263428,I162225,I162233,I263440,I263419,I162250,I263443,I162276,I162167,I162298,I263434,I162324,I162332,I263416,I162349,I162375,I162191,I162397,I162173,I263431,I162437,I162454,I162462,I162479,I162176,I162510,I263422,I162527,I263425,I162553,I162561,I162164,I162182,I162606,I263437,I162623,I162185,I162170,I162179,I162188,I162726,I393495,I162752,I162760,I393486,I393501,I162777,I393507,I162803,I162694,I162825,I393492,I162851,I162859,I162876,I162902,I162718,I162924,I162700,I393489,I162964,I162981,I162989,I163006,I162703,I163037,I393483,I393498,I163054,I163080,I163088,I162691,I162709,I163133,I393504,I163150,I162712,I162697,I162706,I162715,I163253,I401587,I163279,I163287,I401578,I401593,I163304,I401599,I163330,I163221,I163352,I401584,I163378,I163386,I163403,I163429,I163245,I163451,I163227,I401581,I163491,I163508,I163516,I163533,I163230,I163564,I401575,I401590,I163581,I163607,I163615,I163218,I163236,I163660,I401596,I163677,I163239,I163224,I163233,I163242,I163780,I409101,I163806,I163814,I409092,I409107,I163831,I409113,I163857,I163748,I163879,I409098,I163905,I163913,I163930,I163956,I163772,I163978,I163754,I409095,I164018,I164035,I164043,I164060,I163757,I164091,I409089,I409104,I164108,I164134,I164142,I163745,I163763,I164187,I409110,I164204,I163766,I163751,I163760,I163769,I164307,I240036,I164333,I164341,I240048,I240027,I164358,I240051,I164384,I164275,I164406,I240042,I164432,I164440,I240024,I164457,I164483,I164299,I164505,I164281,I240039,I164545,I164562,I164570,I164587,I164284,I164618,I240030,I164635,I240033,I164661,I164669,I164272,I164290,I164714,I240045,I164731,I164293,I164278,I164287,I164296,I164834,I234052,I164860,I164868,I234064,I234043,I164885,I234067,I164911,I164802,I164933,I234058,I164959,I164967,I234040,I164984,I165010,I164826,I165032,I164808,I234055,I165072,I165089,I165097,I165114,I164811,I165145,I234046,I165162,I234049,I165188,I165196,I164799,I164817,I165241,I234061,I165258,I164820,I164805,I164814,I164823,I165361,I165387,I165395,I165412,I165438,I165329,I165460,I165486,I165494,I165511,I165537,I165353,I165559,I165335,I165599,I165616,I165624,I165641,I165338,I165672,I165689,I165715,I165723,I165326,I165344,I165768,I165785,I165347,I165332,I165341,I165350,I165888,I286131,I165914,I165922,I286143,I165939,I286128,I165965,I165856,I165987,I286152,I166013,I166021,I286149,I166038,I166064,I165880,I166086,I165862,I286140,I166126,I166143,I166151,I166168,I165865,I166199,I286137,I166216,I286146,I166242,I166250,I165853,I165871,I166295,I286134,I166312,I165874,I165859,I165868,I165877,I166415,I247108,I166441,I166449,I247120,I247099,I166466,I247123,I166492,I166514,I247114,I166540,I166548,I247096,I166565,I166591,I166613,I247111,I166653,I166670,I166678,I166695,I166726,I247102,I166743,I247105,I166769,I166777,I166822,I247117,I166839,I166942,I166968,I166976,I166993,I167019,I166910,I167041,I167067,I167075,I167092,I167118,I166934,I167140,I166916,I167180,I167197,I167205,I167222,I166919,I167253,I167270,I167296,I167304,I166907,I166925,I167349,I167366,I166928,I166913,I166922,I166931,I167469,I167495,I167503,I167520,I167546,I167437,I167568,I167594,I167602,I167619,I167645,I167461,I167667,I167443,I167707,I167724,I167732,I167749,I167446,I167780,I167797,I167823,I167831,I167434,I167452,I167876,I167893,I167455,I167440,I167449,I167458,I167996,I168022,I168030,I168047,I168073,I167964,I168095,I168121,I168129,I168146,I168172,I167988,I168194,I167970,I168234,I168251,I168259,I168276,I167973,I168307,I168324,I168350,I168358,I167961,I167979,I168403,I168420,I167982,I167967,I167976,I167985,I168523,I669408,I168549,I168557,I669405,I669396,I168574,I669393,I168600,I168491,I168622,I669402,I168648,I168656,I669411,I168673,I168699,I168515,I168721,I168497,I669414,I168761,I168778,I168786,I168803,I168500,I168834,I669399,I168851,I669417,I168877,I168885,I168488,I168506,I168930,I168947,I168509,I168494,I168503,I168512,I169050,I421817,I169076,I169084,I421808,I421823,I169101,I421829,I169127,I169149,I421814,I169175,I169183,I169200,I169226,I169248,I421811,I169288,I169305,I169313,I169330,I169361,I421805,I421820,I169378,I169404,I169412,I169457,I421826,I169474,I169577,I498971,I169603,I169611,I498968,I498986,I169628,I498977,I169654,I169676,I498992,I169702,I169710,I498974,I169727,I169753,I169775,I498980,I169815,I169832,I169840,I169857,I169888,I498995,I169905,I498983,I169931,I169939,I169984,I498989,I170001,I170104,I373843,I170130,I170138,I373834,I373849,I170155,I373855,I170181,I170203,I373840,I170229,I170237,I170254,I170280,I170302,I373837,I170342,I170359,I170367,I170384,I170415,I373831,I373846,I170432,I170458,I170466,I170511,I373852,I170528,I170631,I675188,I170657,I170665,I675185,I675176,I170682,I675173,I170708,I170599,I170730,I675182,I170756,I170764,I675191,I170781,I170807,I170623,I170829,I170605,I675194,I170869,I170886,I170894,I170911,I170608,I170942,I675179,I170959,I675197,I170985,I170993,I170596,I170614,I171038,I171055,I170617,I170602,I170611,I170620,I171158,I525457,I171184,I171192,I525454,I525472,I171209,I525463,I171235,I171126,I171257,I525478,I171283,I171291,I525460,I171308,I171334,I171150,I171356,I171132,I525466,I171396,I171413,I171421,I171438,I171135,I171469,I525481,I171486,I525469,I171512,I171520,I171123,I171141,I171565,I525475,I171582,I171144,I171129,I171138,I171147,I171685,I569963,I171711,I171719,I569960,I171736,I569972,I171762,I171653,I171784,I171810,I171818,I569978,I171835,I171861,I171677,I171883,I171659,I569966,I171923,I171940,I171948,I171965,I171662,I171996,I569975,I569981,I172013,I172039,I172047,I171650,I171668,I172092,I569969,I172109,I171671,I171656,I171665,I171674,I172212,I486051,I172238,I172246,I486048,I486066,I172263,I486057,I172289,I172311,I486072,I172337,I172345,I486054,I172362,I172388,I172410,I486060,I172450,I172467,I172475,I172492,I172523,I486075,I172540,I486063,I172566,I172574,I172619,I486069,I172636,I172739,I726959,I172765,I172773,I726938,I172790,I726965,I172816,I172707,I172838,I726953,I172864,I172872,I726956,I172889,I172915,I172731,I172937,I172713,I726947,I172977,I172994,I173002,I173019,I172716,I173050,I726944,I726941,I173067,I726962,I173093,I173101,I172704,I172722,I173146,I726950,I173163,I172725,I172710,I172719,I172728,I173266,I173292,I173300,I173317,I173343,I173365,I173391,I173399,I173416,I173442,I173464,I173504,I173521,I173529,I173546,I173577,I173594,I173620,I173628,I173673,I173690,I173793,I313734,I173819,I173827,I313719,I313722,I173844,I313737,I173870,I173892,I313731,I173918,I173926,I173943,I173969,I173991,I313728,I174031,I174048,I174056,I174073,I174104,I313743,I174121,I313740,I174147,I174155,I174200,I313725,I174217,I174320,I384825,I174346,I174354,I384816,I384831,I174371,I384837,I174397,I174288,I174419,I384822,I174445,I174453,I174470,I174496,I174312,I174518,I174294,I384819,I174558,I174575,I174583,I174600,I174297,I174631,I384813,I384828,I174648,I174674,I174682,I174285,I174303,I174727,I384834,I174744,I174306,I174291,I174300,I174309,I174847,I632945,I174873,I174881,I632960,I174898,I632963,I174924,I174815,I174946,I632969,I174972,I174980,I632951,I174997,I175023,I174839,I175045,I174821,I632948,I175085,I175102,I175110,I175127,I174824,I175158,I632954,I175175,I632966,I175201,I175209,I174812,I174830,I175254,I632957,I175271,I174833,I174818,I174827,I174836,I175374,I398119,I175400,I175408,I398110,I398125,I175425,I398131,I175451,I175342,I175473,I398116,I175499,I175507,I175524,I175550,I175366,I175572,I175348,I398113,I175612,I175629,I175637,I175654,I175351,I175685,I398107,I398122,I175702,I175728,I175736,I175339,I175357,I175781,I398128,I175798,I175360,I175345,I175354,I175363,I175901,I651255,I175927,I175935,I651237,I651261,I175952,I651252,I175978,I175869,I176000,I651258,I176026,I176034,I651246,I176051,I176077,I175893,I176099,I175875,I176139,I176156,I176164,I176181,I175878,I176212,I651243,I651240,I176229,I651249,I176255,I176263,I175866,I175884,I176308,I176325,I175887,I175872,I175881,I175890,I176428,I377311,I176454,I176462,I377302,I377317,I176479,I377323,I176505,I176396,I176527,I377308,I176553,I176561,I176578,I176604,I176420,I176626,I176402,I377305,I176666,I176683,I176691,I176708,I176405,I176739,I377299,I377314,I176756,I176782,I176790,I176393,I176411,I176835,I377320,I176852,I176414,I176399,I176408,I176417,I176955,I373265,I176981,I176989,I373256,I373271,I177006,I373277,I177032,I176923,I177054,I373262,I177080,I177088,I177105,I177131,I176947,I177153,I176929,I373259,I177193,I177210,I177218,I177235,I176932,I177266,I373253,I373268,I177283,I177309,I177317,I176920,I176938,I177362,I373274,I177379,I176941,I176926,I176935,I176944,I177482,I630055,I177508,I177516,I630070,I177533,I630073,I177559,I177450,I177581,I630079,I177607,I177615,I630061,I177632,I177658,I177474,I177680,I177456,I630058,I177720,I177737,I177745,I177762,I177459,I177793,I630064,I177810,I630076,I177836,I177844,I177447,I177465,I177889,I630067,I177906,I177468,I177453,I177462,I177471,I178009,I704349,I178035,I178043,I704328,I178060,I704355,I178086,I177977,I178108,I704343,I178134,I178142,I704346,I178159,I178185,I178001,I178207,I177983,I704337,I178247,I178264,I178272,I178289,I177986,I178320,I704334,I704331,I178337,I704352,I178363,I178371,I177974,I177992,I178416,I704340,I178433,I177995,I177980,I177989,I177998,I178536,I485405,I178562,I178570,I485402,I485420,I178587,I485411,I178613,I178504,I178635,I485426,I178661,I178669,I485408,I178686,I178712,I178528,I178734,I178510,I485414,I178774,I178791,I178799,I178816,I178513,I178847,I485429,I178864,I485417,I178890,I178898,I178501,I178519,I178943,I485423,I178960,I178522,I178507,I178516,I178525,I179063,I430750,I179089,I179097,I430753,I430747,I179114,I430759,I179140,I179031,I179162,I430762,I179188,I179196,I179213,I179239,I179055,I179261,I179037,I430765,I179301,I179318,I179326,I179343,I179040,I179374,I430756,I179391,I179417,I179425,I179028,I179046,I179470,I430768,I179487,I179049,I179034,I179043,I179052,I179590,I400431,I179616,I179624,I400422,I400437,I179641,I400443,I179667,I179558,I179689,I400428,I179715,I179723,I179740,I179766,I179582,I179788,I179564,I400425,I179828,I179845,I179853,I179870,I179567,I179901,I400419,I400434,I179918,I179944,I179952,I179555,I179573,I179997,I400440,I180014,I179576,I179561,I179570,I179579,I180117,I437074,I180143,I180151,I437077,I437071,I180168,I437083,I180194,I180085,I180216,I437086,I180242,I180250,I180267,I180293,I180109,I180315,I180091,I437089,I180355,I180372,I180380,I180397,I180094,I180428,I437080,I180445,I180471,I180479,I180082,I180100,I180524,I437092,I180541,I180103,I180088,I180097,I180106,I180644,I534501,I180670,I180678,I534498,I534516,I180695,I534507,I180721,I180612,I180743,I534522,I180769,I180777,I534504,I180794,I180820,I180636,I180842,I180618,I534510,I180882,I180899,I180907,I180924,I180621,I180955,I534525,I180972,I534513,I180998,I181006,I180609,I180627,I181051,I534519,I181068,I180630,I180615,I180624,I180633,I181171,I316046,I181197,I181205,I316031,I316034,I181222,I316049,I181248,I181270,I316043,I181296,I181304,I181321,I181347,I181369,I316040,I181409,I181426,I181434,I181451,I181482,I316055,I181499,I316052,I181525,I181533,I181578,I316037,I181595,I181698,I391761,I181724,I181732,I391752,I391767,I181749,I391773,I181775,I181666,I181797,I391758,I181823,I181831,I181848,I181874,I181690,I181896,I181672,I391755,I181936,I181953,I181961,I181978,I181675,I182009,I391749,I391764,I182026,I182052,I182060,I181663,I181681,I182105,I391770,I182122,I181684,I181669,I181678,I181687,I182225,I543596,I182251,I182259,I543593,I182276,I543605,I182302,I182193,I182324,I182350,I182358,I543611,I182375,I182401,I182217,I182423,I182199,I543599,I182463,I182480,I182488,I182505,I182202,I182536,I543608,I543614,I182553,I182579,I182587,I182190,I182208,I182632,I543602,I182649,I182211,I182196,I182205,I182214,I182752,I628321,I182778,I182786,I628336,I182803,I628339,I182829,I182851,I628345,I182877,I182885,I628327,I182902,I182928,I182950,I628324,I182990,I183007,I183015,I183032,I183063,I628330,I183080,I628342,I183106,I183114,I183159,I628333,I183176,I183279,I399275,I183305,I183313,I399266,I399281,I183330,I399287,I183356,I183378,I399272,I183404,I183412,I183429,I183455,I183477,I399269,I183517,I183534,I183542,I183559,I183590,I399263,I399278,I183607,I183633,I183641,I183686,I399284,I183703,I183806,I616183,I183832,I183840,I616198,I183857,I616201,I183883,I183774,I183905,I616207,I183931,I183939,I616189,I183956,I183982,I183798,I184004,I183780,I616186,I184044,I184061,I184069,I184086,I183783,I184117,I616192,I184134,I616204,I184160,I184168,I183771,I183789,I184213,I616195,I184230,I183792,I183777,I183786,I183795,I184333,I575723,I184359,I184367,I575738,I184384,I575741,I184410,I184301,I184432,I575747,I184458,I184466,I575729,I184483,I184509,I184325,I184531,I184307,I575726,I184571,I184588,I184596,I184613,I184310,I184644,I575732,I184661,I575744,I184687,I184695,I184298,I184316,I184740,I575735,I184757,I184319,I184304,I184313,I184322,I184860,I617339,I184886,I184894,I617354,I184911,I617357,I184937,I184828,I184959,I617363,I184985,I184993,I617345,I185010,I185036,I184852,I185058,I184834,I617342,I185098,I185115,I185123,I185140,I184837,I185171,I617348,I185188,I617360,I185214,I185222,I184825,I184843,I185267,I617351,I185284,I184846,I184831,I184840,I184849,I185387,I575145,I185413,I185421,I575160,I185438,I575163,I185464,I185355,I185486,I575169,I185512,I185520,I575151,I185537,I185563,I185379,I185585,I185361,I575148,I185625,I185642,I185650,I185667,I185364,I185698,I575154,I185715,I575166,I185741,I185749,I185352,I185370,I185794,I575157,I185811,I185373,I185358,I185367,I185376,I185914,I329340,I185940,I185948,I329325,I329328,I185965,I329343,I185991,I185882,I186013,I329337,I186039,I186047,I186064,I186090,I185906,I186112,I185888,I329334,I186152,I186169,I186177,I186194,I185891,I186225,I329349,I186242,I329346,I186268,I186276,I185879,I185897,I186321,I329331,I186338,I185900,I185885,I185894,I185903,I186441,I320670,I186467,I186475,I320655,I320658,I186492,I320673,I186518,I186409,I186540,I320667,I186566,I186574,I186591,I186617,I186433,I186639,I186415,I320664,I186679,I186696,I186704,I186721,I186418,I186752,I320679,I186769,I320676,I186795,I186803,I186406,I186424,I186848,I320661,I186865,I186427,I186412,I186421,I186430,I186968,I186994,I187002,I187019,I187045,I186936,I187067,I187093,I187101,I187118,I187144,I186960,I187166,I186942,I187206,I187223,I187231,I187248,I186945,I187279,I187296,I187322,I187330,I186933,I186951,I187375,I187392,I186954,I186939,I186948,I186957,I187495,I468167,I187521,I187529,I468170,I468164,I187546,I468176,I187572,I187463,I187594,I468179,I187620,I187628,I187645,I187671,I187487,I187693,I187469,I468182,I187733,I187750,I187758,I187775,I187472,I187806,I468173,I187823,I187849,I187857,I187460,I187478,I187902,I468185,I187919,I187481,I187466,I187475,I187484,I188022,I290296,I188048,I188056,I290308,I188073,I290293,I188099,I187990,I188121,I290317,I188147,I188155,I290314,I188172,I188198,I188014,I188220,I187996,I290305,I188260,I188277,I188285,I188302,I187999,I188333,I290302,I188350,I290311,I188376,I188384,I187987,I188005,I188429,I290299,I188446,I188008,I187993,I188002,I188011,I188549,I714464,I188575,I188583,I714443,I188600,I714470,I188626,I188517,I188648,I714458,I188674,I188682,I714461,I188699,I188725,I188541,I188747,I188523,I714452,I188787,I188804,I188812,I188829,I188526,I188860,I714449,I714446,I188877,I714467,I188903,I188911,I188514,I188532,I188956,I714455,I188973,I188535,I188520,I188529,I188538,I189076,I189102,I189110,I189127,I189153,I189044,I189175,I189201,I189209,I189226,I189252,I189068,I189274,I189050,I189314,I189331,I189339,I189356,I189053,I189387,I189404,I189430,I189438,I189041,I189059,I189483,I189500,I189062,I189047,I189056,I189065,I189603,I642007,I189629,I189637,I641989,I642013,I189654,I642004,I189680,I189702,I642010,I189728,I189736,I641998,I189753,I189779,I189801,I189841,I189858,I189866,I189883,I189914,I641995,I641992,I189931,I642001,I189957,I189965,I190010,I190027,I190130,I478945,I190156,I190164,I478942,I478960,I190181,I478951,I190207,I190098,I190229,I478966,I190255,I190263,I478948,I190280,I190306,I190122,I190328,I190104,I478954,I190368,I190385,I190393,I190410,I190107,I190441,I478969,I190458,I478957,I190484,I190492,I190095,I190113,I190537,I478963,I190554,I190116,I190101,I190110,I190119,I190657,I619073,I190683,I190691,I619088,I190708,I619091,I190734,I190625,I190756,I619097,I190782,I190790,I619079,I190807,I190833,I190649,I190855,I190631,I619076,I190895,I190912,I190920,I190937,I190634,I190968,I619082,I190985,I619094,I191011,I191019,I190622,I190640,I191064,I619085,I191081,I190643,I190628,I190637,I190646,I191184,I639831,I191210,I191218,I639813,I639837,I191235,I639828,I191261,I191152,I191283,I639834,I191309,I191317,I639822,I191334,I191360,I191176,I191382,I191158,I191422,I191439,I191447,I191464,I191161,I191495,I639819,I639816,I191512,I639825,I191538,I191546,I191149,I191167,I191591,I191608,I191170,I191155,I191164,I191173,I191711,I302174,I191737,I191745,I302159,I302162,I191762,I302177,I191788,I191810,I302171,I191836,I191844,I191861,I191887,I191909,I302168,I191949,I191966,I191974,I191991,I192022,I302183,I192039,I302180,I192065,I192073,I192118,I302165,I192135,I192238,I655607,I192264,I192272,I655589,I655613,I192289,I655604,I192315,I192206,I192337,I655610,I192363,I192371,I655598,I192388,I192414,I192230,I192436,I192212,I192476,I192493,I192501,I192518,I192215,I192549,I655595,I655592,I192566,I655601,I192592,I192600,I192203,I192221,I192645,I192662,I192224,I192209,I192218,I192227,I192765,I535147,I192791,I192799,I535144,I535162,I192816,I535153,I192842,I192733,I192864,I535168,I192890,I192898,I535150,I192915,I192941,I192757,I192963,I192739,I535156,I193003,I193020,I193028,I193045,I192742,I193076,I535171,I193093,I535159,I193119,I193127,I192730,I192748,I193172,I535165,I193189,I192751,I192736,I192745,I192754,I193292,I729934,I193318,I193326,I729913,I193343,I729940,I193369,I193260,I193391,I729928,I193417,I193425,I729931,I193442,I193468,I193284,I193490,I193266,I729922,I193530,I193547,I193555,I193572,I193269,I193603,I729919,I729916,I193620,I729937,I193646,I193654,I193257,I193275,I193699,I729925,I193716,I193278,I193263,I193272,I193281,I193819,I193845,I193853,I193870,I193896,I193787,I193918,I193944,I193952,I193969,I193995,I193811,I194017,I193793,I194057,I194074,I194082,I194099,I193796,I194130,I194147,I194173,I194181,I193784,I193802,I194226,I194243,I193805,I193790,I193799,I193808,I194346,I301596,I194372,I194380,I301581,I301584,I194397,I301599,I194423,I194314,I194445,I301593,I194471,I194479,I194496,I194522,I194338,I194544,I194320,I301590,I194584,I194601,I194609,I194626,I194323,I194657,I301605,I194674,I301602,I194700,I194708,I194311,I194329,I194753,I301587,I194770,I194332,I194317,I194326,I194335,I194873,I194899,I194907,I194924,I194950,I194841,I194972,I194998,I195006,I195023,I195049,I194865,I195071,I194847,I195111,I195128,I195136,I195153,I194850,I195184,I195201,I195227,I195235,I194838,I194856,I195280,I195297,I194859,I194844,I194853,I194862,I195400,I309688,I195426,I195434,I309673,I309676,I195451,I309691,I195477,I195499,I309685,I195525,I195533,I195550,I195576,I195598,I309682,I195638,I195655,I195663,I195680,I195711,I309697,I195728,I309694,I195754,I195762,I195807,I309679,I195824,I195927,I324138,I195953,I195961,I324123,I324126,I195978,I324141,I196004,I195895,I196026,I324135,I196052,I196060,I196077,I196103,I195919,I196125,I195901,I324132,I196165,I196182,I196190,I196207,I195904,I196238,I324147,I196255,I324144,I196281,I196289,I195892,I195910,I196334,I324129,I196351,I195913,I195898,I195907,I195916,I196454,I343212,I196480,I196488,I343197,I343200,I196505,I343215,I196531,I196553,I343209,I196579,I196587,I196604,I196630,I196652,I343206,I196692,I196709,I196717,I196734,I196765,I343221,I196782,I343218,I196808,I196816,I196861,I343203,I196878,I196981,I197007,I197015,I197032,I197058,I196949,I197080,I197106,I197114,I197131,I197157,I196973,I197179,I196955,I197219,I197236,I197244,I197261,I196958,I197292,I197309,I197335,I197343,I196946,I196964,I197388,I197405,I196967,I196952,I196961,I196970,I197508,I709704,I197534,I197542,I709683,I197559,I709710,I197585,I197476,I197607,I709698,I197633,I197641,I709701,I197658,I197684,I197500,I197706,I197482,I709692,I197746,I197763,I197771,I197788,I197485,I197819,I709689,I709686,I197836,I709707,I197862,I197870,I197473,I197491,I197915,I709695,I197932,I197494,I197479,I197488,I197497,I198035,I198061,I198069,I198086,I198112,I198003,I198134,I198160,I198168,I198185,I198211,I198027,I198233,I198009,I198273,I198290,I198298,I198315,I198012,I198346,I198363,I198389,I198397,I198000,I198018,I198442,I198459,I198021,I198006,I198015,I198024,I198562,I483467,I198588,I198596,I483464,I483482,I198613,I483473,I198639,I198661,I483488,I198687,I198695,I483470,I198712,I198738,I198760,I483476,I198800,I198817,I198825,I198842,I198873,I483491,I198890,I483479,I198916,I198924,I198969,I483485,I198986,I199089,I460789,I199115,I199123,I460792,I460786,I199140,I460798,I199166,I199188,I460801,I199214,I199222,I199239,I199265,I199287,I460804,I199327,I199344,I199352,I199369,I199400,I460795,I199417,I199443,I199451,I199496,I460807,I199513,I199616,I199642,I199650,I199667,I199693,I199584,I199715,I199741,I199749,I199766,I199792,I199608,I199814,I199590,I199854,I199871,I199879,I199896,I199593,I199927,I199944,I199970,I199978,I199581,I199599,I200023,I200040,I199602,I199587,I199596,I199605,I200143,I200169,I200177,I200194,I200220,I200111,I200242,I200268,I200276,I200293,I200319,I200135,I200341,I200117,I200381,I200398,I200406,I200423,I200120,I200454,I200471,I200497,I200505,I200108,I200126,I200550,I200567,I200129,I200114,I200123,I200132,I200670,I298031,I200696,I200704,I298043,I200721,I298028,I200747,I200638,I200769,I298052,I200795,I200803,I298049,I200820,I200846,I200662,I200868,I200644,I298040,I200908,I200925,I200933,I200950,I200647,I200981,I298037,I200998,I298046,I201024,I201032,I200635,I200653,I201077,I298034,I201094,I200656,I200641,I200650,I200659,I201197,I420083,I201223,I201231,I420074,I420089,I201248,I420095,I201274,I201296,I420080,I201322,I201330,I201347,I201373,I201395,I420077,I201435,I201452,I201460,I201477,I201508,I420071,I420086,I201525,I201551,I201559,I201604,I420092,I201621,I201724,I608669,I201750,I201758,I608684,I201775,I608687,I201801,I201823,I608693,I201849,I201857,I608675,I201874,I201900,I201922,I608672,I201962,I201979,I201987,I202004,I202035,I608678,I202052,I608690,I202078,I202086,I202131,I608681,I202148,I202251,I470275,I202277,I202285,I470278,I470272,I202302,I470284,I202328,I202219,I202350,I470287,I202376,I202384,I202401,I202427,I202243,I202449,I202225,I470290,I202489,I202506,I202514,I202531,I202228,I202562,I470281,I202579,I202605,I202613,I202216,I202234,I202658,I470293,I202675,I202237,I202222,I202231,I202240,I202778,I677500,I202804,I202812,I677497,I677488,I202829,I677485,I202855,I202746,I202877,I677494,I202903,I202911,I677503,I202928,I202954,I202770,I202976,I202752,I677506,I203016,I203033,I203041,I203058,I202755,I203089,I677491,I203106,I677509,I203132,I203140,I202743,I202761,I203185,I203202,I202764,I202749,I202758,I202767,I203305,I323560,I203331,I203339,I323545,I323548,I203356,I323563,I203382,I203273,I203404,I323557,I203430,I203438,I203455,I203481,I203297,I203503,I203279,I323554,I203543,I203560,I203568,I203585,I203282,I203616,I323569,I203633,I323566,I203659,I203667,I203270,I203288,I203712,I323551,I203729,I203291,I203276,I203285,I203294,I203832,I396963,I203858,I203866,I396954,I396969,I203883,I396975,I203909,I203800,I203931,I396960,I203957,I203965,I203982,I204008,I203824,I204030,I203806,I396957,I204070,I204087,I204095,I204112,I203809,I204143,I396951,I396966,I204160,I204186,I204194,I203797,I203815,I204239,I396972,I204256,I203818,I203803,I203812,I203821,I204359,I204385,I204393,I204410,I204436,I204327,I204458,I204484,I204492,I204509,I204535,I204351,I204557,I204333,I204597,I204614,I204622,I204639,I204336,I204670,I204687,I204713,I204721,I204324,I204342,I204766,I204783,I204345,I204330,I204339,I204348,I204886,I204912,I204920,I204937,I204963,I204854,I204985,I205011,I205019,I205036,I205062,I204878,I205084,I204860,I205124,I205141,I205149,I205166,I204863,I205197,I205214,I205240,I205248,I204851,I204869,I205293,I205310,I204872,I204857,I204866,I204875,I205413,I379623,I205439,I205447,I379614,I379629,I205464,I379635,I205490,I205381,I205512,I379620,I205538,I205546,I205563,I205589,I205405,I205611,I205387,I379617,I205651,I205668,I205676,I205693,I205390,I205724,I379611,I379626,I205741,I205767,I205775,I205378,I205396,I205820,I379632,I205837,I205399,I205384,I205393,I205402,I205940,I450776,I205966,I205974,I450779,I450773,I205991,I450785,I206017,I205908,I206039,I450788,I206065,I206073,I206090,I206116,I205932,I206138,I205914,I450791,I206178,I206195,I206203,I206220,I205917,I206251,I450782,I206268,I206294,I206302,I205905,I205923,I206347,I450794,I206364,I205926,I205911,I205920,I205929,I206467,I604623,I206493,I206501,I604638,I206518,I604641,I206544,I206435,I206566,I604647,I206592,I206600,I604629,I206617,I206643,I206459,I206665,I206441,I604626,I206705,I206722,I206730,I206747,I206444,I206778,I604632,I206795,I604644,I206821,I206829,I206432,I206450,I206874,I604635,I206891,I206453,I206438,I206447,I206456,I206994,I465005,I207020,I207028,I465008,I465002,I207045,I465014,I207071,I206962,I207093,I465017,I207119,I207127,I207144,I207170,I206986,I207192,I206968,I465020,I207232,I207249,I207257,I207274,I206971,I207305,I465011,I207322,I207348,I207356,I206959,I206977,I207401,I465023,I207418,I206980,I206965,I206974,I206983,I207521,I439182,I207547,I207555,I439185,I439179,I207572,I439191,I207598,I207489,I207620,I439194,I207646,I207654,I207671,I207697,I207513,I207719,I207495,I439197,I207759,I207776,I207784,I207801,I207498,I207832,I439188,I207849,I207875,I207883,I207486,I207504,I207928,I439200,I207945,I207507,I207492,I207501,I207510,I208048,I436020,I208074,I208082,I436023,I436017,I208099,I436029,I208125,I208016,I208147,I436032,I208173,I208181,I208198,I208224,I208040,I208246,I208022,I436035,I208286,I208303,I208311,I208328,I208025,I208359,I436026,I208376,I208402,I208410,I208013,I208031,I208455,I436038,I208472,I208034,I208019,I208028,I208037,I208575,I569402,I208601,I208609,I569399,I208626,I569411,I208652,I208543,I208674,I208700,I208708,I569417,I208725,I208751,I208567,I208773,I208549,I569405,I208813,I208830,I208838,I208855,I208552,I208886,I569414,I569420,I208903,I208929,I208937,I208540,I208558,I208982,I569408,I208999,I208561,I208546,I208555,I208564,I209102,I368063,I209128,I209136,I368054,I368069,I209153,I368075,I209179,I209201,I368060,I209227,I209235,I209252,I209278,I209300,I368057,I209340,I209357,I209365,I209382,I209413,I368051,I368066,I209430,I209456,I209464,I209509,I368072,I209526,I209629,I429696,I209655,I209663,I429699,I429693,I209680,I429705,I209706,I209728,I429708,I209754,I209762,I209779,I209805,I209827,I429711,I209867,I209884,I209892,I209909,I209940,I429702,I209957,I209983,I209991,I210036,I429714,I210053,I210156,I606357,I210182,I210190,I606372,I210207,I606375,I210233,I210124,I210255,I606381,I210281,I210289,I606363,I210306,I210332,I210148,I210354,I210130,I606360,I210394,I210411,I210419,I210436,I210133,I210467,I606366,I210484,I606378,I210510,I210518,I210121,I210139,I210563,I606369,I210580,I210142,I210127,I210136,I210145,I210683,I653975,I210709,I210717,I653957,I653981,I210734,I653972,I210760,I210782,I653978,I210808,I210816,I653966,I210833,I210859,I210881,I210921,I210938,I210946,I210963,I210994,I653963,I653960,I211011,I653969,I211037,I211045,I211090,I211107,I211210,I282561,I211236,I211244,I282573,I211261,I282558,I211287,I211178,I211309,I282582,I211335,I211343,I282579,I211360,I211386,I211202,I211408,I211184,I282570,I211448,I211465,I211473,I211490,I211187,I211521,I282567,I211538,I282576,I211564,I211572,I211175,I211193,I211617,I282564,I211634,I211196,I211181,I211190,I211199,I211737,I545279,I211763,I211771,I545276,I211788,I545288,I211814,I211705,I211836,I211862,I211870,I545294,I211887,I211913,I211729,I211935,I211711,I545282,I211975,I211992,I212000,I212017,I211714,I212048,I545291,I545297,I212065,I212091,I212099,I211702,I211720,I212144,I545285,I212161,I211723,I211708,I211717,I211726,I212264,I291486,I212290,I212298,I291498,I212315,I291483,I212341,I212232,I212363,I291507,I212389,I212397,I291504,I212414,I212440,I212256,I212462,I212238,I291495,I212502,I212519,I212527,I212544,I212241,I212575,I291492,I212592,I291501,I212618,I212626,I212229,I212247,I212671,I291489,I212688,I212250,I212235,I212244,I212253,I212791,I346677,I212817,I212825,I346668,I346683,I212842,I346689,I212868,I212759,I212890,I346674,I212916,I212924,I212941,I212967,I212783,I212989,I212765,I346671,I213029,I213046,I213054,I213071,I212768,I213102,I346665,I346680,I213119,I213145,I213153,I212756,I212774,I213198,I346686,I213215,I212777,I212762,I212771,I212780,I213318,I338588,I213344,I213352,I338573,I338576,I213369,I338591,I213395,I213286,I213417,I338585,I213443,I213451,I213468,I213494,I213310,I213516,I213292,I338582,I213556,I213573,I213581,I213598,I213295,I213629,I338597,I213646,I338594,I213672,I213680,I213283,I213301,I213725,I338579,I213742,I213304,I213289,I213298,I213307,I213845,I294461,I213871,I213879,I294473,I213896,I294458,I213922,I213813,I213944,I294482,I213970,I213978,I294479,I213995,I214021,I213837,I214043,I213819,I294470,I214083,I214100,I214108,I214125,I213822,I214156,I294467,I214173,I294476,I214199,I214207,I213810,I213828,I214252,I294464,I214269,I213831,I213816,I213825,I213834,I214372,I333964,I214398,I214406,I333949,I333952,I214423,I333967,I214449,I214340,I214471,I333961,I214497,I214505,I214522,I214548,I214364,I214570,I214346,I333958,I214610,I214627,I214635,I214652,I214349,I214683,I333973,I214700,I333970,I214726,I214734,I214337,I214355,I214779,I333955,I214796,I214358,I214343,I214352,I214361,I214899,I214925,I214933,I214950,I214976,I214998,I215024,I215032,I215049,I215075,I215097,I215137,I215154,I215162,I215179,I215210,I215227,I215253,I215261,I215306,I215323,I215426,I215452,I215460,I215477,I215503,I215394,I215525,I215551,I215559,I215576,I215602,I215418,I215624,I215400,I215664,I215681,I215689,I215706,I215403,I215737,I215754,I215780,I215788,I215391,I215409,I215833,I215850,I215412,I215397,I215406,I215415,I215953,I464478,I215979,I215987,I464481,I464475,I216004,I464487,I216030,I215921,I216052,I464490,I216078,I216086,I216103,I216129,I215945,I216151,I215927,I464493,I216191,I216208,I216216,I216233,I215930,I216264,I464484,I216281,I216307,I216315,I215918,I215936,I216360,I464496,I216377,I215939,I215924,I215933,I215942,I216480,I216506,I216514,I216531,I216557,I216448,I216579,I216605,I216613,I216630,I216656,I216472,I216678,I216454,I216718,I216735,I216743,I216760,I216457,I216791,I216808,I216834,I216842,I216445,I216463,I216887,I216904,I216466,I216451,I216460,I216469,I217007,I700184,I217033,I217041,I700163,I217058,I700190,I217084,I217106,I700178,I217132,I217140,I700181,I217157,I217183,I217205,I700172,I217245,I217262,I217270,I217287,I217318,I700169,I700166,I217335,I700187,I217361,I217369,I217414,I700175,I217431,I217534,I217560,I217568,I217585,I217611,I217633,I217659,I217667,I217684,I217710,I217732,I217772,I217789,I217797,I217814,I217845,I217862,I217888,I217896,I217941,I217958,I218061,I218087,I218095,I218112,I218138,I218029,I218160,I218186,I218194,I218211,I218237,I218053,I218259,I218035,I218299,I218316,I218324,I218341,I218038,I218372,I218389,I218415,I218423,I218026,I218044,I218468,I218485,I218047,I218032,I218041,I218050,I218588,I709109,I218614,I218622,I709088,I218639,I709115,I218665,I218687,I709103,I218713,I218721,I709106,I218738,I218764,I218786,I709097,I218826,I218843,I218851,I218868,I218899,I709094,I709091,I218916,I709112,I218942,I218950,I218995,I709100,I219012,I219115,I380201,I219141,I219149,I380192,I380207,I219166,I380213,I219192,I219083,I219214,I380198,I219240,I219248,I219265,I219291,I219107,I219313,I219089,I380195,I219353,I219370,I219378,I219395,I219092,I219426,I380189,I380204,I219443,I219469,I219477,I219080,I219098,I219522,I380210,I219539,I219101,I219086,I219095,I219104,I219642,I643639,I219668,I219676,I643621,I643645,I219693,I643636,I219719,I219610,I219741,I643642,I219767,I219775,I643630,I219792,I219818,I219634,I219840,I219616,I219880,I219897,I219905,I219922,I219619,I219953,I643627,I643624,I219970,I643633,I219996,I220004,I219607,I219625,I220049,I220066,I219628,I219613,I219622,I219631,I220169,I667674,I220195,I220203,I667671,I667662,I220220,I667659,I220246,I220137,I220268,I667668,I220294,I220302,I667677,I220319,I220345,I220161,I220367,I220143,I667680,I220407,I220424,I220432,I220449,I220146,I220480,I667665,I220497,I667683,I220523,I220531,I220134,I220152,I220576,I220593,I220155,I220140,I220149,I220158,I220696,I237860,I220722,I220730,I237872,I237851,I220747,I237875,I220773,I220795,I237866,I220821,I220829,I237848,I220846,I220872,I220894,I237863,I220934,I220951,I220959,I220976,I221007,I237854,I221024,I237857,I221050,I221058,I221103,I237869,I221120,I221223,I221249,I221257,I221274,I221300,I221322,I221348,I221356,I221373,I221399,I221421,I221461,I221478,I221486,I221503,I221534,I221551,I221577,I221585,I221630,I221647,I221750,I266692,I221776,I221784,I266704,I266683,I221801,I266707,I221827,I221849,I266698,I221875,I221883,I266680,I221900,I221926,I221948,I266695,I221988,I222005,I222013,I222030,I222061,I266686,I222078,I266689,I222104,I222112,I222157,I266701,I222174,I222277,I406789,I222303,I222311,I406780,I406795,I222328,I406801,I222354,I222245,I222376,I406786,I222402,I222410,I222427,I222453,I222269,I222475,I222251,I406783,I222515,I222532,I222540,I222557,I222254,I222588,I406777,I406792,I222605,I222631,I222639,I222242,I222260,I222684,I406798,I222701,I222263,I222248,I222257,I222266,I222804,I626587,I222830,I222838,I626602,I222855,I626605,I222881,I222772,I222903,I626611,I222929,I222937,I626593,I222954,I222980,I222796,I223002,I222778,I626590,I223042,I223059,I223067,I223084,I222781,I223115,I626596,I223132,I626608,I223158,I223166,I222769,I222787,I223211,I626599,I223228,I222790,I222775,I222784,I222793,I223331,I223357,I223365,I223382,I223408,I223299,I223430,I223456,I223464,I223481,I223507,I223323,I223529,I223305,I223569,I223586,I223594,I223611,I223308,I223642,I223659,I223685,I223693,I223296,I223314,I223738,I223755,I223317,I223302,I223311,I223320,I223858,I223884,I223892,I223909,I223935,I223957,I223983,I223991,I224008,I224034,I224056,I224096,I224113,I224121,I224138,I224169,I224186,I224212,I224220,I224265,I224282,I224385,I259620,I224411,I224419,I259632,I259611,I224436,I259635,I224462,I224484,I259626,I224510,I224518,I259608,I224535,I224561,I224583,I259623,I224623,I224640,I224648,I224665,I224696,I259614,I224713,I259617,I224739,I224747,I224792,I259629,I224809,I224912,I271588,I224938,I224946,I271600,I271579,I224963,I271603,I224989,I224880,I225011,I271594,I225037,I225045,I271576,I225062,I225088,I224904,I225110,I224886,I271591,I225150,I225167,I225175,I225192,I224889,I225223,I271582,I225240,I271585,I225266,I225274,I224877,I224895,I225319,I271597,I225336,I224898,I224883,I224892,I224901,I225439,I586127,I225465,I225473,I586142,I225490,I586145,I225516,I225538,I586151,I225564,I225572,I586133,I225589,I225615,I225637,I586130,I225677,I225694,I225702,I225719,I225750,I586136,I225767,I586148,I225793,I225801,I225846,I586139,I225863,I225966,I564914,I225992,I226000,I564911,I226017,I564923,I226043,I225934,I226065,I226091,I226099,I564929,I226116,I226142,I225958,I226164,I225940,I564917,I226204,I226221,I226229,I226246,I225943,I226277,I564926,I564932,I226294,I226320,I226328,I225931,I225949,I226373,I564920,I226390,I225952,I225937,I225946,I225955,I226493,I275396,I226519,I226527,I275408,I275387,I226544,I275411,I226570,I226592,I275402,I226618,I226626,I275384,I226643,I226669,I226691,I275399,I226731,I226748,I226756,I226773,I226804,I275390,I226821,I275393,I226847,I226855,I226900,I275405,I226917,I227020,I227046,I227054,I227071,I227097,I226988,I227119,I227145,I227153,I227170,I227196,I227012,I227218,I226994,I227258,I227275,I227283,I227300,I226997,I227331,I227348,I227374,I227382,I226985,I227003,I227427,I227444,I227006,I226991,I227000,I227009,I227547,I650696,I227573,I227590,I227612,I227629,I650708,I650711,I227646,I650714,I227672,I227680,I650699,I227706,I227714,I650705,I227731,I650693,I227771,I227779,I227824,I650717,I227841,I650702,I227867,I227889,I227906,I227923,I227954,I227971,I228002,I228091,I578038,I228117,I228134,I228156,I228173,I578050,I228190,I578041,I228216,I228224,I578059,I228250,I228258,I578035,I228275,I578053,I228315,I228323,I228368,I578047,I578044,I228385,I578056,I228411,I228433,I228450,I228467,I228498,I228515,I228546,I228635,I351292,I228661,I228678,I228627,I228700,I228717,I351313,I351304,I228734,I228760,I228768,I351298,I228794,I228802,I351295,I228819,I228606,I351289,I228859,I228867,I228600,I228615,I228912,I351301,I228929,I351310,I228955,I228603,I228977,I228994,I229011,I228618,I229042,I229059,I351307,I228609,I229090,I228612,I228624,I228621,I229179,I229205,I229222,I229171,I229244,I229261,I229278,I229304,I229312,I229338,I229346,I229363,I229150,I229403,I229411,I229144,I229159,I229456,I229473,I229499,I229147,I229521,I229538,I229555,I229162,I229586,I229603,I229153,I229634,I229156,I229168,I229165,I229723,I390596,I229749,I229766,I229715,I229788,I229805,I390617,I390608,I229822,I229848,I229856,I390602,I229882,I229890,I390599,I229907,I229694,I390593,I229947,I229955,I229688,I229703,I230000,I390605,I230017,I390614,I230043,I229691,I230065,I230082,I230099,I229706,I230130,I230147,I390611,I229697,I230178,I229700,I229712,I229709,I230267,I432340,I230293,I230310,I230259,I230332,I230349,I432334,I432331,I230366,I432346,I230392,I230400,I230426,I230434,I432328,I230451,I230238,I230491,I230499,I230232,I230247,I230544,I432343,I432337,I230561,I230587,I230235,I230609,I230626,I230643,I230250,I230674,I230691,I432349,I230241,I230722,I230244,I230256,I230253,I230811,I230837,I230854,I230803,I230876,I230893,I230910,I230936,I230944,I230970,I230978,I230995,I230782,I231035,I231043,I230776,I230791,I231088,I231105,I231131,I230779,I231153,I231170,I231187,I230794,I231218,I231235,I230785,I231266,I230788,I230800,I230797,I231355,I231381,I231398,I231420,I231437,I231454,I231480,I231488,I231514,I231522,I231539,I231579,I231587,I231632,I231649,I231675,I231697,I231714,I231731,I231762,I231779,I231810,I231899,I546398,I231925,I231942,I231891,I231964,I231981,I546416,I231998,I546410,I232024,I232032,I546404,I232058,I232066,I546413,I232083,I231870,I546401,I232123,I232131,I231864,I231879,I232176,I546419,I232193,I232219,I231867,I232241,I232258,I232275,I231882,I232306,I232323,I546407,I231873,I232354,I231876,I231888,I231885,I232443,I232469,I232486,I232435,I232508,I232525,I232542,I232568,I232576,I232602,I232610,I232627,I232414,I232667,I232675,I232408,I232423,I232720,I232737,I232763,I232411,I232785,I232802,I232819,I232426,I232850,I232867,I232417,I232898,I232420,I232432,I232429,I232987,I427010,I233013,I233030,I232979,I233052,I233069,I427031,I427022,I233086,I233112,I233120,I427016,I233146,I233154,I427013,I233171,I232958,I427007,I233211,I233219,I232952,I232967,I233264,I427019,I233281,I427028,I233307,I232955,I233329,I233346,I233363,I232970,I233394,I233411,I427025,I232961,I233442,I232964,I232976,I232973,I233531,I233557,I233574,I233596,I233613,I233630,I233656,I233664,I233690,I233698,I233715,I233755,I233763,I233808,I233825,I233851,I233873,I233890,I233907,I233938,I233955,I233986,I234075,I716850,I234101,I234118,I234140,I234157,I716826,I716847,I234174,I716844,I234200,I234208,I716823,I234234,I234242,I716835,I234259,I716838,I234299,I234307,I234352,I716841,I716829,I234369,I716832,I234395,I234417,I234434,I234451,I234482,I234499,I234530,I234619,I333374,I234645,I234662,I234611,I234684,I234701,I333371,I333392,I234718,I333395,I234744,I234752,I333380,I234778,I234786,I333383,I234803,I234590,I333386,I234843,I234851,I234584,I234599,I234896,I333377,I234913,I333389,I234939,I234587,I234961,I234978,I234995,I234602,I235026,I235043,I234593,I235074,I234596,I234608,I234605,I235163,I235189,I235206,I235228,I235245,I235262,I235288,I235296,I235322,I235330,I235347,I235387,I235395,I235440,I235457,I235483,I235505,I235522,I235539,I235570,I235587,I235618,I235707,I668833,I235733,I235750,I235699,I235772,I235789,I668830,I668827,I235806,I668815,I235832,I235840,I668839,I235866,I235874,I668824,I235891,I235678,I668818,I235931,I235939,I235672,I235687,I235984,I668821,I236001,I668836,I236027,I235675,I236049,I236066,I236083,I235690,I236114,I236131,I235681,I236162,I235684,I235696,I235693,I236251,I236277,I236294,I236316,I236333,I236350,I236376,I236384,I236410,I236418,I236435,I236475,I236483,I236528,I236545,I236571,I236593,I236610,I236627,I236658,I236675,I236706,I236795,I236821,I236838,I236787,I236860,I236877,I236894,I236920,I236928,I236954,I236962,I236979,I236766,I237019,I237027,I236760,I236775,I237072,I237089,I237115,I236763,I237137,I237154,I237171,I236778,I237202,I237219,I236769,I237250,I236772,I236784,I236781,I237339,I237365,I237382,I237331,I237404,I237421,I237438,I237464,I237472,I237498,I237506,I237523,I237310,I237563,I237571,I237304,I237319,I237616,I237633,I237659,I237307,I237681,I237698,I237715,I237322,I237746,I237763,I237313,I237794,I237316,I237328,I237325,I237883,I237909,I237926,I237948,I237965,I237982,I238008,I238016,I238042,I238050,I238067,I238107,I238115,I238160,I238177,I238203,I238225,I238242,I238259,I238290,I238307,I238338,I238427,I719825,I238453,I238470,I238419,I238492,I238509,I719801,I719822,I238526,I719819,I238552,I238560,I719798,I238586,I238594,I719810,I238611,I238398,I719813,I238651,I238659,I238392,I238407,I238704,I719816,I719804,I238721,I719807,I238747,I238395,I238769,I238786,I238803,I238410,I238834,I238851,I238401,I238882,I238404,I238416,I238413,I238971,I238997,I239014,I238963,I239036,I239053,I239070,I239096,I239104,I239130,I239138,I239155,I238942,I239195,I239203,I238936,I238951,I239248,I239265,I239291,I238939,I239313,I239330,I239347,I238954,I239378,I239395,I238945,I239426,I238948,I238960,I238957,I239515,I679237,I239541,I239558,I239507,I239580,I239597,I679234,I679231,I239614,I679219,I239640,I239648,I679243,I239674,I239682,I679228,I239699,I239486,I679222,I239739,I239747,I239480,I239495,I239792,I679225,I239809,I679240,I239835,I239483,I239857,I239874,I239891,I239498,I239922,I239939,I239489,I239970,I239492,I239504,I239501,I240059,I507372,I240085,I240102,I240124,I240141,I507387,I507375,I240158,I507366,I240184,I240192,I507378,I240218,I240226,I507369,I240243,I507384,I240283,I240291,I240336,I507393,I507381,I240353,I507390,I240379,I240401,I240418,I240435,I240466,I240483,I240514,I240603,I240629,I240646,I240595,I240668,I240685,I240702,I240728,I240736,I240762,I240770,I240787,I240574,I240827,I240835,I240568,I240583,I240880,I240897,I240923,I240571,I240945,I240962,I240979,I240586,I241010,I241027,I240577,I241058,I240580,I240592,I240589,I241147,I517708,I241173,I241190,I241139,I241212,I241229,I517723,I517711,I241246,I517702,I241272,I241280,I517714,I241306,I241314,I517705,I241331,I241118,I517720,I241371,I241379,I241112,I241127,I241424,I517729,I517717,I241441,I517726,I241467,I241115,I241489,I241506,I241523,I241130,I241554,I241571,I241121,I241602,I241124,I241136,I241133,I241691,I361696,I241717,I241734,I241756,I241773,I361717,I361708,I241790,I241816,I241824,I361702,I241850,I241858,I361699,I241875,I361693,I241915,I241923,I241968,I361705,I241985,I361714,I242011,I242033,I242050,I242067,I242098,I242115,I361711,I242146,I242235,I242261,I242278,I242227,I242300,I242317,I242334,I242360,I242368,I242394,I242402,I242419,I242206,I242459,I242467,I242200,I242215,I242512,I242529,I242555,I242203,I242577,I242594,I242611,I242218,I242642,I242659,I242209,I242690,I242212,I242224,I242221,I242779,I412560,I242805,I242822,I242844,I242861,I412581,I412572,I242878,I242904,I242912,I412566,I242938,I242946,I412563,I242963,I412557,I243003,I243011,I243056,I412569,I243073,I412578,I243099,I243121,I243138,I243155,I243186,I243203,I412575,I243234,I243323,I243349,I243366,I243315,I243388,I243405,I243422,I243448,I243456,I243482,I243490,I243507,I243294,I243547,I243555,I243288,I243303,I243600,I243617,I243643,I243291,I243665,I243682,I243699,I243306,I243730,I243747,I243297,I243778,I243300,I243312,I243309,I243867,I423542,I243893,I243910,I243932,I243949,I423563,I423554,I243966,I243992,I244000,I423548,I244026,I244034,I423545,I244051,I423539,I244091,I244099,I244144,I423551,I244161,I423560,I244187,I244209,I244226,I244243,I244274,I244291,I423557,I244322,I244411,I244437,I244454,I244403,I244476,I244493,I244510,I244536,I244544,I244570,I244578,I244595,I244382,I244635,I244643,I244376,I244391,I244688,I244705,I244731,I244379,I244753,I244770,I244787,I244394,I244818,I244835,I244385,I244866,I244388,I244400,I244397,I244955,I573992,I244981,I244998,I244947,I245020,I245037,I574004,I245054,I573995,I245080,I245088,I574013,I245114,I245122,I573989,I245139,I244926,I574007,I245179,I245187,I244920,I244935,I245232,I574001,I573998,I245249,I574010,I245275,I244923,I245297,I245314,I245331,I244938,I245362,I245379,I244929,I245410,I244932,I244944,I244941,I245499,I245525,I245542,I245491,I245564,I245581,I245598,I245624,I245632,I245658,I245666,I245683,I245470,I245723,I245731,I245464,I245479,I245776,I245793,I245819,I245467,I245841,I245858,I245875,I245482,I245906,I245923,I245473,I245954,I245476,I245488,I245485,I246043,I246069,I246086,I246035,I246108,I246125,I246142,I246168,I246176,I246202,I246210,I246227,I246014,I246267,I246275,I246008,I246023,I246320,I246337,I246363,I246011,I246385,I246402,I246419,I246026,I246450,I246467,I246017,I246498,I246020,I246032,I246029,I246587,I690670,I246613,I246630,I246579,I246652,I246669,I690646,I690667,I246686,I690664,I246712,I246720,I690643,I246746,I246754,I690655,I246771,I246558,I690658,I246811,I246819,I246552,I246567,I246864,I690661,I690649,I246881,I690652,I246907,I246555,I246929,I246946,I246963,I246570,I246994,I247011,I246561,I247042,I246564,I246576,I246573,I247131,I247157,I247174,I247196,I247213,I247230,I247256,I247264,I247290,I247298,I247315,I247355,I247363,I247408,I247425,I247451,I247473,I247490,I247507,I247538,I247555,I247586,I247675,I247701,I247718,I247667,I247740,I247757,I247774,I247800,I247808,I247834,I247842,I247859,I247646,I247899,I247907,I247640,I247655,I247952,I247969,I247995,I247643,I248017,I248034,I248051,I247658,I248082,I248099,I247649,I248130,I247652,I247664,I247661,I248219,I248245,I248262,I248211,I248284,I248301,I248318,I248344,I248352,I248378,I248386,I248403,I248190,I248443,I248451,I248184,I248199,I248496,I248513,I248539,I248187,I248561,I248578,I248595,I248202,I248626,I248643,I248193,I248674,I248196,I248208,I248205,I248763,I248789,I248806,I248755,I248828,I248845,I248862,I248888,I248896,I248922,I248930,I248947,I248734,I248987,I248995,I248728,I248743,I249040,I249057,I249083,I248731,I249105,I249122,I249139,I248746,I249170,I249187,I248737,I249218,I248740,I248752,I248749,I249307,I249333,I249350,I249299,I249372,I249389,I249406,I249432,I249440,I249466,I249474,I249491,I249278,I249531,I249539,I249272,I249287,I249584,I249601,I249627,I249275,I249649,I249666,I249683,I249290,I249714,I249731,I249281,I249762,I249284,I249296,I249293,I249851,I249877,I249894,I249843,I249916,I249933,I249950,I249976,I249984,I250010,I250018,I250035,I249822,I250075,I250083,I249816,I249831,I250128,I250145,I250171,I249819,I250193,I250210,I250227,I249834,I250258,I250275,I249825,I250306,I249828,I249840,I249837,I250395,I250421,I250438,I250387,I250460,I250477,I250494,I250520,I250528,I250554,I250562,I250579,I250366,I250619,I250627,I250360,I250375,I250672,I250689,I250715,I250363,I250737,I250754,I250771,I250378,I250802,I250819,I250369,I250850,I250372,I250384,I250381,I250939,I676347,I250965,I250982,I250931,I251004,I251021,I676344,I676341,I251038,I676329,I251064,I251072,I676353,I251098,I251106,I676338,I251123,I250910,I676332,I251163,I251171,I250904,I250919,I251216,I676335,I251233,I676350,I251259,I250907,I251281,I251298,I251315,I250922,I251346,I251363,I250913,I251394,I250916,I250928,I250925,I251483,I251509,I251526,I251475,I251548,I251565,I251582,I251608,I251616,I251642,I251650,I251667,I251454,I251707,I251715,I251448,I251463,I251760,I251777,I251803,I251451,I251825,I251842,I251859,I251466,I251890,I251907,I251457,I251938,I251460,I251472,I251469,I252027,I289701,I252053,I252070,I252092,I252109,I289704,I289722,I252126,I289710,I252152,I252160,I252186,I252194,I289719,I252211,I289713,I252251,I252259,I252304,I289716,I289698,I252321,I289707,I252347,I252369,I252386,I252403,I252434,I252451,I252482,I252571,I670567,I252597,I252614,I252563,I252636,I252653,I670564,I670561,I252670,I670549,I252696,I252704,I670573,I252730,I252738,I670558,I252755,I252542,I670552,I252795,I252803,I252536,I252551,I252848,I670555,I252865,I670570,I252891,I252539,I252913,I252930,I252947,I252554,I252978,I252995,I252545,I253026,I252548,I252560,I252557,I253115,I253141,I253158,I253107,I253180,I253197,I253214,I253240,I253248,I253274,I253282,I253299,I253086,I253339,I253347,I253080,I253095,I253392,I253409,I253435,I253083,I253457,I253474,I253491,I253098,I253522,I253539,I253089,I253570,I253092,I253104,I253101,I253659,I347824,I253685,I253702,I253651,I253724,I253741,I347845,I347836,I253758,I253784,I253792,I347830,I253818,I253826,I347827,I253843,I253630,I347821,I253883,I253891,I253624,I253639,I253936,I347833,I253953,I347842,I253979,I253627,I254001,I254018,I254035,I253642,I254066,I254083,I347839,I253633,I254114,I253636,I253648,I253645,I254203,I254229,I254246,I254195,I254268,I254285,I254302,I254328,I254336,I254362,I254370,I254387,I254174,I254427,I254435,I254168,I254183,I254480,I254497,I254523,I254171,I254545,I254562,I254579,I254186,I254610,I254627,I254177,I254658,I254180,I254192,I254189,I254747,I659400,I254773,I254790,I254739,I254812,I254829,I659412,I659415,I254846,I659418,I254872,I254880,I659403,I254906,I254914,I659409,I254931,I254718,I659397,I254971,I254979,I254712,I254727,I255024,I659421,I255041,I659406,I255067,I254715,I255089,I255106,I255123,I254730,I255154,I255171,I254721,I255202,I254724,I254736,I254733,I255291,I710900,I255317,I255334,I255283,I255356,I255373,I710876,I710897,I255390,I710894,I255416,I255424,I710873,I255450,I255458,I710885,I255475,I255262,I710888,I255515,I255523,I255256,I255271,I255568,I710891,I710879,I255585,I710882,I255611,I255259,I255633,I255650,I255667,I255274,I255698,I255715,I255265,I255746,I255268,I255280,I255277,I255835,I255861,I255878,I255827,I255900,I255917,I255934,I255960,I255968,I255994,I256002,I256019,I255806,I256059,I256067,I255800,I255815,I256112,I256129,I256155,I255803,I256177,I256194,I256211,I255818,I256242,I256259,I255809,I256290,I255812,I255824,I255821,I256379,I256405,I256422,I256371,I256444,I256461,I256478,I256504,I256512,I256538,I256546,I256563,I256350,I256603,I256611,I256344,I256359,I256656,I256673,I256699,I256347,I256721,I256738,I256755,I256362,I256786,I256803,I256353,I256834,I256356,I256368,I256365,I256923,I565472,I256949,I256966,I256915,I256988,I257005,I565490,I257022,I565484,I257048,I257056,I565478,I257082,I257090,I565487,I257107,I256894,I565475,I257147,I257155,I256888,I256903,I257200,I565493,I257217,I257243,I256891,I257265,I257282,I257299,I256906,I257330,I257347,I565481,I256897,I257378,I256900,I256912,I256909,I257467,I257493,I257510,I257459,I257532,I257549,I257566,I257592,I257600,I257626,I257634,I257651,I257438,I257691,I257699,I257432,I257447,I257744,I257761,I257787,I257435,I257809,I257826,I257843,I257450,I257874,I257891,I257441,I257922,I257444,I257456,I257453,I258011,I258037,I258054,I258003,I258076,I258093,I258110,I258136,I258144,I258170,I258178,I258195,I257982,I258235,I258243,I257976,I257991,I258288,I258305,I258331,I257979,I258353,I258370,I258387,I257994,I258418,I258435,I257985,I258466,I257988,I258000,I257997,I258555,I339154,I258581,I258598,I258547,I258620,I258637,I339151,I339172,I258654,I339175,I258680,I258688,I339160,I258714,I258722,I339163,I258739,I258526,I339166,I258779,I258787,I258520,I258535,I258832,I339157,I258849,I339169,I258875,I258523,I258897,I258914,I258931,I258538,I258962,I258979,I258529,I259010,I258532,I258544,I258541,I259099,I708520,I259125,I259142,I259164,I259181,I708496,I708517,I259198,I708514,I259224,I259232,I708493,I259258,I259266,I708505,I259283,I708508,I259323,I259331,I259376,I708511,I708499,I259393,I708502,I259419,I259441,I259458,I259475,I259506,I259523,I259554,I259643,I259669,I259686,I259708,I259725,I259742,I259768,I259776,I259802,I259810,I259827,I259867,I259875,I259920,I259937,I259963,I259985,I260002,I260019,I260050,I260067,I260098,I260187,I306208,I260213,I260230,I260252,I260269,I306205,I306226,I260286,I306229,I260312,I260320,I306214,I260346,I260354,I306217,I260371,I306220,I260411,I260419,I260464,I306211,I260481,I306223,I260507,I260529,I260546,I260563,I260594,I260611,I260642,I260731,I721610,I260757,I260774,I260796,I260813,I721586,I721607,I260830,I721604,I260856,I260864,I721583,I260890,I260898,I721595,I260915,I721598,I260955,I260963,I261008,I721601,I721589,I261025,I721592,I261051,I261073,I261090,I261107,I261138,I261155,I261186,I261275,I558179,I261301,I261318,I261340,I261357,I558197,I261374,I558191,I261400,I261408,I558185,I261434,I261442,I558194,I261459,I558182,I261499,I261507,I261552,I558200,I261569,I261595,I261617,I261634,I261651,I261682,I261699,I558188,I261730,I261819,I532566,I261845,I261862,I261811,I261884,I261901,I532581,I532569,I261918,I532560,I261944,I261952,I532572,I261978,I261986,I532563,I262003,I261790,I532578,I262043,I262051,I261784,I261799,I262096,I532587,I532575,I262113,I532584,I262139,I261787,I262161,I262178,I262195,I261802,I262226,I262243,I261793,I262274,I261796,I261808,I261805,I262363,I262389,I262406,I262355,I262428,I262445,I262462,I262488,I262496,I262522,I262530,I262547,I262334,I262587,I262595,I262328,I262343,I262640,I262657,I262683,I262331,I262705,I262722,I262739,I262346,I262770,I262787,I262337,I262818,I262340,I262352,I262349,I262907,I311988,I262933,I262950,I262899,I262972,I262989,I311985,I312006,I263006,I312009,I263032,I263040,I311994,I263066,I263074,I311997,I263091,I262878,I312000,I263131,I263139,I262872,I262887,I263184,I311991,I263201,I312003,I263227,I262875,I263249,I263266,I263283,I262890,I263314,I263331,I262881,I263362,I262884,I262896,I262893,I263451,I263477,I263494,I263516,I263533,I263550,I263576,I263584,I263610,I263618,I263635,I263675,I263683,I263728,I263745,I263771,I263793,I263810,I263827,I263858,I263875,I263906,I263995,I264021,I264038,I263987,I264060,I264077,I264094,I264120,I264128,I264154,I264162,I264179,I263966,I264219,I264227,I263960,I263975,I264272,I264289,I264315,I263963,I264337,I264354,I264371,I263978,I264402,I264419,I263969,I264450,I263972,I263984,I263981,I264539,I264565,I264582,I264531,I264604,I264621,I264638,I264664,I264672,I264698,I264706,I264723,I264510,I264763,I264771,I264504,I264519,I264816,I264833,I264859,I264507,I264881,I264898,I264915,I264522,I264946,I264963,I264513,I264994,I264516,I264528,I264525,I265083,I678659,I265109,I265126,I265148,I265165,I678656,I678653,I265182,I678641,I265208,I265216,I678665,I265242,I265250,I678650,I265267,I678644,I265307,I265315,I265360,I678647,I265377,I678662,I265403,I265425,I265442,I265459,I265490,I265507,I265538,I265627,I281966,I265653,I265670,I265619,I265692,I265709,I281969,I281987,I265726,I281975,I265752,I265760,I265786,I265794,I281984,I265811,I265598,I281978,I265851,I265859,I265592,I265607,I265904,I281981,I281963,I265921,I281972,I265947,I265595,I265969,I265986,I266003,I265610,I266034,I266051,I265601,I266082,I265604,I265616,I265613,I266171,I321236,I266197,I266214,I266236,I266253,I321233,I321254,I266270,I321257,I266296,I266304,I321242,I266330,I266338,I321245,I266355,I321248,I266395,I266403,I266448,I321239,I266465,I321251,I266491,I266513,I266530,I266547,I266578,I266595,I266626,I266715,I353026,I266741,I266758,I266780,I266797,I353047,I353038,I266814,I266840,I266848,I353032,I266874,I266882,I353029,I266899,I353023,I266939,I266947,I266992,I353035,I267009,I353044,I267035,I267057,I267074,I267091,I267122,I267139,I353041,I267170,I267259,I458690,I267285,I267302,I267251,I267324,I267341,I458684,I458681,I267358,I458696,I267384,I267392,I267418,I267426,I458678,I267443,I267230,I267483,I267491,I267224,I267239,I267536,I458693,I458687,I267553,I267579,I267227,I267601,I267618,I267635,I267242,I267666,I267683,I458699,I267233,I267714,I267236,I267248,I267245,I267803,I576304,I267829,I267846,I267795,I267868,I267885,I576316,I267902,I576307,I267928,I267936,I576325,I267962,I267970,I576301,I267987,I267774,I576319,I268027,I268035,I267768,I267783,I268080,I576313,I576310,I268097,I576322,I268123,I267771,I268145,I268162,I268179,I267786,I268210,I268227,I267777,I268258,I267780,I267792,I267789,I268347,I268373,I268390,I268339,I268412,I268429,I268446,I268472,I268480,I268506,I268514,I268531,I268318,I268571,I268579,I268312,I268327,I268624,I268641,I268667,I268315,I268689,I268706,I268723,I268330,I268754,I268771,I268321,I268802,I268324,I268336,I268333,I268891,I520938,I268917,I268934,I268883,I268956,I268973,I520953,I520941,I268990,I520932,I269016,I269024,I520944,I269050,I269058,I520935,I269075,I268862,I520950,I269115,I269123,I268856,I268871,I269168,I520959,I520947,I269185,I520956,I269211,I268859,I269233,I269250,I269267,I268874,I269298,I269315,I268865,I269346,I268868,I268880,I268877,I269435,I269461,I269478,I269427,I269500,I269517,I269534,I269560,I269568,I269594,I269602,I269619,I269406,I269659,I269667,I269400,I269415,I269712,I269729,I269755,I269403,I269777,I269794,I269811,I269418,I269842,I269859,I269409,I269890,I269412,I269424,I269421,I269979,I521584,I270005,I270022,I270044,I270061,I521599,I521587,I270078,I521578,I270104,I270112,I521590,I270138,I270146,I521581,I270163,I521596,I270203,I270211,I270256,I521605,I521593,I270273,I521602,I270299,I270321,I270338,I270355,I270386,I270403,I270434,I270523,I428651,I270549,I270566,I270515,I270588,I270605,I428645,I428642,I270622,I428657,I270648,I270656,I270682,I270690,I428639,I270707,I270494,I270747,I270755,I270488,I270503,I270800,I428654,I428648,I270817,I270843,I270491,I270865,I270882,I270899,I270506,I270930,I270947,I428660,I270497,I270978,I270500,I270512,I270509,I271067,I437610,I271093,I271110,I271059,I271132,I271149,I437604,I437601,I271166,I437616,I271192,I271200,I271226,I271234,I437598,I271251,I271038,I271291,I271299,I271032,I271047,I271344,I437613,I437607,I271361,I271387,I271035,I271409,I271426,I271443,I271050,I271474,I271491,I437619,I271041,I271522,I271044,I271056,I271053,I271611,I362274,I271637,I271654,I271676,I271693,I362295,I362286,I271710,I271736,I271744,I362280,I271770,I271778,I362277,I271795,I362271,I271835,I271843,I271888,I362283,I271905,I362292,I271931,I271953,I271970,I271987,I272018,I272035,I362289,I272066,I272155,I272181,I272198,I272147,I272220,I272237,I272254,I272280,I272288,I272314,I272322,I272339,I272126,I272379,I272387,I272120,I272135,I272432,I272449,I272475,I272123,I272497,I272514,I272531,I272138,I272562,I272579,I272129,I272610,I272132,I272144,I272141,I272699,I272725,I272742,I272691,I272764,I272781,I272798,I272824,I272832,I272858,I272866,I272883,I272670,I272923,I272931,I272664,I272679,I272976,I272993,I273019,I272667,I273041,I273058,I273075,I272682,I273106,I273123,I272673,I273154,I272676,I272688,I272685,I273243,I609828,I273269,I273286,I273235,I273308,I273325,I609840,I273342,I609831,I273368,I273376,I609849,I273402,I273410,I609825,I273427,I273214,I609843,I273467,I273475,I273208,I273223,I273520,I609837,I609834,I273537,I609846,I273563,I273211,I273585,I273602,I273619,I273226,I273650,I273667,I273217,I273698,I273220,I273232,I273229,I273787,I344356,I273813,I273830,I273779,I273852,I273869,I344353,I344374,I273886,I344377,I273912,I273920,I344362,I273946,I273954,I344365,I273971,I273758,I344368,I274011,I274019,I273752,I273767,I274064,I344359,I274081,I344371,I274107,I273755,I274129,I274146,I274163,I273770,I274194,I274211,I273761,I274242,I273764,I273776,I273773,I274331,I274357,I274374,I274323,I274396,I274413,I274430,I274456,I274464,I274490,I274498,I274515,I274302,I274555,I274563,I274296,I274311,I274608,I274625,I274651,I274299,I274673,I274690,I274707,I274314,I274738,I274755,I274305,I274786,I274308,I274320,I274317,I274875,I590176,I274901,I274918,I274867,I274940,I274957,I590188,I274974,I590179,I275000,I275008,I590197,I275034,I275042,I590173,I275059,I274846,I590191,I275099,I275107,I274840,I274855,I275152,I590185,I590182,I275169,I590194,I275195,I274843,I275217,I275234,I275251,I274858,I275282,I275299,I274849,I275330,I274852,I274864,I274861,I275419,I275445,I275462,I275484,I275501,I275518,I275544,I275552,I275578,I275586,I275603,I275643,I275651,I275696,I275713,I275739,I275761,I275778,I275795,I275826,I275843,I275874,I275963,I557057,I275989,I276006,I275955,I276028,I276045,I557075,I276062,I557069,I276088,I276096,I557063,I276122,I276130,I557072,I276147,I275934,I557060,I276187,I276195,I275928,I275943,I276240,I557078,I276257,I276283,I275931,I276305,I276322,I276339,I275946,I276370,I276387,I557066,I275937,I276418,I275940,I275952,I275949,I276507,I363430,I276533,I276550,I276499,I276572,I276589,I363451,I363442,I276606,I276632,I276640,I363436,I276666,I276674,I363433,I276691,I276478,I363427,I276731,I276739,I276472,I276487,I276784,I363439,I276801,I363448,I276827,I276475,I276849,I276866,I276883,I276490,I276914,I276931,I363445,I276481,I276962,I276484,I276496,I276493,I277051,I648520,I277077,I277094,I277116,I277133,I648532,I648535,I277150,I648538,I277176,I277184,I648523,I277210,I277218,I648529,I277235,I648517,I277275,I277283,I277328,I648541,I277345,I648526,I277371,I277393,I277410,I277427,I277458,I277475,I277506,I277595,I391174,I277621,I277638,I277587,I277660,I277677,I391195,I391186,I277694,I277720,I277728,I391180,I277754,I277762,I391177,I277779,I277566,I391171,I277819,I277827,I277560,I277575,I277872,I391183,I277889,I391192,I277915,I277563,I277937,I277954,I277971,I277578,I278002,I278019,I391189,I277569,I278050,I277572,I277584,I277581,I278139,I278165,I278182,I278131,I278204,I278221,I278238,I278264,I278272,I278298,I278306,I278323,I278110,I278363,I278371,I278104,I278119,I278416,I278433,I278459,I278107,I278481,I278498,I278515,I278122,I278546,I278563,I278113,I278594,I278116,I278128,I278125,I278683,I278709,I278726,I278675,I278748,I278765,I278782,I278808,I278816,I278842,I278850,I278867,I278654,I278907,I278915,I278648,I278663,I278960,I278977,I279003,I278651,I279025,I279042,I279059,I278666,I279090,I279107,I278657,I279138,I278660,I278672,I278669,I279227,I329906,I279253,I279270,I279219,I279292,I279309,I329903,I329924,I279326,I329927,I279352,I279360,I329912,I279386,I279394,I329915,I279411,I279198,I329918,I279451,I279459,I279192,I279207,I279504,I329909,I279521,I329921,I279547,I279195,I279569,I279586,I279603,I279210,I279634,I279651,I279201,I279682,I279204,I279216,I279213,I279771,I305052,I279797,I279814,I279836,I279853,I305049,I305070,I279870,I305073,I279896,I279904,I305058,I279930,I279938,I305061,I279955,I305064,I279995,I280003,I280048,I305055,I280065,I305067,I280091,I280113,I280130,I280147,I280178,I280195,I280226,I280315,I526106,I280341,I280358,I280307,I280380,I280397,I526121,I526109,I280414,I526100,I280440,I280448,I526112,I280474,I280482,I526103,I280499,I280286,I526118,I280539,I280547,I280280,I280295,I280592,I526127,I526115,I280609,I526124,I280635,I280283,I280657,I280674,I280691,I280298,I280722,I280739,I280289,I280770,I280292,I280304,I280301,I280859,I608094,I280885,I280902,I280924,I280941,I608106,I280958,I608097,I280984,I280992,I608115,I281018,I281026,I608091,I281043,I608109,I281083,I281091,I281136,I608103,I608100,I281153,I608112,I281179,I281201,I281218,I281235,I281266,I281283,I281314,I281400,I281426,I281443,I281392,I281474,I281482,I281499,I281516,I281533,I281550,I281567,I281584,I281389,I281615,I281632,I281649,I281374,I281386,I281694,I281711,I281380,I281742,I281759,I281368,I281790,I281807,I281824,I281850,I281858,I281377,I281889,I281906,I281383,I281937,I281371,I281995,I282021,I282038,I282069,I282077,I282094,I282111,I282128,I282145,I282162,I282179,I282210,I282227,I282244,I282289,I282306,I282337,I282354,I282385,I282402,I282419,I282445,I282453,I282484,I282501,I282532,I282590,I450255,I282616,I282633,I450252,I282664,I282672,I282689,I282706,I450249,I282723,I450264,I282740,I282757,I282774,I282805,I450258,I282822,I450246,I282839,I282884,I282901,I282932,I450267,I282949,I282980,I282997,I450261,I283014,I283040,I283048,I283079,I283096,I283127,I283185,I283211,I283228,I283177,I283259,I283267,I283284,I283301,I283318,I283335,I283352,I283369,I283174,I283400,I283417,I283434,I283159,I283171,I283479,I283496,I283165,I283527,I283544,I283153,I283575,I283592,I283609,I283635,I283643,I283162,I283674,I283691,I283168,I283722,I283156,I283780,I460268,I283806,I283823,I460265,I283854,I283862,I283879,I283896,I460262,I283913,I460277,I283930,I283947,I283964,I283995,I460271,I284012,I460259,I284029,I284074,I284091,I284122,I460280,I284139,I284170,I284187,I460274,I284204,I284230,I284238,I284269,I284286,I284317,I284375,I357656,I284401,I284418,I284367,I357650,I284449,I284457,I357647,I284474,I284491,I357659,I284508,I357662,I284525,I284542,I284559,I284364,I284590,I357671,I284607,I357665,I284624,I284349,I284361,I284669,I284686,I284355,I284717,I357653,I284734,I284343,I284765,I357668,I284782,I284799,I284825,I284833,I284352,I284864,I284881,I284358,I284912,I284346,I284970,I656677,I284996,I285013,I284962,I656692,I285044,I285052,I656701,I285069,I285086,I656680,I285103,I656686,I285120,I285137,I285154,I284959,I285185,I656698,I285202,I656695,I285219,I284944,I284956,I285264,I285281,I284950,I285312,I285329,I284938,I285360,I656689,I285377,I656683,I285394,I285420,I285428,I284947,I285459,I285476,I284953,I285507,I284941,I285565,I730508,I285591,I285608,I285557,I730514,I285639,I285647,I730529,I285664,I285681,I730520,I285698,I730517,I285715,I285732,I285749,I285554,I285780,I285797,I730532,I285814,I285539,I285551,I285859,I285876,I285545,I285907,I730526,I285924,I285533,I285955,I730511,I285972,I730523,I285989,I730535,I286015,I286023,I285542,I286054,I286071,I285548,I286102,I285536,I286160,I380776,I286186,I286203,I380770,I286234,I286242,I380767,I286259,I286276,I380779,I286293,I380782,I286310,I286327,I286344,I286375,I380791,I286392,I380785,I286409,I286454,I286471,I286502,I380773,I286519,I286550,I380788,I286567,I286584,I286610,I286618,I286649,I286666,I286697,I286755,I336264,I286781,I286798,I286747,I336276,I286829,I286837,I336261,I286854,I286871,I336279,I286888,I336270,I286905,I286922,I286939,I286744,I286970,I336282,I286987,I336285,I287004,I286729,I286741,I287049,I287066,I286735,I287097,I287114,I286723,I287145,I336273,I287162,I336267,I287179,I287205,I287213,I286732,I287244,I287261,I286738,I287292,I286726,I287350,I287376,I287393,I287342,I287424,I287432,I287449,I287466,I287483,I287500,I287517,I287534,I287339,I287565,I287582,I287599,I287324,I287336,I287644,I287661,I287330,I287692,I287709,I287318,I287740,I287757,I287774,I287800,I287808,I287327,I287839,I287856,I287333,I287887,I287321,I287945,I473443,I287971,I287988,I473440,I288019,I288027,I288044,I288061,I473437,I288078,I473452,I288095,I288112,I288129,I288160,I473446,I288177,I473434,I288194,I288239,I288256,I288287,I473455,I288304,I288335,I288352,I473449,I288369,I288395,I288403,I288434,I288451,I288482,I288540,I288566,I288583,I288532,I288614,I288622,I288639,I288656,I288673,I288690,I288707,I288724,I288529,I288755,I288772,I288789,I288514,I288526,I288834,I288851,I288520,I288882,I288899,I288508,I288930,I288947,I288964,I288990,I288998,I288517,I289029,I289046,I288523,I289077,I288511,I289135,I664837,I289161,I289178,I289127,I664852,I289209,I289217,I664861,I289234,I289251,I664840,I289268,I664846,I289285,I289302,I289319,I289124,I289350,I664858,I289367,I664855,I289384,I289109,I289121,I289429,I289446,I289115,I289477,I289494,I289103,I289525,I664849,I289542,I664843,I289559,I289585,I289593,I289112,I289624,I289641,I289118,I289672,I289106,I289730,I289756,I289773,I289804,I289812,I289829,I289846,I289863,I289880,I289897,I289914,I289945,I289962,I289979,I290024,I290041,I290072,I290089,I290120,I290137,I290154,I290180,I290188,I290219,I290236,I290267,I290325,I418346,I290351,I290368,I418340,I290399,I290407,I418337,I290424,I290441,I418349,I290458,I418352,I290475,I290492,I290509,I290540,I418361,I290557,I418355,I290574,I290619,I290636,I290667,I418343,I290684,I290715,I418358,I290732,I290749,I290775,I290783,I290814,I290831,I290862,I290920,I668246,I290946,I290963,I290912,I668252,I290994,I291002,I668240,I291019,I291036,I668243,I291053,I668249,I291070,I291087,I291104,I290909,I291135,I291152,I668258,I291169,I290894,I290906,I291214,I291231,I290900,I291262,I668237,I291279,I290888,I291310,I668261,I291327,I291344,I668255,I291370,I291378,I290897,I291409,I291426,I290903,I291457,I290891,I291515,I491877,I291541,I291558,I491865,I291589,I291597,I491862,I291614,I291631,I491874,I291648,I491871,I291665,I291682,I291699,I291730,I491880,I291747,I491883,I291764,I291809,I291826,I291857,I491886,I291874,I291905,I491889,I291922,I491868,I291939,I291965,I291973,I292004,I292021,I292052,I292110,I292136,I292153,I292102,I292184,I292192,I292209,I292226,I292243,I292260,I292277,I292294,I292099,I292325,I292342,I292359,I292084,I292096,I292404,I292421,I292090,I292452,I292469,I292078,I292500,I292517,I292534,I292560,I292568,I292087,I292599,I292616,I292093,I292647,I292081,I292705,I292731,I292748,I292697,I292779,I292787,I292804,I292821,I292838,I292855,I292872,I292889,I292694,I292920,I292937,I292954,I292679,I292691,I292999,I293016,I292685,I293047,I293064,I292673,I293095,I293112,I293129,I293155,I293163,I292682,I293194,I293211,I292688,I293242,I292676,I293300,I293326,I293343,I293292,I293374,I293382,I293399,I293416,I293433,I293450,I293467,I293484,I293289,I293515,I293532,I293549,I293274,I293286,I293594,I293611,I293280,I293642,I293659,I293268,I293690,I293707,I293724,I293750,I293758,I293277,I293789,I293806,I293283,I293837,I293271,I293895,I607531,I293921,I293938,I607513,I293969,I293977,I607519,I293994,I294011,I607534,I294028,I607525,I294045,I294062,I294079,I294110,I607537,I294127,I607516,I294144,I294189,I294206,I294237,I607522,I294254,I294285,I607528,I294302,I294319,I294345,I294353,I294384,I294401,I294432,I294490,I612155,I294516,I294533,I612137,I294564,I294572,I612143,I294589,I294606,I612158,I294623,I612149,I294640,I294657,I294674,I294705,I612161,I294722,I612140,I294739,I294784,I294801,I294832,I612146,I294849,I294880,I612152,I294897,I294914,I294940,I294948,I294979,I294996,I295027,I295085,I657221,I295111,I295128,I657236,I295159,I295167,I657245,I295184,I295201,I657224,I295218,I657230,I295235,I295252,I295269,I295300,I657242,I295317,I657239,I295334,I295379,I295396,I295427,I295444,I295475,I657233,I295492,I657227,I295509,I295535,I295543,I295574,I295591,I295622,I295680,I536451,I295706,I295723,I295672,I536439,I295754,I295762,I536436,I295779,I295796,I536448,I295813,I536445,I295830,I295847,I295864,I295669,I295895,I536454,I295912,I536457,I295929,I295654,I295666,I295974,I295991,I295660,I296022,I536460,I296039,I295648,I296070,I536463,I296087,I536442,I296104,I296130,I296138,I295657,I296169,I296186,I295663,I296217,I295651,I296275,I296301,I296318,I296349,I296357,I296374,I296391,I296408,I296425,I296442,I296459,I296490,I296507,I296524,I296569,I296586,I296617,I296634,I296665,I296682,I296699,I296725,I296733,I296764,I296781,I296812,I296870,I718013,I296896,I296913,I296862,I718019,I296944,I296952,I718034,I296969,I296986,I718025,I297003,I718022,I297020,I297037,I297054,I296859,I297085,I297102,I718037,I297119,I296844,I296856,I297164,I297181,I296850,I297212,I718031,I297229,I296838,I297260,I718016,I297277,I718028,I297294,I718040,I297320,I297328,I296847,I297359,I297376,I296853,I297407,I296841,I297465,I435499,I297491,I297508,I297457,I435496,I297539,I297547,I297564,I297581,I435493,I297598,I435508,I297615,I297632,I297649,I297454,I297680,I435502,I297697,I435490,I297714,I297439,I297451,I297759,I297776,I297445,I297807,I435511,I297824,I297433,I297855,I297872,I435505,I297889,I297915,I297923,I297442,I297954,I297971,I297448,I298002,I297436,I298060,I298086,I298103,I298134,I298142,I298159,I298176,I298193,I298210,I298227,I298244,I298275,I298292,I298309,I298354,I298371,I298402,I298419,I298450,I298467,I298484,I298510,I298518,I298549,I298566,I298597,I298655,I623137,I298681,I298698,I298647,I623119,I298729,I298737,I623125,I298754,I298771,I623140,I298788,I623131,I298805,I298822,I298839,I298644,I298870,I623143,I298887,I623122,I298904,I298629,I298641,I298949,I298966,I298635,I298997,I623128,I299014,I298623,I299045,I623134,I299062,I299079,I299105,I299113,I298632,I299144,I299161,I298638,I299192,I298626,I299250,I462376,I299276,I299293,I462373,I299324,I299332,I299349,I299366,I462370,I299383,I462385,I299400,I299417,I299434,I299465,I462379,I299482,I462367,I299499,I299544,I299561,I299592,I462388,I299609,I299640,I299657,I462382,I299674,I299700,I299708,I299739,I299756,I299787,I299845,I444985,I299871,I299888,I299837,I444982,I299919,I299927,I299944,I299961,I444979,I299978,I444994,I299995,I300012,I300029,I299834,I300060,I444988,I300077,I444976,I300094,I299819,I299831,I300139,I300156,I299825,I300187,I444997,I300204,I299813,I300235,I300252,I444991,I300269,I300295,I300303,I299822,I300334,I300351,I299828,I300382,I299816,I300440,I300466,I300483,I300514,I300522,I300539,I300556,I300573,I300590,I300607,I300624,I300655,I300672,I300689,I300734,I300751,I300782,I300799,I300830,I300847,I300864,I300890,I300898,I300929,I300946,I300977,I301035,I301061,I301069,I301095,I301103,I301120,I301137,I301154,I301171,I301021,I301202,I301219,I301236,I301253,I301018,I301009,I301298,I301012,I301006,I301343,I301360,I301377,I301015,I301408,I301425,I301442,I301468,I301476,I301003,I301027,I301521,I301538,I301555,I301024,I301613,I428118,I301639,I301647,I301673,I301681,I428115,I301698,I428130,I301715,I301732,I428124,I301749,I301780,I301797,I301814,I428121,I301831,I428112,I301876,I301921,I428133,I301938,I301955,I301986,I302003,I302020,I428127,I302046,I302054,I302099,I302116,I302133,I302191,I376721,I302217,I302225,I376733,I302251,I302259,I376724,I302276,I376727,I302293,I302310,I376730,I302327,I302358,I302375,I302392,I302409,I376736,I302454,I302499,I376742,I302516,I302533,I302564,I302581,I376739,I302598,I376745,I302624,I302632,I302677,I302694,I302711,I302769,I302795,I302803,I302829,I302837,I302854,I302871,I302888,I302905,I302755,I302936,I302953,I302970,I302987,I302752,I302743,I303032,I302746,I302740,I303077,I303094,I303111,I302749,I303142,I303159,I303176,I303202,I303210,I302737,I302761,I303255,I303272,I303289,I302758,I303347,I303373,I303381,I303407,I303415,I303432,I303449,I303466,I303483,I303333,I303514,I303531,I303548,I303565,I303330,I303321,I303610,I303324,I303318,I303655,I303672,I303689,I303327,I303720,I303737,I303754,I303780,I303788,I303315,I303339,I303833,I303850,I303867,I303336,I303925,I614449,I303951,I303959,I614455,I303985,I303993,I304010,I614452,I304027,I304044,I614470,I304061,I303911,I304092,I304109,I304126,I614473,I304143,I303908,I303899,I304188,I303902,I303896,I304233,I614458,I304250,I304267,I303905,I304298,I614464,I304315,I614461,I304332,I614467,I304358,I304366,I303893,I303917,I304411,I304428,I304445,I303914,I304503,I304529,I304537,I304563,I304571,I304588,I304605,I304622,I304639,I304489,I304670,I304687,I304704,I304721,I304486,I304477,I304766,I304480,I304474,I304811,I304828,I304845,I304483,I304876,I304893,I304910,I304936,I304944,I304471,I304495,I304989,I305006,I305023,I304492,I305081,I499620,I305107,I305115,I499617,I305141,I305149,I499614,I305166,I499641,I305183,I305200,I499629,I305217,I305248,I305265,I305282,I499635,I305299,I499626,I305344,I305389,I499623,I305406,I305423,I305454,I499638,I305471,I499632,I305488,I305514,I305522,I305567,I305584,I305601,I305659,I547541,I305685,I305693,I547532,I305719,I305727,I547526,I305744,I547538,I305761,I305778,I547529,I305795,I305826,I305843,I305860,I547535,I305877,I547520,I305922,I305967,I305984,I306001,I306032,I547523,I306049,I306066,I306092,I306100,I306145,I306162,I306179,I306237,I515124,I306263,I306271,I515121,I306297,I306305,I515118,I306322,I515145,I306339,I306356,I515133,I306373,I306404,I306421,I306438,I515139,I306455,I515130,I306500,I306545,I515127,I306562,I306579,I306610,I515142,I306627,I515136,I306644,I306670,I306678,I306723,I306740,I306757,I306815,I538380,I306841,I306849,I538377,I306875,I306883,I538374,I306900,I538401,I306917,I306934,I538389,I306951,I306801,I306982,I306999,I307016,I538395,I307033,I538386,I306798,I306789,I307078,I306792,I306786,I307123,I538383,I307140,I307157,I306795,I307188,I538398,I307205,I538392,I307222,I307248,I307256,I306783,I306807,I307301,I307318,I307335,I306804,I307393,I307419,I307427,I307453,I307461,I307478,I307495,I307512,I307529,I307379,I307560,I307577,I307594,I307611,I307376,I307367,I307656,I307370,I307364,I307701,I307718,I307735,I307373,I307766,I307783,I307800,I307826,I307834,I307361,I307385,I307879,I307896,I307913,I307382,I307971,I307997,I308005,I308031,I308039,I308056,I308073,I308090,I308107,I308138,I308155,I308172,I308189,I308234,I308279,I308296,I308313,I308344,I308361,I308378,I308404,I308412,I308457,I308474,I308491,I308549,I636991,I308575,I308583,I636997,I308609,I308617,I308634,I636994,I308651,I308668,I637012,I308685,I308535,I308716,I308733,I308750,I637015,I308767,I308532,I308523,I308812,I308526,I308520,I308857,I637000,I308874,I308891,I308529,I308922,I637006,I308939,I637003,I308956,I637009,I308982,I308990,I308517,I308541,I309035,I309052,I309069,I308538,I309127,I309153,I309161,I309187,I309195,I309212,I309229,I309246,I309263,I309294,I309311,I309328,I309345,I309390,I309435,I309452,I309469,I309500,I309517,I309534,I309560,I309568,I309613,I309630,I309647,I309705,I465535,I309731,I309739,I309765,I309773,I465532,I309790,I465547,I309807,I309824,I465541,I309841,I309872,I309889,I309906,I465538,I309923,I465529,I309968,I310013,I465550,I310030,I310047,I310078,I310095,I310112,I465544,I310138,I310146,I310191,I310208,I310225,I310283,I310309,I310317,I310343,I310351,I310368,I310385,I310402,I310419,I310269,I310450,I310467,I310484,I310501,I310266,I310257,I310546,I310260,I310254,I310591,I310608,I310625,I310263,I310656,I310673,I310690,I310716,I310724,I310251,I310275,I310769,I310786,I310803,I310272,I310861,I680965,I310887,I310895,I680977,I310921,I310929,I680968,I310946,I680956,I310963,I310980,I680953,I310997,I310847,I311028,I311045,I311062,I680959,I311079,I310844,I310835,I311124,I310838,I310832,I311169,I680974,I311186,I311203,I310841,I311234,I680962,I311251,I311268,I680971,I311294,I311302,I310829,I310853,I311347,I311364,I311381,I310850,I311439,I425273,I311465,I311473,I425285,I311499,I311507,I425276,I311524,I425279,I311541,I311558,I425282,I311575,I311425,I311606,I311623,I311640,I311657,I425288,I311422,I311413,I311702,I311416,I311410,I311747,I425294,I311764,I311781,I311419,I311812,I311829,I425291,I311846,I425297,I311872,I311880,I311407,I311431,I311925,I311942,I311959,I311428,I312017,I312043,I312051,I312077,I312085,I312102,I312119,I312136,I312153,I312184,I312201,I312218,I312235,I312280,I312325,I312342,I312359,I312390,I312407,I312424,I312450,I312458,I312503,I312520,I312537,I312595,I312621,I312629,I312655,I312663,I312680,I312697,I312714,I312731,I312762,I312779,I312796,I312813,I312858,I312903,I312920,I312937,I312968,I312985,I313002,I313028,I313036,I313081,I313098,I313115,I313173,I313199,I313207,I313233,I313241,I313258,I313275,I313292,I313309,I313159,I313340,I313357,I313374,I313391,I313156,I313147,I313436,I313150,I313144,I313481,I313498,I313515,I313153,I313546,I313563,I313580,I313606,I313614,I313141,I313165,I313659,I313676,I313693,I313162,I313751,I647447,I313777,I313785,I647441,I313811,I313819,I647450,I313836,I647429,I313853,I313870,I647438,I313887,I313918,I313935,I313952,I647453,I313969,I647432,I314014,I314059,I647435,I314076,I314093,I314124,I647444,I314141,I314158,I314184,I314192,I314237,I314254,I314271,I314329,I314355,I314363,I314389,I314397,I314414,I314431,I314448,I314465,I314315,I314496,I314513,I314530,I314547,I314312,I314303,I314592,I314306,I314300,I314637,I314654,I314671,I314309,I314702,I314719,I314736,I314762,I314770,I314297,I314321,I314815,I314832,I314849,I314318,I314907,I500912,I314933,I314941,I500909,I314967,I314975,I500906,I314992,I500933,I315009,I315026,I500921,I315043,I315074,I315091,I315108,I500927,I315125,I500918,I315170,I315215,I500915,I315232,I315249,I315280,I500930,I315297,I500924,I315314,I315340,I315348,I315393,I315410,I315427,I315485,I446563,I315511,I315519,I315545,I315553,I446560,I315570,I446575,I315587,I315604,I446569,I315621,I315471,I315652,I315669,I315686,I446566,I315703,I446557,I315468,I315459,I315748,I315462,I315456,I315793,I446578,I315810,I315827,I315465,I315858,I315875,I315892,I446572,I315918,I315926,I315453,I315477,I315971,I315988,I316005,I315474,I316063,I316089,I316097,I316123,I316131,I316148,I316165,I316182,I316199,I316230,I316247,I316264,I316281,I316326,I316371,I316388,I316405,I316436,I316453,I316470,I316496,I316504,I316549,I316566,I316583,I316641,I316667,I316675,I316701,I316709,I316726,I316743,I316760,I316777,I316627,I316808,I316825,I316842,I316859,I316624,I316615,I316904,I316618,I316612,I316949,I316966,I316983,I316621,I317014,I317031,I317048,I317074,I317082,I316609,I316633,I317127,I317144,I317161,I316630,I317219,I317245,I317253,I317279,I317287,I317304,I317321,I317338,I317355,I317386,I317403,I317420,I317437,I317482,I317527,I317544,I317561,I317592,I317609,I317626,I317652,I317660,I317705,I317722,I317739,I317797,I573411,I317823,I317831,I573417,I317857,I317865,I317882,I573414,I317899,I317916,I573432,I317933,I317783,I317964,I317981,I317998,I573435,I318015,I317780,I317771,I318060,I317774,I317768,I318105,I573420,I318122,I318139,I317777,I318170,I573426,I318187,I573423,I318204,I573429,I318230,I318238,I317765,I317789,I318283,I318300,I318317,I317786,I318375,I555956,I318401,I318409,I555947,I318435,I318443,I555941,I318460,I555953,I318477,I318494,I555944,I318511,I318361,I318542,I318559,I318576,I555950,I318593,I555935,I318358,I318349,I318638,I318352,I318346,I318683,I318700,I318717,I318355,I318748,I555938,I318765,I318782,I318808,I318816,I318343,I318367,I318861,I318878,I318895,I318364,I318953,I649623,I318979,I318987,I649617,I319013,I319021,I649626,I319038,I649605,I319055,I319072,I649614,I319089,I318939,I319120,I319137,I319154,I649629,I319171,I649608,I318936,I318927,I319216,I318930,I318924,I319261,I649611,I319278,I319295,I318933,I319326,I649620,I319343,I319360,I319386,I319394,I318921,I318945,I319439,I319456,I319473,I318942,I319531,I552590,I319557,I319565,I552581,I319591,I319599,I552575,I319616,I552587,I319633,I319650,I552578,I319667,I319517,I319698,I319715,I319732,I552584,I319749,I552569,I319514,I319505,I319794,I319508,I319502,I319839,I319856,I319873,I319511,I319904,I552572,I319921,I319938,I319964,I319972,I319499,I319523,I320017,I320034,I320051,I319520,I320109,I421227,I320135,I320143,I421239,I320169,I320177,I421230,I320194,I421233,I320211,I320228,I421236,I320245,I320095,I320276,I320293,I320310,I320327,I421242,I320092,I320083,I320372,I320086,I320080,I320417,I421248,I320434,I320451,I320089,I320482,I320499,I421245,I320516,I421251,I320542,I320550,I320077,I320101,I320595,I320612,I320629,I320098,I320687,I320713,I320721,I320747,I320755,I320772,I320789,I320806,I320823,I320854,I320871,I320888,I320905,I320950,I320995,I321012,I321029,I321060,I321077,I321094,I321120,I321128,I321173,I321190,I321207,I321265,I539687,I321291,I321299,I539678,I321325,I321333,I539672,I321350,I539684,I321367,I321384,I539675,I321401,I321432,I321449,I321466,I539681,I321483,I539666,I321528,I321573,I321590,I321607,I321638,I539669,I321655,I321672,I321698,I321706,I321751,I321768,I321785,I321843,I496390,I321869,I321877,I496387,I321903,I321911,I496384,I321928,I496411,I321945,I321962,I496399,I321979,I322010,I322027,I322044,I496405,I322061,I496396,I322106,I322151,I496393,I322168,I322185,I322216,I496408,I322233,I496402,I322250,I322276,I322284,I322329,I322346,I322363,I322421,I619651,I322447,I322455,I619657,I322481,I322489,I322506,I619654,I322523,I322540,I619672,I322557,I322407,I322588,I322605,I322622,I619675,I322639,I322404,I322395,I322684,I322398,I322392,I322729,I619660,I322746,I322763,I322401,I322794,I619666,I322811,I619663,I322828,I619669,I322854,I322862,I322389,I322413,I322907,I322924,I322941,I322410,I322999,I323025,I323033,I323059,I323067,I323084,I323101,I323118,I323135,I322985,I323166,I323183,I323200,I323217,I322982,I322973,I323262,I322976,I322970,I323307,I323324,I323341,I322979,I323372,I323389,I323406,I323432,I323440,I322967,I322991,I323485,I323502,I323519,I322988,I323577,I323603,I323611,I323637,I323645,I323662,I323679,I323696,I323713,I323744,I323761,I323778,I323795,I323840,I323885,I323902,I323919,I323950,I323967,I323984,I324010,I324018,I324063,I324080,I324097,I324155,I427591,I324181,I324189,I324215,I324223,I427588,I324240,I427603,I324257,I324274,I427597,I324291,I324322,I324339,I324356,I427594,I324373,I427585,I324418,I324463,I427606,I324480,I324497,I324528,I324545,I324562,I427600,I324588,I324596,I324641,I324658,I324675,I324733,I375565,I324759,I324767,I375577,I324793,I324801,I375568,I324818,I375571,I324835,I324852,I375574,I324869,I324719,I324900,I324917,I324934,I324951,I375580,I324716,I324707,I324996,I324710,I324704,I325041,I375586,I325058,I325075,I324713,I325106,I325123,I375583,I325140,I375589,I325166,I325174,I324701,I324725,I325219,I325236,I325253,I324722,I325311,I325337,I325345,I325371,I325379,I325396,I325413,I325430,I325447,I325297,I325478,I325495,I325512,I325529,I325294,I325285,I325574,I325288,I325282,I325619,I325636,I325653,I325291,I325684,I325701,I325718,I325744,I325752,I325279,I325303,I325797,I325814,I325831,I325300,I325889,I541931,I325915,I325923,I541922,I325949,I325957,I541916,I325974,I541928,I325991,I326008,I541919,I326025,I325875,I326056,I326073,I326090,I541925,I326107,I541910,I325872,I325863,I326152,I325866,I325860,I326197,I326214,I326231,I325869,I326262,I541913,I326279,I326296,I326322,I326330,I325857,I325881,I326375,I326392,I326409,I325878,I326467,I326493,I326501,I326527,I326535,I326552,I326569,I326586,I326603,I326453,I326634,I326651,I326668,I326685,I326450,I326441,I326730,I326444,I326438,I326775,I326792,I326809,I326447,I326840,I326857,I326874,I326900,I326908,I326435,I326459,I326953,I326970,I326987,I326456,I327045,I327071,I327079,I327105,I327113,I327130,I327147,I327164,I327181,I327031,I327212,I327229,I327246,I327263,I327028,I327019,I327308,I327022,I327016,I327353,I327370,I327387,I327025,I327418,I327435,I327452,I327478,I327486,I327013,I327037,I327531,I327548,I327565,I327034,I327623,I327649,I327657,I327683,I327691,I327708,I327725,I327742,I327759,I327790,I327807,I327824,I327841,I327886,I327931,I327948,I327965,I327996,I328013,I328030,I328056,I328064,I328109,I328126,I328143,I328201,I698973,I328227,I328235,I328261,I328269,I698997,I328286,I698979,I328303,I328320,I698994,I328337,I328187,I328368,I328385,I328402,I698976,I328419,I698985,I328184,I328175,I328464,I328178,I328172,I328509,I698982,I328526,I328543,I328181,I328574,I698991,I328591,I699000,I328608,I698988,I328634,I328642,I328169,I328193,I328687,I328704,I328721,I328190,I328779,I544736,I328805,I328813,I544727,I328839,I328847,I544721,I328864,I544733,I328881,I328898,I544724,I328915,I328765,I328946,I328963,I328980,I544730,I328997,I544715,I328762,I328753,I329042,I328756,I328750,I329087,I329104,I329121,I328759,I329152,I544718,I329169,I329186,I329212,I329220,I328747,I328771,I329265,I329282,I329299,I328768,I329357,I671139,I329383,I329391,I671151,I329417,I329425,I671142,I329442,I671130,I329459,I329476,I671127,I329493,I329524,I329541,I329558,I671133,I329575,I329620,I329665,I671148,I329682,I329699,I329730,I671136,I329747,I329764,I671145,I329790,I329798,I329843,I329860,I329877,I329935,I357069,I329961,I329969,I357081,I329995,I330003,I357072,I330020,I357075,I330037,I330054,I357078,I330071,I330102,I330119,I330136,I330153,I357084,I330198,I330243,I357090,I330260,I330277,I330308,I330325,I357087,I330342,I357093,I330368,I330376,I330421,I330438,I330455,I330513,I330539,I330547,I330573,I330581,I330598,I330615,I330632,I330649,I330499,I330680,I330697,I330714,I330731,I330496,I330487,I330776,I330490,I330484,I330821,I330838,I330855,I330493,I330886,I330903,I330920,I330946,I330954,I330481,I330505,I330999,I331016,I331033,I330502,I331091,I331117,I331125,I331151,I331159,I331176,I331193,I331210,I331227,I331077,I331258,I331275,I331292,I331309,I331074,I331065,I331354,I331068,I331062,I331399,I331416,I331433,I331071,I331464,I331481,I331498,I331524,I331532,I331059,I331083,I331577,I331594,I331611,I331080,I331669,I502204,I331695,I331703,I502201,I331729,I331737,I502198,I331754,I502225,I331771,I331788,I502213,I331805,I331655,I331836,I331853,I331870,I502219,I331887,I502210,I331652,I331643,I331932,I331646,I331640,I331977,I502207,I331994,I332011,I331649,I332042,I502222,I332059,I502216,I332076,I332102,I332110,I331637,I331661,I332155,I332172,I332189,I331658,I332247,I447617,I332273,I332281,I332307,I332315,I447614,I332332,I447629,I332349,I332366,I447623,I332383,I332414,I332431,I332448,I447620,I332465,I447611,I332510,I332555,I447632,I332572,I332589,I332620,I332637,I332654,I447626,I332680,I332688,I332733,I332750,I332767,I332825,I574567,I332851,I332859,I574573,I332885,I332893,I332910,I574570,I332927,I332944,I574588,I332961,I332811,I332992,I333009,I333026,I574591,I333043,I332808,I332799,I333088,I332802,I332796,I333133,I574576,I333150,I333167,I332805,I333198,I574582,I333215,I574579,I333232,I574585,I333258,I333266,I332793,I332817,I333311,I333328,I333345,I332814,I333403,I430226,I333429,I333437,I333463,I333471,I430223,I333488,I430238,I333505,I333522,I430232,I333539,I333570,I333587,I333604,I430229,I333621,I430220,I333666,I333711,I430241,I333728,I333745,I333776,I333793,I333810,I430235,I333836,I333844,I333889,I333906,I333923,I333981,I334007,I334015,I334041,I334049,I334066,I334083,I334100,I334117,I334148,I334165,I334182,I334199,I334244,I334289,I334306,I334323,I334354,I334371,I334388,I334414,I334422,I334467,I334484,I334501,I334559,I334585,I334593,I334619,I334627,I334644,I334661,I334678,I334695,I334545,I334726,I334743,I334760,I334777,I334542,I334533,I334822,I334536,I334530,I334867,I334884,I334901,I334539,I334932,I334949,I334966,I334992,I335000,I334527,I334551,I335045,I335062,I335079,I334548,I335137,I387703,I335163,I335171,I387715,I335197,I335205,I387706,I335222,I387709,I335239,I335256,I387712,I335273,I335123,I335304,I335321,I335338,I335355,I387718,I335120,I335111,I335400,I335114,I335108,I335445,I387724,I335462,I335479,I335117,I335510,I335527,I387721,I335544,I387727,I335570,I335578,I335105,I335129,I335623,I335640,I335657,I335126,I335715,I335741,I335749,I335775,I335783,I335800,I335817,I335834,I335851,I335701,I335882,I335899,I335916,I335933,I335698,I335689,I335978,I335692,I335686,I336023,I336040,I336057,I335695,I336088,I336105,I336122,I336148,I336156,I335683,I335707,I336201,I336218,I336235,I335704,I336293,I336319,I336327,I336353,I336361,I336378,I336395,I336412,I336429,I336460,I336477,I336494,I336511,I336556,I336601,I336618,I336635,I336666,I336683,I336700,I336726,I336734,I336779,I336796,I336813,I336871,I425851,I336897,I336905,I425863,I336931,I336939,I425854,I336956,I425857,I336973,I336990,I425860,I337007,I336857,I337038,I337055,I337072,I337089,I425866,I336854,I336845,I337134,I336848,I336842,I337179,I425872,I337196,I337213,I336851,I337244,I337261,I425869,I337278,I425875,I337304,I337312,I336839,I336863,I337357,I337374,I337391,I336860,I337449,I337475,I337483,I337509,I337517,I337534,I337551,I337568,I337585,I337616,I337633,I337650,I337667,I337712,I337757,I337774,I337791,I337822,I337839,I337856,I337882,I337890,I337935,I337952,I337969,I338027,I338053,I338061,I338087,I338095,I338112,I338129,I338146,I338163,I338013,I338194,I338211,I338228,I338245,I338010,I338001,I338290,I338004,I337998,I338335,I338352,I338369,I338007,I338400,I338417,I338434,I338460,I338468,I337995,I338019,I338513,I338530,I338547,I338016,I338605,I338631,I338639,I338665,I338673,I338690,I338707,I338724,I338741,I338772,I338789,I338806,I338823,I338868,I338913,I338930,I338947,I338978,I338995,I339012,I339038,I339046,I339091,I339108,I339125,I339183,I466589,I339209,I339217,I339243,I339251,I466586,I339268,I466601,I339285,I339302,I466595,I339319,I339350,I339367,I339384,I466592,I339401,I466583,I339446,I339491,I466604,I339508,I339525,I339556,I339573,I339590,I466598,I339616,I339624,I339669,I339686,I339703,I339761,I537734,I339787,I339795,I537731,I339821,I339829,I537728,I339846,I537755,I339863,I339880,I537743,I339897,I339747,I339928,I339945,I339962,I537749,I339979,I537740,I339744,I339735,I340024,I339738,I339732,I340069,I537737,I340086,I340103,I339741,I340134,I537752,I340151,I537746,I340168,I340194,I340202,I339729,I339753,I340247,I340264,I340281,I339750,I340339,I707303,I340365,I340373,I340399,I340407,I707327,I340424,I707309,I340441,I340458,I707324,I340475,I340506,I340523,I340540,I707306,I340557,I707315,I340602,I340647,I707312,I340664,I340681,I340712,I707321,I340729,I707330,I340746,I707318,I340772,I340780,I340825,I340842,I340859,I340917,I484116,I340943,I340951,I484113,I340977,I340985,I484110,I341002,I484137,I341019,I341036,I484125,I341053,I340903,I341084,I341101,I341118,I484131,I341135,I484122,I340900,I340891,I341180,I340894,I340888,I341225,I484119,I341242,I341259,I340897,I341290,I484134,I341307,I484128,I341324,I341350,I341358,I340885,I340909,I341403,I341420,I341437,I340906,I341495,I341521,I341529,I341555,I341563,I341580,I341597,I341614,I341631,I341481,I341662,I341679,I341696,I341713,I341478,I341469,I341758,I341472,I341466,I341803,I341820,I341837,I341475,I341868,I341885,I341902,I341928,I341936,I341463,I341487,I341981,I341998,I342015,I341484,I342073,I472386,I342099,I342107,I342133,I342141,I472383,I342158,I472398,I342175,I342192,I472392,I342209,I342240,I342257,I342274,I472389,I342291,I472380,I342336,I342381,I472401,I342398,I342415,I342446,I342463,I342480,I472395,I342506,I342514,I342559,I342576,I342593,I342651,I342677,I342685,I342711,I342719,I342736,I342753,I342770,I342787,I342818,I342835,I342852,I342869,I342914,I342959,I342976,I342993,I343024,I343041,I343058,I343084,I343092,I343137,I343154,I343171,I343229,I343255,I343263,I343289,I343297,I343314,I343331,I343348,I343365,I343396,I343413,I343430,I343447,I343492,I343537,I343554,I343571,I343602,I343619,I343636,I343662,I343670,I343715,I343732,I343749,I343807,I343833,I343841,I343867,I343875,I343892,I343909,I343926,I343943,I343793,I343974,I343991,I344008,I344025,I343790,I343781,I344070,I343784,I343778,I344115,I344132,I344149,I343787,I344180,I344197,I344214,I344240,I344248,I343775,I343799,I344293,I344310,I344327,I343796,I344385,I560444,I344411,I344419,I560435,I344445,I344453,I560429,I344470,I560441,I344487,I344504,I560432,I344521,I344552,I344569,I344586,I560438,I344603,I560423,I344648,I344693,I344710,I344727,I344758,I560426,I344775,I344792,I344818,I344826,I344871,I344888,I344905,I344963,I369785,I344989,I344997,I369797,I345023,I345031,I369788,I345048,I369791,I345065,I345082,I369794,I345099,I344949,I345130,I345147,I345164,I345181,I369800,I344946,I344937,I345226,I344940,I344934,I345271,I369806,I345288,I345305,I344943,I345336,I345353,I369803,I345370,I369809,I345396,I345404,I344931,I344955,I345449,I345466,I345483,I344952,I345541,I469224,I345567,I345575,I345601,I345609,I469221,I345626,I469236,I345643,I345660,I469230,I345677,I345527,I345708,I345725,I345742,I469227,I345759,I469218,I345524,I345515,I345804,I345518,I345512,I345849,I469239,I345866,I345883,I345521,I345914,I345931,I345948,I469233,I345974,I345982,I345509,I345533,I346027,I346044,I346061,I345530,I346119,I671717,I346145,I346153,I671729,I346179,I346187,I671720,I346204,I671708,I346221,I346238,I671705,I346255,I346105,I346286,I346303,I346320,I671711,I346337,I346102,I346093,I346382,I346096,I346090,I346427,I671726,I346444,I346461,I346099,I346492,I671714,I346509,I346526,I671723,I346552,I346560,I346087,I346111,I346605,I346622,I346639,I346108,I346697,I346723,I346731,I346748,I346765,I346791,I346799,I346825,I346833,I346850,I346867,I346884,I346924,I346932,I346949,I346966,I346983,I347014,I347031,I347057,I347065,I347096,I347127,I347144,I347175,I347275,I541355,I347301,I347309,I347326,I541352,I541370,I347343,I541367,I347369,I347377,I541349,I347403,I347411,I347428,I347445,I347462,I541361,I347502,I347510,I347527,I347544,I347561,I347592,I541364,I347609,I347635,I347643,I347674,I347705,I347722,I347753,I541358,I347853,I347879,I347887,I347904,I347921,I347947,I347955,I347981,I347989,I348006,I348023,I348040,I348080,I348088,I348105,I348122,I348139,I348170,I348187,I348213,I348221,I348252,I348283,I348300,I348331,I348431,I348457,I348465,I348482,I348499,I348525,I348533,I348559,I348567,I348584,I348601,I348618,I348658,I348666,I348683,I348700,I348717,I348748,I348765,I348791,I348799,I348830,I348861,I348878,I348909,I349009,I349035,I349043,I349060,I349077,I349103,I349111,I349137,I349145,I349162,I349179,I349196,I348992,I349236,I349244,I349261,I349278,I349295,I348995,I349326,I349343,I349369,I349377,I348977,I349408,I348986,I349439,I349456,I348998,I349487,I348989,I348980,I348983,I349001,I349587,I349613,I349621,I349638,I349655,I349681,I349689,I349715,I349723,I349740,I349757,I349774,I349570,I349814,I349822,I349839,I349856,I349873,I349573,I349904,I349921,I349947,I349955,I349555,I349986,I349564,I350017,I350034,I349576,I350065,I349567,I349558,I349561,I349579,I350165,I350191,I350199,I350216,I350233,I350259,I350267,I350293,I350301,I350318,I350335,I350352,I350392,I350400,I350417,I350434,I350451,I350482,I350499,I350525,I350533,I350564,I350595,I350612,I350643,I350743,I500284,I350769,I350777,I350794,I500260,I500275,I350811,I500287,I350837,I350845,I500272,I500263,I350871,I350879,I350896,I350913,I350930,I350726,I350970,I350978,I350995,I351012,I351029,I350729,I351060,I500278,I500269,I351077,I500281,I351103,I351111,I350711,I351142,I350720,I351173,I351190,I350732,I351221,I500266,I350723,I350714,I350717,I350735,I351321,I351347,I351355,I351372,I351389,I351415,I351423,I351449,I351457,I351474,I351491,I351508,I351548,I351556,I351573,I351590,I351607,I351638,I351655,I351681,I351689,I351720,I351751,I351768,I351799,I351899,I351925,I351933,I351950,I351967,I351993,I352001,I352027,I352035,I352052,I352069,I352086,I352126,I352134,I352151,I352168,I352185,I352216,I352233,I352259,I352267,I352298,I352329,I352346,I352377,I352477,I352503,I352511,I352528,I352545,I352571,I352579,I352605,I352613,I352630,I352647,I352664,I352704,I352712,I352729,I352746,I352763,I352794,I352811,I352837,I352845,I352876,I352907,I352924,I352955,I353055,I712685,I353081,I353089,I353106,I712670,I712658,I353123,I712673,I353149,I353157,I712676,I353183,I353191,I353208,I353225,I353242,I712664,I353282,I353290,I353307,I353324,I353341,I353372,I712661,I712667,I353389,I712682,I353415,I353423,I353454,I353485,I353502,I353533,I712679,I353633,I583833,I353659,I353667,I353684,I583815,I583827,I353701,I583830,I353727,I353735,I583824,I583821,I353761,I353769,I353786,I353803,I353820,I583839,I353860,I353868,I353885,I353902,I353919,I353950,I583818,I353967,I353993,I354001,I354032,I354063,I354080,I354111,I583836,I354211,I354237,I354245,I354262,I354279,I354305,I354313,I354339,I354347,I354364,I354381,I354398,I354194,I354438,I354446,I354463,I354480,I354497,I354197,I354528,I354545,I354571,I354579,I354179,I354610,I354188,I354641,I354658,I354200,I354689,I354191,I354182,I354185,I354203,I354789,I354815,I354823,I354840,I354857,I354883,I354891,I354917,I354925,I354942,I354959,I354976,I354772,I355016,I355024,I355041,I355058,I355075,I354775,I355106,I355123,I355149,I355157,I354757,I355188,I354766,I355219,I355236,I354778,I355267,I354769,I354760,I354763,I354781,I355367,I355393,I355401,I355418,I355435,I355461,I355469,I355495,I355503,I355520,I355537,I355554,I355594,I355602,I355619,I355636,I355653,I355684,I355701,I355727,I355735,I355766,I355797,I355814,I355845,I355945,I355971,I355979,I355996,I356013,I356039,I356047,I356073,I356081,I356098,I356115,I356132,I356172,I356180,I356197,I356214,I356231,I356262,I356279,I356305,I356313,I356344,I356375,I356392,I356423,I356523,I356549,I356557,I356574,I356591,I356617,I356625,I356651,I356659,I356676,I356693,I356710,I356506,I356750,I356758,I356775,I356792,I356809,I356509,I356840,I356857,I356883,I356891,I356491,I356922,I356500,I356953,I356970,I356512,I357001,I356503,I356494,I356497,I356515,I357101,I357127,I357135,I357152,I357169,I357195,I357203,I357229,I357237,I357254,I357271,I357288,I357328,I357336,I357353,I357370,I357387,I357418,I357435,I357461,I357469,I357500,I357531,I357548,I357579,I357679,I686663,I357705,I357713,I357730,I686651,I686669,I357747,I686660,I357773,I357781,I686675,I686672,I357807,I357815,I357832,I357849,I357866,I686654,I357906,I357914,I357931,I357948,I357965,I357996,I686648,I358013,I686657,I358039,I358047,I358078,I358109,I358126,I358157,I686666,I358257,I358283,I358291,I358308,I358325,I358351,I358359,I358385,I358393,I358410,I358427,I358444,I358484,I358492,I358509,I358526,I358543,I358574,I358591,I358617,I358625,I358656,I358687,I358704,I358735,I358835,I728750,I358861,I358869,I358886,I728735,I728723,I358903,I728738,I358929,I358937,I728741,I358963,I358971,I358988,I359005,I359022,I358818,I728729,I359062,I359070,I359087,I359104,I359121,I358821,I359152,I728726,I728732,I359169,I728747,I359195,I359203,I358803,I359234,I358812,I359265,I359282,I358824,I359313,I728744,I358815,I358806,I358809,I358827,I359413,I624293,I359439,I359447,I359464,I624275,I624287,I359481,I624290,I359507,I359515,I624284,I624281,I359541,I359549,I359566,I359583,I359600,I359396,I624299,I359640,I359648,I359665,I359682,I359699,I359399,I359730,I624278,I359747,I359773,I359781,I359381,I359812,I359390,I359843,I359860,I359402,I359891,I624296,I359393,I359384,I359387,I359405,I359991,I360017,I360025,I360042,I360059,I360085,I360093,I360119,I360127,I360144,I360161,I360178,I359974,I360218,I360226,I360243,I360260,I360277,I359977,I360308,I360325,I360351,I360359,I359959,I360390,I359968,I360421,I360438,I359980,I360469,I359971,I359962,I359965,I359983,I360569,I360595,I360603,I360620,I360637,I360663,I360671,I360697,I360705,I360722,I360739,I360756,I360552,I360796,I360804,I360821,I360838,I360855,I360555,I360886,I360903,I360929,I360937,I360537,I360968,I360546,I360999,I361016,I360558,I361047,I360549,I360540,I360543,I360561,I361147,I361173,I361181,I361198,I361215,I361241,I361249,I361275,I361283,I361300,I361317,I361334,I361130,I361374,I361382,I361399,I361416,I361433,I361133,I361464,I361481,I361507,I361515,I361115,I361546,I361124,I361577,I361594,I361136,I361625,I361127,I361118,I361121,I361139,I361725,I592503,I361751,I361759,I361776,I592485,I592497,I361793,I592500,I361819,I361827,I592494,I592491,I361853,I361861,I361878,I361895,I361912,I592509,I361952,I361960,I361977,I361994,I362011,I362042,I592488,I362059,I362085,I362093,I362124,I362155,I362172,I362203,I592506,I362303,I362329,I362337,I362354,I362371,I362397,I362405,I362431,I362439,I362456,I362473,I362490,I362530,I362538,I362555,I362572,I362589,I362620,I362637,I362663,I362671,I362702,I362733,I362750,I362781,I362881,I362907,I362915,I362932,I362949,I362975,I362983,I363009,I363017,I363034,I363051,I363068,I362864,I363108,I363116,I363133,I363150,I363167,I362867,I363198,I363215,I363241,I363249,I362849,I363280,I362858,I363311,I363328,I362870,I363359,I362861,I362852,I362855,I362873,I363459,I363485,I363493,I363510,I363527,I363553,I363561,I363587,I363595,I363612,I363629,I363646,I363686,I363694,I363711,I363728,I363745,I363776,I363793,I363819,I363827,I363858,I363889,I363906,I363937,I364037,I364063,I364071,I364088,I364105,I364131,I364139,I364165,I364173,I364190,I364207,I364224,I364264,I364272,I364289,I364306,I364323,I364354,I364371,I364397,I364405,I364436,I364467,I364484,I364515,I364615,I364641,I364649,I364666,I364683,I364709,I364717,I364743,I364751,I364768,I364785,I364802,I364598,I364842,I364850,I364867,I364884,I364901,I364601,I364932,I364949,I364975,I364983,I364583,I365014,I364592,I365045,I365062,I364604,I365093,I364595,I364586,I364589,I364607,I365193,I365219,I365227,I365244,I365261,I365287,I365295,I365321,I365329,I365346,I365363,I365380,I365420,I365428,I365445,I365462,I365479,I365510,I365527,I365553,I365561,I365592,I365623,I365640,I365671,I365771,I365797,I365805,I365822,I365839,I365865,I365873,I365899,I365907,I365924,I365941,I365958,I365998,I366006,I366023,I366040,I366057,I366088,I366105,I366131,I366139,I366170,I366201,I366218,I366249,I366349,I658309,I366375,I366383,I366400,I658312,I658321,I366417,I658324,I366443,I366451,I658333,I658315,I366477,I366485,I366502,I366519,I366536,I366332,I366576,I366584,I366601,I366618,I366635,I366335,I366666,I658330,I366683,I658327,I366709,I366717,I366317,I366748,I366326,I366779,I366796,I366338,I366827,I658318,I366329,I366320,I366323,I366341,I366927,I702570,I366953,I366961,I366978,I702555,I702543,I366995,I702558,I367021,I367029,I702561,I367055,I367063,I367080,I367097,I367114,I702549,I367154,I367162,I367179,I367196,I367213,I367244,I702546,I702552,I367261,I702567,I367287,I367295,I367326,I367357,I367374,I367405,I702564,I367505,I549770,I367531,I367539,I367556,I549767,I549785,I367573,I549782,I367599,I367607,I549764,I367633,I367641,I367658,I367675,I367692,I549776,I367732,I367740,I367757,I367774,I367791,I367822,I549779,I367839,I367865,I367873,I367904,I367935,I367952,I367983,I549773,I368083,I368109,I368117,I368134,I368151,I368177,I368185,I368211,I368219,I368236,I368253,I368270,I368310,I368318,I368335,I368352,I368369,I368400,I368417,I368443,I368451,I368482,I368513,I368530,I368561,I368661,I492532,I368687,I368695,I368712,I492508,I492523,I368729,I492535,I368755,I368763,I492520,I492511,I368789,I368797,I368814,I368831,I368848,I368644,I368888,I368896,I368913,I368930,I368947,I368647,I368978,I492526,I492517,I368995,I492529,I369021,I369029,I368629,I369060,I368638,I369091,I369108,I368650,I369139,I492514,I368641,I368632,I368635,I368653,I369239,I369265,I369273,I369290,I369307,I369333,I369341,I369367,I369375,I369392,I369409,I369426,I369466,I369474,I369491,I369508,I369525,I369556,I369573,I369599,I369607,I369638,I369669,I369686,I369717,I369817,I369843,I369851,I369868,I369885,I369911,I369919,I369945,I369953,I369970,I369987,I370004,I370044,I370052,I370069,I370086,I370103,I370134,I370151,I370177,I370185,I370216,I370247,I370264,I370295,I370395,I580365,I370421,I370429,I370446,I580347,I580359,I370463,I580362,I370489,I370497,I580356,I580353,I370523,I370531,I370548,I370565,I370582,I580371,I370622,I370630,I370647,I370664,I370681,I370712,I580350,I370729,I370755,I370763,I370794,I370825,I370842,I370873,I580368,I370973,I370999,I371007,I371024,I371041,I371067,I371075,I371101,I371109,I371126,I371143,I371160,I370956,I371200,I371208,I371225,I371242,I371259,I370959,I371290,I371307,I371333,I371341,I370941,I371372,I370950,I371403,I371420,I370962,I371451,I370953,I370944,I370947,I370965,I371551,I488010,I371577,I371585,I371602,I487986,I488001,I371619,I488013,I371645,I371653,I487998,I487989,I371679,I371687,I371704,I371721,I371738,I371778,I371786,I371803,I371820,I371837,I371868,I488004,I487995,I371885,I488007,I371911,I371919,I371950,I371981,I371998,I372029,I487992,I372129,I476084,I372155,I372163,I372180,I476072,I476090,I372197,I476087,I372223,I372231,I476078,I476075,I372257,I372265,I372282,I372299,I372316,I476069,I372356,I372364,I372381,I372398,I372415,I372446,I372463,I372489,I372497,I372528,I372559,I372576,I372607,I476081,I372707,I372733,I372741,I372758,I372775,I372801,I372809,I372835,I372843,I372860,I372877,I372894,I372690,I372934,I372942,I372959,I372976,I372993,I372693,I373024,I373041,I373067,I373075,I372675,I373106,I372684,I373137,I373154,I372696,I373185,I372687,I372678,I372681,I372699,I373285,I373311,I373319,I373336,I373353,I373379,I373387,I373413,I373421,I373438,I373455,I373472,I373512,I373520,I373537,I373554,I373571,I373602,I373619,I373645,I373653,I373684,I373715,I373732,I373763,I373863,I373889,I373897,I373914,I373931,I373957,I373965,I373991,I373999,I374016,I374033,I374050,I374090,I374098,I374115,I374132,I374149,I374180,I374197,I374223,I374231,I374262,I374293,I374310,I374341,I374441,I374467,I374475,I374492,I374509,I374535,I374543,I374569,I374577,I374594,I374611,I374628,I374424,I374668,I374676,I374693,I374710,I374727,I374427,I374758,I374775,I374801,I374809,I374409,I374840,I374418,I374871,I374888,I374430,I374919,I374421,I374412,I374415,I374433,I375019,I375045,I375053,I375070,I375087,I375113,I375121,I375147,I375155,I375172,I375189,I375206,I375002,I375246,I375254,I375271,I375288,I375305,I375005,I375336,I375353,I375379,I375387,I374987,I375418,I374996,I375449,I375466,I375008,I375497,I374999,I374990,I374993,I375011,I375597,I681531,I375623,I375631,I375648,I681555,I681537,I375665,I681543,I375691,I375699,I681549,I681534,I375725,I375733,I375750,I375767,I375784,I681546,I375824,I375832,I375849,I375866,I375883,I375914,I681552,I681540,I375931,I375957,I375965,I375996,I376027,I376044,I376075,I376175,I376201,I376209,I376226,I376243,I376269,I376277,I376303,I376311,I376328,I376345,I376362,I376158,I376402,I376410,I376427,I376444,I376461,I376161,I376492,I376509,I376535,I376543,I376143,I376574,I376152,I376605,I376622,I376164,I376653,I376155,I376146,I376149,I376167,I376753,I563795,I376779,I376787,I376804,I563792,I563810,I376821,I563807,I376847,I376855,I563789,I376881,I376889,I376906,I376923,I376940,I563801,I376980,I376988,I377005,I377022,I377039,I377070,I563804,I377087,I377113,I377121,I377152,I377183,I377200,I377231,I563798,I377331,I724585,I377357,I377365,I377382,I724570,I724558,I377399,I724573,I377425,I377433,I724576,I377459,I377467,I377484,I377501,I377518,I724564,I377558,I377566,I377583,I377600,I377617,I377648,I724561,I724567,I377665,I724582,I377691,I377699,I377730,I377761,I377778,I377809,I724579,I377909,I377935,I377943,I377960,I377977,I378003,I378011,I378037,I378045,I378062,I378079,I378096,I377892,I378136,I378144,I378161,I378178,I378195,I377895,I378226,I378243,I378269,I378277,I377877,I378308,I377886,I378339,I378356,I377898,I378387,I377889,I377880,I377883,I377901,I378487,I663205,I378513,I378521,I378538,I663208,I663217,I378555,I663220,I378581,I378589,I663229,I663211,I378615,I378623,I378640,I378657,I378674,I378470,I378714,I378722,I378739,I378756,I378773,I378473,I378804,I663226,I378821,I663223,I378847,I378855,I378455,I378886,I378464,I378917,I378934,I378476,I378965,I663214,I378467,I378458,I378461,I378479,I379065,I693050,I379091,I379099,I379116,I693035,I693023,I379133,I693038,I379159,I379167,I693041,I379193,I379201,I379218,I379235,I379252,I379048,I693029,I379292,I379300,I379317,I379334,I379351,I379051,I379382,I693026,I693032,I379399,I693047,I379425,I379433,I379033,I379464,I379042,I379495,I379512,I379054,I379543,I693044,I379045,I379036,I379039,I379057,I379643,I497054,I379669,I379677,I379694,I497030,I497045,I379711,I497057,I379737,I379745,I497042,I497033,I379771,I379779,I379796,I379813,I379830,I379870,I379878,I379895,I379912,I379929,I379960,I497048,I497039,I379977,I497051,I380003,I380011,I380042,I380073,I380090,I380121,I497036,I380221,I572851,I380247,I380255,I380272,I572833,I572845,I380289,I572848,I380315,I380323,I572842,I572839,I380349,I380357,I380374,I380391,I380408,I572857,I380448,I380456,I380473,I380490,I380507,I380538,I572836,I380555,I380581,I380589,I380620,I380651,I380668,I380699,I572854,I380799,I380825,I380833,I380850,I380867,I380893,I380901,I380927,I380935,I380952,I380969,I380986,I381026,I381034,I381051,I381068,I381085,I381116,I381133,I381159,I381167,I381198,I381229,I381246,I381277,I381377,I381403,I381411,I381428,I381445,I381471,I381479,I381505,I381513,I381530,I381547,I381564,I381360,I381604,I381612,I381629,I381646,I381663,I381363,I381694,I381711,I381737,I381745,I381345,I381776,I381354,I381807,I381824,I381366,I381855,I381357,I381348,I381351,I381369,I381955,I381981,I381989,I382006,I382023,I382049,I382057,I382083,I382091,I382108,I382125,I382142,I381938,I382182,I382190,I382207,I382224,I382241,I381941,I382272,I382289,I382315,I382323,I381923,I382354,I381932,I382385,I382402,I381944,I382433,I381935,I381926,I381929,I381947,I382533,I382559,I382567,I382584,I382601,I382627,I382635,I382661,I382669,I382686,I382703,I382720,I382516,I382760,I382768,I382785,I382802,I382819,I382519,I382850,I382867,I382893,I382901,I382501,I382932,I382510,I382963,I382980,I382522,I383011,I382513,I382504,I382507,I382525,I383111,I559307,I383137,I383145,I383162,I559304,I559322,I383179,I559319,I383205,I383213,I559301,I383239,I383247,I383264,I383281,I383298,I383094,I559313,I383338,I383346,I383363,I383380,I383397,I383097,I383428,I559316,I383445,I383471,I383479,I383079,I383510,I383088,I383541,I383558,I383100,I383589,I559310,I383091,I383082,I383085,I383103,I383689,I383715,I383723,I383740,I383757,I383783,I383791,I383817,I383825,I383842,I383859,I383876,I383672,I383916,I383924,I383941,I383958,I383975,I383675,I384006,I384023,I384049,I384057,I383657,I384088,I383666,I384119,I384136,I383678,I384167,I383669,I383660,I383663,I383681,I384267,I384293,I384301,I384318,I384335,I384361,I384369,I384395,I384403,I384420,I384437,I384454,I384250,I384494,I384502,I384519,I384536,I384553,I384253,I384584,I384601,I384627,I384635,I384235,I384666,I384244,I384697,I384714,I384256,I384745,I384247,I384238,I384241,I384259,I384845,I706140,I384871,I384879,I384896,I706125,I706113,I384913,I706128,I384939,I384947,I706131,I384973,I384981,I384998,I385015,I385032,I706119,I385072,I385080,I385097,I385114,I385131,I385162,I706116,I706122,I385179,I706137,I385205,I385213,I385244,I385275,I385292,I385323,I706134,I385423,I454477,I385449,I385457,I385474,I454465,I454483,I385491,I454480,I385517,I385525,I454471,I454468,I385551,I385559,I385576,I385593,I385610,I385406,I454462,I385650,I385658,I385675,I385692,I385709,I385409,I385740,I385757,I385783,I385791,I385391,I385822,I385400,I385853,I385870,I385412,I385901,I454474,I385403,I385394,I385397,I385415,I386001,I386027,I386035,I386052,I386069,I386095,I386103,I386129,I386137,I386154,I386171,I386188,I385984,I386228,I386236,I386253,I386270,I386287,I385987,I386318,I386335,I386361,I386369,I385969,I386400,I385978,I386431,I386448,I385990,I386479,I385981,I385972,I385975,I385993,I386579,I530000,I386605,I386613,I386630,I529976,I529991,I386647,I530003,I386673,I386681,I529988,I529979,I386707,I386715,I386732,I386749,I386766,I386806,I386814,I386831,I386848,I386865,I386896,I529994,I529985,I386913,I529997,I386939,I386947,I386978,I387009,I387026,I387057,I529982,I387157,I387183,I387191,I387208,I387225,I387251,I387259,I387285,I387293,I387310,I387327,I387344,I387140,I387384,I387392,I387409,I387426,I387443,I387143,I387474,I387491,I387517,I387525,I387125,I387556,I387134,I387587,I387604,I387146,I387635,I387137,I387128,I387131,I387149,I387735,I387761,I387769,I387786,I387803,I387829,I387837,I387863,I387871,I387888,I387905,I387922,I387962,I387970,I387987,I388004,I388021,I388052,I388069,I388095,I388103,I388134,I388165,I388182,I388213,I388313,I638725,I388339,I388347,I388364,I638728,I638737,I388381,I638740,I388407,I388415,I638749,I638731,I388441,I388449,I388466,I388483,I388500,I388296,I388540,I388548,I388565,I388582,I388599,I388299,I388630,I638746,I388647,I638743,I388673,I388681,I388281,I388712,I388290,I388743,I388760,I388302,I388791,I638734,I388293,I388284,I388287,I388305,I388891,I388917,I388925,I388942,I388959,I388985,I388993,I389019,I389027,I389044,I389061,I389078,I389118,I389126,I389143,I389160,I389177,I389208,I389225,I389251,I389259,I389290,I389321,I389338,I389369,I389469,I489948,I389495,I389503,I389520,I489924,I489939,I389537,I489951,I389563,I389571,I489936,I489927,I389597,I389605,I389622,I389639,I389656,I389452,I389696,I389704,I389721,I389738,I389755,I389455,I389786,I489942,I489933,I389803,I489945,I389829,I389837,I389437,I389868,I389446,I389899,I389916,I389458,I389947,I489930,I389449,I389440,I389443,I389461,I390047,I390073,I390081,I390098,I390115,I390141,I390149,I390175,I390183,I390200,I390217,I390234,I390030,I390274,I390282,I390299,I390316,I390333,I390033,I390364,I390381,I390407,I390415,I390015,I390446,I390024,I390477,I390494,I390036,I390525,I390027,I390018,I390021,I390039,I390625,I552014,I390651,I390659,I390676,I552011,I552029,I390693,I552026,I390719,I390727,I552008,I390753,I390761,I390778,I390795,I390812,I552020,I390852,I390860,I390877,I390894,I390911,I390942,I552023,I390959,I390985,I390993,I391024,I391055,I391072,I391103,I552017,I391203,I448680,I391229,I391237,I391254,I448668,I448686,I391271,I448683,I391297,I391305,I448674,I448671,I391331,I391339,I391356,I391373,I391390,I448665,I391430,I391438,I391455,I391472,I391489,I391520,I391537,I391563,I391571,I391602,I391633,I391650,I391681,I448677,I391781,I441829,I391807,I391815,I391832,I441817,I441835,I391849,I441832,I391875,I391883,I441823,I441820,I391909,I391917,I391934,I391951,I391968,I441814,I392008,I392016,I392033,I392050,I392067,I392098,I392115,I392141,I392149,I392180,I392211,I392228,I392259,I441826,I392359,I392385,I392393,I392410,I392427,I392453,I392461,I392487,I392495,I392512,I392529,I392546,I392342,I392586,I392594,I392611,I392628,I392645,I392345,I392676,I392693,I392719,I392727,I392327,I392758,I392336,I392789,I392806,I392348,I392837,I392339,I392330,I392333,I392351,I392937,I650149,I392963,I392971,I392988,I650152,I650161,I393005,I650164,I393031,I393039,I650173,I650155,I393065,I393073,I393090,I393107,I393124,I392920,I393164,I393172,I393189,I393206,I393223,I392923,I393254,I650170,I393271,I650167,I393297,I393305,I392905,I393336,I392914,I393367,I393384,I392926,I393415,I650158,I392917,I392908,I392911,I392929,I393515,I393541,I393549,I393566,I393583,I393609,I393617,I393643,I393651,I393668,I393685,I393702,I393742,I393750,I393767,I393784,I393801,I393832,I393849,I393875,I393883,I393914,I393945,I393962,I393993,I394093,I394119,I394127,I394144,I394161,I394187,I394195,I394221,I394229,I394246,I394263,I394280,I394076,I394320,I394328,I394345,I394362,I394379,I394079,I394410,I394427,I394453,I394461,I394061,I394492,I394070,I394523,I394540,I394082,I394571,I394073,I394064,I394067,I394085,I394671,I432870,I394697,I394705,I394722,I432858,I432876,I394739,I432873,I394765,I394773,I432864,I432861,I394799,I394807,I394824,I394841,I394858,I394654,I432855,I394898,I394906,I394923,I394940,I394957,I394657,I394988,I395005,I395031,I395039,I394639,I395070,I394648,I395101,I395118,I394660,I395149,I432867,I394651,I394642,I394645,I394663,I395249,I653413,I395275,I395283,I395300,I653416,I653425,I395317,I653428,I395343,I395351,I653437,I653419,I395377,I395385,I395402,I395419,I395436,I395232,I395476,I395484,I395501,I395518,I395535,I395235,I395566,I653434,I395583,I653431,I395609,I395617,I395217,I395648,I395226,I395679,I395696,I395238,I395727,I653422,I395229,I395220,I395223,I395241,I395827,I395853,I395861,I395878,I395895,I395921,I395929,I395955,I395963,I395980,I395997,I396014,I395810,I396054,I396062,I396079,I396096,I396113,I395813,I396144,I396161,I396187,I396195,I395795,I396226,I395804,I396257,I396274,I395816,I396305,I395807,I395798,I395801,I395819,I396405,I396431,I396439,I396456,I396473,I396499,I396507,I396533,I396541,I396558,I396575,I396592,I396388,I396632,I396640,I396657,I396674,I396691,I396391,I396722,I396739,I396765,I396773,I396373,I396804,I396382,I396835,I396852,I396394,I396883,I396385,I396376,I396379,I396397,I396983,I397009,I397017,I397034,I397051,I397077,I397085,I397111,I397119,I397136,I397153,I397170,I397210,I397218,I397235,I397252,I397269,I397300,I397317,I397343,I397351,I397382,I397413,I397430,I397461,I397561,I683265,I397587,I397595,I397612,I683289,I683271,I397629,I683277,I397655,I397663,I683283,I683268,I397689,I397697,I397714,I397731,I397748,I397544,I683280,I397788,I397796,I397813,I397830,I397847,I397547,I397878,I683286,I683274,I397895,I397921,I397929,I397529,I397960,I397538,I397991,I398008,I397550,I398039,I397541,I397532,I397535,I397553,I398139,I646341,I398165,I398173,I398190,I646344,I646353,I398207,I646356,I398233,I398241,I646365,I646347,I398267,I398275,I398292,I398309,I398326,I398366,I398374,I398391,I398408,I398425,I398456,I646362,I398473,I646359,I398499,I398507,I398538,I398569,I398586,I398617,I646350,I398717,I589613,I398743,I398751,I398768,I589595,I589607,I398785,I589610,I398811,I398819,I589604,I589601,I398845,I398853,I398870,I398887,I398904,I589619,I398944,I398952,I398969,I398986,I399003,I399034,I589598,I399051,I399077,I399085,I399116,I399147,I399164,I399195,I589616,I399295,I399321,I399329,I399346,I399363,I399389,I399397,I399423,I399431,I399448,I399465,I399482,I399522,I399530,I399547,I399564,I399581,I399612,I399629,I399655,I399663,I399694,I399725,I399742,I399773,I399873,I399899,I399907,I399924,I399941,I399967,I399975,I400001,I400009,I400026,I400043,I400060,I400100,I400108,I400125,I400142,I400159,I400190,I400207,I400233,I400241,I400272,I400303,I400320,I400351,I400451,I400477,I400485,I400502,I400519,I400545,I400553,I400579,I400587,I400604,I400621,I400638,I400678,I400686,I400703,I400720,I400737,I400768,I400785,I400811,I400819,I400850,I400881,I400898,I400929,I401029,I474503,I401055,I401063,I401080,I474491,I474509,I401097,I474506,I401123,I401131,I474497,I474494,I401157,I401165,I401182,I401199,I401216,I474488,I401256,I401264,I401281,I401298,I401315,I401346,I401363,I401389,I401397,I401428,I401459,I401476,I401507,I474500,I401607,I401633,I401641,I401658,I401675,I401701,I401709,I401735,I401743,I401760,I401777,I401794,I401834,I401842,I401859,I401876,I401893,I401924,I401941,I401967,I401975,I402006,I402037,I402054,I402085,I402185,I402211,I402219,I402236,I402253,I402279,I402287,I402313,I402321,I402338,I402355,I402372,I402412,I402420,I402437,I402454,I402471,I402502,I402519,I402545,I402553,I402584,I402615,I402632,I402663,I402763,I477138,I402789,I402797,I402814,I477126,I477144,I402831,I477141,I402857,I402865,I477132,I477129,I402891,I402899,I402916,I402933,I402950,I402746,I477123,I402990,I402998,I403015,I403032,I403049,I402749,I403080,I403097,I403123,I403131,I402731,I403162,I402740,I403193,I403210,I402752,I403241,I477135,I402743,I402734,I402737,I402755,I403341,I403367,I403375,I403392,I403409,I403435,I403443,I403469,I403477,I403494,I403511,I403528,I403324,I403568,I403576,I403593,I403610,I403627,I403327,I403658,I403675,I403701,I403709,I403309,I403740,I403318,I403771,I403788,I403330,I403819,I403321,I403312,I403315,I403333,I403919,I697810,I403945,I403953,I403970,I697795,I697783,I403987,I697798,I404013,I404021,I697801,I404047,I404055,I404072,I404089,I404106,I697789,I404146,I404154,I404171,I404188,I404205,I404236,I697786,I697792,I404253,I697807,I404279,I404287,I404318,I404349,I404366,I404397,I697804,I404497,I715065,I404523,I404531,I404548,I715050,I715038,I404565,I715053,I404591,I404599,I715056,I404625,I404633,I404650,I404667,I404684,I404480,I715044,I404724,I404732,I404749,I404766,I404783,I404483,I404814,I715041,I715047,I404831,I715062,I404857,I404865,I404465,I404896,I404474,I404927,I404944,I404486,I404975,I715059,I404477,I404468,I404471,I404489,I405075,I405101,I405109,I405126,I405143,I405169,I405177,I405203,I405211,I405228,I405245,I405262,I405302,I405310,I405327,I405344,I405361,I405392,I405409,I405435,I405443,I405474,I405505,I405522,I405553,I405653,I459747,I405679,I405687,I405704,I459735,I459753,I405721,I459750,I405747,I405755,I459741,I459738,I405781,I405789,I405806,I405823,I405840,I405636,I459732,I405880,I405888,I405905,I405922,I405939,I405639,I405970,I405987,I406013,I406021,I405621,I406052,I405630,I406083,I406100,I405642,I406131,I459744,I405633,I405624,I405627,I405645,I406231,I546965,I406257,I406265,I406282,I546962,I546980,I406299,I546977,I406325,I406333,I546959,I406359,I406367,I406384,I406401,I406418,I406214,I546971,I406458,I406466,I406483,I406500,I406517,I406217,I406548,I546974,I406565,I406591,I406599,I406199,I406630,I406208,I406661,I406678,I406220,I406709,I546968,I406211,I406202,I406205,I406223,I406809,I406835,I406843,I406860,I406877,I406903,I406911,I406937,I406945,I406962,I406979,I406996,I407036,I407044,I407061,I407078,I407095,I407126,I407143,I407169,I407177,I407208,I407239,I407256,I407287,I407387,I503514,I407413,I407421,I407438,I503490,I503505,I407455,I503517,I407481,I407489,I503502,I503493,I407515,I407523,I407540,I407557,I407574,I407614,I407622,I407639,I407656,I407673,I407704,I503508,I503499,I407721,I503511,I407747,I407755,I407786,I407817,I407834,I407865,I503496,I407965,I509328,I407991,I407999,I408016,I509304,I509319,I408033,I509331,I408059,I408067,I509316,I509307,I408093,I408101,I408118,I408135,I408152,I407948,I408192,I408200,I408217,I408234,I408251,I407951,I408282,I509322,I509313,I408299,I509325,I408325,I408333,I407933,I408364,I407942,I408395,I408412,I407954,I408443,I509310,I407945,I407936,I407939,I407957,I408543,I555380,I408569,I408577,I408594,I555377,I555395,I408611,I555392,I408637,I408645,I555374,I408671,I408679,I408696,I408713,I408730,I408526,I555386,I408770,I408778,I408795,I408812,I408829,I408529,I408860,I555389,I408877,I408903,I408911,I408511,I408942,I408520,I408973,I408990,I408532,I409021,I555383,I408523,I408514,I408517,I408535,I409121,I656133,I409147,I409155,I409172,I656136,I656145,I409189,I656148,I409215,I409223,I656157,I656139,I409249,I409257,I409274,I409291,I409308,I409348,I409356,I409373,I409390,I409407,I409438,I656154,I409455,I656151,I409481,I409489,I409520,I409551,I409568,I409599,I656142,I409699,I409725,I409733,I409750,I409767,I409793,I409801,I409827,I409835,I409852,I409869,I409886,I409682,I409926,I409934,I409951,I409968,I409985,I409685,I410016,I410033,I410059,I410067,I409667,I410098,I409676,I410129,I410146,I409688,I410177,I409679,I409670,I409673,I409691,I410277,I693645,I410303,I410311,I410328,I693630,I693618,I410345,I693633,I410371,I410379,I693636,I410405,I410413,I410430,I410447,I410464,I410260,I693624,I410504,I410512,I410529,I410546,I410563,I410263,I410594,I693621,I693627,I410611,I693642,I410637,I410645,I410245,I410676,I410254,I410707,I410724,I410266,I410755,I693639,I410257,I410248,I410251,I410269,I410855,I410881,I410889,I410906,I410923,I410949,I410957,I410983,I410991,I411008,I411025,I411042,I410838,I411082,I411090,I411107,I411124,I411141,I410841,I411172,I411189,I411215,I411223,I410823,I411254,I410832,I411285,I411302,I410844,I411333,I410835,I410826,I410829,I410847,I411433,I411459,I411467,I411484,I411501,I411527,I411535,I411561,I411569,I411586,I411603,I411620,I411660,I411668,I411685,I411702,I411719,I411750,I411767,I411793,I411801,I411832,I411863,I411880,I411911,I412011,I412037,I412045,I412062,I412079,I412105,I412113,I412139,I412147,I412164,I412181,I412198,I411994,I412238,I412246,I412263,I412280,I412297,I411997,I412328,I412345,I412371,I412379,I411979,I412410,I411988,I412441,I412458,I412000,I412489,I411991,I411982,I411985,I412003,I412589,I688346,I412615,I412623,I412640,I688334,I688352,I412657,I688343,I412683,I412691,I688358,I688355,I412717,I412725,I412742,I412759,I412776,I688337,I412816,I412824,I412841,I412858,I412875,I412906,I688331,I412923,I688340,I412949,I412957,I412988,I413019,I413036,I413067,I688349,I413167,I413193,I413201,I413218,I413235,I413261,I413269,I413295,I413303,I413320,I413337,I413354,I413150,I413394,I413402,I413419,I413436,I413453,I413153,I413484,I413501,I413527,I413535,I413135,I413566,I413144,I413597,I413614,I413156,I413645,I413147,I413138,I413141,I413159,I413745,I482196,I413771,I413779,I413796,I482172,I482187,I413813,I482199,I413839,I413847,I482184,I482175,I413873,I413881,I413898,I413915,I413932,I413728,I413972,I413980,I413997,I414014,I414031,I413731,I414062,I482190,I482181,I414079,I482193,I414105,I414113,I413713,I414144,I413722,I414175,I414192,I413734,I414223,I482178,I413725,I413716,I413719,I413737,I414323,I623715,I414349,I414357,I414374,I623697,I623709,I414391,I623712,I414417,I414425,I623706,I623703,I414451,I414459,I414476,I414493,I414510,I414306,I623721,I414550,I414558,I414575,I414592,I414609,I414309,I414640,I623700,I414657,I414683,I414691,I414291,I414722,I414300,I414753,I414770,I414312,I414801,I623718,I414303,I414294,I414297,I414315,I414901,I414927,I414935,I414952,I414969,I414995,I415003,I415029,I415037,I415054,I415071,I415088,I414884,I415128,I415136,I415153,I415170,I415187,I414887,I415218,I415235,I415261,I415269,I414869,I415300,I414878,I415331,I415348,I414890,I415379,I414881,I414872,I414875,I414893,I415479,I449207,I415505,I415513,I415530,I449195,I449213,I415547,I449210,I415573,I415581,I449201,I449198,I415607,I415615,I415632,I415649,I415666,I415462,I449192,I415706,I415714,I415731,I415748,I415765,I415465,I415796,I415813,I415839,I415847,I415447,I415878,I415456,I415909,I415926,I415468,I415957,I449204,I415459,I415450,I415453,I415471,I416057,I556502,I416083,I416091,I416108,I556499,I556517,I416125,I556514,I416151,I416159,I556496,I416185,I416193,I416210,I416227,I416244,I416040,I556508,I416284,I416292,I416309,I416326,I416343,I416043,I416374,I556511,I416391,I416417,I416425,I416025,I416456,I416034,I416487,I416504,I416046,I416535,I556505,I416037,I416028,I416031,I416049,I416635,I416661,I416669,I416686,I416703,I416729,I416737,I416763,I416771,I416788,I416805,I416822,I416618,I416862,I416870,I416887,I416904,I416921,I416621,I416952,I416969,I416995,I417003,I416603,I417034,I416612,I417065,I417082,I416624,I417113,I416615,I416606,I416609,I416627,I417213,I417239,I417247,I417264,I417281,I417307,I417315,I417341,I417349,I417366,I417383,I417400,I417196,I417440,I417448,I417465,I417482,I417499,I417199,I417530,I417547,I417573,I417581,I417181,I417612,I417190,I417643,I417660,I417202,I417691,I417193,I417184,I417187,I417205,I417791,I550892,I417817,I417825,I417842,I550889,I550907,I417859,I550904,I417885,I417893,I550886,I417919,I417927,I417944,I417961,I417978,I417774,I550898,I418018,I418026,I418043,I418060,I418077,I417777,I418108,I550901,I418125,I418151,I418159,I417759,I418190,I417768,I418221,I418238,I417780,I418269,I550895,I417771,I417762,I417765,I417783,I418369,I523540,I418395,I418403,I418420,I523516,I523531,I418437,I523543,I418463,I418471,I523528,I523519,I418497,I418505,I418522,I418539,I418556,I418596,I418604,I418621,I418638,I418655,I418686,I523534,I523525,I418703,I523537,I418729,I418737,I418768,I418799,I418816,I418847,I523522,I418947,I455004,I418973,I418981,I418998,I454992,I455010,I419015,I455007,I419041,I419049,I454998,I454995,I419075,I419083,I419100,I419117,I419134,I454989,I419174,I419182,I419199,I419216,I419233,I419264,I419281,I419307,I419315,I419346,I419377,I419394,I419425,I455001,I419525,I419551,I419559,I419576,I419593,I419619,I419627,I419653,I419661,I419678,I419695,I419712,I419508,I419752,I419760,I419777,I419794,I419811,I419511,I419842,I419859,I419885,I419893,I419493,I419924,I419502,I419955,I419972,I419514,I420003,I419505,I419496,I419499,I419517,I420103,I513204,I420129,I420137,I420154,I513180,I513195,I420171,I513207,I420197,I420205,I513192,I513183,I420231,I420239,I420256,I420273,I420290,I420330,I420338,I420355,I420372,I420389,I420420,I513198,I513189,I420437,I513201,I420463,I420471,I420502,I420533,I420550,I420581,I513186,I420681,I420707,I420715,I420732,I420749,I420775,I420783,I420809,I420817,I420834,I420851,I420868,I420664,I420908,I420916,I420933,I420950,I420967,I420667,I420998,I421015,I421041,I421049,I420649,I421080,I420658,I421111,I421128,I420670,I421159,I420661,I420652,I420655,I420673,I421259,I632385,I421285,I421293,I421310,I632367,I632379,I421327,I632382,I421353,I421361,I632376,I632373,I421387,I421395,I421412,I421429,I421446,I632391,I421486,I421494,I421511,I421528,I421545,I421576,I632370,I421593,I421619,I421627,I421658,I421689,I421706,I421737,I632388,I421837,I664293,I421863,I421871,I421888,I664296,I664305,I421905,I664308,I421931,I421939,I664317,I664299,I421965,I421973,I421990,I422007,I422024,I422064,I422072,I422089,I422106,I422123,I422154,I664314,I422171,I664311,I422197,I422205,I422236,I422267,I422284,I422315,I664302,I422415,I604063,I422441,I422449,I422466,I604045,I604057,I422483,I604060,I422509,I422517,I604054,I604051,I422543,I422551,I422568,I422585,I422602,I422398,I604069,I422642,I422650,I422667,I422684,I422701,I422401,I422732,I604048,I422749,I422775,I422783,I422383,I422814,I422392,I422845,I422862,I422404,I422893,I604066,I422395,I422386,I422389,I422407,I422993,I423019,I423027,I423044,I423061,I423087,I423095,I423121,I423129,I423146,I423163,I423180,I422976,I423220,I423228,I423245,I423262,I423279,I422979,I423310,I423327,I423353,I423361,I422961,I423392,I422970,I423423,I423440,I422982,I423471,I422973,I422964,I422967,I422985,I423571,I542477,I423597,I423605,I423622,I542474,I542492,I423639,I542489,I423665,I423673,I542471,I423699,I423707,I423724,I423741,I423758,I542483,I423798,I423806,I423823,I423840,I423857,I423888,I542486,I423905,I423931,I423939,I423970,I424001,I424018,I424049,I542480,I424149,I452896,I424175,I424183,I424200,I452884,I452902,I424217,I452899,I424243,I424251,I452890,I452887,I424277,I424285,I424302,I424319,I424336,I424132,I452881,I424376,I424384,I424401,I424418,I424435,I424135,I424466,I424483,I424509,I424517,I424117,I424548,I424126,I424579,I424596,I424138,I424627,I452893,I424129,I424120,I424123,I424141,I424727,I424753,I424761,I424778,I424795,I424821,I424829,I424855,I424863,I424880,I424897,I424914,I424710,I424954,I424962,I424979,I424996,I425013,I424713,I425044,I425061,I425087,I425095,I424695,I425126,I424704,I425157,I425174,I424716,I425205,I424707,I424698,I424701,I424719,I425305,I627761,I425331,I425339,I425356,I627743,I627755,I425373,I627758,I425399,I425407,I627752,I627749,I425433,I425441,I425458,I425475,I425492,I627767,I425532,I425540,I425557,I425574,I425591,I425622,I627746,I425639,I425665,I425673,I425704,I425735,I425752,I425783,I627764,I425883,I529354,I425909,I425917,I425934,I529330,I529345,I425951,I529357,I425977,I425985,I529342,I529333,I426011,I426019,I426036,I426053,I426070,I426110,I426118,I426135,I426152,I426169,I426200,I529348,I529339,I426217,I529351,I426243,I426251,I426282,I426313,I426330,I426361,I529336,I426461,I426487,I426495,I426512,I426529,I426555,I426563,I426589,I426597,I426614,I426631,I426648,I426444,I426688,I426696,I426713,I426730,I426747,I426447,I426778,I426795,I426821,I426829,I426429,I426860,I426438,I426891,I426908,I426450,I426939,I426441,I426432,I426435,I426453,I427039,I427065,I427073,I427090,I427107,I427133,I427141,I427167,I427175,I427192,I427209,I427226,I427266,I427274,I427291,I427308,I427325,I427356,I427373,I427399,I427407,I427438,I427469,I427486,I427517,I427614,I427640,I427648,I427665,I427682,I427708,I427739,I427747,I427764,I427790,I427798,I427838,I427874,I427891,I427917,I427925,I427942,I427973,I427990,I428007,I428038,I428069,I428086,I428141,I428167,I428175,I428192,I428209,I428235,I428266,I428274,I428291,I428317,I428325,I428365,I428401,I428418,I428444,I428452,I428469,I428500,I428517,I428534,I428565,I428596,I428613,I428668,I428694,I428702,I428719,I428736,I428762,I428793,I428801,I428818,I428844,I428852,I428892,I428928,I428945,I428971,I428979,I428996,I429027,I429044,I429061,I429092,I429123,I429140,I429195,I429221,I429229,I429246,I429263,I429289,I429320,I429328,I429345,I429371,I429379,I429419,I429455,I429472,I429498,I429506,I429523,I429554,I429571,I429588,I429619,I429650,I429667,I429722,I429748,I429756,I429773,I429790,I429816,I429847,I429855,I429872,I429898,I429906,I429946,I429982,I429999,I430025,I430033,I430050,I430081,I430098,I430115,I430146,I430177,I430194,I430249,I568286,I430275,I430283,I430300,I568295,I568283,I430317,I568280,I430343,I430374,I430382,I568277,I430399,I430425,I430433,I430473,I430509,I568298,I568289,I430526,I568292,I430552,I430560,I430577,I430608,I430625,I430642,I430673,I430704,I430721,I430776,I430802,I430810,I430827,I430844,I430870,I430901,I430909,I430926,I430952,I430960,I431000,I431036,I431053,I431079,I431087,I431104,I431135,I431152,I431169,I431200,I431231,I431248,I431303,I620247,I431329,I431337,I431354,I620229,I431371,I620235,I431397,I431292,I620232,I431428,I431436,I620241,I431453,I431479,I431487,I431295,I620253,I431527,I431286,I431277,I431563,I620244,I620238,I431580,I431606,I431614,I431631,I431280,I431662,I620250,I431679,I431696,I431289,I431727,I431274,I431758,I431775,I431283,I431830,I431856,I431864,I431881,I431898,I431924,I431819,I431955,I431963,I431980,I432006,I432014,I431822,I432054,I431813,I431804,I432090,I432107,I432133,I432141,I432158,I431807,I432189,I432206,I432223,I431816,I432254,I431801,I432285,I432302,I431810,I432357,I432383,I432391,I432408,I432425,I432451,I432482,I432490,I432507,I432533,I432541,I432581,I432617,I432634,I432660,I432668,I432685,I432716,I432733,I432750,I432781,I432812,I432829,I432884,I432910,I432918,I432935,I432952,I432978,I433009,I433017,I433034,I433060,I433068,I433108,I433144,I433161,I433187,I433195,I433212,I433243,I433260,I433277,I433308,I433339,I433356,I433411,I433437,I433445,I433462,I433479,I433505,I433400,I433536,I433544,I433561,I433587,I433595,I433403,I433635,I433394,I433385,I433671,I433688,I433714,I433722,I433739,I433388,I433770,I433787,I433804,I433397,I433835,I433382,I433866,I433883,I433391,I433938,I433964,I433972,I433989,I434006,I434032,I433927,I434063,I434071,I434088,I434114,I434122,I433930,I434162,I433921,I433912,I434198,I434215,I434241,I434249,I434266,I433915,I434297,I434314,I434331,I433924,I434362,I433909,I434393,I434410,I433918,I434465,I434491,I434499,I434516,I434533,I434559,I434454,I434590,I434598,I434615,I434641,I434649,I434457,I434689,I434448,I434439,I434725,I434742,I434768,I434776,I434793,I434442,I434824,I434841,I434858,I434451,I434889,I434436,I434920,I434937,I434445,I434992,I435018,I435026,I435043,I435060,I435086,I434981,I435117,I435125,I435142,I435168,I435176,I434984,I435216,I434975,I434966,I435252,I435269,I435295,I435303,I435320,I434969,I435351,I435368,I435385,I434978,I435416,I434963,I435447,I435464,I434972,I435519,I691848,I435545,I435553,I435570,I691845,I691854,I435587,I691833,I435613,I691836,I435644,I435652,I691851,I435669,I435695,I435703,I691857,I435743,I435779,I691839,I691860,I435796,I691842,I435822,I435830,I435847,I435878,I435895,I435912,I435943,I435974,I435991,I436046,I436072,I436080,I436097,I436114,I436140,I436171,I436179,I436196,I436222,I436230,I436270,I436306,I436323,I436349,I436357,I436374,I436405,I436422,I436439,I436470,I436501,I436518,I436573,I436599,I436607,I436624,I436641,I436667,I436698,I436706,I436723,I436749,I436757,I436797,I436833,I436850,I436876,I436884,I436901,I436932,I436949,I436966,I436997,I437028,I437045,I437100,I727548,I437126,I437134,I437151,I727545,I727554,I437168,I727533,I437194,I727536,I437225,I437233,I727551,I437250,I437276,I437284,I727557,I437324,I437360,I727539,I727560,I437377,I727542,I437403,I437411,I437428,I437459,I437476,I437493,I437524,I437555,I437572,I437627,I520289,I437653,I437661,I437678,I520304,I520286,I437695,I437721,I520295,I437752,I437760,I520313,I437777,I437803,I437811,I520310,I437851,I437887,I520307,I520298,I437904,I520292,I437930,I437938,I437955,I437986,I520301,I438003,I438020,I438051,I438082,I438099,I438154,I519643,I438180,I438188,I438205,I519658,I519640,I438222,I438248,I438143,I519649,I438279,I438287,I519667,I438304,I438330,I438338,I438146,I519664,I438378,I438137,I438128,I438414,I519661,I519652,I438431,I519646,I438457,I438465,I438482,I438131,I438513,I519655,I438530,I438547,I438140,I438578,I438125,I438609,I438626,I438134,I438681,I438707,I438715,I438732,I438749,I438775,I438806,I438814,I438831,I438857,I438865,I438905,I438941,I438958,I438984,I438992,I439009,I439040,I439057,I439074,I439105,I439136,I439153,I439208,I439234,I439242,I439259,I439276,I439302,I439333,I439341,I439358,I439384,I439392,I439432,I439468,I439485,I439511,I439519,I439536,I439567,I439584,I439601,I439632,I439663,I439680,I439735,I695418,I439761,I439769,I439786,I695415,I695424,I439803,I695403,I439829,I439724,I695406,I439860,I439868,I695421,I439885,I439911,I439919,I439727,I695427,I439959,I439718,I439709,I439995,I695409,I695430,I440012,I695412,I440038,I440046,I440063,I439712,I440094,I440111,I440128,I439721,I440159,I439706,I440190,I440207,I439715,I440262,I687776,I440288,I440296,I440313,I687770,I687788,I440330,I687773,I440356,I440251,I687794,I440387,I440395,I687779,I440412,I440438,I440446,I440254,I687791,I440486,I440245,I440236,I440522,I687782,I687797,I440539,I687785,I440565,I440573,I440590,I440239,I440621,I440638,I440655,I440248,I440686,I440233,I440717,I440734,I440242,I440789,I440815,I440823,I440840,I440857,I440883,I440914,I440922,I440939,I440965,I440973,I441013,I441049,I441066,I441092,I441100,I441117,I441148,I441165,I441182,I441213,I441244,I441261,I441316,I441342,I441350,I441367,I441384,I441410,I441305,I441441,I441449,I441466,I441492,I441500,I441308,I441540,I441299,I441290,I441576,I441593,I441619,I441627,I441644,I441293,I441675,I441692,I441709,I441302,I441740,I441287,I441771,I441788,I441296,I441843,I441869,I441877,I441894,I441911,I441937,I441968,I441976,I441993,I442019,I442027,I442067,I442103,I442120,I442146,I442154,I442171,I442202,I442219,I442236,I442267,I442298,I442315,I442370,I442396,I442404,I442421,I442438,I442464,I442359,I442495,I442503,I442520,I442546,I442554,I442362,I442594,I442353,I442344,I442630,I442647,I442673,I442681,I442698,I442347,I442729,I442746,I442763,I442356,I442794,I442341,I442825,I442842,I442350,I442897,I442923,I442931,I442948,I442965,I442991,I443022,I443030,I443047,I443073,I443081,I443121,I443157,I443174,I443200,I443208,I443225,I443256,I443273,I443290,I443321,I443352,I443369,I443424,I443450,I443458,I443475,I443492,I443518,I443549,I443557,I443574,I443600,I443608,I443648,I443684,I443701,I443727,I443735,I443752,I443783,I443800,I443817,I443848,I443879,I443896,I443951,I705533,I443977,I443985,I444002,I705530,I705539,I444019,I705518,I444045,I443940,I705521,I444076,I444084,I705536,I444101,I444127,I444135,I443943,I705542,I444175,I443934,I443925,I444211,I705524,I705545,I444228,I705527,I444254,I444262,I444279,I443928,I444310,I444327,I444344,I443937,I444375,I443922,I444406,I444423,I443931,I444478,I444504,I444512,I444529,I444546,I444572,I444603,I444611,I444628,I444654,I444662,I444702,I444738,I444755,I444781,I444789,I444806,I444837,I444854,I444871,I444902,I444933,I444950,I445005,I445031,I445039,I445056,I445073,I445099,I445130,I445138,I445155,I445181,I445189,I445229,I445265,I445282,I445308,I445316,I445333,I445364,I445381,I445398,I445429,I445460,I445477,I445532,I692443,I445558,I445566,I445583,I692440,I692449,I445600,I692428,I445626,I445521,I692431,I445657,I445665,I692446,I445682,I445708,I445716,I445524,I692452,I445756,I445515,I445506,I445792,I692434,I692455,I445809,I692437,I445835,I445843,I445860,I445509,I445891,I445908,I445925,I445518,I445956,I445503,I445987,I446004,I445512,I446059,I446085,I446093,I446110,I446127,I446153,I446048,I446184,I446192,I446209,I446235,I446243,I446051,I446283,I446042,I446033,I446319,I446336,I446362,I446370,I446387,I446036,I446418,I446435,I446452,I446045,I446483,I446030,I446514,I446531,I446039,I446586,I446612,I446620,I446637,I446654,I446680,I446711,I446719,I446736,I446762,I446770,I446810,I446846,I446863,I446889,I446897,I446914,I446945,I446962,I446979,I447010,I447041,I447058,I447113,I447139,I447147,I447164,I447181,I447207,I447238,I447246,I447263,I447289,I447297,I447337,I447373,I447390,I447416,I447424,I447441,I447472,I447489,I447506,I447537,I447568,I447585,I447640,I447666,I447674,I447691,I447708,I447734,I447765,I447773,I447790,I447816,I447824,I447864,I447900,I447917,I447943,I447951,I447968,I447999,I448016,I448033,I448064,I448095,I448112,I448167,I448193,I448201,I448218,I448235,I448261,I448156,I448292,I448300,I448317,I448343,I448351,I448159,I448391,I448150,I448141,I448427,I448444,I448470,I448478,I448495,I448144,I448526,I448543,I448560,I448153,I448591,I448138,I448622,I448639,I448147,I448694,I448720,I448728,I448745,I448762,I448788,I448819,I448827,I448844,I448870,I448878,I448918,I448954,I448971,I448997,I449005,I449022,I449053,I449070,I449087,I449118,I449149,I449166,I449221,I449247,I449255,I449272,I449289,I449315,I449346,I449354,I449371,I449397,I449405,I449445,I449481,I449498,I449524,I449532,I449549,I449580,I449597,I449614,I449645,I449676,I449693,I449748,I449774,I449782,I449799,I449816,I449842,I449737,I449873,I449881,I449898,I449924,I449932,I449740,I449972,I449731,I449722,I450008,I450025,I450051,I450059,I450076,I449725,I450107,I450124,I450141,I449734,I450172,I449719,I450203,I450220,I449728,I450275,I450301,I450309,I450326,I450343,I450369,I450400,I450408,I450425,I450451,I450459,I450499,I450535,I450552,I450578,I450586,I450603,I450634,I450651,I450668,I450699,I450730,I450747,I450802,I450828,I450836,I450853,I450870,I450896,I450927,I450935,I450952,I450978,I450986,I451026,I451062,I451079,I451105,I451113,I451130,I451161,I451178,I451195,I451226,I451257,I451274,I451329,I717433,I451355,I451363,I451380,I717430,I717439,I451397,I717418,I451423,I717421,I451454,I451462,I717436,I451479,I451505,I451513,I717442,I451553,I451589,I717424,I717445,I451606,I717427,I451632,I451640,I451657,I451688,I451705,I451722,I451753,I451784,I451801,I451856,I451882,I451890,I451907,I451924,I451950,I451981,I451989,I452006,I452032,I452040,I452080,I452116,I452133,I452159,I452167,I452184,I452215,I452232,I452249,I452280,I452311,I452328,I452383,I586723,I452409,I452417,I452434,I586705,I452451,I586711,I452477,I452372,I586708,I452508,I452516,I586717,I452533,I452559,I452567,I452375,I586729,I452607,I452366,I452357,I452643,I586720,I586714,I452660,I452686,I452694,I452711,I452360,I452742,I586726,I452759,I452776,I452369,I452807,I452354,I452838,I452855,I452363,I452910,I452936,I452944,I452961,I452978,I453004,I453035,I453043,I453060,I453086,I453094,I453134,I453170,I453187,I453213,I453221,I453238,I453269,I453286,I453303,I453334,I453365,I453382,I453437,I676925,I453463,I453471,I453488,I676907,I676910,I453505,I676922,I453531,I453426,I676931,I453562,I453570,I676916,I453587,I453613,I453621,I453429,I676928,I453661,I453420,I453411,I453697,I676919,I676913,I453714,I453740,I453748,I453765,I453414,I453796,I453813,I453830,I453423,I453861,I453408,I453892,I453909,I453417,I453964,I453990,I453998,I454015,I454032,I454058,I453953,I454089,I454097,I454114,I454140,I454148,I453956,I454188,I453947,I453938,I454224,I454241,I454267,I454275,I454292,I453941,I454323,I454340,I454357,I453950,I454388,I453935,I454419,I454436,I453944,I454491,I454517,I454525,I454542,I454559,I454585,I454616,I454624,I454641,I454667,I454675,I454715,I454751,I454768,I454794,I454802,I454819,I454850,I454867,I454884,I454915,I454946,I454963,I455018,I455044,I455052,I455069,I455086,I455112,I455143,I455151,I455168,I455194,I455202,I455242,I455278,I455295,I455321,I455329,I455346,I455377,I455394,I455411,I455442,I455473,I455490,I455545,I455571,I455579,I455596,I455613,I455639,I455534,I455670,I455678,I455695,I455721,I455729,I455537,I455769,I455528,I455519,I455805,I455822,I455848,I455856,I455873,I455522,I455904,I455921,I455938,I455531,I455969,I455516,I456000,I456017,I455525,I456072,I456098,I456106,I456123,I456140,I456166,I456197,I456205,I456222,I456248,I456256,I456296,I456332,I456349,I456375,I456383,I456400,I456431,I456448,I456465,I456496,I456527,I456544,I456599,I456625,I456633,I456650,I456667,I456693,I456588,I456724,I456732,I456749,I456775,I456783,I456591,I456823,I456582,I456573,I456859,I456876,I456902,I456910,I456927,I456576,I456958,I456975,I456992,I456585,I457023,I456570,I457054,I457071,I456579,I457126,I457152,I457160,I457177,I457194,I457220,I457251,I457259,I457276,I457302,I457310,I457350,I457386,I457403,I457429,I457437,I457454,I457485,I457502,I457519,I457550,I457581,I457598,I457653,I621981,I457679,I457687,I457704,I621963,I457721,I621969,I457747,I621966,I457778,I457786,I621975,I457803,I457829,I457837,I621987,I457877,I457913,I621978,I621972,I457930,I457956,I457964,I457981,I458012,I621984,I458029,I458046,I458077,I458108,I458125,I458180,I593081,I458206,I458214,I458231,I593063,I458248,I593069,I458274,I593066,I458305,I458313,I593075,I458330,I458356,I458364,I593087,I458404,I458440,I593078,I593072,I458457,I458483,I458491,I458508,I458539,I593084,I458556,I458573,I458604,I458635,I458652,I458707,I458733,I458741,I458758,I458775,I458801,I458832,I458840,I458857,I458883,I458891,I458931,I458967,I458984,I459010,I459018,I459035,I459066,I459083,I459100,I459131,I459162,I459179,I459234,I459260,I459268,I459285,I459302,I459328,I459223,I459359,I459367,I459384,I459410,I459418,I459226,I459458,I459217,I459208,I459494,I459511,I459537,I459545,I459562,I459211,I459593,I459610,I459627,I459220,I459658,I459205,I459689,I459706,I459214,I459761,I459787,I459795,I459812,I459829,I459855,I459886,I459894,I459911,I459937,I459945,I459985,I460021,I460038,I460064,I460072,I460089,I460120,I460137,I460154,I460185,I460216,I460233,I460288,I460314,I460322,I460339,I460356,I460382,I460413,I460421,I460438,I460464,I460472,I460512,I460548,I460565,I460591,I460599,I460616,I460647,I460664,I460681,I460712,I460743,I460760,I460815,I518997,I460841,I460849,I460866,I519012,I518994,I460883,I460909,I519003,I460940,I460948,I519021,I460965,I460991,I460999,I519018,I461039,I461075,I519015,I519006,I461092,I519000,I461118,I461126,I461143,I461174,I519009,I461191,I461208,I461239,I461270,I461287,I461342,I461368,I461376,I461393,I461410,I461436,I461331,I461467,I461475,I461492,I461518,I461526,I461334,I461566,I461325,I461316,I461602,I461619,I461645,I461653,I461670,I461319,I461701,I461718,I461735,I461328,I461766,I461313,I461797,I461814,I461322,I461869,I461895,I461903,I461920,I461937,I461963,I461858,I461994,I462002,I462019,I462045,I462053,I461861,I462093,I461852,I461843,I462129,I462146,I462172,I462180,I462197,I461846,I462228,I462245,I462262,I461855,I462293,I461840,I462324,I462341,I461849,I462396,I508661,I462422,I462430,I462447,I508676,I508658,I462464,I462490,I508667,I462521,I462529,I508685,I462546,I462572,I462580,I508682,I462620,I462656,I508679,I508670,I462673,I508664,I462699,I462707,I462724,I462755,I508673,I462772,I462789,I462820,I462851,I462868,I462923,I462949,I462957,I462974,I462991,I463017,I462912,I463048,I463056,I463073,I463099,I463107,I462915,I463147,I462906,I462897,I463183,I463200,I463226,I463234,I463251,I462900,I463282,I463299,I463316,I462909,I463347,I462894,I463378,I463395,I462903,I463450,I463476,I463484,I463501,I463518,I463544,I463439,I463575,I463583,I463600,I463626,I463634,I463442,I463674,I463433,I463424,I463710,I463727,I463753,I463761,I463778,I463427,I463809,I463826,I463843,I463436,I463874,I463421,I463905,I463922,I463430,I463977,I464003,I464011,I464028,I464045,I464071,I463966,I464102,I464110,I464127,I464153,I464161,I463969,I464201,I463960,I463951,I464237,I464254,I464280,I464288,I464305,I463954,I464336,I464353,I464370,I463963,I464401,I463948,I464432,I464449,I463957,I464504,I644721,I464530,I464538,I464555,I644727,I644709,I464572,I644718,I464598,I644724,I464629,I464637,I644712,I464654,I464680,I464688,I644730,I464728,I464764,I644715,I464781,I644733,I464807,I464815,I464832,I464863,I464880,I464897,I464928,I464959,I464976,I465031,I465057,I465065,I465082,I465099,I465125,I465156,I465164,I465181,I465207,I465215,I465255,I465291,I465308,I465334,I465342,I465359,I465390,I465407,I465424,I465455,I465486,I465503,I465558,I465584,I465592,I465609,I465626,I465652,I465683,I465691,I465708,I465734,I465742,I465782,I465818,I465835,I465861,I465869,I465886,I465917,I465934,I465951,I465982,I466013,I466030,I466085,I466111,I466119,I466136,I466153,I466179,I466074,I466210,I466218,I466235,I466261,I466269,I466077,I466309,I466068,I466059,I466345,I466362,I466388,I466396,I466413,I466062,I466444,I466461,I466478,I466071,I466509,I466056,I466540,I466557,I466065,I466612,I707913,I466638,I466646,I466663,I707910,I707919,I466680,I707898,I466706,I707901,I466737,I466745,I707916,I466762,I466788,I466796,I707922,I466836,I466872,I707904,I707925,I466889,I707907,I466915,I466923,I466940,I466971,I466988,I467005,I467036,I467067,I467084,I467139,I467165,I467173,I467190,I467207,I467233,I467128,I467264,I467272,I467289,I467315,I467323,I467131,I467363,I467122,I467113,I467399,I467416,I467442,I467450,I467467,I467116,I467498,I467515,I467532,I467125,I467563,I467110,I467594,I467611,I467119,I467666,I484759,I467692,I467700,I467717,I484774,I484756,I467734,I467760,I467655,I484765,I467791,I467799,I484783,I467816,I467842,I467850,I467658,I484780,I467890,I467649,I467640,I467926,I484777,I484768,I467943,I484762,I467969,I467977,I467994,I467643,I468025,I484771,I468042,I468059,I467652,I468090,I467637,I468121,I468138,I467646,I468193,I468219,I468227,I468244,I468261,I468287,I468318,I468326,I468343,I468369,I468377,I468417,I468453,I468470,I468496,I468504,I468521,I468552,I468569,I468586,I468617,I468648,I468665,I468720,I468746,I468754,I468771,I468788,I468814,I468845,I468853,I468870,I468896,I468904,I468944,I468980,I468997,I469023,I469031,I469048,I469079,I469096,I469113,I469144,I469175,I469192,I469247,I690063,I469273,I469281,I469298,I690060,I690069,I469315,I690048,I469341,I690051,I469372,I469380,I690066,I469397,I469423,I469431,I690072,I469471,I469507,I690054,I690075,I469524,I690057,I469550,I469558,I469575,I469606,I469623,I469640,I469671,I469702,I469719,I469774,I469800,I469808,I469825,I469842,I469868,I469899,I469907,I469924,I469950,I469958,I469998,I470034,I470051,I470077,I470085,I470102,I470133,I470150,I470167,I470198,I470229,I470246,I470301,I470327,I470335,I470352,I470369,I470395,I470426,I470434,I470451,I470477,I470485,I470525,I470561,I470578,I470604,I470612,I470629,I470660,I470677,I470694,I470725,I470756,I470773,I470828,I669989,I470854,I470862,I470879,I669971,I669974,I470896,I669986,I470922,I669995,I470953,I470961,I669980,I470978,I471004,I471012,I669992,I471052,I471088,I669983,I669977,I471105,I471131,I471139,I471156,I471187,I471204,I471221,I471252,I471283,I471300,I471355,I635275,I471381,I471389,I471406,I635257,I471423,I635263,I471449,I635260,I471480,I471488,I635269,I471505,I471531,I471539,I635281,I471579,I471615,I635272,I635266,I471632,I471658,I471666,I471683,I471714,I635278,I471731,I471748,I471779,I471810,I471827,I471882,I471908,I471916,I471933,I471950,I471976,I472007,I472015,I472032,I472058,I472066,I472106,I472142,I472159,I472185,I472193,I472210,I472241,I472258,I472275,I472306,I472337,I472354,I472409,I472435,I472443,I472460,I472477,I472503,I472534,I472542,I472559,I472585,I472593,I472633,I472669,I472686,I472712,I472720,I472737,I472768,I472785,I472802,I472833,I472864,I472881,I472936,I472962,I472970,I472987,I473004,I473030,I473061,I473069,I473086,I473112,I473120,I473160,I473196,I473213,I473239,I473247,I473264,I473295,I473312,I473329,I473360,I473391,I473408,I473463,I477653,I473489,I473497,I473514,I477668,I477650,I473531,I473557,I477659,I473588,I473596,I477677,I473613,I473639,I473647,I477674,I473687,I473723,I477671,I477662,I473740,I477656,I473766,I473774,I473791,I473822,I477665,I473839,I473856,I473887,I473918,I473935,I473990,I474016,I474024,I474041,I474058,I474084,I473979,I474115,I474123,I474140,I474166,I474174,I473982,I474214,I473973,I473964,I474250,I474267,I474293,I474301,I474318,I473967,I474349,I474366,I474383,I473976,I474414,I473961,I474445,I474462,I473970,I474517,I474543,I474551,I474568,I474585,I474611,I474642,I474650,I474667,I474693,I474701,I474741,I474777,I474794,I474820,I474828,I474845,I474876,I474893,I474910,I474941,I474972,I474989,I475044,I624871,I475070,I475078,I475095,I624853,I475112,I624859,I475138,I475033,I624856,I475169,I475177,I624865,I475194,I475220,I475228,I475036,I624877,I475268,I475027,I475018,I475304,I624868,I624862,I475321,I475347,I475355,I475372,I475021,I475403,I624874,I475420,I475437,I475030,I475468,I475015,I475499,I475516,I475024,I475571,I475597,I475605,I475622,I475639,I475665,I475560,I475696,I475704,I475721,I475747,I475755,I475563,I475795,I475554,I475545,I475831,I475848,I475874,I475882,I475899,I475548,I475930,I475947,I475964,I475557,I475995,I475542,I476026,I476043,I475551,I476098,I476124,I476132,I476149,I476166,I476192,I476223,I476231,I476248,I476274,I476282,I476322,I476358,I476375,I476401,I476409,I476426,I476457,I476474,I476491,I476522,I476553,I476570,I476625,I476651,I476659,I476676,I476693,I476719,I476750,I476758,I476775,I476801,I476809,I476849,I476885,I476902,I476928,I476936,I476953,I476984,I477001,I477018,I477049,I477080,I477097,I477152,I477178,I477186,I477203,I477220,I477246,I477277,I477285,I477302,I477328,I477336,I477376,I477412,I477429,I477455,I477463,I477480,I477511,I477528,I477545,I477576,I477607,I477624,I477685,I584411,I477711,I584393,I477728,I477736,I477753,I584402,I477770,I584414,I477787,I584396,I477804,I584405,I477821,I477852,I477869,I477900,I477917,I584417,I477934,I477965,I478005,I478013,I478030,I478047,I478064,I478095,I584399,I478112,I584408,I478129,I478155,I478177,I478194,I478225,I478270,I478331,I478357,I478374,I478382,I478399,I478416,I478433,I478450,I478467,I478498,I478515,I478546,I478563,I478580,I478611,I478651,I478659,I478676,I478693,I478710,I478741,I478758,I478775,I478801,I478823,I478840,I478871,I478916,I478977,I479003,I479020,I479028,I479045,I479062,I479079,I479096,I479113,I479144,I479161,I479192,I479209,I479226,I479257,I479297,I479305,I479322,I479339,I479356,I479387,I479404,I479421,I479447,I479469,I479486,I479517,I479562,I479623,I479649,I479666,I479674,I479691,I479708,I479725,I479742,I479759,I479790,I479807,I479838,I479855,I479872,I479903,I479943,I479951,I479968,I479985,I480002,I480033,I480050,I480067,I480093,I480115,I480132,I480163,I480208,I480269,I480295,I480312,I480320,I480337,I480354,I480371,I480388,I480405,I480255,I480436,I480453,I480258,I480484,I480501,I480518,I480234,I480549,I480246,I480589,I480597,I480614,I480631,I480648,I480261,I480679,I480696,I480713,I480739,I480249,I480761,I480778,I480243,I480809,I480237,I480240,I480854,I480252,I480915,I480941,I480958,I480966,I480983,I481000,I481017,I481034,I481051,I481082,I481099,I481130,I481147,I481164,I481195,I481235,I481243,I481260,I481277,I481294,I481325,I481342,I481359,I481385,I481407,I481424,I481455,I481500,I481561,I629495,I481587,I629477,I481604,I481612,I481629,I629486,I481646,I629498,I481663,I629480,I481680,I629489,I481697,I481547,I481728,I481745,I481550,I481776,I481793,I629501,I481810,I481526,I481841,I481538,I481881,I481889,I481906,I481923,I481940,I481553,I481971,I629483,I481988,I629492,I482005,I482031,I481541,I482053,I482070,I481535,I482101,I481529,I481532,I482146,I481544,I482207,I482233,I482250,I482258,I482275,I482292,I482309,I482326,I482343,I482374,I482391,I482422,I482439,I482456,I482487,I482527,I482535,I482552,I482569,I482586,I482617,I482634,I482651,I482677,I482699,I482716,I482747,I482792,I482853,I482879,I482896,I482904,I482921,I482938,I482955,I482972,I482989,I483020,I483037,I483068,I483085,I483102,I483133,I483173,I483181,I483198,I483215,I483232,I483263,I483280,I483297,I483323,I483345,I483362,I483393,I483438,I483499,I654519,I483525,I654525,I483542,I483550,I483567,I654522,I483584,I654501,I483601,I654504,I483618,I654510,I483635,I483666,I483683,I483714,I483731,I483748,I483779,I483819,I483827,I483844,I483861,I654513,I483878,I483909,I483926,I654507,I483943,I654516,I483969,I483991,I484008,I484039,I484084,I484145,I484171,I484188,I484196,I484213,I484230,I484247,I484264,I484281,I484312,I484329,I484360,I484377,I484394,I484425,I484465,I484473,I484490,I484507,I484524,I484555,I484572,I484589,I484615,I484637,I484654,I484685,I484730,I484791,I567155,I484817,I567158,I484834,I484842,I484859,I484876,I567167,I484893,I567176,I484910,I567164,I484927,I484958,I484975,I485006,I485023,I567170,I485040,I485071,I485111,I485119,I485136,I485153,I567161,I485170,I485201,I567173,I485218,I485235,I485261,I485283,I485300,I485331,I485376,I485437,I485463,I485480,I485488,I485505,I485522,I485539,I485556,I485573,I485604,I485621,I485652,I485669,I485686,I485717,I485757,I485765,I485782,I485799,I485816,I485847,I485864,I485881,I485907,I485929,I485946,I485977,I486022,I486083,I486109,I486126,I486134,I486151,I486168,I486185,I486202,I486219,I486250,I486267,I486298,I486315,I486332,I486363,I486403,I486411,I486428,I486445,I486462,I486493,I486510,I486527,I486553,I486575,I486592,I486623,I486668,I486729,I486755,I486772,I486780,I486797,I486814,I486831,I486848,I486865,I486896,I486913,I486944,I486961,I486978,I487009,I487049,I487057,I487074,I487091,I487108,I487139,I487156,I487173,I487199,I487221,I487238,I487269,I487314,I487375,I487401,I487418,I487426,I487443,I487460,I487477,I487494,I487511,I487361,I487542,I487559,I487364,I487590,I487607,I487624,I487340,I487655,I487352,I487695,I487703,I487720,I487737,I487754,I487367,I487785,I487802,I487819,I487845,I487355,I487867,I487884,I487349,I487915,I487343,I487346,I487960,I487358,I488021,I488047,I488064,I488072,I488089,I488106,I488123,I488140,I488157,I488188,I488205,I488236,I488253,I488270,I488301,I488341,I488349,I488366,I488383,I488400,I488431,I488448,I488465,I488491,I488513,I488530,I488561,I488606,I488667,I601173,I488693,I601155,I488710,I488718,I488735,I601164,I488752,I601176,I488769,I601158,I488786,I601167,I488803,I488653,I488834,I488851,I488656,I488882,I488899,I601179,I488916,I488632,I488947,I488644,I488987,I488995,I489012,I489029,I489046,I488659,I489077,I601161,I489094,I601170,I489111,I489137,I488647,I489159,I489176,I488641,I489207,I488635,I488638,I489252,I488650,I489313,I489339,I489356,I489364,I489381,I489398,I489415,I489432,I489449,I489480,I489497,I489528,I489545,I489562,I489593,I489633,I489641,I489658,I489675,I489692,I489723,I489740,I489757,I489783,I489805,I489822,I489853,I489898,I489959,I649079,I489985,I649085,I490002,I490010,I490027,I649082,I490044,I649061,I490061,I649064,I490078,I649070,I490095,I490126,I490143,I490174,I490191,I490208,I490239,I490279,I490287,I490304,I490321,I649073,I490338,I490369,I490386,I649067,I490403,I649076,I490429,I490451,I490468,I490499,I490544,I490605,I490631,I490648,I490656,I490673,I490690,I490707,I490724,I490741,I490591,I490772,I490789,I490594,I490820,I490837,I490854,I490570,I490885,I490582,I490925,I490933,I490950,I490967,I490984,I490597,I491015,I491032,I491049,I491075,I490585,I491097,I491114,I490579,I491145,I490573,I490576,I491190,I490588,I491251,I491277,I491294,I491302,I491319,I491336,I491353,I491370,I491387,I491237,I491418,I491435,I491240,I491466,I491483,I491500,I491216,I491531,I491228,I491571,I491579,I491596,I491613,I491630,I491243,I491661,I491678,I491695,I491721,I491231,I491743,I491760,I491225,I491791,I491219,I491222,I491836,I491234,I491897,I697188,I491923,I697212,I491940,I491948,I491965,I697194,I491982,I697203,I491999,I492016,I697209,I492033,I492064,I492081,I492112,I492129,I697206,I492146,I492177,I492217,I492225,I492242,I492259,I697200,I492276,I492307,I697191,I492324,I697215,I492341,I697197,I492367,I492389,I492406,I492437,I492482,I492543,I492569,I492586,I492594,I492611,I492628,I492645,I492662,I492679,I492710,I492727,I492758,I492775,I492792,I492823,I492863,I492871,I492888,I492905,I492922,I492953,I492970,I492987,I493013,I493035,I493052,I493083,I493128,I493189,I635853,I493215,I635835,I493232,I493240,I493257,I635844,I493274,I635856,I493291,I635838,I493308,I635847,I493325,I493356,I493373,I493404,I493421,I635859,I493438,I493469,I493509,I493517,I493534,I493551,I493568,I493599,I635841,I493616,I635850,I493633,I493659,I493681,I493698,I493729,I493774,I493835,I613311,I493861,I613293,I493878,I493886,I493903,I613302,I493920,I613314,I493937,I613296,I493954,I613305,I493971,I493821,I494002,I494019,I493824,I494050,I494067,I613317,I494084,I493800,I494115,I493812,I494155,I494163,I494180,I494197,I494214,I493827,I494245,I613299,I494262,I613308,I494279,I494305,I493815,I494327,I494344,I493809,I494375,I493803,I493806,I494420,I493818,I494481,I494507,I494524,I494532,I494549,I494566,I494583,I494600,I494617,I494648,I494665,I494696,I494713,I494730,I494761,I494801,I494809,I494826,I494843,I494860,I494891,I494908,I494925,I494951,I494973,I494990,I495021,I495066,I495127,I495153,I495170,I495178,I495195,I495212,I495229,I495246,I495263,I495113,I495294,I495311,I495116,I495342,I495359,I495376,I495092,I495407,I495104,I495447,I495455,I495472,I495489,I495506,I495119,I495537,I495554,I495571,I495597,I495107,I495619,I495636,I495101,I495667,I495095,I495098,I495712,I495110,I495773,I495799,I495816,I495824,I495841,I495858,I495875,I495892,I495909,I495759,I495940,I495957,I495762,I495988,I496005,I496022,I495738,I496053,I495750,I496093,I496101,I496118,I496135,I496152,I495765,I496183,I496200,I496217,I496243,I495753,I496265,I496282,I495747,I496313,I495741,I495744,I496358,I495756,I496419,I496445,I496462,I496470,I496487,I496504,I496521,I496538,I496555,I496586,I496603,I496634,I496651,I496668,I496699,I496739,I496747,I496764,I496781,I496798,I496829,I496846,I496863,I496889,I496911,I496928,I496959,I497004,I497065,I497091,I497108,I497116,I497133,I497150,I497167,I497184,I497201,I497232,I497249,I497280,I497297,I497314,I497345,I497385,I497393,I497410,I497427,I497444,I497475,I497492,I497509,I497535,I497557,I497574,I497605,I497650,I497711,I497737,I497754,I497762,I497779,I497796,I497813,I497830,I497847,I497878,I497895,I497926,I497943,I497960,I497991,I498031,I498039,I498056,I498073,I498090,I498121,I498138,I498155,I498181,I498203,I498220,I498251,I498296,I498357,I640919,I498383,I640925,I498400,I498408,I498425,I640922,I498442,I640901,I498459,I640904,I498476,I640910,I498493,I498343,I498524,I498541,I498346,I498572,I498589,I498606,I498322,I498637,I498334,I498677,I498685,I498702,I498719,I640913,I498736,I498349,I498767,I498784,I640907,I498801,I640916,I498827,I498337,I498849,I498866,I498331,I498897,I498325,I498328,I498942,I498340,I499003,I499029,I499046,I499054,I499071,I499088,I499105,I499122,I499139,I499170,I499187,I499218,I499235,I499252,I499283,I499323,I499331,I499348,I499365,I499382,I499413,I499430,I499447,I499473,I499495,I499512,I499543,I499588,I499649,I499675,I499692,I499700,I499717,I499734,I499751,I499768,I499785,I499816,I499833,I499864,I499881,I499898,I499929,I499969,I499977,I499994,I500011,I500028,I500059,I500076,I500093,I500119,I500141,I500158,I500189,I500234,I500295,I710278,I500321,I710302,I500338,I500346,I500363,I710284,I500380,I710293,I500397,I500414,I710299,I500431,I500462,I500479,I500510,I500527,I710296,I500544,I500575,I500615,I500623,I500640,I500657,I710290,I500674,I500705,I710281,I500722,I710305,I500739,I710287,I500765,I500787,I500804,I500835,I500880,I500941,I600595,I500967,I600577,I500984,I500992,I501009,I600586,I501026,I600598,I501043,I600580,I501060,I600589,I501077,I501108,I501125,I501156,I501173,I600601,I501190,I501221,I501261,I501269,I501286,I501303,I501320,I501351,I600583,I501368,I600592,I501385,I501411,I501433,I501450,I501481,I501526,I501587,I501613,I501630,I501638,I501655,I501672,I501689,I501706,I501723,I501754,I501771,I501802,I501819,I501836,I501867,I501907,I501915,I501932,I501949,I501966,I501997,I502014,I502031,I502057,I502079,I502096,I502127,I502172,I502233,I502259,I502276,I502284,I502301,I502318,I502335,I502352,I502369,I502400,I502417,I502448,I502465,I502482,I502513,I502553,I502561,I502578,I502595,I502612,I502643,I502660,I502677,I502703,I502725,I502742,I502773,I502818,I502879,I502905,I502922,I502930,I502947,I502964,I502981,I502998,I503015,I502865,I503046,I503063,I502868,I503094,I503111,I503128,I502844,I503159,I502856,I503199,I503207,I503224,I503241,I503258,I502871,I503289,I503306,I503323,I503349,I502859,I503371,I503388,I502853,I503419,I502847,I502850,I503464,I502862,I503525,I545837,I503551,I545840,I503568,I503576,I503593,I503610,I545849,I503627,I545858,I503644,I545846,I503661,I503692,I503709,I503740,I503757,I545852,I503774,I503805,I503845,I503853,I503870,I503887,I545843,I503904,I503935,I545855,I503952,I503969,I503995,I504017,I504034,I504065,I504110,I504171,I504197,I504214,I504222,I504239,I504256,I504273,I504290,I504307,I504157,I504338,I504355,I504160,I504386,I504403,I504420,I504136,I504451,I504148,I504491,I504499,I504516,I504533,I504550,I504163,I504581,I504598,I504615,I504641,I504151,I504663,I504680,I504145,I504711,I504139,I504142,I504756,I504154,I504817,I504843,I504860,I504868,I504885,I504902,I504919,I504936,I504953,I504984,I505001,I505032,I505049,I505066,I505097,I505137,I505145,I505162,I505179,I505196,I505227,I505244,I505261,I505287,I505309,I505326,I505357,I505402,I505463,I505489,I505506,I505514,I505531,I505548,I505565,I505582,I505599,I505449,I505630,I505647,I505452,I505678,I505695,I505712,I505428,I505743,I505440,I505783,I505791,I505808,I505825,I505842,I505455,I505873,I505890,I505907,I505933,I505443,I505955,I505972,I505437,I506003,I505431,I505434,I506048,I505446,I506109,I506135,I506152,I506160,I506177,I506194,I506211,I506228,I506245,I506095,I506276,I506293,I506098,I506324,I506341,I506358,I506074,I506389,I506086,I506429,I506437,I506454,I506471,I506488,I506101,I506519,I506536,I506553,I506579,I506089,I506601,I506618,I506083,I506649,I506077,I506080,I506694,I506092,I506755,I694808,I506781,I694832,I506798,I506806,I506823,I694814,I506840,I694823,I506857,I506874,I694829,I506891,I506922,I506939,I506970,I506987,I694826,I507004,I507035,I507075,I507083,I507100,I507117,I694820,I507134,I507165,I694811,I507182,I694835,I507199,I694817,I507225,I507247,I507264,I507295,I507340,I507401,I507427,I507444,I507452,I507469,I507486,I507503,I507520,I507537,I507568,I507585,I507616,I507633,I507650,I507681,I507721,I507729,I507746,I507763,I507780,I507811,I507828,I507845,I507871,I507893,I507910,I507941,I507986,I508047,I571695,I508073,I571677,I508090,I508098,I508115,I571686,I508132,I571698,I508149,I571680,I508166,I571689,I508183,I508033,I508214,I508231,I508036,I508262,I508279,I571701,I508296,I508012,I508327,I508024,I508367,I508375,I508392,I508409,I508426,I508039,I508457,I571683,I508474,I571692,I508491,I508517,I508027,I508539,I508556,I508021,I508587,I508015,I508018,I508632,I508030,I508693,I508719,I508736,I508744,I508761,I508778,I508795,I508812,I508829,I508860,I508877,I508908,I508925,I508942,I508973,I509013,I509021,I509038,I509055,I509072,I509103,I509120,I509137,I509163,I509185,I509202,I509233,I509278,I509339,I571117,I509365,I571099,I509382,I509390,I509407,I571108,I509424,I571120,I509441,I571102,I509458,I571111,I509475,I509506,I509523,I509554,I509571,I571123,I509588,I509619,I509659,I509667,I509684,I509701,I509718,I509749,I571105,I509766,I571114,I509783,I509809,I509831,I509848,I509879,I509924,I509985,I715633,I510011,I715657,I510028,I510036,I510053,I715639,I510070,I715648,I510087,I510104,I715654,I510121,I509971,I510152,I510169,I509974,I510200,I510217,I715651,I510234,I509950,I510265,I509962,I510305,I510313,I510330,I510347,I715645,I510364,I509977,I510395,I715636,I510412,I715660,I510429,I715642,I510455,I509965,I510477,I510494,I509959,I510525,I509953,I509956,I510570,I509968,I510631,I510657,I510674,I510682,I510699,I510716,I510733,I510750,I510767,I510798,I510815,I510846,I510863,I510880,I510911,I510951,I510959,I510976,I510993,I511010,I511041,I511058,I511075,I511101,I511123,I511140,I511171,I511216,I511277,I511303,I511320,I511328,I511345,I511362,I511379,I511396,I511413,I511263,I511444,I511461,I511266,I511492,I511509,I511526,I511242,I511557,I511254,I511597,I511605,I511622,I511639,I511656,I511269,I511687,I511704,I511721,I511747,I511257,I511769,I511786,I511251,I511817,I511245,I511248,I511862,I511260,I511923,I511949,I511966,I511974,I511991,I512008,I512025,I512042,I512059,I511909,I512090,I512107,I511912,I512138,I512155,I512172,I511888,I512203,I511900,I512243,I512251,I512268,I512285,I512302,I511915,I512333,I512350,I512367,I512393,I511903,I512415,I512432,I511897,I512463,I511891,I511894,I512508,I511906,I512569,I512595,I512612,I512620,I512637,I512654,I512671,I512688,I512705,I512736,I512753,I512784,I512801,I512818,I512849,I512889,I512897,I512914,I512931,I512948,I512979,I512996,I513013,I513039,I513061,I513078,I513109,I513154,I513215,I513241,I513258,I513266,I513283,I513300,I513317,I513334,I513351,I513382,I513399,I513430,I513447,I513464,I513495,I513535,I513543,I513560,I513577,I513594,I513625,I513642,I513659,I513685,I513707,I513724,I513755,I513800,I513861,I513887,I513904,I513912,I513929,I513946,I513963,I513980,I513997,I513847,I514028,I514045,I513850,I514076,I514093,I514110,I513826,I514141,I513838,I514181,I514189,I514206,I514223,I514240,I513853,I514271,I514288,I514305,I514331,I513841,I514353,I514370,I513835,I514401,I513829,I513832,I514446,I513844,I514507,I514533,I514550,I514558,I514575,I514592,I514609,I514626,I514643,I514674,I514691,I514722,I514739,I514756,I514787,I514827,I514835,I514852,I514869,I514886,I514917,I514934,I514951,I514977,I514999,I515016,I515047,I515092,I515153,I691238,I515179,I691262,I515196,I515204,I515221,I691244,I515238,I691253,I515255,I515272,I691259,I515289,I515320,I515337,I515368,I515385,I691256,I515402,I515433,I515473,I515481,I515498,I515515,I691250,I515532,I515563,I691241,I515580,I691265,I515597,I691247,I515623,I515645,I515662,I515693,I515738,I515799,I515825,I515842,I515850,I515867,I515884,I515901,I515918,I515935,I515966,I515983,I516014,I516031,I516048,I516079,I516119,I516127,I516144,I516161,I516178,I516209,I516226,I516243,I516269,I516291,I516308,I516339,I516384,I516445,I516471,I516488,I516496,I516513,I516530,I516547,I516564,I516581,I516612,I516629,I516660,I516677,I516694,I516725,I516765,I516773,I516790,I516807,I516824,I516855,I516872,I516889,I516915,I516937,I516954,I516985,I517030,I517091,I517117,I517134,I517142,I517159,I517176,I517193,I517210,I517227,I517258,I517275,I517306,I517323,I517340,I517371,I517411,I517419,I517436,I517453,I517470,I517501,I517518,I517535,I517561,I517583,I517600,I517631,I517676,I517737,I517763,I517780,I517788,I517805,I517822,I517839,I517856,I517873,I517904,I517921,I517952,I517969,I517986,I518017,I518057,I518065,I518082,I518099,I518116,I518147,I518164,I518181,I518207,I518229,I518246,I518277,I518322,I518383,I518409,I518426,I518434,I518451,I518468,I518485,I518502,I518519,I518369,I518550,I518567,I518372,I518598,I518615,I518632,I518348,I518663,I518360,I518703,I518711,I518728,I518745,I518762,I518375,I518793,I518810,I518827,I518853,I518363,I518875,I518892,I518357,I518923,I518351,I518354,I518968,I518366,I519029,I519055,I519072,I519080,I519097,I519114,I519131,I519148,I519165,I519196,I519213,I519244,I519261,I519278,I519309,I519349,I519357,I519374,I519391,I519408,I519439,I519456,I519473,I519499,I519521,I519538,I519569,I519614,I519675,I519701,I519718,I519726,I519743,I519760,I519777,I519794,I519811,I519842,I519859,I519890,I519907,I519924,I519955,I519995,I520003,I520020,I520037,I520054,I520085,I520102,I520119,I520145,I520167,I520184,I520215,I520260,I520321,I520347,I520364,I520372,I520389,I520406,I520423,I520440,I520457,I520488,I520505,I520536,I520553,I520570,I520601,I520641,I520649,I520666,I520683,I520700,I520731,I520748,I520765,I520791,I520813,I520830,I520861,I520906,I520967,I520993,I521010,I521018,I521035,I521052,I521069,I521086,I521103,I521134,I521151,I521182,I521199,I521216,I521247,I521287,I521295,I521312,I521329,I521346,I521377,I521394,I521411,I521437,I521459,I521476,I521507,I521552,I521613,I521639,I521656,I521664,I521681,I521698,I521715,I521732,I521749,I521780,I521797,I521828,I521845,I521862,I521893,I521933,I521941,I521958,I521975,I521992,I522023,I522040,I522057,I522083,I522105,I522122,I522153,I522198,I522259,I651799,I522285,I651805,I522302,I522310,I522327,I651802,I522344,I651781,I522361,I651784,I522378,I651790,I522395,I522245,I522426,I522443,I522248,I522474,I522491,I522508,I522224,I522539,I522236,I522579,I522587,I522604,I522621,I651793,I522638,I522251,I522669,I522686,I651787,I522703,I651796,I522729,I522239,I522751,I522768,I522233,I522799,I522227,I522230,I522844,I522242,I522905,I522931,I522948,I522956,I522973,I522990,I523007,I523024,I523041,I522891,I523072,I523089,I522894,I523120,I523137,I523154,I522870,I523185,I522882,I523225,I523233,I523250,I523267,I523284,I522897,I523315,I523332,I523349,I523375,I522885,I523397,I523414,I522879,I523445,I522873,I522876,I523490,I522888,I523551,I523577,I523594,I523602,I523619,I523636,I523653,I523670,I523687,I523718,I523735,I523766,I523783,I523800,I523831,I523871,I523879,I523896,I523913,I523930,I523961,I523978,I523995,I524021,I524043,I524060,I524091,I524136,I524197,I524223,I524240,I524248,I524265,I524282,I524299,I524316,I524333,I524183,I524364,I524381,I524186,I524412,I524429,I524446,I524162,I524477,I524174,I524517,I524525,I524542,I524559,I524576,I524189,I524607,I524624,I524641,I524667,I524177,I524689,I524706,I524171,I524737,I524165,I524168,I524782,I524180,I524843,I524869,I524886,I524894,I524911,I524928,I524945,I524962,I524979,I525010,I525027,I525058,I525075,I525092,I525123,I525163,I525171,I525188,I525205,I525222,I525253,I525270,I525287,I525313,I525335,I525352,I525383,I525428,I525489,I525515,I525532,I525540,I525557,I525574,I525591,I525608,I525625,I525656,I525673,I525704,I525721,I525738,I525769,I525809,I525817,I525834,I525851,I525868,I525899,I525916,I525933,I525959,I525981,I525998,I526029,I526074,I526135,I526161,I526178,I526186,I526203,I526220,I526237,I526254,I526271,I526302,I526319,I526350,I526367,I526384,I526415,I526455,I526463,I526480,I526497,I526514,I526545,I526562,I526579,I526605,I526627,I526644,I526675,I526720,I526781,I526807,I526824,I526832,I526849,I526866,I526883,I526900,I526917,I526767,I526948,I526965,I526770,I526996,I527013,I527030,I526746,I527061,I526758,I527101,I527109,I527126,I527143,I527160,I526773,I527191,I527208,I527225,I527251,I526761,I527273,I527290,I526755,I527321,I526749,I526752,I527366,I526764,I527427,I527453,I527470,I527478,I527495,I527512,I527529,I527546,I527563,I527594,I527611,I527642,I527659,I527676,I527707,I527747,I527755,I527772,I527789,I527806,I527837,I527854,I527871,I527897,I527919,I527936,I527967,I528012,I528073,I528099,I528116,I528124,I528141,I528158,I528175,I528192,I528209,I528059,I528240,I528257,I528062,I528288,I528305,I528322,I528038,I528353,I528050,I528393,I528401,I528418,I528435,I528452,I528065,I528483,I528500,I528517,I528543,I528053,I528565,I528582,I528047,I528613,I528041,I528044,I528658,I528056,I528719,I528745,I528762,I528770,I528787,I528804,I528821,I528838,I528855,I528886,I528903,I528934,I528951,I528968,I528999,I529039,I529047,I529064,I529081,I529098,I529129,I529146,I529163,I529189,I529211,I529228,I529259,I529304,I529365,I529391,I529408,I529416,I529433,I529450,I529467,I529484,I529501,I529532,I529549,I529580,I529597,I529614,I529645,I529685,I529693,I529710,I529727,I529744,I529775,I529792,I529809,I529835,I529857,I529874,I529905,I529950,I530011,I530037,I530054,I530062,I530079,I530096,I530113,I530130,I530147,I530178,I530195,I530226,I530243,I530260,I530291,I530331,I530339,I530356,I530373,I530390,I530421,I530438,I530455,I530481,I530503,I530520,I530551,I530596,I530657,I530683,I530700,I530708,I530725,I530742,I530759,I530776,I530793,I530824,I530841,I530872,I530889,I530906,I530937,I530977,I530985,I531002,I531019,I531036,I531067,I531084,I531101,I531127,I531149,I531166,I531197,I531242,I531303,I544154,I531329,I544157,I531346,I531354,I531371,I531388,I544166,I531405,I544175,I531422,I544163,I531439,I531470,I531487,I531518,I531535,I544169,I531552,I531583,I531623,I531631,I531648,I531665,I544160,I531682,I531713,I544172,I531730,I531747,I531773,I531795,I531812,I531843,I531888,I531949,I647991,I531975,I647997,I531992,I532000,I532017,I647994,I532034,I647973,I532051,I647976,I532068,I647982,I532085,I532116,I532133,I532164,I532181,I532198,I532229,I532269,I532277,I532294,I532311,I647985,I532328,I532359,I532376,I647979,I532393,I647988,I532419,I532441,I532458,I532489,I532534,I532595,I716228,I532621,I716252,I532638,I532646,I532663,I716234,I532680,I716243,I532697,I532714,I716249,I532731,I532762,I532779,I532810,I532827,I716246,I532844,I532875,I532915,I532923,I532940,I532957,I716240,I532974,I533005,I716231,I533022,I716255,I533039,I716237,I533065,I533087,I533104,I533135,I533180,I533241,I533267,I533284,I533292,I533309,I533326,I533343,I533360,I533377,I533227,I533408,I533425,I533230,I533456,I533473,I533490,I533206,I533521,I533218,I533561,I533569,I533586,I533603,I533620,I533233,I533651,I533668,I533685,I533711,I533221,I533733,I533750,I533215,I533781,I533209,I533212,I533826,I533224,I533887,I533913,I533930,I533938,I533955,I533972,I533989,I534006,I534023,I533873,I534054,I534071,I533876,I534102,I534119,I534136,I533852,I534167,I533864,I534207,I534215,I534232,I534249,I534266,I533879,I534297,I534314,I534331,I534357,I533867,I534379,I534396,I533861,I534427,I533855,I533858,I534472,I533870,I534533,I534559,I534576,I534584,I534601,I534618,I534635,I534652,I534669,I534700,I534717,I534748,I534765,I534782,I534813,I534853,I534861,I534878,I534895,I534912,I534943,I534960,I534977,I535003,I535025,I535042,I535073,I535118,I535179,I535205,I535222,I535230,I535247,I535264,I535281,I535298,I535315,I535346,I535363,I535394,I535411,I535428,I535459,I535499,I535507,I535524,I535541,I535558,I535589,I535606,I535623,I535649,I535671,I535688,I535719,I535764,I535825,I535851,I535868,I535876,I535893,I535910,I535927,I535944,I535961,I535811,I535992,I536009,I535814,I536040,I536057,I536074,I535790,I536105,I535802,I536145,I536153,I536170,I536187,I536204,I535817,I536235,I536252,I536269,I536295,I535805,I536317,I536334,I535799,I536365,I535793,I535796,I536410,I535808,I536471,I536497,I536514,I536522,I536539,I536556,I536573,I536590,I536607,I536638,I536655,I536686,I536703,I536720,I536751,I536791,I536799,I536816,I536833,I536850,I536881,I536898,I536915,I536941,I536963,I536980,I537011,I537056,I537117,I662135,I537143,I662141,I537160,I537168,I537185,I662138,I537202,I662117,I537219,I662120,I537236,I662126,I537253,I537103,I537284,I537301,I537106,I537332,I537349,I537366,I537082,I537397,I537094,I537437,I537445,I537462,I537479,I662129,I537496,I537109,I537527,I537544,I662123,I537561,I662132,I537587,I537097,I537609,I537626,I537091,I537657,I537085,I537088,I537702,I537100,I537763,I687224,I537789,I687221,I537806,I537814,I537831,I687218,I537848,I687209,I537865,I687230,I537882,I537899,I537930,I537947,I537978,I537995,I687233,I538012,I538043,I538083,I538091,I538108,I538125,I687212,I538142,I538173,I687215,I538190,I687236,I538207,I687227,I538233,I538255,I538272,I538303,I538348,I538409,I538435,I538452,I538460,I538477,I538494,I538511,I538528,I538545,I538576,I538593,I538624,I538641,I538658,I538689,I538729,I538737,I538754,I538771,I538788,I538819,I538836,I538853,I538879,I538901,I538918,I538949,I538994,I539055,I539081,I539098,I539106,I539123,I539140,I539157,I539174,I539191,I539041,I539222,I539239,I539044,I539270,I539287,I539304,I539020,I539335,I539032,I539375,I539383,I539400,I539417,I539434,I539047,I539465,I539482,I539499,I539525,I539035,I539547,I539564,I539029,I539595,I539023,I539026,I539640,I539038,I539695,I539721,I539738,I539760,I539786,I539794,I539811,I539828,I539845,I539862,I539879,I539896,I539927,I539958,I539975,I539992,I540009,I540040,I540085,I540102,I540119,I540145,I540153,I540184,I540201,I540256,I540282,I540299,I540321,I540347,I540355,I540372,I540389,I540406,I540423,I540440,I540457,I540488,I540519,I540536,I540553,I540570,I540601,I540646,I540663,I540680,I540706,I540714,I540745,I540762,I540817,I540843,I540860,I540882,I540908,I540916,I540933,I540950,I540967,I540984,I541001,I541018,I541049,I541080,I541097,I541114,I541131,I541162,I541207,I541224,I541241,I541267,I541275,I541306,I541323,I541378,I541404,I541421,I541443,I541469,I541477,I541494,I541511,I541528,I541545,I541562,I541579,I541610,I541641,I541658,I541675,I541692,I541723,I541768,I541785,I541802,I541828,I541836,I541867,I541884,I541939,I541965,I541982,I542004,I542030,I542038,I542055,I542072,I542089,I542106,I542123,I542140,I542171,I542202,I542219,I542236,I542253,I542284,I542329,I542346,I542363,I542389,I542397,I542428,I542445,I542500,I615042,I542526,I542543,I542565,I615033,I542591,I542599,I615030,I542616,I542633,I615039,I542650,I615048,I542667,I542684,I615027,I542701,I542732,I542763,I615036,I542780,I542797,I542814,I542845,I542890,I615051,I542907,I542924,I615045,I542950,I542958,I542989,I543006,I543061,I543087,I543104,I543053,I543126,I543152,I543160,I543177,I543194,I543211,I543228,I543245,I543262,I543035,I543293,I543038,I543324,I543341,I543358,I543375,I543047,I543406,I543050,I543044,I543451,I543468,I543485,I543511,I543519,I543032,I543550,I543567,I543041,I543622,I543648,I543665,I543687,I543713,I543721,I543738,I543755,I543772,I543789,I543806,I543823,I543854,I543885,I543902,I543919,I543936,I543967,I544012,I544029,I544046,I544072,I544080,I544111,I544128,I544183,I544209,I544226,I544248,I544274,I544282,I544299,I544316,I544333,I544350,I544367,I544384,I544415,I544446,I544463,I544480,I544497,I544528,I544573,I544590,I544607,I544633,I544641,I544672,I544689,I544744,I544770,I544787,I544809,I544835,I544843,I544860,I544877,I544894,I544911,I544928,I544945,I544976,I545007,I545024,I545041,I545058,I545089,I545134,I545151,I545168,I545194,I545202,I545233,I545250,I545305,I584986,I545331,I545348,I545370,I584977,I545396,I545404,I584974,I545421,I545438,I584983,I545455,I584992,I545472,I545489,I584971,I545506,I545537,I545568,I584980,I545585,I545602,I545619,I545650,I545695,I584995,I545712,I545729,I584989,I545755,I545763,I545794,I545811,I545866,I545892,I545909,I545931,I545957,I545965,I545982,I545999,I546016,I546033,I546050,I546067,I546098,I546129,I546146,I546163,I546180,I546211,I546256,I546273,I546290,I546316,I546324,I546355,I546372,I546427,I546453,I546470,I546492,I546518,I546526,I546543,I546560,I546577,I546594,I546611,I546628,I546659,I546690,I546707,I546724,I546741,I546772,I546817,I546834,I546851,I546877,I546885,I546916,I546933,I546988,I547014,I547031,I547053,I547079,I547087,I547104,I547121,I547138,I547155,I547172,I547189,I547220,I547251,I547268,I547285,I547302,I547333,I547378,I547395,I547412,I547438,I547446,I547477,I547494,I547549,I547575,I547592,I547614,I547640,I547648,I547665,I547682,I547699,I547716,I547733,I547750,I547781,I547812,I547829,I547846,I547863,I547894,I547939,I547956,I547973,I547999,I548007,I548038,I548055,I548110,I548136,I548153,I548102,I548175,I548201,I548209,I548226,I548243,I548260,I548277,I548294,I548311,I548084,I548342,I548087,I548373,I548390,I548407,I548424,I548096,I548455,I548099,I548093,I548500,I548517,I548534,I548560,I548568,I548081,I548599,I548616,I548090,I548671,I548697,I548714,I548736,I548762,I548770,I548787,I548804,I548821,I548838,I548855,I548872,I548903,I548934,I548951,I548968,I548985,I549016,I549061,I549078,I549095,I549121,I549129,I549160,I549177,I549232,I672286,I549258,I549275,I549297,I672283,I549323,I549331,I672289,I549348,I549365,I672298,I549382,I672292,I549399,I549416,I672304,I549433,I549464,I549495,I672301,I549512,I549529,I549546,I549577,I549622,I672295,I549639,I672307,I549656,I549682,I549690,I549721,I549738,I549793,I549819,I549836,I549858,I549884,I549892,I549909,I549926,I549943,I549960,I549977,I549994,I550025,I550056,I550073,I550090,I550107,I550138,I550183,I550200,I550217,I550243,I550251,I550282,I550299,I550354,I550380,I550397,I550346,I550419,I550445,I550453,I550470,I550487,I550504,I550521,I550538,I550555,I550328,I550586,I550331,I550617,I550634,I550651,I550668,I550340,I550699,I550343,I550337,I550744,I550761,I550778,I550804,I550812,I550325,I550843,I550860,I550334,I550915,I550941,I550958,I550980,I551006,I551014,I551031,I551048,I551065,I551082,I551099,I551116,I551147,I551178,I551195,I551212,I551229,I551260,I551305,I551322,I551339,I551365,I551373,I551404,I551421,I551476,I551502,I551519,I551468,I551541,I551567,I551575,I551592,I551609,I551626,I551643,I551660,I551677,I551450,I551708,I551453,I551739,I551756,I551773,I551790,I551462,I551821,I551465,I551459,I551866,I551883,I551900,I551926,I551934,I551447,I551965,I551982,I551456,I552037,I627180,I552063,I552080,I552102,I627171,I552128,I552136,I627168,I552153,I552170,I627177,I552187,I627186,I552204,I552221,I627165,I552238,I552269,I552300,I627174,I552317,I552334,I552351,I552382,I552427,I627189,I552444,I552461,I627183,I552487,I552495,I552526,I552543,I552598,I552624,I552641,I552663,I552689,I552697,I552714,I552731,I552748,I552765,I552782,I552799,I552830,I552861,I552878,I552895,I552912,I552943,I552988,I553005,I553022,I553048,I553056,I553087,I553104,I553159,I553185,I553202,I553151,I553224,I553250,I553258,I553275,I553292,I553309,I553326,I553343,I553360,I553133,I553391,I553136,I553422,I553439,I553456,I553473,I553145,I553504,I553148,I553142,I553549,I553566,I553583,I553609,I553617,I553130,I553648,I553665,I553139,I553720,I553746,I553763,I553712,I553785,I553811,I553819,I553836,I553853,I553870,I553887,I553904,I553921,I553694,I553952,I553697,I553983,I554000,I554017,I554034,I553706,I554065,I553709,I553703,I554110,I554127,I554144,I554170,I554178,I553691,I554209,I554226,I553700,I554281,I554307,I554324,I554346,I554372,I554380,I554397,I554414,I554431,I554448,I554465,I554482,I554513,I554544,I554561,I554578,I554595,I554626,I554671,I554688,I554705,I554731,I554739,I554770,I554787,I554842,I672864,I554868,I554885,I554834,I554907,I672861,I554933,I554941,I672867,I554958,I554975,I672876,I554992,I672870,I555009,I555026,I672882,I555043,I554816,I555074,I554819,I555105,I672879,I555122,I555139,I555156,I554828,I555187,I554831,I554825,I555232,I672873,I555249,I672885,I555266,I555292,I555300,I554813,I555331,I555348,I554822,I555403,I606950,I555429,I555446,I555468,I606941,I555494,I555502,I606938,I555519,I555536,I606947,I555553,I606956,I555570,I555587,I606935,I555604,I555635,I555666,I606944,I555683,I555700,I555717,I555748,I555793,I606959,I555810,I555827,I606953,I555853,I555861,I555892,I555909,I555964,I640363,I555990,I556007,I556029,I640369,I556055,I556063,I640378,I556080,I556097,I640357,I556114,I640360,I556131,I556148,I640372,I556165,I556196,I556227,I640366,I556244,I556261,I556278,I556309,I556354,I640381,I556371,I556388,I640375,I556414,I556422,I556453,I556470,I556525,I556551,I556568,I556590,I556616,I556624,I556641,I556658,I556675,I556692,I556709,I556726,I556757,I556788,I556805,I556822,I556839,I556870,I556915,I556932,I556949,I556975,I556983,I557014,I557031,I557086,I557112,I557129,I557151,I557177,I557185,I557202,I557219,I557236,I557253,I557270,I557287,I557318,I557349,I557366,I557383,I557400,I557431,I557476,I557493,I557510,I557536,I557544,I557575,I557592,I557647,I557673,I557690,I557639,I557712,I557738,I557746,I557763,I557780,I557797,I557814,I557831,I557848,I557621,I557879,I557624,I557910,I557927,I557944,I557961,I557633,I557992,I557636,I557630,I558037,I558054,I558071,I558097,I558105,I557618,I558136,I558153,I557627,I558208,I558234,I558251,I558273,I558299,I558307,I558324,I558341,I558358,I558375,I558392,I558409,I558440,I558471,I558488,I558505,I558522,I558553,I558598,I558615,I558632,I558658,I558666,I558697,I558714,I558769,I558795,I558812,I558761,I558834,I558860,I558868,I558885,I558902,I558919,I558936,I558953,I558970,I558743,I559001,I558746,I559032,I559049,I559066,I559083,I558755,I559114,I558758,I558752,I559159,I559176,I559193,I559219,I559227,I558740,I559258,I559275,I558749,I559330,I559356,I559373,I559395,I559421,I559429,I559446,I559463,I559480,I559497,I559514,I559531,I559562,I559593,I559610,I559627,I559644,I559675,I559720,I559737,I559754,I559780,I559788,I559819,I559836,I559891,I559917,I559934,I559883,I559956,I559982,I559990,I560007,I560024,I560041,I560058,I560075,I560092,I559865,I560123,I559868,I560154,I560171,I560188,I560205,I559877,I560236,I559880,I559874,I560281,I560298,I560315,I560341,I560349,I559862,I560380,I560397,I559871,I560452,I560478,I560495,I560517,I560543,I560551,I560568,I560585,I560602,I560619,I560636,I560653,I560684,I560715,I560732,I560749,I560766,I560797,I560842,I560859,I560876,I560902,I560910,I560941,I560958,I561013,I561039,I561056,I561005,I561078,I561104,I561112,I561129,I561146,I561163,I561180,I561197,I561214,I560987,I561245,I560990,I561276,I561293,I561310,I561327,I560999,I561358,I561002,I560996,I561403,I561420,I561437,I561463,I561471,I560984,I561502,I561519,I560993,I561574,I561600,I561617,I561566,I561639,I561665,I561673,I561690,I561707,I561724,I561741,I561758,I561775,I561548,I561806,I561551,I561837,I561854,I561871,I561888,I561560,I561919,I561563,I561557,I561964,I561981,I561998,I562024,I562032,I561545,I562063,I562080,I561554,I562135,I562161,I562178,I562127,I562200,I562226,I562234,I562251,I562268,I562285,I562302,I562319,I562336,I562109,I562367,I562112,I562398,I562415,I562432,I562449,I562121,I562480,I562124,I562118,I562525,I562542,I562559,I562585,I562593,I562106,I562624,I562641,I562115,I562696,I562722,I562739,I562761,I562787,I562795,I562812,I562829,I562846,I562863,I562880,I562897,I562928,I562959,I562976,I562993,I563010,I563041,I563086,I563103,I563120,I563146,I563154,I563185,I563202,I563257,I563283,I563300,I563249,I563322,I563348,I563356,I563373,I563390,I563407,I563424,I563441,I563458,I563231,I563489,I563234,I563520,I563537,I563554,I563571,I563243,I563602,I563246,I563240,I563647,I563664,I563681,I563707,I563715,I563228,I563746,I563763,I563237,I563818,I725763,I563844,I563861,I563883,I725757,I563909,I563917,I725748,I563934,I563951,I725775,I563968,I725760,I725769,I563985,I564002,I725754,I564019,I564050,I564081,I725772,I564098,I564115,I564132,I564163,I564208,I725766,I564225,I564242,I725751,I564268,I564276,I564307,I564324,I564379,I699583,I564405,I564422,I564371,I564444,I699577,I564470,I564478,I699568,I564495,I564512,I699595,I564529,I699580,I699589,I564546,I564563,I699574,I564580,I564353,I564611,I564356,I564642,I699592,I564659,I564676,I564693,I564365,I564724,I564368,I564362,I564769,I699586,I564786,I564803,I699571,I564829,I564837,I564350,I564868,I564885,I564359,I564940,I637584,I564966,I564983,I565005,I637575,I565031,I565039,I637572,I565056,I565073,I637581,I565090,I637590,I565107,I565124,I637569,I565141,I565172,I565203,I637578,I565220,I565237,I565254,I565285,I565330,I637593,I565347,I565364,I637587,I565390,I565398,I565429,I565446,I565501,I565527,I565544,I565566,I565592,I565600,I565617,I565634,I565651,I565668,I565685,I565702,I565733,I565764,I565781,I565798,I565815,I565846,I565891,I565908,I565925,I565951,I565959,I565990,I566007,I566062,I566088,I566105,I566054,I566127,I566153,I566161,I566178,I566195,I566212,I566229,I566246,I566263,I566036,I566294,I566039,I566325,I566342,I566359,I566376,I566048,I566407,I566051,I566045,I566452,I566469,I566486,I566512,I566520,I566033,I566551,I566568,I566042,I566623,I566649,I566666,I566615,I566688,I566714,I566722,I566739,I566756,I566773,I566790,I566807,I566824,I566597,I566855,I566600,I566886,I566903,I566920,I566937,I566609,I566968,I566612,I566606,I567013,I567030,I567047,I567073,I567081,I566594,I567112,I567129,I566603,I567184,I567210,I567227,I567249,I567275,I567283,I567300,I567317,I567334,I567351,I567368,I567385,I567416,I567447,I567464,I567481,I567498,I567529,I567574,I567591,I567608,I567634,I567642,I567673,I567690,I567745,I567771,I567788,I567810,I567836,I567844,I567861,I567878,I567895,I567912,I567929,I567946,I567977,I568008,I568025,I568042,I568059,I568090,I568135,I568152,I568169,I568195,I568203,I568234,I568251,I568306,I568332,I568349,I568371,I568397,I568405,I568422,I568439,I568456,I568473,I568490,I568507,I568538,I568569,I568586,I568603,I568620,I568651,I568696,I568713,I568730,I568756,I568764,I568795,I568812,I568867,I568893,I568910,I568932,I568958,I568966,I568983,I569000,I569017,I569034,I569051,I569068,I569099,I569130,I569147,I569164,I569181,I569212,I569257,I569274,I569291,I569317,I569325,I569356,I569373,I569428,I569454,I569471,I569493,I569519,I569527,I569544,I569561,I569578,I569595,I569612,I569629,I569660,I569691,I569708,I569725,I569742,I569773,I569818,I569835,I569852,I569878,I569886,I569917,I569934,I569989,I570015,I570032,I570054,I570080,I570088,I570105,I570122,I570139,I570156,I570173,I570190,I570221,I570252,I570269,I570286,I570303,I570334,I570379,I570396,I570413,I570439,I570447,I570478,I570495,I570553,I570579,I570587,I570536,I570627,I570635,I570652,I570669,I570524,I570709,I570545,I570731,I570748,I570774,I570782,I570799,I570816,I570833,I570850,I570521,I570542,I570895,I570533,I570926,I570943,I570969,I570977,I570539,I571008,I571025,I571042,I571059,I570530,I570527,I571131,I694240,I571157,I571165,I694222,I694213,I571205,I571213,I694228,I571230,I694216,I571247,I571287,I571309,I694225,I571326,I571352,I571360,I571377,I694234,I571394,I571411,I571428,I571473,I694237,I571504,I571521,I694231,I694219,I571547,I571555,I571586,I571603,I571620,I571637,I571709,I571735,I571743,I571783,I571791,I571808,I571825,I571865,I571887,I571904,I571930,I571938,I571955,I571972,I571989,I572006,I572051,I572082,I572099,I572125,I572133,I572164,I572181,I572198,I572215,I572287,I572313,I572321,I572361,I572369,I572386,I572403,I572443,I572465,I572482,I572508,I572516,I572533,I572550,I572567,I572584,I572629,I572660,I572677,I572703,I572711,I572742,I572759,I572776,I572793,I572865,I572891,I572899,I572939,I572947,I572964,I572981,I573021,I573043,I573060,I573086,I573094,I573111,I573128,I573145,I573162,I573207,I573238,I573255,I573281,I573289,I573320,I573337,I573354,I573371,I573443,I573469,I573477,I573517,I573525,I573542,I573559,I573599,I573621,I573638,I573664,I573672,I573689,I573706,I573723,I573740,I573785,I573816,I573833,I573859,I573867,I573898,I573915,I573932,I573949,I574021,I574047,I574055,I574095,I574103,I574120,I574137,I574177,I574199,I574216,I574242,I574250,I574267,I574284,I574301,I574318,I574363,I574394,I574411,I574437,I574445,I574476,I574493,I574510,I574527,I574599,I574625,I574633,I574673,I574681,I574698,I574715,I574755,I574777,I574794,I574820,I574828,I574845,I574862,I574879,I574896,I574941,I574972,I574989,I575015,I575023,I575054,I575071,I575088,I575105,I575177,I575203,I575211,I575251,I575259,I575276,I575293,I575333,I575355,I575372,I575398,I575406,I575423,I575440,I575457,I575474,I575519,I575550,I575567,I575593,I575601,I575632,I575649,I575666,I575683,I575755,I575781,I575789,I575829,I575837,I575854,I575871,I575911,I575933,I575950,I575976,I575984,I576001,I576018,I576035,I576052,I576097,I576128,I576145,I576171,I576179,I576210,I576227,I576244,I576261,I576333,I576359,I576367,I576407,I576415,I576432,I576449,I576489,I576511,I576528,I576554,I576562,I576579,I576596,I576613,I576630,I576675,I576706,I576723,I576749,I576757,I576788,I576805,I576822,I576839,I576911,I726370,I576937,I576945,I726352,I726343,I576985,I576993,I726358,I577010,I726346,I577027,I577067,I577089,I726355,I577106,I577132,I577140,I577157,I726364,I577174,I577191,I577208,I577253,I726367,I577284,I577301,I726361,I726349,I577327,I577335,I577366,I577383,I577400,I577417,I577489,I577515,I577523,I577563,I577571,I577588,I577605,I577645,I577667,I577684,I577710,I577718,I577735,I577752,I577769,I577786,I577831,I577862,I577879,I577905,I577913,I577944,I577961,I577978,I577995,I578067,I578093,I578101,I578141,I578149,I578166,I578183,I578223,I578245,I578262,I578288,I578296,I578313,I578330,I578347,I578364,I578409,I578440,I578457,I578483,I578491,I578522,I578539,I578556,I578573,I578645,I578671,I578679,I578719,I578727,I578744,I578761,I578801,I578823,I578840,I578866,I578874,I578891,I578908,I578925,I578942,I578987,I579018,I579035,I579061,I579069,I579100,I579117,I579134,I579151,I579223,I579249,I579257,I579206,I579297,I579305,I579322,I579339,I579194,I579379,I579215,I579401,I579418,I579444,I579452,I579469,I579486,I579503,I579520,I579191,I579212,I579565,I579203,I579596,I579613,I579639,I579647,I579209,I579678,I579695,I579712,I579729,I579200,I579197,I579801,I579827,I579835,I579784,I579875,I579883,I579900,I579917,I579772,I579957,I579793,I579979,I579996,I580022,I580030,I580047,I580064,I580081,I580098,I579769,I579790,I580143,I579781,I580174,I580191,I580217,I580225,I579787,I580256,I580273,I580290,I580307,I579778,I579775,I580379,I713280,I580405,I580413,I713262,I713253,I580453,I580461,I713268,I580478,I713256,I580495,I580535,I580557,I713265,I580574,I580600,I580608,I580625,I713274,I580642,I580659,I580676,I580721,I713277,I580752,I580769,I713271,I713259,I580795,I580803,I580834,I580851,I580868,I580885,I580957,I723395,I580983,I580991,I723377,I723368,I581031,I581039,I723383,I581056,I723371,I581073,I581113,I581135,I723380,I581152,I581178,I581186,I581203,I723389,I581220,I581237,I581254,I581299,I723392,I581330,I581347,I723386,I723374,I581373,I581381,I581412,I581429,I581446,I581463,I581535,I581561,I581569,I581609,I581617,I581634,I581651,I581691,I581713,I581730,I581756,I581764,I581781,I581798,I581815,I581832,I581877,I581908,I581925,I581951,I581959,I581990,I582007,I582024,I582041,I582113,I582139,I582147,I582096,I582187,I582195,I582212,I582229,I582084,I582269,I582105,I582291,I582308,I582334,I582342,I582359,I582376,I582393,I582410,I582081,I582102,I582455,I582093,I582486,I582503,I582529,I582537,I582099,I582568,I582585,I582602,I582619,I582090,I582087,I582691,I582717,I582725,I582765,I582773,I582790,I582807,I582847,I582869,I582886,I582912,I582920,I582937,I582954,I582971,I582988,I583033,I583064,I583081,I583107,I583115,I583146,I583163,I583180,I583197,I583269,I583295,I583303,I583252,I583343,I583351,I583368,I583385,I583240,I583425,I583261,I583447,I583464,I583490,I583498,I583515,I583532,I583549,I583566,I583237,I583258,I583611,I583249,I583642,I583659,I583685,I583693,I583255,I583724,I583741,I583758,I583775,I583246,I583243,I583847,I583873,I583881,I583921,I583929,I583946,I583963,I584003,I584025,I584042,I584068,I584076,I584093,I584110,I584127,I584144,I584189,I584220,I584237,I584263,I584271,I584302,I584319,I584336,I584353,I584425,I721015,I584451,I584459,I720997,I720988,I584499,I584507,I721003,I584524,I720991,I584541,I584581,I584603,I721000,I584620,I584646,I584654,I584671,I721009,I584688,I584705,I584722,I584767,I721012,I584798,I584815,I721006,I720994,I584841,I584849,I584880,I584897,I584914,I584931,I585003,I585029,I585037,I585077,I585085,I585102,I585119,I585159,I585181,I585198,I585224,I585232,I585249,I585266,I585283,I585300,I585345,I585376,I585393,I585419,I585427,I585458,I585475,I585492,I585509,I585581,I585607,I585615,I585655,I585663,I585680,I585697,I585737,I585759,I585776,I585802,I585810,I585827,I585844,I585861,I585878,I585923,I585954,I585971,I585997,I586005,I586036,I586053,I586070,I586087,I586159,I586185,I586193,I586233,I586241,I586258,I586275,I586315,I586337,I586354,I586380,I586388,I586405,I586422,I586439,I586456,I586501,I586532,I586549,I586575,I586583,I586614,I586631,I586648,I586665,I586737,I586763,I586771,I586811,I586819,I586836,I586853,I586893,I586915,I586932,I586958,I586966,I586983,I587000,I587017,I587034,I587079,I587110,I587127,I587153,I587161,I587192,I587209,I587226,I587243,I587315,I587341,I587349,I587389,I587397,I587414,I587431,I587471,I587493,I587510,I587536,I587544,I587561,I587578,I587595,I587612,I587657,I587688,I587705,I587731,I587739,I587770,I587787,I587804,I587821,I587893,I659962,I587919,I587927,I659956,I659941,I587967,I587975,I659947,I587992,I659959,I588009,I588049,I588071,I588088,I588114,I588122,I588139,I659965,I588156,I659953,I588173,I588190,I588235,I659944,I588266,I588283,I659950,I588309,I588317,I588348,I588365,I588382,I588399,I588471,I588497,I588505,I588545,I588553,I588570,I588587,I588627,I588649,I588666,I588692,I588700,I588717,I588734,I588751,I588768,I588813,I588844,I588861,I588887,I588895,I588926,I588943,I588960,I588977,I589049,I589075,I589083,I589123,I589131,I589148,I589165,I589205,I589227,I589244,I589270,I589278,I589295,I589312,I589329,I589346,I589391,I589422,I589439,I589465,I589473,I589504,I589521,I589538,I589555,I589627,I589653,I589661,I589701,I589709,I589726,I589743,I589783,I589805,I589822,I589848,I589856,I589873,I589890,I589907,I589924,I589969,I590000,I590017,I590043,I590051,I590082,I590099,I590116,I590133,I590205,I590231,I590239,I590279,I590287,I590304,I590321,I590361,I590383,I590400,I590426,I590434,I590451,I590468,I590485,I590502,I590547,I590578,I590595,I590621,I590629,I590660,I590677,I590694,I590711,I590783,I729345,I590809,I590817,I729327,I729318,I590857,I590865,I729333,I590882,I729321,I590899,I590939,I590961,I729330,I590978,I591004,I591012,I591029,I729339,I591046,I591063,I591080,I591125,I729342,I591156,I591173,I729336,I729324,I591199,I591207,I591238,I591255,I591272,I591289,I591361,I696620,I591387,I591395,I696602,I591344,I696593,I591435,I591443,I696608,I591460,I696596,I591477,I591332,I591517,I591353,I591539,I696605,I591556,I591582,I591590,I591607,I696614,I591624,I591641,I591658,I591329,I591350,I591703,I696617,I591341,I591734,I591751,I696611,I696599,I591777,I591785,I591347,I591816,I591833,I591850,I591867,I591338,I591335,I591939,I591965,I591973,I592013,I592021,I592038,I592055,I592095,I592117,I592134,I592160,I592168,I592185,I592202,I592219,I592236,I592281,I592312,I592329,I592355,I592363,I592394,I592411,I592428,I592445,I592517,I592543,I592551,I592591,I592599,I592616,I592633,I592673,I592695,I592712,I592738,I592746,I592763,I592780,I592797,I592814,I592859,I592890,I592907,I592933,I592941,I592972,I592989,I593006,I593023,I593095,I593121,I593129,I593169,I593177,I593194,I593211,I593251,I593273,I593290,I593316,I593324,I593341,I593358,I593375,I593392,I593437,I593468,I593485,I593511,I593519,I593550,I593567,I593584,I593601,I593673,I593699,I593707,I593747,I593755,I593772,I593789,I593829,I593851,I593868,I593894,I593902,I593919,I593936,I593953,I593970,I594015,I594046,I594063,I594089,I594097,I594128,I594145,I594162,I594179,I594251,I594277,I594285,I594325,I594333,I594350,I594367,I594407,I594429,I594446,I594472,I594480,I594497,I594514,I594531,I594548,I594593,I594624,I594641,I594667,I594675,I594706,I594723,I594740,I594757,I594829,I594855,I594863,I594903,I594911,I594928,I594945,I594985,I595007,I595024,I595050,I595058,I595075,I595092,I595109,I595126,I595171,I595202,I595219,I595245,I595253,I595284,I595301,I595318,I595335,I595407,I595433,I595441,I595481,I595489,I595506,I595523,I595563,I595585,I595602,I595628,I595636,I595653,I595670,I595687,I595704,I595749,I595780,I595797,I595823,I595831,I595862,I595879,I595896,I595913,I595985,I596011,I596019,I596059,I596067,I596084,I596101,I596141,I596163,I596180,I596206,I596214,I596231,I596248,I596265,I596282,I596327,I596358,I596375,I596401,I596409,I596440,I596457,I596474,I596491,I596563,I596589,I596597,I596546,I596637,I596645,I596662,I596679,I596534,I596719,I596555,I596741,I596758,I596784,I596792,I596809,I596826,I596843,I596860,I596531,I596552,I596905,I596543,I596936,I596953,I596979,I596987,I596549,I597018,I597035,I597052,I597069,I596540,I596537,I597141,I597167,I597175,I597215,I597223,I597240,I597257,I597297,I597319,I597336,I597362,I597370,I597387,I597404,I597421,I597438,I597483,I597514,I597531,I597557,I597565,I597596,I597613,I597630,I597647,I597719,I597745,I597753,I597793,I597801,I597818,I597835,I597875,I597897,I597914,I597940,I597948,I597965,I597982,I597999,I598016,I598061,I598092,I598109,I598135,I598143,I598174,I598191,I598208,I598225,I598297,I598323,I598331,I598280,I598371,I598379,I598396,I598413,I598268,I598453,I598289,I598475,I598492,I598518,I598526,I598543,I598560,I598577,I598594,I598265,I598286,I598639,I598277,I598670,I598687,I598713,I598721,I598283,I598752,I598769,I598786,I598803,I598274,I598271,I598875,I598901,I598909,I598949,I598957,I598974,I598991,I599031,I599053,I599070,I599096,I599104,I599121,I599138,I599155,I599172,I599217,I599248,I599265,I599291,I599299,I599330,I599347,I599364,I599381,I599453,I599479,I599487,I599527,I599535,I599552,I599569,I599609,I599631,I599648,I599674,I599682,I599699,I599716,I599733,I599750,I599795,I599826,I599843,I599869,I599877,I599908,I599925,I599942,I599959,I600031,I600057,I600065,I600014,I600105,I600113,I600130,I600147,I600002,I600187,I600023,I600209,I600226,I600252,I600260,I600277,I600294,I600311,I600328,I599999,I600020,I600373,I600011,I600404,I600421,I600447,I600455,I600017,I600486,I600503,I600520,I600537,I600008,I600005,I600609,I600635,I600643,I600683,I600691,I600708,I600725,I600765,I600787,I600804,I600830,I600838,I600855,I600872,I600889,I600906,I600951,I600982,I600999,I601025,I601033,I601064,I601081,I601098,I601115,I601187,I655066,I601213,I601221,I655060,I655045,I601261,I601269,I655051,I601286,I655063,I601303,I601343,I601365,I601382,I601408,I601416,I601433,I655069,I601450,I655057,I601467,I601484,I601529,I655048,I601560,I601577,I655054,I601603,I601611,I601642,I601659,I601676,I601693,I601765,I601791,I601799,I601748,I601839,I601847,I601864,I601881,I601736,I601921,I601757,I601943,I601960,I601986,I601994,I602011,I602028,I602045,I602062,I601733,I601754,I602107,I601745,I602138,I602155,I602181,I602189,I601751,I602220,I602237,I602254,I602271,I601742,I601739,I602343,I602369,I602377,I602417,I602425,I602442,I602459,I602499,I602521,I602538,I602564,I602572,I602589,I602606,I602623,I602640,I602685,I602716,I602733,I602759,I602767,I602798,I602815,I602832,I602849,I602921,I602947,I602955,I602904,I602995,I603003,I603020,I603037,I602892,I603077,I602913,I603099,I603116,I603142,I603150,I603167,I603184,I603201,I603218,I602889,I602910,I603263,I602901,I603294,I603311,I603337,I603345,I602907,I603376,I603393,I603410,I603427,I602898,I602895,I603499,I696025,I603525,I603533,I696007,I695998,I603573,I603581,I696013,I603598,I696001,I603615,I603655,I603677,I696010,I603694,I603720,I603728,I603745,I696019,I603762,I603779,I603796,I603841,I696022,I603872,I603889,I696016,I696004,I603915,I603923,I603954,I603971,I603988,I604005,I604077,I604103,I604111,I604151,I604159,I604176,I604193,I604233,I604255,I604272,I604298,I604306,I604323,I604340,I604357,I604374,I604419,I604450,I604467,I604493,I604501,I604532,I604549,I604566,I604583,I604655,I604681,I604689,I604729,I604737,I604754,I604771,I604811,I604833,I604850,I604876,I604884,I604901,I604918,I604935,I604952,I604997,I605028,I605045,I605071,I605079,I605110,I605127,I605144,I605161,I605233,I605259,I605267,I605307,I605315,I605332,I605349,I605389,I605411,I605428,I605454,I605462,I605479,I605496,I605513,I605530,I605575,I605606,I605623,I605649,I605657,I605688,I605705,I605722,I605739,I605811,I605837,I605845,I605885,I605893,I605910,I605927,I605967,I605989,I606006,I606032,I606040,I606057,I606074,I606091,I606108,I606153,I606184,I606201,I606227,I606235,I606266,I606283,I606300,I606317,I606389,I665402,I606415,I606423,I665396,I665381,I606463,I606471,I665387,I606488,I665399,I606505,I606545,I606567,I606584,I606610,I606618,I606635,I665405,I606652,I665393,I606669,I606686,I606731,I665384,I606762,I606779,I665390,I606805,I606813,I606844,I606861,I606878,I606895,I606967,I606993,I607001,I607041,I607049,I607066,I607083,I607123,I607145,I607162,I607188,I607196,I607213,I607230,I607247,I607264,I607309,I607340,I607357,I607383,I607391,I607422,I607439,I607456,I607473,I607545,I607571,I607579,I607619,I607627,I607644,I607661,I607701,I607723,I607740,I607766,I607774,I607791,I607808,I607825,I607842,I607887,I607918,I607935,I607961,I607969,I608000,I608017,I608034,I608051,I608123,I608149,I608157,I608197,I608205,I608222,I608239,I608279,I608301,I608318,I608344,I608352,I608369,I608386,I608403,I608420,I608465,I608496,I608513,I608539,I608547,I608578,I608595,I608612,I608629,I608701,I608727,I608735,I608775,I608783,I608800,I608817,I608857,I608879,I608896,I608922,I608930,I608947,I608964,I608981,I608998,I609043,I609074,I609091,I609117,I609125,I609156,I609173,I609190,I609207,I609279,I609305,I609313,I609262,I609353,I609361,I609378,I609395,I609250,I609435,I609271,I609457,I609474,I609500,I609508,I609525,I609542,I609559,I609576,I609247,I609268,I609621,I609259,I609652,I609669,I609695,I609703,I609265,I609734,I609751,I609768,I609785,I609256,I609253,I609857,I609883,I609891,I609931,I609939,I609956,I609973,I610013,I610035,I610052,I610078,I610086,I610103,I610120,I610137,I610154,I610199,I610230,I610247,I610273,I610281,I610312,I610329,I610346,I610363,I610435,I610461,I610469,I610418,I610509,I610517,I610534,I610551,I610406,I610591,I610427,I610613,I610630,I610656,I610664,I610681,I610698,I610715,I610732,I610403,I610424,I610777,I610415,I610808,I610825,I610851,I610859,I610421,I610890,I610907,I610924,I610941,I610412,I610409,I611013,I611039,I611047,I610996,I611087,I611095,I611112,I611129,I610984,I611169,I611005,I611191,I611208,I611234,I611242,I611259,I611276,I611293,I611310,I610981,I611002,I611355,I610993,I611386,I611403,I611429,I611437,I610999,I611468,I611485,I611502,I611519,I610990,I610987,I611591,I611617,I611625,I611665,I611673,I611690,I611707,I611747,I611769,I611786,I611812,I611820,I611837,I611854,I611871,I611888,I611933,I611964,I611981,I612007,I612015,I612046,I612063,I612080,I612097,I612169,I612195,I612203,I612243,I612251,I612268,I612285,I612325,I612347,I612364,I612390,I612398,I612415,I612432,I612449,I612466,I612511,I612542,I612559,I612585,I612593,I612624,I612641,I612658,I612675,I612747,I612773,I612781,I612821,I612829,I612846,I612863,I612903,I612925,I612942,I612968,I612976,I612993,I613010,I613027,I613044,I613089,I613120,I613137,I613163,I613171,I613202,I613219,I613236,I613253,I613325,I613351,I613359,I613399,I613407,I613424,I613441,I613481,I613503,I613520,I613546,I613554,I613571,I613588,I613605,I613622,I613667,I613698,I613715,I613741,I613749,I613780,I613797,I613814,I613831,I613903,I613929,I613937,I613886,I613977,I613985,I614002,I614019,I613874,I614059,I613895,I614081,I614098,I614124,I614132,I614149,I614166,I614183,I614200,I613871,I613892,I614245,I613883,I614276,I614293,I614319,I614327,I613889,I614358,I614375,I614392,I614409,I613880,I613877,I614481,I657786,I614507,I614515,I657780,I657765,I614555,I614563,I657771,I614580,I657783,I614597,I614637,I614659,I614676,I614702,I614710,I614727,I657789,I614744,I657777,I614761,I614778,I614823,I657768,I614854,I614871,I657774,I614897,I614905,I614936,I614953,I614970,I614987,I615059,I615085,I615093,I615133,I615141,I615158,I615175,I615215,I615237,I615254,I615280,I615288,I615305,I615322,I615339,I615356,I615401,I615432,I615449,I615475,I615483,I615514,I615531,I615548,I615565,I615637,I615663,I615671,I615711,I615719,I615736,I615753,I615793,I615815,I615832,I615858,I615866,I615883,I615900,I615917,I615934,I615979,I616010,I616027,I616053,I616061,I616092,I616109,I616126,I616143,I616215,I616241,I616249,I616289,I616297,I616314,I616331,I616371,I616393,I616410,I616436,I616444,I616461,I616478,I616495,I616512,I616557,I616588,I616605,I616631,I616639,I616670,I616687,I616704,I616721,I616793,I616819,I616827,I616867,I616875,I616892,I616909,I616949,I616971,I616988,I617014,I617022,I617039,I617056,I617073,I617090,I617135,I617166,I617183,I617209,I617217,I617248,I617265,I617282,I617299,I617371,I617397,I617405,I617445,I617453,I617470,I617487,I617527,I617549,I617566,I617592,I617600,I617617,I617634,I617651,I617668,I617713,I617744,I617761,I617787,I617795,I617826,I617843,I617860,I617877,I617949,I617975,I617983,I618023,I618031,I618048,I618065,I618105,I618127,I618144,I618170,I618178,I618195,I618212,I618229,I618246,I618291,I618322,I618339,I618365,I618373,I618404,I618421,I618438,I618455,I618527,I644186,I618553,I618561,I644180,I644165,I618601,I618609,I644171,I618626,I644183,I618643,I618683,I618705,I618722,I618748,I618756,I618773,I644189,I618790,I644177,I618807,I618824,I618869,I644168,I618900,I618917,I644174,I618943,I618951,I618982,I618999,I619016,I619033,I619105,I619131,I619139,I619179,I619187,I619204,I619221,I619261,I619283,I619300,I619326,I619334,I619351,I619368,I619385,I619402,I619447,I619478,I619495,I619521,I619529,I619560,I619577,I619594,I619611,I619683,I619709,I619717,I619757,I619765,I619782,I619799,I619839,I619861,I619878,I619904,I619912,I619929,I619946,I619963,I619980,I620025,I620056,I620073,I620099,I620107,I620138,I620155,I620172,I620189,I620261,I620287,I620295,I620335,I620343,I620360,I620377,I620417,I620439,I620456,I620482,I620490,I620507,I620524,I620541,I620558,I620603,I620634,I620651,I620677,I620685,I620716,I620733,I620750,I620767,I620839,I620865,I620873,I620913,I620921,I620938,I620955,I620995,I621017,I621034,I621060,I621068,I621085,I621102,I621119,I621136,I621181,I621212,I621229,I621255,I621263,I621294,I621311,I621328,I621345,I621417,I701975,I621443,I621451,I701957,I701948,I621491,I621499,I701963,I621516,I701951,I621533,I621573,I621595,I701960,I621612,I621638,I621646,I621663,I701969,I621680,I621697,I621714,I621759,I701972,I621790,I621807,I701966,I701954,I621833,I621841,I621872,I621889,I621906,I621923,I621995,I622021,I622029,I622069,I622077,I622094,I622111,I622151,I622173,I622190,I622216,I622224,I622241,I622258,I622275,I622292,I622337,I622368,I622385,I622411,I622419,I622450,I622467,I622484,I622501,I622573,I622599,I622607,I622647,I622655,I622672,I622689,I622729,I622751,I622768,I622794,I622802,I622819,I622836,I622853,I622870,I622915,I622946,I622963,I622989,I622997,I623028,I623045,I623062,I623079,I623151,I623177,I623185,I623225,I623233,I623250,I623267,I623307,I623329,I623346,I623372,I623380,I623397,I623414,I623431,I623448,I623493,I623524,I623541,I623567,I623575,I623606,I623623,I623640,I623657,I623729,I728155,I623755,I623763,I728137,I728128,I623803,I623811,I728143,I623828,I728131,I623845,I623885,I623907,I728140,I623924,I623950,I623958,I623975,I728149,I623992,I624009,I624026,I624071,I728152,I624102,I624119,I728146,I728134,I624145,I624153,I624184,I624201,I624218,I624235,I624307,I624333,I624341,I624381,I624389,I624406,I624423,I624463,I624485,I624502,I624528,I624536,I624553,I624570,I624587,I624604,I624649,I624680,I624697,I624723,I624731,I624762,I624779,I624796,I624813,I624885,I624911,I624919,I624959,I624967,I624984,I625001,I625041,I625063,I625080,I625106,I625114,I625131,I625148,I625165,I625182,I625227,I625258,I625275,I625301,I625309,I625340,I625357,I625374,I625391,I625463,I625489,I625497,I625446,I625537,I625545,I625562,I625579,I625434,I625619,I625455,I625641,I625658,I625684,I625692,I625709,I625726,I625743,I625760,I625431,I625452,I625805,I625443,I625836,I625853,I625879,I625887,I625449,I625918,I625935,I625952,I625969,I625440,I625437,I626041,I626067,I626075,I626115,I626123,I626140,I626157,I626197,I626219,I626236,I626262,I626270,I626287,I626304,I626321,I626338,I626383,I626414,I626431,I626457,I626465,I626496,I626513,I626530,I626547,I626619,I626645,I626653,I626693,I626701,I626718,I626735,I626775,I626797,I626814,I626840,I626848,I626865,I626882,I626899,I626916,I626961,I626992,I627009,I627035,I627043,I627074,I627091,I627108,I627125,I627197,I627223,I627231,I627271,I627279,I627296,I627313,I627353,I627375,I627392,I627418,I627426,I627443,I627460,I627477,I627494,I627539,I627570,I627587,I627613,I627621,I627652,I627669,I627686,I627703,I627775,I627801,I627809,I627849,I627857,I627874,I627891,I627931,I627953,I627970,I627996,I628004,I628021,I628038,I628055,I628072,I628117,I628148,I628165,I628191,I628199,I628230,I628247,I628264,I628281,I628353,I628379,I628387,I628427,I628435,I628452,I628469,I628509,I628531,I628548,I628574,I628582,I628599,I628616,I628633,I628650,I628695,I628726,I628743,I628769,I628777,I628808,I628825,I628842,I628859,I628931,I628957,I628965,I629005,I629013,I629030,I629047,I629087,I629109,I629126,I629152,I629160,I629177,I629194,I629211,I629228,I629273,I629304,I629321,I629347,I629355,I629386,I629403,I629420,I629437,I629509,I629535,I629543,I629583,I629591,I629608,I629625,I629665,I629687,I629704,I629730,I629738,I629755,I629772,I629789,I629806,I629851,I629882,I629899,I629925,I629933,I629964,I629981,I629998,I630015,I630087,I630113,I630121,I630161,I630169,I630186,I630203,I630243,I630265,I630282,I630308,I630316,I630333,I630350,I630367,I630384,I630429,I630460,I630477,I630503,I630511,I630542,I630559,I630576,I630593,I630665,I630691,I630699,I630739,I630747,I630764,I630781,I630821,I630843,I630860,I630886,I630894,I630911,I630928,I630945,I630962,I631007,I631038,I631055,I631081,I631089,I631120,I631137,I631154,I631171,I631243,I631269,I631277,I631317,I631325,I631342,I631359,I631399,I631421,I631438,I631464,I631472,I631489,I631506,I631523,I631540,I631585,I631616,I631633,I631659,I631667,I631698,I631715,I631732,I631749,I631821,I631847,I631855,I631895,I631903,I631920,I631937,I631977,I631999,I632016,I632042,I632050,I632067,I632084,I632101,I632118,I632163,I632194,I632211,I632237,I632245,I632276,I632293,I632310,I632327,I632399,I632425,I632433,I632473,I632481,I632498,I632515,I632555,I632577,I632594,I632620,I632628,I632645,I632662,I632679,I632696,I632741,I632772,I632789,I632815,I632823,I632854,I632871,I632888,I632905,I632977,I633003,I633011,I633051,I633059,I633076,I633093,I633133,I633155,I633172,I633198,I633206,I633223,I633240,I633257,I633274,I633319,I633350,I633367,I633393,I633401,I633432,I633449,I633466,I633483,I633555,I660506,I633581,I633589,I660500,I660485,I633629,I633637,I660491,I633654,I660503,I633671,I633711,I633733,I633750,I633776,I633784,I633801,I660509,I633818,I660497,I633835,I633852,I633897,I660488,I633928,I633945,I660494,I633971,I633979,I634010,I634027,I634044,I634061,I634133,I634159,I634167,I634207,I634215,I634232,I634249,I634289,I634311,I634328,I634354,I634362,I634379,I634396,I634413,I634430,I634475,I634506,I634523,I634549,I634557,I634588,I634605,I634622,I634639,I634711,I634737,I634745,I634694,I634785,I634793,I634810,I634827,I634682,I634867,I634703,I634889,I634906,I634932,I634940,I634957,I634974,I634991,I635008,I634679,I634700,I635053,I634691,I635084,I635101,I635127,I635135,I634697,I635166,I635183,I635200,I635217,I634688,I634685,I635289,I635315,I635323,I635363,I635371,I635388,I635405,I635445,I635467,I635484,I635510,I635518,I635535,I635552,I635569,I635586,I635631,I635662,I635679,I635705,I635713,I635744,I635761,I635778,I635795,I635867,I635893,I635901,I635941,I635949,I635966,I635983,I636023,I636045,I636062,I636088,I636096,I636113,I636130,I636147,I636164,I636209,I636240,I636257,I636283,I636291,I636322,I636339,I636356,I636373,I636445,I636471,I636479,I636519,I636527,I636544,I636561,I636601,I636623,I636640,I636666,I636674,I636691,I636708,I636725,I636742,I636787,I636818,I636835,I636861,I636869,I636900,I636917,I636934,I636951,I637023,I637049,I637057,I637097,I637105,I637122,I637139,I637179,I637201,I637218,I637244,I637252,I637269,I637286,I637303,I637320,I637365,I637396,I637413,I637439,I637447,I637478,I637495,I637512,I637529,I637601,I637627,I637635,I637675,I637683,I637700,I637717,I637757,I637779,I637796,I637822,I637830,I637847,I637864,I637881,I637898,I637943,I637974,I637991,I638017,I638025,I638056,I638073,I638090,I638107,I638179,I638205,I638213,I638253,I638261,I638278,I638295,I638335,I638357,I638374,I638400,I638408,I638425,I638442,I638459,I638476,I638521,I638552,I638569,I638595,I638603,I638634,I638651,I638668,I638685,I638757,I638783,I638791,I638817,I638834,I638856,I638873,I638890,I638907,I638924,I638955,I638972,I638989,I639006,I639051,I639068,I639085,I639144,I639170,I639178,I639195,I639212,I639243,I639301,I639327,I639335,I639361,I639378,I639400,I639417,I639434,I639451,I639468,I639499,I639516,I639533,I639550,I639595,I639612,I639629,I639688,I639714,I639722,I639739,I639756,I639787,I639845,I639871,I639879,I639905,I639922,I639944,I639961,I639978,I639995,I640012,I640043,I640060,I640077,I640094,I640139,I640156,I640173,I640232,I640258,I640266,I640283,I640300,I640331,I640389,I640415,I640423,I640449,I640466,I640488,I640505,I640522,I640539,I640556,I640587,I640604,I640621,I640638,I640683,I640700,I640717,I640776,I640802,I640810,I640827,I640844,I640875,I640933,I640959,I640967,I640993,I641010,I641032,I641049,I641066,I641083,I641100,I641131,I641148,I641165,I641182,I641227,I641244,I641261,I641320,I641346,I641354,I641371,I641388,I641419,I641477,I641503,I641511,I641537,I641554,I641576,I641593,I641610,I641627,I641644,I641675,I641692,I641709,I641726,I641771,I641788,I641805,I641864,I641890,I641898,I641915,I641932,I641963,I642021,I642047,I642055,I642081,I642098,I642120,I642137,I642154,I642171,I642188,I642219,I642236,I642253,I642270,I642315,I642332,I642349,I642408,I642434,I642442,I642459,I642476,I642507,I642565,I642591,I642599,I642625,I642642,I642664,I642681,I642698,I642715,I642732,I642763,I642780,I642797,I642814,I642859,I642876,I642893,I642952,I642978,I642986,I643003,I643020,I643051,I643109,I643135,I643143,I643169,I643186,I643208,I643225,I643242,I643259,I643276,I643307,I643324,I643341,I643358,I643403,I643420,I643437,I643496,I643522,I643530,I643547,I643564,I643595,I643653,I643679,I643687,I643713,I643730,I643752,I643769,I643786,I643803,I643820,I643851,I643868,I643885,I643902,I643947,I643964,I643981,I644040,I644066,I644074,I644091,I644108,I644139,I644197,I722205,I644223,I644231,I722190,I722184,I644257,I644274,I644296,I722178,I644313,I722199,I644330,I722187,I644347,I644364,I644395,I722196,I644412,I722202,I644429,I722193,I644446,I644491,I722181,I644508,I644525,I644584,I644610,I644618,I644635,I644652,I644683,I644741,I644767,I644775,I644801,I644818,I644840,I644857,I644874,I644891,I644908,I644939,I644956,I644973,I644990,I645035,I645052,I645069,I645128,I645154,I645162,I645179,I645196,I645227,I645285,I645311,I645319,I645345,I645362,I645384,I645401,I645418,I645435,I645452,I645483,I645500,I645517,I645534,I645579,I645596,I645613,I645672,I645698,I645706,I645723,I645740,I645771,I645829,I645855,I645863,I645889,I645906,I645928,I645945,I645962,I645979,I645996,I646027,I646044,I646061,I646078,I646123,I646140,I646157,I646216,I646242,I646250,I646267,I646284,I646315,I646373,I646399,I646407,I646433,I646450,I646472,I646489,I646506,I646523,I646540,I646571,I646588,I646605,I646622,I646667,I646684,I646701,I646760,I646786,I646794,I646811,I646828,I646859,I646917,I646943,I646951,I646977,I646994,I647016,I647033,I647050,I647067,I647084,I647115,I647132,I647149,I647166,I647211,I647228,I647245,I647304,I647330,I647338,I647355,I647372,I647403,I647461,I647487,I647495,I647521,I647538,I647560,I647577,I647594,I647611,I647628,I647659,I647676,I647693,I647710,I647755,I647772,I647789,I647848,I647874,I647882,I647899,I647916,I647947,I648005,I648031,I648039,I648065,I648082,I648104,I648121,I648138,I648155,I648172,I648203,I648220,I648237,I648254,I648299,I648316,I648333,I648392,I648418,I648426,I648443,I648460,I648491,I648549,I648575,I648583,I648609,I648626,I648648,I648665,I648682,I648699,I648716,I648747,I648764,I648781,I648798,I648843,I648860,I648877,I648936,I648962,I648970,I648987,I649004,I649035,I649093,I649119,I649127,I649153,I649170,I649192,I649209,I649226,I649243,I649260,I649291,I649308,I649325,I649342,I649387,I649404,I649421,I649480,I649506,I649514,I649531,I649548,I649579,I649637,I649663,I649671,I649697,I649714,I649736,I649753,I649770,I649787,I649804,I649835,I649852,I649869,I649886,I649931,I649948,I649965,I650024,I650050,I650058,I650075,I650092,I650123,I650181,I650207,I650215,I650241,I650258,I650280,I650297,I650314,I650331,I650348,I650379,I650396,I650413,I650430,I650475,I650492,I650509,I650568,I650594,I650602,I650619,I650636,I650667,I650725,I650751,I650759,I650785,I650802,I650824,I650841,I650858,I650875,I650892,I650923,I650940,I650957,I650974,I651019,I651036,I651053,I651112,I651138,I651146,I651163,I651180,I651211,I651269,I731725,I651295,I651303,I731710,I731704,I651329,I651346,I651368,I731698,I651385,I731719,I651402,I731707,I651419,I651436,I651467,I731716,I651484,I731722,I651501,I731713,I651518,I651563,I731701,I651580,I651597,I651656,I651682,I651690,I651707,I651724,I651755,I651813,I651839,I651847,I651873,I651890,I651912,I651929,I651946,I651963,I651980,I652011,I652028,I652045,I652062,I652107,I652124,I652141,I652200,I652226,I652234,I652251,I652268,I652299,I652357,I652383,I652391,I652417,I652434,I652456,I652473,I652490,I652507,I652524,I652555,I652572,I652589,I652606,I652651,I652668,I652685,I652744,I652770,I652778,I652795,I652812,I652843,I652901,I652927,I652935,I652961,I652978,I653000,I653017,I653034,I653051,I653068,I653099,I653116,I653133,I653150,I653195,I653212,I653229,I653288,I653314,I653322,I653339,I653356,I653387,I653445,I653471,I653479,I653505,I653522,I653544,I653561,I653578,I653595,I653612,I653643,I653660,I653677,I653694,I653739,I653756,I653773,I653832,I653858,I653866,I653883,I653900,I653931,I653989,I654015,I654023,I654049,I654066,I654088,I654105,I654122,I654139,I654156,I654187,I654204,I654221,I654238,I654283,I654300,I654317,I654376,I654402,I654410,I654427,I654444,I654475,I654533,I654559,I654567,I654593,I654610,I654632,I654649,I654666,I654683,I654700,I654731,I654748,I654765,I654782,I654827,I654844,I654861,I654920,I654946,I654954,I654971,I654988,I655019,I655077,I655103,I655111,I655137,I655154,I655176,I655193,I655210,I655227,I655244,I655275,I655292,I655309,I655326,I655371,I655388,I655405,I655464,I655490,I655498,I655515,I655532,I655563,I655621,I655647,I655655,I655681,I655698,I655720,I655737,I655754,I655771,I655788,I655819,I655836,I655853,I655870,I655915,I655932,I655949,I656008,I656034,I656042,I656059,I656076,I656107,I656165,I656191,I656199,I656225,I656242,I656264,I656281,I656298,I656315,I656332,I656363,I656380,I656397,I656414,I656459,I656476,I656493,I656552,I656578,I656586,I656603,I656620,I656651,I656709,I656735,I656743,I656769,I656786,I656808,I656825,I656842,I656859,I656876,I656907,I656924,I656941,I656958,I657003,I657020,I657037,I657096,I657122,I657130,I657147,I657164,I657195,I657253,I657279,I657287,I657313,I657330,I657352,I657369,I657386,I657403,I657420,I657451,I657468,I657485,I657502,I657547,I657564,I657581,I657640,I657666,I657674,I657691,I657708,I657739,I657797,I657823,I657831,I657857,I657874,I657896,I657913,I657930,I657947,I657964,I657995,I658012,I658029,I658046,I658091,I658108,I658125,I658184,I658210,I658218,I658235,I658252,I658283,I658341,I658367,I658375,I658401,I658418,I658440,I658457,I658474,I658491,I658508,I658539,I658556,I658573,I658590,I658635,I658652,I658669,I658728,I658754,I658762,I658779,I658796,I658827,I658885,I658911,I658919,I658945,I658962,I658984,I659001,I659018,I659035,I659052,I659083,I659100,I659117,I659134,I659179,I659196,I659213,I659272,I659298,I659306,I659323,I659340,I659371,I659429,I659455,I659463,I659489,I659506,I659528,I659545,I659562,I659579,I659596,I659627,I659644,I659661,I659678,I659723,I659740,I659757,I659816,I659842,I659850,I659867,I659884,I659915,I659973,I659999,I660007,I660033,I660050,I660072,I660089,I660106,I660123,I660140,I660171,I660188,I660205,I660222,I660267,I660284,I660301,I660360,I660386,I660394,I660411,I660428,I660459,I660517,I660543,I660551,I660577,I660594,I660616,I660633,I660650,I660667,I660684,I660715,I660732,I660749,I660766,I660811,I660828,I660845,I660904,I660930,I660938,I660955,I660972,I661003,I661061,I661087,I661095,I661121,I661138,I661160,I661177,I661194,I661211,I661228,I661259,I661276,I661293,I661310,I661355,I661372,I661389,I661448,I661474,I661482,I661499,I661516,I661547,I661605,I731130,I661631,I661639,I731115,I731109,I661665,I661682,I661704,I731103,I661721,I731124,I661738,I731112,I661755,I661772,I661803,I731121,I661820,I731127,I661837,I731118,I661854,I661899,I731106,I661916,I661933,I661992,I662018,I662026,I662043,I662060,I662091,I662149,I723990,I662175,I662183,I723975,I723969,I662209,I662226,I662248,I723963,I662265,I723984,I662282,I723972,I662299,I662316,I662347,I723981,I662364,I723987,I662381,I723978,I662398,I662443,I723966,I662460,I662477,I662536,I662562,I662570,I662587,I662604,I662635,I662693,I662719,I662727,I662753,I662770,I662792,I662809,I662826,I662843,I662860,I662891,I662908,I662925,I662942,I662987,I663004,I663021,I663080,I663106,I663114,I663131,I663148,I663179,I663237,I663263,I663271,I663297,I663314,I663336,I663353,I663370,I663387,I663404,I663435,I663452,I663469,I663486,I663531,I663548,I663565,I663624,I663650,I663658,I663675,I663692,I663723,I663781,I663807,I663815,I663841,I663858,I663773,I663880,I663897,I663914,I663931,I663948,I663752,I663979,I663996,I664013,I664030,I663755,I663770,I664075,I664092,I664109,I663767,I663764,I663761,I664168,I664194,I664202,I664219,I664236,I663749,I664267,I663758,I664325,I664351,I664359,I664385,I664402,I664424,I664441,I664458,I664475,I664492,I664523,I664540,I664557,I664574,I664619,I664636,I664653,I664712,I664738,I664746,I664763,I664780,I664811,I664869,I664895,I664903,I664929,I664946,I664968,I664985,I665002,I665019,I665036,I665067,I665084,I665101,I665118,I665163,I665180,I665197,I665256,I665282,I665290,I665307,I665324,I665355,I665413,I665439,I665447,I665473,I665490,I665512,I665529,I665546,I665563,I665580,I665611,I665628,I665645,I665662,I665707,I665724,I665741,I665800,I665826,I665834,I665851,I665868,I665899,I665957,I665983,I665991,I666008,I666034,I666042,I666059,I666076,I666093,I666110,I666141,I666158,I666175,I666206,I666223,I666263,I666271,I666302,I666319,I666336,I666353,I666384,I666415,I666441,I666463,I666535,I666561,I666569,I666586,I666612,I666620,I666637,I666654,I666671,I666688,I666719,I666736,I666753,I666784,I666801,I666841,I666849,I666880,I666897,I666914,I666931,I666962,I666993,I667019,I667041,I667113,I667139,I667147,I667164,I667190,I667198,I667215,I667232,I667249,I667266,I667297,I667314,I667331,I667362,I667379,I667419,I667427,I667458,I667475,I667492,I667509,I667540,I667571,I667597,I667619,I667691,I667717,I667725,I667742,I667768,I667776,I667793,I667810,I667827,I667844,I667875,I667892,I667909,I667940,I667957,I667997,I668005,I668036,I668053,I668070,I668087,I668118,I668149,I668175,I668197,I668269,I668295,I668303,I668320,I668346,I668354,I668371,I668388,I668405,I668422,I668453,I668470,I668487,I668518,I668535,I668575,I668583,I668614,I668631,I668648,I668665,I668696,I668727,I668753,I668775,I668847,I668873,I668881,I668898,I668924,I668932,I668949,I668966,I668983,I669000,I669031,I669048,I669065,I669096,I669113,I669153,I669161,I669192,I669209,I669226,I669243,I669274,I669305,I669331,I669353,I669425,I669451,I669459,I669476,I669502,I669510,I669527,I669544,I669561,I669578,I669609,I669626,I669643,I669674,I669691,I669731,I669739,I669770,I669787,I669804,I669821,I669852,I669883,I669909,I669931,I670003,I670029,I670037,I670054,I670080,I670088,I670105,I670122,I670139,I670156,I670187,I670204,I670221,I670252,I670269,I670309,I670317,I670348,I670365,I670382,I670399,I670430,I670461,I670487,I670509,I670581,I670607,I670615,I670632,I670658,I670666,I670683,I670700,I670717,I670734,I670765,I670782,I670799,I670830,I670847,I670887,I670895,I670926,I670943,I670960,I670977,I671008,I671039,I671065,I671087,I671159,I671185,I671193,I671210,I671236,I671244,I671261,I671278,I671295,I671312,I671343,I671360,I671377,I671408,I671425,I671465,I671473,I671504,I671521,I671538,I671555,I671586,I671617,I671643,I671665,I671737,I671763,I671771,I671788,I671814,I671822,I671839,I671856,I671873,I671890,I671921,I671938,I671955,I671986,I672003,I672043,I672051,I672082,I672099,I672116,I672133,I672164,I672195,I672221,I672243,I672315,I672341,I672349,I672366,I672392,I672400,I672417,I672434,I672451,I672468,I672499,I672516,I672533,I672564,I672581,I672621,I672629,I672660,I672677,I672694,I672711,I672742,I672773,I672799,I672821,I672893,I672919,I672927,I672944,I672970,I672978,I672995,I673012,I673029,I673046,I673077,I673094,I673111,I673142,I673159,I673199,I673207,I673238,I673255,I673272,I673289,I673320,I673351,I673377,I673399,I673471,I673497,I673505,I673522,I673548,I673556,I673573,I673590,I673607,I673624,I673655,I673672,I673689,I673720,I673737,I673777,I673785,I673816,I673833,I673850,I673867,I673898,I673929,I673955,I673977,I674049,I674075,I674083,I674100,I674126,I674134,I674151,I674168,I674185,I674202,I674233,I674250,I674267,I674298,I674315,I674355,I674363,I674394,I674411,I674428,I674445,I674476,I674507,I674533,I674555,I674627,I674653,I674661,I674678,I674704,I674712,I674729,I674746,I674763,I674780,I674619,I674811,I674828,I674845,I674598,I674876,I674893,I674604,I674933,I674941,I674613,I674972,I674989,I675006,I675023,I674616,I675054,I674595,I675085,I675111,I674610,I675133,I674607,I674601,I675205,I675231,I675239,I675256,I675282,I675290,I675307,I675324,I675341,I675358,I675389,I675406,I675423,I675454,I675471,I675511,I675519,I675550,I675567,I675584,I675601,I675632,I675663,I675689,I675711,I675783,I675809,I675817,I675834,I675860,I675868,I675885,I675902,I675919,I675936,I675967,I675984,I676001,I676032,I676049,I676089,I676097,I676128,I676145,I676162,I676179,I676210,I676241,I676267,I676289,I676361,I676387,I676395,I676412,I676438,I676446,I676463,I676480,I676497,I676514,I676545,I676562,I676579,I676610,I676627,I676667,I676675,I676706,I676723,I676740,I676757,I676788,I676819,I676845,I676867,I676939,I676965,I676973,I676990,I677016,I677024,I677041,I677058,I677075,I677092,I677123,I677140,I677157,I677188,I677205,I677245,I677253,I677284,I677301,I677318,I677335,I677366,I677397,I677423,I677445,I677517,I677543,I677551,I677568,I677594,I677602,I677619,I677636,I677653,I677670,I677701,I677718,I677735,I677766,I677783,I677823,I677831,I677862,I677879,I677896,I677913,I677944,I677975,I678001,I678023,I678095,I678121,I678129,I678146,I678172,I678180,I678197,I678214,I678231,I678248,I678279,I678296,I678313,I678344,I678361,I678401,I678409,I678440,I678457,I678474,I678491,I678522,I678553,I678579,I678601,I678673,I725177,I678699,I678707,I725168,I678724,I725153,I678750,I678758,I678775,I725156,I678792,I725165,I678809,I678826,I725162,I678857,I725174,I678874,I678891,I678922,I725159,I678939,I678979,I678987,I679018,I725180,I679035,I679052,I679069,I679100,I679131,I725171,I679157,I679179,I679251,I679277,I679285,I679302,I679328,I679336,I679353,I679370,I679387,I679404,I679435,I679452,I679469,I679500,I679517,I679557,I679565,I679596,I679613,I679630,I679647,I679678,I679709,I679735,I679757,I679829,I679855,I679863,I679880,I679906,I679914,I679931,I679948,I679965,I679982,I680013,I680030,I680047,I680078,I680095,I680135,I680143,I680174,I680191,I680208,I680225,I680256,I680287,I680313,I680335,I680407,I680433,I680441,I680458,I680484,I680492,I680509,I680526,I680543,I680560,I680591,I680608,I680625,I680656,I680673,I680713,I680721,I680752,I680769,I680786,I680803,I680834,I680865,I680891,I680913,I680985,I681011,I681019,I681036,I681062,I681070,I681087,I681104,I681121,I681138,I681169,I681186,I681203,I681234,I681251,I681291,I681299,I681330,I681347,I681364,I681381,I681412,I681443,I681469,I681491,I681563,I681589,I681597,I681614,I681640,I681648,I681665,I681682,I681699,I681716,I681747,I681764,I681781,I681812,I681829,I681869,I681877,I681908,I681925,I681942,I681959,I681990,I682021,I682047,I682069,I682141,I682167,I682175,I682192,I682218,I682226,I682243,I682260,I682277,I682294,I682325,I682342,I682359,I682390,I682407,I682447,I682455,I682486,I682503,I682520,I682537,I682568,I682599,I682625,I682647,I682719,I682745,I682753,I682770,I682796,I682804,I682821,I682838,I682855,I682872,I682711,I682903,I682920,I682937,I682690,I682968,I682985,I682696,I683025,I683033,I682705,I683064,I683081,I683098,I683115,I682708,I683146,I682687,I683177,I683203,I682702,I683225,I682699,I682693,I683297,I683323,I683331,I683348,I683374,I683382,I683399,I683416,I683433,I683450,I683481,I683498,I683515,I683546,I683563,I683603,I683611,I683642,I683659,I683676,I683693,I683724,I683755,I683781,I683803,I683878,I683904,I683912,I683929,I683955,I683963,I683980,I683997,I683864,I684028,I683867,I684059,I684076,I684093,I684110,I684127,I683852,I684158,I683855,I683849,I683846,I684217,I684234,I684260,I683870,I684282,I684308,I684316,I684333,I683861,I684364,I683843,I683858,I684439,I684465,I684473,I684490,I684516,I684524,I684541,I684558,I684589,I684620,I684637,I684654,I684671,I684688,I684719,I684778,I684795,I684821,I684843,I684869,I684877,I684894,I684925,I685000,I703153,I685026,I685034,I703147,I685051,I703165,I685077,I685085,I685102,I703150,I703141,I685119,I685150,I703156,I685181,I703159,I685198,I703162,I685215,I685232,I703144,I685249,I685280,I685339,I703138,I685356,I685382,I685404,I685430,I685438,I685455,I685486,I685561,I685587,I685595,I685612,I685638,I685646,I685663,I685680,I685711,I685742,I685759,I685776,I685793,I685810,I685841,I685900,I685917,I685943,I685965,I685991,I685999,I686016,I686047,I686122,I686148,I686156,I686173,I686199,I686207,I686224,I686241,I686272,I686303,I686320,I686337,I686354,I686371,I686402,I686461,I686478,I686504,I686526,I686552,I686560,I686577,I686608,I686683,I686709,I686717,I686734,I686760,I686768,I686785,I686802,I686833,I686864,I686881,I686898,I686915,I686932,I686963,I687022,I687039,I687065,I687087,I687113,I687121,I687138,I687169,I687244,I687270,I687278,I687295,I687321,I687329,I687346,I687363,I687394,I687425,I687442,I687459,I687476,I687493,I687524,I687583,I687600,I687626,I687648,I687674,I687682,I687699,I687730,I687805,I687831,I687839,I687856,I687882,I687890,I687907,I687924,I687955,I687986,I688003,I688020,I688037,I688054,I688085,I688144,I688161,I688187,I688209,I688235,I688243,I688260,I688291,I688366,I688392,I688400,I688417,I688443,I688451,I688468,I688485,I688516,I688547,I688564,I688581,I688598,I688615,I688646,I688705,I688722,I688748,I688770,I688796,I688804,I688821,I688852,I688927,I688953,I688961,I688978,I689004,I689012,I689029,I689046,I688913,I689077,I688916,I689108,I689125,I689142,I689159,I689176,I688901,I689207,I688904,I688898,I688895,I689266,I689283,I689309,I688919,I689331,I689357,I689365,I689382,I688910,I689413,I688892,I688907,I689488,I689514,I689531,I689539,I689584,I689601,I689618,I689635,I689652,I689669,I689686,I689717,I689734,I689779,I689796,I689813,I689844,I689870,I689878,I689909,I689926,I689943,I689969,I689977,I689994,I690083,I690109,I690126,I690134,I690179,I690196,I690213,I690230,I690247,I690264,I690281,I690312,I690329,I690374,I690391,I690408,I690439,I690465,I690473,I690504,I690521,I690538,I690564,I690572,I690589,I690678,I690704,I690721,I690729,I690774,I690791,I690808,I690825,I690842,I690859,I690876,I690907,I690924,I690969,I690986,I691003,I691034,I691060,I691068,I691099,I691116,I691133,I691159,I691167,I691184,I691273,I691299,I691316,I691324,I691369,I691386,I691403,I691420,I691437,I691454,I691471,I691502,I691519,I691564,I691581,I691598,I691629,I691655,I691663,I691694,I691711,I691728,I691754,I691762,I691779,I691868,I691894,I691911,I691919,I691964,I691981,I691998,I692015,I692032,I692049,I692066,I692097,I692114,I692159,I692176,I692193,I692224,I692250,I692258,I692289,I692306,I692323,I692349,I692357,I692374,I692463,I692489,I692506,I692514,I692559,I692576,I692593,I692610,I692627,I692644,I692661,I692692,I692709,I692754,I692771,I692788,I692819,I692845,I692853,I692884,I692901,I692918,I692944,I692952,I692969,I693058,I693084,I693101,I693109,I693154,I693171,I693188,I693205,I693222,I693239,I693256,I693287,I693304,I693349,I693366,I693383,I693414,I693440,I693448,I693479,I693496,I693513,I693539,I693547,I693564,I693653,I693679,I693696,I693704,I693749,I693766,I693783,I693800,I693817,I693834,I693851,I693882,I693899,I693944,I693961,I693978,I694009,I694035,I694043,I694074,I694091,I694108,I694134,I694142,I694159,I694248,I694274,I694291,I694299,I694344,I694361,I694378,I694395,I694412,I694429,I694446,I694477,I694494,I694539,I694556,I694573,I694604,I694630,I694638,I694669,I694686,I694703,I694729,I694737,I694754,I694843,I694869,I694886,I694894,I694939,I694956,I694973,I694990,I695007,I695024,I695041,I695072,I695089,I695134,I695151,I695168,I695199,I695225,I695233,I695264,I695281,I695298,I695324,I695332,I695349,I695438,I695464,I695481,I695489,I695534,I695551,I695568,I695585,I695602,I695619,I695636,I695667,I695684,I695729,I695746,I695763,I695794,I695820,I695828,I695859,I695876,I695893,I695919,I695927,I695944,I696033,I696059,I696076,I696084,I696129,I696146,I696163,I696180,I696197,I696214,I696231,I696262,I696279,I696324,I696341,I696358,I696389,I696415,I696423,I696454,I696471,I696488,I696514,I696522,I696539,I696628,I696654,I696671,I696679,I696724,I696741,I696758,I696775,I696792,I696809,I696826,I696857,I696874,I696919,I696936,I696953,I696984,I697010,I697018,I697049,I697066,I697083,I697109,I697117,I697134,I697223,I697249,I697266,I697274,I697319,I697336,I697353,I697370,I697387,I697404,I697421,I697452,I697469,I697514,I697531,I697548,I697579,I697605,I697613,I697644,I697661,I697678,I697704,I697712,I697729,I697818,I697844,I697861,I697869,I697914,I697931,I697948,I697965,I697982,I697999,I698016,I698047,I698064,I698109,I698126,I698143,I698174,I698200,I698208,I698239,I698256,I698273,I698299,I698307,I698324,I698413,I698439,I698456,I698464,I698509,I698526,I698543,I698560,I698577,I698594,I698611,I698642,I698659,I698704,I698721,I698738,I698769,I698795,I698803,I698834,I698851,I698868,I698894,I698902,I698919,I699008,I699034,I699051,I699059,I699104,I699121,I699138,I699155,I699172,I699189,I699206,I699237,I699254,I699299,I699316,I699333,I699364,I699390,I699398,I699429,I699446,I699463,I699489,I699497,I699514,I699603,I699629,I699646,I699654,I699699,I699716,I699733,I699750,I699767,I699784,I699801,I699832,I699849,I699894,I699911,I699928,I699959,I699985,I699993,I700024,I700041,I700058,I700084,I700092,I700109,I700198,I700224,I700241,I700249,I700294,I700311,I700328,I700345,I700362,I700379,I700396,I700427,I700444,I700489,I700506,I700523,I700554,I700580,I700588,I700619,I700636,I700653,I700679,I700687,I700704,I700793,I700819,I700836,I700844,I700889,I700906,I700923,I700940,I700957,I700974,I700991,I701022,I701039,I701084,I701101,I701118,I701149,I701175,I701183,I701214,I701231,I701248,I701274,I701282,I701299,I701388,I701414,I701431,I701439,I701484,I701501,I701518,I701535,I701552,I701569,I701586,I701617,I701634,I701679,I701696,I701713,I701744,I701770,I701778,I701809,I701826,I701843,I701869,I701877,I701894,I701983,I702009,I702026,I702034,I702079,I702096,I702113,I702130,I702147,I702164,I702181,I702212,I702229,I702274,I702291,I702308,I702339,I702365,I702373,I702404,I702421,I702438,I702464,I702472,I702489,I702578,I702604,I702621,I702629,I702674,I702691,I702708,I702725,I702742,I702759,I702776,I702807,I702824,I702869,I702886,I702903,I702934,I702960,I702968,I702999,I703016,I703033,I703059,I703067,I703084,I703173,I703199,I703216,I703224,I703269,I703286,I703303,I703320,I703337,I703354,I703371,I703402,I703419,I703464,I703481,I703498,I703529,I703555,I703563,I703594,I703611,I703628,I703654,I703662,I703679,I703768,I703794,I703811,I703819,I703864,I703881,I703898,I703915,I703932,I703949,I703966,I703997,I704014,I704059,I704076,I704093,I704124,I704150,I704158,I704189,I704206,I704223,I704249,I704257,I704274,I704363,I704389,I704406,I704414,I704459,I704476,I704493,I704510,I704527,I704544,I704561,I704592,I704609,I704654,I704671,I704688,I704719,I704745,I704753,I704784,I704801,I704818,I704844,I704852,I704869,I704958,I704984,I705001,I705009,I705054,I705071,I705088,I705105,I705122,I705139,I705156,I705187,I705204,I705249,I705266,I705283,I705314,I705340,I705348,I705379,I705396,I705413,I705439,I705447,I705464,I705553,I705579,I705596,I705604,I705649,I705666,I705683,I705700,I705717,I705734,I705751,I705782,I705799,I705844,I705861,I705878,I705909,I705935,I705943,I705974,I705991,I706008,I706034,I706042,I706059,I706148,I706174,I706191,I706199,I706244,I706261,I706278,I706295,I706312,I706329,I706346,I706377,I706394,I706439,I706456,I706473,I706504,I706530,I706538,I706569,I706586,I706603,I706629,I706637,I706654,I706743,I706769,I706786,I706794,I706839,I706856,I706873,I706890,I706907,I706924,I706941,I706972,I706989,I707034,I707051,I707068,I707099,I707125,I707133,I707164,I707181,I707198,I707224,I707232,I707249,I707338,I707364,I707381,I707389,I707434,I707451,I707468,I707485,I707502,I707519,I707536,I707567,I707584,I707629,I707646,I707663,I707694,I707720,I707728,I707759,I707776,I707793,I707819,I707827,I707844,I707933,I707959,I707976,I707984,I708029,I708046,I708063,I708080,I708097,I708114,I708131,I708162,I708179,I708224,I708241,I708258,I708289,I708315,I708323,I708354,I708371,I708388,I708414,I708422,I708439,I708528,I708554,I708571,I708579,I708624,I708641,I708658,I708675,I708692,I708709,I708726,I708757,I708774,I708819,I708836,I708853,I708884,I708910,I708918,I708949,I708966,I708983,I709009,I709017,I709034,I709123,I709149,I709166,I709174,I709219,I709236,I709253,I709270,I709287,I709304,I709321,I709352,I709369,I709414,I709431,I709448,I709479,I709505,I709513,I709544,I709561,I709578,I709604,I709612,I709629,I709718,I709744,I709761,I709769,I709814,I709831,I709848,I709865,I709882,I709899,I709916,I709947,I709964,I710009,I710026,I710043,I710074,I710100,I710108,I710139,I710156,I710173,I710199,I710207,I710224,I710313,I710339,I710356,I710364,I710409,I710426,I710443,I710460,I710477,I710494,I710511,I710542,I710559,I710604,I710621,I710638,I710669,I710695,I710703,I710734,I710751,I710768,I710794,I710802,I710819,I710908,I710934,I710951,I710959,I711004,I711021,I711038,I711055,I711072,I711089,I711106,I711137,I711154,I711199,I711216,I711233,I711264,I711290,I711298,I711329,I711346,I711363,I711389,I711397,I711414,I711503,I711529,I711546,I711554,I711599,I711616,I711633,I711650,I711667,I711684,I711701,I711732,I711749,I711794,I711811,I711828,I711859,I711885,I711893,I711924,I711941,I711958,I711984,I711992,I712009,I712098,I712124,I712141,I712149,I712194,I712211,I712228,I712245,I712262,I712279,I712296,I712327,I712344,I712389,I712406,I712423,I712454,I712480,I712488,I712519,I712536,I712553,I712579,I712587,I712604,I712693,I712719,I712736,I712744,I712789,I712806,I712823,I712840,I712857,I712874,I712891,I712922,I712939,I712984,I713001,I713018,I713049,I713075,I713083,I713114,I713131,I713148,I713174,I713182,I713199,I713288,I713314,I713331,I713339,I713384,I713401,I713418,I713435,I713452,I713469,I713486,I713517,I713534,I713579,I713596,I713613,I713644,I713670,I713678,I713709,I713726,I713743,I713769,I713777,I713794,I713883,I713909,I713926,I713934,I713979,I713996,I714013,I714030,I714047,I714064,I714081,I714112,I714129,I714174,I714191,I714208,I714239,I714265,I714273,I714304,I714321,I714338,I714364,I714372,I714389,I714478,I714504,I714521,I714529,I714574,I714591,I714608,I714625,I714642,I714659,I714676,I714707,I714724,I714769,I714786,I714803,I714834,I714860,I714868,I714899,I714916,I714933,I714959,I714967,I714984,I715073,I715099,I715116,I715124,I715169,I715186,I715203,I715220,I715237,I715254,I715271,I715302,I715319,I715364,I715381,I715398,I715429,I715455,I715463,I715494,I715511,I715528,I715554,I715562,I715579,I715668,I715694,I715711,I715719,I715764,I715781,I715798,I715815,I715832,I715849,I715866,I715897,I715914,I715959,I715976,I715993,I716024,I716050,I716058,I716089,I716106,I716123,I716149,I716157,I716174,I716263,I716289,I716306,I716314,I716359,I716376,I716393,I716410,I716427,I716444,I716461,I716492,I716509,I716554,I716571,I716588,I716619,I716645,I716653,I716684,I716701,I716718,I716744,I716752,I716769,I716858,I716884,I716901,I716909,I716954,I716971,I716988,I717005,I717022,I717039,I717056,I717087,I717104,I717149,I717166,I717183,I717214,I717240,I717248,I717279,I717296,I717313,I717339,I717347,I717364,I717453,I717479,I717496,I717504,I717549,I717566,I717583,I717600,I717617,I717634,I717651,I717682,I717699,I717744,I717761,I717778,I717809,I717835,I717843,I717874,I717891,I717908,I717934,I717942,I717959,I718048,I718074,I718091,I718099,I718144,I718161,I718178,I718195,I718212,I718229,I718246,I718277,I718294,I718339,I718356,I718373,I718404,I718430,I718438,I718469,I718486,I718503,I718529,I718537,I718554,I718643,I718669,I718686,I718694,I718739,I718756,I718773,I718790,I718807,I718824,I718841,I718872,I718889,I718934,I718951,I718968,I718999,I719025,I719033,I719064,I719081,I719098,I719124,I719132,I719149,I719238,I719264,I719281,I719289,I719334,I719351,I719368,I719385,I719402,I719419,I719436,I719467,I719484,I719529,I719546,I719563,I719594,I719620,I719628,I719659,I719676,I719693,I719719,I719727,I719744,I719833,I719859,I719876,I719884,I719929,I719946,I719963,I719980,I719997,I720014,I720031,I720062,I720079,I720124,I720141,I720158,I720189,I720215,I720223,I720254,I720271,I720288,I720314,I720322,I720339,I720428,I720454,I720471,I720479,I720524,I720541,I720558,I720575,I720592,I720609,I720626,I720657,I720674,I720719,I720736,I720753,I720784,I720810,I720818,I720849,I720866,I720883,I720909,I720917,I720934,I721023,I721049,I721066,I721074,I721119,I721136,I721153,I721170,I721187,I721204,I721221,I721252,I721269,I721314,I721331,I721348,I721379,I721405,I721413,I721444,I721461,I721478,I721504,I721512,I721529,I721618,I721644,I721661,I721669,I721714,I721731,I721748,I721765,I721782,I721799,I721816,I721847,I721864,I721909,I721926,I721943,I721974,I722000,I722008,I722039,I722056,I722073,I722099,I722107,I722124,I722213,I722239,I722256,I722264,I722309,I722326,I722343,I722360,I722377,I722394,I722411,I722442,I722459,I722504,I722521,I722538,I722569,I722595,I722603,I722634,I722651,I722668,I722694,I722702,I722719,I722808,I722834,I722851,I722859,I722904,I722921,I722938,I722955,I722972,I722989,I723006,I723037,I723054,I723099,I723116,I723133,I723164,I723190,I723198,I723229,I723246,I723263,I723289,I723297,I723314,I723403,I723429,I723446,I723454,I723499,I723516,I723533,I723550,I723567,I723584,I723601,I723632,I723649,I723694,I723711,I723728,I723759,I723785,I723793,I723824,I723841,I723858,I723884,I723892,I723909,I723998,I724024,I724041,I724049,I724094,I724111,I724128,I724145,I724162,I724179,I724196,I724227,I724244,I724289,I724306,I724323,I724354,I724380,I724388,I724419,I724436,I724453,I724479,I724487,I724504,I724593,I724619,I724636,I724644,I724689,I724706,I724723,I724740,I724757,I724774,I724791,I724822,I724839,I724884,I724901,I724918,I724949,I724975,I724983,I725014,I725031,I725048,I725074,I725082,I725099,I725188,I725214,I725231,I725239,I725284,I725301,I725318,I725335,I725352,I725369,I725386,I725417,I725434,I725479,I725496,I725513,I725544,I725570,I725578,I725609,I725626,I725643,I725669,I725677,I725694,I725783,I725809,I725826,I725834,I725879,I725896,I725913,I725930,I725947,I725964,I725981,I726012,I726029,I726074,I726091,I726108,I726139,I726165,I726173,I726204,I726221,I726238,I726264,I726272,I726289,I726378,I726404,I726421,I726429,I726474,I726491,I726508,I726525,I726542,I726559,I726576,I726607,I726624,I726669,I726686,I726703,I726734,I726760,I726768,I726799,I726816,I726833,I726859,I726867,I726884,I726973,I726999,I727016,I727024,I727069,I727086,I727103,I727120,I727137,I727154,I727171,I727202,I727219,I727264,I727281,I727298,I727329,I727355,I727363,I727394,I727411,I727428,I727454,I727462,I727479,I727568,I727594,I727611,I727619,I727664,I727681,I727698,I727715,I727732,I727749,I727766,I727797,I727814,I727859,I727876,I727893,I727924,I727950,I727958,I727989,I728006,I728023,I728049,I728057,I728074,I728163,I728189,I728206,I728214,I728259,I728276,I728293,I728310,I728327,I728344,I728361,I728392,I728409,I728454,I728471,I728488,I728519,I728545,I728553,I728584,I728601,I728618,I728644,I728652,I728669,I728758,I728784,I728801,I728809,I728854,I728871,I728888,I728905,I728922,I728939,I728956,I728987,I729004,I729049,I729066,I729083,I729114,I729140,I729148,I729179,I729196,I729213,I729239,I729247,I729264,I729353,I729379,I729396,I729404,I729449,I729466,I729483,I729500,I729517,I729534,I729551,I729582,I729599,I729644,I729661,I729678,I729709,I729735,I729743,I729774,I729791,I729808,I729834,I729842,I729859,I729948,I729974,I729991,I729999,I730044,I730061,I730078,I730095,I730112,I730129,I730146,I730177,I730194,I730239,I730256,I730273,I730304,I730330,I730338,I730369,I730386,I730403,I730429,I730437,I730454,I730543,I730569,I730586,I730594,I730639,I730656,I730673,I730690,I730707,I730724,I730741,I730772,I730789,I730834,I730851,I730868,I730899,I730925,I730933,I730964,I730981,I730998,I731024,I731032,I731049,I731138,I731164,I731181,I731189,I731234,I731251,I731268,I731285,I731302,I731319,I731336,I731367,I731384,I731429,I731446,I731463,I731494,I731520,I731528,I731559,I731576,I731593,I731619,I731627,I731644,I731733,I731759,I731776,I731784,I731829,I731846,I731863,I731880,I731897,I731914,I731931,I731962,I731979,I732024,I732041,I732058,I732089,I732115,I732123,I732154,I732171,I732188,I732214,I732222,I732239;
not I_0 (I2546,I2514);
DFFARX1 I_1 (I399865,I2507,I2546,I2572,);
nand I_2 (I2580,I2572,I399844);
not I_3 (I2597,I2580);
DFFARX1 I_4 (I2597,I2507,I2546,I2538,);
DFFARX1 I_5 (I399853,I2507,I2546,I2637,);
not I_6 (I2645,I2637);
not I_7 (I2662,I399859);
not I_8 (I2679,I399856);
nand I_9 (I2696,I2645,I2679);
nor I_10 (I2713,I2696,I399859);
DFFARX1 I_11 (I2713,I2507,I2546,I2517,);
nor I_12 (I2744,I399856,I399859);
nand I_13 (I2761,I2637,I2744);
nor I_14 (I2778,I399847,I399841);
nor I_15 (I2520,I2696,I399847);
not I_16 (I2809,I399847);
not I_17 (I2826,I399862);
nand I_18 (I2843,I2826,I399844);
nand I_19 (I2860,I2662,I2843);
not I_20 (I2877,I2860);
nor I_21 (I2894,I399862,I399841);
nor I_22 (I2529,I2877,I2894);
nor I_23 (I2925,I399850,I399862);
and I_24 (I2942,I2925,I2778);
nor I_25 (I2959,I2860,I2942);
DFFARX1 I_26 (I2959,I2507,I2546,I2535,);
nor I_27 (I2990,I2580,I2942);
DFFARX1 I_28 (I2990,I2507,I2546,I2532,);
nor I_29 (I3021,I399850,I399841);
DFFARX1 I_30 (I3021,I2507,I2546,I3047,);
nor I_31 (I3055,I3047,I399856);
nand I_32 (I3072,I3055,I2662);
nand I_33 (I2526,I3072,I2761);
nand I_34 (I2523,I3055,I2809);
not I_35 (I3141,I2514);
DFFARX1 I_36 (I567722,I2507,I3141,I3167,);
nand I_37 (I3175,I3167,I567734);
not I_38 (I3192,I3175);
DFFARX1 I_39 (I3192,I2507,I3141,I3133,);
DFFARX1 I_40 (I567719,I2507,I3141,I3232,);
not I_41 (I3240,I3232);
not I_42 (I3257,I567722);
not I_43 (I3274,I567716);
nand I_44 (I3291,I3240,I3274);
nor I_45 (I3308,I3291,I567722);
DFFARX1 I_46 (I3308,I2507,I3141,I3112,);
nor I_47 (I3339,I567716,I567722);
nand I_48 (I3356,I3232,I3339);
nor I_49 (I3373,I567725,I567719);
nor I_50 (I3115,I3291,I567725);
not I_51 (I3404,I567725);
not I_52 (I3421,I567731);
nand I_53 (I3438,I3421,I567716);
nand I_54 (I3455,I3257,I3438);
not I_55 (I3472,I3455);
nor I_56 (I3489,I567731,I567719);
nor I_57 (I3124,I3472,I3489);
nor I_58 (I3520,I567728,I567731);
and I_59 (I3537,I3520,I3373);
nor I_60 (I3554,I3455,I3537);
DFFARX1 I_61 (I3554,I2507,I3141,I3130,);
nor I_62 (I3585,I3175,I3537);
DFFARX1 I_63 (I3585,I2507,I3141,I3127,);
nor I_64 (I3616,I567728,I567737);
DFFARX1 I_65 (I3616,I2507,I3141,I3642,);
nor I_66 (I3650,I3642,I567716);
nand I_67 (I3667,I3650,I3257);
nand I_68 (I3121,I3667,I3356);
nand I_69 (I3118,I3650,I3404);
not I_70 (I3736,I2514);
DFFARX1 I_71 (I628902,I2507,I3736,I3762,);
nand I_72 (I3770,I3762,I628902);
not I_73 (I3787,I3770);
DFFARX1 I_74 (I3787,I2507,I3736,I3728,);
DFFARX1 I_75 (I628917,I2507,I3736,I3827,);
not I_76 (I3835,I3827);
not I_77 (I3852,I628914);
not I_78 (I3869,I628923);
nand I_79 (I3886,I3835,I3869);
nor I_80 (I3903,I3886,I628914);
DFFARX1 I_81 (I3903,I2507,I3736,I3707,);
nor I_82 (I3934,I628923,I628914);
nand I_83 (I3951,I3827,I3934);
nor I_84 (I3968,I628911,I628920);
nor I_85 (I3710,I3886,I628911);
not I_86 (I3999,I628911);
not I_87 (I4016,I628908);
nand I_88 (I4033,I4016,I628899);
nand I_89 (I4050,I3852,I4033);
not I_90 (I4067,I4050);
nor I_91 (I4084,I628908,I628920);
nor I_92 (I3719,I4067,I4084);
nor I_93 (I4115,I628905,I628908);
and I_94 (I4132,I4115,I3968);
nor I_95 (I4149,I4050,I4132);
DFFARX1 I_96 (I4149,I2507,I3736,I3725,);
nor I_97 (I4180,I3770,I4132);
DFFARX1 I_98 (I4180,I2507,I3736,I3722,);
nor I_99 (I4211,I628905,I628899);
DFFARX1 I_100 (I4211,I2507,I3736,I4237,);
nor I_101 (I4245,I4237,I628923);
nand I_102 (I4262,I4245,I3852);
nand I_103 (I3716,I4262,I3951);
nand I_104 (I3713,I4245,I3999);
not I_105 (I4331,I2514);
DFFARX1 I_106 (I577460,I2507,I4331,I4357,);
nand I_107 (I4365,I4357,I577460);
not I_108 (I4382,I4365);
DFFARX1 I_109 (I4382,I2507,I4331,I4323,);
DFFARX1 I_110 (I577475,I2507,I4331,I4422,);
not I_111 (I4430,I4422);
not I_112 (I4447,I577472);
not I_113 (I4464,I577481);
nand I_114 (I4481,I4430,I4464);
nor I_115 (I4498,I4481,I577472);
DFFARX1 I_116 (I4498,I2507,I4331,I4302,);
nor I_117 (I4529,I577481,I577472);
nand I_118 (I4546,I4422,I4529);
nor I_119 (I4563,I577469,I577478);
nor I_120 (I4305,I4481,I577469);
not I_121 (I4594,I577469);
not I_122 (I4611,I577466);
nand I_123 (I4628,I4611,I577457);
nand I_124 (I4645,I4447,I4628);
not I_125 (I4662,I4645);
nor I_126 (I4679,I577466,I577478);
nor I_127 (I4314,I4662,I4679);
nor I_128 (I4710,I577463,I577466);
and I_129 (I4727,I4710,I4563);
nor I_130 (I4744,I4645,I4727);
DFFARX1 I_131 (I4744,I2507,I4331,I4320,);
nor I_132 (I4775,I4365,I4727);
DFFARX1 I_133 (I4775,I2507,I4331,I4317,);
nor I_134 (I4806,I577463,I577457);
DFFARX1 I_135 (I4806,I2507,I4331,I4832,);
nor I_136 (I4840,I4832,I577481);
nand I_137 (I4857,I4840,I4447);
nand I_138 (I4311,I4857,I4546);
nand I_139 (I4308,I4840,I4594);
not I_140 (I4926,I2514);
DFFARX1 I_141 (I457633,I2507,I4926,I4952,);
nand I_142 (I4960,I4952,I457624);
not I_143 (I4977,I4960);
DFFARX1 I_144 (I4977,I2507,I4926,I4918,);
DFFARX1 I_145 (I457630,I2507,I4926,I5017,);
not I_146 (I5025,I5017);
not I_147 (I5042,I457624);
not I_148 (I5059,I457636);
nand I_149 (I5076,I5025,I5059);
nor I_150 (I5093,I5076,I457624);
DFFARX1 I_151 (I5093,I2507,I4926,I4897,);
nor I_152 (I5124,I457636,I457624);
nand I_153 (I5141,I5017,I5124);
nor I_154 (I5158,I457645,I457642);
nor I_155 (I4900,I5076,I457645);
not I_156 (I5189,I457645);
not I_157 (I5206,I457630);
nand I_158 (I5223,I5206,I457627);
nand I_159 (I5240,I5042,I5223);
not I_160 (I5257,I5240);
nor I_161 (I5274,I457630,I457642);
nor I_162 (I4909,I5257,I5274);
nor I_163 (I5305,I457627,I457630);
and I_164 (I5322,I5305,I5158);
nor I_165 (I5339,I5240,I5322);
DFFARX1 I_166 (I5339,I2507,I4926,I4915,);
nor I_167 (I5370,I4960,I5322);
DFFARX1 I_168 (I5370,I2507,I4926,I4912,);
nor I_169 (I5401,I457627,I457639);
DFFARX1 I_170 (I5401,I2507,I4926,I5427,);
nor I_171 (I5435,I5427,I457636);
nand I_172 (I5452,I5435,I5042);
nand I_173 (I4906,I5452,I5141);
nand I_174 (I4903,I5435,I5189);
not I_175 (I5521,I2514);
DFFARX1 I_176 (I456052,I2507,I5521,I5547,);
nand I_177 (I5555,I5547,I456043);
not I_178 (I5572,I5555);
DFFARX1 I_179 (I5572,I2507,I5521,I5513,);
DFFARX1 I_180 (I456049,I2507,I5521,I5612,);
not I_181 (I5620,I5612);
not I_182 (I5637,I456043);
not I_183 (I5654,I456055);
nand I_184 (I5671,I5620,I5654);
nor I_185 (I5688,I5671,I456043);
DFFARX1 I_186 (I5688,I2507,I5521,I5492,);
nor I_187 (I5719,I456055,I456043);
nand I_188 (I5736,I5612,I5719);
nor I_189 (I5753,I456064,I456061);
nor I_190 (I5495,I5671,I456064);
not I_191 (I5784,I456064);
not I_192 (I5801,I456049);
nand I_193 (I5818,I5801,I456046);
nand I_194 (I5835,I5637,I5818);
not I_195 (I5852,I5835);
nor I_196 (I5869,I456049,I456061);
nor I_197 (I5504,I5852,I5869);
nor I_198 (I5900,I456046,I456049);
and I_199 (I5917,I5900,I5753);
nor I_200 (I5934,I5835,I5917);
DFFARX1 I_201 (I5934,I2507,I5521,I5510,);
nor I_202 (I5965,I5555,I5917);
DFFARX1 I_203 (I5965,I2507,I5521,I5507,);
nor I_204 (I5996,I456046,I456058);
DFFARX1 I_205 (I5996,I2507,I5521,I6022,);
nor I_206 (I6030,I6022,I456055);
nand I_207 (I6047,I6030,I5637);
nand I_208 (I5501,I6047,I5736);
nand I_209 (I5498,I6030,I5784);
not I_210 (I6116,I2514);
DFFARX1 I_211 (I489299,I2507,I6116,I6142,);
nand I_212 (I6150,I6142,I489290);
not I_213 (I6167,I6150);
DFFARX1 I_214 (I6167,I2507,I6116,I6108,);
DFFARX1 I_215 (I489293,I2507,I6116,I6207,);
not I_216 (I6215,I6207);
not I_217 (I6232,I489305);
not I_218 (I6249,I489284);
nand I_219 (I6266,I6215,I6249);
nor I_220 (I6283,I6266,I489305);
DFFARX1 I_221 (I6283,I2507,I6116,I6087,);
nor I_222 (I6314,I489284,I489305);
nand I_223 (I6331,I6207,I6314);
nor I_224 (I6348,I489296,I489302);
nor I_225 (I6090,I6266,I489296);
not I_226 (I6379,I489296);
not I_227 (I6396,I489287);
nand I_228 (I6413,I6396,I489278);
nand I_229 (I6430,I6232,I6413);
not I_230 (I6447,I6430);
nor I_231 (I6464,I489287,I489302);
nor I_232 (I6099,I6447,I6464);
nor I_233 (I6495,I489278,I489287);
and I_234 (I6512,I6495,I6348);
nor I_235 (I6529,I6430,I6512);
DFFARX1 I_236 (I6529,I2507,I6116,I6105,);
nor I_237 (I6560,I6150,I6512);
DFFARX1 I_238 (I6560,I2507,I6116,I6102,);
nor I_239 (I6591,I489278,I489281);
DFFARX1 I_240 (I6591,I2507,I6116,I6617,);
nor I_241 (I6625,I6617,I489284);
nand I_242 (I6642,I6625,I6232);
nand I_243 (I6096,I6642,I6331);
nand I_244 (I6093,I6625,I6379);
not I_245 (I6714,I2514);
DFFARX1 I_246 (I501576,I2507,I6714,I6740,);
DFFARX1 I_247 (I6740,I2507,I6714,I6757,);
not I_248 (I6765,I6757);
nand I_249 (I6782,I501552,I501579);
and I_250 (I6799,I6782,I501564);
DFFARX1 I_251 (I6799,I2507,I6714,I6825,);
DFFARX1 I_252 (I6825,I2507,I6714,I6706,);
DFFARX1 I_253 (I6825,I2507,I6714,I6697,);
DFFARX1 I_254 (I501570,I2507,I6714,I6870,);
nand I_255 (I6878,I6870,I501555);
not I_256 (I6895,I6878);
nor I_257 (I6694,I6740,I6895);
DFFARX1 I_258 (I501573,I2507,I6714,I6935,);
not I_259 (I6943,I6935);
nor I_260 (I6700,I6943,I6765);
nand I_261 (I6688,I6943,I6878);
nand I_262 (I6988,I501558,I501561);
and I_263 (I7005,I6988,I501552);
DFFARX1 I_264 (I7005,I2507,I6714,I7031,);
nor I_265 (I7039,I7031,I6740);
DFFARX1 I_266 (I7039,I2507,I6714,I6682,);
not I_267 (I7070,I7031);
nor I_268 (I7087,I501567,I501561);
not I_269 (I7104,I7087);
nor I_270 (I7121,I6878,I7104);
nor I_271 (I7138,I7070,I7121);
DFFARX1 I_272 (I7138,I2507,I6714,I6703,);
nor I_273 (I7169,I7031,I7104);
nor I_274 (I6691,I6895,I7169);
nor I_275 (I6685,I7031,I7087);
not I_276 (I7241,I2514);
DFFARX1 I_277 (I591931,I2507,I7241,I7267,);
DFFARX1 I_278 (I7267,I2507,I7241,I7284,);
not I_279 (I7292,I7284);
nand I_280 (I7309,I591919,I591910);
and I_281 (I7326,I7309,I591907);
DFFARX1 I_282 (I7326,I2507,I7241,I7352,);
DFFARX1 I_283 (I7352,I2507,I7241,I7233,);
DFFARX1 I_284 (I7352,I2507,I7241,I7224,);
DFFARX1 I_285 (I591913,I2507,I7241,I7397,);
nand I_286 (I7405,I7397,I591925);
not I_287 (I7422,I7405);
nor I_288 (I7221,I7267,I7422);
DFFARX1 I_289 (I591922,I2507,I7241,I7462,);
not I_290 (I7470,I7462);
nor I_291 (I7227,I7470,I7292);
nand I_292 (I7215,I7470,I7405);
nand I_293 (I7515,I591916,I591910);
and I_294 (I7532,I7515,I591928);
DFFARX1 I_295 (I7532,I2507,I7241,I7558,);
nor I_296 (I7566,I7558,I7267);
DFFARX1 I_297 (I7566,I2507,I7241,I7209,);
not I_298 (I7597,I7558);
nor I_299 (I7614,I591907,I591910);
not I_300 (I7631,I7614);
nor I_301 (I7648,I7405,I7631);
nor I_302 (I7665,I7597,I7648);
DFFARX1 I_303 (I7665,I2507,I7241,I7230,);
nor I_304 (I7696,I7558,I7631);
nor I_305 (I7218,I7422,I7696);
nor I_306 (I7212,I7558,I7614);
not I_307 (I7768,I2514);
DFFARX1 I_308 (I517080,I2507,I7768,I7794,);
DFFARX1 I_309 (I7794,I2507,I7768,I7811,);
not I_310 (I7819,I7811);
nand I_311 (I7836,I517056,I517083);
and I_312 (I7853,I7836,I517068);
DFFARX1 I_313 (I7853,I2507,I7768,I7879,);
DFFARX1 I_314 (I7879,I2507,I7768,I7760,);
DFFARX1 I_315 (I7879,I2507,I7768,I7751,);
DFFARX1 I_316 (I517074,I2507,I7768,I7924,);
nand I_317 (I7932,I7924,I517059);
not I_318 (I7949,I7932);
nor I_319 (I7748,I7794,I7949);
DFFARX1 I_320 (I517077,I2507,I7768,I7989,);
not I_321 (I7997,I7989);
nor I_322 (I7754,I7997,I7819);
nand I_323 (I7742,I7997,I7932);
nand I_324 (I8042,I517062,I517065);
and I_325 (I8059,I8042,I517056);
DFFARX1 I_326 (I8059,I2507,I7768,I8085,);
nor I_327 (I8093,I8085,I7794);
DFFARX1 I_328 (I8093,I2507,I7768,I7736,);
not I_329 (I8124,I8085);
nor I_330 (I8141,I517071,I517065);
not I_331 (I8158,I8141);
nor I_332 (I8175,I7932,I8158);
nor I_333 (I8192,I8124,I8175);
DFFARX1 I_334 (I8192,I2507,I7768,I7757,);
nor I_335 (I8223,I8085,I8158);
nor I_336 (I7745,I7949,I8223);
nor I_337 (I7739,I8085,I8141);
not I_338 (I8295,I2514);
DFFARX1 I_339 (I225431,I2507,I8295,I8321,);
DFFARX1 I_340 (I8321,I2507,I8295,I8338,);
not I_341 (I8346,I8338);
nand I_342 (I8363,I225428,I225422);
and I_343 (I8380,I8363,I225416);
DFFARX1 I_344 (I8380,I2507,I8295,I8406,);
DFFARX1 I_345 (I8406,I2507,I8295,I8287,);
DFFARX1 I_346 (I8406,I2507,I8295,I8278,);
DFFARX1 I_347 (I225404,I2507,I8295,I8451,);
nand I_348 (I8459,I8451,I225413);
not I_349 (I8476,I8459);
nor I_350 (I8275,I8321,I8476);
DFFARX1 I_351 (I225410,I2507,I8295,I8516,);
not I_352 (I8524,I8516);
nor I_353 (I8281,I8524,I8346);
nand I_354 (I8269,I8524,I8459);
nand I_355 (I8569,I225407,I225425);
and I_356 (I8586,I8569,I225404);
DFFARX1 I_357 (I8586,I2507,I8295,I8612,);
nor I_358 (I8620,I8612,I8321);
DFFARX1 I_359 (I8620,I2507,I8295,I8263,);
not I_360 (I8651,I8612);
nor I_361 (I8668,I225419,I225425);
not I_362 (I8685,I8668);
nor I_363 (I8702,I8459,I8685);
nor I_364 (I8719,I8651,I8702);
DFFARX1 I_365 (I8719,I2507,I8295,I8284,);
nor I_366 (I8750,I8612,I8685);
nor I_367 (I8272,I8476,I8750);
nor I_368 (I8266,I8612,I8668);
not I_369 (I8822,I2514);
DFFARX1 I_370 (I667096,I2507,I8822,I8848,);
DFFARX1 I_371 (I8848,I2507,I8822,I8865,);
not I_372 (I8873,I8865);
nand I_373 (I8890,I667099,I667093);
and I_374 (I8907,I8890,I667102);
DFFARX1 I_375 (I8907,I2507,I8822,I8933,);
DFFARX1 I_376 (I8933,I2507,I8822,I8814,);
DFFARX1 I_377 (I8933,I2507,I8822,I8805,);
DFFARX1 I_378 (I667090,I2507,I8822,I8978,);
nand I_379 (I8986,I8978,I667105);
not I_380 (I9003,I8986);
nor I_381 (I8802,I8848,I9003);
DFFARX1 I_382 (I667081,I2507,I8822,I9043,);
not I_383 (I9051,I9043);
nor I_384 (I8808,I9051,I8873);
nand I_385 (I8796,I9051,I8986);
nand I_386 (I9096,I667084,I667084);
and I_387 (I9113,I9096,I667081);
DFFARX1 I_388 (I9113,I2507,I8822,I9139,);
nor I_389 (I9147,I9139,I8848);
DFFARX1 I_390 (I9147,I2507,I8822,I8790,);
not I_391 (I9178,I9139);
nor I_392 (I9195,I667087,I667084);
not I_393 (I9212,I9195);
nor I_394 (I9229,I8986,I9212);
nor I_395 (I9246,I9178,I9229);
DFFARX1 I_396 (I9246,I2507,I8822,I8811,);
nor I_397 (I9277,I9139,I9212);
nor I_398 (I8799,I9003,I9277);
nor I_399 (I8793,I9139,I9195);
not I_400 (I9349,I2514);
DFFARX1 I_401 (I646885,I2507,I9349,I9375,);
DFFARX1 I_402 (I9375,I2507,I9349,I9392,);
not I_403 (I9400,I9392);
nand I_404 (I9417,I646903,I646897);
and I_405 (I9434,I9417,I646906);
DFFARX1 I_406 (I9434,I2507,I9349,I9460,);
DFFARX1 I_407 (I9460,I2507,I9349,I9341,);
DFFARX1 I_408 (I9460,I2507,I9349,I9332,);
DFFARX1 I_409 (I646891,I2507,I9349,I9505,);
nand I_410 (I9513,I9505,I646900);
not I_411 (I9530,I9513);
nor I_412 (I9329,I9375,I9530);
DFFARX1 I_413 (I646888,I2507,I9349,I9570,);
not I_414 (I9578,I9570);
nor I_415 (I9335,I9578,I9400);
nand I_416 (I9323,I9578,I9513);
nand I_417 (I9623,I646909,I646894);
and I_418 (I9640,I9623,I646888);
DFFARX1 I_419 (I9640,I2507,I9349,I9666,);
nor I_420 (I9674,I9666,I9375);
DFFARX1 I_421 (I9674,I2507,I9349,I9317,);
not I_422 (I9705,I9666);
nor I_423 (I9722,I646885,I646894);
not I_424 (I9739,I9722);
nor I_425 (I9756,I9513,I9739);
nor I_426 (I9773,I9705,I9756);
DFFARX1 I_427 (I9773,I2507,I9349,I9338,);
nor I_428 (I9804,I9666,I9739);
nor I_429 (I9326,I9530,I9804);
nor I_430 (I9320,I9666,I9722);
not I_431 (I9876,I2514);
DFFARX1 I_432 (I140155,I2507,I9876,I9902,);
DFFARX1 I_433 (I9902,I2507,I9876,I9919,);
not I_434 (I9927,I9919);
nand I_435 (I9944,I140173,I140158);
and I_436 (I9961,I9944,I140161);
DFFARX1 I_437 (I9961,I2507,I9876,I9987,);
DFFARX1 I_438 (I9987,I2507,I9876,I9868,);
DFFARX1 I_439 (I9987,I2507,I9876,I9859,);
DFFARX1 I_440 (I140149,I2507,I9876,I10032,);
nand I_441 (I10040,I10032,I140152);
not I_442 (I10057,I10040);
nor I_443 (I9856,I9902,I10057);
DFFARX1 I_444 (I140164,I2507,I9876,I10097,);
not I_445 (I10105,I10097);
nor I_446 (I9862,I10105,I9927);
nand I_447 (I9850,I10105,I10040);
nand I_448 (I10150,I140170,I140167);
and I_449 (I10167,I10150,I140152);
DFFARX1 I_450 (I10167,I2507,I9876,I10193,);
nor I_451 (I10201,I10193,I9902);
DFFARX1 I_452 (I10201,I2507,I9876,I9844,);
not I_453 (I10232,I10193);
nor I_454 (I10249,I140149,I140167);
not I_455 (I10266,I10249);
nor I_456 (I10283,I10040,I10266);
nor I_457 (I10300,I10232,I10283);
DFFARX1 I_458 (I10300,I2507,I9876,I9865,);
nor I_459 (I10331,I10193,I10266);
nor I_460 (I9853,I10057,I10331);
nor I_461 (I9847,I10193,I10249);
not I_462 (I10403,I2514);
DFFARX1 I_463 (I722773,I2507,I10403,I10429,);
DFFARX1 I_464 (I10429,I2507,I10403,I10446,);
not I_465 (I10454,I10446);
nand I_466 (I10471,I722776,I722782);
and I_467 (I10488,I10471,I722791);
DFFARX1 I_468 (I10488,I2507,I10403,I10514,);
DFFARX1 I_469 (I10514,I2507,I10403,I10395,);
DFFARX1 I_470 (I10514,I2507,I10403,I10386,);
DFFARX1 I_471 (I722794,I2507,I10403,I10559,);
nand I_472 (I10567,I10559,I722785);
not I_473 (I10584,I10567);
nor I_474 (I10383,I10429,I10584);
DFFARX1 I_475 (I722773,I2507,I10403,I10624,);
not I_476 (I10632,I10624);
nor I_477 (I10389,I10632,I10454);
nand I_478 (I10377,I10632,I10567);
nand I_479 (I10677,I722800,I722779);
and I_480 (I10694,I10677,I722788);
DFFARX1 I_481 (I10694,I2507,I10403,I10720,);
nor I_482 (I10728,I10720,I10429);
DFFARX1 I_483 (I10728,I2507,I10403,I10371,);
not I_484 (I10759,I10720);
nor I_485 (I10776,I722797,I722779);
not I_486 (I10793,I10776);
nor I_487 (I10810,I10567,I10793);
nor I_488 (I10827,I10759,I10810);
DFFARX1 I_489 (I10827,I2507,I10403,I10392,);
nor I_490 (I10858,I10720,I10793);
nor I_491 (I10380,I10584,I10858);
nor I_492 (I10374,I10720,I10776);
not I_493 (I10930,I2514);
DFFARX1 I_494 (I589041,I2507,I10930,I10956,);
DFFARX1 I_495 (I10956,I2507,I10930,I10973,);
not I_496 (I10981,I10973);
nand I_497 (I10998,I589029,I589020);
and I_498 (I11015,I10998,I589017);
DFFARX1 I_499 (I11015,I2507,I10930,I11041,);
DFFARX1 I_500 (I11041,I2507,I10930,I10922,);
DFFARX1 I_501 (I11041,I2507,I10930,I10913,);
DFFARX1 I_502 (I589023,I2507,I10930,I11086,);
nand I_503 (I11094,I11086,I589035);
not I_504 (I11111,I11094);
nor I_505 (I10910,I10956,I11111);
DFFARX1 I_506 (I589032,I2507,I10930,I11151,);
not I_507 (I11159,I11151);
nor I_508 (I10916,I11159,I10981);
nand I_509 (I10904,I11159,I11094);
nand I_510 (I11204,I589026,I589020);
and I_511 (I11221,I11204,I589038);
DFFARX1 I_512 (I11221,I2507,I10930,I11247,);
nor I_513 (I11255,I11247,I10956);
DFFARX1 I_514 (I11255,I2507,I10930,I10898,);
not I_515 (I11286,I11247);
nor I_516 (I11303,I589017,I589020);
not I_517 (I11320,I11303);
nor I_518 (I11337,I11094,I11320);
nor I_519 (I11354,I11286,I11337);
DFFARX1 I_520 (I11354,I2507,I10930,I10919,);
nor I_521 (I11385,I11247,I11320);
nor I_522 (I10907,I11111,I11385);
nor I_523 (I10901,I11247,I11303);
not I_524 (I11457,I2514);
DFFARX1 I_525 (I1724,I2507,I11457,I11483,);
DFFARX1 I_526 (I11483,I2507,I11457,I11500,);
not I_527 (I11508,I11500);
nand I_528 (I11525,I1604,I1732);
and I_529 (I11542,I11525,I1956);
DFFARX1 I_530 (I11542,I2507,I11457,I11568,);
DFFARX1 I_531 (I11568,I2507,I11457,I11449,);
DFFARX1 I_532 (I11568,I2507,I11457,I11440,);
DFFARX1 I_533 (I1636,I2507,I11457,I11613,);
nand I_534 (I11621,I11613,I2132);
not I_535 (I11638,I11621);
nor I_536 (I11437,I11483,I11638);
DFFARX1 I_537 (I1588,I2507,I11457,I11678,);
not I_538 (I11686,I11678);
nor I_539 (I11443,I11686,I11508);
nand I_540 (I11431,I11686,I11621);
nand I_541 (I11731,I1908,I1524);
and I_542 (I11748,I11731,I2020);
DFFARX1 I_543 (I11748,I2507,I11457,I11774,);
nor I_544 (I11782,I11774,I11483);
DFFARX1 I_545 (I11782,I2507,I11457,I11425,);
not I_546 (I11813,I11774);
nor I_547 (I11830,I1652,I1524);
not I_548 (I11847,I11830);
nor I_549 (I11864,I11621,I11847);
nor I_550 (I11881,I11813,I11864);
DFFARX1 I_551 (I11881,I2507,I11457,I11446,);
nor I_552 (I11912,I11774,I11847);
nor I_553 (I11434,I11638,I11912);
nor I_554 (I11428,I11774,I11830);
not I_555 (I11984,I2514);
DFFARX1 I_556 (I266136,I2507,I11984,I12010,);
DFFARX1 I_557 (I12010,I2507,I11984,I12027,);
not I_558 (I12035,I12027);
nand I_559 (I12052,I266136,I266139);
and I_560 (I12069,I12052,I266160);
DFFARX1 I_561 (I12069,I2507,I11984,I12095,);
DFFARX1 I_562 (I12095,I2507,I11984,I11976,);
DFFARX1 I_563 (I12095,I2507,I11984,I11967,);
DFFARX1 I_564 (I266148,I2507,I11984,I12140,);
nand I_565 (I12148,I12140,I266151);
not I_566 (I12165,I12148);
nor I_567 (I11964,I12010,I12165);
DFFARX1 I_568 (I266157,I2507,I11984,I12205,);
not I_569 (I12213,I12205);
nor I_570 (I11970,I12213,I12035);
nand I_571 (I11958,I12213,I12148);
nand I_572 (I12258,I266154,I266142);
and I_573 (I12275,I12258,I266145);
DFFARX1 I_574 (I12275,I2507,I11984,I12301,);
nor I_575 (I12309,I12301,I12010);
DFFARX1 I_576 (I12309,I2507,I11984,I11952,);
not I_577 (I12340,I12301);
nor I_578 (I12357,I266163,I266142);
not I_579 (I12374,I12357);
nor I_580 (I12391,I12148,I12374);
nor I_581 (I12408,I12340,I12391);
DFFARX1 I_582 (I12408,I2507,I11984,I11973,);
nor I_583 (I12439,I12301,I12374);
nor I_584 (I11961,I12165,I12439);
nor I_585 (I11955,I12301,I12357);
not I_586 (I12511,I2514);
DFFARX1 I_587 (I585573,I2507,I12511,I12537,);
DFFARX1 I_588 (I12537,I2507,I12511,I12554,);
not I_589 (I12562,I12554);
nand I_590 (I12579,I585561,I585552);
and I_591 (I12596,I12579,I585549);
DFFARX1 I_592 (I12596,I2507,I12511,I12622,);
DFFARX1 I_593 (I12622,I2507,I12511,I12503,);
DFFARX1 I_594 (I12622,I2507,I12511,I12494,);
DFFARX1 I_595 (I585555,I2507,I12511,I12667,);
nand I_596 (I12675,I12667,I585567);
not I_597 (I12692,I12675);
nor I_598 (I12491,I12537,I12692);
DFFARX1 I_599 (I585564,I2507,I12511,I12732,);
not I_600 (I12740,I12732);
nor I_601 (I12497,I12740,I12562);
nand I_602 (I12485,I12740,I12675);
nand I_603 (I12785,I585558,I585552);
and I_604 (I12802,I12785,I585570);
DFFARX1 I_605 (I12802,I2507,I12511,I12828,);
nor I_606 (I12836,I12828,I12537);
DFFARX1 I_607 (I12836,I2507,I12511,I12479,);
not I_608 (I12867,I12828);
nor I_609 (I12884,I585549,I585552);
not I_610 (I12901,I12884);
nor I_611 (I12918,I12675,I12901);
nor I_612 (I12935,I12867,I12918);
DFFARX1 I_613 (I12935,I2507,I12511,I12500,);
nor I_614 (I12966,I12828,I12901);
nor I_615 (I12488,I12692,I12966);
nor I_616 (I12482,I12828,I12884);
not I_617 (I13038,I2514);
DFFARX1 I_618 (I641445,I2507,I13038,I13064,);
DFFARX1 I_619 (I13064,I2507,I13038,I13081,);
not I_620 (I13089,I13081);
nand I_621 (I13106,I641463,I641457);
and I_622 (I13123,I13106,I641466);
DFFARX1 I_623 (I13123,I2507,I13038,I13149,);
DFFARX1 I_624 (I13149,I2507,I13038,I13030,);
DFFARX1 I_625 (I13149,I2507,I13038,I13021,);
DFFARX1 I_626 (I641451,I2507,I13038,I13194,);
nand I_627 (I13202,I13194,I641460);
not I_628 (I13219,I13202);
nor I_629 (I13018,I13064,I13219);
DFFARX1 I_630 (I641448,I2507,I13038,I13259,);
not I_631 (I13267,I13259);
nor I_632 (I13024,I13267,I13089);
nand I_633 (I13012,I13267,I13202);
nand I_634 (I13312,I641469,I641454);
and I_635 (I13329,I13312,I641448);
DFFARX1 I_636 (I13329,I2507,I13038,I13355,);
nor I_637 (I13363,I13355,I13064);
DFFARX1 I_638 (I13363,I2507,I13038,I13006,);
not I_639 (I13394,I13355);
nor I_640 (I13411,I641445,I641454);
not I_641 (I13428,I13411);
nor I_642 (I13445,I13202,I13428);
nor I_643 (I13462,I13394,I13445);
DFFARX1 I_644 (I13462,I2507,I13038,I13027,);
nor I_645 (I13493,I13355,I13428);
nor I_646 (I13015,I13219,I13493);
nor I_647 (I13009,I13355,I13411);
not I_648 (I13565,I2514);
DFFARX1 I_649 (I261240,I2507,I13565,I13591,);
DFFARX1 I_650 (I13591,I2507,I13565,I13608,);
not I_651 (I13616,I13608);
nand I_652 (I13633,I261240,I261243);
and I_653 (I13650,I13633,I261264);
DFFARX1 I_654 (I13650,I2507,I13565,I13676,);
DFFARX1 I_655 (I13676,I2507,I13565,I13557,);
DFFARX1 I_656 (I13676,I2507,I13565,I13548,);
DFFARX1 I_657 (I261252,I2507,I13565,I13721,);
nand I_658 (I13729,I13721,I261255);
not I_659 (I13746,I13729);
nor I_660 (I13545,I13591,I13746);
DFFARX1 I_661 (I261261,I2507,I13565,I13786,);
not I_662 (I13794,I13786);
nor I_663 (I13551,I13794,I13616);
nand I_664 (I13539,I13794,I13729);
nand I_665 (I13839,I261258,I261246);
and I_666 (I13856,I13839,I261249);
DFFARX1 I_667 (I13856,I2507,I13565,I13882,);
nor I_668 (I13890,I13882,I13591);
DFFARX1 I_669 (I13890,I2507,I13565,I13533,);
not I_670 (I13921,I13882);
nor I_671 (I13938,I261267,I261246);
not I_672 (I13955,I13938);
nor I_673 (I13972,I13729,I13955);
nor I_674 (I13989,I13921,I13972);
DFFARX1 I_675 (I13989,I2507,I13565,I13554,);
nor I_676 (I14020,I13882,I13955);
nor I_677 (I13542,I13746,I14020);
nor I_678 (I13536,I13882,I13938);
not I_679 (I14092,I2514);
DFFARX1 I_680 (I711468,I2507,I14092,I14118,);
DFFARX1 I_681 (I14118,I2507,I14092,I14135,);
not I_682 (I14143,I14135);
nand I_683 (I14160,I711471,I711477);
and I_684 (I14177,I14160,I711486);
DFFARX1 I_685 (I14177,I2507,I14092,I14203,);
DFFARX1 I_686 (I14203,I2507,I14092,I14084,);
DFFARX1 I_687 (I14203,I2507,I14092,I14075,);
DFFARX1 I_688 (I711489,I2507,I14092,I14248,);
nand I_689 (I14256,I14248,I711480);
not I_690 (I14273,I14256);
nor I_691 (I14072,I14118,I14273);
DFFARX1 I_692 (I711468,I2507,I14092,I14313,);
not I_693 (I14321,I14313);
nor I_694 (I14078,I14321,I14143);
nand I_695 (I14066,I14321,I14256);
nand I_696 (I14366,I711495,I711474);
and I_697 (I14383,I14366,I711483);
DFFARX1 I_698 (I14383,I2507,I14092,I14409,);
nor I_699 (I14417,I14409,I14118);
DFFARX1 I_700 (I14417,I2507,I14092,I14060,);
not I_701 (I14448,I14409);
nor I_702 (I14465,I711492,I711474);
not I_703 (I14482,I14465);
nor I_704 (I14499,I14256,I14482);
nor I_705 (I14516,I14448,I14499);
DFFARX1 I_706 (I14516,I2507,I14092,I14081,);
nor I_707 (I14547,I14409,I14482);
nor I_708 (I14069,I14273,I14547);
nor I_709 (I14063,I14409,I14465);
not I_710 (I14619,I2514);
DFFARX1 I_711 (I220688,I2507,I14619,I14645,);
DFFARX1 I_712 (I14645,I2507,I14619,I14662,);
not I_713 (I14670,I14662);
nand I_714 (I14687,I220685,I220679);
and I_715 (I14704,I14687,I220673);
DFFARX1 I_716 (I14704,I2507,I14619,I14730,);
DFFARX1 I_717 (I14730,I2507,I14619,I14611,);
DFFARX1 I_718 (I14730,I2507,I14619,I14602,);
DFFARX1 I_719 (I220661,I2507,I14619,I14775,);
nand I_720 (I14783,I14775,I220670);
not I_721 (I14800,I14783);
nor I_722 (I14599,I14645,I14800);
DFFARX1 I_723 (I220667,I2507,I14619,I14840,);
not I_724 (I14848,I14840);
nor I_725 (I14605,I14848,I14670);
nand I_726 (I14593,I14848,I14783);
nand I_727 (I14893,I220664,I220682);
and I_728 (I14910,I14893,I220661);
DFFARX1 I_729 (I14910,I2507,I14619,I14936,);
nor I_730 (I14944,I14936,I14645);
DFFARX1 I_731 (I14944,I2507,I14619,I14587,);
not I_732 (I14975,I14936);
nor I_733 (I14992,I220676,I220682);
not I_734 (I15009,I14992);
nor I_735 (I15026,I14783,I15009);
nor I_736 (I15043,I14975,I15026);
DFFARX1 I_737 (I15043,I2507,I14619,I14608,);
nor I_738 (I15074,I14936,I15009);
nor I_739 (I14596,I14800,I15074);
nor I_740 (I14590,I14936,I14992);
not I_741 (I15146,I2514);
DFFARX1 I_742 (I195392,I2507,I15146,I15172,);
DFFARX1 I_743 (I15172,I2507,I15146,I15189,);
not I_744 (I15197,I15189);
nand I_745 (I15214,I195389,I195383);
and I_746 (I15231,I15214,I195377);
DFFARX1 I_747 (I15231,I2507,I15146,I15257,);
DFFARX1 I_748 (I15257,I2507,I15146,I15138,);
DFFARX1 I_749 (I15257,I2507,I15146,I15129,);
DFFARX1 I_750 (I195365,I2507,I15146,I15302,);
nand I_751 (I15310,I15302,I195374);
not I_752 (I15327,I15310);
nor I_753 (I15126,I15172,I15327);
DFFARX1 I_754 (I195371,I2507,I15146,I15367,);
not I_755 (I15375,I15367);
nor I_756 (I15132,I15375,I15197);
nand I_757 (I15120,I15375,I15310);
nand I_758 (I15420,I195368,I195386);
and I_759 (I15437,I15420,I195365);
DFFARX1 I_760 (I15437,I2507,I15146,I15463,);
nor I_761 (I15471,I15463,I15172);
DFFARX1 I_762 (I15471,I2507,I15146,I15114,);
not I_763 (I15502,I15463);
nor I_764 (I15519,I195380,I195386);
not I_765 (I15536,I15519);
nor I_766 (I15553,I15310,I15536);
nor I_767 (I15570,I15502,I15553);
DFFARX1 I_768 (I15570,I2507,I15146,I15135,);
nor I_769 (I15601,I15463,I15536);
nor I_770 (I15123,I15327,I15601);
nor I_771 (I15117,I15463,I15519);
not I_772 (I15673,I2514);
DFFARX1 I_773 (I594243,I2507,I15673,I15699,);
DFFARX1 I_774 (I15699,I2507,I15673,I15716,);
not I_775 (I15724,I15716);
nand I_776 (I15741,I594231,I594222);
and I_777 (I15758,I15741,I594219);
DFFARX1 I_778 (I15758,I2507,I15673,I15784,);
DFFARX1 I_779 (I15784,I2507,I15673,I15665,);
DFFARX1 I_780 (I15784,I2507,I15673,I15656,);
DFFARX1 I_781 (I594225,I2507,I15673,I15829,);
nand I_782 (I15837,I15829,I594237);
not I_783 (I15854,I15837);
nor I_784 (I15653,I15699,I15854);
DFFARX1 I_785 (I594234,I2507,I15673,I15894,);
not I_786 (I15902,I15894);
nor I_787 (I15659,I15902,I15724);
nand I_788 (I15647,I15902,I15837);
nand I_789 (I15947,I594228,I594222);
and I_790 (I15964,I15947,I594240);
DFFARX1 I_791 (I15964,I2507,I15673,I15990,);
nor I_792 (I15998,I15990,I15699);
DFFARX1 I_793 (I15998,I2507,I15673,I15641,);
not I_794 (I16029,I15990);
nor I_795 (I16046,I594219,I594222);
not I_796 (I16063,I16046);
nor I_797 (I16080,I15837,I16063);
nor I_798 (I16097,I16029,I16080);
DFFARX1 I_799 (I16097,I2507,I15673,I15662,);
nor I_800 (I16128,I15990,I16063);
nor I_801 (I15650,I15854,I16128);
nor I_802 (I15644,I15990,I16046);
not I_803 (I16200,I2514);
DFFARX1 I_804 (I44102,I2507,I16200,I16226,);
DFFARX1 I_805 (I16226,I2507,I16200,I16243,);
not I_806 (I16251,I16243);
nand I_807 (I16268,I44102,I44117);
and I_808 (I16285,I16268,I44120);
DFFARX1 I_809 (I16285,I2507,I16200,I16311,);
DFFARX1 I_810 (I16311,I2507,I16200,I16192,);
DFFARX1 I_811 (I16311,I2507,I16200,I16183,);
DFFARX1 I_812 (I44114,I2507,I16200,I16356,);
nand I_813 (I16364,I16356,I44123);
not I_814 (I16381,I16364);
nor I_815 (I16180,I16226,I16381);
DFFARX1 I_816 (I44099,I2507,I16200,I16421,);
not I_817 (I16429,I16421);
nor I_818 (I16186,I16429,I16251);
nand I_819 (I16174,I16429,I16364);
nand I_820 (I16474,I44099,I44105);
and I_821 (I16491,I16474,I44108);
DFFARX1 I_822 (I16491,I2507,I16200,I16517,);
nor I_823 (I16525,I16517,I16226);
DFFARX1 I_824 (I16525,I2507,I16200,I16168,);
not I_825 (I16556,I16517);
nor I_826 (I16573,I44111,I44105);
not I_827 (I16590,I16573);
nor I_828 (I16607,I16364,I16590);
nor I_829 (I16624,I16556,I16607);
DFFARX1 I_830 (I16624,I2507,I16200,I16189,);
nor I_831 (I16655,I16517,I16590);
nor I_832 (I16177,I16381,I16655);
nor I_833 (I16171,I16517,I16573);
not I_834 (I16727,I2514);
DFFARX1 I_835 (I364011,I2507,I16727,I16753,);
DFFARX1 I_836 (I16753,I2507,I16727,I16770,);
not I_837 (I16778,I16770);
nand I_838 (I16795,I364026,I364029);
and I_839 (I16812,I16795,I364008);
DFFARX1 I_840 (I16812,I2507,I16727,I16838,);
DFFARX1 I_841 (I16838,I2507,I16727,I16719,);
DFFARX1 I_842 (I16838,I2507,I16727,I16710,);
DFFARX1 I_843 (I364014,I2507,I16727,I16883,);
nand I_844 (I16891,I16883,I364020);
not I_845 (I16908,I16891);
nor I_846 (I16707,I16753,I16908);
DFFARX1 I_847 (I364008,I2507,I16727,I16948,);
not I_848 (I16956,I16948);
nor I_849 (I16713,I16956,I16778);
nand I_850 (I16701,I16956,I16891);
nand I_851 (I17001,I364023,I364005);
and I_852 (I17018,I17001,I364017);
DFFARX1 I_853 (I17018,I2507,I16727,I17044,);
nor I_854 (I17052,I17044,I16753);
DFFARX1 I_855 (I17052,I2507,I16727,I16695,);
not I_856 (I17083,I17044);
nor I_857 (I17100,I364005,I364005);
not I_858 (I17117,I17100);
nor I_859 (I17134,I16891,I17117);
nor I_860 (I17151,I17083,I17134);
DFFARX1 I_861 (I17151,I2507,I16727,I16716,);
nor I_862 (I17182,I17044,I17117);
nor I_863 (I16704,I16908,I17182);
nor I_864 (I16698,I17044,I17100);
not I_865 (I17254,I2514);
DFFARX1 I_866 (I580949,I2507,I17254,I17280,);
DFFARX1 I_867 (I17280,I2507,I17254,I17297,);
not I_868 (I17305,I17297);
nand I_869 (I17322,I580937,I580928);
and I_870 (I17339,I17322,I580925);
DFFARX1 I_871 (I17339,I2507,I17254,I17365,);
DFFARX1 I_872 (I17365,I2507,I17254,I17246,);
DFFARX1 I_873 (I17365,I2507,I17254,I17237,);
DFFARX1 I_874 (I580931,I2507,I17254,I17410,);
nand I_875 (I17418,I17410,I580943);
not I_876 (I17435,I17418);
nor I_877 (I17234,I17280,I17435);
DFFARX1 I_878 (I580940,I2507,I17254,I17475,);
not I_879 (I17483,I17475);
nor I_880 (I17240,I17483,I17305);
nand I_881 (I17228,I17483,I17418);
nand I_882 (I17528,I580934,I580928);
and I_883 (I17545,I17528,I580946);
DFFARX1 I_884 (I17545,I2507,I17254,I17571,);
nor I_885 (I17579,I17571,I17280);
DFFARX1 I_886 (I17579,I2507,I17254,I17222,);
not I_887 (I17610,I17571);
nor I_888 (I17627,I580925,I580928);
not I_889 (I17644,I17627);
nor I_890 (I17661,I17418,I17644);
nor I_891 (I17678,I17610,I17661);
DFFARX1 I_892 (I17678,I2507,I17254,I17243,);
nor I_893 (I17709,I17571,I17644);
nor I_894 (I17231,I17435,I17709);
nor I_895 (I17225,I17571,I17627);
not I_896 (I17781,I2514);
DFFARX1 I_897 (I679812,I2507,I17781,I17807,);
DFFARX1 I_898 (I17807,I2507,I17781,I17824,);
not I_899 (I17832,I17824);
nand I_900 (I17849,I679815,I679809);
and I_901 (I17866,I17849,I679818);
DFFARX1 I_902 (I17866,I2507,I17781,I17892,);
DFFARX1 I_903 (I17892,I2507,I17781,I17773,);
DFFARX1 I_904 (I17892,I2507,I17781,I17764,);
DFFARX1 I_905 (I679806,I2507,I17781,I17937,);
nand I_906 (I17945,I17937,I679821);
not I_907 (I17962,I17945);
nor I_908 (I17761,I17807,I17962);
DFFARX1 I_909 (I679797,I2507,I17781,I18002,);
not I_910 (I18010,I18002);
nor I_911 (I17767,I18010,I17832);
nand I_912 (I17755,I18010,I17945);
nand I_913 (I18055,I679800,I679800);
and I_914 (I18072,I18055,I679797);
DFFARX1 I_915 (I18072,I2507,I17781,I18098,);
nor I_916 (I18106,I18098,I17807);
DFFARX1 I_917 (I18106,I2507,I17781,I17749,);
not I_918 (I18137,I18098);
nor I_919 (I18154,I679803,I679800);
not I_920 (I18171,I18154);
nor I_921 (I18188,I17945,I18171);
nor I_922 (I18205,I18137,I18188);
DFFARX1 I_923 (I18205,I2507,I17781,I17770,);
nor I_924 (I18236,I18098,I18171);
nor I_925 (I17758,I17962,I18236);
nor I_926 (I17752,I18098,I18154);
not I_927 (I18308,I2514);
DFFARX1 I_928 (I704923,I2507,I18308,I18334,);
DFFARX1 I_929 (I18334,I2507,I18308,I18351,);
not I_930 (I18359,I18351);
nand I_931 (I18376,I704926,I704932);
and I_932 (I18393,I18376,I704941);
DFFARX1 I_933 (I18393,I2507,I18308,I18419,);
DFFARX1 I_934 (I18419,I2507,I18308,I18300,);
DFFARX1 I_935 (I18419,I2507,I18308,I18291,);
DFFARX1 I_936 (I704944,I2507,I18308,I18464,);
nand I_937 (I18472,I18464,I704935);
not I_938 (I18489,I18472);
nor I_939 (I18288,I18334,I18489);
DFFARX1 I_940 (I704923,I2507,I18308,I18529,);
not I_941 (I18537,I18529);
nor I_942 (I18294,I18537,I18359);
nand I_943 (I18282,I18537,I18472);
nand I_944 (I18582,I704950,I704929);
and I_945 (I18599,I18582,I704938);
DFFARX1 I_946 (I18599,I2507,I18308,I18625,);
nor I_947 (I18633,I18625,I18334);
DFFARX1 I_948 (I18633,I2507,I18308,I18276,);
not I_949 (I18664,I18625);
nor I_950 (I18681,I704947,I704929);
not I_951 (I18698,I18681);
nor I_952 (I18715,I18472,I18698);
nor I_953 (I18732,I18664,I18715);
DFFARX1 I_954 (I18732,I2507,I18308,I18297,);
nor I_955 (I18763,I18625,I18698);
nor I_956 (I18285,I18489,I18763);
nor I_957 (I18279,I18625,I18681);
not I_958 (I18835,I2514);
DFFARX1 I_959 (I287922,I2507,I18835,I18861,);
DFFARX1 I_960 (I18861,I2507,I18835,I18878,);
not I_961 (I18886,I18878);
nand I_962 (I18903,I287928,I287916);
and I_963 (I18920,I18903,I287913);
DFFARX1 I_964 (I18920,I2507,I18835,I18946,);
DFFARX1 I_965 (I18946,I2507,I18835,I18827,);
DFFARX1 I_966 (I18946,I2507,I18835,I18818,);
DFFARX1 I_967 (I287925,I2507,I18835,I18991,);
nand I_968 (I18999,I18991,I287919);
not I_969 (I19016,I18999);
nor I_970 (I18815,I18861,I19016);
DFFARX1 I_971 (I287937,I2507,I18835,I19056,);
not I_972 (I19064,I19056);
nor I_973 (I18821,I19064,I18886);
nand I_974 (I18809,I19064,I18999);
nand I_975 (I19109,I287931,I287934);
and I_976 (I19126,I19109,I287916);
DFFARX1 I_977 (I19126,I2507,I18835,I19152,);
nor I_978 (I19160,I19152,I18861);
DFFARX1 I_979 (I19160,I2507,I18835,I18803,);
not I_980 (I19191,I19152);
nor I_981 (I19208,I287913,I287934);
not I_982 (I19225,I19208);
nor I_983 (I19242,I18999,I19225);
nor I_984 (I19259,I19191,I19242);
DFFARX1 I_985 (I19259,I2507,I18835,I18824,);
nor I_986 (I19290,I19152,I19225);
nor I_987 (I18812,I19016,I19290);
nor I_988 (I18806,I19152,I19208);
not I_989 (I19362,I2514);
DFFARX1 I_990 (I38305,I2507,I19362,I19388,);
DFFARX1 I_991 (I19388,I2507,I19362,I19405,);
not I_992 (I19413,I19405);
nand I_993 (I19430,I38305,I38320);
and I_994 (I19447,I19430,I38323);
DFFARX1 I_995 (I19447,I2507,I19362,I19473,);
DFFARX1 I_996 (I19473,I2507,I19362,I19354,);
DFFARX1 I_997 (I19473,I2507,I19362,I19345,);
DFFARX1 I_998 (I38317,I2507,I19362,I19518,);
nand I_999 (I19526,I19518,I38326);
not I_1000 (I19543,I19526);
nor I_1001 (I19342,I19388,I19543);
DFFARX1 I_1002 (I38302,I2507,I19362,I19583,);
not I_1003 (I19591,I19583);
nor I_1004 (I19348,I19591,I19413);
nand I_1005 (I19336,I19591,I19526);
nand I_1006 (I19636,I38302,I38308);
and I_1007 (I19653,I19636,I38311);
DFFARX1 I_1008 (I19653,I2507,I19362,I19679,);
nor I_1009 (I19687,I19679,I19388);
DFFARX1 I_1010 (I19687,I2507,I19362,I19330,);
not I_1011 (I19718,I19679);
nor I_1012 (I19735,I38314,I38308);
not I_1013 (I19752,I19735);
nor I_1014 (I19769,I19526,I19752);
nor I_1015 (I19786,I19718,I19769);
DFFARX1 I_1016 (I19786,I2507,I19362,I19351,);
nor I_1017 (I19817,I19679,I19752);
nor I_1018 (I19339,I19543,I19817);
nor I_1019 (I19333,I19679,I19735);
not I_1020 (I19889,I2514);
DFFARX1 I_1021 (I588463,I2507,I19889,I19915,);
DFFARX1 I_1022 (I19915,I2507,I19889,I19932,);
not I_1023 (I19940,I19932);
nand I_1024 (I19957,I588451,I588442);
and I_1025 (I19974,I19957,I588439);
DFFARX1 I_1026 (I19974,I2507,I19889,I20000,);
DFFARX1 I_1027 (I20000,I2507,I19889,I19881,);
DFFARX1 I_1028 (I20000,I2507,I19889,I19872,);
DFFARX1 I_1029 (I588445,I2507,I19889,I20045,);
nand I_1030 (I20053,I20045,I588457);
not I_1031 (I20070,I20053);
nor I_1032 (I19869,I19915,I20070);
DFFARX1 I_1033 (I588454,I2507,I19889,I20110,);
not I_1034 (I20118,I20110);
nor I_1035 (I19875,I20118,I19940);
nand I_1036 (I19863,I20118,I20053);
nand I_1037 (I20163,I588448,I588442);
and I_1038 (I20180,I20163,I588460);
DFFARX1 I_1039 (I20180,I2507,I19889,I20206,);
nor I_1040 (I20214,I20206,I19915);
DFFARX1 I_1041 (I20214,I2507,I19889,I19857,);
not I_1042 (I20245,I20206);
nor I_1043 (I20262,I588439,I588442);
not I_1044 (I20279,I20262);
nor I_1045 (I20296,I20053,I20279);
nor I_1046 (I20313,I20245,I20296);
DFFARX1 I_1047 (I20313,I2507,I19889,I19878,);
nor I_1048 (I20344,I20206,I20279);
nor I_1049 (I19866,I20070,I20344);
nor I_1050 (I19860,I20206,I20262);
not I_1051 (I20416,I2514);
DFFARX1 I_1052 (I48318,I2507,I20416,I20442,);
DFFARX1 I_1053 (I20442,I2507,I20416,I20459,);
not I_1054 (I20467,I20459);
nand I_1055 (I20484,I48318,I48333);
and I_1056 (I20501,I20484,I48336);
DFFARX1 I_1057 (I20501,I2507,I20416,I20527,);
DFFARX1 I_1058 (I20527,I2507,I20416,I20408,);
DFFARX1 I_1059 (I20527,I2507,I20416,I20399,);
DFFARX1 I_1060 (I48330,I2507,I20416,I20572,);
nand I_1061 (I20580,I20572,I48339);
not I_1062 (I20597,I20580);
nor I_1063 (I20396,I20442,I20597);
DFFARX1 I_1064 (I48315,I2507,I20416,I20637,);
not I_1065 (I20645,I20637);
nor I_1066 (I20402,I20645,I20467);
nand I_1067 (I20390,I20645,I20580);
nand I_1068 (I20690,I48315,I48321);
and I_1069 (I20707,I20690,I48324);
DFFARX1 I_1070 (I20707,I2507,I20416,I20733,);
nor I_1071 (I20741,I20733,I20442);
DFFARX1 I_1072 (I20741,I2507,I20416,I20384,);
not I_1073 (I20772,I20733);
nor I_1074 (I20789,I48327,I48321);
not I_1075 (I20806,I20789);
nor I_1076 (I20823,I20580,I20806);
nor I_1077 (I20840,I20772,I20823);
DFFARX1 I_1078 (I20840,I2507,I20416,I20405,);
nor I_1079 (I20871,I20733,I20806);
nor I_1080 (I20393,I20597,I20871);
nor I_1081 (I20387,I20733,I20789);
not I_1082 (I20943,I2514);
DFFARX1 I_1083 (I243832,I2507,I20943,I20969,);
DFFARX1 I_1084 (I20969,I2507,I20943,I20986,);
not I_1085 (I20994,I20986);
nand I_1086 (I21011,I243832,I243835);
and I_1087 (I21028,I21011,I243856);
DFFARX1 I_1088 (I21028,I2507,I20943,I21054,);
DFFARX1 I_1089 (I21054,I2507,I20943,I20935,);
DFFARX1 I_1090 (I21054,I2507,I20943,I20926,);
DFFARX1 I_1091 (I243844,I2507,I20943,I21099,);
nand I_1092 (I21107,I21099,I243847);
not I_1093 (I21124,I21107);
nor I_1094 (I20923,I20969,I21124);
DFFARX1 I_1095 (I243853,I2507,I20943,I21164,);
not I_1096 (I21172,I21164);
nor I_1097 (I20929,I21172,I20994);
nand I_1098 (I20917,I21172,I21107);
nand I_1099 (I21217,I243850,I243838);
and I_1100 (I21234,I21217,I243841);
DFFARX1 I_1101 (I21234,I2507,I20943,I21260,);
nor I_1102 (I21268,I21260,I20969);
DFFARX1 I_1103 (I21268,I2507,I20943,I20911,);
not I_1104 (I21299,I21260);
nor I_1105 (I21316,I243859,I243838);
not I_1106 (I21333,I21316);
nor I_1107 (I21350,I21107,I21333);
nor I_1108 (I21367,I21299,I21350);
DFFARX1 I_1109 (I21367,I2507,I20943,I20932,);
nor I_1110 (I21398,I21260,I21333);
nor I_1111 (I20920,I21124,I21398);
nor I_1112 (I20914,I21260,I21316);
not I_1113 (I21470,I2514);
DFFARX1 I_1114 (I403893,I2507,I21470,I21496,);
DFFARX1 I_1115 (I21496,I2507,I21470,I21513,);
not I_1116 (I21521,I21513);
nand I_1117 (I21538,I403908,I403911);
and I_1118 (I21555,I21538,I403890);
DFFARX1 I_1119 (I21555,I2507,I21470,I21581,);
DFFARX1 I_1120 (I21581,I2507,I21470,I21462,);
DFFARX1 I_1121 (I21581,I2507,I21470,I21453,);
DFFARX1 I_1122 (I403896,I2507,I21470,I21626,);
nand I_1123 (I21634,I21626,I403902);
not I_1124 (I21651,I21634);
nor I_1125 (I21450,I21496,I21651);
DFFARX1 I_1126 (I403890,I2507,I21470,I21691,);
not I_1127 (I21699,I21691);
nor I_1128 (I21456,I21699,I21521);
nand I_1129 (I21444,I21699,I21634);
nand I_1130 (I21744,I403905,I403887);
and I_1131 (I21761,I21744,I403899);
DFFARX1 I_1132 (I21761,I2507,I21470,I21787,);
nor I_1133 (I21795,I21787,I21496);
DFFARX1 I_1134 (I21795,I2507,I21470,I21438,);
not I_1135 (I21826,I21787);
nor I_1136 (I21843,I403887,I403887);
not I_1137 (I21860,I21843);
nor I_1138 (I21877,I21634,I21860);
nor I_1139 (I21894,I21826,I21877);
DFFARX1 I_1140 (I21894,I2507,I21470,I21459,);
nor I_1141 (I21925,I21787,I21860);
nor I_1142 (I21447,I21651,I21925);
nor I_1143 (I21441,I21787,I21843);
not I_1144 (I21997,I2514);
DFFARX1 I_1145 (I540233,I2507,I21997,I22023,);
DFFARX1 I_1146 (I22023,I2507,I21997,I22040,);
not I_1147 (I22048,I22040);
nand I_1148 (I22065,I540227,I540248);
and I_1149 (I22082,I22065,I540233);
DFFARX1 I_1150 (I22082,I2507,I21997,I22108,);
DFFARX1 I_1151 (I22108,I2507,I21997,I21989,);
DFFARX1 I_1152 (I22108,I2507,I21997,I21980,);
DFFARX1 I_1153 (I540230,I2507,I21997,I22153,);
nand I_1154 (I22161,I22153,I540239);
not I_1155 (I22178,I22161);
nor I_1156 (I21977,I22023,I22178);
DFFARX1 I_1157 (I540227,I2507,I21997,I22218,);
not I_1158 (I22226,I22218);
nor I_1159 (I21983,I22226,I22048);
nand I_1160 (I21971,I22226,I22161);
nand I_1161 (I22271,I540230,I540245);
and I_1162 (I22288,I22271,I540236);
DFFARX1 I_1163 (I22288,I2507,I21997,I22314,);
nor I_1164 (I22322,I22314,I22023);
DFFARX1 I_1165 (I22322,I2507,I21997,I21965,);
not I_1166 (I22353,I22314);
nor I_1167 (I22370,I540242,I540245);
not I_1168 (I22387,I22370);
nor I_1169 (I22404,I22161,I22387);
nor I_1170 (I22421,I22353,I22404);
DFFARX1 I_1171 (I22421,I2507,I21997,I21986,);
nor I_1172 (I22452,I22314,I22387);
nor I_1173 (I21974,I22178,I22452);
nor I_1174 (I21968,I22314,I22370);
not I_1175 (I22524,I2514);
DFFARX1 I_1176 (I605803,I2507,I22524,I22550,);
DFFARX1 I_1177 (I22550,I2507,I22524,I22567,);
not I_1178 (I22575,I22567);
nand I_1179 (I22592,I605791,I605782);
and I_1180 (I22609,I22592,I605779);
DFFARX1 I_1181 (I22609,I2507,I22524,I22635,);
DFFARX1 I_1182 (I22635,I2507,I22524,I22516,);
DFFARX1 I_1183 (I22635,I2507,I22524,I22507,);
DFFARX1 I_1184 (I605785,I2507,I22524,I22680,);
nand I_1185 (I22688,I22680,I605797);
not I_1186 (I22705,I22688);
nor I_1187 (I22504,I22550,I22705);
DFFARX1 I_1188 (I605794,I2507,I22524,I22745,);
not I_1189 (I22753,I22745);
nor I_1190 (I22510,I22753,I22575);
nand I_1191 (I22498,I22753,I22688);
nand I_1192 (I22798,I605788,I605782);
and I_1193 (I22815,I22798,I605800);
DFFARX1 I_1194 (I22815,I2507,I22524,I22841,);
nor I_1195 (I22849,I22841,I22550);
DFFARX1 I_1196 (I22849,I2507,I22524,I22492,);
not I_1197 (I22880,I22841);
nor I_1198 (I22897,I605779,I605782);
not I_1199 (I22914,I22897);
nor I_1200 (I22931,I22688,I22914);
nor I_1201 (I22948,I22880,I22931);
DFFARX1 I_1202 (I22948,I2507,I22524,I22513,);
nor I_1203 (I22979,I22841,I22914);
nor I_1204 (I22501,I22705,I22979);
nor I_1205 (I22495,I22841,I22897);
not I_1206 (I23051,I2514);
DFFARX1 I_1207 (I182744,I2507,I23051,I23077,);
DFFARX1 I_1208 (I23077,I2507,I23051,I23094,);
not I_1209 (I23102,I23094);
nand I_1210 (I23119,I182741,I182735);
and I_1211 (I23136,I23119,I182729);
DFFARX1 I_1212 (I23136,I2507,I23051,I23162,);
DFFARX1 I_1213 (I23162,I2507,I23051,I23043,);
DFFARX1 I_1214 (I23162,I2507,I23051,I23034,);
DFFARX1 I_1215 (I182717,I2507,I23051,I23207,);
nand I_1216 (I23215,I23207,I182726);
not I_1217 (I23232,I23215);
nor I_1218 (I23031,I23077,I23232);
DFFARX1 I_1219 (I182723,I2507,I23051,I23272,);
not I_1220 (I23280,I23272);
nor I_1221 (I23037,I23280,I23102);
nand I_1222 (I23025,I23280,I23215);
nand I_1223 (I23325,I182720,I182738);
and I_1224 (I23342,I23325,I182717);
DFFARX1 I_1225 (I23342,I2507,I23051,I23368,);
nor I_1226 (I23376,I23368,I23077);
DFFARX1 I_1227 (I23376,I2507,I23051,I23019,);
not I_1228 (I23407,I23368);
nor I_1229 (I23424,I182732,I182738);
not I_1230 (I23441,I23424);
nor I_1231 (I23458,I23215,I23441);
nor I_1232 (I23475,I23407,I23458);
DFFARX1 I_1233 (I23475,I2507,I23051,I23040,);
nor I_1234 (I23506,I23368,I23441);
nor I_1235 (I23028,I23232,I23506);
nor I_1236 (I23022,I23368,I23424);
not I_1237 (I23578,I2514);
DFFARX1 I_1238 (I332230,I2507,I23578,I23604,);
DFFARX1 I_1239 (I23604,I2507,I23578,I23621,);
not I_1240 (I23629,I23621);
nand I_1241 (I23646,I332215,I332233);
and I_1242 (I23663,I23646,I332227);
DFFARX1 I_1243 (I23663,I2507,I23578,I23689,);
DFFARX1 I_1244 (I23689,I2507,I23578,I23570,);
DFFARX1 I_1245 (I23689,I2507,I23578,I23561,);
DFFARX1 I_1246 (I332224,I2507,I23578,I23734,);
nand I_1247 (I23742,I23734,I332215);
not I_1248 (I23759,I23742);
nor I_1249 (I23558,I23604,I23759);
DFFARX1 I_1250 (I332218,I2507,I23578,I23799,);
not I_1251 (I23807,I23799);
nor I_1252 (I23564,I23807,I23629);
nand I_1253 (I23552,I23807,I23742);
nand I_1254 (I23852,I332239,I332221);
and I_1255 (I23869,I23852,I332236);
DFFARX1 I_1256 (I23869,I2507,I23578,I23895,);
nor I_1257 (I23903,I23895,I23604);
DFFARX1 I_1258 (I23903,I2507,I23578,I23546,);
not I_1259 (I23934,I23895);
nor I_1260 (I23951,I332218,I332221);
not I_1261 (I23968,I23951);
nor I_1262 (I23985,I23742,I23968);
nor I_1263 (I24002,I23934,I23985);
DFFARX1 I_1264 (I24002,I2507,I23578,I23567,);
nor I_1265 (I24033,I23895,I23968);
nor I_1266 (I23555,I23759,I24033);
nor I_1267 (I23549,I23895,I23951);
not I_1268 (I24105,I2514);
DFFARX1 I_1269 (I58858,I2507,I24105,I24131,);
DFFARX1 I_1270 (I24131,I2507,I24105,I24148,);
not I_1271 (I24156,I24148);
nand I_1272 (I24173,I58858,I58873);
and I_1273 (I24190,I24173,I58876);
DFFARX1 I_1274 (I24190,I2507,I24105,I24216,);
DFFARX1 I_1275 (I24216,I2507,I24105,I24097,);
DFFARX1 I_1276 (I24216,I2507,I24105,I24088,);
DFFARX1 I_1277 (I58870,I2507,I24105,I24261,);
nand I_1278 (I24269,I24261,I58879);
not I_1279 (I24286,I24269);
nor I_1280 (I24085,I24131,I24286);
DFFARX1 I_1281 (I58855,I2507,I24105,I24326,);
not I_1282 (I24334,I24326);
nor I_1283 (I24091,I24334,I24156);
nand I_1284 (I24079,I24334,I24269);
nand I_1285 (I24379,I58855,I58861);
and I_1286 (I24396,I24379,I58864);
DFFARX1 I_1287 (I24396,I2507,I24105,I24422,);
nor I_1288 (I24430,I24422,I24131);
DFFARX1 I_1289 (I24430,I2507,I24105,I24073,);
not I_1290 (I24461,I24422);
nor I_1291 (I24478,I58867,I58861);
not I_1292 (I24495,I24478);
nor I_1293 (I24512,I24269,I24495);
nor I_1294 (I24529,I24461,I24512);
DFFARX1 I_1295 (I24529,I2507,I24105,I24094,);
nor I_1296 (I24560,I24422,I24495);
nor I_1297 (I24082,I24286,I24560);
nor I_1298 (I24076,I24422,I24478);
not I_1299 (I24632,I2514);
DFFARX1 I_1300 (I612739,I2507,I24632,I24658,);
DFFARX1 I_1301 (I24658,I2507,I24632,I24675,);
not I_1302 (I24683,I24675);
nand I_1303 (I24700,I612727,I612718);
and I_1304 (I24717,I24700,I612715);
DFFARX1 I_1305 (I24717,I2507,I24632,I24743,);
DFFARX1 I_1306 (I24743,I2507,I24632,I24624,);
DFFARX1 I_1307 (I24743,I2507,I24632,I24615,);
DFFARX1 I_1308 (I612721,I2507,I24632,I24788,);
nand I_1309 (I24796,I24788,I612733);
not I_1310 (I24813,I24796);
nor I_1311 (I24612,I24658,I24813);
DFFARX1 I_1312 (I612730,I2507,I24632,I24853,);
not I_1313 (I24861,I24853);
nor I_1314 (I24618,I24861,I24683);
nand I_1315 (I24606,I24861,I24796);
nand I_1316 (I24906,I612724,I612718);
and I_1317 (I24923,I24906,I612736);
DFFARX1 I_1318 (I24923,I2507,I24632,I24949,);
nor I_1319 (I24957,I24949,I24658);
DFFARX1 I_1320 (I24957,I2507,I24632,I24600,);
not I_1321 (I24988,I24949);
nor I_1322 (I25005,I612715,I612718);
not I_1323 (I25022,I25005);
nor I_1324 (I25039,I24796,I25022);
nor I_1325 (I25056,I24988,I25039);
DFFARX1 I_1326 (I25056,I2507,I24632,I24621,);
nor I_1327 (I25087,I24949,I25022);
nor I_1328 (I24609,I24813,I25087);
nor I_1329 (I24603,I24949,I25005);
not I_1330 (I25159,I2514);
DFFARX1 I_1331 (I531292,I2507,I25159,I25185,);
DFFARX1 I_1332 (I25185,I2507,I25159,I25202,);
not I_1333 (I25210,I25202);
nand I_1334 (I25227,I531268,I531295);
and I_1335 (I25244,I25227,I531280);
DFFARX1 I_1336 (I25244,I2507,I25159,I25270,);
DFFARX1 I_1337 (I25270,I2507,I25159,I25151,);
DFFARX1 I_1338 (I25270,I2507,I25159,I25142,);
DFFARX1 I_1339 (I531286,I2507,I25159,I25315,);
nand I_1340 (I25323,I25315,I531271);
not I_1341 (I25340,I25323);
nor I_1342 (I25139,I25185,I25340);
DFFARX1 I_1343 (I531289,I2507,I25159,I25380,);
not I_1344 (I25388,I25380);
nor I_1345 (I25145,I25388,I25210);
nand I_1346 (I25133,I25388,I25323);
nand I_1347 (I25433,I531274,I531277);
and I_1348 (I25450,I25433,I531268);
DFFARX1 I_1349 (I25450,I2507,I25159,I25476,);
nor I_1350 (I25484,I25476,I25185);
DFFARX1 I_1351 (I25484,I2507,I25159,I25127,);
not I_1352 (I25515,I25476);
nor I_1353 (I25532,I531283,I531277);
not I_1354 (I25549,I25532);
nor I_1355 (I25566,I25323,I25549);
nor I_1356 (I25583,I25515,I25566);
DFFARX1 I_1357 (I25583,I2507,I25159,I25148,);
nor I_1358 (I25614,I25476,I25549);
nor I_1359 (I25136,I25340,I25614);
nor I_1360 (I25130,I25476,I25532);
not I_1361 (I25686,I2514);
DFFARX1 I_1362 (I568844,I2507,I25686,I25712,);
DFFARX1 I_1363 (I25712,I2507,I25686,I25729,);
not I_1364 (I25737,I25729);
nand I_1365 (I25754,I568838,I568859);
and I_1366 (I25771,I25754,I568844);
DFFARX1 I_1367 (I25771,I2507,I25686,I25797,);
DFFARX1 I_1368 (I25797,I2507,I25686,I25678,);
DFFARX1 I_1369 (I25797,I2507,I25686,I25669,);
DFFARX1 I_1370 (I568841,I2507,I25686,I25842,);
nand I_1371 (I25850,I25842,I568850);
not I_1372 (I25867,I25850);
nor I_1373 (I25666,I25712,I25867);
DFFARX1 I_1374 (I568838,I2507,I25686,I25907,);
not I_1375 (I25915,I25907);
nor I_1376 (I25672,I25915,I25737);
nand I_1377 (I25660,I25915,I25850);
nand I_1378 (I25960,I568841,I568856);
and I_1379 (I25977,I25960,I568847);
DFFARX1 I_1380 (I25977,I2507,I25686,I26003,);
nor I_1381 (I26011,I26003,I25712);
DFFARX1 I_1382 (I26011,I2507,I25686,I25654,);
not I_1383 (I26042,I26003);
nor I_1384 (I26059,I568853,I568856);
not I_1385 (I26076,I26059);
nor I_1386 (I26093,I25850,I26076);
nor I_1387 (I26110,I26042,I26093);
DFFARX1 I_1388 (I26110,I2507,I25686,I25675,);
nor I_1389 (I26141,I26003,I26076);
nor I_1390 (I25663,I25867,I26141);
nor I_1391 (I25657,I26003,I26059);
not I_1392 (I26213,I2514);
DFFARX1 I_1393 (I1876,I2507,I26213,I26239,);
DFFARX1 I_1394 (I26239,I2507,I26213,I26256,);
not I_1395 (I26264,I26256);
nand I_1396 (I26281,I1460,I2468);
and I_1397 (I26298,I26281,I2244);
DFFARX1 I_1398 (I26298,I2507,I26213,I26324,);
DFFARX1 I_1399 (I26324,I2507,I26213,I26205,);
DFFARX1 I_1400 (I26324,I2507,I26213,I26196,);
DFFARX1 I_1401 (I2036,I2507,I26213,I26369,);
nand I_1402 (I26377,I26369,I1620);
not I_1403 (I26394,I26377);
nor I_1404 (I26193,I26239,I26394);
DFFARX1 I_1405 (I1844,I2507,I26213,I26434,);
not I_1406 (I26442,I26434);
nor I_1407 (I26199,I26442,I26264);
nand I_1408 (I26187,I26442,I26377);
nand I_1409 (I26487,I2396,I1676);
and I_1410 (I26504,I26487,I1420);
DFFARX1 I_1411 (I26504,I2507,I26213,I26530,);
nor I_1412 (I26538,I26530,I26239);
DFFARX1 I_1413 (I26538,I2507,I26213,I26181,);
not I_1414 (I26569,I26530);
nor I_1415 (I26586,I1716,I1676);
not I_1416 (I26603,I26586);
nor I_1417 (I26620,I26377,I26603);
nor I_1418 (I26637,I26569,I26620);
DFFARX1 I_1419 (I26637,I2507,I26213,I26202,);
nor I_1420 (I26668,I26530,I26603);
nor I_1421 (I26190,I26394,I26668);
nor I_1422 (I26184,I26530,I26586);
not I_1423 (I26740,I2514);
DFFARX1 I_1424 (I443404,I2507,I26740,I26766,);
DFFARX1 I_1425 (I26766,I2507,I26740,I26783,);
not I_1426 (I26791,I26783);
nand I_1427 (I26808,I443395,I443416);
and I_1428 (I26825,I26808,I443398);
DFFARX1 I_1429 (I26825,I2507,I26740,I26851,);
DFFARX1 I_1430 (I26851,I2507,I26740,I26732,);
DFFARX1 I_1431 (I26851,I2507,I26740,I26723,);
DFFARX1 I_1432 (I443398,I2507,I26740,I26896,);
nand I_1433 (I26904,I26896,I443413);
not I_1434 (I26921,I26904);
nor I_1435 (I26720,I26766,I26921);
DFFARX1 I_1436 (I443407,I2507,I26740,I26961,);
not I_1437 (I26969,I26961);
nor I_1438 (I26726,I26969,I26791);
nand I_1439 (I26714,I26969,I26904);
nand I_1440 (I27014,I443401,I443410);
and I_1441 (I27031,I27014,I443395);
DFFARX1 I_1442 (I27031,I2507,I26740,I27057,);
nor I_1443 (I27065,I27057,I26766);
DFFARX1 I_1444 (I27065,I2507,I26740,I26708,);
not I_1445 (I27096,I27057);
nor I_1446 (I27113,I443401,I443410);
not I_1447 (I27130,I27113);
nor I_1448 (I27147,I26904,I27130);
nor I_1449 (I27164,I27096,I27147);
DFFARX1 I_1450 (I27164,I2507,I26740,I26729,);
nor I_1451 (I27195,I27057,I27130);
nor I_1452 (I26717,I26921,I27195);
nor I_1453 (I26711,I27057,I27113);
not I_1454 (I27267,I2514);
DFFARX1 I_1455 (I209621,I2507,I27267,I27293,);
DFFARX1 I_1456 (I27293,I2507,I27267,I27310,);
not I_1457 (I27318,I27310);
nand I_1458 (I27335,I209618,I209612);
and I_1459 (I27352,I27335,I209606);
DFFARX1 I_1460 (I27352,I2507,I27267,I27378,);
DFFARX1 I_1461 (I27378,I2507,I27267,I27259,);
DFFARX1 I_1462 (I27378,I2507,I27267,I27250,);
DFFARX1 I_1463 (I209594,I2507,I27267,I27423,);
nand I_1464 (I27431,I27423,I209603);
not I_1465 (I27448,I27431);
nor I_1466 (I27247,I27293,I27448);
DFFARX1 I_1467 (I209600,I2507,I27267,I27488,);
not I_1468 (I27496,I27488);
nor I_1469 (I27253,I27496,I27318);
nand I_1470 (I27241,I27496,I27431);
nand I_1471 (I27541,I209597,I209615);
and I_1472 (I27558,I27541,I209594);
DFFARX1 I_1473 (I27558,I2507,I27267,I27584,);
nor I_1474 (I27592,I27584,I27293);
DFFARX1 I_1475 (I27592,I2507,I27267,I27235,);
not I_1476 (I27623,I27584);
nor I_1477 (I27640,I209609,I209615);
not I_1478 (I27657,I27640);
nor I_1479 (I27674,I27431,I27657);
nor I_1480 (I27691,I27623,I27674);
DFFARX1 I_1481 (I27691,I2507,I27267,I27256,);
nor I_1482 (I27722,I27584,I27657);
nor I_1483 (I27244,I27448,I27722);
nor I_1484 (I27238,I27584,I27640);
not I_1485 (I27794,I2514);
DFFARX1 I_1486 (I652325,I2507,I27794,I27820,);
DFFARX1 I_1487 (I27820,I2507,I27794,I27837,);
not I_1488 (I27845,I27837);
nand I_1489 (I27862,I652343,I652337);
and I_1490 (I27879,I27862,I652346);
DFFARX1 I_1491 (I27879,I2507,I27794,I27905,);
DFFARX1 I_1492 (I27905,I2507,I27794,I27786,);
DFFARX1 I_1493 (I27905,I2507,I27794,I27777,);
DFFARX1 I_1494 (I652331,I2507,I27794,I27950,);
nand I_1495 (I27958,I27950,I652340);
not I_1496 (I27975,I27958);
nor I_1497 (I27774,I27820,I27975);
DFFARX1 I_1498 (I652328,I2507,I27794,I28015,);
not I_1499 (I28023,I28015);
nor I_1500 (I27780,I28023,I27845);
nand I_1501 (I27768,I28023,I27958);
nand I_1502 (I28068,I652349,I652334);
and I_1503 (I28085,I28068,I652328);
DFFARX1 I_1504 (I28085,I2507,I27794,I28111,);
nor I_1505 (I28119,I28111,I27820);
DFFARX1 I_1506 (I28119,I2507,I27794,I27762,);
not I_1507 (I28150,I28111);
nor I_1508 (I28167,I652325,I652334);
not I_1509 (I28184,I28167);
nor I_1510 (I28201,I27958,I28184);
nor I_1511 (I28218,I28150,I28201);
DFFARX1 I_1512 (I28218,I2507,I27794,I27783,);
nor I_1513 (I28249,I28111,I28184);
nor I_1514 (I27771,I27975,I28249);
nor I_1515 (I27765,I28111,I28167);
not I_1516 (I28321,I2514);
DFFARX1 I_1517 (I94340,I2507,I28321,I28347,);
DFFARX1 I_1518 (I28347,I2507,I28321,I28364,);
not I_1519 (I28372,I28364);
nand I_1520 (I28389,I94358,I94343);
and I_1521 (I28406,I28389,I94346);
DFFARX1 I_1522 (I28406,I2507,I28321,I28432,);
DFFARX1 I_1523 (I28432,I2507,I28321,I28313,);
DFFARX1 I_1524 (I28432,I2507,I28321,I28304,);
DFFARX1 I_1525 (I94334,I2507,I28321,I28477,);
nand I_1526 (I28485,I28477,I94337);
not I_1527 (I28502,I28485);
nor I_1528 (I28301,I28347,I28502);
DFFARX1 I_1529 (I94349,I2507,I28321,I28542,);
not I_1530 (I28550,I28542);
nor I_1531 (I28307,I28550,I28372);
nand I_1532 (I28295,I28550,I28485);
nand I_1533 (I28595,I94355,I94352);
and I_1534 (I28612,I28595,I94337);
DFFARX1 I_1535 (I28612,I2507,I28321,I28638,);
nor I_1536 (I28646,I28638,I28347);
DFFARX1 I_1537 (I28646,I2507,I28321,I28289,);
not I_1538 (I28677,I28638);
nor I_1539 (I28694,I94334,I94352);
not I_1540 (I28711,I28694);
nor I_1541 (I28728,I28485,I28711);
nor I_1542 (I28745,I28677,I28728);
DFFARX1 I_1543 (I28745,I2507,I28321,I28310,);
nor I_1544 (I28776,I28638,I28711);
nor I_1545 (I28298,I28502,I28776);
nor I_1546 (I28292,I28638,I28694);
not I_1547 (I28848,I2514);
DFFARX1 I_1548 (I299227,I2507,I28848,I28874,);
DFFARX1 I_1549 (I28874,I2507,I28848,I28891,);
not I_1550 (I28899,I28891);
nand I_1551 (I28916,I299233,I299221);
and I_1552 (I28933,I28916,I299218);
DFFARX1 I_1553 (I28933,I2507,I28848,I28959,);
DFFARX1 I_1554 (I28959,I2507,I28848,I28840,);
DFFARX1 I_1555 (I28959,I2507,I28848,I28831,);
DFFARX1 I_1556 (I299230,I2507,I28848,I29004,);
nand I_1557 (I29012,I29004,I299224);
not I_1558 (I29029,I29012);
nor I_1559 (I28828,I28874,I29029);
DFFARX1 I_1560 (I299242,I2507,I28848,I29069,);
not I_1561 (I29077,I29069);
nor I_1562 (I28834,I29077,I28899);
nand I_1563 (I28822,I29077,I29012);
nand I_1564 (I29122,I299236,I299239);
and I_1565 (I29139,I29122,I299221);
DFFARX1 I_1566 (I29139,I2507,I28848,I29165,);
nor I_1567 (I29173,I29165,I28874);
DFFARX1 I_1568 (I29173,I2507,I28848,I28816,);
not I_1569 (I29204,I29165);
nor I_1570 (I29221,I299218,I299239);
not I_1571 (I29238,I29221);
nor I_1572 (I29255,I29012,I29238);
nor I_1573 (I29272,I29204,I29255);
DFFARX1 I_1574 (I29272,I2507,I28848,I28837,);
nor I_1575 (I29303,I29165,I29238);
nor I_1576 (I28825,I29029,I29303);
nor I_1577 (I28819,I29165,I29221);
not I_1578 (I29375,I2514);
DFFARX1 I_1579 (I155030,I2507,I29375,I29401,);
DFFARX1 I_1580 (I29401,I2507,I29375,I29418,);
not I_1581 (I29426,I29418);
nand I_1582 (I29443,I155048,I155033);
and I_1583 (I29460,I29443,I155036);
DFFARX1 I_1584 (I29460,I2507,I29375,I29486,);
DFFARX1 I_1585 (I29486,I2507,I29375,I29367,);
DFFARX1 I_1586 (I29486,I2507,I29375,I29358,);
DFFARX1 I_1587 (I155024,I2507,I29375,I29531,);
nand I_1588 (I29539,I29531,I155027);
not I_1589 (I29556,I29539);
nor I_1590 (I29355,I29401,I29556);
DFFARX1 I_1591 (I155039,I2507,I29375,I29596,);
not I_1592 (I29604,I29596);
nor I_1593 (I29361,I29604,I29426);
nand I_1594 (I29349,I29604,I29539);
nand I_1595 (I29649,I155045,I155042);
and I_1596 (I29666,I29649,I155027);
DFFARX1 I_1597 (I29666,I2507,I29375,I29692,);
nor I_1598 (I29700,I29692,I29401);
DFFARX1 I_1599 (I29700,I2507,I29375,I29343,);
not I_1600 (I29731,I29692);
nor I_1601 (I29748,I155024,I155042);
not I_1602 (I29765,I29748);
nor I_1603 (I29782,I29539,I29765);
nor I_1604 (I29799,I29731,I29782);
DFFARX1 I_1605 (I29799,I2507,I29375,I29364,);
nor I_1606 (I29830,I29692,I29765);
nor I_1607 (I29352,I29556,I29830);
nor I_1608 (I29346,I29692,I29748);
not I_1609 (I29902,I2514);
DFFARX1 I_1610 (I317202,I2507,I29902,I29928,);
DFFARX1 I_1611 (I29928,I2507,I29902,I29945,);
not I_1612 (I29953,I29945);
nand I_1613 (I29970,I317187,I317205);
and I_1614 (I29987,I29970,I317199);
DFFARX1 I_1615 (I29987,I2507,I29902,I30013,);
DFFARX1 I_1616 (I30013,I2507,I29902,I29894,);
DFFARX1 I_1617 (I30013,I2507,I29902,I29885,);
DFFARX1 I_1618 (I317196,I2507,I29902,I30058,);
nand I_1619 (I30066,I30058,I317187);
not I_1620 (I30083,I30066);
nor I_1621 (I29882,I29928,I30083);
DFFARX1 I_1622 (I317190,I2507,I29902,I30123,);
not I_1623 (I30131,I30123);
nor I_1624 (I29888,I30131,I29953);
nand I_1625 (I29876,I30131,I30066);
nand I_1626 (I30176,I317211,I317193);
and I_1627 (I30193,I30176,I317208);
DFFARX1 I_1628 (I30193,I2507,I29902,I30219,);
nor I_1629 (I30227,I30219,I29928);
DFFARX1 I_1630 (I30227,I2507,I29902,I29870,);
not I_1631 (I30258,I30219);
nor I_1632 (I30275,I317190,I317193);
not I_1633 (I30292,I30275);
nor I_1634 (I30309,I30066,I30292);
nor I_1635 (I30326,I30258,I30309);
DFFARX1 I_1636 (I30326,I2507,I29902,I29891,);
nor I_1637 (I30357,I30219,I30292);
nor I_1638 (I29879,I30083,I30357);
nor I_1639 (I29873,I30219,I30275);
not I_1640 (I30429,I2514);
DFFARX1 I_1641 (I528708,I2507,I30429,I30455,);
DFFARX1 I_1642 (I30455,I2507,I30429,I30472,);
not I_1643 (I30480,I30472);
nand I_1644 (I30497,I528684,I528711);
and I_1645 (I30514,I30497,I528696);
DFFARX1 I_1646 (I30514,I2507,I30429,I30540,);
DFFARX1 I_1647 (I30540,I2507,I30429,I30421,);
DFFARX1 I_1648 (I30540,I2507,I30429,I30412,);
DFFARX1 I_1649 (I528702,I2507,I30429,I30585,);
nand I_1650 (I30593,I30585,I528687);
not I_1651 (I30610,I30593);
nor I_1652 (I30409,I30455,I30610);
DFFARX1 I_1653 (I528705,I2507,I30429,I30650,);
not I_1654 (I30658,I30650);
nor I_1655 (I30415,I30658,I30480);
nand I_1656 (I30403,I30658,I30593);
nand I_1657 (I30703,I528690,I528693);
and I_1658 (I30720,I30703,I528684);
DFFARX1 I_1659 (I30720,I2507,I30429,I30746,);
nor I_1660 (I30754,I30746,I30455);
DFFARX1 I_1661 (I30754,I2507,I30429,I30397,);
not I_1662 (I30785,I30746);
nor I_1663 (I30802,I528699,I528693);
not I_1664 (I30819,I30802);
nor I_1665 (I30836,I30593,I30819);
nor I_1666 (I30853,I30785,I30836);
DFFARX1 I_1667 (I30853,I2507,I30429,I30418,);
nor I_1668 (I30884,I30746,I30819);
nor I_1669 (I30406,I30610,I30884);
nor I_1670 (I30400,I30746,I30802);
not I_1671 (I30956,I2514);
DFFARX1 I_1672 (I497700,I2507,I30956,I30982,);
DFFARX1 I_1673 (I30982,I2507,I30956,I30999,);
not I_1674 (I31007,I30999);
nand I_1675 (I31024,I497676,I497703);
and I_1676 (I31041,I31024,I497688);
DFFARX1 I_1677 (I31041,I2507,I30956,I31067,);
DFFARX1 I_1678 (I31067,I2507,I30956,I30948,);
DFFARX1 I_1679 (I31067,I2507,I30956,I30939,);
DFFARX1 I_1680 (I497694,I2507,I30956,I31112,);
nand I_1681 (I31120,I31112,I497679);
not I_1682 (I31137,I31120);
nor I_1683 (I30936,I30982,I31137);
DFFARX1 I_1684 (I497697,I2507,I30956,I31177,);
not I_1685 (I31185,I31177);
nor I_1686 (I30942,I31185,I31007);
nand I_1687 (I30930,I31185,I31120);
nand I_1688 (I31230,I497682,I497685);
and I_1689 (I31247,I31230,I497676);
DFFARX1 I_1690 (I31247,I2507,I30956,I31273,);
nor I_1691 (I31281,I31273,I30982);
DFFARX1 I_1692 (I31281,I2507,I30956,I30924,);
not I_1693 (I31312,I31273);
nor I_1694 (I31329,I497691,I497685);
not I_1695 (I31346,I31329);
nor I_1696 (I31363,I31120,I31346);
nor I_1697 (I31380,I31312,I31363);
DFFARX1 I_1698 (I31380,I2507,I30956,I30945,);
nor I_1699 (I31411,I31273,I31346);
nor I_1700 (I30933,I31137,I31411);
nor I_1701 (I30927,I31273,I31329);
not I_1702 (I31483,I2514);
DFFARX1 I_1703 (I621409,I2507,I31483,I31509,);
DFFARX1 I_1704 (I31509,I2507,I31483,I31526,);
not I_1705 (I31534,I31526);
nand I_1706 (I31551,I621397,I621388);
and I_1707 (I31568,I31551,I621385);
DFFARX1 I_1708 (I31568,I2507,I31483,I31594,);
DFFARX1 I_1709 (I31594,I2507,I31483,I31475,);
DFFARX1 I_1710 (I31594,I2507,I31483,I31466,);
DFFARX1 I_1711 (I621391,I2507,I31483,I31639,);
nand I_1712 (I31647,I31639,I621403);
not I_1713 (I31664,I31647);
nor I_1714 (I31463,I31509,I31664);
DFFARX1 I_1715 (I621400,I2507,I31483,I31704,);
not I_1716 (I31712,I31704);
nor I_1717 (I31469,I31712,I31534);
nand I_1718 (I31457,I31712,I31647);
nand I_1719 (I31757,I621394,I621388);
and I_1720 (I31774,I31757,I621406);
DFFARX1 I_1721 (I31774,I2507,I31483,I31800,);
nor I_1722 (I31808,I31800,I31509);
DFFARX1 I_1723 (I31808,I2507,I31483,I31451,);
not I_1724 (I31839,I31800);
nor I_1725 (I31856,I621385,I621388);
not I_1726 (I31873,I31856);
nor I_1727 (I31890,I31647,I31873);
nor I_1728 (I31907,I31839,I31890);
DFFARX1 I_1729 (I31907,I2507,I31483,I31472,);
nor I_1730 (I31938,I31800,I31873);
nor I_1731 (I31460,I31664,I31938);
nor I_1732 (I31454,I31800,I31856);
not I_1733 (I32010,I2514);
DFFARX1 I_1734 (I684428,I2507,I32010,I32036,);
DFFARX1 I_1735 (I32036,I2507,I32010,I32053,);
not I_1736 (I32061,I32053);
nand I_1737 (I32078,I684419,I684425);
and I_1738 (I32095,I32078,I684404);
DFFARX1 I_1739 (I32095,I2507,I32010,I32121,);
DFFARX1 I_1740 (I32121,I2507,I32010,I32002,);
DFFARX1 I_1741 (I32121,I2507,I32010,I31993,);
DFFARX1 I_1742 (I684422,I2507,I32010,I32166,);
nand I_1743 (I32174,I32166,I684404);
not I_1744 (I32191,I32174);
nor I_1745 (I31990,I32036,I32191);
DFFARX1 I_1746 (I684416,I2507,I32010,I32231,);
not I_1747 (I32239,I32231);
nor I_1748 (I31996,I32239,I32061);
nand I_1749 (I31984,I32239,I32174);
nand I_1750 (I32284,I684410,I684431);
and I_1751 (I32301,I32284,I684413);
DFFARX1 I_1752 (I32301,I2507,I32010,I32327,);
nor I_1753 (I32335,I32327,I32036);
DFFARX1 I_1754 (I32335,I2507,I32010,I31978,);
not I_1755 (I32366,I32327);
nor I_1756 (I32383,I684407,I684431);
not I_1757 (I32400,I32383);
nor I_1758 (I32417,I32174,I32400);
nor I_1759 (I32434,I32366,I32417);
DFFARX1 I_1760 (I32434,I2507,I32010,I31999,);
nor I_1761 (I32465,I32327,I32400);
nor I_1762 (I31987,I32191,I32465);
nor I_1763 (I31981,I32327,I32383);
not I_1764 (I32537,I2514);
DFFARX1 I_1765 (I700758,I2507,I32537,I32563,);
DFFARX1 I_1766 (I32563,I2507,I32537,I32580,);
not I_1767 (I32588,I32580);
nand I_1768 (I32605,I700761,I700767);
and I_1769 (I32622,I32605,I700776);
DFFARX1 I_1770 (I32622,I2507,I32537,I32648,);
DFFARX1 I_1771 (I32648,I2507,I32537,I32529,);
DFFARX1 I_1772 (I32648,I2507,I32537,I32520,);
DFFARX1 I_1773 (I700779,I2507,I32537,I32693,);
nand I_1774 (I32701,I32693,I700770);
not I_1775 (I32718,I32701);
nor I_1776 (I32517,I32563,I32718);
DFFARX1 I_1777 (I700758,I2507,I32537,I32758,);
not I_1778 (I32766,I32758);
nor I_1779 (I32523,I32766,I32588);
nand I_1780 (I32511,I32766,I32701);
nand I_1781 (I32811,I700785,I700764);
and I_1782 (I32828,I32811,I700773);
DFFARX1 I_1783 (I32828,I2507,I32537,I32854,);
nor I_1784 (I32862,I32854,I32563);
DFFARX1 I_1785 (I32862,I2507,I32537,I32505,);
not I_1786 (I32893,I32854);
nor I_1787 (I32910,I700782,I700764);
not I_1788 (I32927,I32910);
nor I_1789 (I32944,I32701,I32927);
nor I_1790 (I32961,I32893,I32944);
DFFARX1 I_1791 (I32961,I2507,I32537,I32526,);
nor I_1792 (I32992,I32854,I32927);
nor I_1793 (I32514,I32718,I32992);
nor I_1794 (I32508,I32854,I32910);
not I_1795 (I33064,I2514);
DFFARX1 I_1796 (I512558,I2507,I33064,I33090,);
DFFARX1 I_1797 (I33090,I2507,I33064,I33107,);
not I_1798 (I33115,I33107);
nand I_1799 (I33132,I512534,I512561);
and I_1800 (I33149,I33132,I512546);
DFFARX1 I_1801 (I33149,I2507,I33064,I33175,);
DFFARX1 I_1802 (I33175,I2507,I33064,I33056,);
DFFARX1 I_1803 (I33175,I2507,I33064,I33047,);
DFFARX1 I_1804 (I512552,I2507,I33064,I33220,);
nand I_1805 (I33228,I33220,I512537);
not I_1806 (I33245,I33228);
nor I_1807 (I33044,I33090,I33245);
DFFARX1 I_1808 (I512555,I2507,I33064,I33285,);
not I_1809 (I33293,I33285);
nor I_1810 (I33050,I33293,I33115);
nand I_1811 (I33038,I33293,I33228);
nand I_1812 (I33338,I512540,I512543);
and I_1813 (I33355,I33338,I512534);
DFFARX1 I_1814 (I33355,I2507,I33064,I33381,);
nor I_1815 (I33389,I33381,I33090);
DFFARX1 I_1816 (I33389,I2507,I33064,I33032,);
not I_1817 (I33420,I33381);
nor I_1818 (I33437,I512549,I512543);
not I_1819 (I33454,I33437);
nor I_1820 (I33471,I33228,I33454);
nor I_1821 (I33488,I33420,I33471);
DFFARX1 I_1822 (I33488,I2507,I33064,I33053,);
nor I_1823 (I33519,I33381,I33454);
nor I_1824 (I33041,I33245,I33519);
nor I_1825 (I33035,I33381,I33437);
not I_1826 (I33591,I2514);
DFFARX1 I_1827 (I686087,I2507,I33591,I33617,);
not I_1828 (I33625,I33617);
nand I_1829 (I33642,I686093,I686111);
and I_1830 (I33659,I33642,I686108);
DFFARX1 I_1831 (I33659,I2507,I33591,I33685,);
DFFARX1 I_1832 (I686105,I2507,I33591,I33702,);
and I_1833 (I33710,I33702,I686099);
nor I_1834 (I33727,I33685,I33710);
DFFARX1 I_1835 (I33727,I2507,I33591,I33559,);
nand I_1836 (I33758,I33702,I686099);
nand I_1837 (I33775,I33625,I33758);
not I_1838 (I33571,I33775);
DFFARX1 I_1839 (I686087,I2507,I33591,I33815,);
DFFARX1 I_1840 (I33815,I2507,I33591,I33580,);
nand I_1841 (I33837,I686102,I686090);
and I_1842 (I33854,I33837,I686114);
DFFARX1 I_1843 (I33854,I2507,I33591,I33880,);
DFFARX1 I_1844 (I33880,I2507,I33591,I33897,);
not I_1845 (I33583,I33897);
not I_1846 (I33919,I33880);
nand I_1847 (I33568,I33919,I33758);
nor I_1848 (I33950,I686096,I686090);
not I_1849 (I33967,I33950);
nor I_1850 (I33984,I33919,I33967);
nor I_1851 (I34001,I33625,I33984);
DFFARX1 I_1852 (I34001,I2507,I33591,I33577,);
nor I_1853 (I34032,I33685,I33967);
nor I_1854 (I33565,I33880,I34032);
nor I_1855 (I33574,I33815,I33950);
nor I_1856 (I33562,I33685,I33950);
not I_1857 (I34118,I2514);
DFFARX1 I_1858 (I633529,I2507,I34118,I34144,);
not I_1859 (I34152,I34144);
nand I_1860 (I34169,I633544,I633523);
and I_1861 (I34186,I34169,I633526);
DFFARX1 I_1862 (I34186,I2507,I34118,I34212,);
DFFARX1 I_1863 (I633547,I2507,I34118,I34229,);
and I_1864 (I34237,I34229,I633526);
nor I_1865 (I34254,I34212,I34237);
DFFARX1 I_1866 (I34254,I2507,I34118,I34086,);
nand I_1867 (I34285,I34229,I633526);
nand I_1868 (I34302,I34152,I34285);
not I_1869 (I34098,I34302);
DFFARX1 I_1870 (I633523,I2507,I34118,I34342,);
DFFARX1 I_1871 (I34342,I2507,I34118,I34107,);
nand I_1872 (I34364,I633535,I633532);
and I_1873 (I34381,I34364,I633538);
DFFARX1 I_1874 (I34381,I2507,I34118,I34407,);
DFFARX1 I_1875 (I34407,I2507,I34118,I34424,);
not I_1876 (I34110,I34424);
not I_1877 (I34446,I34407);
nand I_1878 (I34095,I34446,I34285);
nor I_1879 (I34477,I633541,I633532);
not I_1880 (I34494,I34477);
nor I_1881 (I34511,I34446,I34494);
nor I_1882 (I34528,I34152,I34511);
DFFARX1 I_1883 (I34528,I2507,I34118,I34104,);
nor I_1884 (I34559,I34212,I34494);
nor I_1885 (I34092,I34407,I34559);
nor I_1886 (I34101,I34342,I34477);
nor I_1887 (I34089,I34212,I34477);
not I_1888 (I34645,I2514);
DFFARX1 I_1889 (I221742,I2507,I34645,I34671,);
not I_1890 (I34679,I34671);
nand I_1891 (I34696,I221724,I221739);
and I_1892 (I34713,I34696,I221715);
DFFARX1 I_1893 (I34713,I2507,I34645,I34739,);
DFFARX1 I_1894 (I221718,I2507,I34645,I34756,);
and I_1895 (I34764,I34756,I221733);
nor I_1896 (I34781,I34739,I34764);
DFFARX1 I_1897 (I34781,I2507,I34645,I34613,);
nand I_1898 (I34812,I34756,I221733);
nand I_1899 (I34829,I34679,I34812);
not I_1900 (I34625,I34829);
DFFARX1 I_1901 (I221736,I2507,I34645,I34869,);
DFFARX1 I_1902 (I34869,I2507,I34645,I34634,);
nand I_1903 (I34891,I221715,I221727);
and I_1904 (I34908,I34891,I221721);
DFFARX1 I_1905 (I34908,I2507,I34645,I34934,);
DFFARX1 I_1906 (I34934,I2507,I34645,I34951,);
not I_1907 (I34637,I34951);
not I_1908 (I34973,I34934);
nand I_1909 (I34622,I34973,I34812);
nor I_1910 (I35004,I221730,I221727);
not I_1911 (I35021,I35004);
nor I_1912 (I35038,I34973,I35021);
nor I_1913 (I35055,I34679,I35038);
DFFARX1 I_1914 (I35055,I2507,I34645,I34631,);
nor I_1915 (I35086,I34739,I35021);
nor I_1916 (I34619,I34934,I35086);
nor I_1917 (I34628,I34869,I35004);
nor I_1918 (I34616,I34739,I35004);
not I_1919 (I35172,I2514);
DFFARX1 I_1920 (I12503,I2507,I35172,I35198,);
not I_1921 (I35206,I35198);
nand I_1922 (I35223,I12491,I12497);
and I_1923 (I35240,I35223,I12500);
DFFARX1 I_1924 (I35240,I2507,I35172,I35266,);
DFFARX1 I_1925 (I12482,I2507,I35172,I35283,);
and I_1926 (I35291,I35283,I12488);
nor I_1927 (I35308,I35266,I35291);
DFFARX1 I_1928 (I35308,I2507,I35172,I35140,);
nand I_1929 (I35339,I35283,I12488);
nand I_1930 (I35356,I35206,I35339);
not I_1931 (I35152,I35356);
DFFARX1 I_1932 (I12482,I2507,I35172,I35396,);
DFFARX1 I_1933 (I35396,I2507,I35172,I35161,);
nand I_1934 (I35418,I12485,I12479);
and I_1935 (I35435,I35418,I12494);
DFFARX1 I_1936 (I35435,I2507,I35172,I35461,);
DFFARX1 I_1937 (I35461,I2507,I35172,I35478,);
not I_1938 (I35164,I35478);
not I_1939 (I35500,I35461);
nand I_1940 (I35149,I35500,I35339);
nor I_1941 (I35531,I12479,I12479);
not I_1942 (I35548,I35531);
nor I_1943 (I35565,I35500,I35548);
nor I_1944 (I35582,I35206,I35565);
DFFARX1 I_1945 (I35582,I2507,I35172,I35158,);
nor I_1946 (I35613,I35266,I35548);
nor I_1947 (I35146,I35461,I35613);
nor I_1948 (I35155,I35396,I35531);
nor I_1949 (I35143,I35266,I35531);
not I_1950 (I35699,I2514);
DFFARX1 I_1951 (I658859,I2507,I35699,I35725,);
not I_1952 (I35733,I35725);
nand I_1953 (I35750,I658853,I658874);
and I_1954 (I35767,I35750,I658865);
DFFARX1 I_1955 (I35767,I2507,I35699,I35793,);
DFFARX1 I_1956 (I658856,I2507,I35699,I35810,);
and I_1957 (I35818,I35810,I658868);
nor I_1958 (I35835,I35793,I35818);
DFFARX1 I_1959 (I35835,I2507,I35699,I35667,);
nand I_1960 (I35866,I35810,I658868);
nand I_1961 (I35883,I35733,I35866);
not I_1962 (I35679,I35883);
DFFARX1 I_1963 (I658856,I2507,I35699,I35923,);
DFFARX1 I_1964 (I35923,I2507,I35699,I35688,);
nand I_1965 (I35945,I658877,I658862);
and I_1966 (I35962,I35945,I658853);
DFFARX1 I_1967 (I35962,I2507,I35699,I35988,);
DFFARX1 I_1968 (I35988,I2507,I35699,I36005,);
not I_1969 (I35691,I36005);
not I_1970 (I36027,I35988);
nand I_1971 (I35676,I36027,I35866);
nor I_1972 (I36058,I658871,I658862);
not I_1973 (I36075,I36058);
nor I_1974 (I36092,I36027,I36075);
nor I_1975 (I36109,I35733,I36092);
DFFARX1 I_1976 (I36109,I2507,I35699,I35685,);
nor I_1977 (I36140,I35793,I36075);
nor I_1978 (I35673,I35988,I36140);
nor I_1979 (I35682,I35923,I36058);
nor I_1980 (I35670,I35793,I36058);
not I_1981 (I36226,I2514);
DFFARX1 I_1982 (I26205,I2507,I36226,I36252,);
not I_1983 (I36260,I36252);
nand I_1984 (I36277,I26193,I26199);
and I_1985 (I36294,I36277,I26202);
DFFARX1 I_1986 (I36294,I2507,I36226,I36320,);
DFFARX1 I_1987 (I26184,I2507,I36226,I36337,);
and I_1988 (I36345,I36337,I26190);
nor I_1989 (I36362,I36320,I36345);
DFFARX1 I_1990 (I36362,I2507,I36226,I36194,);
nand I_1991 (I36393,I36337,I26190);
nand I_1992 (I36410,I36260,I36393);
not I_1993 (I36206,I36410);
DFFARX1 I_1994 (I26184,I2507,I36226,I36450,);
DFFARX1 I_1995 (I36450,I2507,I36226,I36215,);
nand I_1996 (I36472,I26187,I26181);
and I_1997 (I36489,I36472,I26196);
DFFARX1 I_1998 (I36489,I2507,I36226,I36515,);
DFFARX1 I_1999 (I36515,I2507,I36226,I36532,);
not I_2000 (I36218,I36532);
not I_2001 (I36554,I36515);
nand I_2002 (I36203,I36554,I36393);
nor I_2003 (I36585,I26181,I26181);
not I_2004 (I36602,I36585);
nor I_2005 (I36619,I36554,I36602);
nor I_2006 (I36636,I36260,I36619);
DFFARX1 I_2007 (I36636,I2507,I36226,I36212,);
nor I_2008 (I36667,I36320,I36602);
nor I_2009 (I36200,I36515,I36667);
nor I_2010 (I36209,I36450,I36585);
nor I_2011 (I36197,I36320,I36585);
not I_2012 (I36753,I2514);
DFFARX1 I_2013 (I154441,I2507,I36753,I36779,);
not I_2014 (I36787,I36779);
nand I_2015 (I36804,I154435,I154429);
and I_2016 (I36821,I36804,I154450);
DFFARX1 I_2017 (I36821,I2507,I36753,I36847,);
DFFARX1 I_2018 (I154447,I2507,I36753,I36864,);
and I_2019 (I36872,I36864,I154444);
nor I_2020 (I36889,I36847,I36872);
DFFARX1 I_2021 (I36889,I2507,I36753,I36721,);
nand I_2022 (I36920,I36864,I154444);
nand I_2023 (I36937,I36787,I36920);
not I_2024 (I36733,I36937);
DFFARX1 I_2025 (I154429,I2507,I36753,I36977,);
DFFARX1 I_2026 (I36977,I2507,I36753,I36742,);
nand I_2027 (I36999,I154432,I154432);
and I_2028 (I37016,I36999,I154453);
DFFARX1 I_2029 (I37016,I2507,I36753,I37042,);
DFFARX1 I_2030 (I37042,I2507,I36753,I37059,);
not I_2031 (I36745,I37059);
not I_2032 (I37081,I37042);
nand I_2033 (I36730,I37081,I36920);
nor I_2034 (I37112,I154438,I154432);
not I_2035 (I37129,I37112);
nor I_2036 (I37146,I37081,I37129);
nor I_2037 (I37163,I36787,I37146);
DFFARX1 I_2038 (I37163,I2507,I36753,I36739,);
nor I_2039 (I37194,I36847,I37129);
nor I_2040 (I36727,I37042,I37194);
nor I_2041 (I36736,I36977,I37112);
nor I_2042 (I36724,I36847,I37112);
not I_2043 (I37280,I2514);
DFFARX1 I_2044 (I158606,I2507,I37280,I37306,);
not I_2045 (I37314,I37306);
nand I_2046 (I37331,I158600,I158594);
and I_2047 (I37348,I37331,I158615);
DFFARX1 I_2048 (I37348,I2507,I37280,I37374,);
DFFARX1 I_2049 (I158612,I2507,I37280,I37391,);
and I_2050 (I37399,I37391,I158609);
nor I_2051 (I37416,I37374,I37399);
DFFARX1 I_2052 (I37416,I2507,I37280,I37248,);
nand I_2053 (I37447,I37391,I158609);
nand I_2054 (I37464,I37314,I37447);
not I_2055 (I37260,I37464);
DFFARX1 I_2056 (I158594,I2507,I37280,I37504,);
DFFARX1 I_2057 (I37504,I2507,I37280,I37269,);
nand I_2058 (I37526,I158597,I158597);
and I_2059 (I37543,I37526,I158618);
DFFARX1 I_2060 (I37543,I2507,I37280,I37569,);
DFFARX1 I_2061 (I37569,I2507,I37280,I37586,);
not I_2062 (I37272,I37586);
not I_2063 (I37608,I37569);
nand I_2064 (I37257,I37608,I37447);
nor I_2065 (I37639,I158603,I158597);
not I_2066 (I37656,I37639);
nor I_2067 (I37673,I37608,I37656);
nor I_2068 (I37690,I37314,I37673);
DFFARX1 I_2069 (I37690,I2507,I37280,I37266,);
nor I_2070 (I37721,I37374,I37656);
nor I_2071 (I37254,I37569,I37721);
nor I_2072 (I37263,I37504,I37639);
nor I_2073 (I37251,I37374,I37639);
not I_2074 (I37807,I2514);
DFFARX1 I_2075 (I224377,I2507,I37807,I37833,);
not I_2076 (I37841,I37833);
nand I_2077 (I37858,I224359,I224374);
and I_2078 (I37875,I37858,I224350);
DFFARX1 I_2079 (I37875,I2507,I37807,I37901,);
DFFARX1 I_2080 (I224353,I2507,I37807,I37918,);
and I_2081 (I37926,I37918,I224368);
nor I_2082 (I37943,I37901,I37926);
DFFARX1 I_2083 (I37943,I2507,I37807,I37775,);
nand I_2084 (I37974,I37918,I224368);
nand I_2085 (I37991,I37841,I37974);
not I_2086 (I37787,I37991);
DFFARX1 I_2087 (I224371,I2507,I37807,I38031,);
DFFARX1 I_2088 (I38031,I2507,I37807,I37796,);
nand I_2089 (I38053,I224350,I224362);
and I_2090 (I38070,I38053,I224356);
DFFARX1 I_2091 (I38070,I2507,I37807,I38096,);
DFFARX1 I_2092 (I38096,I2507,I37807,I38113,);
not I_2093 (I37799,I38113);
not I_2094 (I38135,I38096);
nand I_2095 (I37784,I38135,I37974);
nor I_2096 (I38166,I224365,I224362);
not I_2097 (I38183,I38166);
nor I_2098 (I38200,I38135,I38183);
nor I_2099 (I38217,I37841,I38200);
DFFARX1 I_2100 (I38217,I2507,I37807,I37793,);
nor I_2101 (I38248,I37901,I38183);
nor I_2102 (I37781,I38096,I38248);
nor I_2103 (I37790,I38031,I38166);
nor I_2104 (I37778,I37901,I38166);
not I_2105 (I38334,I2514);
DFFARX1 I_2106 (I314884,I2507,I38334,I38360,);
not I_2107 (I38368,I38360);
nand I_2108 (I38385,I314896,I314881);
and I_2109 (I38402,I38385,I314875);
DFFARX1 I_2110 (I38402,I2507,I38334,I38428,);
DFFARX1 I_2111 (I314890,I2507,I38334,I38445,);
and I_2112 (I38453,I38445,I314878);
nor I_2113 (I38470,I38428,I38453);
DFFARX1 I_2114 (I38470,I2507,I38334,I38302,);
nand I_2115 (I38501,I38445,I314878);
nand I_2116 (I38518,I38368,I38501);
not I_2117 (I38314,I38518);
DFFARX1 I_2118 (I314887,I2507,I38334,I38558,);
DFFARX1 I_2119 (I38558,I2507,I38334,I38323,);
nand I_2120 (I38580,I314893,I314899);
and I_2121 (I38597,I38580,I314875);
DFFARX1 I_2122 (I38597,I2507,I38334,I38623,);
DFFARX1 I_2123 (I38623,I2507,I38334,I38640,);
not I_2124 (I38326,I38640);
not I_2125 (I38662,I38623);
nand I_2126 (I38311,I38662,I38501);
nor I_2127 (I38693,I314878,I314899);
not I_2128 (I38710,I38693);
nor I_2129 (I38727,I38662,I38710);
nor I_2130 (I38744,I38368,I38727);
DFFARX1 I_2131 (I38744,I2507,I38334,I38320,);
nor I_2132 (I38775,I38428,I38710);
nor I_2133 (I38308,I38623,I38775);
nor I_2134 (I38317,I38558,I38693);
nor I_2135 (I38305,I38428,I38693);
not I_2136 (I38861,I2514);
DFFARX1 I_2137 (I337426,I2507,I38861,I38887,);
not I_2138 (I38895,I38887);
nand I_2139 (I38912,I337438,I337423);
and I_2140 (I38929,I38912,I337417);
DFFARX1 I_2141 (I38929,I2507,I38861,I38955,);
DFFARX1 I_2142 (I337432,I2507,I38861,I38972,);
and I_2143 (I38980,I38972,I337420);
nor I_2144 (I38997,I38955,I38980);
DFFARX1 I_2145 (I38997,I2507,I38861,I38829,);
nand I_2146 (I39028,I38972,I337420);
nand I_2147 (I39045,I38895,I39028);
not I_2148 (I38841,I39045);
DFFARX1 I_2149 (I337429,I2507,I38861,I39085,);
DFFARX1 I_2150 (I39085,I2507,I38861,I38850,);
nand I_2151 (I39107,I337435,I337441);
and I_2152 (I39124,I39107,I337417);
DFFARX1 I_2153 (I39124,I2507,I38861,I39150,);
DFFARX1 I_2154 (I39150,I2507,I38861,I39167,);
not I_2155 (I38853,I39167);
not I_2156 (I39189,I39150);
nand I_2157 (I38838,I39189,I39028);
nor I_2158 (I39220,I337420,I337441);
not I_2159 (I39237,I39220);
nor I_2160 (I39254,I39189,I39237);
nor I_2161 (I39271,I38895,I39254);
DFFARX1 I_2162 (I39271,I2507,I38861,I38847,);
nor I_2163 (I39302,I38955,I39237);
nor I_2164 (I38835,I39150,I39302);
nor I_2165 (I38844,I39085,I39220);
nor I_2166 (I38832,I38955,I39220);
not I_2167 (I39388,I2514);
DFFARX1 I_2168 (I478305,I2507,I39388,I39414,);
not I_2169 (I39422,I39414);
nand I_2170 (I39439,I478323,I478317);
and I_2171 (I39456,I39439,I478296);
DFFARX1 I_2172 (I39456,I2507,I39388,I39482,);
DFFARX1 I_2173 (I478314,I2507,I39388,I39499,);
and I_2174 (I39507,I39499,I478299);
nor I_2175 (I39524,I39482,I39507);
DFFARX1 I_2176 (I39524,I2507,I39388,I39356,);
nand I_2177 (I39555,I39499,I478299);
nand I_2178 (I39572,I39422,I39555);
not I_2179 (I39368,I39572);
DFFARX1 I_2180 (I478311,I2507,I39388,I39612,);
DFFARX1 I_2181 (I39612,I2507,I39388,I39377,);
nand I_2182 (I39634,I478320,I478308);
and I_2183 (I39651,I39634,I478302);
DFFARX1 I_2184 (I39651,I2507,I39388,I39677,);
DFFARX1 I_2185 (I39677,I2507,I39388,I39694,);
not I_2186 (I39380,I39694);
not I_2187 (I39716,I39677);
nand I_2188 (I39365,I39716,I39555);
nor I_2189 (I39747,I478296,I478308);
not I_2190 (I39764,I39747);
nor I_2191 (I39781,I39716,I39764);
nor I_2192 (I39798,I39422,I39781);
DFFARX1 I_2193 (I39798,I2507,I39388,I39374,);
nor I_2194 (I39829,I39482,I39764);
nor I_2195 (I39362,I39677,I39829);
nor I_2196 (I39371,I39612,I39747);
nor I_2197 (I39359,I39482,I39747);
not I_2198 (I39915,I2514);
DFFARX1 I_2199 (I102676,I2507,I39915,I39941,);
not I_2200 (I39949,I39941);
nand I_2201 (I39966,I102670,I102664);
and I_2202 (I39983,I39966,I102685);
DFFARX1 I_2203 (I39983,I2507,I39915,I40009,);
DFFARX1 I_2204 (I102682,I2507,I39915,I40026,);
and I_2205 (I40034,I40026,I102679);
nor I_2206 (I40051,I40009,I40034);
DFFARX1 I_2207 (I40051,I2507,I39915,I39883,);
nand I_2208 (I40082,I40026,I102679);
nand I_2209 (I40099,I39949,I40082);
not I_2210 (I39895,I40099);
DFFARX1 I_2211 (I102664,I2507,I39915,I40139,);
DFFARX1 I_2212 (I40139,I2507,I39915,I39904,);
nand I_2213 (I40161,I102667,I102667);
and I_2214 (I40178,I40161,I102688);
DFFARX1 I_2215 (I40178,I2507,I39915,I40204,);
DFFARX1 I_2216 (I40204,I2507,I39915,I40221,);
not I_2217 (I39907,I40221);
not I_2218 (I40243,I40204);
nand I_2219 (I39892,I40243,I40082);
nor I_2220 (I40274,I102673,I102667);
not I_2221 (I40291,I40274);
nor I_2222 (I40308,I40243,I40291);
nor I_2223 (I40325,I39949,I40308);
DFFARX1 I_2224 (I40325,I2507,I39915,I39901,);
nor I_2225 (I40356,I40009,I40291);
nor I_2226 (I39889,I40204,I40356);
nor I_2227 (I39898,I40139,I40274);
nor I_2228 (I39886,I40009,I40274);
not I_2229 (I40442,I2514);
DFFARX1 I_2230 (I105056,I2507,I40442,I40468,);
not I_2231 (I40476,I40468);
nand I_2232 (I40493,I105050,I105044);
and I_2233 (I40510,I40493,I105065);
DFFARX1 I_2234 (I40510,I2507,I40442,I40536,);
DFFARX1 I_2235 (I105062,I2507,I40442,I40553,);
and I_2236 (I40561,I40553,I105059);
nor I_2237 (I40578,I40536,I40561);
DFFARX1 I_2238 (I40578,I2507,I40442,I40410,);
nand I_2239 (I40609,I40553,I105059);
nand I_2240 (I40626,I40476,I40609);
not I_2241 (I40422,I40626);
DFFARX1 I_2242 (I105044,I2507,I40442,I40666,);
DFFARX1 I_2243 (I40666,I2507,I40442,I40431,);
nand I_2244 (I40688,I105047,I105047);
and I_2245 (I40705,I40688,I105068);
DFFARX1 I_2246 (I40705,I2507,I40442,I40731,);
DFFARX1 I_2247 (I40731,I2507,I40442,I40748,);
not I_2248 (I40434,I40748);
not I_2249 (I40770,I40731);
nand I_2250 (I40419,I40770,I40609);
nor I_2251 (I40801,I105053,I105047);
not I_2252 (I40818,I40801);
nor I_2253 (I40835,I40770,I40818);
nor I_2254 (I40852,I40476,I40835);
DFFARX1 I_2255 (I40852,I2507,I40442,I40428,);
nor I_2256 (I40883,I40536,I40818);
nor I_2257 (I40416,I40731,I40883);
nor I_2258 (I40425,I40666,I40801);
nor I_2259 (I40413,I40536,I40801);
not I_2260 (I40969,I2514);
DFFARX1 I_2261 (I366907,I2507,I40969,I40995,);
not I_2262 (I41003,I40995);
nand I_2263 (I41020,I366898,I366916);
and I_2264 (I41037,I41020,I366895);
DFFARX1 I_2265 (I41037,I2507,I40969,I41063,);
DFFARX1 I_2266 (I366898,I2507,I40969,I41080,);
and I_2267 (I41088,I41080,I366901);
nor I_2268 (I41105,I41063,I41088);
DFFARX1 I_2269 (I41105,I2507,I40969,I40937,);
nand I_2270 (I41136,I41080,I366901);
nand I_2271 (I41153,I41003,I41136);
not I_2272 (I40949,I41153);
DFFARX1 I_2273 (I366895,I2507,I40969,I41193,);
DFFARX1 I_2274 (I41193,I2507,I40969,I40958,);
nand I_2275 (I41215,I366913,I366904);
and I_2276 (I41232,I41215,I366919);
DFFARX1 I_2277 (I41232,I2507,I40969,I41258,);
DFFARX1 I_2278 (I41258,I2507,I40969,I41275,);
not I_2279 (I40961,I41275);
not I_2280 (I41297,I41258);
nand I_2281 (I40946,I41297,I41136);
nor I_2282 (I41328,I366910,I366904);
not I_2283 (I41345,I41328);
nor I_2284 (I41362,I41297,I41345);
nor I_2285 (I41379,I41003,I41362);
DFFARX1 I_2286 (I41379,I2507,I40969,I40955,);
nor I_2287 (I41410,I41063,I41345);
nor I_2288 (I40943,I41258,I41410);
nor I_2289 (I40952,I41193,I41328);
nor I_2290 (I40940,I41063,I41328);
not I_2291 (I41496,I2514);
DFFARX1 I_2292 (I112791,I2507,I41496,I41522,);
not I_2293 (I41530,I41522);
nand I_2294 (I41547,I112785,I112779);
and I_2295 (I41564,I41547,I112800);
DFFARX1 I_2296 (I41564,I2507,I41496,I41590,);
DFFARX1 I_2297 (I112797,I2507,I41496,I41607,);
and I_2298 (I41615,I41607,I112794);
nor I_2299 (I41632,I41590,I41615);
DFFARX1 I_2300 (I41632,I2507,I41496,I41464,);
nand I_2301 (I41663,I41607,I112794);
nand I_2302 (I41680,I41530,I41663);
not I_2303 (I41476,I41680);
DFFARX1 I_2304 (I112779,I2507,I41496,I41720,);
DFFARX1 I_2305 (I41720,I2507,I41496,I41485,);
nand I_2306 (I41742,I112782,I112782);
and I_2307 (I41759,I41742,I112803);
DFFARX1 I_2308 (I41759,I2507,I41496,I41785,);
DFFARX1 I_2309 (I41785,I2507,I41496,I41802,);
not I_2310 (I41488,I41802);
not I_2311 (I41824,I41785);
nand I_2312 (I41473,I41824,I41663);
nor I_2313 (I41855,I112788,I112782);
not I_2314 (I41872,I41855);
nor I_2315 (I41889,I41824,I41872);
nor I_2316 (I41906,I41530,I41889);
DFFARX1 I_2317 (I41906,I2507,I41496,I41482,);
nor I_2318 (I41937,I41590,I41872);
nor I_2319 (I41470,I41785,I41937);
nor I_2320 (I41479,I41720,I41855);
nor I_2321 (I41467,I41590,I41855);
not I_2322 (I42023,I2514);
DFFARX1 I_2323 (I199081,I2507,I42023,I42049,);
not I_2324 (I42057,I42049);
nand I_2325 (I42074,I199063,I199078);
and I_2326 (I42091,I42074,I199054);
DFFARX1 I_2327 (I42091,I2507,I42023,I42117,);
DFFARX1 I_2328 (I199057,I2507,I42023,I42134,);
and I_2329 (I42142,I42134,I199072);
nor I_2330 (I42159,I42117,I42142);
DFFARX1 I_2331 (I42159,I2507,I42023,I41991,);
nand I_2332 (I42190,I42134,I199072);
nand I_2333 (I42207,I42057,I42190);
not I_2334 (I42003,I42207);
DFFARX1 I_2335 (I199075,I2507,I42023,I42247,);
DFFARX1 I_2336 (I42247,I2507,I42023,I42012,);
nand I_2337 (I42269,I199054,I199066);
and I_2338 (I42286,I42269,I199060);
DFFARX1 I_2339 (I42286,I2507,I42023,I42312,);
DFFARX1 I_2340 (I42312,I2507,I42023,I42329,);
not I_2341 (I42015,I42329);
not I_2342 (I42351,I42312);
nand I_2343 (I42000,I42351,I42190);
nor I_2344 (I42382,I199069,I199066);
not I_2345 (I42399,I42382);
nor I_2346 (I42416,I42351,I42399);
nor I_2347 (I42433,I42057,I42416);
DFFARX1 I_2348 (I42433,I2507,I42023,I42009,);
nor I_2349 (I42464,I42117,I42399);
nor I_2350 (I41997,I42312,I42464);
nor I_2351 (I42006,I42247,I42382);
nor I_2352 (I41994,I42117,I42382);
not I_2353 (I42550,I2514);
DFFARX1 I_2354 (I189595,I2507,I42550,I42576,);
not I_2355 (I42584,I42576);
nand I_2356 (I42601,I189577,I189592);
and I_2357 (I42618,I42601,I189568);
DFFARX1 I_2358 (I42618,I2507,I42550,I42644,);
DFFARX1 I_2359 (I189571,I2507,I42550,I42661,);
and I_2360 (I42669,I42661,I189586);
nor I_2361 (I42686,I42644,I42669);
DFFARX1 I_2362 (I42686,I2507,I42550,I42518,);
nand I_2363 (I42717,I42661,I189586);
nand I_2364 (I42734,I42584,I42717);
not I_2365 (I42530,I42734);
DFFARX1 I_2366 (I189589,I2507,I42550,I42774,);
DFFARX1 I_2367 (I42774,I2507,I42550,I42539,);
nand I_2368 (I42796,I189568,I189580);
and I_2369 (I42813,I42796,I189574);
DFFARX1 I_2370 (I42813,I2507,I42550,I42839,);
DFFARX1 I_2371 (I42839,I2507,I42550,I42856,);
not I_2372 (I42542,I42856);
not I_2373 (I42878,I42839);
nand I_2374 (I42527,I42878,I42717);
nor I_2375 (I42909,I189583,I189580);
not I_2376 (I42926,I42909);
nor I_2377 (I42943,I42878,I42926);
nor I_2378 (I42960,I42584,I42943);
DFFARX1 I_2379 (I42960,I2507,I42550,I42536,);
nor I_2380 (I42991,I42644,I42926);
nor I_2381 (I42524,I42839,I42991);
nor I_2382 (I42533,I42774,I42909);
nor I_2383 (I42521,I42644,I42909);
not I_2384 (I43077,I2514);
DFFARX1 I_2385 (I587867,I2507,I43077,I43103,);
not I_2386 (I43111,I43103);
nand I_2387 (I43128,I587882,I587861);
and I_2388 (I43145,I43128,I587864);
DFFARX1 I_2389 (I43145,I2507,I43077,I43171,);
DFFARX1 I_2390 (I587885,I2507,I43077,I43188,);
and I_2391 (I43196,I43188,I587864);
nor I_2392 (I43213,I43171,I43196);
DFFARX1 I_2393 (I43213,I2507,I43077,I43045,);
nand I_2394 (I43244,I43188,I587864);
nand I_2395 (I43261,I43111,I43244);
not I_2396 (I43057,I43261);
DFFARX1 I_2397 (I587861,I2507,I43077,I43301,);
DFFARX1 I_2398 (I43301,I2507,I43077,I43066,);
nand I_2399 (I43323,I587873,I587870);
and I_2400 (I43340,I43323,I587876);
DFFARX1 I_2401 (I43340,I2507,I43077,I43366,);
DFFARX1 I_2402 (I43366,I2507,I43077,I43383,);
not I_2403 (I43069,I43383);
not I_2404 (I43405,I43366);
nand I_2405 (I43054,I43405,I43244);
nor I_2406 (I43436,I587879,I587870);
not I_2407 (I43453,I43436);
nor I_2408 (I43470,I43405,I43453);
nor I_2409 (I43487,I43111,I43470);
DFFARX1 I_2410 (I43487,I2507,I43077,I43063,);
nor I_2411 (I43518,I43171,I43453);
nor I_2412 (I43051,I43366,I43518);
nor I_2413 (I43060,I43301,I43436);
nor I_2414 (I43048,I43171,I43436);
not I_2415 (I43604,I2514);
DFFARX1 I_2416 (I342050,I2507,I43604,I43630,);
not I_2417 (I43638,I43630);
nand I_2418 (I43655,I342062,I342047);
and I_2419 (I43672,I43655,I342041);
DFFARX1 I_2420 (I43672,I2507,I43604,I43698,);
DFFARX1 I_2421 (I342056,I2507,I43604,I43715,);
and I_2422 (I43723,I43715,I342044);
nor I_2423 (I43740,I43698,I43723);
DFFARX1 I_2424 (I43740,I2507,I43604,I43572,);
nand I_2425 (I43771,I43715,I342044);
nand I_2426 (I43788,I43638,I43771);
not I_2427 (I43584,I43788);
DFFARX1 I_2428 (I342053,I2507,I43604,I43828,);
DFFARX1 I_2429 (I43828,I2507,I43604,I43593,);
nand I_2430 (I43850,I342059,I342065);
and I_2431 (I43867,I43850,I342041);
DFFARX1 I_2432 (I43867,I2507,I43604,I43893,);
DFFARX1 I_2433 (I43893,I2507,I43604,I43910,);
not I_2434 (I43596,I43910);
not I_2435 (I43932,I43893);
nand I_2436 (I43581,I43932,I43771);
nor I_2437 (I43963,I342044,I342065);
not I_2438 (I43980,I43963);
nor I_2439 (I43997,I43932,I43980);
nor I_2440 (I44014,I43638,I43997);
DFFARX1 I_2441 (I44014,I2507,I43604,I43590,);
nor I_2442 (I44045,I43698,I43980);
nor I_2443 (I43578,I43893,I44045);
nor I_2444 (I43587,I43828,I43963);
nor I_2445 (I43575,I43698,I43963);
not I_2446 (I44131,I2514);
DFFARX1 I_2447 (I365173,I2507,I44131,I44157,);
not I_2448 (I44165,I44157);
nand I_2449 (I44182,I365164,I365182);
and I_2450 (I44199,I44182,I365161);
DFFARX1 I_2451 (I44199,I2507,I44131,I44225,);
DFFARX1 I_2452 (I365164,I2507,I44131,I44242,);
and I_2453 (I44250,I44242,I365167);
nor I_2454 (I44267,I44225,I44250);
DFFARX1 I_2455 (I44267,I2507,I44131,I44099,);
nand I_2456 (I44298,I44242,I365167);
nand I_2457 (I44315,I44165,I44298);
not I_2458 (I44111,I44315);
DFFARX1 I_2459 (I365161,I2507,I44131,I44355,);
DFFARX1 I_2460 (I44355,I2507,I44131,I44120,);
nand I_2461 (I44377,I365179,I365170);
and I_2462 (I44394,I44377,I365185);
DFFARX1 I_2463 (I44394,I2507,I44131,I44420,);
DFFARX1 I_2464 (I44420,I2507,I44131,I44437,);
not I_2465 (I44123,I44437);
not I_2466 (I44459,I44420);
nand I_2467 (I44108,I44459,I44298);
nor I_2468 (I44490,I365176,I365170);
not I_2469 (I44507,I44490);
nor I_2470 (I44524,I44459,I44507);
nor I_2471 (I44541,I44165,I44524);
DFFARX1 I_2472 (I44541,I2507,I44131,I44117,);
nor I_2473 (I44572,I44225,I44507);
nor I_2474 (I44105,I44420,I44572);
nor I_2475 (I44114,I44355,I44490);
nor I_2476 (I44102,I44225,I44490);
not I_2477 (I44658,I2514);
DFFARX1 I_2478 (I5507,I2507,I44658,I44684,);
not I_2479 (I44692,I44684);
nand I_2480 (I44709,I5492,I5492);
and I_2481 (I44726,I44709,I5513);
DFFARX1 I_2482 (I44726,I2507,I44658,I44752,);
DFFARX1 I_2483 (I5495,I2507,I44658,I44769,);
and I_2484 (I44777,I44769,I5504);
nor I_2485 (I44794,I44752,I44777);
DFFARX1 I_2486 (I44794,I2507,I44658,I44626,);
nand I_2487 (I44825,I44769,I5504);
nand I_2488 (I44842,I44692,I44825);
not I_2489 (I44638,I44842);
DFFARX1 I_2490 (I5498,I2507,I44658,I44882,);
DFFARX1 I_2491 (I44882,I2507,I44658,I44647,);
nand I_2492 (I44904,I5501,I5510);
and I_2493 (I44921,I44904,I5495);
DFFARX1 I_2494 (I44921,I2507,I44658,I44947,);
DFFARX1 I_2495 (I44947,I2507,I44658,I44964,);
not I_2496 (I44650,I44964);
not I_2497 (I44986,I44947);
nand I_2498 (I44635,I44986,I44825);
nor I_2499 (I45017,I5498,I5510);
not I_2500 (I45034,I45017);
nor I_2501 (I45051,I44986,I45034);
nor I_2502 (I45068,I44692,I45051);
DFFARX1 I_2503 (I45068,I2507,I44658,I44644,);
nor I_2504 (I45099,I44752,I45034);
nor I_2505 (I44632,I44947,I45099);
nor I_2506 (I44641,I44882,I45017);
nor I_2507 (I44629,I44752,I45017);
not I_2508 (I45185,I2514);
DFFARX1 I_2509 (I429175,I2507,I45185,I45211,);
not I_2510 (I45219,I45211);
nand I_2511 (I45236,I429172,I429187);
and I_2512 (I45253,I45236,I429169);
DFFARX1 I_2513 (I45253,I2507,I45185,I45279,);
DFFARX1 I_2514 (I429166,I2507,I45185,I45296,);
and I_2515 (I45304,I45296,I429166);
nor I_2516 (I45321,I45279,I45304);
DFFARX1 I_2517 (I45321,I2507,I45185,I45153,);
nand I_2518 (I45352,I45296,I429166);
nand I_2519 (I45369,I45219,I45352);
not I_2520 (I45165,I45369);
DFFARX1 I_2521 (I429169,I2507,I45185,I45409,);
DFFARX1 I_2522 (I45409,I2507,I45185,I45174,);
nand I_2523 (I45431,I429181,I429172);
and I_2524 (I45448,I45431,I429184);
DFFARX1 I_2525 (I45448,I2507,I45185,I45474,);
DFFARX1 I_2526 (I45474,I2507,I45185,I45491,);
not I_2527 (I45177,I45491);
not I_2528 (I45513,I45474);
nand I_2529 (I45162,I45513,I45352);
nor I_2530 (I45544,I429178,I429172);
not I_2531 (I45561,I45544);
nor I_2532 (I45578,I45513,I45561);
nor I_2533 (I45595,I45219,I45578);
DFFARX1 I_2534 (I45595,I2507,I45185,I45171,);
nor I_2535 (I45626,I45279,I45561);
nor I_2536 (I45159,I45474,I45626);
nor I_2537 (I45168,I45409,I45544);
nor I_2538 (I45156,I45279,I45544);
not I_2539 (I45712,I2514);
DFFARX1 I_2540 (I642539,I2507,I45712,I45738,);
not I_2541 (I45746,I45738);
nand I_2542 (I45763,I642533,I642554);
and I_2543 (I45780,I45763,I642545);
DFFARX1 I_2544 (I45780,I2507,I45712,I45806,);
DFFARX1 I_2545 (I642536,I2507,I45712,I45823,);
and I_2546 (I45831,I45823,I642548);
nor I_2547 (I45848,I45806,I45831);
DFFARX1 I_2548 (I45848,I2507,I45712,I45680,);
nand I_2549 (I45879,I45823,I642548);
nand I_2550 (I45896,I45746,I45879);
not I_2551 (I45692,I45896);
DFFARX1 I_2552 (I642536,I2507,I45712,I45936,);
DFFARX1 I_2553 (I45936,I2507,I45712,I45701,);
nand I_2554 (I45958,I642557,I642542);
and I_2555 (I45975,I45958,I642533);
DFFARX1 I_2556 (I45975,I2507,I45712,I46001,);
DFFARX1 I_2557 (I46001,I2507,I45712,I46018,);
not I_2558 (I45704,I46018);
not I_2559 (I46040,I46001);
nand I_2560 (I45689,I46040,I45879);
nor I_2561 (I46071,I642551,I642542);
not I_2562 (I46088,I46071);
nor I_2563 (I46105,I46040,I46088);
nor I_2564 (I46122,I45746,I46105);
DFFARX1 I_2565 (I46122,I2507,I45712,I45698,);
nor I_2566 (I46153,I45806,I46088);
nor I_2567 (I45686,I46001,I46153);
nor I_2568 (I45695,I45936,I46071);
nor I_2569 (I45683,I45806,I46071);
not I_2570 (I46239,I2514);
DFFARX1 I_2571 (I214891,I2507,I46239,I46265,);
not I_2572 (I46273,I46265);
nand I_2573 (I46290,I214873,I214888);
and I_2574 (I46307,I46290,I214864);
DFFARX1 I_2575 (I46307,I2507,I46239,I46333,);
DFFARX1 I_2576 (I214867,I2507,I46239,I46350,);
and I_2577 (I46358,I46350,I214882);
nor I_2578 (I46375,I46333,I46358);
DFFARX1 I_2579 (I46375,I2507,I46239,I46207,);
nand I_2580 (I46406,I46350,I214882);
nand I_2581 (I46423,I46273,I46406);
not I_2582 (I46219,I46423);
DFFARX1 I_2583 (I214885,I2507,I46239,I46463,);
DFFARX1 I_2584 (I46463,I2507,I46239,I46228,);
nand I_2585 (I46485,I214864,I214876);
and I_2586 (I46502,I46485,I214870);
DFFARX1 I_2587 (I46502,I2507,I46239,I46528,);
DFFARX1 I_2588 (I46528,I2507,I46239,I46545,);
not I_2589 (I46231,I46545);
not I_2590 (I46567,I46528);
nand I_2591 (I46216,I46567,I46406);
nor I_2592 (I46598,I214879,I214876);
not I_2593 (I46615,I46598);
nor I_2594 (I46632,I46567,I46615);
nor I_2595 (I46649,I46273,I46632);
DFFARX1 I_2596 (I46649,I2507,I46239,I46225,);
nor I_2597 (I46680,I46333,I46615);
nor I_2598 (I46213,I46528,I46680);
nor I_2599 (I46222,I46463,I46598);
nor I_2600 (I46210,I46333,I46598);
not I_2601 (I46766,I2514);
DFFARX1 I_2602 (I27259,I2507,I46766,I46792,);
not I_2603 (I46800,I46792);
nand I_2604 (I46817,I27247,I27253);
and I_2605 (I46834,I46817,I27256);
DFFARX1 I_2606 (I46834,I2507,I46766,I46860,);
DFFARX1 I_2607 (I27238,I2507,I46766,I46877,);
and I_2608 (I46885,I46877,I27244);
nor I_2609 (I46902,I46860,I46885);
DFFARX1 I_2610 (I46902,I2507,I46766,I46734,);
nand I_2611 (I46933,I46877,I27244);
nand I_2612 (I46950,I46800,I46933);
not I_2613 (I46746,I46950);
DFFARX1 I_2614 (I27238,I2507,I46766,I46990,);
DFFARX1 I_2615 (I46990,I2507,I46766,I46755,);
nand I_2616 (I47012,I27241,I27235);
and I_2617 (I47029,I47012,I27250);
DFFARX1 I_2618 (I47029,I2507,I46766,I47055,);
DFFARX1 I_2619 (I47055,I2507,I46766,I47072,);
not I_2620 (I46758,I47072);
not I_2621 (I47094,I47055);
nand I_2622 (I46743,I47094,I46933);
nor I_2623 (I47125,I27235,I27235);
not I_2624 (I47142,I47125);
nor I_2625 (I47159,I47094,I47142);
nor I_2626 (I47176,I46800,I47159);
DFFARX1 I_2627 (I47176,I2507,I46766,I46752,);
nor I_2628 (I47207,I46860,I47142);
nor I_2629 (I46740,I47055,I47207);
nor I_2630 (I46749,I46990,I47125);
nor I_2631 (I46737,I46860,I47125);
not I_2632 (I47293,I2514);
DFFARX1 I_2633 (I139566,I2507,I47293,I47319,);
not I_2634 (I47327,I47319);
nand I_2635 (I47344,I139560,I139554);
and I_2636 (I47361,I47344,I139575);
DFFARX1 I_2637 (I47361,I2507,I47293,I47387,);
DFFARX1 I_2638 (I139572,I2507,I47293,I47404,);
and I_2639 (I47412,I47404,I139569);
nor I_2640 (I47429,I47387,I47412);
DFFARX1 I_2641 (I47429,I2507,I47293,I47261,);
nand I_2642 (I47460,I47404,I139569);
nand I_2643 (I47477,I47327,I47460);
not I_2644 (I47273,I47477);
DFFARX1 I_2645 (I139554,I2507,I47293,I47517,);
DFFARX1 I_2646 (I47517,I2507,I47293,I47282,);
nand I_2647 (I47539,I139557,I139557);
and I_2648 (I47556,I47539,I139578);
DFFARX1 I_2649 (I47556,I2507,I47293,I47582,);
DFFARX1 I_2650 (I47582,I2507,I47293,I47599,);
not I_2651 (I47285,I47599);
not I_2652 (I47621,I47582);
nand I_2653 (I47270,I47621,I47460);
nor I_2654 (I47652,I139563,I139557);
not I_2655 (I47669,I47652);
nor I_2656 (I47686,I47621,I47669);
nor I_2657 (I47703,I47327,I47686);
DFFARX1 I_2658 (I47703,I2507,I47293,I47279,);
nor I_2659 (I47734,I47387,I47669);
nor I_2660 (I47267,I47582,I47734);
nor I_2661 (I47276,I47517,I47652);
nor I_2662 (I47264,I47387,I47652);
not I_2663 (I47820,I2514);
DFFARX1 I_2664 (I173785,I2507,I47820,I47846,);
not I_2665 (I47854,I47846);
nand I_2666 (I47871,I173767,I173782);
and I_2667 (I47888,I47871,I173758);
DFFARX1 I_2668 (I47888,I2507,I47820,I47914,);
DFFARX1 I_2669 (I173761,I2507,I47820,I47931,);
and I_2670 (I47939,I47931,I173776);
nor I_2671 (I47956,I47914,I47939);
DFFARX1 I_2672 (I47956,I2507,I47820,I47788,);
nand I_2673 (I47987,I47931,I173776);
nand I_2674 (I48004,I47854,I47987);
not I_2675 (I47800,I48004);
DFFARX1 I_2676 (I173779,I2507,I47820,I48044,);
DFFARX1 I_2677 (I48044,I2507,I47820,I47809,);
nand I_2678 (I48066,I173758,I173770);
and I_2679 (I48083,I48066,I173764);
DFFARX1 I_2680 (I48083,I2507,I47820,I48109,);
DFFARX1 I_2681 (I48109,I2507,I47820,I48126,);
not I_2682 (I47812,I48126);
not I_2683 (I48148,I48109);
nand I_2684 (I47797,I48148,I47987);
nor I_2685 (I48179,I173773,I173770);
not I_2686 (I48196,I48179);
nor I_2687 (I48213,I48148,I48196);
nor I_2688 (I48230,I47854,I48213);
DFFARX1 I_2689 (I48230,I2507,I47820,I47806,);
nor I_2690 (I48261,I47914,I48196);
nor I_2691 (I47794,I48109,I48261);
nor I_2692 (I47803,I48044,I48179);
nor I_2693 (I47791,I47914,I48179);
not I_2694 (I48347,I2514);
DFFARX1 I_2695 (I372109,I2507,I48347,I48373,);
not I_2696 (I48381,I48373);
nand I_2697 (I48398,I372100,I372118);
and I_2698 (I48415,I48398,I372097);
DFFARX1 I_2699 (I48415,I2507,I48347,I48441,);
DFFARX1 I_2700 (I372100,I2507,I48347,I48458,);
and I_2701 (I48466,I48458,I372103);
nor I_2702 (I48483,I48441,I48466);
DFFARX1 I_2703 (I48483,I2507,I48347,I48315,);
nand I_2704 (I48514,I48458,I372103);
nand I_2705 (I48531,I48381,I48514);
not I_2706 (I48327,I48531);
DFFARX1 I_2707 (I372097,I2507,I48347,I48571,);
DFFARX1 I_2708 (I48571,I2507,I48347,I48336,);
nand I_2709 (I48593,I372115,I372106);
and I_2710 (I48610,I48593,I372121);
DFFARX1 I_2711 (I48610,I2507,I48347,I48636,);
DFFARX1 I_2712 (I48636,I2507,I48347,I48653,);
not I_2713 (I48339,I48653);
not I_2714 (I48675,I48636);
nand I_2715 (I48324,I48675,I48514);
nor I_2716 (I48706,I372112,I372106);
not I_2717 (I48723,I48706);
nor I_2718 (I48740,I48675,I48723);
nor I_2719 (I48757,I48381,I48740);
DFFARX1 I_2720 (I48757,I2507,I48347,I48333,);
nor I_2721 (I48788,I48441,I48723);
nor I_2722 (I48321,I48636,I48788);
nor I_2723 (I48330,I48571,I48706);
nor I_2724 (I48318,I48441,I48706);
not I_2725 (I48874,I2514);
DFFARX1 I_2726 (I32002,I2507,I48874,I48900,);
not I_2727 (I48908,I48900);
nand I_2728 (I48925,I31990,I31996);
and I_2729 (I48942,I48925,I31999);
DFFARX1 I_2730 (I48942,I2507,I48874,I48968,);
DFFARX1 I_2731 (I31981,I2507,I48874,I48985,);
and I_2732 (I48993,I48985,I31987);
nor I_2733 (I49010,I48968,I48993);
DFFARX1 I_2734 (I49010,I2507,I48874,I48842,);
nand I_2735 (I49041,I48985,I31987);
nand I_2736 (I49058,I48908,I49041);
not I_2737 (I48854,I49058);
DFFARX1 I_2738 (I31981,I2507,I48874,I49098,);
DFFARX1 I_2739 (I49098,I2507,I48874,I48863,);
nand I_2740 (I49120,I31984,I31978);
and I_2741 (I49137,I49120,I31993);
DFFARX1 I_2742 (I49137,I2507,I48874,I49163,);
DFFARX1 I_2743 (I49163,I2507,I48874,I49180,);
not I_2744 (I48866,I49180);
not I_2745 (I49202,I49163);
nand I_2746 (I48851,I49202,I49041);
nor I_2747 (I49233,I31978,I31978);
not I_2748 (I49250,I49233);
nor I_2749 (I49267,I49202,I49250);
nor I_2750 (I49284,I48908,I49267);
DFFARX1 I_2751 (I49284,I2507,I48874,I48860,);
nor I_2752 (I49315,I48968,I49250);
nor I_2753 (I48848,I49163,I49315);
nor I_2754 (I48857,I49098,I49233);
nor I_2755 (I48845,I48968,I49233);
not I_2756 (I49401,I2514);
DFFARX1 I_2757 (I260170,I2507,I49401,I49427,);
not I_2758 (I49435,I49427);
nand I_2759 (I49452,I260164,I260155);
and I_2760 (I49469,I49452,I260176);
DFFARX1 I_2761 (I49469,I2507,I49401,I49495,);
DFFARX1 I_2762 (I260158,I2507,I49401,I49512,);
and I_2763 (I49520,I49512,I260152);
nor I_2764 (I49537,I49495,I49520);
DFFARX1 I_2765 (I49537,I2507,I49401,I49369,);
nand I_2766 (I49568,I49512,I260152);
nand I_2767 (I49585,I49435,I49568);
not I_2768 (I49381,I49585);
DFFARX1 I_2769 (I260152,I2507,I49401,I49625,);
DFFARX1 I_2770 (I49625,I2507,I49401,I49390,);
nand I_2771 (I49647,I260179,I260161);
and I_2772 (I49664,I49647,I260167);
DFFARX1 I_2773 (I49664,I2507,I49401,I49690,);
DFFARX1 I_2774 (I49690,I2507,I49401,I49707,);
not I_2775 (I49393,I49707);
not I_2776 (I49729,I49690);
nand I_2777 (I49378,I49729,I49568);
nor I_2778 (I49760,I260173,I260161);
not I_2779 (I49777,I49760);
nor I_2780 (I49794,I49729,I49777);
nor I_2781 (I49811,I49435,I49794);
DFFARX1 I_2782 (I49811,I2507,I49401,I49387,);
nor I_2783 (I49842,I49495,I49777);
nor I_2784 (I49375,I49690,I49842);
nor I_2785 (I49384,I49625,I49760);
nor I_2786 (I49372,I49495,I49760);
not I_2787 (I49928,I2514);
DFFARX1 I_2788 (I666524,I2507,I49928,I49954,);
not I_2789 (I49962,I49954);
nand I_2790 (I49979,I666527,I666521);
and I_2791 (I49996,I49979,I666518);
DFFARX1 I_2792 (I49996,I2507,I49928,I50022,);
DFFARX1 I_2793 (I666503,I2507,I49928,I50039,);
and I_2794 (I50047,I50039,I666512);
nor I_2795 (I50064,I50022,I50047);
DFFARX1 I_2796 (I50064,I2507,I49928,I49896,);
nand I_2797 (I50095,I50039,I666512);
nand I_2798 (I50112,I49962,I50095);
not I_2799 (I49908,I50112);
DFFARX1 I_2800 (I666503,I2507,I49928,I50152,);
DFFARX1 I_2801 (I50152,I2507,I49928,I49917,);
nand I_2802 (I50174,I666506,I666509);
and I_2803 (I50191,I50174,I666515);
DFFARX1 I_2804 (I50191,I2507,I49928,I50217,);
DFFARX1 I_2805 (I50217,I2507,I49928,I50234,);
not I_2806 (I49920,I50234);
not I_2807 (I50256,I50217);
nand I_2808 (I49905,I50256,I50095);
nor I_2809 (I50287,I666506,I666509);
not I_2810 (I50304,I50287);
nor I_2811 (I50321,I50256,I50304);
nor I_2812 (I50338,I49962,I50321);
DFFARX1 I_2813 (I50338,I2507,I49928,I49914,);
nor I_2814 (I50369,I50022,I50304);
nor I_2815 (I49902,I50217,I50369);
nor I_2816 (I49911,I50152,I50287);
nor I_2817 (I49899,I50022,I50287);
not I_2818 (I50455,I2514);
DFFARX1 I_2819 (I597693,I2507,I50455,I50481,);
not I_2820 (I50489,I50481);
nand I_2821 (I50506,I597708,I597687);
and I_2822 (I50523,I50506,I597690);
DFFARX1 I_2823 (I50523,I2507,I50455,I50549,);
DFFARX1 I_2824 (I597711,I2507,I50455,I50566,);
and I_2825 (I50574,I50566,I597690);
nor I_2826 (I50591,I50549,I50574);
DFFARX1 I_2827 (I50591,I2507,I50455,I50423,);
nand I_2828 (I50622,I50566,I597690);
nand I_2829 (I50639,I50489,I50622);
not I_2830 (I50435,I50639);
DFFARX1 I_2831 (I597687,I2507,I50455,I50679,);
DFFARX1 I_2832 (I50679,I2507,I50455,I50444,);
nand I_2833 (I50701,I597699,I597696);
and I_2834 (I50718,I50701,I597702);
DFFARX1 I_2835 (I50718,I2507,I50455,I50744,);
DFFARX1 I_2836 (I50744,I2507,I50455,I50761,);
not I_2837 (I50447,I50761);
not I_2838 (I50783,I50744);
nand I_2839 (I50432,I50783,I50622);
nor I_2840 (I50814,I597705,I597696);
not I_2841 (I50831,I50814);
nor I_2842 (I50848,I50783,I50831);
nor I_2843 (I50865,I50489,I50848);
DFFARX1 I_2844 (I50865,I2507,I50455,I50441,);
nor I_2845 (I50896,I50549,I50831);
nor I_2846 (I50429,I50744,I50896);
nor I_2847 (I50438,I50679,I50814);
nor I_2848 (I50426,I50549,I50814);
not I_2849 (I50982,I2514);
DFFARX1 I_2850 (I111601,I2507,I50982,I51008,);
not I_2851 (I51016,I51008);
nand I_2852 (I51033,I111595,I111589);
and I_2853 (I51050,I51033,I111610);
DFFARX1 I_2854 (I51050,I2507,I50982,I51076,);
DFFARX1 I_2855 (I111607,I2507,I50982,I51093,);
and I_2856 (I51101,I51093,I111604);
nor I_2857 (I51118,I51076,I51101);
DFFARX1 I_2858 (I51118,I2507,I50982,I50950,);
nand I_2859 (I51149,I51093,I111604);
nand I_2860 (I51166,I51016,I51149);
not I_2861 (I50962,I51166);
DFFARX1 I_2862 (I111589,I2507,I50982,I51206,);
DFFARX1 I_2863 (I51206,I2507,I50982,I50971,);
nand I_2864 (I51228,I111592,I111592);
and I_2865 (I51245,I51228,I111613);
DFFARX1 I_2866 (I51245,I2507,I50982,I51271,);
DFFARX1 I_2867 (I51271,I2507,I50982,I51288,);
not I_2868 (I50974,I51288);
not I_2869 (I51310,I51271);
nand I_2870 (I50959,I51310,I51149);
nor I_2871 (I51341,I111598,I111592);
not I_2872 (I51358,I51341);
nor I_2873 (I51375,I51310,I51358);
nor I_2874 (I51392,I51016,I51375);
DFFARX1 I_2875 (I51392,I2507,I50982,I50968,);
nor I_2876 (I51423,I51076,I51358);
nor I_2877 (I50956,I51271,I51423);
nor I_2878 (I50965,I51206,I51341);
nor I_2879 (I50953,I51076,I51341);
not I_2880 (I51509,I2514);
DFFARX1 I_2881 (I97916,I2507,I51509,I51535,);
not I_2882 (I51543,I51535);
nand I_2883 (I51560,I97910,I97904);
and I_2884 (I51577,I51560,I97925);
DFFARX1 I_2885 (I51577,I2507,I51509,I51603,);
DFFARX1 I_2886 (I97922,I2507,I51509,I51620,);
and I_2887 (I51628,I51620,I97919);
nor I_2888 (I51645,I51603,I51628);
DFFARX1 I_2889 (I51645,I2507,I51509,I51477,);
nand I_2890 (I51676,I51620,I97919);
nand I_2891 (I51693,I51543,I51676);
not I_2892 (I51489,I51693);
DFFARX1 I_2893 (I97904,I2507,I51509,I51733,);
DFFARX1 I_2894 (I51733,I2507,I51509,I51498,);
nand I_2895 (I51755,I97907,I97907);
and I_2896 (I51772,I51755,I97928);
DFFARX1 I_2897 (I51772,I2507,I51509,I51798,);
DFFARX1 I_2898 (I51798,I2507,I51509,I51815,);
not I_2899 (I51501,I51815);
not I_2900 (I51837,I51798);
nand I_2901 (I51486,I51837,I51676);
nor I_2902 (I51868,I97913,I97907);
not I_2903 (I51885,I51868);
nor I_2904 (I51902,I51837,I51885);
nor I_2905 (I51919,I51543,I51902);
DFFARX1 I_2906 (I51919,I2507,I51509,I51495,);
nor I_2907 (I51950,I51603,I51885);
nor I_2908 (I51483,I51798,I51950);
nor I_2909 (I51492,I51733,I51868);
nor I_2910 (I51480,I51603,I51868);
not I_2911 (I52036,I2514);
DFFARX1 I_2912 (I10395,I2507,I52036,I52062,);
not I_2913 (I52070,I52062);
nand I_2914 (I52087,I10383,I10389);
and I_2915 (I52104,I52087,I10392);
DFFARX1 I_2916 (I52104,I2507,I52036,I52130,);
DFFARX1 I_2917 (I10374,I2507,I52036,I52147,);
and I_2918 (I52155,I52147,I10380);
nor I_2919 (I52172,I52130,I52155);
DFFARX1 I_2920 (I52172,I2507,I52036,I52004,);
nand I_2921 (I52203,I52147,I10380);
nand I_2922 (I52220,I52070,I52203);
not I_2923 (I52016,I52220);
DFFARX1 I_2924 (I10374,I2507,I52036,I52260,);
DFFARX1 I_2925 (I52260,I2507,I52036,I52025,);
nand I_2926 (I52282,I10377,I10371);
and I_2927 (I52299,I52282,I10386);
DFFARX1 I_2928 (I52299,I2507,I52036,I52325,);
DFFARX1 I_2929 (I52325,I2507,I52036,I52342,);
not I_2930 (I52028,I52342);
not I_2931 (I52364,I52325);
nand I_2932 (I52013,I52364,I52203);
nor I_2933 (I52395,I10371,I10371);
not I_2934 (I52412,I52395);
nor I_2935 (I52429,I52364,I52412);
nor I_2936 (I52446,I52070,I52429);
DFFARX1 I_2937 (I52446,I2507,I52036,I52022,);
nor I_2938 (I52477,I52130,I52412);
nor I_2939 (I52010,I52325,I52477);
nor I_2940 (I52019,I52260,I52395);
nor I_2941 (I52007,I52130,I52395);
not I_2942 (I52563,I2514);
DFFARX1 I_2943 (I112196,I2507,I52563,I52589,);
not I_2944 (I52597,I52589);
nand I_2945 (I52614,I112190,I112184);
and I_2946 (I52631,I52614,I112205);
DFFARX1 I_2947 (I52631,I2507,I52563,I52657,);
DFFARX1 I_2948 (I112202,I2507,I52563,I52674,);
and I_2949 (I52682,I52674,I112199);
nor I_2950 (I52699,I52657,I52682);
DFFARX1 I_2951 (I52699,I2507,I52563,I52531,);
nand I_2952 (I52730,I52674,I112199);
nand I_2953 (I52747,I52597,I52730);
not I_2954 (I52543,I52747);
DFFARX1 I_2955 (I112184,I2507,I52563,I52787,);
DFFARX1 I_2956 (I52787,I2507,I52563,I52552,);
nand I_2957 (I52809,I112187,I112187);
and I_2958 (I52826,I52809,I112208);
DFFARX1 I_2959 (I52826,I2507,I52563,I52852,);
DFFARX1 I_2960 (I52852,I2507,I52563,I52869,);
not I_2961 (I52555,I52869);
not I_2962 (I52891,I52852);
nand I_2963 (I52540,I52891,I52730);
nor I_2964 (I52922,I112193,I112187);
not I_2965 (I52939,I52922);
nor I_2966 (I52956,I52891,I52939);
nor I_2967 (I52973,I52597,I52956);
DFFARX1 I_2968 (I52973,I2507,I52563,I52549,);
nor I_2969 (I53004,I52657,I52939);
nor I_2970 (I52537,I52852,I53004);
nor I_2971 (I52546,I52787,I52922);
nor I_2972 (I52534,I52657,I52922);
not I_2973 (I53090,I2514);
DFFARX1 I_2974 (I127666,I2507,I53090,I53116,);
not I_2975 (I53124,I53116);
nand I_2976 (I53141,I127660,I127654);
and I_2977 (I53158,I53141,I127675);
DFFARX1 I_2978 (I53158,I2507,I53090,I53184,);
DFFARX1 I_2979 (I127672,I2507,I53090,I53201,);
and I_2980 (I53209,I53201,I127669);
nor I_2981 (I53226,I53184,I53209);
DFFARX1 I_2982 (I53226,I2507,I53090,I53058,);
nand I_2983 (I53257,I53201,I127669);
nand I_2984 (I53274,I53124,I53257);
not I_2985 (I53070,I53274);
DFFARX1 I_2986 (I127654,I2507,I53090,I53314,);
DFFARX1 I_2987 (I53314,I2507,I53090,I53079,);
nand I_2988 (I53336,I127657,I127657);
and I_2989 (I53353,I53336,I127678);
DFFARX1 I_2990 (I53353,I2507,I53090,I53379,);
DFFARX1 I_2991 (I53379,I2507,I53090,I53396,);
not I_2992 (I53082,I53396);
not I_2993 (I53418,I53379);
nand I_2994 (I53067,I53418,I53257);
nor I_2995 (I53449,I127663,I127657);
not I_2996 (I53466,I53449);
nor I_2997 (I53483,I53418,I53466);
nor I_2998 (I53500,I53124,I53483);
DFFARX1 I_2999 (I53500,I2507,I53090,I53076,);
nor I_3000 (I53531,I53184,I53466);
nor I_3001 (I53064,I53379,I53531);
nor I_3002 (I53073,I53314,I53449);
nor I_3003 (I53061,I53184,I53449);
not I_3004 (I53617,I2514);
DFFARX1 I_3005 (I236234,I2507,I53617,I53643,);
not I_3006 (I53651,I53643);
nand I_3007 (I53668,I236228,I236219);
and I_3008 (I53685,I53668,I236240);
DFFARX1 I_3009 (I53685,I2507,I53617,I53711,);
DFFARX1 I_3010 (I236222,I2507,I53617,I53728,);
and I_3011 (I53736,I53728,I236216);
nor I_3012 (I53753,I53711,I53736);
DFFARX1 I_3013 (I53753,I2507,I53617,I53585,);
nand I_3014 (I53784,I53728,I236216);
nand I_3015 (I53801,I53651,I53784);
not I_3016 (I53597,I53801);
DFFARX1 I_3017 (I236216,I2507,I53617,I53841,);
DFFARX1 I_3018 (I53841,I2507,I53617,I53606,);
nand I_3019 (I53863,I236243,I236225);
and I_3020 (I53880,I53863,I236231);
DFFARX1 I_3021 (I53880,I2507,I53617,I53906,);
DFFARX1 I_3022 (I53906,I2507,I53617,I53923,);
not I_3023 (I53609,I53923);
not I_3024 (I53945,I53906);
nand I_3025 (I53594,I53945,I53784);
nor I_3026 (I53976,I236237,I236225);
not I_3027 (I53993,I53976);
nor I_3028 (I54010,I53945,I53993);
nor I_3029 (I54027,I53651,I54010);
DFFARX1 I_3030 (I54027,I2507,I53617,I53603,);
nor I_3031 (I54058,I53711,I53993);
nor I_3032 (I53591,I53906,I54058);
nor I_3033 (I53600,I53841,I53976);
nor I_3034 (I53588,I53711,I53976);
not I_3035 (I54144,I2514);
DFFARX1 I_3036 (I181163,I2507,I54144,I54170,);
not I_3037 (I54178,I54170);
nand I_3038 (I54195,I181145,I181160);
and I_3039 (I54212,I54195,I181136);
DFFARX1 I_3040 (I54212,I2507,I54144,I54238,);
DFFARX1 I_3041 (I181139,I2507,I54144,I54255,);
and I_3042 (I54263,I54255,I181154);
nor I_3043 (I54280,I54238,I54263);
DFFARX1 I_3044 (I54280,I2507,I54144,I54112,);
nand I_3045 (I54311,I54255,I181154);
nand I_3046 (I54328,I54178,I54311);
not I_3047 (I54124,I54328);
DFFARX1 I_3048 (I181157,I2507,I54144,I54368,);
DFFARX1 I_3049 (I54368,I2507,I54144,I54133,);
nand I_3050 (I54390,I181136,I181148);
and I_3051 (I54407,I54390,I181142);
DFFARX1 I_3052 (I54407,I2507,I54144,I54433,);
DFFARX1 I_3053 (I54433,I2507,I54144,I54450,);
not I_3054 (I54136,I54450);
not I_3055 (I54472,I54433);
nand I_3056 (I54121,I54472,I54311);
nor I_3057 (I54503,I181151,I181148);
not I_3058 (I54520,I54503);
nor I_3059 (I54537,I54472,I54520);
nor I_3060 (I54554,I54178,I54537);
DFFARX1 I_3061 (I54554,I2507,I54144,I54130,);
nor I_3062 (I54585,I54238,I54520);
nor I_3063 (I54118,I54433,I54585);
nor I_3064 (I54127,I54368,I54503);
nor I_3065 (I54115,I54238,I54503);
not I_3066 (I54671,I2514);
DFFARX1 I_3067 (I312572,I2507,I54671,I54697,);
not I_3068 (I54705,I54697);
nand I_3069 (I54722,I312584,I312569);
and I_3070 (I54739,I54722,I312563);
DFFARX1 I_3071 (I54739,I2507,I54671,I54765,);
DFFARX1 I_3072 (I312578,I2507,I54671,I54782,);
and I_3073 (I54790,I54782,I312566);
nor I_3074 (I54807,I54765,I54790);
DFFARX1 I_3075 (I54807,I2507,I54671,I54639,);
nand I_3076 (I54838,I54782,I312566);
nand I_3077 (I54855,I54705,I54838);
not I_3078 (I54651,I54855);
DFFARX1 I_3079 (I312575,I2507,I54671,I54895,);
DFFARX1 I_3080 (I54895,I2507,I54671,I54660,);
nand I_3081 (I54917,I312581,I312587);
and I_3082 (I54934,I54917,I312563);
DFFARX1 I_3083 (I54934,I2507,I54671,I54960,);
DFFARX1 I_3084 (I54960,I2507,I54671,I54977,);
not I_3085 (I54663,I54977);
not I_3086 (I54999,I54960);
nand I_3087 (I54648,I54999,I54838);
nor I_3088 (I55030,I312566,I312587);
not I_3089 (I55047,I55030);
nor I_3090 (I55064,I54999,I55047);
nor I_3091 (I55081,I54705,I55064);
DFFARX1 I_3092 (I55081,I2507,I54671,I54657,);
nor I_3093 (I55112,I54765,I55047);
nor I_3094 (I54645,I54960,I55112);
nor I_3095 (I54654,I54895,I55030);
nor I_3096 (I54642,I54765,I55030);
not I_3097 (I55198,I2514);
DFFARX1 I_3098 (I689465,I2507,I55198,I55224,);
not I_3099 (I55232,I55224);
nand I_3100 (I55249,I689459,I689480);
and I_3101 (I55266,I55249,I689456);
DFFARX1 I_3102 (I55266,I2507,I55198,I55292,);
DFFARX1 I_3103 (I689477,I2507,I55198,I55309,);
and I_3104 (I55317,I55309,I689474);
nor I_3105 (I55334,I55292,I55317);
DFFARX1 I_3106 (I55334,I2507,I55198,I55166,);
nand I_3107 (I55365,I55309,I689474);
nand I_3108 (I55382,I55232,I55365);
not I_3109 (I55178,I55382);
DFFARX1 I_3110 (I689462,I2507,I55198,I55422,);
DFFARX1 I_3111 (I55422,I2507,I55198,I55187,);
nand I_3112 (I55444,I689471,I689468);
and I_3113 (I55461,I55444,I689453);
DFFARX1 I_3114 (I55461,I2507,I55198,I55487,);
DFFARX1 I_3115 (I55487,I2507,I55198,I55504,);
not I_3116 (I55190,I55504);
not I_3117 (I55526,I55487);
nand I_3118 (I55175,I55526,I55365);
nor I_3119 (I55557,I689453,I689468);
not I_3120 (I55574,I55557);
nor I_3121 (I55591,I55526,I55574);
nor I_3122 (I55608,I55232,I55591);
DFFARX1 I_3123 (I55608,I2507,I55198,I55184,);
nor I_3124 (I55639,I55292,I55574);
nor I_3125 (I55172,I55487,I55639);
nor I_3126 (I55181,I55422,I55557);
nor I_3127 (I55169,I55292,I55557);
not I_3128 (I55725,I2514);
DFFARX1 I_3129 (I451836,I2507,I55725,I55751,);
not I_3130 (I55759,I55751);
nand I_3131 (I55776,I451833,I451848);
and I_3132 (I55793,I55776,I451830);
DFFARX1 I_3133 (I55793,I2507,I55725,I55819,);
DFFARX1 I_3134 (I451827,I2507,I55725,I55836,);
and I_3135 (I55844,I55836,I451827);
nor I_3136 (I55861,I55819,I55844);
DFFARX1 I_3137 (I55861,I2507,I55725,I55693,);
nand I_3138 (I55892,I55836,I451827);
nand I_3139 (I55909,I55759,I55892);
not I_3140 (I55705,I55909);
DFFARX1 I_3141 (I451830,I2507,I55725,I55949,);
DFFARX1 I_3142 (I55949,I2507,I55725,I55714,);
nand I_3143 (I55971,I451842,I451833);
and I_3144 (I55988,I55971,I451845);
DFFARX1 I_3145 (I55988,I2507,I55725,I56014,);
DFFARX1 I_3146 (I56014,I2507,I55725,I56031,);
not I_3147 (I55717,I56031);
not I_3148 (I56053,I56014);
nand I_3149 (I55702,I56053,I55892);
nor I_3150 (I56084,I451839,I451833);
not I_3151 (I56101,I56084);
nor I_3152 (I56118,I56053,I56101);
nor I_3153 (I56135,I55759,I56118);
DFFARX1 I_3154 (I56135,I2507,I55725,I55711,);
nor I_3155 (I56166,I55819,I56101);
nor I_3156 (I55699,I56014,I56166);
nor I_3157 (I55708,I55949,I56084);
nor I_3158 (I55696,I55819,I56084);
not I_3159 (I56252,I2514);
DFFARX1 I_3160 (I442877,I2507,I56252,I56278,);
not I_3161 (I56286,I56278);
nand I_3162 (I56303,I442874,I442889);
and I_3163 (I56320,I56303,I442871);
DFFARX1 I_3164 (I56320,I2507,I56252,I56346,);
DFFARX1 I_3165 (I442868,I2507,I56252,I56363,);
and I_3166 (I56371,I56363,I442868);
nor I_3167 (I56388,I56346,I56371);
DFFARX1 I_3168 (I56388,I2507,I56252,I56220,);
nand I_3169 (I56419,I56363,I442868);
nand I_3170 (I56436,I56286,I56419);
not I_3171 (I56232,I56436);
DFFARX1 I_3172 (I442871,I2507,I56252,I56476,);
DFFARX1 I_3173 (I56476,I2507,I56252,I56241,);
nand I_3174 (I56498,I442883,I442874);
and I_3175 (I56515,I56498,I442886);
DFFARX1 I_3176 (I56515,I2507,I56252,I56541,);
DFFARX1 I_3177 (I56541,I2507,I56252,I56558,);
not I_3178 (I56244,I56558);
not I_3179 (I56580,I56541);
nand I_3180 (I56229,I56580,I56419);
nor I_3181 (I56611,I442880,I442874);
not I_3182 (I56628,I56611);
nor I_3183 (I56645,I56580,I56628);
nor I_3184 (I56662,I56286,I56645);
DFFARX1 I_3185 (I56662,I2507,I56252,I56238,);
nor I_3186 (I56693,I56346,I56628);
nor I_3187 (I56226,I56541,I56693);
nor I_3188 (I56235,I56476,I56611);
nor I_3189 (I56223,I56346,I56611);
not I_3190 (I56779,I2514);
DFFARX1 I_3191 (I191703,I2507,I56779,I56805,);
not I_3192 (I56813,I56805);
nand I_3193 (I56830,I191685,I191700);
and I_3194 (I56847,I56830,I191676);
DFFARX1 I_3195 (I56847,I2507,I56779,I56873,);
DFFARX1 I_3196 (I191679,I2507,I56779,I56890,);
and I_3197 (I56898,I56890,I191694);
nor I_3198 (I56915,I56873,I56898);
DFFARX1 I_3199 (I56915,I2507,I56779,I56747,);
nand I_3200 (I56946,I56890,I191694);
nand I_3201 (I56963,I56813,I56946);
not I_3202 (I56759,I56963);
DFFARX1 I_3203 (I191697,I2507,I56779,I57003,);
DFFARX1 I_3204 (I57003,I2507,I56779,I56768,);
nand I_3205 (I57025,I191676,I191688);
and I_3206 (I57042,I57025,I191682);
DFFARX1 I_3207 (I57042,I2507,I56779,I57068,);
DFFARX1 I_3208 (I57068,I2507,I56779,I57085,);
not I_3209 (I56771,I57085);
not I_3210 (I57107,I57068);
nand I_3211 (I56756,I57107,I56946);
nor I_3212 (I57138,I191691,I191688);
not I_3213 (I57155,I57138);
nor I_3214 (I57172,I57107,I57155);
nor I_3215 (I57189,I56813,I57172);
DFFARX1 I_3216 (I57189,I2507,I56779,I56765,);
nor I_3217 (I57220,I56873,I57155);
nor I_3218 (I56753,I57068,I57220);
nor I_3219 (I56762,I57003,I57138);
nor I_3220 (I56750,I56873,I57138);
not I_3221 (I57306,I2514);
DFFARX1 I_3222 (I402165,I2507,I57306,I57332,);
not I_3223 (I57340,I57332);
nand I_3224 (I57357,I402156,I402174);
and I_3225 (I57374,I57357,I402153);
DFFARX1 I_3226 (I57374,I2507,I57306,I57400,);
DFFARX1 I_3227 (I402156,I2507,I57306,I57417,);
and I_3228 (I57425,I57417,I402159);
nor I_3229 (I57442,I57400,I57425);
DFFARX1 I_3230 (I57442,I2507,I57306,I57274,);
nand I_3231 (I57473,I57417,I402159);
nand I_3232 (I57490,I57340,I57473);
not I_3233 (I57286,I57490);
DFFARX1 I_3234 (I402153,I2507,I57306,I57530,);
DFFARX1 I_3235 (I57530,I2507,I57306,I57295,);
nand I_3236 (I57552,I402171,I402162);
and I_3237 (I57569,I57552,I402177);
DFFARX1 I_3238 (I57569,I2507,I57306,I57595,);
DFFARX1 I_3239 (I57595,I2507,I57306,I57612,);
not I_3240 (I57298,I57612);
not I_3241 (I57634,I57595);
nand I_3242 (I57283,I57634,I57473);
nor I_3243 (I57665,I402168,I402162);
not I_3244 (I57682,I57665);
nor I_3245 (I57699,I57634,I57682);
nor I_3246 (I57716,I57340,I57699);
DFFARX1 I_3247 (I57716,I2507,I57306,I57292,);
nor I_3248 (I57747,I57400,I57682);
nor I_3249 (I57280,I57595,I57747);
nor I_3250 (I57289,I57530,I57665);
nor I_3251 (I57277,I57400,I57665);
not I_3252 (I57833,I2514);
DFFARX1 I_3253 (I210675,I2507,I57833,I57859,);
not I_3254 (I57867,I57859);
nand I_3255 (I57884,I210657,I210672);
and I_3256 (I57901,I57884,I210648);
DFFARX1 I_3257 (I57901,I2507,I57833,I57927,);
DFFARX1 I_3258 (I210651,I2507,I57833,I57944,);
and I_3259 (I57952,I57944,I210666);
nor I_3260 (I57969,I57927,I57952);
DFFARX1 I_3261 (I57969,I2507,I57833,I57801,);
nand I_3262 (I58000,I57944,I210666);
nand I_3263 (I58017,I57867,I58000);
not I_3264 (I57813,I58017);
DFFARX1 I_3265 (I210669,I2507,I57833,I58057,);
DFFARX1 I_3266 (I58057,I2507,I57833,I57822,);
nand I_3267 (I58079,I210648,I210660);
and I_3268 (I58096,I58079,I210654);
DFFARX1 I_3269 (I58096,I2507,I57833,I58122,);
DFFARX1 I_3270 (I58122,I2507,I57833,I58139,);
not I_3271 (I57825,I58139);
not I_3272 (I58161,I58122);
nand I_3273 (I57810,I58161,I58000);
nor I_3274 (I58192,I210663,I210660);
not I_3275 (I58209,I58192);
nor I_3276 (I58226,I58161,I58209);
nor I_3277 (I58243,I57867,I58226);
DFFARX1 I_3278 (I58243,I2507,I57833,I57819,);
nor I_3279 (I58274,I57927,I58209);
nor I_3280 (I57807,I58122,I58274);
nor I_3281 (I57816,I58057,I58192);
nor I_3282 (I57804,I57927,I58192);
not I_3283 (I58360,I2514);
DFFARX1 I_3284 (I436553,I2507,I58360,I58386,);
not I_3285 (I58394,I58386);
nand I_3286 (I58411,I436550,I436565);
and I_3287 (I58428,I58411,I436547);
DFFARX1 I_3288 (I58428,I2507,I58360,I58454,);
DFFARX1 I_3289 (I436544,I2507,I58360,I58471,);
and I_3290 (I58479,I58471,I436544);
nor I_3291 (I58496,I58454,I58479);
DFFARX1 I_3292 (I58496,I2507,I58360,I58328,);
nand I_3293 (I58527,I58471,I436544);
nand I_3294 (I58544,I58394,I58527);
not I_3295 (I58340,I58544);
DFFARX1 I_3296 (I436547,I2507,I58360,I58584,);
DFFARX1 I_3297 (I58584,I2507,I58360,I58349,);
nand I_3298 (I58606,I436559,I436550);
and I_3299 (I58623,I58606,I436562);
DFFARX1 I_3300 (I58623,I2507,I58360,I58649,);
DFFARX1 I_3301 (I58649,I2507,I58360,I58666,);
not I_3302 (I58352,I58666);
not I_3303 (I58688,I58649);
nand I_3304 (I58337,I58688,I58527);
nor I_3305 (I58719,I436556,I436550);
not I_3306 (I58736,I58719);
nor I_3307 (I58753,I58688,I58736);
nor I_3308 (I58770,I58394,I58753);
DFFARX1 I_3309 (I58770,I2507,I58360,I58346,);
nor I_3310 (I58801,I58454,I58736);
nor I_3311 (I58334,I58649,I58801);
nor I_3312 (I58343,I58584,I58719);
nor I_3313 (I58331,I58454,I58719);
not I_3314 (I58887,I2514);
DFFARX1 I_3315 (I598849,I2507,I58887,I58913,);
not I_3316 (I58921,I58913);
nand I_3317 (I58938,I598864,I598843);
and I_3318 (I58955,I58938,I598846);
DFFARX1 I_3319 (I58955,I2507,I58887,I58981,);
DFFARX1 I_3320 (I598867,I2507,I58887,I58998,);
and I_3321 (I59006,I58998,I598846);
nor I_3322 (I59023,I58981,I59006);
DFFARX1 I_3323 (I59023,I2507,I58887,I58855,);
nand I_3324 (I59054,I58998,I598846);
nand I_3325 (I59071,I58921,I59054);
not I_3326 (I58867,I59071);
DFFARX1 I_3327 (I598843,I2507,I58887,I59111,);
DFFARX1 I_3328 (I59111,I2507,I58887,I58876,);
nand I_3329 (I59133,I598855,I598852);
and I_3330 (I59150,I59133,I598858);
DFFARX1 I_3331 (I59150,I2507,I58887,I59176,);
DFFARX1 I_3332 (I59176,I2507,I58887,I59193,);
not I_3333 (I58879,I59193);
not I_3334 (I59215,I59176);
nand I_3335 (I58864,I59215,I59054);
nor I_3336 (I59246,I598861,I598852);
not I_3337 (I59263,I59246);
nor I_3338 (I59280,I59215,I59263);
nor I_3339 (I59297,I58921,I59280);
DFFARX1 I_3340 (I59297,I2507,I58887,I58873,);
nor I_3341 (I59328,I58981,I59263);
nor I_3342 (I58861,I59176,I59328);
nor I_3343 (I58870,I59111,I59246);
nor I_3344 (I58858,I58981,I59246);
not I_3345 (I59414,I2514);
DFFARX1 I_3346 (I108626,I2507,I59414,I59440,);
not I_3347 (I59448,I59440);
nand I_3348 (I59465,I108620,I108614);
and I_3349 (I59482,I59465,I108635);
DFFARX1 I_3350 (I59482,I2507,I59414,I59508,);
DFFARX1 I_3351 (I108632,I2507,I59414,I59525,);
and I_3352 (I59533,I59525,I108629);
nor I_3353 (I59550,I59508,I59533);
DFFARX1 I_3354 (I59550,I2507,I59414,I59382,);
nand I_3355 (I59581,I59525,I108629);
nand I_3356 (I59598,I59448,I59581);
not I_3357 (I59394,I59598);
DFFARX1 I_3358 (I108614,I2507,I59414,I59638,);
DFFARX1 I_3359 (I59638,I2507,I59414,I59403,);
nand I_3360 (I59660,I108617,I108617);
and I_3361 (I59677,I59660,I108638);
DFFARX1 I_3362 (I59677,I2507,I59414,I59703,);
DFFARX1 I_3363 (I59703,I2507,I59414,I59720,);
not I_3364 (I59406,I59720);
not I_3365 (I59742,I59703);
nand I_3366 (I59391,I59742,I59581);
nor I_3367 (I59773,I108623,I108617);
not I_3368 (I59790,I59773);
nor I_3369 (I59807,I59742,I59790);
nor I_3370 (I59824,I59448,I59807);
DFFARX1 I_3371 (I59824,I2507,I59414,I59400,);
nor I_3372 (I59855,I59508,I59790);
nor I_3373 (I59388,I59703,I59855);
nor I_3374 (I59397,I59638,I59773);
nor I_3375 (I59385,I59508,I59773);
not I_3376 (I59941,I2514);
DFFARX1 I_3377 (I93751,I2507,I59941,I59967,);
not I_3378 (I59975,I59967);
nand I_3379 (I59992,I93745,I93739);
and I_3380 (I60009,I59992,I93760);
DFFARX1 I_3381 (I60009,I2507,I59941,I60035,);
DFFARX1 I_3382 (I93757,I2507,I59941,I60052,);
and I_3383 (I60060,I60052,I93754);
nor I_3384 (I60077,I60035,I60060);
DFFARX1 I_3385 (I60077,I2507,I59941,I59909,);
nand I_3386 (I60108,I60052,I93754);
nand I_3387 (I60125,I59975,I60108);
not I_3388 (I59921,I60125);
DFFARX1 I_3389 (I93739,I2507,I59941,I60165,);
DFFARX1 I_3390 (I60165,I2507,I59941,I59930,);
nand I_3391 (I60187,I93742,I93742);
and I_3392 (I60204,I60187,I93763);
DFFARX1 I_3393 (I60204,I2507,I59941,I60230,);
DFFARX1 I_3394 (I60230,I2507,I59941,I60247,);
not I_3395 (I59933,I60247);
not I_3396 (I60269,I60230);
nand I_3397 (I59918,I60269,I60108);
nor I_3398 (I60300,I93748,I93742);
not I_3399 (I60317,I60300);
nor I_3400 (I60334,I60269,I60317);
nor I_3401 (I60351,I59975,I60334);
DFFARX1 I_3402 (I60351,I2507,I59941,I59927,);
nor I_3403 (I60382,I60035,I60317);
nor I_3404 (I59915,I60230,I60382);
nor I_3405 (I59924,I60165,I60300);
nor I_3406 (I59912,I60035,I60300);
not I_3407 (I60468,I2514);
DFFARX1 I_3408 (I84835,I2507,I60468,I60494,);
not I_3409 (I60502,I60494);
nand I_3410 (I60519,I84832,I84814);
and I_3411 (I60536,I60519,I84820);
DFFARX1 I_3412 (I60536,I2507,I60468,I60562,);
DFFARX1 I_3413 (I84829,I2507,I60468,I60579,);
and I_3414 (I60587,I60579,I84823);
nor I_3415 (I60604,I60562,I60587);
DFFARX1 I_3416 (I60604,I2507,I60468,I60436,);
nand I_3417 (I60635,I60579,I84823);
nand I_3418 (I60652,I60502,I60635);
not I_3419 (I60448,I60652);
DFFARX1 I_3420 (I84838,I2507,I60468,I60692,);
DFFARX1 I_3421 (I60692,I2507,I60468,I60457,);
nand I_3422 (I60714,I84826,I84817);
and I_3423 (I60731,I60714,I84814);
DFFARX1 I_3424 (I60731,I2507,I60468,I60757,);
DFFARX1 I_3425 (I60757,I2507,I60468,I60774,);
not I_3426 (I60460,I60774);
not I_3427 (I60796,I60757);
nand I_3428 (I60445,I60796,I60635);
nor I_3429 (I60827,I84841,I84817);
not I_3430 (I60844,I60827);
nor I_3431 (I60861,I60796,I60844);
nor I_3432 (I60878,I60502,I60861);
DFFARX1 I_3433 (I60878,I2507,I60468,I60454,);
nor I_3434 (I60909,I60562,I60844);
nor I_3435 (I60442,I60757,I60909);
nor I_3436 (I60451,I60692,I60827);
nor I_3437 (I60439,I60562,I60827);
not I_3438 (I60995,I2514);
DFFARX1 I_3439 (I17773,I2507,I60995,I61021,);
not I_3440 (I61029,I61021);
nand I_3441 (I61046,I17761,I17767);
and I_3442 (I61063,I61046,I17770);
DFFARX1 I_3443 (I61063,I2507,I60995,I61089,);
DFFARX1 I_3444 (I17752,I2507,I60995,I61106,);
and I_3445 (I61114,I61106,I17758);
nor I_3446 (I61131,I61089,I61114);
DFFARX1 I_3447 (I61131,I2507,I60995,I60963,);
nand I_3448 (I61162,I61106,I17758);
nand I_3449 (I61179,I61029,I61162);
not I_3450 (I60975,I61179);
DFFARX1 I_3451 (I17752,I2507,I60995,I61219,);
DFFARX1 I_3452 (I61219,I2507,I60995,I60984,);
nand I_3453 (I61241,I17755,I17749);
and I_3454 (I61258,I61241,I17764);
DFFARX1 I_3455 (I61258,I2507,I60995,I61284,);
DFFARX1 I_3456 (I61284,I2507,I60995,I61301,);
not I_3457 (I60987,I61301);
not I_3458 (I61323,I61284);
nand I_3459 (I60972,I61323,I61162);
nor I_3460 (I61354,I17749,I17749);
not I_3461 (I61371,I61354);
nor I_3462 (I61388,I61323,I61371);
nor I_3463 (I61405,I61029,I61388);
DFFARX1 I_3464 (I61405,I2507,I60995,I60981,);
nor I_3465 (I61436,I61089,I61371);
nor I_3466 (I60969,I61284,I61436);
nor I_3467 (I60978,I61219,I61354);
nor I_3468 (I60966,I61089,I61354);
not I_3469 (I61522,I2514);
DFFARX1 I_3470 (I7233,I2507,I61522,I61548,);
not I_3471 (I61556,I61548);
nand I_3472 (I61573,I7221,I7227);
and I_3473 (I61590,I61573,I7230);
DFFARX1 I_3474 (I61590,I2507,I61522,I61616,);
DFFARX1 I_3475 (I7212,I2507,I61522,I61633,);
and I_3476 (I61641,I61633,I7218);
nor I_3477 (I61658,I61616,I61641);
DFFARX1 I_3478 (I61658,I2507,I61522,I61490,);
nand I_3479 (I61689,I61633,I7218);
nand I_3480 (I61706,I61556,I61689);
not I_3481 (I61502,I61706);
DFFARX1 I_3482 (I7212,I2507,I61522,I61746,);
DFFARX1 I_3483 (I61746,I2507,I61522,I61511,);
nand I_3484 (I61768,I7215,I7209);
and I_3485 (I61785,I61768,I7224);
DFFARX1 I_3486 (I61785,I2507,I61522,I61811,);
DFFARX1 I_3487 (I61811,I2507,I61522,I61828,);
not I_3488 (I61514,I61828);
not I_3489 (I61850,I61811);
nand I_3490 (I61499,I61850,I61689);
nor I_3491 (I61881,I7209,I7209);
not I_3492 (I61898,I61881);
nor I_3493 (I61915,I61850,I61898);
nor I_3494 (I61932,I61556,I61915);
DFFARX1 I_3495 (I61932,I2507,I61522,I61508,);
nor I_3496 (I61963,I61616,I61898);
nor I_3497 (I61496,I61811,I61963);
nor I_3498 (I61505,I61746,I61881);
nor I_3499 (I61493,I61616,I61881);
not I_3500 (I62049,I2514);
DFFARX1 I_3501 (I602317,I2507,I62049,I62075,);
not I_3502 (I62083,I62075);
nand I_3503 (I62100,I602332,I602311);
and I_3504 (I62117,I62100,I602314);
DFFARX1 I_3505 (I62117,I2507,I62049,I62143,);
DFFARX1 I_3506 (I602335,I2507,I62049,I62160,);
and I_3507 (I62168,I62160,I602314);
nor I_3508 (I62185,I62143,I62168);
DFFARX1 I_3509 (I62185,I2507,I62049,I62017,);
nand I_3510 (I62216,I62160,I602314);
nand I_3511 (I62233,I62083,I62216);
not I_3512 (I62029,I62233);
DFFARX1 I_3513 (I602311,I2507,I62049,I62273,);
DFFARX1 I_3514 (I62273,I2507,I62049,I62038,);
nand I_3515 (I62295,I602323,I602320);
and I_3516 (I62312,I62295,I602326);
DFFARX1 I_3517 (I62312,I2507,I62049,I62338,);
DFFARX1 I_3518 (I62338,I2507,I62049,I62355,);
not I_3519 (I62041,I62355);
not I_3520 (I62377,I62338);
nand I_3521 (I62026,I62377,I62216);
nor I_3522 (I62408,I602329,I602320);
not I_3523 (I62425,I62408);
nor I_3524 (I62442,I62377,I62425);
nor I_3525 (I62459,I62083,I62442);
DFFARX1 I_3526 (I62459,I2507,I62049,I62035,);
nor I_3527 (I62490,I62143,I62425);
nor I_3528 (I62023,I62338,I62490);
nor I_3529 (I62032,I62273,I62408);
nor I_3530 (I62020,I62143,I62408);
not I_3531 (I62576,I2514);
DFFARX1 I_3532 (I405055,I2507,I62576,I62602,);
not I_3533 (I62610,I62602);
nand I_3534 (I62627,I405046,I405064);
and I_3535 (I62644,I62627,I405043);
DFFARX1 I_3536 (I62644,I2507,I62576,I62670,);
DFFARX1 I_3537 (I405046,I2507,I62576,I62687,);
and I_3538 (I62695,I62687,I405049);
nor I_3539 (I62712,I62670,I62695);
DFFARX1 I_3540 (I62712,I2507,I62576,I62544,);
nand I_3541 (I62743,I62687,I405049);
nand I_3542 (I62760,I62610,I62743);
not I_3543 (I62556,I62760);
DFFARX1 I_3544 (I405043,I2507,I62576,I62800,);
DFFARX1 I_3545 (I62800,I2507,I62576,I62565,);
nand I_3546 (I62822,I405061,I405052);
and I_3547 (I62839,I62822,I405067);
DFFARX1 I_3548 (I62839,I2507,I62576,I62865,);
DFFARX1 I_3549 (I62865,I2507,I62576,I62882,);
not I_3550 (I62568,I62882);
not I_3551 (I62904,I62865);
nand I_3552 (I62553,I62904,I62743);
nor I_3553 (I62935,I405058,I405052);
not I_3554 (I62952,I62935);
nor I_3555 (I62969,I62904,I62952);
nor I_3556 (I62986,I62610,I62969);
DFFARX1 I_3557 (I62986,I2507,I62576,I62562,);
nor I_3558 (I63017,I62670,I62952);
nor I_3559 (I62550,I62865,I63017);
nor I_3560 (I62559,I62800,I62935);
nor I_3561 (I62547,I62670,I62935);
not I_3562 (I63103,I2514);
DFFARX1 I_3563 (I605207,I2507,I63103,I63129,);
not I_3564 (I63137,I63129);
nand I_3565 (I63154,I605222,I605201);
and I_3566 (I63171,I63154,I605204);
DFFARX1 I_3567 (I63171,I2507,I63103,I63197,);
DFFARX1 I_3568 (I605225,I2507,I63103,I63214,);
and I_3569 (I63222,I63214,I605204);
nor I_3570 (I63239,I63197,I63222);
DFFARX1 I_3571 (I63239,I2507,I63103,I63071,);
nand I_3572 (I63270,I63214,I605204);
nand I_3573 (I63287,I63137,I63270);
not I_3574 (I63083,I63287);
DFFARX1 I_3575 (I605201,I2507,I63103,I63327,);
DFFARX1 I_3576 (I63327,I2507,I63103,I63092,);
nand I_3577 (I63349,I605213,I605210);
and I_3578 (I63366,I63349,I605216);
DFFARX1 I_3579 (I63366,I2507,I63103,I63392,);
DFFARX1 I_3580 (I63392,I2507,I63103,I63409,);
not I_3581 (I63095,I63409);
not I_3582 (I63431,I63392);
nand I_3583 (I63080,I63431,I63270);
nor I_3584 (I63462,I605219,I605210);
not I_3585 (I63479,I63462);
nor I_3586 (I63496,I63431,I63479);
nor I_3587 (I63513,I63137,I63496);
DFFARX1 I_3588 (I63513,I2507,I63103,I63089,);
nor I_3589 (I63544,I63197,I63479);
nor I_3590 (I63077,I63392,I63544);
nor I_3591 (I63086,I63327,I63462);
nor I_3592 (I63074,I63197,I63462);
not I_3593 (I63630,I2514);
DFFARX1 I_3594 (I226485,I2507,I63630,I63656,);
not I_3595 (I63664,I63656);
nand I_3596 (I63681,I226467,I226482);
and I_3597 (I63698,I63681,I226458);
DFFARX1 I_3598 (I63698,I2507,I63630,I63724,);
DFFARX1 I_3599 (I226461,I2507,I63630,I63741,);
and I_3600 (I63749,I63741,I226476);
nor I_3601 (I63766,I63724,I63749);
DFFARX1 I_3602 (I63766,I2507,I63630,I63598,);
nand I_3603 (I63797,I63741,I226476);
nand I_3604 (I63814,I63664,I63797);
not I_3605 (I63610,I63814);
DFFARX1 I_3606 (I226479,I2507,I63630,I63854,);
DFFARX1 I_3607 (I63854,I2507,I63630,I63619,);
nand I_3608 (I63876,I226458,I226470);
and I_3609 (I63893,I63876,I226464);
DFFARX1 I_3610 (I63893,I2507,I63630,I63919,);
DFFARX1 I_3611 (I63919,I2507,I63630,I63936,);
not I_3612 (I63622,I63936);
not I_3613 (I63958,I63919);
nand I_3614 (I63607,I63958,I63797);
nor I_3615 (I63989,I226473,I226470);
not I_3616 (I64006,I63989);
nor I_3617 (I64023,I63958,I64006);
nor I_3618 (I64040,I63664,I64023);
DFFARX1 I_3619 (I64040,I2507,I63630,I63616,);
nor I_3620 (I64071,I63724,I64006);
nor I_3621 (I63604,I63919,I64071);
nor I_3622 (I63613,I63854,I63989);
nor I_3623 (I63601,I63724,I63989);
not I_3624 (I64157,I2514);
DFFARX1 I_3625 (I611565,I2507,I64157,I64183,);
not I_3626 (I64191,I64183);
nand I_3627 (I64208,I611580,I611559);
and I_3628 (I64225,I64208,I611562);
DFFARX1 I_3629 (I64225,I2507,I64157,I64251,);
DFFARX1 I_3630 (I611583,I2507,I64157,I64268,);
and I_3631 (I64276,I64268,I611562);
nor I_3632 (I64293,I64251,I64276);
DFFARX1 I_3633 (I64293,I2507,I64157,I64125,);
nand I_3634 (I64324,I64268,I611562);
nand I_3635 (I64341,I64191,I64324);
not I_3636 (I64137,I64341);
DFFARX1 I_3637 (I611559,I2507,I64157,I64381,);
DFFARX1 I_3638 (I64381,I2507,I64157,I64146,);
nand I_3639 (I64403,I611571,I611568);
and I_3640 (I64420,I64403,I611574);
DFFARX1 I_3641 (I64420,I2507,I64157,I64446,);
DFFARX1 I_3642 (I64446,I2507,I64157,I64463,);
not I_3643 (I64149,I64463);
not I_3644 (I64485,I64446);
nand I_3645 (I64134,I64485,I64324);
nor I_3646 (I64516,I611577,I611568);
not I_3647 (I64533,I64516);
nor I_3648 (I64550,I64485,I64533);
nor I_3649 (I64567,I64191,I64550);
DFFARX1 I_3650 (I64567,I2507,I64157,I64143,);
nor I_3651 (I64598,I64251,I64533);
nor I_3652 (I64131,I64446,I64598);
nor I_3653 (I64140,I64381,I64516);
nor I_3654 (I64128,I64251,I64516);
not I_3655 (I64684,I2514);
DFFARX1 I_3656 (I241674,I2507,I64684,I64710,);
not I_3657 (I64718,I64710);
nand I_3658 (I64735,I241668,I241659);
and I_3659 (I64752,I64735,I241680);
DFFARX1 I_3660 (I64752,I2507,I64684,I64778,);
DFFARX1 I_3661 (I241662,I2507,I64684,I64795,);
and I_3662 (I64803,I64795,I241656);
nor I_3663 (I64820,I64778,I64803);
DFFARX1 I_3664 (I64820,I2507,I64684,I64652,);
nand I_3665 (I64851,I64795,I241656);
nand I_3666 (I64868,I64718,I64851);
not I_3667 (I64664,I64868);
DFFARX1 I_3668 (I241656,I2507,I64684,I64908,);
DFFARX1 I_3669 (I64908,I2507,I64684,I64673,);
nand I_3670 (I64930,I241683,I241665);
and I_3671 (I64947,I64930,I241671);
DFFARX1 I_3672 (I64947,I2507,I64684,I64973,);
DFFARX1 I_3673 (I64973,I2507,I64684,I64990,);
not I_3674 (I64676,I64990);
not I_3675 (I65012,I64973);
nand I_3676 (I64661,I65012,I64851);
nor I_3677 (I65043,I241677,I241665);
not I_3678 (I65060,I65043);
nor I_3679 (I65077,I65012,I65060);
nor I_3680 (I65094,I64718,I65077);
DFFARX1 I_3681 (I65094,I2507,I64684,I64670,);
nor I_3682 (I65125,I64778,I65060);
nor I_3683 (I64658,I64973,I65125);
nor I_3684 (I64667,I64908,I65043);
nor I_3685 (I64655,I64778,I65043);
not I_3686 (I65211,I2514);
DFFARX1 I_3687 (I280842,I2507,I65211,I65237,);
not I_3688 (I65245,I65237);
nand I_3689 (I65262,I280836,I280827);
and I_3690 (I65279,I65262,I280848);
DFFARX1 I_3691 (I65279,I2507,I65211,I65305,);
DFFARX1 I_3692 (I280830,I2507,I65211,I65322,);
and I_3693 (I65330,I65322,I280824);
nor I_3694 (I65347,I65305,I65330);
DFFARX1 I_3695 (I65347,I2507,I65211,I65179,);
nand I_3696 (I65378,I65322,I280824);
nand I_3697 (I65395,I65245,I65378);
not I_3698 (I65191,I65395);
DFFARX1 I_3699 (I280824,I2507,I65211,I65435,);
DFFARX1 I_3700 (I65435,I2507,I65211,I65200,);
nand I_3701 (I65457,I280851,I280833);
and I_3702 (I65474,I65457,I280839);
DFFARX1 I_3703 (I65474,I2507,I65211,I65500,);
DFFARX1 I_3704 (I65500,I2507,I65211,I65517,);
not I_3705 (I65203,I65517);
not I_3706 (I65539,I65500);
nand I_3707 (I65188,I65539,I65378);
nor I_3708 (I65570,I280845,I280833);
not I_3709 (I65587,I65570);
nor I_3710 (I65604,I65539,I65587);
nor I_3711 (I65621,I65245,I65604);
DFFARX1 I_3712 (I65621,I2507,I65211,I65197,);
nor I_3713 (I65652,I65305,I65587);
nor I_3714 (I65185,I65500,I65652);
nor I_3715 (I65194,I65435,I65570);
nor I_3716 (I65182,I65305,I65570);
not I_3717 (I65738,I2514);
DFFARX1 I_3718 (I645259,I2507,I65738,I65764,);
not I_3719 (I65772,I65764);
nand I_3720 (I65789,I645253,I645274);
and I_3721 (I65806,I65789,I645265);
DFFARX1 I_3722 (I65806,I2507,I65738,I65832,);
DFFARX1 I_3723 (I645256,I2507,I65738,I65849,);
and I_3724 (I65857,I65849,I645268);
nor I_3725 (I65874,I65832,I65857);
DFFARX1 I_3726 (I65874,I2507,I65738,I65706,);
nand I_3727 (I65905,I65849,I645268);
nand I_3728 (I65922,I65772,I65905);
not I_3729 (I65718,I65922);
DFFARX1 I_3730 (I645256,I2507,I65738,I65962,);
DFFARX1 I_3731 (I65962,I2507,I65738,I65727,);
nand I_3732 (I65984,I645277,I645262);
and I_3733 (I66001,I65984,I645253);
DFFARX1 I_3734 (I66001,I2507,I65738,I66027,);
DFFARX1 I_3735 (I66027,I2507,I65738,I66044,);
not I_3736 (I65730,I66044);
not I_3737 (I66066,I66027);
nand I_3738 (I65715,I66066,I65905);
nor I_3739 (I66097,I645271,I645262);
not I_3740 (I66114,I66097);
nor I_3741 (I66131,I66066,I66114);
nor I_3742 (I66148,I65772,I66131);
DFFARX1 I_3743 (I66148,I2507,I65738,I65724,);
nor I_3744 (I66179,I65832,I66114);
nor I_3745 (I65712,I66027,I66179);
nor I_3746 (I65721,I65962,I66097);
nor I_3747 (I65709,I65832,I66097);
not I_3748 (I66265,I2514);
DFFARX1 I_3749 (I209094,I2507,I66265,I66291,);
not I_3750 (I66299,I66291);
nand I_3751 (I66316,I209076,I209091);
and I_3752 (I66333,I66316,I209067);
DFFARX1 I_3753 (I66333,I2507,I66265,I66359,);
DFFARX1 I_3754 (I209070,I2507,I66265,I66376,);
and I_3755 (I66384,I66376,I209085);
nor I_3756 (I66401,I66359,I66384);
DFFARX1 I_3757 (I66401,I2507,I66265,I66233,);
nand I_3758 (I66432,I66376,I209085);
nand I_3759 (I66449,I66299,I66432);
not I_3760 (I66245,I66449);
DFFARX1 I_3761 (I209088,I2507,I66265,I66489,);
DFFARX1 I_3762 (I66489,I2507,I66265,I66254,);
nand I_3763 (I66511,I209067,I209079);
and I_3764 (I66528,I66511,I209073);
DFFARX1 I_3765 (I66528,I2507,I66265,I66554,);
DFFARX1 I_3766 (I66554,I2507,I66265,I66571,);
not I_3767 (I66257,I66571);
not I_3768 (I66593,I66554);
nand I_3769 (I66242,I66593,I66432);
nor I_3770 (I66624,I209082,I209079);
not I_3771 (I66641,I66624);
nor I_3772 (I66658,I66593,I66641);
nor I_3773 (I66675,I66299,I66658);
DFFARX1 I_3774 (I66675,I2507,I66265,I66251,);
nor I_3775 (I66706,I66359,I66641);
nor I_3776 (I66239,I66554,I66706);
nor I_3777 (I66248,I66489,I66624);
nor I_3778 (I66236,I66359,I66624);
not I_3779 (I66792,I2514);
DFFARX1 I_3780 (I662667,I2507,I66792,I66818,);
not I_3781 (I66826,I66818);
nand I_3782 (I66843,I662661,I662682);
and I_3783 (I66860,I66843,I662673);
DFFARX1 I_3784 (I66860,I2507,I66792,I66886,);
DFFARX1 I_3785 (I662664,I2507,I66792,I66903,);
and I_3786 (I66911,I66903,I662676);
nor I_3787 (I66928,I66886,I66911);
DFFARX1 I_3788 (I66928,I2507,I66792,I66760,);
nand I_3789 (I66959,I66903,I662676);
nand I_3790 (I66976,I66826,I66959);
not I_3791 (I66772,I66976);
DFFARX1 I_3792 (I662664,I2507,I66792,I67016,);
DFFARX1 I_3793 (I67016,I2507,I66792,I66781,);
nand I_3794 (I67038,I662685,I662670);
and I_3795 (I67055,I67038,I662661);
DFFARX1 I_3796 (I67055,I2507,I66792,I67081,);
DFFARX1 I_3797 (I67081,I2507,I66792,I67098,);
not I_3798 (I66784,I67098);
not I_3799 (I67120,I67081);
nand I_3800 (I66769,I67120,I66959);
nor I_3801 (I67151,I662679,I662670);
not I_3802 (I67168,I67151);
nor I_3803 (I67185,I67120,I67168);
nor I_3804 (I67202,I66826,I67185);
DFFARX1 I_3805 (I67202,I2507,I66792,I66778,);
nor I_3806 (I67233,I66886,I67168);
nor I_3807 (I66766,I67081,I67233);
nor I_3808 (I66775,I67016,I67151);
nor I_3809 (I66763,I66886,I67151);
not I_3810 (I67319,I2514);
DFFARX1 I_3811 (I296246,I2507,I67319,I67345,);
not I_3812 (I67353,I67345);
nand I_3813 (I67370,I296267,I296261);
and I_3814 (I67387,I67370,I296243);
DFFARX1 I_3815 (I67387,I2507,I67319,I67413,);
DFFARX1 I_3816 (I296246,I2507,I67319,I67430,);
and I_3817 (I67438,I67430,I296255);
nor I_3818 (I67455,I67413,I67438);
DFFARX1 I_3819 (I67455,I2507,I67319,I67287,);
nand I_3820 (I67486,I67430,I296255);
nand I_3821 (I67503,I67353,I67486);
not I_3822 (I67299,I67503);
DFFARX1 I_3823 (I296252,I2507,I67319,I67543,);
DFFARX1 I_3824 (I67543,I2507,I67319,I67308,);
nand I_3825 (I67565,I296258,I296249);
and I_3826 (I67582,I67565,I296243);
DFFARX1 I_3827 (I67582,I2507,I67319,I67608,);
DFFARX1 I_3828 (I67608,I2507,I67319,I67625,);
not I_3829 (I67311,I67625);
not I_3830 (I67647,I67608);
nand I_3831 (I67296,I67647,I67486);
nor I_3832 (I67678,I296264,I296249);
not I_3833 (I67695,I67678);
nor I_3834 (I67712,I67647,I67695);
nor I_3835 (I67729,I67353,I67712);
DFFARX1 I_3836 (I67729,I2507,I67319,I67305,);
nor I_3837 (I67760,I67413,I67695);
nor I_3838 (I67293,I67608,I67760);
nor I_3839 (I67302,I67543,I67678);
nor I_3840 (I67290,I67413,I67678);
not I_3841 (I67846,I2514);
DFFARX1 I_3842 (I645803,I2507,I67846,I67872,);
not I_3843 (I67880,I67872);
nand I_3844 (I67897,I645797,I645818);
and I_3845 (I67914,I67897,I645809);
DFFARX1 I_3846 (I67914,I2507,I67846,I67940,);
DFFARX1 I_3847 (I645800,I2507,I67846,I67957,);
and I_3848 (I67965,I67957,I645812);
nor I_3849 (I67982,I67940,I67965);
DFFARX1 I_3850 (I67982,I2507,I67846,I67814,);
nand I_3851 (I68013,I67957,I645812);
nand I_3852 (I68030,I67880,I68013);
not I_3853 (I67826,I68030);
DFFARX1 I_3854 (I645800,I2507,I67846,I68070,);
DFFARX1 I_3855 (I68070,I2507,I67846,I67835,);
nand I_3856 (I68092,I645821,I645806);
and I_3857 (I68109,I68092,I645797);
DFFARX1 I_3858 (I68109,I2507,I67846,I68135,);
DFFARX1 I_3859 (I68135,I2507,I67846,I68152,);
not I_3860 (I67838,I68152);
not I_3861 (I68174,I68135);
nand I_3862 (I67823,I68174,I68013);
nor I_3863 (I68205,I645815,I645806);
not I_3864 (I68222,I68205);
nor I_3865 (I68239,I68174,I68222);
nor I_3866 (I68256,I67880,I68239);
DFFARX1 I_3867 (I68256,I2507,I67846,I67832,);
nor I_3868 (I68287,I67940,I68222);
nor I_3869 (I67820,I68135,I68287);
nor I_3870 (I67829,I68070,I68205);
nor I_3871 (I67817,I67940,I68205);
not I_3872 (I68373,I2514);
DFFARX1 I_3873 (I480889,I2507,I68373,I68399,);
not I_3874 (I68407,I68399);
nand I_3875 (I68424,I480907,I480901);
and I_3876 (I68441,I68424,I480880);
DFFARX1 I_3877 (I68441,I2507,I68373,I68467,);
DFFARX1 I_3878 (I480898,I2507,I68373,I68484,);
and I_3879 (I68492,I68484,I480883);
nor I_3880 (I68509,I68467,I68492);
DFFARX1 I_3881 (I68509,I2507,I68373,I68341,);
nand I_3882 (I68540,I68484,I480883);
nand I_3883 (I68557,I68407,I68540);
not I_3884 (I68353,I68557);
DFFARX1 I_3885 (I480895,I2507,I68373,I68597,);
DFFARX1 I_3886 (I68597,I2507,I68373,I68362,);
nand I_3887 (I68619,I480904,I480892);
and I_3888 (I68636,I68619,I480886);
DFFARX1 I_3889 (I68636,I2507,I68373,I68662,);
DFFARX1 I_3890 (I68662,I2507,I68373,I68679,);
not I_3891 (I68365,I68679);
not I_3892 (I68701,I68662);
nand I_3893 (I68350,I68701,I68540);
nor I_3894 (I68732,I480880,I480892);
not I_3895 (I68749,I68732);
nor I_3896 (I68766,I68701,I68749);
nor I_3897 (I68783,I68407,I68766);
DFFARX1 I_3898 (I68783,I2507,I68373,I68359,);
nor I_3899 (I68814,I68467,I68749);
nor I_3900 (I68347,I68662,I68814);
nor I_3901 (I68356,I68597,I68732);
nor I_3902 (I68344,I68467,I68732);
not I_3903 (I68900,I2514);
DFFARX1 I_3904 (I90181,I2507,I68900,I68926,);
not I_3905 (I68934,I68926);
nand I_3906 (I68951,I90175,I90169);
and I_3907 (I68968,I68951,I90190);
DFFARX1 I_3908 (I68968,I2507,I68900,I68994,);
DFFARX1 I_3909 (I90187,I2507,I68900,I69011,);
and I_3910 (I69019,I69011,I90184);
nor I_3911 (I69036,I68994,I69019);
DFFARX1 I_3912 (I69036,I2507,I68900,I68868,);
nand I_3913 (I69067,I69011,I90184);
nand I_3914 (I69084,I68934,I69067);
not I_3915 (I68880,I69084);
DFFARX1 I_3916 (I90169,I2507,I68900,I69124,);
DFFARX1 I_3917 (I69124,I2507,I68900,I68889,);
nand I_3918 (I69146,I90172,I90172);
and I_3919 (I69163,I69146,I90193);
DFFARX1 I_3920 (I69163,I2507,I68900,I69189,);
DFFARX1 I_3921 (I69189,I2507,I68900,I69206,);
not I_3922 (I68892,I69206);
not I_3923 (I69228,I69189);
nand I_3924 (I68877,I69228,I69067);
nor I_3925 (I69259,I90178,I90172);
not I_3926 (I69276,I69259);
nor I_3927 (I69293,I69228,I69276);
nor I_3928 (I69310,I68934,I69293);
DFFARX1 I_3929 (I69310,I2507,I68900,I68886,);
nor I_3930 (I69341,I68994,I69276);
nor I_3931 (I68874,I69189,I69341);
nor I_3932 (I68883,I69124,I69259);
nor I_3933 (I68871,I68994,I69259);
not I_3934 (I69427,I2514);
DFFARX1 I_3935 (I698390,I2507,I69427,I69453,);
not I_3936 (I69461,I69453);
nand I_3937 (I69478,I698384,I698405);
and I_3938 (I69495,I69478,I698381);
DFFARX1 I_3939 (I69495,I2507,I69427,I69521,);
DFFARX1 I_3940 (I698402,I2507,I69427,I69538,);
and I_3941 (I69546,I69538,I698399);
nor I_3942 (I69563,I69521,I69546);
DFFARX1 I_3943 (I69563,I2507,I69427,I69395,);
nand I_3944 (I69594,I69538,I698399);
nand I_3945 (I69611,I69461,I69594);
not I_3946 (I69407,I69611);
DFFARX1 I_3947 (I698387,I2507,I69427,I69651,);
DFFARX1 I_3948 (I69651,I2507,I69427,I69416,);
nand I_3949 (I69673,I698396,I698393);
and I_3950 (I69690,I69673,I698378);
DFFARX1 I_3951 (I69690,I2507,I69427,I69716,);
DFFARX1 I_3952 (I69716,I2507,I69427,I69733,);
not I_3953 (I69419,I69733);
not I_3954 (I69755,I69716);
nand I_3955 (I69404,I69755,I69594);
nor I_3956 (I69786,I698378,I698393);
not I_3957 (I69803,I69786);
nor I_3958 (I69820,I69755,I69803);
nor I_3959 (I69837,I69461,I69820);
DFFARX1 I_3960 (I69837,I2507,I69427,I69413,);
nor I_3961 (I69868,I69521,I69803);
nor I_3962 (I69401,I69716,I69868);
nor I_3963 (I69410,I69651,I69786);
nor I_3964 (I69398,I69521,I69786);
not I_3965 (I69954,I2514);
DFFARX1 I_3966 (I401009,I2507,I69954,I69980,);
not I_3967 (I69988,I69980);
nand I_3968 (I70005,I401000,I401018);
and I_3969 (I70022,I70005,I400997);
DFFARX1 I_3970 (I70022,I2507,I69954,I70048,);
DFFARX1 I_3971 (I401000,I2507,I69954,I70065,);
and I_3972 (I70073,I70065,I401003);
nor I_3973 (I70090,I70048,I70073);
DFFARX1 I_3974 (I70090,I2507,I69954,I69922,);
nand I_3975 (I70121,I70065,I401003);
nand I_3976 (I70138,I69988,I70121);
not I_3977 (I69934,I70138);
DFFARX1 I_3978 (I400997,I2507,I69954,I70178,);
DFFARX1 I_3979 (I70178,I2507,I69954,I69943,);
nand I_3980 (I70200,I401015,I401006);
and I_3981 (I70217,I70200,I401021);
DFFARX1 I_3982 (I70217,I2507,I69954,I70243,);
DFFARX1 I_3983 (I70243,I2507,I69954,I70260,);
not I_3984 (I69946,I70260);
not I_3985 (I70282,I70243);
nand I_3986 (I69931,I70282,I70121);
nor I_3987 (I70313,I401012,I401006);
not I_3988 (I70330,I70313);
nor I_3989 (I70347,I70282,I70330);
nor I_3990 (I70364,I69988,I70347);
DFFARX1 I_3991 (I70364,I2507,I69954,I69940,);
nor I_3992 (I70395,I70048,I70330);
nor I_3993 (I69928,I70243,I70395);
nor I_3994 (I69937,I70178,I70313);
nor I_3995 (I69925,I70048,I70313);
not I_3996 (I70481,I2514);
DFFARX1 I_3997 (I170096,I2507,I70481,I70507,);
not I_3998 (I70515,I70507);
nand I_3999 (I70532,I170078,I170093);
and I_4000 (I70549,I70532,I170069);
DFFARX1 I_4001 (I70549,I2507,I70481,I70575,);
DFFARX1 I_4002 (I170072,I2507,I70481,I70592,);
and I_4003 (I70600,I70592,I170087);
nor I_4004 (I70617,I70575,I70600);
DFFARX1 I_4005 (I70617,I2507,I70481,I70449,);
nand I_4006 (I70648,I70592,I170087);
nand I_4007 (I70665,I70515,I70648);
not I_4008 (I70461,I70665);
DFFARX1 I_4009 (I170090,I2507,I70481,I70705,);
DFFARX1 I_4010 (I70705,I2507,I70481,I70470,);
nand I_4011 (I70727,I170069,I170081);
and I_4012 (I70744,I70727,I170075);
DFFARX1 I_4013 (I70744,I2507,I70481,I70770,);
DFFARX1 I_4014 (I70770,I2507,I70481,I70787,);
not I_4015 (I70473,I70787);
not I_4016 (I70809,I70770);
nand I_4017 (I70458,I70809,I70648);
nor I_4018 (I70840,I170084,I170081);
not I_4019 (I70857,I70840);
nor I_4020 (I70874,I70809,I70857);
nor I_4021 (I70891,I70515,I70874);
DFFARX1 I_4022 (I70891,I2507,I70481,I70467,);
nor I_4023 (I70922,I70575,I70857);
nor I_4024 (I70455,I70770,I70922);
nor I_4025 (I70464,I70705,I70840);
nor I_4026 (I70452,I70575,I70840);
not I_4027 (I71008,I2514);
DFFARX1 I_4028 (I703745,I2507,I71008,I71034,);
not I_4029 (I71042,I71034);
nand I_4030 (I71059,I703739,I703760);
and I_4031 (I71076,I71059,I703736);
DFFARX1 I_4032 (I71076,I2507,I71008,I71102,);
DFFARX1 I_4033 (I703757,I2507,I71008,I71119,);
and I_4034 (I71127,I71119,I703754);
nor I_4035 (I71144,I71102,I71127);
DFFARX1 I_4036 (I71144,I2507,I71008,I70976,);
nand I_4037 (I71175,I71119,I703754);
nand I_4038 (I71192,I71042,I71175);
not I_4039 (I70988,I71192);
DFFARX1 I_4040 (I703742,I2507,I71008,I71232,);
DFFARX1 I_4041 (I71232,I2507,I71008,I70997,);
nand I_4042 (I71254,I703751,I703748);
and I_4043 (I71271,I71254,I703733);
DFFARX1 I_4044 (I71271,I2507,I71008,I71297,);
DFFARX1 I_4045 (I71297,I2507,I71008,I71314,);
not I_4046 (I71000,I71314);
not I_4047 (I71336,I71297);
nand I_4048 (I70985,I71336,I71175);
nor I_4049 (I71367,I703733,I703748);
not I_4050 (I71384,I71367);
nor I_4051 (I71401,I71336,I71384);
nor I_4052 (I71418,I71042,I71401);
DFFARX1 I_4053 (I71418,I2507,I71008,I70994,);
nor I_4054 (I71449,I71102,I71384);
nor I_4055 (I70982,I71297,I71449);
nor I_4056 (I70991,I71232,I71367);
nor I_4057 (I70979,I71102,I71367);
not I_4058 (I71535,I2514);
DFFARX1 I_4059 (I407367,I2507,I71535,I71561,);
not I_4060 (I71569,I71561);
nand I_4061 (I71586,I407358,I407376);
and I_4062 (I71603,I71586,I407355);
DFFARX1 I_4063 (I71603,I2507,I71535,I71629,);
DFFARX1 I_4064 (I407358,I2507,I71535,I71646,);
and I_4065 (I71654,I71646,I407361);
nor I_4066 (I71671,I71629,I71654);
DFFARX1 I_4067 (I71671,I2507,I71535,I71503,);
nand I_4068 (I71702,I71646,I407361);
nand I_4069 (I71719,I71569,I71702);
not I_4070 (I71515,I71719);
DFFARX1 I_4071 (I407355,I2507,I71535,I71759,);
DFFARX1 I_4072 (I71759,I2507,I71535,I71524,);
nand I_4073 (I71781,I407373,I407364);
and I_4074 (I71798,I71781,I407379);
DFFARX1 I_4075 (I71798,I2507,I71535,I71824,);
DFFARX1 I_4076 (I71824,I2507,I71535,I71841,);
not I_4077 (I71527,I71841);
not I_4078 (I71863,I71824);
nand I_4079 (I71512,I71863,I71702);
nor I_4080 (I71894,I407370,I407364);
not I_4081 (I71911,I71894);
nor I_4082 (I71928,I71863,I71911);
nor I_4083 (I71945,I71569,I71928);
DFFARX1 I_4084 (I71945,I2507,I71535,I71521,);
nor I_4085 (I71976,I71629,I71911);
nor I_4086 (I71509,I71824,I71976);
nor I_4087 (I71518,I71759,I71894);
nor I_4088 (I71506,I71629,I71894);
not I_4089 (I72062,I2514);
DFFARX1 I_4090 (I152656,I2507,I72062,I72088,);
not I_4091 (I72096,I72088);
nand I_4092 (I72113,I152650,I152644);
and I_4093 (I72130,I72113,I152665);
DFFARX1 I_4094 (I72130,I2507,I72062,I72156,);
DFFARX1 I_4095 (I152662,I2507,I72062,I72173,);
and I_4096 (I72181,I72173,I152659);
nor I_4097 (I72198,I72156,I72181);
DFFARX1 I_4098 (I72198,I2507,I72062,I72030,);
nand I_4099 (I72229,I72173,I152659);
nand I_4100 (I72246,I72096,I72229);
not I_4101 (I72042,I72246);
DFFARX1 I_4102 (I152644,I2507,I72062,I72286,);
DFFARX1 I_4103 (I72286,I2507,I72062,I72051,);
nand I_4104 (I72308,I152647,I152647);
and I_4105 (I72325,I72308,I152668);
DFFARX1 I_4106 (I72325,I2507,I72062,I72351,);
DFFARX1 I_4107 (I72351,I2507,I72062,I72368,);
not I_4108 (I72054,I72368);
not I_4109 (I72390,I72351);
nand I_4110 (I72039,I72390,I72229);
nor I_4111 (I72421,I152653,I152647);
not I_4112 (I72438,I72421);
nor I_4113 (I72455,I72390,I72438);
nor I_4114 (I72472,I72096,I72455);
DFFARX1 I_4115 (I72472,I2507,I72062,I72048,);
nor I_4116 (I72503,I72156,I72438);
nor I_4117 (I72036,I72351,I72503);
nor I_4118 (I72045,I72286,I72421);
nor I_4119 (I72033,I72156,I72421);
not I_4120 (I72589,I2514);
DFFARX1 I_4121 (I141946,I2507,I72589,I72615,);
not I_4122 (I72623,I72615);
nand I_4123 (I72640,I141940,I141934);
and I_4124 (I72657,I72640,I141955);
DFFARX1 I_4125 (I72657,I2507,I72589,I72683,);
DFFARX1 I_4126 (I141952,I2507,I72589,I72700,);
and I_4127 (I72708,I72700,I141949);
nor I_4128 (I72725,I72683,I72708);
DFFARX1 I_4129 (I72725,I2507,I72589,I72557,);
nand I_4130 (I72756,I72700,I141949);
nand I_4131 (I72773,I72623,I72756);
not I_4132 (I72569,I72773);
DFFARX1 I_4133 (I141934,I2507,I72589,I72813,);
DFFARX1 I_4134 (I72813,I2507,I72589,I72578,);
nand I_4135 (I72835,I141937,I141937);
and I_4136 (I72852,I72835,I141958);
DFFARX1 I_4137 (I72852,I2507,I72589,I72878,);
DFFARX1 I_4138 (I72878,I2507,I72589,I72895,);
not I_4139 (I72581,I72895);
not I_4140 (I72917,I72878);
nand I_4141 (I72566,I72917,I72756);
nor I_4142 (I72948,I141943,I141937);
not I_4143 (I72965,I72948);
nor I_4144 (I72982,I72917,I72965);
nor I_4145 (I72999,I72623,I72982);
DFFARX1 I_4146 (I72999,I2507,I72589,I72575,);
nor I_4147 (I73030,I72683,I72965);
nor I_4148 (I72563,I72878,I73030);
nor I_4149 (I72572,I72813,I72948);
nor I_4150 (I72560,I72683,I72948);
not I_4151 (I73116,I2514);
DFFARX1 I_4152 (I661579,I2507,I73116,I73142,);
not I_4153 (I73150,I73142);
nand I_4154 (I73167,I661573,I661594);
and I_4155 (I73184,I73167,I661585);
DFFARX1 I_4156 (I73184,I2507,I73116,I73210,);
DFFARX1 I_4157 (I661576,I2507,I73116,I73227,);
and I_4158 (I73235,I73227,I661588);
nor I_4159 (I73252,I73210,I73235);
DFFARX1 I_4160 (I73252,I2507,I73116,I73084,);
nand I_4161 (I73283,I73227,I661588);
nand I_4162 (I73300,I73150,I73283);
not I_4163 (I73096,I73300);
DFFARX1 I_4164 (I661576,I2507,I73116,I73340,);
DFFARX1 I_4165 (I73340,I2507,I73116,I73105,);
nand I_4166 (I73362,I661597,I661582);
and I_4167 (I73379,I73362,I661573);
DFFARX1 I_4168 (I73379,I2507,I73116,I73405,);
DFFARX1 I_4169 (I73405,I2507,I73116,I73422,);
not I_4170 (I73108,I73422);
not I_4171 (I73444,I73405);
nand I_4172 (I73093,I73444,I73283);
nor I_4173 (I73475,I661591,I661582);
not I_4174 (I73492,I73475);
nor I_4175 (I73509,I73444,I73492);
nor I_4176 (I73526,I73150,I73509);
DFFARX1 I_4177 (I73526,I2507,I73116,I73102,);
nor I_4178 (I73557,I73210,I73492);
nor I_4179 (I73090,I73405,I73557);
nor I_4180 (I73099,I73340,I73475);
nor I_4181 (I73087,I73210,I73475);
not I_4182 (I73643,I2514);
DFFARX1 I_4183 (I1444,I2507,I73643,I73669,);
not I_4184 (I73677,I73669);
nand I_4185 (I73694,I1572,I1492);
and I_4186 (I73711,I73694,I1476);
DFFARX1 I_4187 (I73711,I2507,I73643,I73737,);
DFFARX1 I_4188 (I2116,I2507,I73643,I73754,);
and I_4189 (I73762,I73754,I1820);
nor I_4190 (I73779,I73737,I73762);
DFFARX1 I_4191 (I73779,I2507,I73643,I73611,);
nand I_4192 (I73810,I73754,I1820);
nand I_4193 (I73827,I73677,I73810);
not I_4194 (I73623,I73827);
DFFARX1 I_4195 (I1940,I2507,I73643,I73867,);
DFFARX1 I_4196 (I73867,I2507,I73643,I73632,);
nand I_4197 (I73889,I2324,I1428);
and I_4198 (I73906,I73889,I1924);
DFFARX1 I_4199 (I73906,I2507,I73643,I73932,);
DFFARX1 I_4200 (I73932,I2507,I73643,I73949,);
not I_4201 (I73635,I73949);
not I_4202 (I73971,I73932);
nand I_4203 (I73620,I73971,I73810);
nor I_4204 (I74002,I1780,I1428);
not I_4205 (I74019,I74002);
nor I_4206 (I74036,I73971,I74019);
nor I_4207 (I74053,I73677,I74036);
DFFARX1 I_4208 (I74053,I2507,I73643,I73629,);
nor I_4209 (I74084,I73737,I74019);
nor I_4210 (I73617,I73932,I74084);
nor I_4211 (I73626,I73867,I74002);
nor I_4212 (I73614,I73737,I74002);
not I_4213 (I74170,I2514);
DFFARX1 I_4214 (I358237,I2507,I74170,I74196,);
not I_4215 (I74204,I74196);
nand I_4216 (I74221,I358228,I358246);
and I_4217 (I74238,I74221,I358225);
DFFARX1 I_4218 (I74238,I2507,I74170,I74264,);
DFFARX1 I_4219 (I358228,I2507,I74170,I74281,);
and I_4220 (I74289,I74281,I358231);
nor I_4221 (I74306,I74264,I74289);
DFFARX1 I_4222 (I74306,I2507,I74170,I74138,);
nand I_4223 (I74337,I74281,I358231);
nand I_4224 (I74354,I74204,I74337);
not I_4225 (I74150,I74354);
DFFARX1 I_4226 (I358225,I2507,I74170,I74394,);
DFFARX1 I_4227 (I74394,I2507,I74170,I74159,);
nand I_4228 (I74416,I358243,I358234);
and I_4229 (I74433,I74416,I358249);
DFFARX1 I_4230 (I74433,I2507,I74170,I74459,);
DFFARX1 I_4231 (I74459,I2507,I74170,I74476,);
not I_4232 (I74162,I74476);
not I_4233 (I74498,I74459);
nand I_4234 (I74147,I74498,I74337);
nor I_4235 (I74529,I358240,I358234);
not I_4236 (I74546,I74529);
nor I_4237 (I74563,I74498,I74546);
nor I_4238 (I74580,I74204,I74563);
DFFARX1 I_4239 (I74580,I2507,I74170,I74156,);
nor I_4240 (I74611,I74264,I74546);
nor I_4241 (I74144,I74459,I74611);
nor I_4242 (I74153,I74394,I74529);
nor I_4243 (I74141,I74264,I74529);
not I_4244 (I74697,I2514);
DFFARX1 I_4245 (I493163,I2507,I74697,I74723,);
not I_4246 (I74731,I74723);
nand I_4247 (I74748,I493181,I493175);
and I_4248 (I74765,I74748,I493154);
DFFARX1 I_4249 (I74765,I2507,I74697,I74791,);
DFFARX1 I_4250 (I493172,I2507,I74697,I74808,);
and I_4251 (I74816,I74808,I493157);
nor I_4252 (I74833,I74791,I74816);
DFFARX1 I_4253 (I74833,I2507,I74697,I74665,);
nand I_4254 (I74864,I74808,I493157);
nand I_4255 (I74881,I74731,I74864);
not I_4256 (I74677,I74881);
DFFARX1 I_4257 (I493169,I2507,I74697,I74921,);
DFFARX1 I_4258 (I74921,I2507,I74697,I74686,);
nand I_4259 (I74943,I493178,I493166);
and I_4260 (I74960,I74943,I493160);
DFFARX1 I_4261 (I74960,I2507,I74697,I74986,);
DFFARX1 I_4262 (I74986,I2507,I74697,I75003,);
not I_4263 (I74689,I75003);
not I_4264 (I75025,I74986);
nand I_4265 (I74674,I75025,I74864);
nor I_4266 (I75056,I493154,I493166);
not I_4267 (I75073,I75056);
nor I_4268 (I75090,I75025,I75073);
nor I_4269 (I75107,I74731,I75090);
DFFARX1 I_4270 (I75107,I2507,I74697,I74683,);
nor I_4271 (I75138,I74791,I75073);
nor I_4272 (I74671,I74986,I75138);
nor I_4273 (I74680,I74921,I75056);
nor I_4274 (I74668,I74791,I75056);
not I_4275 (I75224,I2514);
DFFARX1 I_4276 (I265066,I2507,I75224,I75250,);
not I_4277 (I75258,I75250);
nand I_4278 (I75275,I265060,I265051);
and I_4279 (I75292,I75275,I265072);
DFFARX1 I_4280 (I75292,I2507,I75224,I75318,);
DFFARX1 I_4281 (I265054,I2507,I75224,I75335,);
and I_4282 (I75343,I75335,I265048);
nor I_4283 (I75360,I75318,I75343);
DFFARX1 I_4284 (I75360,I2507,I75224,I75192,);
nand I_4285 (I75391,I75335,I265048);
nand I_4286 (I75408,I75258,I75391);
not I_4287 (I75204,I75408);
DFFARX1 I_4288 (I265048,I2507,I75224,I75448,);
DFFARX1 I_4289 (I75448,I2507,I75224,I75213,);
nand I_4290 (I75470,I265075,I265057);
and I_4291 (I75487,I75470,I265063);
DFFARX1 I_4292 (I75487,I2507,I75224,I75513,);
DFFARX1 I_4293 (I75513,I2507,I75224,I75530,);
not I_4294 (I75216,I75530);
not I_4295 (I75552,I75513);
nand I_4296 (I75201,I75552,I75391);
nor I_4297 (I75583,I265069,I265057);
not I_4298 (I75600,I75583);
nor I_4299 (I75617,I75552,I75600);
nor I_4300 (I75634,I75258,I75617);
DFFARX1 I_4301 (I75634,I2507,I75224,I75210,);
nor I_4302 (I75665,I75318,I75600);
nor I_4303 (I75198,I75513,I75665);
nor I_4304 (I75207,I75448,I75583);
nor I_4305 (I75195,I75318,I75583);
not I_4306 (I75751,I2514);
DFFARX1 I_4307 (I386559,I2507,I75751,I75777,);
not I_4308 (I75785,I75777);
nand I_4309 (I75802,I386550,I386568);
and I_4310 (I75819,I75802,I386547);
DFFARX1 I_4311 (I75819,I2507,I75751,I75845,);
DFFARX1 I_4312 (I386550,I2507,I75751,I75862,);
and I_4313 (I75870,I75862,I386553);
nor I_4314 (I75887,I75845,I75870);
DFFARX1 I_4315 (I75887,I2507,I75751,I75719,);
nand I_4316 (I75918,I75862,I386553);
nand I_4317 (I75935,I75785,I75918);
not I_4318 (I75731,I75935);
DFFARX1 I_4319 (I386547,I2507,I75751,I75975,);
DFFARX1 I_4320 (I75975,I2507,I75751,I75740,);
nand I_4321 (I75997,I386565,I386556);
and I_4322 (I76014,I75997,I386571);
DFFARX1 I_4323 (I76014,I2507,I75751,I76040,);
DFFARX1 I_4324 (I76040,I2507,I75751,I76057,);
not I_4325 (I75743,I76057);
not I_4326 (I76079,I76040);
nand I_4327 (I75728,I76079,I75918);
nor I_4328 (I76110,I386562,I386556);
not I_4329 (I76127,I76110);
nor I_4330 (I76144,I76079,I76127);
nor I_4331 (I76161,I75785,I76144);
DFFARX1 I_4332 (I76161,I2507,I75751,I75737,);
nor I_4333 (I76192,I75845,I76127);
nor I_4334 (I75725,I76040,I76192);
nor I_4335 (I75734,I75975,I76110);
nor I_4336 (I75722,I75845,I76110);
not I_4337 (I76278,I2514);
DFFARX1 I_4338 (I701365,I2507,I76278,I76304,);
not I_4339 (I76312,I76304);
nand I_4340 (I76329,I701359,I701380);
and I_4341 (I76346,I76329,I701356);
DFFARX1 I_4342 (I76346,I2507,I76278,I76372,);
DFFARX1 I_4343 (I701377,I2507,I76278,I76389,);
and I_4344 (I76397,I76389,I701374);
nor I_4345 (I76414,I76372,I76397);
DFFARX1 I_4346 (I76414,I2507,I76278,I76246,);
nand I_4347 (I76445,I76389,I701374);
nand I_4348 (I76462,I76312,I76445);
not I_4349 (I76258,I76462);
DFFARX1 I_4350 (I701362,I2507,I76278,I76502,);
DFFARX1 I_4351 (I76502,I2507,I76278,I76267,);
nand I_4352 (I76524,I701371,I701368);
and I_4353 (I76541,I76524,I701353);
DFFARX1 I_4354 (I76541,I2507,I76278,I76567,);
DFFARX1 I_4355 (I76567,I2507,I76278,I76584,);
not I_4356 (I76270,I76584);
not I_4357 (I76606,I76567);
nand I_4358 (I76255,I76606,I76445);
nor I_4359 (I76637,I701353,I701368);
not I_4360 (I76654,I76637);
nor I_4361 (I76671,I76606,I76654);
nor I_4362 (I76688,I76312,I76671);
DFFARX1 I_4363 (I76688,I2507,I76278,I76264,);
nor I_4364 (I76719,I76372,I76654);
nor I_4365 (I76252,I76567,I76719);
nor I_4366 (I76261,I76502,I76637);
nor I_4367 (I76249,I76372,I76637);
not I_4368 (I76805,I2514);
DFFARX1 I_4369 (I125881,I2507,I76805,I76831,);
not I_4370 (I76839,I76831);
nand I_4371 (I76856,I125875,I125869);
and I_4372 (I76873,I76856,I125890);
DFFARX1 I_4373 (I76873,I2507,I76805,I76899,);
DFFARX1 I_4374 (I125887,I2507,I76805,I76916,);
and I_4375 (I76924,I76916,I125884);
nor I_4376 (I76941,I76899,I76924);
DFFARX1 I_4377 (I76941,I2507,I76805,I76773,);
nand I_4378 (I76972,I76916,I125884);
nand I_4379 (I76989,I76839,I76972);
not I_4380 (I76785,I76989);
DFFARX1 I_4381 (I125869,I2507,I76805,I77029,);
DFFARX1 I_4382 (I77029,I2507,I76805,I76794,);
nand I_4383 (I77051,I125872,I125872);
and I_4384 (I77068,I77051,I125893);
DFFARX1 I_4385 (I77068,I2507,I76805,I77094,);
DFFARX1 I_4386 (I77094,I2507,I76805,I77111,);
not I_4387 (I76797,I77111);
not I_4388 (I77133,I77094);
nand I_4389 (I76782,I77133,I76972);
nor I_4390 (I77164,I125878,I125872);
not I_4391 (I77181,I77164);
nor I_4392 (I77198,I77133,I77181);
nor I_4393 (I77215,I76839,I77198);
DFFARX1 I_4394 (I77215,I2507,I76805,I76791,);
nor I_4395 (I77246,I76899,I77181);
nor I_4396 (I76779,I77094,I77246);
nor I_4397 (I76788,I77029,I77164);
nor I_4398 (I76776,I76899,I77164);
not I_4399 (I77332,I2514);
DFFARX1 I_4400 (I388871,I2507,I77332,I77358,);
not I_4401 (I77366,I77358);
nand I_4402 (I77383,I388862,I388880);
and I_4403 (I77400,I77383,I388859);
DFFARX1 I_4404 (I77400,I2507,I77332,I77426,);
DFFARX1 I_4405 (I388862,I2507,I77332,I77443,);
and I_4406 (I77451,I77443,I388865);
nor I_4407 (I77468,I77426,I77451);
DFFARX1 I_4408 (I77468,I2507,I77332,I77300,);
nand I_4409 (I77499,I77443,I388865);
nand I_4410 (I77516,I77366,I77499);
not I_4411 (I77312,I77516);
DFFARX1 I_4412 (I388859,I2507,I77332,I77556,);
DFFARX1 I_4413 (I77556,I2507,I77332,I77321,);
nand I_4414 (I77578,I388877,I388868);
and I_4415 (I77595,I77578,I388883);
DFFARX1 I_4416 (I77595,I2507,I77332,I77621,);
DFFARX1 I_4417 (I77621,I2507,I77332,I77638,);
not I_4418 (I77324,I77638);
not I_4419 (I77660,I77621);
nand I_4420 (I77309,I77660,I77499);
nor I_4421 (I77691,I388874,I388868);
not I_4422 (I77708,I77691);
nor I_4423 (I77725,I77660,I77708);
nor I_4424 (I77742,I77366,I77725);
DFFARX1 I_4425 (I77742,I2507,I77332,I77318,);
nor I_4426 (I77773,I77426,I77708);
nor I_4427 (I77306,I77621,I77773);
nor I_4428 (I77315,I77556,I77691);
nor I_4429 (I77303,I77426,I77691);
not I_4430 (I77859,I2514);
DFFARX1 I_4431 (I172204,I2507,I77859,I77885,);
not I_4432 (I77893,I77885);
nand I_4433 (I77910,I172186,I172201);
and I_4434 (I77927,I77910,I172177);
DFFARX1 I_4435 (I77927,I2507,I77859,I77953,);
DFFARX1 I_4436 (I172180,I2507,I77859,I77970,);
and I_4437 (I77978,I77970,I172195);
nor I_4438 (I77995,I77953,I77978);
DFFARX1 I_4439 (I77995,I2507,I77859,I77827,);
nand I_4440 (I78026,I77970,I172195);
nand I_4441 (I78043,I77893,I78026);
not I_4442 (I77839,I78043);
DFFARX1 I_4443 (I172198,I2507,I77859,I78083,);
DFFARX1 I_4444 (I78083,I2507,I77859,I77848,);
nand I_4445 (I78105,I172177,I172189);
and I_4446 (I78122,I78105,I172183);
DFFARX1 I_4447 (I78122,I2507,I77859,I78148,);
DFFARX1 I_4448 (I78148,I2507,I77859,I78165,);
not I_4449 (I77851,I78165);
not I_4450 (I78187,I78148);
nand I_4451 (I77836,I78187,I78026);
nor I_4452 (I78218,I172192,I172189);
not I_4453 (I78235,I78218);
nor I_4454 (I78252,I78187,I78235);
nor I_4455 (I78269,I77893,I78252);
DFFARX1 I_4456 (I78269,I2507,I77859,I77845,);
nor I_4457 (I78300,I77953,I78235);
nor I_4458 (I77833,I78148,I78300);
nor I_4459 (I77842,I78083,I78218);
nor I_4460 (I77830,I77953,I78218);
not I_4461 (I78386,I2514);
DFFARX1 I_4462 (I216999,I2507,I78386,I78412,);
not I_4463 (I78420,I78412);
nand I_4464 (I78437,I216981,I216996);
and I_4465 (I78454,I78437,I216972);
DFFARX1 I_4466 (I78454,I2507,I78386,I78480,);
DFFARX1 I_4467 (I216975,I2507,I78386,I78497,);
and I_4468 (I78505,I78497,I216990);
nor I_4469 (I78522,I78480,I78505);
DFFARX1 I_4470 (I78522,I2507,I78386,I78354,);
nand I_4471 (I78553,I78497,I216990);
nand I_4472 (I78570,I78420,I78553);
not I_4473 (I78366,I78570);
DFFARX1 I_4474 (I216993,I2507,I78386,I78610,);
DFFARX1 I_4475 (I78610,I2507,I78386,I78375,);
nand I_4476 (I78632,I216972,I216984);
and I_4477 (I78649,I78632,I216978);
DFFARX1 I_4478 (I78649,I2507,I78386,I78675,);
DFFARX1 I_4479 (I78675,I2507,I78386,I78692,);
not I_4480 (I78378,I78692);
not I_4481 (I78714,I78675);
nand I_4482 (I78363,I78714,I78553);
nor I_4483 (I78745,I216987,I216984);
not I_4484 (I78762,I78745);
nor I_4485 (I78779,I78714,I78762);
nor I_4486 (I78796,I78420,I78779);
DFFARX1 I_4487 (I78796,I2507,I78386,I78372,);
nor I_4488 (I78827,I78480,I78762);
nor I_4489 (I78360,I78675,I78827);
nor I_4490 (I78369,I78610,I78745);
nor I_4491 (I78357,I78480,I78745);
not I_4492 (I78913,I2514);
DFFARX1 I_4493 (I661035,I2507,I78913,I78939,);
not I_4494 (I78947,I78939);
nand I_4495 (I78964,I661029,I661050);
and I_4496 (I78981,I78964,I661041);
DFFARX1 I_4497 (I78981,I2507,I78913,I79007,);
DFFARX1 I_4498 (I661032,I2507,I78913,I79024,);
and I_4499 (I79032,I79024,I661044);
nor I_4500 (I79049,I79007,I79032);
DFFARX1 I_4501 (I79049,I2507,I78913,I78881,);
nand I_4502 (I79080,I79024,I661044);
nand I_4503 (I79097,I78947,I79080);
not I_4504 (I78893,I79097);
DFFARX1 I_4505 (I661032,I2507,I78913,I79137,);
DFFARX1 I_4506 (I79137,I2507,I78913,I78902,);
nand I_4507 (I79159,I661053,I661038);
and I_4508 (I79176,I79159,I661029);
DFFARX1 I_4509 (I79176,I2507,I78913,I79202,);
DFFARX1 I_4510 (I79202,I2507,I78913,I79219,);
not I_4511 (I78905,I79219);
not I_4512 (I79241,I79202);
nand I_4513 (I78890,I79241,I79080);
nor I_4514 (I79272,I661047,I661038);
not I_4515 (I79289,I79272);
nor I_4516 (I79306,I79241,I79289);
nor I_4517 (I79323,I78947,I79306);
DFFARX1 I_4518 (I79323,I2507,I78913,I78899,);
nor I_4519 (I79354,I79007,I79289);
nor I_4520 (I78887,I79202,I79354);
nor I_4521 (I78896,I79137,I79272);
nor I_4522 (I78884,I79007,I79272);
not I_4523 (I79440,I2514);
DFFARX1 I_4524 (I616767,I2507,I79440,I79466,);
not I_4525 (I79474,I79466);
nand I_4526 (I79491,I616782,I616761);
and I_4527 (I79508,I79491,I616764);
DFFARX1 I_4528 (I79508,I2507,I79440,I79534,);
DFFARX1 I_4529 (I616785,I2507,I79440,I79551,);
and I_4530 (I79559,I79551,I616764);
nor I_4531 (I79576,I79534,I79559);
DFFARX1 I_4532 (I79576,I2507,I79440,I79408,);
nand I_4533 (I79607,I79551,I616764);
nand I_4534 (I79624,I79474,I79607);
not I_4535 (I79420,I79624);
DFFARX1 I_4536 (I616761,I2507,I79440,I79664,);
DFFARX1 I_4537 (I79664,I2507,I79440,I79429,);
nand I_4538 (I79686,I616773,I616770);
and I_4539 (I79703,I79686,I616776);
DFFARX1 I_4540 (I79703,I2507,I79440,I79729,);
DFFARX1 I_4541 (I79729,I2507,I79440,I79746,);
not I_4542 (I79432,I79746);
not I_4543 (I79768,I79729);
nand I_4544 (I79417,I79768,I79607);
nor I_4545 (I79799,I616779,I616770);
not I_4546 (I79816,I79799);
nor I_4547 (I79833,I79768,I79816);
nor I_4548 (I79850,I79474,I79833);
DFFARX1 I_4549 (I79850,I2507,I79440,I79426,);
nor I_4550 (I79881,I79534,I79816);
nor I_4551 (I79414,I79729,I79881);
nor I_4552 (I79423,I79664,I79799);
nor I_4553 (I79411,I79534,I79799);
not I_4554 (I79967,I2514);
DFFARX1 I_4555 (I9341,I2507,I79967,I79993,);
not I_4556 (I80001,I79993);
nand I_4557 (I80018,I9329,I9335);
and I_4558 (I80035,I80018,I9338);
DFFARX1 I_4559 (I80035,I2507,I79967,I80061,);
DFFARX1 I_4560 (I9320,I2507,I79967,I80078,);
and I_4561 (I80086,I80078,I9326);
nor I_4562 (I80103,I80061,I80086);
DFFARX1 I_4563 (I80103,I2507,I79967,I79935,);
nand I_4564 (I80134,I80078,I9326);
nand I_4565 (I80151,I80001,I80134);
not I_4566 (I79947,I80151);
DFFARX1 I_4567 (I9320,I2507,I79967,I80191,);
DFFARX1 I_4568 (I80191,I2507,I79967,I79956,);
nand I_4569 (I80213,I9323,I9317);
and I_4570 (I80230,I80213,I9332);
DFFARX1 I_4571 (I80230,I2507,I79967,I80256,);
DFFARX1 I_4572 (I80256,I2507,I79967,I80273,);
not I_4573 (I79959,I80273);
not I_4574 (I80295,I80256);
nand I_4575 (I79944,I80295,I80134);
nor I_4576 (I80326,I9317,I9317);
not I_4577 (I80343,I80326);
nor I_4578 (I80360,I80295,I80343);
nor I_4579 (I80377,I80001,I80360);
DFFARX1 I_4580 (I80377,I2507,I79967,I79953,);
nor I_4581 (I80408,I80061,I80343);
nor I_4582 (I79941,I80256,I80408);
nor I_4583 (I79950,I80191,I80326);
nor I_4584 (I79938,I80061,I80326);
not I_4585 (I80494,I2514);
DFFARX1 I_4586 (I582665,I2507,I80494,I80520,);
not I_4587 (I80528,I80520);
nand I_4588 (I80545,I582680,I582659);
and I_4589 (I80562,I80545,I582662);
DFFARX1 I_4590 (I80562,I2507,I80494,I80588,);
DFFARX1 I_4591 (I582683,I2507,I80494,I80605,);
and I_4592 (I80613,I80605,I582662);
nor I_4593 (I80630,I80588,I80613);
DFFARX1 I_4594 (I80630,I2507,I80494,I80462,);
nand I_4595 (I80661,I80605,I582662);
nand I_4596 (I80678,I80528,I80661);
not I_4597 (I80474,I80678);
DFFARX1 I_4598 (I582659,I2507,I80494,I80718,);
DFFARX1 I_4599 (I80718,I2507,I80494,I80483,);
nand I_4600 (I80740,I582671,I582668);
and I_4601 (I80757,I80740,I582674);
DFFARX1 I_4602 (I80757,I2507,I80494,I80783,);
DFFARX1 I_4603 (I80783,I2507,I80494,I80800,);
not I_4604 (I80486,I80800);
not I_4605 (I80822,I80783);
nand I_4606 (I80471,I80822,I80661);
nor I_4607 (I80853,I582677,I582668);
not I_4608 (I80870,I80853);
nor I_4609 (I80887,I80822,I80870);
nor I_4610 (I80904,I80528,I80887);
DFFARX1 I_4611 (I80904,I2507,I80494,I80480,);
nor I_4612 (I80935,I80588,I80870);
nor I_4613 (I80468,I80783,I80935);
nor I_4614 (I80477,I80718,I80853);
nor I_4615 (I80465,I80588,I80853);
not I_4616 (I81021,I2514);
DFFARX1 I_4617 (I183271,I2507,I81021,I81047,);
not I_4618 (I81055,I81047);
nand I_4619 (I81072,I183253,I183268);
and I_4620 (I81089,I81072,I183244);
DFFARX1 I_4621 (I81089,I2507,I81021,I81115,);
DFFARX1 I_4622 (I183247,I2507,I81021,I81132,);
and I_4623 (I81140,I81132,I183262);
nor I_4624 (I81157,I81115,I81140);
DFFARX1 I_4625 (I81157,I2507,I81021,I80989,);
nand I_4626 (I81188,I81132,I183262);
nand I_4627 (I81205,I81055,I81188);
not I_4628 (I81001,I81205);
DFFARX1 I_4629 (I183265,I2507,I81021,I81245,);
DFFARX1 I_4630 (I81245,I2507,I81021,I81010,);
nand I_4631 (I81267,I183244,I183256);
and I_4632 (I81284,I81267,I183250);
DFFARX1 I_4633 (I81284,I2507,I81021,I81310,);
DFFARX1 I_4634 (I81310,I2507,I81021,I81327,);
not I_4635 (I81013,I81327);
not I_4636 (I81349,I81310);
nand I_4637 (I80998,I81349,I81188);
nor I_4638 (I81380,I183259,I183256);
not I_4639 (I81397,I81380);
nor I_4640 (I81414,I81349,I81397);
nor I_4641 (I81431,I81055,I81414);
DFFARX1 I_4642 (I81431,I2507,I81021,I81007,);
nor I_4643 (I81462,I81115,I81397);
nor I_4644 (I80995,I81310,I81462);
nor I_4645 (I81004,I81245,I81380);
nor I_4646 (I80992,I81115,I81380);
not I_4647 (I81548,I2514);
DFFARX1 I_4648 (I470808,I2507,I81548,I81574,);
not I_4649 (I81582,I81574);
nand I_4650 (I81599,I470805,I470820);
and I_4651 (I81616,I81599,I470802);
DFFARX1 I_4652 (I81616,I2507,I81548,I81642,);
DFFARX1 I_4653 (I470799,I2507,I81548,I81659,);
and I_4654 (I81667,I81659,I470799);
nor I_4655 (I81684,I81642,I81667);
DFFARX1 I_4656 (I81684,I2507,I81548,I81516,);
nand I_4657 (I81715,I81659,I470799);
nand I_4658 (I81732,I81582,I81715);
not I_4659 (I81528,I81732);
DFFARX1 I_4660 (I470802,I2507,I81548,I81772,);
DFFARX1 I_4661 (I81772,I2507,I81548,I81537,);
nand I_4662 (I81794,I470814,I470805);
and I_4663 (I81811,I81794,I470817);
DFFARX1 I_4664 (I81811,I2507,I81548,I81837,);
DFFARX1 I_4665 (I81837,I2507,I81548,I81854,);
not I_4666 (I81540,I81854);
not I_4667 (I81876,I81837);
nand I_4668 (I81525,I81876,I81715);
nor I_4669 (I81907,I470811,I470805);
not I_4670 (I81924,I81907);
nor I_4671 (I81941,I81876,I81924);
nor I_4672 (I81958,I81582,I81941);
DFFARX1 I_4673 (I81958,I2507,I81548,I81534,);
nor I_4674 (I81989,I81642,I81924);
nor I_4675 (I81522,I81837,I81989);
nor I_4676 (I81531,I81772,I81907);
nor I_4677 (I81519,I81642,I81907);
not I_4678 (I82075,I2514);
DFFARX1 I_4679 (I457106,I2507,I82075,I82101,);
not I_4680 (I82109,I82101);
nand I_4681 (I82126,I457103,I457118);
and I_4682 (I82143,I82126,I457100);
DFFARX1 I_4683 (I82143,I2507,I82075,I82169,);
DFFARX1 I_4684 (I457097,I2507,I82075,I82186,);
and I_4685 (I82194,I82186,I457097);
nor I_4686 (I82211,I82169,I82194);
DFFARX1 I_4687 (I82211,I2507,I82075,I82043,);
nand I_4688 (I82242,I82186,I457097);
nand I_4689 (I82259,I82109,I82242);
not I_4690 (I82055,I82259);
DFFARX1 I_4691 (I457100,I2507,I82075,I82299,);
DFFARX1 I_4692 (I82299,I2507,I82075,I82064,);
nand I_4693 (I82321,I457112,I457103);
and I_4694 (I82338,I82321,I457115);
DFFARX1 I_4695 (I82338,I2507,I82075,I82364,);
DFFARX1 I_4696 (I82364,I2507,I82075,I82381,);
not I_4697 (I82067,I82381);
not I_4698 (I82403,I82364);
nand I_4699 (I82052,I82403,I82242);
nor I_4700 (I82434,I457109,I457103);
not I_4701 (I82451,I82434);
nor I_4702 (I82468,I82403,I82451);
nor I_4703 (I82485,I82109,I82468);
DFFARX1 I_4704 (I82485,I2507,I82075,I82061,);
nor I_4705 (I82516,I82169,I82451);
nor I_4706 (I82049,I82364,I82516);
nor I_4707 (I82058,I82299,I82434);
nor I_4708 (I82046,I82169,I82434);
not I_4709 (I82602,I2514);
DFFARX1 I_4710 (I506729,I2507,I82602,I82628,);
not I_4711 (I82636,I82628);
nand I_4712 (I82653,I506747,I506741);
and I_4713 (I82670,I82653,I506720);
DFFARX1 I_4714 (I82670,I2507,I82602,I82696,);
DFFARX1 I_4715 (I506738,I2507,I82602,I82713,);
and I_4716 (I82721,I82713,I506723);
nor I_4717 (I82738,I82696,I82721);
DFFARX1 I_4718 (I82738,I2507,I82602,I82570,);
nand I_4719 (I82769,I82713,I506723);
nand I_4720 (I82786,I82636,I82769);
not I_4721 (I82582,I82786);
DFFARX1 I_4722 (I506735,I2507,I82602,I82826,);
DFFARX1 I_4723 (I82826,I2507,I82602,I82591,);
nand I_4724 (I82848,I506744,I506732);
and I_4725 (I82865,I82848,I506726);
DFFARX1 I_4726 (I82865,I2507,I82602,I82891,);
DFFARX1 I_4727 (I82891,I2507,I82602,I82908,);
not I_4728 (I82594,I82908);
not I_4729 (I82930,I82891);
nand I_4730 (I82579,I82930,I82769);
nor I_4731 (I82961,I506720,I506732);
not I_4732 (I82978,I82961);
nor I_4733 (I82995,I82930,I82978);
nor I_4734 (I83012,I82636,I82995);
DFFARX1 I_4735 (I83012,I2507,I82602,I82588,);
nor I_4736 (I83043,I82696,I82978);
nor I_4737 (I82576,I82891,I83043);
nor I_4738 (I82585,I82826,I82961);
nor I_4739 (I82573,I82696,I82961);
not I_4740 (I83129,I2514);
DFFARX1 I_4741 (I342628,I2507,I83129,I83155,);
not I_4742 (I83163,I83155);
nand I_4743 (I83180,I342640,I342625);
and I_4744 (I83197,I83180,I342619);
DFFARX1 I_4745 (I83197,I2507,I83129,I83223,);
DFFARX1 I_4746 (I342634,I2507,I83129,I83240,);
and I_4747 (I83248,I83240,I342622);
nor I_4748 (I83265,I83223,I83248);
DFFARX1 I_4749 (I83265,I2507,I83129,I83097,);
nand I_4750 (I83296,I83240,I342622);
nand I_4751 (I83313,I83163,I83296);
not I_4752 (I83109,I83313);
DFFARX1 I_4753 (I342631,I2507,I83129,I83353,);
DFFARX1 I_4754 (I83353,I2507,I83129,I83118,);
nand I_4755 (I83375,I342637,I342643);
and I_4756 (I83392,I83375,I342619);
DFFARX1 I_4757 (I83392,I2507,I83129,I83418,);
DFFARX1 I_4758 (I83418,I2507,I83129,I83435,);
not I_4759 (I83121,I83435);
not I_4760 (I83457,I83418);
nand I_4761 (I83106,I83457,I83296);
nor I_4762 (I83488,I342622,I342643);
not I_4763 (I83505,I83488);
nor I_4764 (I83522,I83457,I83505);
nor I_4765 (I83539,I83163,I83522);
DFFARX1 I_4766 (I83539,I2507,I83129,I83115,);
nor I_4767 (I83570,I83223,I83505);
nor I_4768 (I83103,I83418,I83570);
nor I_4769 (I83112,I83353,I83488);
nor I_4770 (I83100,I83223,I83488);
not I_4771 (I83659,I2514);
DFFARX1 I_4772 (I458157,I2507,I83659,I83685,);
not I_4773 (I83693,I83685);
DFFARX1 I_4774 (I458157,I2507,I83659,I83719,);
not I_4775 (I83727,I458154);
or I_4776 (I83744,I458166,I458154);
nor I_4777 (I83761,I83719,I458166);
nand I_4778 (I83636,I83727,I83761);
nor I_4779 (I83792,I458160,I458166);
nand I_4780 (I83630,I83792,I83727);
not I_4781 (I83823,I458172);
nand I_4782 (I83840,I83727,I83823);
nor I_4783 (I83857,I458163,I458151);
not I_4784 (I83874,I83857);
nor I_4785 (I83891,I83874,I83840);
nor I_4786 (I83908,I83792,I83891);
DFFARX1 I_4787 (I83908,I2507,I83659,I83645,);
nor I_4788 (I83642,I83857,I83744);
DFFARX1 I_4789 (I83857,I2507,I83659,I83648,);
nor I_4790 (I83967,I83823,I458163);
nor I_4791 (I83984,I83967,I458154);
nor I_4792 (I84001,I458154,I458151);
DFFARX1 I_4793 (I84001,I2507,I83659,I84027,);
nor I_4794 (I83627,I84027,I83984);
DFFARX1 I_4795 (I84027,I2507,I83659,I84058,);
nand I_4796 (I84066,I84058,I458169);
nor I_4797 (I83651,I83693,I84066);
not I_4798 (I84097,I84027);
nand I_4799 (I84114,I84097,I458169);
nor I_4800 (I84131,I83693,I84114);
nor I_4801 (I83633,I83719,I84131);
nor I_4802 (I84162,I458154,I458160);
nor I_4803 (I84179,I83719,I84162);
DFFARX1 I_4804 (I84179,I2507,I83659,I83624,);
and I_4805 (I83639,I83792,I458154);
not I_4806 (I84254,I2514);
DFFARX1 I_4807 (I196428,I2507,I84254,I84280,);
not I_4808 (I84288,I84280);
DFFARX1 I_4809 (I196425,I2507,I84254,I84314,);
not I_4810 (I84322,I196422);
or I_4811 (I84339,I196434,I196422);
nor I_4812 (I84356,I84314,I196434);
nand I_4813 (I84231,I84322,I84356);
nor I_4814 (I84387,I196443,I196434);
nand I_4815 (I84225,I84387,I84322);
not I_4816 (I84418,I196440);
nand I_4817 (I84435,I84322,I84418);
nor I_4818 (I84452,I196419,I196419);
not I_4819 (I84469,I84452);
nor I_4820 (I84486,I84469,I84435);
nor I_4821 (I84503,I84387,I84486);
DFFARX1 I_4822 (I84503,I2507,I84254,I84240,);
nor I_4823 (I84237,I84452,I84339);
DFFARX1 I_4824 (I84452,I2507,I84254,I84243,);
nor I_4825 (I84562,I84418,I196419);
nor I_4826 (I84579,I84562,I196422);
nor I_4827 (I84596,I196431,I196446);
DFFARX1 I_4828 (I84596,I2507,I84254,I84622,);
nor I_4829 (I84222,I84622,I84579);
DFFARX1 I_4830 (I84622,I2507,I84254,I84653,);
nand I_4831 (I84661,I84653,I196437);
nor I_4832 (I84246,I84288,I84661);
not I_4833 (I84692,I84622);
nand I_4834 (I84709,I84692,I196437);
nor I_4835 (I84726,I84288,I84709);
nor I_4836 (I84228,I84314,I84726);
nor I_4837 (I84757,I196431,I196443);
nor I_4838 (I84774,I84314,I84757);
DFFARX1 I_4839 (I84774,I2507,I84254,I84219,);
and I_4840 (I84234,I84387,I196431);
not I_4841 (I84849,I2514);
DFFARX1 I_4842 (I674020,I2507,I84849,I84875,);
not I_4843 (I84883,I84875);
DFFARX1 I_4844 (I674017,I2507,I84849,I84909,);
not I_4845 (I84917,I674035);
or I_4846 (I84934,I674029,I674035);
nor I_4847 (I84951,I84909,I674029);
nand I_4848 (I84826,I84917,I84951);
nor I_4849 (I84982,I674023,I674029);
nand I_4850 (I84820,I84982,I84917);
not I_4851 (I85013,I674020);
nand I_4852 (I85030,I84917,I85013);
nor I_4853 (I85047,I674026,I674032);
not I_4854 (I85064,I85047);
nor I_4855 (I85081,I85064,I85030);
nor I_4856 (I85098,I84982,I85081);
DFFARX1 I_4857 (I85098,I2507,I84849,I84835,);
nor I_4858 (I84832,I85047,I84934);
DFFARX1 I_4859 (I85047,I2507,I84849,I84838,);
nor I_4860 (I85157,I85013,I674026);
nor I_4861 (I85174,I85157,I674035);
nor I_4862 (I85191,I674038,I674017);
DFFARX1 I_4863 (I85191,I2507,I84849,I85217,);
nor I_4864 (I84817,I85217,I85174);
DFFARX1 I_4865 (I85217,I2507,I84849,I85248,);
nand I_4866 (I85256,I85248,I674041);
nor I_4867 (I84841,I84883,I85256);
not I_4868 (I85287,I85217);
nand I_4869 (I85304,I85287,I674041);
nor I_4870 (I85321,I84883,I85304);
nor I_4871 (I84823,I84909,I85321);
nor I_4872 (I85352,I674038,I674023);
nor I_4873 (I85369,I84909,I85352);
DFFARX1 I_4874 (I85369,I2507,I84849,I84814,);
and I_4875 (I84829,I84982,I674038);
not I_4876 (I85444,I2514);
DFFARX1 I_4877 (I228080,I2507,I85444,I85470,);
not I_4878 (I85478,I85470);
DFFARX1 I_4879 (I228074,I2507,I85444,I85504,);
not I_4880 (I85512,I228071);
or I_4881 (I85529,I228062,I228071);
nor I_4882 (I85546,I85504,I228062);
nand I_4883 (I85421,I85512,I85546);
nor I_4884 (I85577,I228065,I228062);
nand I_4885 (I85415,I85577,I85512);
not I_4886 (I85608,I228068);
nand I_4887 (I85625,I85512,I85608);
nor I_4888 (I85642,I228056,I228083);
not I_4889 (I85659,I85642);
nor I_4890 (I85676,I85659,I85625);
nor I_4891 (I85693,I85577,I85676);
DFFARX1 I_4892 (I85693,I2507,I85444,I85430,);
nor I_4893 (I85427,I85642,I85529);
DFFARX1 I_4894 (I85642,I2507,I85444,I85433,);
nor I_4895 (I85752,I85608,I228056);
nor I_4896 (I85769,I85752,I228071);
nor I_4897 (I85786,I228059,I228056);
DFFARX1 I_4898 (I85786,I2507,I85444,I85812,);
nor I_4899 (I85412,I85812,I85769);
DFFARX1 I_4900 (I85812,I2507,I85444,I85843,);
nand I_4901 (I85851,I85843,I228077);
nor I_4902 (I85436,I85478,I85851);
not I_4903 (I85882,I85812);
nand I_4904 (I85899,I85882,I228077);
nor I_4905 (I85916,I85478,I85899);
nor I_4906 (I85418,I85504,I85916);
nor I_4907 (I85947,I228059,I228065);
nor I_4908 (I85964,I85504,I85947);
DFFARX1 I_4909 (I85964,I2507,I85444,I85409,);
and I_4910 (I85424,I85577,I228059);
not I_4911 (I86039,I2514);
DFFARX1 I_4912 (I201171,I2507,I86039,I86065,);
not I_4913 (I86073,I86065);
DFFARX1 I_4914 (I201168,I2507,I86039,I86099,);
not I_4915 (I86107,I201165);
or I_4916 (I86124,I201177,I201165);
nor I_4917 (I86141,I86099,I201177);
nand I_4918 (I86016,I86107,I86141);
nor I_4919 (I86172,I201186,I201177);
nand I_4920 (I86010,I86172,I86107);
not I_4921 (I86203,I201183);
nand I_4922 (I86220,I86107,I86203);
nor I_4923 (I86237,I201162,I201162);
not I_4924 (I86254,I86237);
nor I_4925 (I86271,I86254,I86220);
nor I_4926 (I86288,I86172,I86271);
DFFARX1 I_4927 (I86288,I2507,I86039,I86025,);
nor I_4928 (I86022,I86237,I86124);
DFFARX1 I_4929 (I86237,I2507,I86039,I86028,);
nor I_4930 (I86347,I86203,I201162);
nor I_4931 (I86364,I86347,I201165);
nor I_4932 (I86381,I201174,I201189);
DFFARX1 I_4933 (I86381,I2507,I86039,I86407,);
nor I_4934 (I86007,I86407,I86364);
DFFARX1 I_4935 (I86407,I2507,I86039,I86438,);
nand I_4936 (I86446,I86438,I201180);
nor I_4937 (I86031,I86073,I86446);
not I_4938 (I86477,I86407);
nand I_4939 (I86494,I86477,I201180);
nor I_4940 (I86511,I86073,I86494);
nor I_4941 (I86013,I86099,I86511);
nor I_4942 (I86542,I201174,I201186);
nor I_4943 (I86559,I86099,I86542);
DFFARX1 I_4944 (I86559,I2507,I86039,I86004,);
and I_4945 (I86019,I86172,I201174);
not I_4946 (I86634,I2514);
DFFARX1 I_4947 (I471859,I2507,I86634,I86660,);
not I_4948 (I86668,I86660);
DFFARX1 I_4949 (I471859,I2507,I86634,I86694,);
not I_4950 (I86702,I471856);
or I_4951 (I86719,I471868,I471856);
nor I_4952 (I86736,I86694,I471868);
nand I_4953 (I86611,I86702,I86736);
nor I_4954 (I86767,I471862,I471868);
nand I_4955 (I86605,I86767,I86702);
not I_4956 (I86798,I471874);
nand I_4957 (I86815,I86702,I86798);
nor I_4958 (I86832,I471865,I471853);
not I_4959 (I86849,I86832);
nor I_4960 (I86866,I86849,I86815);
nor I_4961 (I86883,I86767,I86866);
DFFARX1 I_4962 (I86883,I2507,I86634,I86620,);
nor I_4963 (I86617,I86832,I86719);
DFFARX1 I_4964 (I86832,I2507,I86634,I86623,);
nor I_4965 (I86942,I86798,I471865);
nor I_4966 (I86959,I86942,I471856);
nor I_4967 (I86976,I471856,I471853);
DFFARX1 I_4968 (I86976,I2507,I86634,I87002,);
nor I_4969 (I86602,I87002,I86959);
DFFARX1 I_4970 (I87002,I2507,I86634,I87033,);
nand I_4971 (I87041,I87033,I471871);
nor I_4972 (I86626,I86668,I87041);
not I_4973 (I87072,I87002);
nand I_4974 (I87089,I87072,I471871);
nor I_4975 (I87106,I86668,I87089);
nor I_4976 (I86608,I86694,I87106);
nor I_4977 (I87137,I471856,I471862);
nor I_4978 (I87154,I86694,I87137);
DFFARX1 I_4979 (I87154,I2507,I86634,I86599,);
and I_4980 (I86614,I86767,I471856);
not I_4981 (I87229,I2514);
DFFARX1 I_4982 (I2260,I2507,I87229,I87255,);
not I_4983 (I87263,I87255);
DFFARX1 I_4984 (I2460,I2507,I87229,I87289,);
not I_4985 (I87297,I2092);
or I_4986 (I87314,I1988,I2092);
nor I_4987 (I87331,I87289,I1988);
nand I_4988 (I87206,I87297,I87331);
nor I_4989 (I87362,I1868,I1988);
nand I_4990 (I87200,I87362,I87297);
not I_4991 (I87393,I2452);
nand I_4992 (I87410,I87297,I87393);
nor I_4993 (I87427,I1692,I1772);
not I_4994 (I87444,I87427);
nor I_4995 (I87461,I87444,I87410);
nor I_4996 (I87478,I87362,I87461);
DFFARX1 I_4997 (I87478,I2507,I87229,I87215,);
nor I_4998 (I87212,I87427,I87314);
DFFARX1 I_4999 (I87427,I2507,I87229,I87218,);
nor I_5000 (I87537,I87393,I1692);
nor I_5001 (I87554,I87537,I2092);
nor I_5002 (I87571,I1388,I1964);
DFFARX1 I_5003 (I87571,I2507,I87229,I87597,);
nor I_5004 (I87197,I87597,I87554);
DFFARX1 I_5005 (I87597,I2507,I87229,I87628,);
nand I_5006 (I87636,I87628,I2284);
nor I_5007 (I87221,I87263,I87636);
not I_5008 (I87667,I87597);
nand I_5009 (I87684,I87667,I2284);
nor I_5010 (I87701,I87263,I87684);
nor I_5011 (I87203,I87289,I87701);
nor I_5012 (I87732,I1388,I1868);
nor I_5013 (I87749,I87289,I87732);
DFFARX1 I_5014 (I87749,I2507,I87229,I87194,);
and I_5015 (I87209,I87362,I1388);
not I_5016 (I87824,I2514);
DFFARX1 I_5017 (I617920,I2507,I87824,I87850,);
not I_5018 (I87858,I87850);
DFFARX1 I_5019 (I617917,I2507,I87824,I87884,);
not I_5020 (I87892,I617926);
or I_5021 (I87909,I617917,I617926);
nor I_5022 (I87926,I87884,I617917);
nand I_5023 (I87801,I87892,I87926);
nor I_5024 (I87957,I617929,I617917);
nand I_5025 (I87795,I87957,I87892);
not I_5026 (I87988,I617923);
nand I_5027 (I88005,I87892,I87988);
nor I_5028 (I88022,I617920,I617938);
not I_5029 (I88039,I88022);
nor I_5030 (I88056,I88039,I88005);
nor I_5031 (I88073,I87957,I88056);
DFFARX1 I_5032 (I88073,I2507,I87824,I87810,);
nor I_5033 (I87807,I88022,I87909);
DFFARX1 I_5034 (I88022,I2507,I87824,I87813,);
nor I_5035 (I88132,I87988,I617920);
nor I_5036 (I88149,I88132,I617926);
nor I_5037 (I88166,I617941,I617935);
DFFARX1 I_5038 (I88166,I2507,I87824,I88192,);
nor I_5039 (I87792,I88192,I88149);
DFFARX1 I_5040 (I88192,I2507,I87824,I88223,);
nand I_5041 (I88231,I88223,I617932);
nor I_5042 (I87816,I87858,I88231);
not I_5043 (I88262,I88192);
nand I_5044 (I88279,I88262,I617932);
nor I_5045 (I88296,I87858,I88279);
nor I_5046 (I87798,I87884,I88296);
nor I_5047 (I88327,I617941,I617929);
nor I_5048 (I88344,I87884,I88327);
DFFARX1 I_5049 (I88344,I2507,I87824,I87789,);
and I_5050 (I87804,I87957,I617941);
not I_5051 (I88416,I2514);
DFFARX1 I_5052 (I603467,I2507,I88416,I88442,);
DFFARX1 I_5053 (I88442,I2507,I88416,I88459,);
not I_5054 (I88408,I88459);
not I_5055 (I88481,I88442);
DFFARX1 I_5056 (I603467,I2507,I88416,I88507,);
not I_5057 (I88515,I88507);
and I_5058 (I88532,I88481,I603470);
not I_5059 (I88549,I603482);
nand I_5060 (I88566,I88549,I603470);
not I_5061 (I88583,I603488);
nor I_5062 (I88600,I88583,I603479);
nand I_5063 (I88617,I88600,I603485);
nor I_5064 (I88634,I88617,I88566);
DFFARX1 I_5065 (I88634,I2507,I88416,I88384,);
not I_5066 (I88665,I88617);
not I_5067 (I88682,I603479);
nand I_5068 (I88699,I88682,I603470);
nor I_5069 (I88716,I603479,I603482);
nand I_5070 (I88396,I88532,I88716);
nand I_5071 (I88390,I88481,I603479);
nand I_5072 (I88761,I88583,I603476);
DFFARX1 I_5073 (I88761,I2507,I88416,I88405,);
DFFARX1 I_5074 (I88761,I2507,I88416,I88399,);
not I_5075 (I88806,I603476);
nor I_5076 (I88823,I88806,I603473);
and I_5077 (I88840,I88823,I603491);
or I_5078 (I88857,I88840,I603470);
DFFARX1 I_5079 (I88857,I2507,I88416,I88883,);
nand I_5080 (I88891,I88883,I88549);
nor I_5081 (I88393,I88891,I88699);
nor I_5082 (I88387,I88883,I88515);
DFFARX1 I_5083 (I88883,I2507,I88416,I88945,);
not I_5084 (I88953,I88945);
nor I_5085 (I88402,I88953,I88665);
not I_5086 (I89011,I2514);
DFFARX1 I_5087 (I554255,I2507,I89011,I89037,);
DFFARX1 I_5088 (I89037,I2507,I89011,I89054,);
not I_5089 (I89003,I89054);
not I_5090 (I89076,I89037);
DFFARX1 I_5091 (I554264,I2507,I89011,I89102,);
not I_5092 (I89110,I89102);
and I_5093 (I89127,I89076,I554258);
not I_5094 (I89144,I554252);
nand I_5095 (I89161,I89144,I554258);
not I_5096 (I89178,I554267);
nor I_5097 (I89195,I89178,I554255);
nand I_5098 (I89212,I89195,I554261);
nor I_5099 (I89229,I89212,I89161);
DFFARX1 I_5100 (I89229,I2507,I89011,I88979,);
not I_5101 (I89260,I89212);
not I_5102 (I89277,I554255);
nand I_5103 (I89294,I89277,I554258);
nor I_5104 (I89311,I554255,I554252);
nand I_5105 (I88991,I89127,I89311);
nand I_5106 (I88985,I89076,I554255);
nand I_5107 (I89356,I89178,I554258);
DFFARX1 I_5108 (I89356,I2507,I89011,I89000,);
DFFARX1 I_5109 (I89356,I2507,I89011,I88994,);
not I_5110 (I89401,I554258);
nor I_5111 (I89418,I89401,I554273);
and I_5112 (I89435,I89418,I554270);
or I_5113 (I89452,I89435,I554252);
DFFARX1 I_5114 (I89452,I2507,I89011,I89478,);
nand I_5115 (I89486,I89478,I89144);
nor I_5116 (I88988,I89486,I89294);
nor I_5117 (I88982,I89478,I89110);
DFFARX1 I_5118 (I89478,I2507,I89011,I89540,);
not I_5119 (I89548,I89540);
nor I_5120 (I88997,I89548,I89260);
not I_5121 (I89606,I2514);
DFFARX1 I_5122 (I367485,I2507,I89606,I89632,);
DFFARX1 I_5123 (I89632,I2507,I89606,I89649,);
not I_5124 (I89598,I89649);
not I_5125 (I89671,I89632);
DFFARX1 I_5126 (I367482,I2507,I89606,I89697,);
not I_5127 (I89705,I89697);
and I_5128 (I89722,I89671,I367488);
not I_5129 (I89739,I367473);
nand I_5130 (I89756,I89739,I367488);
not I_5131 (I89773,I367476);
nor I_5132 (I89790,I89773,I367497);
nand I_5133 (I89807,I89790,I367494);
nor I_5134 (I89824,I89807,I89756);
DFFARX1 I_5135 (I89824,I2507,I89606,I89574,);
not I_5136 (I89855,I89807);
not I_5137 (I89872,I367497);
nand I_5138 (I89889,I89872,I367488);
nor I_5139 (I89906,I367497,I367473);
nand I_5140 (I89586,I89722,I89906);
nand I_5141 (I89580,I89671,I367497);
nand I_5142 (I89951,I89773,I367473);
DFFARX1 I_5143 (I89951,I2507,I89606,I89595,);
DFFARX1 I_5144 (I89951,I2507,I89606,I89589,);
not I_5145 (I89996,I367473);
nor I_5146 (I90013,I89996,I367479);
and I_5147 (I90030,I90013,I367491);
or I_5148 (I90047,I90030,I367476);
DFFARX1 I_5149 (I90047,I2507,I89606,I90073,);
nand I_5150 (I90081,I90073,I89739);
nor I_5151 (I89583,I90081,I89889);
nor I_5152 (I89577,I90073,I89705);
DFFARX1 I_5153 (I90073,I2507,I89606,I90135,);
not I_5154 (I90143,I90135);
nor I_5155 (I89592,I90143,I89855);
not I_5156 (I90201,I2514);
DFFARX1 I_5157 (I594797,I2507,I90201,I90227,);
DFFARX1 I_5158 (I90227,I2507,I90201,I90244,);
not I_5159 (I90193,I90244);
not I_5160 (I90266,I90227);
DFFARX1 I_5161 (I594797,I2507,I90201,I90292,);
not I_5162 (I90300,I90292);
and I_5163 (I90317,I90266,I594800);
not I_5164 (I90334,I594812);
nand I_5165 (I90351,I90334,I594800);
not I_5166 (I90368,I594818);
nor I_5167 (I90385,I90368,I594809);
nand I_5168 (I90402,I90385,I594815);
nor I_5169 (I90419,I90402,I90351);
DFFARX1 I_5170 (I90419,I2507,I90201,I90169,);
not I_5171 (I90450,I90402);
not I_5172 (I90467,I594809);
nand I_5173 (I90484,I90467,I594800);
nor I_5174 (I90501,I594809,I594812);
nand I_5175 (I90181,I90317,I90501);
nand I_5176 (I90175,I90266,I594809);
nand I_5177 (I90546,I90368,I594806);
DFFARX1 I_5178 (I90546,I2507,I90201,I90190,);
DFFARX1 I_5179 (I90546,I2507,I90201,I90184,);
not I_5180 (I90591,I594806);
nor I_5181 (I90608,I90591,I594803);
and I_5182 (I90625,I90608,I594821);
or I_5183 (I90642,I90625,I594800);
DFFARX1 I_5184 (I90642,I2507,I90201,I90668,);
nand I_5185 (I90676,I90668,I90334);
nor I_5186 (I90178,I90676,I90484);
nor I_5187 (I90172,I90668,I90300);
DFFARX1 I_5188 (I90668,I2507,I90201,I90730,);
not I_5189 (I90738,I90730);
nor I_5190 (I90187,I90738,I90450);
not I_5191 (I90796,I2514);
DFFARX1 I_5192 (I531929,I2507,I90796,I90822,);
DFFARX1 I_5193 (I90822,I2507,I90796,I90839,);
not I_5194 (I90788,I90839);
not I_5195 (I90861,I90822);
DFFARX1 I_5196 (I531938,I2507,I90796,I90887,);
not I_5197 (I90895,I90887);
and I_5198 (I90912,I90861,I531926);
not I_5199 (I90929,I531917);
nand I_5200 (I90946,I90929,I531926);
not I_5201 (I90963,I531923);
nor I_5202 (I90980,I90963,I531941);
nand I_5203 (I90997,I90980,I531914);
nor I_5204 (I91014,I90997,I90946);
DFFARX1 I_5205 (I91014,I2507,I90796,I90764,);
not I_5206 (I91045,I90997);
not I_5207 (I91062,I531941);
nand I_5208 (I91079,I91062,I531926);
nor I_5209 (I91096,I531941,I531917);
nand I_5210 (I90776,I90912,I91096);
nand I_5211 (I90770,I90861,I531941);
nand I_5212 (I91141,I90963,I531920);
DFFARX1 I_5213 (I91141,I2507,I90796,I90785,);
DFFARX1 I_5214 (I91141,I2507,I90796,I90779,);
not I_5215 (I91186,I531920);
nor I_5216 (I91203,I91186,I531932);
and I_5217 (I91220,I91203,I531914);
or I_5218 (I91237,I91220,I531935);
DFFARX1 I_5219 (I91237,I2507,I90796,I91263,);
nand I_5220 (I91271,I91263,I90929);
nor I_5221 (I90773,I91271,I91079);
nor I_5222 (I90767,I91263,I90895);
DFFARX1 I_5223 (I91263,I2507,I90796,I91325,);
not I_5224 (I91333,I91325);
nor I_5225 (I90782,I91333,I91045);
not I_5226 (I91391,I2514);
DFFARX1 I_5227 (I2268,I2507,I91391,I91417,);
DFFARX1 I_5228 (I91417,I2507,I91391,I91434,);
not I_5229 (I91383,I91434);
not I_5230 (I91456,I91417);
DFFARX1 I_5231 (I2380,I2507,I91391,I91482,);
not I_5232 (I91490,I91482);
and I_5233 (I91507,I91456,I2404);
not I_5234 (I91524,I2476);
nand I_5235 (I91541,I91524,I2404);
not I_5236 (I91558,I2332);
nor I_5237 (I91575,I91558,I1548);
nand I_5238 (I91592,I91575,I1788);
nor I_5239 (I91609,I91592,I91541);
DFFARX1 I_5240 (I91609,I2507,I91391,I91359,);
not I_5241 (I91640,I91592);
not I_5242 (I91657,I1548);
nand I_5243 (I91674,I91657,I2404);
nor I_5244 (I91691,I1548,I2476);
nand I_5245 (I91371,I91507,I91691);
nand I_5246 (I91365,I91456,I1548);
nand I_5247 (I91736,I91558,I1516);
DFFARX1 I_5248 (I91736,I2507,I91391,I91380,);
DFFARX1 I_5249 (I91736,I2507,I91391,I91374,);
not I_5250 (I91781,I1516);
nor I_5251 (I91798,I91781,I2228);
and I_5252 (I91815,I91798,I1436);
or I_5253 (I91832,I91815,I2028);
DFFARX1 I_5254 (I91832,I2507,I91391,I91858,);
nand I_5255 (I91866,I91858,I91524);
nor I_5256 (I91368,I91866,I91674);
nor I_5257 (I91362,I91858,I91490);
DFFARX1 I_5258 (I91858,I2507,I91391,I91920,);
not I_5259 (I91928,I91920);
nor I_5260 (I91377,I91928,I91640);
not I_5261 (I91986,I2514);
DFFARX1 I_5262 (I615605,I2507,I91986,I92012,);
DFFARX1 I_5263 (I92012,I2507,I91986,I92029,);
not I_5264 (I91978,I92029);
not I_5265 (I92051,I92012);
DFFARX1 I_5266 (I615605,I2507,I91986,I92077,);
not I_5267 (I92085,I92077);
and I_5268 (I92102,I92051,I615608);
not I_5269 (I92119,I615620);
nand I_5270 (I92136,I92119,I615608);
not I_5271 (I92153,I615626);
nor I_5272 (I92170,I92153,I615617);
nand I_5273 (I92187,I92170,I615623);
nor I_5274 (I92204,I92187,I92136);
DFFARX1 I_5275 (I92204,I2507,I91986,I91954,);
not I_5276 (I92235,I92187);
not I_5277 (I92252,I615617);
nand I_5278 (I92269,I92252,I615608);
nor I_5279 (I92286,I615617,I615620);
nand I_5280 (I91966,I92102,I92286);
nand I_5281 (I91960,I92051,I615617);
nand I_5282 (I92331,I92153,I615614);
DFFARX1 I_5283 (I92331,I2507,I91986,I91975,);
DFFARX1 I_5284 (I92331,I2507,I91986,I91969,);
not I_5285 (I92376,I615614);
nor I_5286 (I92393,I92376,I615611);
and I_5287 (I92410,I92393,I615629);
or I_5288 (I92427,I92410,I615608);
DFFARX1 I_5289 (I92427,I2507,I91986,I92453,);
nand I_5290 (I92461,I92453,I92119);
nor I_5291 (I91963,I92461,I92269);
nor I_5292 (I91957,I92453,I92085);
DFFARX1 I_5293 (I92453,I2507,I91986,I92515,);
not I_5294 (I92523,I92515);
nor I_5295 (I91972,I92523,I92235);
not I_5296 (I92581,I2514);
DFFARX1 I_5297 (I340322,I2507,I92581,I92607,);
DFFARX1 I_5298 (I92607,I2507,I92581,I92624,);
not I_5299 (I92573,I92624);
not I_5300 (I92646,I92607);
DFFARX1 I_5301 (I340313,I2507,I92581,I92672,);
not I_5302 (I92680,I92672);
and I_5303 (I92697,I92646,I340331);
not I_5304 (I92714,I340328);
nand I_5305 (I92731,I92714,I340331);
not I_5306 (I92748,I340307);
nor I_5307 (I92765,I92748,I340310);
nand I_5308 (I92782,I92765,I340319);
nor I_5309 (I92799,I92782,I92731);
DFFARX1 I_5310 (I92799,I2507,I92581,I92549,);
not I_5311 (I92830,I92782);
not I_5312 (I92847,I340310);
nand I_5313 (I92864,I92847,I340331);
nor I_5314 (I92881,I340310,I340328);
nand I_5315 (I92561,I92697,I92881);
nand I_5316 (I92555,I92646,I340310);
nand I_5317 (I92926,I92748,I340325);
DFFARX1 I_5318 (I92926,I2507,I92581,I92570,);
DFFARX1 I_5319 (I92926,I2507,I92581,I92564,);
not I_5320 (I92971,I340325);
nor I_5321 (I92988,I92971,I340307);
and I_5322 (I93005,I92988,I340316);
or I_5323 (I93022,I93005,I340310);
DFFARX1 I_5324 (I93022,I2507,I92581,I93048,);
nand I_5325 (I93056,I93048,I92714);
nor I_5326 (I92558,I93056,I92864);
nor I_5327 (I92552,I93048,I92680);
DFFARX1 I_5328 (I93048,I2507,I92581,I93110,);
not I_5329 (I93118,I93110);
nor I_5330 (I92567,I93118,I92830);
not I_5331 (I93176,I2514);
DFFARX1 I_5332 (I665928,I2507,I93176,I93202,);
DFFARX1 I_5333 (I93202,I2507,I93176,I93219,);
not I_5334 (I93168,I93219);
not I_5335 (I93241,I93202);
DFFARX1 I_5336 (I665940,I2507,I93176,I93267,);
not I_5337 (I93275,I93267);
and I_5338 (I93292,I93241,I665934);
not I_5339 (I93309,I665946);
nand I_5340 (I93326,I93309,I665934);
not I_5341 (I93343,I665931);
nor I_5342 (I93360,I93343,I665943);
nand I_5343 (I93377,I93360,I665925);
nor I_5344 (I93394,I93377,I93326);
DFFARX1 I_5345 (I93394,I2507,I93176,I93144,);
not I_5346 (I93425,I93377);
not I_5347 (I93442,I665943);
nand I_5348 (I93459,I93442,I665934);
nor I_5349 (I93476,I665943,I665946);
nand I_5350 (I93156,I93292,I93476);
nand I_5351 (I93150,I93241,I665943);
nand I_5352 (I93521,I93343,I665937);
DFFARX1 I_5353 (I93521,I2507,I93176,I93165,);
DFFARX1 I_5354 (I93521,I2507,I93176,I93159,);
not I_5355 (I93566,I665937);
nor I_5356 (I93583,I93566,I665928);
and I_5357 (I93600,I93583,I665925);
or I_5358 (I93617,I93600,I665949);
DFFARX1 I_5359 (I93617,I2507,I93176,I93643,);
nand I_5360 (I93651,I93643,I93309);
nor I_5361 (I93153,I93651,I93459);
nor I_5362 (I93147,I93643,I93275);
DFFARX1 I_5363 (I93643,I2507,I93176,I93705,);
not I_5364 (I93713,I93705);
nor I_5365 (I93162,I93713,I93425);
not I_5366 (I93771,I2514);
DFFARX1 I_5367 (I719224,I2507,I93771,I93797,);
DFFARX1 I_5368 (I93797,I2507,I93771,I93814,);
not I_5369 (I93763,I93814);
not I_5370 (I93836,I93797);
DFFARX1 I_5371 (I719215,I2507,I93771,I93862,);
not I_5372 (I93870,I93862);
and I_5373 (I93887,I93836,I719209);
not I_5374 (I93904,I719203);
nand I_5375 (I93921,I93904,I719209);
not I_5376 (I93938,I719230);
nor I_5377 (I93955,I93938,I719203);
nand I_5378 (I93972,I93955,I719227);
nor I_5379 (I93989,I93972,I93921);
DFFARX1 I_5380 (I93989,I2507,I93771,I93739,);
not I_5381 (I94020,I93972);
not I_5382 (I94037,I719203);
nand I_5383 (I94054,I94037,I719209);
nor I_5384 (I94071,I719203,I719203);
nand I_5385 (I93751,I93887,I94071);
nand I_5386 (I93745,I93836,I719203);
nand I_5387 (I94116,I93938,I719212);
DFFARX1 I_5388 (I94116,I2507,I93771,I93760,);
DFFARX1 I_5389 (I94116,I2507,I93771,I93754,);
not I_5390 (I94161,I719212);
nor I_5391 (I94178,I94161,I719218);
and I_5392 (I94195,I94178,I719221);
or I_5393 (I94212,I94195,I719206);
DFFARX1 I_5394 (I94212,I2507,I93771,I94238,);
nand I_5395 (I94246,I94238,I93904);
nor I_5396 (I93748,I94246,I94054);
nor I_5397 (I93742,I94238,I93870);
DFFARX1 I_5398 (I94238,I2507,I93771,I94300,);
not I_5399 (I94308,I94300);
nor I_5400 (I93757,I94308,I94020);
not I_5401 (I94366,I2514);
DFFARX1 I_5402 (I53067,I2507,I94366,I94392,);
DFFARX1 I_5403 (I94392,I2507,I94366,I94409,);
not I_5404 (I94358,I94409);
not I_5405 (I94431,I94392);
DFFARX1 I_5406 (I53061,I2507,I94366,I94457,);
not I_5407 (I94465,I94457);
and I_5408 (I94482,I94431,I53058);
not I_5409 (I94499,I53079);
nand I_5410 (I94516,I94499,I53058);
not I_5411 (I94533,I53073);
nor I_5412 (I94550,I94533,I53064);
nand I_5413 (I94567,I94550,I53070);
nor I_5414 (I94584,I94567,I94516);
DFFARX1 I_5415 (I94584,I2507,I94366,I94334,);
not I_5416 (I94615,I94567);
not I_5417 (I94632,I53064);
nand I_5418 (I94649,I94632,I53058);
nor I_5419 (I94666,I53064,I53079);
nand I_5420 (I94346,I94482,I94666);
nand I_5421 (I94340,I94431,I53064);
nand I_5422 (I94711,I94533,I53058);
DFFARX1 I_5423 (I94711,I2507,I94366,I94355,);
DFFARX1 I_5424 (I94711,I2507,I94366,I94349,);
not I_5425 (I94756,I53058);
nor I_5426 (I94773,I94756,I53076);
and I_5427 (I94790,I94773,I53082);
or I_5428 (I94807,I94790,I53061);
DFFARX1 I_5429 (I94807,I2507,I94366,I94833,);
nand I_5430 (I94841,I94833,I94499);
nor I_5431 (I94343,I94841,I94649);
nor I_5432 (I94337,I94833,I94465);
DFFARX1 I_5433 (I94833,I2507,I94366,I94895,);
not I_5434 (I94903,I94895);
nor I_5435 (I94352,I94903,I94615);
not I_5436 (I94961,I2514);
DFFARX1 I_5437 (I510611,I2507,I94961,I94987,);
DFFARX1 I_5438 (I94987,I2507,I94961,I95004,);
not I_5439 (I94953,I95004);
not I_5440 (I95026,I94987);
DFFARX1 I_5441 (I510620,I2507,I94961,I95052,);
not I_5442 (I95060,I95052);
and I_5443 (I95077,I95026,I510608);
not I_5444 (I95094,I510599);
nand I_5445 (I95111,I95094,I510608);
not I_5446 (I95128,I510605);
nor I_5447 (I95145,I95128,I510623);
nand I_5448 (I95162,I95145,I510596);
nor I_5449 (I95179,I95162,I95111);
DFFARX1 I_5450 (I95179,I2507,I94961,I94929,);
not I_5451 (I95210,I95162);
not I_5452 (I95227,I510623);
nand I_5453 (I95244,I95227,I510608);
nor I_5454 (I95261,I510623,I510599);
nand I_5455 (I94941,I95077,I95261);
nand I_5456 (I94935,I95026,I510623);
nand I_5457 (I95306,I95128,I510602);
DFFARX1 I_5458 (I95306,I2507,I94961,I94950,);
DFFARX1 I_5459 (I95306,I2507,I94961,I94944,);
not I_5460 (I95351,I510602);
nor I_5461 (I95368,I95351,I510614);
and I_5462 (I95385,I95368,I510596);
or I_5463 (I95402,I95385,I510617);
DFFARX1 I_5464 (I95402,I2507,I94961,I95428,);
nand I_5465 (I95436,I95428,I95094);
nor I_5466 (I94938,I95436,I95244);
nor I_5467 (I94932,I95428,I95060);
DFFARX1 I_5468 (I95428,I2507,I94961,I95490,);
not I_5469 (I95498,I95490);
nor I_5470 (I94947,I95498,I95210);
not I_5471 (I95556,I2514);
DFFARX1 I_5472 (I355347,I2507,I95556,I95582,);
DFFARX1 I_5473 (I95582,I2507,I95556,I95599,);
not I_5474 (I95548,I95599);
not I_5475 (I95621,I95582);
DFFARX1 I_5476 (I355344,I2507,I95556,I95647,);
not I_5477 (I95655,I95647);
and I_5478 (I95672,I95621,I355350);
not I_5479 (I95689,I355335);
nand I_5480 (I95706,I95689,I355350);
not I_5481 (I95723,I355338);
nor I_5482 (I95740,I95723,I355359);
nand I_5483 (I95757,I95740,I355356);
nor I_5484 (I95774,I95757,I95706);
DFFARX1 I_5485 (I95774,I2507,I95556,I95524,);
not I_5486 (I95805,I95757);
not I_5487 (I95822,I355359);
nand I_5488 (I95839,I95822,I355350);
nor I_5489 (I95856,I355359,I355335);
nand I_5490 (I95536,I95672,I95856);
nand I_5491 (I95530,I95621,I355359);
nand I_5492 (I95901,I95723,I355335);
DFFARX1 I_5493 (I95901,I2507,I95556,I95545,);
DFFARX1 I_5494 (I95901,I2507,I95556,I95539,);
not I_5495 (I95946,I355335);
nor I_5496 (I95963,I95946,I355341);
and I_5497 (I95980,I95963,I355353);
or I_5498 (I95997,I95980,I355338);
DFFARX1 I_5499 (I95997,I2507,I95556,I96023,);
nand I_5500 (I96031,I96023,I95689);
nor I_5501 (I95533,I96031,I95839);
nor I_5502 (I95527,I96023,I95655);
DFFARX1 I_5503 (I96023,I2507,I95556,I96085,);
not I_5504 (I96093,I96085);
nor I_5505 (I95542,I96093,I95805);
not I_5506 (I96151,I2514);
DFFARX1 I_5507 (I223823,I2507,I96151,I96177,);
DFFARX1 I_5508 (I96177,I2507,I96151,I96194,);
not I_5509 (I96143,I96194);
not I_5510 (I96216,I96177);
DFFARX1 I_5511 (I223838,I2507,I96151,I96242,);
not I_5512 (I96250,I96242);
and I_5513 (I96267,I96216,I223835);
not I_5514 (I96284,I223823);
nand I_5515 (I96301,I96284,I223835);
not I_5516 (I96318,I223832);
nor I_5517 (I96335,I96318,I223847);
nand I_5518 (I96352,I96335,I223844);
nor I_5519 (I96369,I96352,I96301);
DFFARX1 I_5520 (I96369,I2507,I96151,I96119,);
not I_5521 (I96400,I96352);
not I_5522 (I96417,I223847);
nand I_5523 (I96434,I96417,I223835);
nor I_5524 (I96451,I223847,I223823);
nand I_5525 (I96131,I96267,I96451);
nand I_5526 (I96125,I96216,I223847);
nand I_5527 (I96496,I96318,I223841);
DFFARX1 I_5528 (I96496,I2507,I96151,I96140,);
DFFARX1 I_5529 (I96496,I2507,I96151,I96134,);
not I_5530 (I96541,I223841);
nor I_5531 (I96558,I96541,I223829);
and I_5532 (I96575,I96558,I223850);
or I_5533 (I96592,I96575,I223826);
DFFARX1 I_5534 (I96592,I2507,I96151,I96618,);
nand I_5535 (I96626,I96618,I96284);
nor I_5536 (I96128,I96626,I96434);
nor I_5537 (I96122,I96618,I96250);
DFFARX1 I_5538 (I96618,I2507,I96151,I96680,);
not I_5539 (I96688,I96680);
nor I_5540 (I96137,I96688,I96400);
not I_5541 (I96746,I2514);
DFFARX1 I_5542 (I231344,I2507,I96746,I96772,);
DFFARX1 I_5543 (I96772,I2507,I96746,I96789,);
not I_5544 (I96738,I96789);
not I_5545 (I96811,I96772);
DFFARX1 I_5546 (I231332,I2507,I96746,I96837,);
not I_5547 (I96845,I96837);
and I_5548 (I96862,I96811,I231341);
not I_5549 (I96879,I231338);
nand I_5550 (I96896,I96879,I231341);
not I_5551 (I96913,I231329);
nor I_5552 (I96930,I96913,I231335);
nand I_5553 (I96947,I96930,I231320);
nor I_5554 (I96964,I96947,I96896);
DFFARX1 I_5555 (I96964,I2507,I96746,I96714,);
not I_5556 (I96995,I96947);
not I_5557 (I97012,I231335);
nand I_5558 (I97029,I97012,I231341);
nor I_5559 (I97046,I231335,I231338);
nand I_5560 (I96726,I96862,I97046);
nand I_5561 (I96720,I96811,I231335);
nand I_5562 (I97091,I96913,I231320);
DFFARX1 I_5563 (I97091,I2507,I96746,I96735,);
DFFARX1 I_5564 (I97091,I2507,I96746,I96729,);
not I_5565 (I97136,I231320);
nor I_5566 (I97153,I97136,I231326);
and I_5567 (I97170,I97153,I231323);
or I_5568 (I97187,I97170,I231347);
DFFARX1 I_5569 (I97187,I2507,I96746,I97213,);
nand I_5570 (I97221,I97213,I96879);
nor I_5571 (I96723,I97221,I97029);
nor I_5572 (I96717,I97213,I96845);
DFFARX1 I_5573 (I97213,I2507,I96746,I97275,);
not I_5574 (I97283,I97275);
nor I_5575 (I96732,I97283,I96995);
not I_5576 (I97341,I2514);
DFFARX1 I_5577 (I221188,I2507,I97341,I97367,);
DFFARX1 I_5578 (I97367,I2507,I97341,I97384,);
not I_5579 (I97333,I97384);
not I_5580 (I97406,I97367);
DFFARX1 I_5581 (I221203,I2507,I97341,I97432,);
not I_5582 (I97440,I97432);
and I_5583 (I97457,I97406,I221200);
not I_5584 (I97474,I221188);
nand I_5585 (I97491,I97474,I221200);
not I_5586 (I97508,I221197);
nor I_5587 (I97525,I97508,I221212);
nand I_5588 (I97542,I97525,I221209);
nor I_5589 (I97559,I97542,I97491);
DFFARX1 I_5590 (I97559,I2507,I97341,I97309,);
not I_5591 (I97590,I97542);
not I_5592 (I97607,I221212);
nand I_5593 (I97624,I97607,I221200);
nor I_5594 (I97641,I221212,I221188);
nand I_5595 (I97321,I97457,I97641);
nand I_5596 (I97315,I97406,I221212);
nand I_5597 (I97686,I97508,I221206);
DFFARX1 I_5598 (I97686,I2507,I97341,I97330,);
DFFARX1 I_5599 (I97686,I2507,I97341,I97324,);
not I_5600 (I97731,I221206);
nor I_5601 (I97748,I97731,I221194);
and I_5602 (I97765,I97748,I221215);
or I_5603 (I97782,I97765,I221191);
DFFARX1 I_5604 (I97782,I2507,I97341,I97808,);
nand I_5605 (I97816,I97808,I97474);
nor I_5606 (I97318,I97816,I97624);
nor I_5607 (I97312,I97808,I97440);
DFFARX1 I_5608 (I97808,I2507,I97341,I97870,);
not I_5609 (I97878,I97870);
nor I_5610 (I97327,I97878,I97590);
not I_5611 (I97936,I2514);
DFFARX1 I_5612 (I682112,I2507,I97936,I97962,);
DFFARX1 I_5613 (I97962,I2507,I97936,I97979,);
not I_5614 (I97928,I97979);
not I_5615 (I98001,I97962);
DFFARX1 I_5616 (I682124,I2507,I97936,I98027,);
not I_5617 (I98035,I98027);
and I_5618 (I98052,I98001,I682118);
not I_5619 (I98069,I682130);
nand I_5620 (I98086,I98069,I682118);
not I_5621 (I98103,I682115);
nor I_5622 (I98120,I98103,I682127);
nand I_5623 (I98137,I98120,I682109);
nor I_5624 (I98154,I98137,I98086);
DFFARX1 I_5625 (I98154,I2507,I97936,I97904,);
not I_5626 (I98185,I98137);
not I_5627 (I98202,I682127);
nand I_5628 (I98219,I98202,I682118);
nor I_5629 (I98236,I682127,I682130);
nand I_5630 (I97916,I98052,I98236);
nand I_5631 (I97910,I98001,I682127);
nand I_5632 (I98281,I98103,I682121);
DFFARX1 I_5633 (I98281,I2507,I97936,I97925,);
DFFARX1 I_5634 (I98281,I2507,I97936,I97919,);
not I_5635 (I98326,I682121);
nor I_5636 (I98343,I98326,I682112);
and I_5637 (I98360,I98343,I682109);
or I_5638 (I98377,I98360,I682133);
DFFARX1 I_5639 (I98377,I2507,I97936,I98403,);
nand I_5640 (I98411,I98403,I98069);
nor I_5641 (I97913,I98411,I98219);
nor I_5642 (I97907,I98403,I98035);
DFFARX1 I_5643 (I98403,I2507,I97936,I98465,);
not I_5644 (I98473,I98465);
nor I_5645 (I97922,I98473,I98185);
not I_5646 (I98531,I2514);
DFFARX1 I_5647 (I472913,I2507,I98531,I98557,);
DFFARX1 I_5648 (I98557,I2507,I98531,I98574,);
not I_5649 (I98523,I98574);
not I_5650 (I98596,I98557);
DFFARX1 I_5651 (I472907,I2507,I98531,I98622,);
not I_5652 (I98630,I98622);
and I_5653 (I98647,I98596,I472925);
not I_5654 (I98664,I472913);
nand I_5655 (I98681,I98664,I472925);
not I_5656 (I98698,I472907);
nor I_5657 (I98715,I98698,I472919);
nand I_5658 (I98732,I98715,I472910);
nor I_5659 (I98749,I98732,I98681);
DFFARX1 I_5660 (I98749,I2507,I98531,I98499,);
not I_5661 (I98780,I98732);
not I_5662 (I98797,I472919);
nand I_5663 (I98814,I98797,I472925);
nor I_5664 (I98831,I472919,I472913);
nand I_5665 (I98511,I98647,I98831);
nand I_5666 (I98505,I98596,I472919);
nand I_5667 (I98876,I98698,I472922);
DFFARX1 I_5668 (I98876,I2507,I98531,I98520,);
DFFARX1 I_5669 (I98876,I2507,I98531,I98514,);
not I_5670 (I98921,I472922);
nor I_5671 (I98938,I98921,I472928);
and I_5672 (I98955,I98938,I472910);
or I_5673 (I98972,I98955,I472916);
DFFARX1 I_5674 (I98972,I2507,I98531,I98998,);
nand I_5675 (I99006,I98998,I98664);
nor I_5676 (I98508,I99006,I98814);
nor I_5677 (I98502,I98998,I98630);
DFFARX1 I_5678 (I98998,I2507,I98531,I99060,);
not I_5679 (I99068,I99060);
nor I_5680 (I98517,I99068,I98780);
not I_5681 (I99126,I2514);
DFFARX1 I_5682 (I618495,I2507,I99126,I99152,);
DFFARX1 I_5683 (I99152,I2507,I99126,I99169,);
not I_5684 (I99118,I99169);
not I_5685 (I99191,I99152);
DFFARX1 I_5686 (I618495,I2507,I99126,I99217,);
not I_5687 (I99225,I99217);
and I_5688 (I99242,I99191,I618498);
not I_5689 (I99259,I618510);
nand I_5690 (I99276,I99259,I618498);
not I_5691 (I99293,I618516);
nor I_5692 (I99310,I99293,I618507);
nand I_5693 (I99327,I99310,I618513);
nor I_5694 (I99344,I99327,I99276);
DFFARX1 I_5695 (I99344,I2507,I99126,I99094,);
not I_5696 (I99375,I99327);
not I_5697 (I99392,I618507);
nand I_5698 (I99409,I99392,I618498);
nor I_5699 (I99426,I618507,I618510);
nand I_5700 (I99106,I99242,I99426);
nand I_5701 (I99100,I99191,I618507);
nand I_5702 (I99471,I99293,I618504);
DFFARX1 I_5703 (I99471,I2507,I99126,I99115,);
DFFARX1 I_5704 (I99471,I2507,I99126,I99109,);
not I_5705 (I99516,I618504);
nor I_5706 (I99533,I99516,I618501);
and I_5707 (I99550,I99533,I618519);
or I_5708 (I99567,I99550,I618498);
DFFARX1 I_5709 (I99567,I2507,I99126,I99593,);
nand I_5710 (I99601,I99593,I99259);
nor I_5711 (I99103,I99601,I99409);
nor I_5712 (I99097,I99593,I99225);
DFFARX1 I_5713 (I99593,I2507,I99126,I99655,);
not I_5714 (I99663,I99655);
nor I_5715 (I99112,I99663,I99375);
not I_5716 (I99721,I2514);
DFFARX1 I_5717 (I562670,I2507,I99721,I99747,);
DFFARX1 I_5718 (I99747,I2507,I99721,I99764,);
not I_5719 (I99713,I99764);
not I_5720 (I99786,I99747);
DFFARX1 I_5721 (I562679,I2507,I99721,I99812,);
not I_5722 (I99820,I99812);
and I_5723 (I99837,I99786,I562673);
not I_5724 (I99854,I562667);
nand I_5725 (I99871,I99854,I562673);
not I_5726 (I99888,I562682);
nor I_5727 (I99905,I99888,I562670);
nand I_5728 (I99922,I99905,I562676);
nor I_5729 (I99939,I99922,I99871);
DFFARX1 I_5730 (I99939,I2507,I99721,I99689,);
not I_5731 (I99970,I99922);
not I_5732 (I99987,I562670);
nand I_5733 (I100004,I99987,I562673);
nor I_5734 (I100021,I562670,I562667);
nand I_5735 (I99701,I99837,I100021);
nand I_5736 (I99695,I99786,I562670);
nand I_5737 (I100066,I99888,I562673);
DFFARX1 I_5738 (I100066,I2507,I99721,I99710,);
DFFARX1 I_5739 (I100066,I2507,I99721,I99704,);
not I_5740 (I100111,I562673);
nor I_5741 (I100128,I100111,I562688);
and I_5742 (I100145,I100128,I562685);
or I_5743 (I100162,I100145,I562667);
DFFARX1 I_5744 (I100162,I2507,I99721,I100188,);
nand I_5745 (I100196,I100188,I99854);
nor I_5746 (I99698,I100196,I100004);
nor I_5747 (I99692,I100188,I99820);
DFFARX1 I_5748 (I100188,I2507,I99721,I100250,);
not I_5749 (I100258,I100250);
nor I_5750 (I99707,I100258,I99970);
not I_5751 (I100316,I2514);
DFFARX1 I_5752 (I622541,I2507,I100316,I100342,);
DFFARX1 I_5753 (I100342,I2507,I100316,I100359,);
not I_5754 (I100308,I100359);
not I_5755 (I100381,I100342);
DFFARX1 I_5756 (I622541,I2507,I100316,I100407,);
not I_5757 (I100415,I100407);
and I_5758 (I100432,I100381,I622544);
not I_5759 (I100449,I622556);
nand I_5760 (I100466,I100449,I622544);
not I_5761 (I100483,I622562);
nor I_5762 (I100500,I100483,I622553);
nand I_5763 (I100517,I100500,I622559);
nor I_5764 (I100534,I100517,I100466);
DFFARX1 I_5765 (I100534,I2507,I100316,I100284,);
not I_5766 (I100565,I100517);
not I_5767 (I100582,I622553);
nand I_5768 (I100599,I100582,I622544);
nor I_5769 (I100616,I622553,I622556);
nand I_5770 (I100296,I100432,I100616);
nand I_5771 (I100290,I100381,I622553);
nand I_5772 (I100661,I100483,I622550);
DFFARX1 I_5773 (I100661,I2507,I100316,I100305,);
DFFARX1 I_5774 (I100661,I2507,I100316,I100299,);
not I_5775 (I100706,I622550);
nor I_5776 (I100723,I100706,I622547);
and I_5777 (I100740,I100723,I622565);
or I_5778 (I100757,I100740,I622544);
DFFARX1 I_5779 (I100757,I2507,I100316,I100783,);
nand I_5780 (I100791,I100783,I100449);
nor I_5781 (I100293,I100791,I100599);
nor I_5782 (I100287,I100783,I100415);
DFFARX1 I_5783 (I100783,I2507,I100316,I100845,);
not I_5784 (I100853,I100845);
nor I_5785 (I100302,I100853,I100565);
not I_5786 (I100911,I2514);
DFFARX1 I_5787 (I444455,I2507,I100911,I100937,);
DFFARX1 I_5788 (I100937,I2507,I100911,I100954,);
not I_5789 (I100903,I100954);
not I_5790 (I100976,I100937);
DFFARX1 I_5791 (I444449,I2507,I100911,I101002,);
not I_5792 (I101010,I101002);
and I_5793 (I101027,I100976,I444467);
not I_5794 (I101044,I444455);
nand I_5795 (I101061,I101044,I444467);
not I_5796 (I101078,I444449);
nor I_5797 (I101095,I101078,I444461);
nand I_5798 (I101112,I101095,I444452);
nor I_5799 (I101129,I101112,I101061);
DFFARX1 I_5800 (I101129,I2507,I100911,I100879,);
not I_5801 (I101160,I101112);
not I_5802 (I101177,I444461);
nand I_5803 (I101194,I101177,I444467);
nor I_5804 (I101211,I444461,I444455);
nand I_5805 (I100891,I101027,I101211);
nand I_5806 (I100885,I100976,I444461);
nand I_5807 (I101256,I101078,I444464);
DFFARX1 I_5808 (I101256,I2507,I100911,I100900,);
DFFARX1 I_5809 (I101256,I2507,I100911,I100894,);
not I_5810 (I101301,I444464);
nor I_5811 (I101318,I101301,I444470);
and I_5812 (I101335,I101318,I444452);
or I_5813 (I101352,I101335,I444458);
DFFARX1 I_5814 (I101352,I2507,I100911,I101378,);
nand I_5815 (I101386,I101378,I101044);
nor I_5816 (I100888,I101386,I101194);
nor I_5817 (I100882,I101378,I101010);
DFFARX1 I_5818 (I101378,I2507,I100911,I101440,);
not I_5819 (I101448,I101440);
nor I_5820 (I100897,I101448,I101160);
not I_5821 (I101506,I2514);
DFFARX1 I_5822 (I572255,I2507,I101506,I101532,);
DFFARX1 I_5823 (I101532,I2507,I101506,I101549,);
not I_5824 (I101498,I101549);
not I_5825 (I101571,I101532);
DFFARX1 I_5826 (I572255,I2507,I101506,I101597,);
not I_5827 (I101605,I101597);
and I_5828 (I101622,I101571,I572258);
not I_5829 (I101639,I572270);
nand I_5830 (I101656,I101639,I572258);
not I_5831 (I101673,I572276);
nor I_5832 (I101690,I101673,I572267);
nand I_5833 (I101707,I101690,I572273);
nor I_5834 (I101724,I101707,I101656);
DFFARX1 I_5835 (I101724,I2507,I101506,I101474,);
not I_5836 (I101755,I101707);
not I_5837 (I101772,I572267);
nand I_5838 (I101789,I101772,I572258);
nor I_5839 (I101806,I572267,I572270);
nand I_5840 (I101486,I101622,I101806);
nand I_5841 (I101480,I101571,I572267);
nand I_5842 (I101851,I101673,I572264);
DFFARX1 I_5843 (I101851,I2507,I101506,I101495,);
DFFARX1 I_5844 (I101851,I2507,I101506,I101489,);
not I_5845 (I101896,I572264);
nor I_5846 (I101913,I101896,I572261);
and I_5847 (I101930,I101913,I572279);
or I_5848 (I101947,I101930,I572258);
DFFARX1 I_5849 (I101947,I2507,I101506,I101973,);
nand I_5850 (I101981,I101973,I101639);
nor I_5851 (I101483,I101981,I101789);
nor I_5852 (I101477,I101973,I101605);
DFFARX1 I_5853 (I101973,I2507,I101506,I102035,);
not I_5854 (I102043,I102035);
nor I_5855 (I101492,I102043,I101755);
not I_5856 (I102101,I2514);
DFFARX1 I_5857 (I720414,I2507,I102101,I102127,);
DFFARX1 I_5858 (I102127,I2507,I102101,I102144,);
not I_5859 (I102093,I102144);
not I_5860 (I102166,I102127);
DFFARX1 I_5861 (I720405,I2507,I102101,I102192,);
not I_5862 (I102200,I102192);
and I_5863 (I102217,I102166,I720399);
not I_5864 (I102234,I720393);
nand I_5865 (I102251,I102234,I720399);
not I_5866 (I102268,I720420);
nor I_5867 (I102285,I102268,I720393);
nand I_5868 (I102302,I102285,I720417);
nor I_5869 (I102319,I102302,I102251);
DFFARX1 I_5870 (I102319,I2507,I102101,I102069,);
not I_5871 (I102350,I102302);
not I_5872 (I102367,I720393);
nand I_5873 (I102384,I102367,I720399);
nor I_5874 (I102401,I720393,I720393);
nand I_5875 (I102081,I102217,I102401);
nand I_5876 (I102075,I102166,I720393);
nand I_5877 (I102446,I102268,I720402);
DFFARX1 I_5878 (I102446,I2507,I102101,I102090,);
DFFARX1 I_5879 (I102446,I2507,I102101,I102084,);
not I_5880 (I102491,I720402);
nor I_5881 (I102508,I102491,I720408);
and I_5882 (I102525,I102508,I720411);
or I_5883 (I102542,I102525,I720396);
DFFARX1 I_5884 (I102542,I2507,I102101,I102568,);
nand I_5885 (I102576,I102568,I102234);
nor I_5886 (I102078,I102576,I102384);
nor I_5887 (I102072,I102568,I102200);
DFFARX1 I_5888 (I102568,I2507,I102101,I102630,);
not I_5889 (I102638,I102630);
nor I_5890 (I102087,I102638,I102350);
not I_5891 (I102696,I2514);
DFFARX1 I_5892 (I39365,I2507,I102696,I102722,);
DFFARX1 I_5893 (I102722,I2507,I102696,I102739,);
not I_5894 (I102688,I102739);
not I_5895 (I102761,I102722);
DFFARX1 I_5896 (I39359,I2507,I102696,I102787,);
not I_5897 (I102795,I102787);
and I_5898 (I102812,I102761,I39356);
not I_5899 (I102829,I39377);
nand I_5900 (I102846,I102829,I39356);
not I_5901 (I102863,I39371);
nor I_5902 (I102880,I102863,I39362);
nand I_5903 (I102897,I102880,I39368);
nor I_5904 (I102914,I102897,I102846);
DFFARX1 I_5905 (I102914,I2507,I102696,I102664,);
not I_5906 (I102945,I102897);
not I_5907 (I102962,I39362);
nand I_5908 (I102979,I102962,I39356);
nor I_5909 (I102996,I39362,I39377);
nand I_5910 (I102676,I102812,I102996);
nand I_5911 (I102670,I102761,I39362);
nand I_5912 (I103041,I102863,I39356);
DFFARX1 I_5913 (I103041,I2507,I102696,I102685,);
DFFARX1 I_5914 (I103041,I2507,I102696,I102679,);
not I_5915 (I103086,I39356);
nor I_5916 (I103103,I103086,I39374);
and I_5917 (I103120,I103103,I39380);
or I_5918 (I103137,I103120,I39359);
DFFARX1 I_5919 (I103137,I2507,I102696,I103163,);
nand I_5920 (I103171,I103163,I102829);
nor I_5921 (I102673,I103171,I102979);
nor I_5922 (I102667,I103163,I102795);
DFFARX1 I_5923 (I103163,I2507,I102696,I103225,);
not I_5924 (I103233,I103225);
nor I_5925 (I102682,I103233,I102945);
not I_5926 (I103291,I2514);
DFFARX1 I_5927 (I494461,I2507,I103291,I103317,);
DFFARX1 I_5928 (I103317,I2507,I103291,I103334,);
not I_5929 (I103283,I103334);
not I_5930 (I103356,I103317);
DFFARX1 I_5931 (I494470,I2507,I103291,I103382,);
not I_5932 (I103390,I103382);
and I_5933 (I103407,I103356,I494458);
not I_5934 (I103424,I494449);
nand I_5935 (I103441,I103424,I494458);
not I_5936 (I103458,I494455);
nor I_5937 (I103475,I103458,I494473);
nand I_5938 (I103492,I103475,I494446);
nor I_5939 (I103509,I103492,I103441);
DFFARX1 I_5940 (I103509,I2507,I103291,I103259,);
not I_5941 (I103540,I103492);
not I_5942 (I103557,I494473);
nand I_5943 (I103574,I103557,I494458);
nor I_5944 (I103591,I494473,I494449);
nand I_5945 (I103271,I103407,I103591);
nand I_5946 (I103265,I103356,I494473);
nand I_5947 (I103636,I103458,I494452);
DFFARX1 I_5948 (I103636,I2507,I103291,I103280,);
DFFARX1 I_5949 (I103636,I2507,I103291,I103274,);
not I_5950 (I103681,I494452);
nor I_5951 (I103698,I103681,I494464);
and I_5952 (I103715,I103698,I494446);
or I_5953 (I103732,I103715,I494467);
DFFARX1 I_5954 (I103732,I2507,I103291,I103758,);
nand I_5955 (I103766,I103758,I103424);
nor I_5956 (I103268,I103766,I103574);
nor I_5957 (I103262,I103758,I103390);
DFFARX1 I_5958 (I103758,I2507,I103291,I103820,);
not I_5959 (I103828,I103820);
nor I_5960 (I103277,I103828,I103540);
not I_5961 (I103886,I2514);
DFFARX1 I_5962 (I479603,I2507,I103886,I103912,);
DFFARX1 I_5963 (I103912,I2507,I103886,I103929,);
not I_5964 (I103878,I103929);
not I_5965 (I103951,I103912);
DFFARX1 I_5966 (I479612,I2507,I103886,I103977,);
not I_5967 (I103985,I103977);
and I_5968 (I104002,I103951,I479600);
not I_5969 (I104019,I479591);
nand I_5970 (I104036,I104019,I479600);
not I_5971 (I104053,I479597);
nor I_5972 (I104070,I104053,I479615);
nand I_5973 (I104087,I104070,I479588);
nor I_5974 (I104104,I104087,I104036);
DFFARX1 I_5975 (I104104,I2507,I103886,I103854,);
not I_5976 (I104135,I104087);
not I_5977 (I104152,I479615);
nand I_5978 (I104169,I104152,I479600);
nor I_5979 (I104186,I479615,I479591);
nand I_5980 (I103866,I104002,I104186);
nand I_5981 (I103860,I103951,I479615);
nand I_5982 (I104231,I104053,I479594);
DFFARX1 I_5983 (I104231,I2507,I103886,I103875,);
DFFARX1 I_5984 (I104231,I2507,I103886,I103869,);
not I_5985 (I104276,I479594);
nor I_5986 (I104293,I104276,I479606);
and I_5987 (I104310,I104293,I479588);
or I_5988 (I104327,I104310,I479609);
DFFARX1 I_5989 (I104327,I2507,I103886,I104353,);
nand I_5990 (I104361,I104353,I104019);
nor I_5991 (I103863,I104361,I104169);
nor I_5992 (I103857,I104353,I103985);
DFFARX1 I_5993 (I104353,I2507,I103886,I104415,);
not I_5994 (I104423,I104415);
nor I_5995 (I103872,I104423,I104135);
not I_5996 (I104481,I2514);
DFFARX1 I_5997 (I218553,I2507,I104481,I104507,);
DFFARX1 I_5998 (I104507,I2507,I104481,I104524,);
not I_5999 (I104473,I104524);
not I_6000 (I104546,I104507);
DFFARX1 I_6001 (I218568,I2507,I104481,I104572,);
not I_6002 (I104580,I104572);
and I_6003 (I104597,I104546,I218565);
not I_6004 (I104614,I218553);
nand I_6005 (I104631,I104614,I218565);
not I_6006 (I104648,I218562);
nor I_6007 (I104665,I104648,I218577);
nand I_6008 (I104682,I104665,I218574);
nor I_6009 (I104699,I104682,I104631);
DFFARX1 I_6010 (I104699,I2507,I104481,I104449,);
not I_6011 (I104730,I104682);
not I_6012 (I104747,I218577);
nand I_6013 (I104764,I104747,I218565);
nor I_6014 (I104781,I218577,I218553);
nand I_6015 (I104461,I104597,I104781);
nand I_6016 (I104455,I104546,I218577);
nand I_6017 (I104826,I104648,I218571);
DFFARX1 I_6018 (I104826,I2507,I104481,I104470,);
DFFARX1 I_6019 (I104826,I2507,I104481,I104464,);
not I_6020 (I104871,I218571);
nor I_6021 (I104888,I104871,I218559);
and I_6022 (I104905,I104888,I218580);
or I_6023 (I104922,I104905,I218556);
DFFARX1 I_6024 (I104922,I2507,I104481,I104948,);
nand I_6025 (I104956,I104948,I104614);
nor I_6026 (I104458,I104956,I104764);
nor I_6027 (I104452,I104948,I104580);
DFFARX1 I_6028 (I104948,I2507,I104481,I105010,);
not I_6029 (I105018,I105010);
nor I_6030 (I104467,I105018,I104730);
not I_6031 (I105076,I2514);
DFFARX1 I_6032 (I295065,I2507,I105076,I105102,);
DFFARX1 I_6033 (I105102,I2507,I105076,I105119,);
not I_6034 (I105068,I105119);
not I_6035 (I105141,I105102);
DFFARX1 I_6036 (I295059,I2507,I105076,I105167,);
not I_6037 (I105175,I105167);
and I_6038 (I105192,I105141,I295074);
not I_6039 (I105209,I295071);
nand I_6040 (I105226,I105209,I295074);
not I_6041 (I105243,I295062);
nor I_6042 (I105260,I105243,I295053);
nand I_6043 (I105277,I105260,I295056);
nor I_6044 (I105294,I105277,I105226);
DFFARX1 I_6045 (I105294,I2507,I105076,I105044,);
not I_6046 (I105325,I105277);
not I_6047 (I105342,I295053);
nand I_6048 (I105359,I105342,I295074);
nor I_6049 (I105376,I295053,I295071);
nand I_6050 (I105056,I105192,I105376);
nand I_6051 (I105050,I105141,I295053);
nand I_6052 (I105421,I105243,I295077);
DFFARX1 I_6053 (I105421,I2507,I105076,I105065,);
DFFARX1 I_6054 (I105421,I2507,I105076,I105059,);
not I_6055 (I105466,I295077);
nor I_6056 (I105483,I105466,I295068);
and I_6057 (I105500,I105483,I295053);
or I_6058 (I105517,I105500,I295056);
DFFARX1 I_6059 (I105517,I2507,I105076,I105543,);
nand I_6060 (I105551,I105543,I105209);
nor I_6061 (I105053,I105551,I105359);
nor I_6062 (I105047,I105543,I105175);
DFFARX1 I_6063 (I105543,I2507,I105076,I105605,);
not I_6064 (I105613,I105605);
nor I_6065 (I105062,I105613,I105325);
not I_6066 (I105671,I2514);
DFFARX1 I_6067 (I233520,I2507,I105671,I105697,);
DFFARX1 I_6068 (I105697,I2507,I105671,I105714,);
not I_6069 (I105663,I105714);
not I_6070 (I105736,I105697);
DFFARX1 I_6071 (I233508,I2507,I105671,I105762,);
not I_6072 (I105770,I105762);
and I_6073 (I105787,I105736,I233517);
not I_6074 (I105804,I233514);
nand I_6075 (I105821,I105804,I233517);
not I_6076 (I105838,I233505);
nor I_6077 (I105855,I105838,I233511);
nand I_6078 (I105872,I105855,I233496);
nor I_6079 (I105889,I105872,I105821);
DFFARX1 I_6080 (I105889,I2507,I105671,I105639,);
not I_6081 (I105920,I105872);
not I_6082 (I105937,I233511);
nand I_6083 (I105954,I105937,I233517);
nor I_6084 (I105971,I233511,I233514);
nand I_6085 (I105651,I105787,I105971);
nand I_6086 (I105645,I105736,I233511);
nand I_6087 (I106016,I105838,I233496);
DFFARX1 I_6088 (I106016,I2507,I105671,I105660,);
DFFARX1 I_6089 (I106016,I2507,I105671,I105654,);
not I_6090 (I106061,I233496);
nor I_6091 (I106078,I106061,I233502);
and I_6092 (I106095,I106078,I233499);
or I_6093 (I106112,I106095,I233523);
DFFARX1 I_6094 (I106112,I2507,I105671,I106138,);
nand I_6095 (I106146,I106138,I105804);
nor I_6096 (I105648,I106146,I105954);
nor I_6097 (I105642,I106138,I105770);
DFFARX1 I_6098 (I106138,I2507,I105671,I106200,);
not I_6099 (I106208,I106200);
nor I_6100 (I105657,I106208,I105920);
not I_6101 (I106266,I2514);
DFFARX1 I_6102 (I438658,I2507,I106266,I106292,);
DFFARX1 I_6103 (I106292,I2507,I106266,I106309,);
not I_6104 (I106258,I106309);
not I_6105 (I106331,I106292);
DFFARX1 I_6106 (I438652,I2507,I106266,I106357,);
not I_6107 (I106365,I106357);
and I_6108 (I106382,I106331,I438670);
not I_6109 (I106399,I438658);
nand I_6110 (I106416,I106399,I438670);
not I_6111 (I106433,I438652);
nor I_6112 (I106450,I106433,I438664);
nand I_6113 (I106467,I106450,I438655);
nor I_6114 (I106484,I106467,I106416);
DFFARX1 I_6115 (I106484,I2507,I106266,I106234,);
not I_6116 (I106515,I106467);
not I_6117 (I106532,I438664);
nand I_6118 (I106549,I106532,I438670);
nor I_6119 (I106566,I438664,I438658);
nand I_6120 (I106246,I106382,I106566);
nand I_6121 (I106240,I106331,I438664);
nand I_6122 (I106611,I106433,I438667);
DFFARX1 I_6123 (I106611,I2507,I106266,I106255,);
DFFARX1 I_6124 (I106611,I2507,I106266,I106249,);
not I_6125 (I106656,I438667);
nor I_6126 (I106673,I106656,I438673);
and I_6127 (I106690,I106673,I438655);
or I_6128 (I106707,I106690,I438661);
DFFARX1 I_6129 (I106707,I2507,I106266,I106733,);
nand I_6130 (I106741,I106733,I106399);
nor I_6131 (I106243,I106741,I106549);
nor I_6132 (I106237,I106733,I106365);
DFFARX1 I_6133 (I106733,I2507,I106266,I106795,);
not I_6134 (I106803,I106795);
nor I_6135 (I106252,I106803,I106515);
not I_6136 (I106861,I2514);
DFFARX1 I_6137 (I355925,I2507,I106861,I106887,);
DFFARX1 I_6138 (I106887,I2507,I106861,I106904,);
not I_6139 (I106853,I106904);
not I_6140 (I106926,I106887);
DFFARX1 I_6141 (I355922,I2507,I106861,I106952,);
not I_6142 (I106960,I106952);
and I_6143 (I106977,I106926,I355928);
not I_6144 (I106994,I355913);
nand I_6145 (I107011,I106994,I355928);
not I_6146 (I107028,I355916);
nor I_6147 (I107045,I107028,I355937);
nand I_6148 (I107062,I107045,I355934);
nor I_6149 (I107079,I107062,I107011);
DFFARX1 I_6150 (I107079,I2507,I106861,I106829,);
not I_6151 (I107110,I107062);
not I_6152 (I107127,I355937);
nand I_6153 (I107144,I107127,I355928);
nor I_6154 (I107161,I355937,I355913);
nand I_6155 (I106841,I106977,I107161);
nand I_6156 (I106835,I106926,I355937);
nand I_6157 (I107206,I107028,I355913);
DFFARX1 I_6158 (I107206,I2507,I106861,I106850,);
DFFARX1 I_6159 (I107206,I2507,I106861,I106844,);
not I_6160 (I107251,I355913);
nor I_6161 (I107268,I107251,I355919);
and I_6162 (I107285,I107268,I355931);
or I_6163 (I107302,I107285,I355916);
DFFARX1 I_6164 (I107302,I2507,I106861,I107328,);
nand I_6165 (I107336,I107328,I106994);
nor I_6166 (I106838,I107336,I107144);
nor I_6167 (I106832,I107328,I106960);
DFFARX1 I_6168 (I107328,I2507,I106861,I107390,);
not I_6169 (I107398,I107390);
nor I_6170 (I106847,I107398,I107110);
not I_6171 (I107456,I2514);
DFFARX1 I_6172 (I530637,I2507,I107456,I107482,);
DFFARX1 I_6173 (I107482,I2507,I107456,I107499,);
not I_6174 (I107448,I107499);
not I_6175 (I107521,I107482);
DFFARX1 I_6176 (I530646,I2507,I107456,I107547,);
not I_6177 (I107555,I107547);
and I_6178 (I107572,I107521,I530634);
not I_6179 (I107589,I530625);
nand I_6180 (I107606,I107589,I530634);
not I_6181 (I107623,I530631);
nor I_6182 (I107640,I107623,I530649);
nand I_6183 (I107657,I107640,I530622);
nor I_6184 (I107674,I107657,I107606);
DFFARX1 I_6185 (I107674,I2507,I107456,I107424,);
not I_6186 (I107705,I107657);
not I_6187 (I107722,I530649);
nand I_6188 (I107739,I107722,I530634);
nor I_6189 (I107756,I530649,I530625);
nand I_6190 (I107436,I107572,I107756);
nand I_6191 (I107430,I107521,I530649);
nand I_6192 (I107801,I107623,I530628);
DFFARX1 I_6193 (I107801,I2507,I107456,I107445,);
DFFARX1 I_6194 (I107801,I2507,I107456,I107439,);
not I_6195 (I107846,I530628);
nor I_6196 (I107863,I107846,I530640);
and I_6197 (I107880,I107863,I530622);
or I_6198 (I107897,I107880,I530643);
DFFARX1 I_6199 (I107897,I2507,I107456,I107923,);
nand I_6200 (I107931,I107923,I107589);
nor I_6201 (I107433,I107931,I107739);
nor I_6202 (I107427,I107923,I107555);
DFFARX1 I_6203 (I107923,I2507,I107456,I107985,);
not I_6204 (I107993,I107985);
nor I_6205 (I107442,I107993,I107705);
not I_6206 (I108051,I2514);
DFFARX1 I_6207 (I652887,I2507,I108051,I108077,);
DFFARX1 I_6208 (I108077,I2507,I108051,I108094,);
not I_6209 (I108043,I108094);
not I_6210 (I108116,I108077);
DFFARX1 I_6211 (I652872,I2507,I108051,I108142,);
not I_6212 (I108150,I108142);
and I_6213 (I108167,I108116,I652890);
not I_6214 (I108184,I652872);
nand I_6215 (I108201,I108184,I652890);
not I_6216 (I108218,I652893);
nor I_6217 (I108235,I108218,I652884);
nand I_6218 (I108252,I108235,I652881);
nor I_6219 (I108269,I108252,I108201);
DFFARX1 I_6220 (I108269,I2507,I108051,I108019,);
not I_6221 (I108300,I108252);
not I_6222 (I108317,I652884);
nand I_6223 (I108334,I108317,I652890);
nor I_6224 (I108351,I652884,I652872);
nand I_6225 (I108031,I108167,I108351);
nand I_6226 (I108025,I108116,I652884);
nand I_6227 (I108396,I108218,I652878);
DFFARX1 I_6228 (I108396,I2507,I108051,I108040,);
DFFARX1 I_6229 (I108396,I2507,I108051,I108034,);
not I_6230 (I108441,I652878);
nor I_6231 (I108458,I108441,I652869);
and I_6232 (I108475,I108458,I652875);
or I_6233 (I108492,I108475,I652869);
DFFARX1 I_6234 (I108492,I2507,I108051,I108518,);
nand I_6235 (I108526,I108518,I108184);
nor I_6236 (I108028,I108526,I108334);
nor I_6237 (I108022,I108518,I108150);
DFFARX1 I_6238 (I108518,I2507,I108051,I108580,);
not I_6239 (I108588,I108580);
nor I_6240 (I108037,I108588,I108300);
not I_6241 (I108646,I2514);
DFFARX1 I_6242 (I578613,I2507,I108646,I108672,);
DFFARX1 I_6243 (I108672,I2507,I108646,I108689,);
not I_6244 (I108638,I108689);
not I_6245 (I108711,I108672);
DFFARX1 I_6246 (I578613,I2507,I108646,I108737,);
not I_6247 (I108745,I108737);
and I_6248 (I108762,I108711,I578616);
not I_6249 (I108779,I578628);
nand I_6250 (I108796,I108779,I578616);
not I_6251 (I108813,I578634);
nor I_6252 (I108830,I108813,I578625);
nand I_6253 (I108847,I108830,I578631);
nor I_6254 (I108864,I108847,I108796);
DFFARX1 I_6255 (I108864,I2507,I108646,I108614,);
not I_6256 (I108895,I108847);
not I_6257 (I108912,I578625);
nand I_6258 (I108929,I108912,I578616);
nor I_6259 (I108946,I578625,I578628);
nand I_6260 (I108626,I108762,I108946);
nand I_6261 (I108620,I108711,I578625);
nand I_6262 (I108991,I108813,I578622);
DFFARX1 I_6263 (I108991,I2507,I108646,I108635,);
DFFARX1 I_6264 (I108991,I2507,I108646,I108629,);
not I_6265 (I109036,I578622);
nor I_6266 (I109053,I109036,I578619);
and I_6267 (I109070,I109053,I578637);
or I_6268 (I109087,I109070,I578616);
DFFARX1 I_6269 (I109087,I2507,I108646,I109113,);
nand I_6270 (I109121,I109113,I108779);
nor I_6271 (I108623,I109121,I108929);
nor I_6272 (I108617,I109113,I108745);
DFFARX1 I_6273 (I109113,I2507,I108646,I109175,);
not I_6274 (I109183,I109175);
nor I_6275 (I108632,I109183,I108895);
not I_6276 (I109241,I2514);
DFFARX1 I_6277 (I514487,I2507,I109241,I109267,);
DFFARX1 I_6278 (I109267,I2507,I109241,I109284,);
not I_6279 (I109233,I109284);
not I_6280 (I109306,I109267);
DFFARX1 I_6281 (I514496,I2507,I109241,I109332,);
not I_6282 (I109340,I109332);
and I_6283 (I109357,I109306,I514484);
not I_6284 (I109374,I514475);
nand I_6285 (I109391,I109374,I514484);
not I_6286 (I109408,I514481);
nor I_6287 (I109425,I109408,I514499);
nand I_6288 (I109442,I109425,I514472);
nor I_6289 (I109459,I109442,I109391);
DFFARX1 I_6290 (I109459,I2507,I109241,I109209,);
not I_6291 (I109490,I109442);
not I_6292 (I109507,I514499);
nand I_6293 (I109524,I109507,I514484);
nor I_6294 (I109541,I514499,I514475);
nand I_6295 (I109221,I109357,I109541);
nand I_6296 (I109215,I109306,I514499);
nand I_6297 (I109586,I109408,I514478);
DFFARX1 I_6298 (I109586,I2507,I109241,I109230,);
DFFARX1 I_6299 (I109586,I2507,I109241,I109224,);
not I_6300 (I109631,I514478);
nor I_6301 (I109648,I109631,I514490);
and I_6302 (I109665,I109648,I514472);
or I_6303 (I109682,I109665,I514493);
DFFARX1 I_6304 (I109682,I2507,I109241,I109708,);
nand I_6305 (I109716,I109708,I109374);
nor I_6306 (I109218,I109716,I109524);
nor I_6307 (I109212,I109708,I109340);
DFFARX1 I_6308 (I109708,I2507,I109241,I109770,);
not I_6309 (I109778,I109770);
nor I_6310 (I109227,I109778,I109490);
not I_6311 (I109836,I2514);
DFFARX1 I_6312 (I712084,I2507,I109836,I109862,);
DFFARX1 I_6313 (I109862,I2507,I109836,I109879,);
not I_6314 (I109828,I109879);
not I_6315 (I109901,I109862);
DFFARX1 I_6316 (I712075,I2507,I109836,I109927,);
not I_6317 (I109935,I109927);
and I_6318 (I109952,I109901,I712069);
not I_6319 (I109969,I712063);
nand I_6320 (I109986,I109969,I712069);
not I_6321 (I110003,I712090);
nor I_6322 (I110020,I110003,I712063);
nand I_6323 (I110037,I110020,I712087);
nor I_6324 (I110054,I110037,I109986);
DFFARX1 I_6325 (I110054,I2507,I109836,I109804,);
not I_6326 (I110085,I110037);
not I_6327 (I110102,I712063);
nand I_6328 (I110119,I110102,I712069);
nor I_6329 (I110136,I712063,I712063);
nand I_6330 (I109816,I109952,I110136);
nand I_6331 (I109810,I109901,I712063);
nand I_6332 (I110181,I110003,I712072);
DFFARX1 I_6333 (I110181,I2507,I109836,I109825,);
DFFARX1 I_6334 (I110181,I2507,I109836,I109819,);
not I_6335 (I110226,I712072);
nor I_6336 (I110243,I110226,I712078);
and I_6337 (I110260,I110243,I712081);
or I_6338 (I110277,I110260,I712066);
DFFARX1 I_6339 (I110277,I2507,I109836,I110303,);
nand I_6340 (I110311,I110303,I109969);
nor I_6341 (I109813,I110311,I110119);
nor I_6342 (I109807,I110303,I109935);
DFFARX1 I_6343 (I110303,I2507,I109836,I110365,);
not I_6344 (I110373,I110365);
nor I_6345 (I109822,I110373,I110085);
not I_6346 (I110431,I2514);
DFFARX1 I_6347 (I599421,I2507,I110431,I110457,);
DFFARX1 I_6348 (I110457,I2507,I110431,I110474,);
not I_6349 (I110423,I110474);
not I_6350 (I110496,I110457);
DFFARX1 I_6351 (I599421,I2507,I110431,I110522,);
not I_6352 (I110530,I110522);
and I_6353 (I110547,I110496,I599424);
not I_6354 (I110564,I599436);
nand I_6355 (I110581,I110564,I599424);
not I_6356 (I110598,I599442);
nor I_6357 (I110615,I110598,I599433);
nand I_6358 (I110632,I110615,I599439);
nor I_6359 (I110649,I110632,I110581);
DFFARX1 I_6360 (I110649,I2507,I110431,I110399,);
not I_6361 (I110680,I110632);
not I_6362 (I110697,I599433);
nand I_6363 (I110714,I110697,I599424);
nor I_6364 (I110731,I599433,I599436);
nand I_6365 (I110411,I110547,I110731);
nand I_6366 (I110405,I110496,I599433);
nand I_6367 (I110776,I110598,I599430);
DFFARX1 I_6368 (I110776,I2507,I110431,I110420,);
DFFARX1 I_6369 (I110776,I2507,I110431,I110414,);
not I_6370 (I110821,I599430);
nor I_6371 (I110838,I110821,I599427);
and I_6372 (I110855,I110838,I599445);
or I_6373 (I110872,I110855,I599424);
DFFARX1 I_6374 (I110872,I2507,I110431,I110898,);
nand I_6375 (I110906,I110898,I110564);
nor I_6376 (I110408,I110906,I110714);
nor I_6377 (I110402,I110898,I110530);
DFFARX1 I_6378 (I110898,I2507,I110431,I110960,);
not I_6379 (I110968,I110960);
nor I_6380 (I110417,I110968,I110680);
not I_6381 (I111026,I2514);
DFFARX1 I_6382 (I217499,I2507,I111026,I111052,);
DFFARX1 I_6383 (I111052,I2507,I111026,I111069,);
not I_6384 (I111018,I111069);
not I_6385 (I111091,I111052);
DFFARX1 I_6386 (I217514,I2507,I111026,I111117,);
not I_6387 (I111125,I111117);
and I_6388 (I111142,I111091,I217511);
not I_6389 (I111159,I217499);
nand I_6390 (I111176,I111159,I217511);
not I_6391 (I111193,I217508);
nor I_6392 (I111210,I111193,I217523);
nand I_6393 (I111227,I111210,I217520);
nor I_6394 (I111244,I111227,I111176);
DFFARX1 I_6395 (I111244,I2507,I111026,I110994,);
not I_6396 (I111275,I111227);
not I_6397 (I111292,I217523);
nand I_6398 (I111309,I111292,I217511);
nor I_6399 (I111326,I217523,I217499);
nand I_6400 (I111006,I111142,I111326);
nand I_6401 (I111000,I111091,I217523);
nand I_6402 (I111371,I111193,I217517);
DFFARX1 I_6403 (I111371,I2507,I111026,I111015,);
DFFARX1 I_6404 (I111371,I2507,I111026,I111009,);
not I_6405 (I111416,I217517);
nor I_6406 (I111433,I111416,I217505);
and I_6407 (I111450,I111433,I217526);
or I_6408 (I111467,I111450,I217502);
DFFARX1 I_6409 (I111467,I2507,I111026,I111493,);
nand I_6410 (I111501,I111493,I111159);
nor I_6411 (I111003,I111501,I111309);
nor I_6412 (I110997,I111493,I111125);
DFFARX1 I_6413 (I111493,I2507,I111026,I111555,);
not I_6414 (I111563,I111555);
nor I_6415 (I111012,I111563,I111275);
not I_6416 (I111621,I2514);
DFFARX1 I_6417 (I72039,I2507,I111621,I111647,);
DFFARX1 I_6418 (I111647,I2507,I111621,I111664,);
not I_6419 (I111613,I111664);
not I_6420 (I111686,I111647);
DFFARX1 I_6421 (I72033,I2507,I111621,I111712,);
not I_6422 (I111720,I111712);
and I_6423 (I111737,I111686,I72030);
not I_6424 (I111754,I72051);
nand I_6425 (I111771,I111754,I72030);
not I_6426 (I111788,I72045);
nor I_6427 (I111805,I111788,I72036);
nand I_6428 (I111822,I111805,I72042);
nor I_6429 (I111839,I111822,I111771);
DFFARX1 I_6430 (I111839,I2507,I111621,I111589,);
not I_6431 (I111870,I111822);
not I_6432 (I111887,I72036);
nand I_6433 (I111904,I111887,I72030);
nor I_6434 (I111921,I72036,I72051);
nand I_6435 (I111601,I111737,I111921);
nand I_6436 (I111595,I111686,I72036);
nand I_6437 (I111966,I111788,I72030);
DFFARX1 I_6438 (I111966,I2507,I111621,I111610,);
DFFARX1 I_6439 (I111966,I2507,I111621,I111604,);
not I_6440 (I112011,I72030);
nor I_6441 (I112028,I112011,I72048);
and I_6442 (I112045,I112028,I72054);
or I_6443 (I112062,I112045,I72033);
DFFARX1 I_6444 (I112062,I2507,I111621,I112088,);
nand I_6445 (I112096,I112088,I111754);
nor I_6446 (I111598,I112096,I111904);
nor I_6447 (I111592,I112088,I111720);
DFFARX1 I_6448 (I112088,I2507,I111621,I112150,);
not I_6449 (I112158,I112150);
nor I_6450 (I111607,I112158,I111870);
not I_6451 (I112216,I2514);
DFFARX1 I_6452 (I277040,I2507,I112216,I112242,);
DFFARX1 I_6453 (I112242,I2507,I112216,I112259,);
not I_6454 (I112208,I112259);
not I_6455 (I112281,I112242);
DFFARX1 I_6456 (I277028,I2507,I112216,I112307,);
not I_6457 (I112315,I112307);
and I_6458 (I112332,I112281,I277037);
not I_6459 (I112349,I277034);
nand I_6460 (I112366,I112349,I277037);
not I_6461 (I112383,I277025);
nor I_6462 (I112400,I112383,I277031);
nand I_6463 (I112417,I112400,I277016);
nor I_6464 (I112434,I112417,I112366);
DFFARX1 I_6465 (I112434,I2507,I112216,I112184,);
not I_6466 (I112465,I112417);
not I_6467 (I112482,I277031);
nand I_6468 (I112499,I112482,I277037);
nor I_6469 (I112516,I277031,I277034);
nand I_6470 (I112196,I112332,I112516);
nand I_6471 (I112190,I112281,I277031);
nand I_6472 (I112561,I112383,I277016);
DFFARX1 I_6473 (I112561,I2507,I112216,I112205,);
DFFARX1 I_6474 (I112561,I2507,I112216,I112199,);
not I_6475 (I112606,I277016);
nor I_6476 (I112623,I112606,I277022);
and I_6477 (I112640,I112623,I277019);
or I_6478 (I112657,I112640,I277043);
DFFARX1 I_6479 (I112657,I2507,I112216,I112683,);
nand I_6480 (I112691,I112683,I112349);
nor I_6481 (I112193,I112691,I112499);
nor I_6482 (I112187,I112683,I112315);
DFFARX1 I_6483 (I112683,I2507,I112216,I112745,);
not I_6484 (I112753,I112745);
nor I_6485 (I112202,I112753,I112465);
not I_6486 (I112811,I2514);
DFFARX1 I_6487 (I630633,I2507,I112811,I112837,);
DFFARX1 I_6488 (I112837,I2507,I112811,I112854,);
not I_6489 (I112803,I112854);
not I_6490 (I112876,I112837);
DFFARX1 I_6491 (I630633,I2507,I112811,I112902,);
not I_6492 (I112910,I112902);
and I_6493 (I112927,I112876,I630636);
not I_6494 (I112944,I630648);
nand I_6495 (I112961,I112944,I630636);
not I_6496 (I112978,I630654);
nor I_6497 (I112995,I112978,I630645);
nand I_6498 (I113012,I112995,I630651);
nor I_6499 (I113029,I113012,I112961);
DFFARX1 I_6500 (I113029,I2507,I112811,I112779,);
not I_6501 (I113060,I113012);
not I_6502 (I113077,I630645);
nand I_6503 (I113094,I113077,I630636);
nor I_6504 (I113111,I630645,I630648);
nand I_6505 (I112791,I112927,I113111);
nand I_6506 (I112785,I112876,I630645);
nand I_6507 (I113156,I112978,I630642);
DFFARX1 I_6508 (I113156,I2507,I112811,I112800,);
DFFARX1 I_6509 (I113156,I2507,I112811,I112794,);
not I_6510 (I113201,I630642);
nor I_6511 (I113218,I113201,I630639);
and I_6512 (I113235,I113218,I630657);
or I_6513 (I113252,I113235,I630636);
DFFARX1 I_6514 (I113252,I2507,I112811,I113278,);
nand I_6515 (I113286,I113278,I112944);
nor I_6516 (I112788,I113286,I113094);
nor I_6517 (I112782,I113278,I112910);
DFFARX1 I_6518 (I113278,I2507,I112811,I113340,);
not I_6519 (I113348,I113340);
nor I_6520 (I112797,I113348,I113060);
not I_6521 (I113406,I2514);
DFFARX1 I_6522 (I469751,I2507,I113406,I113432,);
DFFARX1 I_6523 (I113432,I2507,I113406,I113449,);
not I_6524 (I113398,I113449);
not I_6525 (I113471,I113432);
DFFARX1 I_6526 (I469745,I2507,I113406,I113497,);
not I_6527 (I113505,I113497);
and I_6528 (I113522,I113471,I469763);
not I_6529 (I113539,I469751);
nand I_6530 (I113556,I113539,I469763);
not I_6531 (I113573,I469745);
nor I_6532 (I113590,I113573,I469757);
nand I_6533 (I113607,I113590,I469748);
nor I_6534 (I113624,I113607,I113556);
DFFARX1 I_6535 (I113624,I2507,I113406,I113374,);
not I_6536 (I113655,I113607);
not I_6537 (I113672,I469757);
nand I_6538 (I113689,I113672,I469763);
nor I_6539 (I113706,I469757,I469751);
nand I_6540 (I113386,I113522,I113706);
nand I_6541 (I113380,I113471,I469757);
nand I_6542 (I113751,I113573,I469760);
DFFARX1 I_6543 (I113751,I2507,I113406,I113395,);
DFFARX1 I_6544 (I113751,I2507,I113406,I113389,);
not I_6545 (I113796,I469760);
nor I_6546 (I113813,I113796,I469766);
and I_6547 (I113830,I113813,I469748);
or I_6548 (I113847,I113830,I469754);
DFFARX1 I_6549 (I113847,I2507,I113406,I113873,);
nand I_6550 (I113881,I113873,I113539);
nor I_6551 (I113383,I113881,I113689);
nor I_6552 (I113377,I113873,I113505);
DFFARX1 I_6553 (I113873,I2507,I113406,I113935,);
not I_6554 (I113943,I113935);
nor I_6555 (I113392,I113943,I113655);
not I_6556 (I114001,I2514);
DFFARX1 I_6557 (I684992,I2507,I114001,I114027,);
DFFARX1 I_6558 (I114027,I2507,I114001,I114044,);
not I_6559 (I113993,I114044);
not I_6560 (I114066,I114027);
DFFARX1 I_6561 (I684965,I2507,I114001,I114092,);
not I_6562 (I114100,I114092);
and I_6563 (I114117,I114066,I684989);
not I_6564 (I114134,I684986);
nand I_6565 (I114151,I114134,I684989);
not I_6566 (I114168,I684965);
nor I_6567 (I114185,I114168,I684983);
nand I_6568 (I114202,I114185,I684971);
nor I_6569 (I114219,I114202,I114151);
DFFARX1 I_6570 (I114219,I2507,I114001,I113969,);
not I_6571 (I114250,I114202);
not I_6572 (I114267,I684983);
nand I_6573 (I114284,I114267,I684989);
nor I_6574 (I114301,I684983,I684986);
nand I_6575 (I113981,I114117,I114301);
nand I_6576 (I113975,I114066,I684983);
nand I_6577 (I114346,I114168,I684977);
DFFARX1 I_6578 (I114346,I2507,I114001,I113990,);
DFFARX1 I_6579 (I114346,I2507,I114001,I113984,);
not I_6580 (I114391,I684977);
nor I_6581 (I114408,I114391,I684980);
and I_6582 (I114425,I114408,I684968);
or I_6583 (I114442,I114425,I684974);
DFFARX1 I_6584 (I114442,I2507,I114001,I114468,);
nand I_6585 (I114476,I114468,I114134);
nor I_6586 (I113978,I114476,I114284);
nor I_6587 (I113972,I114468,I114100);
DFFARX1 I_6588 (I114468,I2507,I114001,I114530,);
not I_6589 (I114538,I114530);
nor I_6590 (I113987,I114538,I114250);
not I_6591 (I114596,I2514);
DFFARX1 I_6592 (I347255,I2507,I114596,I114622,);
DFFARX1 I_6593 (I114622,I2507,I114596,I114639,);
not I_6594 (I114588,I114639);
not I_6595 (I114661,I114622);
DFFARX1 I_6596 (I347252,I2507,I114596,I114687,);
not I_6597 (I114695,I114687);
and I_6598 (I114712,I114661,I347258);
not I_6599 (I114729,I347243);
nand I_6600 (I114746,I114729,I347258);
not I_6601 (I114763,I347246);
nor I_6602 (I114780,I114763,I347267);
nand I_6603 (I114797,I114780,I347264);
nor I_6604 (I114814,I114797,I114746);
DFFARX1 I_6605 (I114814,I2507,I114596,I114564,);
not I_6606 (I114845,I114797);
not I_6607 (I114862,I347267);
nand I_6608 (I114879,I114862,I347258);
nor I_6609 (I114896,I347267,I347243);
nand I_6610 (I114576,I114712,I114896);
nand I_6611 (I114570,I114661,I347267);
nand I_6612 (I114941,I114763,I347243);
DFFARX1 I_6613 (I114941,I2507,I114596,I114585,);
DFFARX1 I_6614 (I114941,I2507,I114596,I114579,);
not I_6615 (I114986,I347243);
nor I_6616 (I115003,I114986,I347249);
and I_6617 (I115020,I115003,I347261);
or I_6618 (I115037,I115020,I347246);
DFFARX1 I_6619 (I115037,I2507,I114596,I115063,);
nand I_6620 (I115071,I115063,I114729);
nor I_6621 (I114573,I115071,I114879);
nor I_6622 (I114567,I115063,I114695);
DFFARX1 I_6623 (I115063,I2507,I114596,I115125,);
not I_6624 (I115133,I115125);
nor I_6625 (I114582,I115133,I114845);
not I_6626 (I115191,I2514);
DFFARX1 I_6627 (I300420,I2507,I115191,I115217,);
DFFARX1 I_6628 (I115217,I2507,I115191,I115234,);
not I_6629 (I115183,I115234);
not I_6630 (I115256,I115217);
DFFARX1 I_6631 (I300414,I2507,I115191,I115282,);
not I_6632 (I115290,I115282);
and I_6633 (I115307,I115256,I300429);
not I_6634 (I115324,I300426);
nand I_6635 (I115341,I115324,I300429);
not I_6636 (I115358,I300417);
nor I_6637 (I115375,I115358,I300408);
nand I_6638 (I115392,I115375,I300411);
nor I_6639 (I115409,I115392,I115341);
DFFARX1 I_6640 (I115409,I2507,I115191,I115159,);
not I_6641 (I115440,I115392);
not I_6642 (I115457,I300408);
nand I_6643 (I115474,I115457,I300429);
nor I_6644 (I115491,I300408,I300426);
nand I_6645 (I115171,I115307,I115491);
nand I_6646 (I115165,I115256,I300408);
nand I_6647 (I115536,I115358,I300432);
DFFARX1 I_6648 (I115536,I2507,I115191,I115180,);
DFFARX1 I_6649 (I115536,I2507,I115191,I115174,);
not I_6650 (I115581,I300432);
nor I_6651 (I115598,I115581,I300423);
and I_6652 (I115615,I115598,I300408);
or I_6653 (I115632,I115615,I300411);
DFFARX1 I_6654 (I115632,I2507,I115191,I115658,);
nand I_6655 (I115666,I115658,I115324);
nor I_6656 (I115168,I115666,I115474);
nor I_6657 (I115162,I115658,I115290);
DFFARX1 I_6658 (I115658,I2507,I115191,I115720,);
not I_6659 (I115728,I115720);
nor I_6660 (I115177,I115728,I115440);
not I_6661 (I115786,I2514);
DFFARX1 I_6662 (I369219,I2507,I115786,I115812,);
DFFARX1 I_6663 (I115812,I2507,I115786,I115829,);
not I_6664 (I115778,I115829);
not I_6665 (I115851,I115812);
DFFARX1 I_6666 (I369216,I2507,I115786,I115877,);
not I_6667 (I115885,I115877);
and I_6668 (I115902,I115851,I369222);
not I_6669 (I115919,I369207);
nand I_6670 (I115936,I115919,I369222);
not I_6671 (I115953,I369210);
nor I_6672 (I115970,I115953,I369231);
nand I_6673 (I115987,I115970,I369228);
nor I_6674 (I116004,I115987,I115936);
DFFARX1 I_6675 (I116004,I2507,I115786,I115754,);
not I_6676 (I116035,I115987);
not I_6677 (I116052,I369231);
nand I_6678 (I116069,I116052,I369222);
nor I_6679 (I116086,I369231,I369207);
nand I_6680 (I115766,I115902,I116086);
nand I_6681 (I115760,I115851,I369231);
nand I_6682 (I116131,I115953,I369207);
DFFARX1 I_6683 (I116131,I2507,I115786,I115775,);
DFFARX1 I_6684 (I116131,I2507,I115786,I115769,);
not I_6685 (I116176,I369207);
nor I_6686 (I116193,I116176,I369213);
and I_6687 (I116210,I116193,I369225);
or I_6688 (I116227,I116210,I369210);
DFFARX1 I_6689 (I116227,I2507,I115786,I116253,);
nand I_6690 (I116261,I116253,I115919);
nor I_6691 (I115763,I116261,I116069);
nor I_6692 (I115757,I116253,I115885);
DFFARX1 I_6693 (I116253,I2507,I115786,I116315,);
not I_6694 (I116323,I116315);
nor I_6695 (I115772,I116323,I116035);
not I_6696 (I116381,I2514);
DFFARX1 I_6697 (I675754,I2507,I116381,I116407,);
DFFARX1 I_6698 (I116407,I2507,I116381,I116424,);
not I_6699 (I116373,I116424);
not I_6700 (I116446,I116407);
DFFARX1 I_6701 (I675766,I2507,I116381,I116472,);
not I_6702 (I116480,I116472);
and I_6703 (I116497,I116446,I675760);
not I_6704 (I116514,I675772);
nand I_6705 (I116531,I116514,I675760);
not I_6706 (I116548,I675757);
nor I_6707 (I116565,I116548,I675769);
nand I_6708 (I116582,I116565,I675751);
nor I_6709 (I116599,I116582,I116531);
DFFARX1 I_6710 (I116599,I2507,I116381,I116349,);
not I_6711 (I116630,I116582);
not I_6712 (I116647,I675769);
nand I_6713 (I116664,I116647,I675760);
nor I_6714 (I116681,I675769,I675772);
nand I_6715 (I116361,I116497,I116681);
nand I_6716 (I116355,I116446,I675769);
nand I_6717 (I116726,I116548,I675763);
DFFARX1 I_6718 (I116726,I2507,I116381,I116370,);
DFFARX1 I_6719 (I116726,I2507,I116381,I116364,);
not I_6720 (I116771,I675763);
nor I_6721 (I116788,I116771,I675754);
and I_6722 (I116805,I116788,I675751);
or I_6723 (I116822,I116805,I675775);
DFFARX1 I_6724 (I116822,I2507,I116381,I116848,);
nand I_6725 (I116856,I116848,I116514);
nor I_6726 (I116358,I116856,I116664);
nor I_6727 (I116352,I116848,I116480);
DFFARX1 I_6728 (I116848,I2507,I116381,I116910,);
not I_6729 (I116918,I116910);
nor I_6730 (I116367,I116918,I116630);
not I_6731 (I116976,I2514);
DFFARX1 I_6732 (I576879,I2507,I116976,I117002,);
DFFARX1 I_6733 (I117002,I2507,I116976,I117019,);
not I_6734 (I116968,I117019);
not I_6735 (I117041,I117002);
DFFARX1 I_6736 (I576879,I2507,I116976,I117067,);
not I_6737 (I117075,I117067);
and I_6738 (I117092,I117041,I576882);
not I_6739 (I117109,I576894);
nand I_6740 (I117126,I117109,I576882);
not I_6741 (I117143,I576900);
nor I_6742 (I117160,I117143,I576891);
nand I_6743 (I117177,I117160,I576897);
nor I_6744 (I117194,I117177,I117126);
DFFARX1 I_6745 (I117194,I2507,I116976,I116944,);
not I_6746 (I117225,I117177);
not I_6747 (I117242,I576891);
nand I_6748 (I117259,I117242,I576882);
nor I_6749 (I117276,I576891,I576894);
nand I_6750 (I116956,I117092,I117276);
nand I_6751 (I116950,I117041,I576891);
nand I_6752 (I117321,I117143,I576888);
DFFARX1 I_6753 (I117321,I2507,I116976,I116965,);
DFFARX1 I_6754 (I117321,I2507,I116976,I116959,);
not I_6755 (I117366,I576888);
nor I_6756 (I117383,I117366,I576885);
and I_6757 (I117400,I117383,I576903);
or I_6758 (I117417,I117400,I576882);
DFFARX1 I_6759 (I117417,I2507,I116976,I117443,);
nand I_6760 (I117451,I117443,I117109);
nor I_6761 (I116953,I117451,I117259);
nor I_6762 (I116947,I117443,I117075);
DFFARX1 I_6763 (I117443,I2507,I116976,I117505,);
not I_6764 (I117513,I117505);
nor I_6765 (I116962,I117513,I117225);
not I_6766 (I117571,I2514);
DFFARX1 I_6767 (I353613,I2507,I117571,I117597,);
DFFARX1 I_6768 (I117597,I2507,I117571,I117614,);
not I_6769 (I117563,I117614);
not I_6770 (I117636,I117597);
DFFARX1 I_6771 (I353610,I2507,I117571,I117662,);
not I_6772 (I117670,I117662);
and I_6773 (I117687,I117636,I353616);
not I_6774 (I117704,I353601);
nand I_6775 (I117721,I117704,I353616);
not I_6776 (I117738,I353604);
nor I_6777 (I117755,I117738,I353625);
nand I_6778 (I117772,I117755,I353622);
nor I_6779 (I117789,I117772,I117721);
DFFARX1 I_6780 (I117789,I2507,I117571,I117539,);
not I_6781 (I117820,I117772);
not I_6782 (I117837,I353625);
nand I_6783 (I117854,I117837,I353616);
nor I_6784 (I117871,I353625,I353601);
nand I_6785 (I117551,I117687,I117871);
nand I_6786 (I117545,I117636,I353625);
nand I_6787 (I117916,I117738,I353601);
DFFARX1 I_6788 (I117916,I2507,I117571,I117560,);
DFFARX1 I_6789 (I117916,I2507,I117571,I117554,);
not I_6790 (I117961,I353601);
nor I_6791 (I117978,I117961,I353607);
and I_6792 (I117995,I117978,I353619);
or I_6793 (I118012,I117995,I353604);
DFFARX1 I_6794 (I118012,I2507,I117571,I118038,);
nand I_6795 (I118046,I118038,I117704);
nor I_6796 (I117548,I118046,I117854);
nor I_6797 (I117542,I118038,I117670);
DFFARX1 I_6798 (I118038,I2507,I117571,I118100,);
not I_6799 (I118108,I118100);
nor I_6800 (I117557,I118108,I117820);
not I_6801 (I118166,I2514);
DFFARX1 I_6802 (I65715,I2507,I118166,I118192,);
DFFARX1 I_6803 (I118192,I2507,I118166,I118209,);
not I_6804 (I118158,I118209);
not I_6805 (I118231,I118192);
DFFARX1 I_6806 (I65709,I2507,I118166,I118257,);
not I_6807 (I118265,I118257);
and I_6808 (I118282,I118231,I65706);
not I_6809 (I118299,I65727);
nand I_6810 (I118316,I118299,I65706);
not I_6811 (I118333,I65721);
nor I_6812 (I118350,I118333,I65712);
nand I_6813 (I118367,I118350,I65718);
nor I_6814 (I118384,I118367,I118316);
DFFARX1 I_6815 (I118384,I2507,I118166,I118134,);
not I_6816 (I118415,I118367);
not I_6817 (I118432,I65712);
nand I_6818 (I118449,I118432,I65706);
nor I_6819 (I118466,I65712,I65727);
nand I_6820 (I118146,I118282,I118466);
nand I_6821 (I118140,I118231,I65712);
nand I_6822 (I118511,I118333,I65706);
DFFARX1 I_6823 (I118511,I2507,I118166,I118155,);
DFFARX1 I_6824 (I118511,I2507,I118166,I118149,);
not I_6825 (I118556,I65706);
nor I_6826 (I118573,I118556,I65724);
and I_6827 (I118590,I118573,I65730);
or I_6828 (I118607,I118590,I65709);
DFFARX1 I_6829 (I118607,I2507,I118166,I118633,);
nand I_6830 (I118641,I118633,I118299);
nor I_6831 (I118143,I118641,I118449);
nor I_6832 (I118137,I118633,I118265);
DFFARX1 I_6833 (I118633,I2507,I118166,I118695,);
not I_6834 (I118703,I118695);
nor I_6835 (I118152,I118703,I118415);
not I_6836 (I118761,I2514);
DFFARX1 I_6837 (I548645,I2507,I118761,I118787,);
DFFARX1 I_6838 (I118787,I2507,I118761,I118804,);
not I_6839 (I118753,I118804);
not I_6840 (I118826,I118787);
DFFARX1 I_6841 (I548654,I2507,I118761,I118852,);
not I_6842 (I118860,I118852);
and I_6843 (I118877,I118826,I548648);
not I_6844 (I118894,I548642);
nand I_6845 (I118911,I118894,I548648);
not I_6846 (I118928,I548657);
nor I_6847 (I118945,I118928,I548645);
nand I_6848 (I118962,I118945,I548651);
nor I_6849 (I118979,I118962,I118911);
DFFARX1 I_6850 (I118979,I2507,I118761,I118729,);
not I_6851 (I119010,I118962);
not I_6852 (I119027,I548645);
nand I_6853 (I119044,I119027,I548648);
nor I_6854 (I119061,I548645,I548642);
nand I_6855 (I118741,I118877,I119061);
nand I_6856 (I118735,I118826,I548645);
nand I_6857 (I119106,I118928,I548648);
DFFARX1 I_6858 (I119106,I2507,I118761,I118750,);
DFFARX1 I_6859 (I119106,I2507,I118761,I118744,);
not I_6860 (I119151,I548648);
nor I_6861 (I119168,I119151,I548663);
and I_6862 (I119185,I119168,I548660);
or I_6863 (I119202,I119185,I548642);
DFFARX1 I_6864 (I119202,I2507,I118761,I119228,);
nand I_6865 (I119236,I119228,I118894);
nor I_6866 (I118738,I119236,I119044);
nor I_6867 (I118732,I119228,I118860);
DFFARX1 I_6868 (I119228,I2507,I118761,I119290,);
not I_6869 (I119298,I119290);
nor I_6870 (I118747,I119298,I119010);
not I_6871 (I119356,I2514);
DFFARX1 I_6872 (I30948,I2507,I119356,I119382,);
DFFARX1 I_6873 (I119382,I2507,I119356,I119399,);
not I_6874 (I119348,I119399);
not I_6875 (I119421,I119382);
DFFARX1 I_6876 (I30924,I2507,I119356,I119447,);
not I_6877 (I119455,I119447);
and I_6878 (I119472,I119421,I30939);
not I_6879 (I119489,I30927);
nand I_6880 (I119506,I119489,I30939);
not I_6881 (I119523,I30930);
nor I_6882 (I119540,I119523,I30942);
nand I_6883 (I119557,I119540,I30933);
nor I_6884 (I119574,I119557,I119506);
DFFARX1 I_6885 (I119574,I2507,I119356,I119324,);
not I_6886 (I119605,I119557);
not I_6887 (I119622,I30942);
nand I_6888 (I119639,I119622,I30939);
nor I_6889 (I119656,I30942,I30927);
nand I_6890 (I119336,I119472,I119656);
nand I_6891 (I119330,I119421,I30942);
nand I_6892 (I119701,I119523,I30936);
DFFARX1 I_6893 (I119701,I2507,I119356,I119345,);
DFFARX1 I_6894 (I119701,I2507,I119356,I119339,);
not I_6895 (I119746,I30936);
nor I_6896 (I119763,I119746,I30927);
and I_6897 (I119780,I119763,I30924);
or I_6898 (I119797,I119780,I30945);
DFFARX1 I_6899 (I119797,I2507,I119356,I119823,);
nand I_6900 (I119831,I119823,I119489);
nor I_6901 (I119333,I119831,I119639);
nor I_6902 (I119327,I119823,I119455);
DFFARX1 I_6903 (I119823,I2507,I119356,I119885,);
not I_6904 (I119893,I119885);
nor I_6905 (I119342,I119893,I119605);
not I_6906 (I119951,I2514);
DFFARX1 I_6907 (I252016,I2507,I119951,I119977,);
DFFARX1 I_6908 (I119977,I2507,I119951,I119994,);
not I_6909 (I119943,I119994);
not I_6910 (I120016,I119977);
DFFARX1 I_6911 (I252004,I2507,I119951,I120042,);
not I_6912 (I120050,I120042);
and I_6913 (I120067,I120016,I252013);
not I_6914 (I120084,I252010);
nand I_6915 (I120101,I120084,I252013);
not I_6916 (I120118,I252001);
nor I_6917 (I120135,I120118,I252007);
nand I_6918 (I120152,I120135,I251992);
nor I_6919 (I120169,I120152,I120101);
DFFARX1 I_6920 (I120169,I2507,I119951,I119919,);
not I_6921 (I120200,I120152);
not I_6922 (I120217,I252007);
nand I_6923 (I120234,I120217,I252013);
nor I_6924 (I120251,I252007,I252010);
nand I_6925 (I119931,I120067,I120251);
nand I_6926 (I119925,I120016,I252007);
nand I_6927 (I120296,I120118,I251992);
DFFARX1 I_6928 (I120296,I2507,I119951,I119940,);
DFFARX1 I_6929 (I120296,I2507,I119951,I119934,);
not I_6930 (I120341,I251992);
nor I_6931 (I120358,I120341,I251998);
and I_6932 (I120375,I120358,I251995);
or I_6933 (I120392,I120375,I252019);
DFFARX1 I_6934 (I120392,I2507,I119951,I120418,);
nand I_6935 (I120426,I120418,I120084);
nor I_6936 (I119928,I120426,I120234);
nor I_6937 (I119922,I120418,I120050);
DFFARX1 I_6938 (I120418,I2507,I119951,I120480,);
not I_6939 (I120488,I120480);
nor I_6940 (I119937,I120488,I120200);
not I_6941 (I120546,I2514);
DFFARX1 I_6942 (I638147,I2507,I120546,I120572,);
DFFARX1 I_6943 (I120572,I2507,I120546,I120589,);
not I_6944 (I120538,I120589);
not I_6945 (I120611,I120572);
DFFARX1 I_6946 (I638147,I2507,I120546,I120637,);
not I_6947 (I120645,I120637);
and I_6948 (I120662,I120611,I638150);
not I_6949 (I120679,I638162);
nand I_6950 (I120696,I120679,I638150);
not I_6951 (I120713,I638168);
nor I_6952 (I120730,I120713,I638159);
nand I_6953 (I120747,I120730,I638165);
nor I_6954 (I120764,I120747,I120696);
DFFARX1 I_6955 (I120764,I2507,I120546,I120514,);
not I_6956 (I120795,I120747);
not I_6957 (I120812,I638159);
nand I_6958 (I120829,I120812,I638150);
nor I_6959 (I120846,I638159,I638162);
nand I_6960 (I120526,I120662,I120846);
nand I_6961 (I120520,I120611,I638159);
nand I_6962 (I120891,I120713,I638156);
DFFARX1 I_6963 (I120891,I2507,I120546,I120535,);
DFFARX1 I_6964 (I120891,I2507,I120546,I120529,);
not I_6965 (I120936,I638156);
nor I_6966 (I120953,I120936,I638153);
and I_6967 (I120970,I120953,I638171);
or I_6968 (I120987,I120970,I638150);
DFFARX1 I_6969 (I120987,I2507,I120546,I121013,);
nand I_6970 (I121021,I121013,I120679);
nor I_6971 (I120523,I121021,I120829);
nor I_6972 (I120517,I121013,I120645);
DFFARX1 I_6973 (I121013,I2507,I120546,I121075,);
not I_6974 (I121083,I121075);
nor I_6975 (I120532,I121083,I120795);
not I_6976 (I121141,I2514);
DFFARX1 I_6977 (I595375,I2507,I121141,I121167,);
DFFARX1 I_6978 (I121167,I2507,I121141,I121184,);
not I_6979 (I121133,I121184);
not I_6980 (I121206,I121167);
DFFARX1 I_6981 (I595375,I2507,I121141,I121232,);
not I_6982 (I121240,I121232);
and I_6983 (I121257,I121206,I595378);
not I_6984 (I121274,I595390);
nand I_6985 (I121291,I121274,I595378);
not I_6986 (I121308,I595396);
nor I_6987 (I121325,I121308,I595387);
nand I_6988 (I121342,I121325,I595393);
nor I_6989 (I121359,I121342,I121291);
DFFARX1 I_6990 (I121359,I2507,I121141,I121109,);
not I_6991 (I121390,I121342);
not I_6992 (I121407,I595387);
nand I_6993 (I121424,I121407,I595378);
nor I_6994 (I121441,I595387,I595390);
nand I_6995 (I121121,I121257,I121441);
nand I_6996 (I121115,I121206,I595387);
nand I_6997 (I121486,I121308,I595384);
DFFARX1 I_6998 (I121486,I2507,I121141,I121130,);
DFFARX1 I_6999 (I121486,I2507,I121141,I121124,);
not I_7000 (I121531,I595384);
nor I_7001 (I121548,I121531,I595381);
and I_7002 (I121565,I121548,I595399);
or I_7003 (I121582,I121565,I595378);
DFFARX1 I_7004 (I121582,I2507,I121141,I121608,);
nand I_7005 (I121616,I121608,I121274);
nor I_7006 (I121118,I121616,I121424);
nor I_7007 (I121112,I121608,I121240);
DFFARX1 I_7008 (I121608,I2507,I121141,I121670,);
not I_7009 (I121678,I121670);
nor I_7010 (I121127,I121678,I121390);
not I_7011 (I121736,I2514);
DFFARX1 I_7012 (I631789,I2507,I121736,I121762,);
DFFARX1 I_7013 (I121762,I2507,I121736,I121779,);
not I_7014 (I121728,I121779);
not I_7015 (I121801,I121762);
DFFARX1 I_7016 (I631789,I2507,I121736,I121827,);
not I_7017 (I121835,I121827);
and I_7018 (I121852,I121801,I631792);
not I_7019 (I121869,I631804);
nand I_7020 (I121886,I121869,I631792);
not I_7021 (I121903,I631810);
nor I_7022 (I121920,I121903,I631801);
nand I_7023 (I121937,I121920,I631807);
nor I_7024 (I121954,I121937,I121886);
DFFARX1 I_7025 (I121954,I2507,I121736,I121704,);
not I_7026 (I121985,I121937);
not I_7027 (I122002,I631801);
nand I_7028 (I122019,I122002,I631792);
nor I_7029 (I122036,I631801,I631804);
nand I_7030 (I121716,I121852,I122036);
nand I_7031 (I121710,I121801,I631801);
nand I_7032 (I122081,I121903,I631798);
DFFARX1 I_7033 (I122081,I2507,I121736,I121725,);
DFFARX1 I_7034 (I122081,I2507,I121736,I121719,);
not I_7035 (I122126,I631798);
nor I_7036 (I122143,I122126,I631795);
and I_7037 (I122160,I122143,I631813);
or I_7038 (I122177,I122160,I631792);
DFFARX1 I_7039 (I122177,I2507,I121736,I122203,);
nand I_7040 (I122211,I122203,I121869);
nor I_7041 (I121713,I122211,I122019);
nor I_7042 (I121707,I122203,I121835);
DFFARX1 I_7043 (I122203,I2507,I121736,I122265,);
not I_7044 (I122273,I122265);
nor I_7045 (I121722,I122273,I121985);
not I_7046 (I122331,I2514);
DFFARX1 I_7047 (I476602,I2507,I122331,I122357,);
DFFARX1 I_7048 (I122357,I2507,I122331,I122374,);
not I_7049 (I122323,I122374);
not I_7050 (I122396,I122357);
DFFARX1 I_7051 (I476596,I2507,I122331,I122422,);
not I_7052 (I122430,I122422);
and I_7053 (I122447,I122396,I476614);
not I_7054 (I122464,I476602);
nand I_7055 (I122481,I122464,I476614);
not I_7056 (I122498,I476596);
nor I_7057 (I122515,I122498,I476608);
nand I_7058 (I122532,I122515,I476599);
nor I_7059 (I122549,I122532,I122481);
DFFARX1 I_7060 (I122549,I2507,I122331,I122299,);
not I_7061 (I122580,I122532);
not I_7062 (I122597,I476608);
nand I_7063 (I122614,I122597,I476614);
nor I_7064 (I122631,I476608,I476602);
nand I_7065 (I122311,I122447,I122631);
nand I_7066 (I122305,I122396,I476608);
nand I_7067 (I122676,I122498,I476611);
DFFARX1 I_7068 (I122676,I2507,I122331,I122320,);
DFFARX1 I_7069 (I122676,I2507,I122331,I122314,);
not I_7070 (I122721,I476611);
nor I_7071 (I122738,I122721,I476617);
and I_7072 (I122755,I122738,I476599);
or I_7073 (I122772,I122755,I476605);
DFFARX1 I_7074 (I122772,I2507,I122331,I122798,);
nand I_7075 (I122806,I122798,I122464);
nor I_7076 (I122308,I122806,I122614);
nor I_7077 (I122302,I122798,I122430);
DFFARX1 I_7078 (I122798,I2507,I122331,I122860,);
not I_7079 (I122868,I122860);
nor I_7080 (I122317,I122868,I122580);
not I_7081 (I122926,I2514);
DFFARX1 I_7082 (I634101,I2507,I122926,I122952,);
DFFARX1 I_7083 (I122952,I2507,I122926,I122969,);
not I_7084 (I122918,I122969);
not I_7085 (I122991,I122952);
DFFARX1 I_7086 (I634101,I2507,I122926,I123017,);
not I_7087 (I123025,I123017);
and I_7088 (I123042,I122991,I634104);
not I_7089 (I123059,I634116);
nand I_7090 (I123076,I123059,I634104);
not I_7091 (I123093,I634122);
nor I_7092 (I123110,I123093,I634113);
nand I_7093 (I123127,I123110,I634119);
nor I_7094 (I123144,I123127,I123076);
DFFARX1 I_7095 (I123144,I2507,I122926,I122894,);
not I_7096 (I123175,I123127);
not I_7097 (I123192,I634113);
nand I_7098 (I123209,I123192,I634104);
nor I_7099 (I123226,I634113,I634116);
nand I_7100 (I122906,I123042,I123226);
nand I_7101 (I122900,I122991,I634113);
nand I_7102 (I123271,I123093,I634110);
DFFARX1 I_7103 (I123271,I2507,I122926,I122915,);
DFFARX1 I_7104 (I123271,I2507,I122926,I122909,);
not I_7105 (I123316,I634110);
nor I_7106 (I123333,I123316,I634107);
and I_7107 (I123350,I123333,I634125);
or I_7108 (I123367,I123350,I634104);
DFFARX1 I_7109 (I123367,I2507,I122926,I123393,);
nand I_7110 (I123401,I123393,I123059);
nor I_7111 (I122903,I123401,I123209);
nor I_7112 (I122897,I123393,I123025);
DFFARX1 I_7113 (I123393,I2507,I122926,I123455,);
not I_7114 (I123463,I123455);
nor I_7115 (I122912,I123463,I123175);
not I_7116 (I123521,I2514);
DFFARX1 I_7117 (I440766,I2507,I123521,I123547,);
DFFARX1 I_7118 (I123547,I2507,I123521,I123564,);
not I_7119 (I123513,I123564);
not I_7120 (I123586,I123547);
DFFARX1 I_7121 (I440760,I2507,I123521,I123612,);
not I_7122 (I123620,I123612);
and I_7123 (I123637,I123586,I440778);
not I_7124 (I123654,I440766);
nand I_7125 (I123671,I123654,I440778);
not I_7126 (I123688,I440760);
nor I_7127 (I123705,I123688,I440772);
nand I_7128 (I123722,I123705,I440763);
nor I_7129 (I123739,I123722,I123671);
DFFARX1 I_7130 (I123739,I2507,I123521,I123489,);
not I_7131 (I123770,I123722);
not I_7132 (I123787,I440772);
nand I_7133 (I123804,I123787,I440778);
nor I_7134 (I123821,I440772,I440766);
nand I_7135 (I123501,I123637,I123821);
nand I_7136 (I123495,I123586,I440772);
nand I_7137 (I123866,I123688,I440775);
DFFARX1 I_7138 (I123866,I2507,I123521,I123510,);
DFFARX1 I_7139 (I123866,I2507,I123521,I123504,);
not I_7140 (I123911,I440775);
nor I_7141 (I123928,I123911,I440781);
and I_7142 (I123945,I123928,I440763);
or I_7143 (I123962,I123945,I440769);
DFFARX1 I_7144 (I123962,I2507,I123521,I123988,);
nand I_7145 (I123996,I123988,I123654);
nor I_7146 (I123498,I123996,I123804);
nor I_7147 (I123492,I123988,I123620);
DFFARX1 I_7148 (I123988,I2507,I123521,I124050,);
not I_7149 (I124058,I124050);
nor I_7150 (I123507,I124058,I123770);
not I_7151 (I124116,I2514);
DFFARX1 I_7152 (I620807,I2507,I124116,I124142,);
DFFARX1 I_7153 (I124142,I2507,I124116,I124159,);
not I_7154 (I124108,I124159);
not I_7155 (I124181,I124142);
DFFARX1 I_7156 (I620807,I2507,I124116,I124207,);
not I_7157 (I124215,I124207);
and I_7158 (I124232,I124181,I620810);
not I_7159 (I124249,I620822);
nand I_7160 (I124266,I124249,I620810);
not I_7161 (I124283,I620828);
nor I_7162 (I124300,I124283,I620819);
nand I_7163 (I124317,I124300,I620825);
nor I_7164 (I124334,I124317,I124266);
DFFARX1 I_7165 (I124334,I2507,I124116,I124084,);
not I_7166 (I124365,I124317);
not I_7167 (I124382,I620819);
nand I_7168 (I124399,I124382,I620810);
nor I_7169 (I124416,I620819,I620822);
nand I_7170 (I124096,I124232,I124416);
nand I_7171 (I124090,I124181,I620819);
nand I_7172 (I124461,I124283,I620816);
DFFARX1 I_7173 (I124461,I2507,I124116,I124105,);
DFFARX1 I_7174 (I124461,I2507,I124116,I124099,);
not I_7175 (I124506,I620816);
nor I_7176 (I124523,I124506,I620813);
and I_7177 (I124540,I124523,I620831);
or I_7178 (I124557,I124540,I620810);
DFFARX1 I_7179 (I124557,I2507,I124116,I124583,);
nand I_7180 (I124591,I124583,I124249);
nor I_7181 (I124093,I124591,I124399);
nor I_7182 (I124087,I124583,I124215);
DFFARX1 I_7183 (I124583,I2507,I124116,I124645,);
not I_7184 (I124653,I124645);
nor I_7185 (I124102,I124653,I124365);
not I_7186 (I124711,I2514);
DFFARX1 I_7187 (I75201,I2507,I124711,I124737,);
DFFARX1 I_7188 (I124737,I2507,I124711,I124754,);
not I_7189 (I124703,I124754);
not I_7190 (I124776,I124737);
DFFARX1 I_7191 (I75195,I2507,I124711,I124802,);
not I_7192 (I124810,I124802);
and I_7193 (I124827,I124776,I75192);
not I_7194 (I124844,I75213);
nand I_7195 (I124861,I124844,I75192);
not I_7196 (I124878,I75207);
nor I_7197 (I124895,I124878,I75198);
nand I_7198 (I124912,I124895,I75204);
nor I_7199 (I124929,I124912,I124861);
DFFARX1 I_7200 (I124929,I2507,I124711,I124679,);
not I_7201 (I124960,I124912);
not I_7202 (I124977,I75198);
nand I_7203 (I124994,I124977,I75192);
nor I_7204 (I125011,I75198,I75213);
nand I_7205 (I124691,I124827,I125011);
nand I_7206 (I124685,I124776,I75198);
nand I_7207 (I125056,I124878,I75192);
DFFARX1 I_7208 (I125056,I2507,I124711,I124700,);
DFFARX1 I_7209 (I125056,I2507,I124711,I124694,);
not I_7210 (I125101,I75192);
nor I_7211 (I125118,I125101,I75210);
and I_7212 (I125135,I125118,I75216);
or I_7213 (I125152,I125135,I75195);
DFFARX1 I_7214 (I125152,I2507,I124711,I125178,);
nand I_7215 (I125186,I125178,I124844);
nor I_7216 (I124688,I125186,I124994);
nor I_7217 (I124682,I125178,I124810);
DFFARX1 I_7218 (I125178,I2507,I124711,I125240,);
not I_7219 (I125248,I125240);
nor I_7220 (I124697,I125248,I124960);
not I_7221 (I125306,I2514);
DFFARX1 I_7222 (I515779,I2507,I125306,I125332,);
DFFARX1 I_7223 (I125332,I2507,I125306,I125349,);
not I_7224 (I125298,I125349);
not I_7225 (I125371,I125332);
DFFARX1 I_7226 (I515788,I2507,I125306,I125397,);
not I_7227 (I125405,I125397);
and I_7228 (I125422,I125371,I515776);
not I_7229 (I125439,I515767);
nand I_7230 (I125456,I125439,I515776);
not I_7231 (I125473,I515773);
nor I_7232 (I125490,I125473,I515791);
nand I_7233 (I125507,I125490,I515764);
nor I_7234 (I125524,I125507,I125456);
DFFARX1 I_7235 (I125524,I2507,I125306,I125274,);
not I_7236 (I125555,I125507);
not I_7237 (I125572,I515791);
nand I_7238 (I125589,I125572,I515776);
nor I_7239 (I125606,I515791,I515767);
nand I_7240 (I125286,I125422,I125606);
nand I_7241 (I125280,I125371,I515791);
nand I_7242 (I125651,I125473,I515770);
DFFARX1 I_7243 (I125651,I2507,I125306,I125295,);
DFFARX1 I_7244 (I125651,I2507,I125306,I125289,);
not I_7245 (I125696,I515770);
nor I_7246 (I125713,I125696,I515782);
and I_7247 (I125730,I125713,I515764);
or I_7248 (I125747,I125730,I515785);
DFFARX1 I_7249 (I125747,I2507,I125306,I125773,);
nand I_7250 (I125781,I125773,I125439);
nor I_7251 (I125283,I125781,I125589);
nor I_7252 (I125277,I125773,I125405);
DFFARX1 I_7253 (I125773,I2507,I125306,I125835,);
not I_7254 (I125843,I125835);
nor I_7255 (I125292,I125843,I125555);
not I_7256 (I125901,I2514);
DFFARX1 I_7257 (I17246,I2507,I125901,I125927,);
DFFARX1 I_7258 (I125927,I2507,I125901,I125944,);
not I_7259 (I125893,I125944);
not I_7260 (I125966,I125927);
DFFARX1 I_7261 (I17222,I2507,I125901,I125992,);
not I_7262 (I126000,I125992);
and I_7263 (I126017,I125966,I17237);
not I_7264 (I126034,I17225);
nand I_7265 (I126051,I126034,I17237);
not I_7266 (I126068,I17228);
nor I_7267 (I126085,I126068,I17240);
nand I_7268 (I126102,I126085,I17231);
nor I_7269 (I126119,I126102,I126051);
DFFARX1 I_7270 (I126119,I2507,I125901,I125869,);
not I_7271 (I126150,I126102);
not I_7272 (I126167,I17240);
nand I_7273 (I126184,I126167,I17237);
nor I_7274 (I126201,I17240,I17225);
nand I_7275 (I125881,I126017,I126201);
nand I_7276 (I125875,I125966,I17240);
nand I_7277 (I126246,I126068,I17234);
DFFARX1 I_7278 (I126246,I2507,I125901,I125890,);
DFFARX1 I_7279 (I126246,I2507,I125901,I125884,);
not I_7280 (I126291,I17234);
nor I_7281 (I126308,I126291,I17225);
and I_7282 (I126325,I126308,I17222);
or I_7283 (I126342,I126325,I17243);
DFFARX1 I_7284 (I126342,I2507,I125901,I126368,);
nand I_7285 (I126376,I126368,I126034);
nor I_7286 (I125878,I126376,I126184);
nor I_7287 (I125872,I126368,I126000);
DFFARX1 I_7288 (I126368,I2507,I125901,I126430,);
not I_7289 (I126438,I126430);
nor I_7290 (I125887,I126438,I126150);
not I_7291 (I126496,I2514);
DFFARX1 I_7292 (I595953,I2507,I126496,I126522,);
DFFARX1 I_7293 (I126522,I2507,I126496,I126539,);
not I_7294 (I126488,I126539);
not I_7295 (I126561,I126522);
DFFARX1 I_7296 (I595953,I2507,I126496,I126587,);
not I_7297 (I126595,I126587);
and I_7298 (I126612,I126561,I595956);
not I_7299 (I126629,I595968);
nand I_7300 (I126646,I126629,I595956);
not I_7301 (I126663,I595974);
nor I_7302 (I126680,I126663,I595965);
nand I_7303 (I126697,I126680,I595971);
nor I_7304 (I126714,I126697,I126646);
DFFARX1 I_7305 (I126714,I2507,I126496,I126464,);
not I_7306 (I126745,I126697);
not I_7307 (I126762,I595965);
nand I_7308 (I126779,I126762,I595956);
nor I_7309 (I126796,I595965,I595968);
nand I_7310 (I126476,I126612,I126796);
nand I_7311 (I126470,I126561,I595965);
nand I_7312 (I126841,I126663,I595962);
DFFARX1 I_7313 (I126841,I2507,I126496,I126485,);
DFFARX1 I_7314 (I126841,I2507,I126496,I126479,);
not I_7315 (I126886,I595962);
nor I_7316 (I126903,I126886,I595959);
and I_7317 (I126920,I126903,I595977);
or I_7318 (I126937,I126920,I595956);
DFFARX1 I_7319 (I126937,I2507,I126496,I126963,);
nand I_7320 (I126971,I126963,I126629);
nor I_7321 (I126473,I126971,I126779);
nor I_7322 (I126467,I126963,I126595);
DFFARX1 I_7323 (I126963,I2507,I126496,I127025,);
not I_7324 (I127033,I127025);
nor I_7325 (I126482,I127033,I126745);
not I_7326 (I127091,I2514);
DFFARX1 I_7327 (I34095,I2507,I127091,I127117,);
DFFARX1 I_7328 (I127117,I2507,I127091,I127134,);
not I_7329 (I127083,I127134);
not I_7330 (I127156,I127117);
DFFARX1 I_7331 (I34089,I2507,I127091,I127182,);
not I_7332 (I127190,I127182);
and I_7333 (I127207,I127156,I34086);
not I_7334 (I127224,I34107);
nand I_7335 (I127241,I127224,I34086);
not I_7336 (I127258,I34101);
nor I_7337 (I127275,I127258,I34092);
nand I_7338 (I127292,I127275,I34098);
nor I_7339 (I127309,I127292,I127241);
DFFARX1 I_7340 (I127309,I2507,I127091,I127059,);
not I_7341 (I127340,I127292);
not I_7342 (I127357,I34092);
nand I_7343 (I127374,I127357,I34086);
nor I_7344 (I127391,I34092,I34107);
nand I_7345 (I127071,I127207,I127391);
nand I_7346 (I127065,I127156,I34092);
nand I_7347 (I127436,I127258,I34086);
DFFARX1 I_7348 (I127436,I2507,I127091,I127080,);
DFFARX1 I_7349 (I127436,I2507,I127091,I127074,);
not I_7350 (I127481,I34086);
nor I_7351 (I127498,I127481,I34104);
and I_7352 (I127515,I127498,I34110);
or I_7353 (I127532,I127515,I34089);
DFFARX1 I_7354 (I127532,I2507,I127091,I127558,);
nand I_7355 (I127566,I127558,I127224);
nor I_7356 (I127068,I127566,I127374);
nor I_7357 (I127062,I127558,I127190);
DFFARX1 I_7358 (I127558,I2507,I127091,I127620,);
not I_7359 (I127628,I127620);
nor I_7360 (I127077,I127628,I127340);
not I_7361 (I127686,I2514);
DFFARX1 I_7362 (I593641,I2507,I127686,I127712,);
DFFARX1 I_7363 (I127712,I2507,I127686,I127729,);
not I_7364 (I127678,I127729);
not I_7365 (I127751,I127712);
DFFARX1 I_7366 (I593641,I2507,I127686,I127777,);
not I_7367 (I127785,I127777);
and I_7368 (I127802,I127751,I593644);
not I_7369 (I127819,I593656);
nand I_7370 (I127836,I127819,I593644);
not I_7371 (I127853,I593662);
nor I_7372 (I127870,I127853,I593653);
nand I_7373 (I127887,I127870,I593659);
nor I_7374 (I127904,I127887,I127836);
DFFARX1 I_7375 (I127904,I2507,I127686,I127654,);
not I_7376 (I127935,I127887);
not I_7377 (I127952,I593653);
nand I_7378 (I127969,I127952,I593644);
nor I_7379 (I127986,I593653,I593656);
nand I_7380 (I127666,I127802,I127986);
nand I_7381 (I127660,I127751,I593653);
nand I_7382 (I128031,I127853,I593650);
DFFARX1 I_7383 (I128031,I2507,I127686,I127675,);
DFFARX1 I_7384 (I128031,I2507,I127686,I127669,);
not I_7385 (I128076,I593650);
nor I_7386 (I128093,I128076,I593647);
and I_7387 (I128110,I128093,I593665);
or I_7388 (I128127,I128110,I593644);
DFFARX1 I_7389 (I128127,I2507,I127686,I128153,);
nand I_7390 (I128161,I128153,I127819);
nor I_7391 (I127663,I128161,I127969);
nor I_7392 (I127657,I128153,I127785);
DFFARX1 I_7393 (I128153,I2507,I127686,I128215,);
not I_7394 (I128223,I128215);
nor I_7395 (I127672,I128223,I127935);
not I_7396 (I128281,I2514);
DFFARX1 I_7397 (I597109,I2507,I128281,I128307,);
DFFARX1 I_7398 (I128307,I2507,I128281,I128324,);
not I_7399 (I128273,I128324);
not I_7400 (I128346,I128307);
DFFARX1 I_7401 (I597109,I2507,I128281,I128372,);
not I_7402 (I128380,I128372);
and I_7403 (I128397,I128346,I597112);
not I_7404 (I128414,I597124);
nand I_7405 (I128431,I128414,I597112);
not I_7406 (I128448,I597130);
nor I_7407 (I128465,I128448,I597121);
nand I_7408 (I128482,I128465,I597127);
nor I_7409 (I128499,I128482,I128431);
DFFARX1 I_7410 (I128499,I2507,I128281,I128249,);
not I_7411 (I128530,I128482);
not I_7412 (I128547,I597121);
nand I_7413 (I128564,I128547,I597112);
nor I_7414 (I128581,I597121,I597124);
nand I_7415 (I128261,I128397,I128581);
nand I_7416 (I128255,I128346,I597121);
nand I_7417 (I128626,I128448,I597118);
DFFARX1 I_7418 (I128626,I2507,I128281,I128270,);
DFFARX1 I_7419 (I128626,I2507,I128281,I128264,);
not I_7420 (I128671,I597118);
nor I_7421 (I128688,I128671,I597115);
and I_7422 (I128705,I128688,I597133);
or I_7423 (I128722,I128705,I597112);
DFFARX1 I_7424 (I128722,I2507,I128281,I128748,);
nand I_7425 (I128756,I128748,I128414);
nor I_7426 (I128258,I128756,I128564);
nor I_7427 (I128252,I128748,I128380);
DFFARX1 I_7428 (I128748,I2507,I128281,I128810,);
not I_7429 (I128818,I128810);
nor I_7430 (I128267,I128818,I128530);
not I_7431 (I128876,I2514);
DFFARX1 I_7432 (I305642,I2507,I128876,I128902,);
DFFARX1 I_7433 (I128902,I2507,I128876,I128919,);
not I_7434 (I128868,I128919);
not I_7435 (I128941,I128902);
DFFARX1 I_7436 (I305633,I2507,I128876,I128967,);
not I_7437 (I128975,I128967);
and I_7438 (I128992,I128941,I305651);
not I_7439 (I129009,I305648);
nand I_7440 (I129026,I129009,I305651);
not I_7441 (I129043,I305627);
nor I_7442 (I129060,I129043,I305630);
nand I_7443 (I129077,I129060,I305639);
nor I_7444 (I129094,I129077,I129026);
DFFARX1 I_7445 (I129094,I2507,I128876,I128844,);
not I_7446 (I129125,I129077);
not I_7447 (I129142,I305630);
nand I_7448 (I129159,I129142,I305651);
nor I_7449 (I129176,I305630,I305648);
nand I_7450 (I128856,I128992,I129176);
nand I_7451 (I128850,I128941,I305630);
nand I_7452 (I129221,I129043,I305645);
DFFARX1 I_7453 (I129221,I2507,I128876,I128865,);
DFFARX1 I_7454 (I129221,I2507,I128876,I128859,);
not I_7455 (I129266,I305645);
nor I_7456 (I129283,I129266,I305627);
and I_7457 (I129300,I129283,I305636);
or I_7458 (I129317,I129300,I305630);
DFFARX1 I_7459 (I129317,I2507,I128876,I129343,);
nand I_7460 (I129351,I129343,I129009);
nor I_7461 (I128853,I129351,I129159);
nor I_7462 (I128847,I129343,I128975);
DFFARX1 I_7463 (I129343,I2507,I128876,I129405,);
not I_7464 (I129413,I129405);
nor I_7465 (I128862,I129413,I129125);
not I_7466 (I129471,I2514);
DFFARX1 I_7467 (I411413,I2507,I129471,I129497,);
DFFARX1 I_7468 (I129497,I2507,I129471,I129514,);
not I_7469 (I129463,I129514);
not I_7470 (I129536,I129497);
DFFARX1 I_7471 (I411410,I2507,I129471,I129562,);
not I_7472 (I129570,I129562);
and I_7473 (I129587,I129536,I411416);
not I_7474 (I129604,I411401);
nand I_7475 (I129621,I129604,I411416);
not I_7476 (I129638,I411404);
nor I_7477 (I129655,I129638,I411425);
nand I_7478 (I129672,I129655,I411422);
nor I_7479 (I129689,I129672,I129621);
DFFARX1 I_7480 (I129689,I2507,I129471,I129439,);
not I_7481 (I129720,I129672);
not I_7482 (I129737,I411425);
nand I_7483 (I129754,I129737,I411416);
nor I_7484 (I129771,I411425,I411401);
nand I_7485 (I129451,I129587,I129771);
nand I_7486 (I129445,I129536,I411425);
nand I_7487 (I129816,I129638,I411401);
DFFARX1 I_7488 (I129816,I2507,I129471,I129460,);
DFFARX1 I_7489 (I129816,I2507,I129471,I129454,);
not I_7490 (I129861,I411401);
nor I_7491 (I129878,I129861,I411407);
and I_7492 (I129895,I129878,I411419);
or I_7493 (I129912,I129895,I411404);
DFFARX1 I_7494 (I129912,I2507,I129471,I129938,);
nand I_7495 (I129946,I129938,I129604);
nor I_7496 (I129448,I129946,I129754);
nor I_7497 (I129442,I129938,I129570);
DFFARX1 I_7498 (I129938,I2507,I129471,I130000,);
not I_7499 (I130008,I130000);
nor I_7500 (I129457,I130008,I129720);
not I_7501 (I130066,I2514);
DFFARX1 I_7502 (I87212,I2507,I130066,I130092,);
DFFARX1 I_7503 (I130092,I2507,I130066,I130109,);
not I_7504 (I130058,I130109);
not I_7505 (I130131,I130092);
DFFARX1 I_7506 (I87197,I2507,I130066,I130157,);
not I_7507 (I130165,I130157);
and I_7508 (I130182,I130131,I87218);
not I_7509 (I130199,I87209);
nand I_7510 (I130216,I130199,I87218);
not I_7511 (I130233,I87194);
nor I_7512 (I130250,I130233,I87206);
nand I_7513 (I130267,I130250,I87221);
nor I_7514 (I130284,I130267,I130216);
DFFARX1 I_7515 (I130284,I2507,I130066,I130034,);
not I_7516 (I130315,I130267);
not I_7517 (I130332,I87206);
nand I_7518 (I130349,I130332,I87218);
nor I_7519 (I130366,I87206,I87209);
nand I_7520 (I130046,I130182,I130366);
nand I_7521 (I130040,I130131,I87206);
nand I_7522 (I130411,I130233,I87200);
DFFARX1 I_7523 (I130411,I2507,I130066,I130055,);
DFFARX1 I_7524 (I130411,I2507,I130066,I130049,);
not I_7525 (I130456,I87200);
nor I_7526 (I130473,I130456,I87203);
and I_7527 (I130490,I130473,I87194);
or I_7528 (I130507,I130490,I87215);
DFFARX1 I_7529 (I130507,I2507,I130066,I130533,);
nand I_7530 (I130541,I130533,I130199);
nor I_7531 (I130043,I130541,I130349);
nor I_7532 (I130037,I130533,I130165);
DFFARX1 I_7533 (I130533,I2507,I130066,I130595,);
not I_7534 (I130603,I130595);
nor I_7535 (I130052,I130603,I130315);
not I_7536 (I130661,I2514);
DFFARX1 I_7537 (I309110,I2507,I130661,I130687,);
DFFARX1 I_7538 (I130687,I2507,I130661,I130704,);
not I_7539 (I130653,I130704);
not I_7540 (I130726,I130687);
DFFARX1 I_7541 (I309101,I2507,I130661,I130752,);
not I_7542 (I130760,I130752);
and I_7543 (I130777,I130726,I309119);
not I_7544 (I130794,I309116);
nand I_7545 (I130811,I130794,I309119);
not I_7546 (I130828,I309095);
nor I_7547 (I130845,I130828,I309098);
nand I_7548 (I130862,I130845,I309107);
nor I_7549 (I130879,I130862,I130811);
DFFARX1 I_7550 (I130879,I2507,I130661,I130629,);
not I_7551 (I130910,I130862);
not I_7552 (I130927,I309098);
nand I_7553 (I130944,I130927,I309119);
nor I_7554 (I130961,I309098,I309116);
nand I_7555 (I130641,I130777,I130961);
nand I_7556 (I130635,I130726,I309098);
nand I_7557 (I131006,I130828,I309113);
DFFARX1 I_7558 (I131006,I2507,I130661,I130650,);
DFFARX1 I_7559 (I131006,I2507,I130661,I130644,);
not I_7560 (I131051,I309113);
nor I_7561 (I131068,I131051,I309095);
and I_7562 (I131085,I131068,I309104);
or I_7563 (I131102,I131085,I309098);
DFFARX1 I_7564 (I131102,I2507,I130661,I131128,);
nand I_7565 (I131136,I131128,I130794);
nor I_7566 (I130638,I131136,I130944);
nor I_7567 (I130632,I131128,I130760);
DFFARX1 I_7568 (I131128,I2507,I130661,I131190,);
not I_7569 (I131198,I131190);
nor I_7570 (I130647,I131198,I130910);
not I_7571 (I131256,I2514);
DFFARX1 I_7572 (I468697,I2507,I131256,I131282,);
DFFARX1 I_7573 (I131282,I2507,I131256,I131299,);
not I_7574 (I131248,I131299);
not I_7575 (I131321,I131282);
DFFARX1 I_7576 (I468691,I2507,I131256,I131347,);
not I_7577 (I131355,I131347);
and I_7578 (I131372,I131321,I468709);
not I_7579 (I131389,I468697);
nand I_7580 (I131406,I131389,I468709);
not I_7581 (I131423,I468691);
nor I_7582 (I131440,I131423,I468703);
nand I_7583 (I131457,I131440,I468694);
nor I_7584 (I131474,I131457,I131406);
DFFARX1 I_7585 (I131474,I2507,I131256,I131224,);
not I_7586 (I131505,I131457);
not I_7587 (I131522,I468703);
nand I_7588 (I131539,I131522,I468709);
nor I_7589 (I131556,I468703,I468697);
nand I_7590 (I131236,I131372,I131556);
nand I_7591 (I131230,I131321,I468703);
nand I_7592 (I131601,I131423,I468706);
DFFARX1 I_7593 (I131601,I2507,I131256,I131245,);
DFFARX1 I_7594 (I131601,I2507,I131256,I131239,);
not I_7595 (I131646,I468706);
nor I_7596 (I131663,I131646,I468712);
and I_7597 (I131680,I131663,I468694);
or I_7598 (I131697,I131680,I468700);
DFFARX1 I_7599 (I131697,I2507,I131256,I131723,);
nand I_7600 (I131731,I131723,I131389);
nor I_7601 (I131233,I131731,I131539);
nor I_7602 (I131227,I131723,I131355);
DFFARX1 I_7603 (I131723,I2507,I131256,I131785,);
not I_7604 (I131793,I131785);
nor I_7605 (I131242,I131793,I131505);
not I_7606 (I131851,I2514);
DFFARX1 I_7607 (I524823,I2507,I131851,I131877,);
DFFARX1 I_7608 (I131877,I2507,I131851,I131894,);
not I_7609 (I131843,I131894);
not I_7610 (I131916,I131877);
DFFARX1 I_7611 (I524832,I2507,I131851,I131942,);
not I_7612 (I131950,I131942);
and I_7613 (I131967,I131916,I524820);
not I_7614 (I131984,I524811);
nand I_7615 (I132001,I131984,I524820);
not I_7616 (I132018,I524817);
nor I_7617 (I132035,I132018,I524835);
nand I_7618 (I132052,I132035,I524808);
nor I_7619 (I132069,I132052,I132001);
DFFARX1 I_7620 (I132069,I2507,I131851,I131819,);
not I_7621 (I132100,I132052);
not I_7622 (I132117,I524835);
nand I_7623 (I132134,I132117,I524820);
nor I_7624 (I132151,I524835,I524811);
nand I_7625 (I131831,I131967,I132151);
nand I_7626 (I131825,I131916,I524835);
nand I_7627 (I132196,I132018,I524814);
DFFARX1 I_7628 (I132196,I2507,I131851,I131840,);
DFFARX1 I_7629 (I132196,I2507,I131851,I131834,);
not I_7630 (I132241,I524814);
nor I_7631 (I132258,I132241,I524826);
and I_7632 (I132275,I132258,I524808);
or I_7633 (I132292,I132275,I524829);
DFFARX1 I_7634 (I132292,I2507,I131851,I132318,);
nand I_7635 (I132326,I132318,I131984);
nor I_7636 (I131828,I132326,I132134);
nor I_7637 (I131822,I132318,I131950);
DFFARX1 I_7638 (I132318,I2507,I131851,I132380,);
not I_7639 (I132388,I132380);
nor I_7640 (I131837,I132388,I132100);
not I_7641 (I132446,I2514);
DFFARX1 I_7642 (I418927,I2507,I132446,I132472,);
DFFARX1 I_7643 (I132472,I2507,I132446,I132489,);
not I_7644 (I132438,I132489);
not I_7645 (I132511,I132472);
DFFARX1 I_7646 (I418924,I2507,I132446,I132537,);
not I_7647 (I132545,I132537);
and I_7648 (I132562,I132511,I418930);
not I_7649 (I132579,I418915);
nand I_7650 (I132596,I132579,I418930);
not I_7651 (I132613,I418918);
nor I_7652 (I132630,I132613,I418939);
nand I_7653 (I132647,I132630,I418936);
nor I_7654 (I132664,I132647,I132596);
DFFARX1 I_7655 (I132664,I2507,I132446,I132414,);
not I_7656 (I132695,I132647);
not I_7657 (I132712,I418939);
nand I_7658 (I132729,I132712,I418930);
nor I_7659 (I132746,I418939,I418915);
nand I_7660 (I132426,I132562,I132746);
nand I_7661 (I132420,I132511,I418939);
nand I_7662 (I132791,I132613,I418915);
DFFARX1 I_7663 (I132791,I2507,I132446,I132435,);
DFFARX1 I_7664 (I132791,I2507,I132446,I132429,);
not I_7665 (I132836,I418915);
nor I_7666 (I132853,I132836,I418921);
and I_7667 (I132870,I132853,I418933);
or I_7668 (I132887,I132870,I418918);
DFFARX1 I_7669 (I132887,I2507,I132446,I132913,);
nand I_7670 (I132921,I132913,I132579);
nor I_7671 (I132423,I132921,I132729);
nor I_7672 (I132417,I132913,I132545);
DFFARX1 I_7673 (I132913,I2507,I132446,I132975,);
not I_7674 (I132983,I132975);
nor I_7675 (I132432,I132983,I132695);
not I_7676 (I133041,I2514);
DFFARX1 I_7677 (I504797,I2507,I133041,I133067,);
DFFARX1 I_7678 (I133067,I2507,I133041,I133084,);
not I_7679 (I133033,I133084);
not I_7680 (I133106,I133067);
DFFARX1 I_7681 (I504806,I2507,I133041,I133132,);
not I_7682 (I133140,I133132);
and I_7683 (I133157,I133106,I504794);
not I_7684 (I133174,I504785);
nand I_7685 (I133191,I133174,I504794);
not I_7686 (I133208,I504791);
nor I_7687 (I133225,I133208,I504809);
nand I_7688 (I133242,I133225,I504782);
nor I_7689 (I133259,I133242,I133191);
DFFARX1 I_7690 (I133259,I2507,I133041,I133009,);
not I_7691 (I133290,I133242);
not I_7692 (I133307,I504809);
nand I_7693 (I133324,I133307,I504794);
nor I_7694 (I133341,I504809,I504785);
nand I_7695 (I133021,I133157,I133341);
nand I_7696 (I133015,I133106,I504809);
nand I_7697 (I133386,I133208,I504788);
DFFARX1 I_7698 (I133386,I2507,I133041,I133030,);
DFFARX1 I_7699 (I133386,I2507,I133041,I133024,);
not I_7700 (I133431,I504788);
nor I_7701 (I133448,I133431,I504800);
and I_7702 (I133465,I133448,I504782);
or I_7703 (I133482,I133465,I504803);
DFFARX1 I_7704 (I133482,I2507,I133041,I133508,);
nand I_7705 (I133516,I133508,I133174);
nor I_7706 (I133018,I133516,I133324);
nor I_7707 (I133012,I133508,I133140);
DFFARX1 I_7708 (I133508,I2507,I133041,I133570,);
not I_7709 (I133578,I133570);
nor I_7710 (I133027,I133578,I133290);
not I_7711 (I133636,I2514);
DFFARX1 I_7712 (I451306,I2507,I133636,I133662,);
DFFARX1 I_7713 (I133662,I2507,I133636,I133679,);
not I_7714 (I133628,I133679);
not I_7715 (I133701,I133662);
DFFARX1 I_7716 (I451300,I2507,I133636,I133727,);
not I_7717 (I133735,I133727);
and I_7718 (I133752,I133701,I451318);
not I_7719 (I133769,I451306);
nand I_7720 (I133786,I133769,I451318);
not I_7721 (I133803,I451300);
nor I_7722 (I133820,I133803,I451312);
nand I_7723 (I133837,I133820,I451303);
nor I_7724 (I133854,I133837,I133786);
DFFARX1 I_7725 (I133854,I2507,I133636,I133604,);
not I_7726 (I133885,I133837);
not I_7727 (I133902,I451312);
nand I_7728 (I133919,I133902,I451318);
nor I_7729 (I133936,I451312,I451306);
nand I_7730 (I133616,I133752,I133936);
nand I_7731 (I133610,I133701,I451312);
nand I_7732 (I133981,I133803,I451315);
DFFARX1 I_7733 (I133981,I2507,I133636,I133625,);
DFFARX1 I_7734 (I133981,I2507,I133636,I133619,);
not I_7735 (I134026,I451315);
nor I_7736 (I134043,I134026,I451321);
and I_7737 (I134060,I134043,I451303);
or I_7738 (I134077,I134060,I451309);
DFFARX1 I_7739 (I134077,I2507,I133636,I134103,);
nand I_7740 (I134111,I134103,I133769);
nor I_7741 (I133613,I134111,I133919);
nor I_7742 (I133607,I134103,I133735);
DFFARX1 I_7743 (I134103,I2507,I133636,I134165,);
not I_7744 (I134173,I134165);
nor I_7745 (I133622,I134173,I133885);
not I_7746 (I134231,I2514);
DFFARX1 I_7747 (I673442,I2507,I134231,I134257,);
DFFARX1 I_7748 (I134257,I2507,I134231,I134274,);
not I_7749 (I134223,I134274);
not I_7750 (I134296,I134257);
DFFARX1 I_7751 (I673454,I2507,I134231,I134322,);
not I_7752 (I134330,I134322);
and I_7753 (I134347,I134296,I673448);
not I_7754 (I134364,I673460);
nand I_7755 (I134381,I134364,I673448);
not I_7756 (I134398,I673445);
nor I_7757 (I134415,I134398,I673457);
nand I_7758 (I134432,I134415,I673439);
nor I_7759 (I134449,I134432,I134381);
DFFARX1 I_7760 (I134449,I2507,I134231,I134199,);
not I_7761 (I134480,I134432);
not I_7762 (I134497,I673457);
nand I_7763 (I134514,I134497,I673448);
nor I_7764 (I134531,I673457,I673460);
nand I_7765 (I134211,I134347,I134531);
nand I_7766 (I134205,I134296,I673457);
nand I_7767 (I134576,I134398,I673451);
DFFARX1 I_7768 (I134576,I2507,I134231,I134220,);
DFFARX1 I_7769 (I134576,I2507,I134231,I134214,);
not I_7770 (I134621,I673451);
nor I_7771 (I134638,I134621,I673442);
and I_7772 (I134655,I134638,I673439);
or I_7773 (I134672,I134655,I673463);
DFFARX1 I_7774 (I134672,I2507,I134231,I134698,);
nand I_7775 (I134706,I134698,I134364);
nor I_7776 (I134208,I134706,I134514);
nor I_7777 (I134202,I134698,I134330);
DFFARX1 I_7778 (I134698,I2507,I134231,I134760,);
not I_7779 (I134768,I134760);
nor I_7780 (I134217,I134768,I134480);
not I_7781 (I134826,I2514);
DFFARX1 I_7782 (I643095,I2507,I134826,I134852,);
DFFARX1 I_7783 (I134852,I2507,I134826,I134869,);
not I_7784 (I134818,I134869);
not I_7785 (I134891,I134852);
DFFARX1 I_7786 (I643080,I2507,I134826,I134917,);
not I_7787 (I134925,I134917);
and I_7788 (I134942,I134891,I643098);
not I_7789 (I134959,I643080);
nand I_7790 (I134976,I134959,I643098);
not I_7791 (I134993,I643101);
nor I_7792 (I135010,I134993,I643092);
nand I_7793 (I135027,I135010,I643089);
nor I_7794 (I135044,I135027,I134976);
DFFARX1 I_7795 (I135044,I2507,I134826,I134794,);
not I_7796 (I135075,I135027);
not I_7797 (I135092,I643092);
nand I_7798 (I135109,I135092,I643098);
nor I_7799 (I135126,I643092,I643080);
nand I_7800 (I134806,I134942,I135126);
nand I_7801 (I134800,I134891,I643092);
nand I_7802 (I135171,I134993,I643086);
DFFARX1 I_7803 (I135171,I2507,I134826,I134815,);
DFFARX1 I_7804 (I135171,I2507,I134826,I134809,);
not I_7805 (I135216,I643086);
nor I_7806 (I135233,I135216,I643077);
and I_7807 (I135250,I135233,I643083);
or I_7808 (I135267,I135250,I643077);
DFFARX1 I_7809 (I135267,I2507,I134826,I135293,);
nand I_7810 (I135301,I135293,I134959);
nor I_7811 (I134803,I135301,I135109);
nor I_7812 (I134797,I135293,I134925);
DFFARX1 I_7813 (I135293,I2507,I134826,I135355,);
not I_7814 (I135363,I135355);
nor I_7815 (I134812,I135363,I135075);
not I_7816 (I135421,I2514);
DFFARX1 I_7817 (I293875,I2507,I135421,I135447,);
DFFARX1 I_7818 (I135447,I2507,I135421,I135464,);
not I_7819 (I135413,I135464);
not I_7820 (I135486,I135447);
DFFARX1 I_7821 (I293869,I2507,I135421,I135512,);
not I_7822 (I135520,I135512);
and I_7823 (I135537,I135486,I293884);
not I_7824 (I135554,I293881);
nand I_7825 (I135571,I135554,I293884);
not I_7826 (I135588,I293872);
nor I_7827 (I135605,I135588,I293863);
nand I_7828 (I135622,I135605,I293866);
nor I_7829 (I135639,I135622,I135571);
DFFARX1 I_7830 (I135639,I2507,I135421,I135389,);
not I_7831 (I135670,I135622);
not I_7832 (I135687,I293863);
nand I_7833 (I135704,I135687,I293884);
nor I_7834 (I135721,I293863,I293881);
nand I_7835 (I135401,I135537,I135721);
nand I_7836 (I135395,I135486,I293863);
nand I_7837 (I135766,I135588,I293887);
DFFARX1 I_7838 (I135766,I2507,I135421,I135410,);
DFFARX1 I_7839 (I135766,I2507,I135421,I135404,);
not I_7840 (I135811,I293887);
nor I_7841 (I135828,I135811,I293878);
and I_7842 (I135845,I135828,I293863);
or I_7843 (I135862,I135845,I293866);
DFFARX1 I_7844 (I135862,I2507,I135421,I135888,);
nand I_7845 (I135896,I135888,I135554);
nor I_7846 (I135398,I135896,I135704);
nor I_7847 (I135392,I135888,I135520);
DFFARX1 I_7848 (I135888,I2507,I135421,I135950,);
not I_7849 (I135958,I135950);
nor I_7850 (I135407,I135958,I135670);
not I_7851 (I136016,I2514);
DFFARX1 I_7852 (I166380,I2507,I136016,I136042,);
DFFARX1 I_7853 (I136042,I2507,I136016,I136059,);
not I_7854 (I136008,I136059);
not I_7855 (I136081,I136042);
DFFARX1 I_7856 (I166395,I2507,I136016,I136107,);
not I_7857 (I136115,I136107);
and I_7858 (I136132,I136081,I166392);
not I_7859 (I136149,I166380);
nand I_7860 (I136166,I136149,I166392);
not I_7861 (I136183,I166389);
nor I_7862 (I136200,I136183,I166404);
nand I_7863 (I136217,I136200,I166401);
nor I_7864 (I136234,I136217,I136166);
DFFARX1 I_7865 (I136234,I2507,I136016,I135984,);
not I_7866 (I136265,I136217);
not I_7867 (I136282,I166404);
nand I_7868 (I136299,I136282,I166392);
nor I_7869 (I136316,I166404,I166380);
nand I_7870 (I135996,I136132,I136316);
nand I_7871 (I135990,I136081,I166404);
nand I_7872 (I136361,I136183,I166398);
DFFARX1 I_7873 (I136361,I2507,I136016,I136005,);
DFFARX1 I_7874 (I136361,I2507,I136016,I135999,);
not I_7875 (I136406,I166398);
nor I_7876 (I136423,I136406,I166386);
and I_7877 (I136440,I136423,I166407);
or I_7878 (I136457,I136440,I166383);
DFFARX1 I_7879 (I136457,I2507,I136016,I136483,);
nand I_7880 (I136491,I136483,I136149);
nor I_7881 (I135993,I136491,I136299);
nor I_7882 (I135987,I136483,I136115);
DFFARX1 I_7883 (I136483,I2507,I136016,I136545,);
not I_7884 (I136553,I136545);
nor I_7885 (I136002,I136553,I136265);
not I_7886 (I136611,I2514);
DFFARX1 I_7887 (I626009,I2507,I136611,I136637,);
DFFARX1 I_7888 (I136637,I2507,I136611,I136654,);
not I_7889 (I136603,I136654);
not I_7890 (I136676,I136637);
DFFARX1 I_7891 (I626009,I2507,I136611,I136702,);
not I_7892 (I136710,I136702);
and I_7893 (I136727,I136676,I626012);
not I_7894 (I136744,I626024);
nand I_7895 (I136761,I136744,I626012);
not I_7896 (I136778,I626030);
nor I_7897 (I136795,I136778,I626021);
nand I_7898 (I136812,I136795,I626027);
nor I_7899 (I136829,I136812,I136761);
DFFARX1 I_7900 (I136829,I2507,I136611,I136579,);
not I_7901 (I136860,I136812);
not I_7902 (I136877,I626021);
nand I_7903 (I136894,I136877,I626012);
nor I_7904 (I136911,I626021,I626024);
nand I_7905 (I136591,I136727,I136911);
nand I_7906 (I136585,I136676,I626021);
nand I_7907 (I136956,I136778,I626018);
DFFARX1 I_7908 (I136956,I2507,I136611,I136600,);
DFFARX1 I_7909 (I136956,I2507,I136611,I136594,);
not I_7910 (I137001,I626018);
nor I_7911 (I137018,I137001,I626015);
and I_7912 (I137035,I137018,I626033);
or I_7913 (I137052,I137035,I626012);
DFFARX1 I_7914 (I137052,I2507,I136611,I137078,);
nand I_7915 (I137086,I137078,I136744);
nor I_7916 (I136588,I137086,I136894);
nor I_7917 (I136582,I137078,I136710);
DFFARX1 I_7918 (I137078,I2507,I136611,I137140,);
not I_7919 (I137148,I137140);
nor I_7920 (I136597,I137148,I136860);
not I_7921 (I137206,I2514);
DFFARX1 I_7922 (I486709,I2507,I137206,I137232,);
DFFARX1 I_7923 (I137232,I2507,I137206,I137249,);
not I_7924 (I137198,I137249);
not I_7925 (I137271,I137232);
DFFARX1 I_7926 (I486718,I2507,I137206,I137297,);
not I_7927 (I137305,I137297);
and I_7928 (I137322,I137271,I486706);
not I_7929 (I137339,I486697);
nand I_7930 (I137356,I137339,I486706);
not I_7931 (I137373,I486703);
nor I_7932 (I137390,I137373,I486721);
nand I_7933 (I137407,I137390,I486694);
nor I_7934 (I137424,I137407,I137356);
DFFARX1 I_7935 (I137424,I2507,I137206,I137174,);
not I_7936 (I137455,I137407);
not I_7937 (I137472,I486721);
nand I_7938 (I137489,I137472,I486706);
nor I_7939 (I137506,I486721,I486697);
nand I_7940 (I137186,I137322,I137506);
nand I_7941 (I137180,I137271,I486721);
nand I_7942 (I137551,I137373,I486700);
DFFARX1 I_7943 (I137551,I2507,I137206,I137195,);
DFFARX1 I_7944 (I137551,I2507,I137206,I137189,);
not I_7945 (I137596,I486700);
nor I_7946 (I137613,I137596,I486712);
and I_7947 (I137630,I137613,I486694);
or I_7948 (I137647,I137630,I486715);
DFFARX1 I_7949 (I137647,I2507,I137206,I137673,);
nand I_7950 (I137681,I137673,I137339);
nor I_7951 (I137183,I137681,I137489);
nor I_7952 (I137177,I137673,I137305);
DFFARX1 I_7953 (I137673,I2507,I137206,I137735,);
not I_7954 (I137743,I137735);
nor I_7955 (I137192,I137743,I137455);
not I_7956 (I137801,I2514);
DFFARX1 I_7957 (I370375,I2507,I137801,I137827,);
DFFARX1 I_7958 (I137827,I2507,I137801,I137844,);
not I_7959 (I137793,I137844);
not I_7960 (I137866,I137827);
DFFARX1 I_7961 (I370372,I2507,I137801,I137892,);
not I_7962 (I137900,I137892);
and I_7963 (I137917,I137866,I370378);
not I_7964 (I137934,I370363);
nand I_7965 (I137951,I137934,I370378);
not I_7966 (I137968,I370366);
nor I_7967 (I137985,I137968,I370387);
nand I_7968 (I138002,I137985,I370384);
nor I_7969 (I138019,I138002,I137951);
DFFARX1 I_7970 (I138019,I2507,I137801,I137769,);
not I_7971 (I138050,I138002);
not I_7972 (I138067,I370387);
nand I_7973 (I138084,I138067,I370378);
nor I_7974 (I138101,I370387,I370363);
nand I_7975 (I137781,I137917,I138101);
nand I_7976 (I137775,I137866,I370387);
nand I_7977 (I138146,I137968,I370363);
DFFARX1 I_7978 (I138146,I2507,I137801,I137790,);
DFFARX1 I_7979 (I138146,I2507,I137801,I137784,);
not I_7980 (I138191,I370363);
nor I_7981 (I138208,I138191,I370369);
and I_7982 (I138225,I138208,I370381);
or I_7983 (I138242,I138225,I370366);
DFFARX1 I_7984 (I138242,I2507,I137801,I138268,);
nand I_7985 (I138276,I138268,I137934);
nor I_7986 (I137778,I138276,I138084);
nor I_7987 (I137772,I138268,I137900);
DFFARX1 I_7988 (I138268,I2507,I137801,I138330,);
not I_7989 (I138338,I138330);
nor I_7990 (I137787,I138338,I138050);
not I_7991 (I138396,I2514);
DFFARX1 I_7992 (I527407,I2507,I138396,I138422,);
DFFARX1 I_7993 (I138422,I2507,I138396,I138439,);
not I_7994 (I138388,I138439);
not I_7995 (I138461,I138422);
DFFARX1 I_7996 (I527416,I2507,I138396,I138487,);
not I_7997 (I138495,I138487);
and I_7998 (I138512,I138461,I527404);
not I_7999 (I138529,I527395);
nand I_8000 (I138546,I138529,I527404);
not I_8001 (I138563,I527401);
nor I_8002 (I138580,I138563,I527419);
nand I_8003 (I138597,I138580,I527392);
nor I_8004 (I138614,I138597,I138546);
DFFARX1 I_8005 (I138614,I2507,I138396,I138364,);
not I_8006 (I138645,I138597);
not I_8007 (I138662,I527419);
nand I_8008 (I138679,I138662,I527404);
nor I_8009 (I138696,I527419,I527395);
nand I_8010 (I138376,I138512,I138696);
nand I_8011 (I138370,I138461,I527419);
nand I_8012 (I138741,I138563,I527398);
DFFARX1 I_8013 (I138741,I2507,I138396,I138385,);
DFFARX1 I_8014 (I138741,I2507,I138396,I138379,);
not I_8015 (I138786,I527398);
nor I_8016 (I138803,I138786,I527410);
and I_8017 (I138820,I138803,I527392);
or I_8018 (I138837,I138820,I527413);
DFFARX1 I_8019 (I138837,I2507,I138396,I138863,);
nand I_8020 (I138871,I138863,I138529);
nor I_8021 (I138373,I138871,I138679);
nor I_8022 (I138367,I138863,I138495);
DFFARX1 I_8023 (I138863,I2507,I138396,I138925,);
not I_8024 (I138933,I138925);
nor I_8025 (I138382,I138933,I138645);
not I_8026 (I138991,I2514);
DFFARX1 I_8027 (I69404,I2507,I138991,I139017,);
DFFARX1 I_8028 (I139017,I2507,I138991,I139034,);
not I_8029 (I138983,I139034);
not I_8030 (I139056,I139017);
DFFARX1 I_8031 (I69398,I2507,I138991,I139082,);
not I_8032 (I139090,I139082);
and I_8033 (I139107,I139056,I69395);
not I_8034 (I139124,I69416);
nand I_8035 (I139141,I139124,I69395);
not I_8036 (I139158,I69410);
nor I_8037 (I139175,I139158,I69401);
nand I_8038 (I139192,I139175,I69407);
nor I_8039 (I139209,I139192,I139141);
DFFARX1 I_8040 (I139209,I2507,I138991,I138959,);
not I_8041 (I139240,I139192);
not I_8042 (I139257,I69401);
nand I_8043 (I139274,I139257,I69395);
nor I_8044 (I139291,I69401,I69416);
nand I_8045 (I138971,I139107,I139291);
nand I_8046 (I138965,I139056,I69401);
nand I_8047 (I139336,I139158,I69395);
DFFARX1 I_8048 (I139336,I2507,I138991,I138980,);
DFFARX1 I_8049 (I139336,I2507,I138991,I138974,);
not I_8050 (I139381,I69395);
nor I_8051 (I139398,I139381,I69413);
and I_8052 (I139415,I139398,I69419);
or I_8053 (I139432,I139415,I69398);
DFFARX1 I_8054 (I139432,I2507,I138991,I139458,);
nand I_8055 (I139466,I139458,I139124);
nor I_8056 (I138968,I139466,I139274);
nor I_8057 (I138962,I139458,I139090);
DFFARX1 I_8058 (I139458,I2507,I138991,I139520,);
not I_8059 (I139528,I139520);
nor I_8060 (I138977,I139528,I139240);
not I_8061 (I139586,I2514);
DFFARX1 I_8062 (I321826,I2507,I139586,I139612,);
DFFARX1 I_8063 (I139612,I2507,I139586,I139629,);
not I_8064 (I139578,I139629);
not I_8065 (I139651,I139612);
DFFARX1 I_8066 (I321817,I2507,I139586,I139677,);
not I_8067 (I139685,I139677);
and I_8068 (I139702,I139651,I321835);
not I_8069 (I139719,I321832);
nand I_8070 (I139736,I139719,I321835);
not I_8071 (I139753,I321811);
nor I_8072 (I139770,I139753,I321814);
nand I_8073 (I139787,I139770,I321823);
nor I_8074 (I139804,I139787,I139736);
DFFARX1 I_8075 (I139804,I2507,I139586,I139554,);
not I_8076 (I139835,I139787);
not I_8077 (I139852,I321814);
nand I_8078 (I139869,I139852,I321835);
nor I_8079 (I139886,I321814,I321832);
nand I_8080 (I139566,I139702,I139886);
nand I_8081 (I139560,I139651,I321814);
nand I_8082 (I139931,I139753,I321829);
DFFARX1 I_8083 (I139931,I2507,I139586,I139575,);
DFFARX1 I_8084 (I139931,I2507,I139586,I139569,);
not I_8085 (I139976,I321829);
nor I_8086 (I139993,I139976,I321811);
and I_8087 (I140010,I139993,I321820);
or I_8088 (I140027,I140010,I321814);
DFFARX1 I_8089 (I140027,I2507,I139586,I140053,);
nand I_8090 (I140061,I140053,I139719);
nor I_8091 (I139563,I140061,I139869);
nor I_8092 (I139557,I140053,I139685);
DFFARX1 I_8093 (I140053,I2507,I139586,I140115,);
not I_8094 (I140123,I140115);
nor I_8095 (I139572,I140123,I139835);
not I_8096 (I140181,I2514);
DFFARX1 I_8097 (I680378,I2507,I140181,I140207,);
DFFARX1 I_8098 (I140207,I2507,I140181,I140224,);
not I_8099 (I140173,I140224);
not I_8100 (I140246,I140207);
DFFARX1 I_8101 (I680390,I2507,I140181,I140272,);
not I_8102 (I140280,I140272);
and I_8103 (I140297,I140246,I680384);
not I_8104 (I140314,I680396);
nand I_8105 (I140331,I140314,I680384);
not I_8106 (I140348,I680381);
nor I_8107 (I140365,I140348,I680393);
nand I_8108 (I140382,I140365,I680375);
nor I_8109 (I140399,I140382,I140331);
DFFARX1 I_8110 (I140399,I2507,I140181,I140149,);
not I_8111 (I140430,I140382);
not I_8112 (I140447,I680393);
nand I_8113 (I140464,I140447,I680384);
nor I_8114 (I140481,I680393,I680396);
nand I_8115 (I140161,I140297,I140481);
nand I_8116 (I140155,I140246,I680393);
nand I_8117 (I140526,I140348,I680387);
DFFARX1 I_8118 (I140526,I2507,I140181,I140170,);
DFFARX1 I_8119 (I140526,I2507,I140181,I140164,);
not I_8120 (I140571,I680387);
nor I_8121 (I140588,I140571,I680378);
and I_8122 (I140605,I140588,I680375);
or I_8123 (I140622,I140605,I680399);
DFFARX1 I_8124 (I140622,I2507,I140181,I140648,);
nand I_8125 (I140656,I140648,I140314);
nor I_8126 (I140158,I140656,I140464);
nor I_8127 (I140152,I140648,I140280);
DFFARX1 I_8128 (I140648,I2507,I140181,I140710,);
not I_8129 (I140718,I140710);
nor I_8130 (I140167,I140718,I140430);
not I_8131 (I140776,I2514);
DFFARX1 I_8132 (I227536,I2507,I140776,I140802,);
DFFARX1 I_8133 (I140802,I2507,I140776,I140819,);
not I_8134 (I140768,I140819);
not I_8135 (I140841,I140802);
DFFARX1 I_8136 (I227524,I2507,I140776,I140867,);
not I_8137 (I140875,I140867);
and I_8138 (I140892,I140841,I227533);
not I_8139 (I140909,I227530);
nand I_8140 (I140926,I140909,I227533);
not I_8141 (I140943,I227521);
nor I_8142 (I140960,I140943,I227527);
nand I_8143 (I140977,I140960,I227512);
nor I_8144 (I140994,I140977,I140926);
DFFARX1 I_8145 (I140994,I2507,I140776,I140744,);
not I_8146 (I141025,I140977);
not I_8147 (I141042,I227527);
nand I_8148 (I141059,I141042,I227533);
nor I_8149 (I141076,I227527,I227530);
nand I_8150 (I140756,I140892,I141076);
nand I_8151 (I140750,I140841,I227527);
nand I_8152 (I141121,I140943,I227512);
DFFARX1 I_8153 (I141121,I2507,I140776,I140765,);
DFFARX1 I_8154 (I141121,I2507,I140776,I140759,);
not I_8155 (I141166,I227512);
nor I_8156 (I141183,I141166,I227518);
and I_8157 (I141200,I141183,I227515);
or I_8158 (I141217,I141200,I227539);
DFFARX1 I_8159 (I141217,I2507,I140776,I141243,);
nand I_8160 (I141251,I141243,I140909);
nor I_8161 (I140753,I141251,I141059);
nor I_8162 (I140747,I141243,I140875);
DFFARX1 I_8163 (I141243,I2507,I140776,I141305,);
not I_8164 (I141313,I141305);
nor I_8165 (I140762,I141313,I141025);
not I_8166 (I141371,I2514);
DFFARX1 I_8167 (I685553,I2507,I141371,I141397,);
DFFARX1 I_8168 (I141397,I2507,I141371,I141414,);
not I_8169 (I141363,I141414);
not I_8170 (I141436,I141397);
DFFARX1 I_8171 (I685526,I2507,I141371,I141462,);
not I_8172 (I141470,I141462);
and I_8173 (I141487,I141436,I685550);
not I_8174 (I141504,I685547);
nand I_8175 (I141521,I141504,I685550);
not I_8176 (I141538,I685526);
nor I_8177 (I141555,I141538,I685544);
nand I_8178 (I141572,I141555,I685532);
nor I_8179 (I141589,I141572,I141521);
DFFARX1 I_8180 (I141589,I2507,I141371,I141339,);
not I_8181 (I141620,I141572);
not I_8182 (I141637,I685544);
nand I_8183 (I141654,I141637,I685550);
nor I_8184 (I141671,I685544,I685547);
nand I_8185 (I141351,I141487,I141671);
nand I_8186 (I141345,I141436,I685544);
nand I_8187 (I141716,I141538,I685538);
DFFARX1 I_8188 (I141716,I2507,I141371,I141360,);
DFFARX1 I_8189 (I141716,I2507,I141371,I141354,);
not I_8190 (I141761,I685538);
nor I_8191 (I141778,I141761,I685541);
and I_8192 (I141795,I141778,I685529);
or I_8193 (I141812,I141795,I685535);
DFFARX1 I_8194 (I141812,I2507,I141371,I141838,);
nand I_8195 (I141846,I141838,I141504);
nor I_8196 (I141348,I141846,I141654);
nor I_8197 (I141342,I141838,I141470);
DFFARX1 I_8198 (I141838,I2507,I141371,I141900,);
not I_8199 (I141908,I141900);
nor I_8200 (I141357,I141908,I141620);
not I_8201 (I141966,I2514);
DFFARX1 I_8202 (I631211,I2507,I141966,I141992,);
DFFARX1 I_8203 (I141992,I2507,I141966,I142009,);
not I_8204 (I141958,I142009);
not I_8205 (I142031,I141992);
DFFARX1 I_8206 (I631211,I2507,I141966,I142057,);
not I_8207 (I142065,I142057);
and I_8208 (I142082,I142031,I631214);
not I_8209 (I142099,I631226);
nand I_8210 (I142116,I142099,I631214);
not I_8211 (I142133,I631232);
nor I_8212 (I142150,I142133,I631223);
nand I_8213 (I142167,I142150,I631229);
nor I_8214 (I142184,I142167,I142116);
DFFARX1 I_8215 (I142184,I2507,I141966,I141934,);
not I_8216 (I142215,I142167);
not I_8217 (I142232,I631223);
nand I_8218 (I142249,I142232,I631214);
nor I_8219 (I142266,I631223,I631226);
nand I_8220 (I141946,I142082,I142266);
nand I_8221 (I141940,I142031,I631223);
nand I_8222 (I142311,I142133,I631220);
DFFARX1 I_8223 (I142311,I2507,I141966,I141955,);
DFFARX1 I_8224 (I142311,I2507,I141966,I141949,);
not I_8225 (I142356,I631220);
nor I_8226 (I142373,I142356,I631217);
and I_8227 (I142390,I142373,I631235);
or I_8228 (I142407,I142390,I631214);
DFFARX1 I_8229 (I142407,I2507,I141966,I142433,);
nand I_8230 (I142441,I142433,I142099);
nor I_8231 (I141943,I142441,I142249);
nor I_8232 (I141937,I142433,I142065);
DFFARX1 I_8233 (I142433,I2507,I141966,I142495,);
not I_8234 (I142503,I142495);
nor I_8235 (I141952,I142503,I142215);
not I_8236 (I142561,I2514);
DFFARX1 I_8237 (I516425,I2507,I142561,I142587,);
DFFARX1 I_8238 (I142587,I2507,I142561,I142604,);
not I_8239 (I142553,I142604);
not I_8240 (I142626,I142587);
DFFARX1 I_8241 (I516434,I2507,I142561,I142652,);
not I_8242 (I142660,I142652);
and I_8243 (I142677,I142626,I516422);
not I_8244 (I142694,I516413);
nand I_8245 (I142711,I142694,I516422);
not I_8246 (I142728,I516419);
nor I_8247 (I142745,I142728,I516437);
nand I_8248 (I142762,I142745,I516410);
nor I_8249 (I142779,I142762,I142711);
DFFARX1 I_8250 (I142779,I2507,I142561,I142529,);
not I_8251 (I142810,I142762);
not I_8252 (I142827,I516437);
nand I_8253 (I142844,I142827,I516422);
nor I_8254 (I142861,I516437,I516413);
nand I_8255 (I142541,I142677,I142861);
nand I_8256 (I142535,I142626,I516437);
nand I_8257 (I142906,I142728,I516416);
DFFARX1 I_8258 (I142906,I2507,I142561,I142550,);
DFFARX1 I_8259 (I142906,I2507,I142561,I142544,);
not I_8260 (I142951,I516416);
nor I_8261 (I142968,I142951,I516428);
and I_8262 (I142985,I142968,I516410);
or I_8263 (I143002,I142985,I516431);
DFFARX1 I_8264 (I143002,I2507,I142561,I143028,);
nand I_8265 (I143036,I143028,I142694);
nor I_8266 (I142538,I143036,I142844);
nor I_8267 (I142532,I143028,I142660);
DFFARX1 I_8268 (I143028,I2507,I142561,I143090,);
not I_8269 (I143098,I143090);
nor I_8270 (I142547,I143098,I142810);
not I_8271 (I143156,I2514);
DFFARX1 I_8272 (I279760,I2507,I143156,I143182,);
DFFARX1 I_8273 (I143182,I2507,I143156,I143199,);
not I_8274 (I143148,I143199);
not I_8275 (I143221,I143182);
DFFARX1 I_8276 (I279748,I2507,I143156,I143247,);
not I_8277 (I143255,I143247);
and I_8278 (I143272,I143221,I279757);
not I_8279 (I143289,I279754);
nand I_8280 (I143306,I143289,I279757);
not I_8281 (I143323,I279745);
nor I_8282 (I143340,I143323,I279751);
nand I_8283 (I143357,I143340,I279736);
nor I_8284 (I143374,I143357,I143306);
DFFARX1 I_8285 (I143374,I2507,I143156,I143124,);
not I_8286 (I143405,I143357);
not I_8287 (I143422,I279751);
nand I_8288 (I143439,I143422,I279757);
nor I_8289 (I143456,I279751,I279754);
nand I_8290 (I143136,I143272,I143456);
nand I_8291 (I143130,I143221,I279751);
nand I_8292 (I143501,I143323,I279736);
DFFARX1 I_8293 (I143501,I2507,I143156,I143145,);
DFFARX1 I_8294 (I143501,I2507,I143156,I143139,);
not I_8295 (I143546,I279736);
nor I_8296 (I143563,I143546,I279742);
and I_8297 (I143580,I143563,I279739);
or I_8298 (I143597,I143580,I279763);
DFFARX1 I_8299 (I143597,I2507,I143156,I143623,);
nand I_8300 (I143631,I143623,I143289);
nor I_8301 (I143133,I143631,I143439);
nor I_8302 (I143127,I143623,I143255);
DFFARX1 I_8303 (I143623,I2507,I143156,I143685,);
not I_8304 (I143693,I143685);
nor I_8305 (I143142,I143693,I143405);
not I_8306 (I143751,I2514);
DFFARX1 I_8307 (I482833,I2507,I143751,I143777,);
DFFARX1 I_8308 (I143777,I2507,I143751,I143794,);
not I_8309 (I143743,I143794);
not I_8310 (I143816,I143777);
DFFARX1 I_8311 (I482842,I2507,I143751,I143842,);
not I_8312 (I143850,I143842);
and I_8313 (I143867,I143816,I482830);
not I_8314 (I143884,I482821);
nand I_8315 (I143901,I143884,I482830);
not I_8316 (I143918,I482827);
nor I_8317 (I143935,I143918,I482845);
nand I_8318 (I143952,I143935,I482818);
nor I_8319 (I143969,I143952,I143901);
DFFARX1 I_8320 (I143969,I2507,I143751,I143719,);
not I_8321 (I144000,I143952);
not I_8322 (I144017,I482845);
nand I_8323 (I144034,I144017,I482830);
nor I_8324 (I144051,I482845,I482821);
nand I_8325 (I143731,I143867,I144051);
nand I_8326 (I143725,I143816,I482845);
nand I_8327 (I144096,I143918,I482824);
DFFARX1 I_8328 (I144096,I2507,I143751,I143740,);
DFFARX1 I_8329 (I144096,I2507,I143751,I143734,);
not I_8330 (I144141,I482824);
nor I_8331 (I144158,I144141,I482836);
and I_8332 (I144175,I144158,I482818);
or I_8333 (I144192,I144175,I482839);
DFFARX1 I_8334 (I144192,I2507,I143751,I144218,);
nand I_8335 (I144226,I144218,I143884);
nor I_8336 (I143728,I144226,I144034);
nor I_8337 (I143722,I144218,I143850);
DFFARX1 I_8338 (I144218,I2507,I143751,I144280,);
not I_8339 (I144288,I144280);
nor I_8340 (I143737,I144288,I144000);
not I_8341 (I144346,I2514);
DFFARX1 I_8342 (I365751,I2507,I144346,I144372,);
DFFARX1 I_8343 (I144372,I2507,I144346,I144389,);
not I_8344 (I144338,I144389);
not I_8345 (I144411,I144372);
DFFARX1 I_8346 (I365748,I2507,I144346,I144437,);
not I_8347 (I144445,I144437);
and I_8348 (I144462,I144411,I365754);
not I_8349 (I144479,I365739);
nand I_8350 (I144496,I144479,I365754);
not I_8351 (I144513,I365742);
nor I_8352 (I144530,I144513,I365763);
nand I_8353 (I144547,I144530,I365760);
nor I_8354 (I144564,I144547,I144496);
DFFARX1 I_8355 (I144564,I2507,I144346,I144314,);
not I_8356 (I144595,I144547);
not I_8357 (I144612,I365763);
nand I_8358 (I144629,I144612,I365754);
nor I_8359 (I144646,I365763,I365739);
nand I_8360 (I144326,I144462,I144646);
nand I_8361 (I144320,I144411,I365763);
nand I_8362 (I144691,I144513,I365739);
DFFARX1 I_8363 (I144691,I2507,I144346,I144335,);
DFFARX1 I_8364 (I144691,I2507,I144346,I144329,);
not I_8365 (I144736,I365739);
nor I_8366 (I144753,I144736,I365745);
and I_8367 (I144770,I144753,I365757);
or I_8368 (I144787,I144770,I365742);
DFFARX1 I_8369 (I144787,I2507,I144346,I144813,);
nand I_8370 (I144821,I144813,I144479);
nor I_8371 (I144323,I144821,I144629);
nor I_8372 (I144317,I144813,I144445);
DFFARX1 I_8373 (I144813,I2507,I144346,I144875,);
not I_8374 (I144883,I144875);
nor I_8375 (I144332,I144883,I144595);
not I_8376 (I144941,I2514);
DFFARX1 I_8377 (I169015,I2507,I144941,I144967,);
DFFARX1 I_8378 (I144967,I2507,I144941,I144984,);
not I_8379 (I144933,I144984);
not I_8380 (I145006,I144967);
DFFARX1 I_8381 (I169030,I2507,I144941,I145032,);
not I_8382 (I145040,I145032);
and I_8383 (I145057,I145006,I169027);
not I_8384 (I145074,I169015);
nand I_8385 (I145091,I145074,I169027);
not I_8386 (I145108,I169024);
nor I_8387 (I145125,I145108,I169039);
nand I_8388 (I145142,I145125,I169036);
nor I_8389 (I145159,I145142,I145091);
DFFARX1 I_8390 (I145159,I2507,I144941,I144909,);
not I_8391 (I145190,I145142);
not I_8392 (I145207,I169039);
nand I_8393 (I145224,I145207,I169027);
nor I_8394 (I145241,I169039,I169015);
nand I_8395 (I144921,I145057,I145241);
nand I_8396 (I144915,I145006,I169039);
nand I_8397 (I145286,I145108,I169033);
DFFARX1 I_8398 (I145286,I2507,I144941,I144930,);
DFFARX1 I_8399 (I145286,I2507,I144941,I144924,);
not I_8400 (I145331,I169033);
nor I_8401 (I145348,I145331,I169021);
and I_8402 (I145365,I145348,I169042);
or I_8403 (I145382,I145365,I169018);
DFFARX1 I_8404 (I145382,I2507,I144941,I145408,);
nand I_8405 (I145416,I145408,I145074);
nor I_8406 (I144918,I145416,I145224);
nor I_8407 (I144912,I145408,I145040);
DFFARX1 I_8408 (I145408,I2507,I144941,I145470,);
not I_8409 (I145478,I145470);
nor I_8410 (I144927,I145478,I145190);
not I_8411 (I145536,I2514);
DFFARX1 I_8412 (I581503,I2507,I145536,I145562,);
DFFARX1 I_8413 (I145562,I2507,I145536,I145579,);
not I_8414 (I145528,I145579);
not I_8415 (I145601,I145562);
DFFARX1 I_8416 (I581503,I2507,I145536,I145627,);
not I_8417 (I145635,I145627);
and I_8418 (I145652,I145601,I581506);
not I_8419 (I145669,I581518);
nand I_8420 (I145686,I145669,I581506);
not I_8421 (I145703,I581524);
nor I_8422 (I145720,I145703,I581515);
nand I_8423 (I145737,I145720,I581521);
nor I_8424 (I145754,I145737,I145686);
DFFARX1 I_8425 (I145754,I2507,I145536,I145504,);
not I_8426 (I145785,I145737);
not I_8427 (I145802,I581515);
nand I_8428 (I145819,I145802,I581506);
nor I_8429 (I145836,I581515,I581518);
nand I_8430 (I145516,I145652,I145836);
nand I_8431 (I145510,I145601,I581515);
nand I_8432 (I145881,I145703,I581512);
DFFARX1 I_8433 (I145881,I2507,I145536,I145525,);
DFFARX1 I_8434 (I145881,I2507,I145536,I145519,);
not I_8435 (I145926,I581512);
nor I_8436 (I145943,I145926,I581509);
and I_8437 (I145960,I145943,I581527);
or I_8438 (I145977,I145960,I581506);
DFFARX1 I_8439 (I145977,I2507,I145536,I146003,);
nand I_8440 (I146011,I146003,I145669);
nor I_8441 (I145513,I146011,I145819);
nor I_8442 (I145507,I146003,I145635);
DFFARX1 I_8443 (I146003,I2507,I145536,I146065,);
not I_8444 (I146073,I146065);
nor I_8445 (I145522,I146073,I145785);
not I_8446 (I146131,I2514);
DFFARX1 I_8447 (I348411,I2507,I146131,I146157,);
DFFARX1 I_8448 (I146157,I2507,I146131,I146174,);
not I_8449 (I146123,I146174);
not I_8450 (I146196,I146157);
DFFARX1 I_8451 (I348408,I2507,I146131,I146222,);
not I_8452 (I146230,I146222);
and I_8453 (I146247,I146196,I348414);
not I_8454 (I146264,I348399);
nand I_8455 (I146281,I146264,I348414);
not I_8456 (I146298,I348402);
nor I_8457 (I146315,I146298,I348423);
nand I_8458 (I146332,I146315,I348420);
nor I_8459 (I146349,I146332,I146281);
DFFARX1 I_8460 (I146349,I2507,I146131,I146099,);
not I_8461 (I146380,I146332);
not I_8462 (I146397,I348423);
nand I_8463 (I146414,I146397,I348414);
nor I_8464 (I146431,I348423,I348399);
nand I_8465 (I146111,I146247,I146431);
nand I_8466 (I146105,I146196,I348423);
nand I_8467 (I146476,I146298,I348399);
DFFARX1 I_8468 (I146476,I2507,I146131,I146120,);
DFFARX1 I_8469 (I146476,I2507,I146131,I146114,);
not I_8470 (I146521,I348399);
nor I_8471 (I146538,I146521,I348405);
and I_8472 (I146555,I146538,I348417);
or I_8473 (I146572,I146555,I348402);
DFFARX1 I_8474 (I146572,I2507,I146131,I146598,);
nand I_8475 (I146606,I146598,I146264);
nor I_8476 (I146108,I146606,I146414);
nor I_8477 (I146102,I146598,I146230);
DFFARX1 I_8478 (I146598,I2507,I146131,I146660,);
not I_8479 (I146668,I146660);
nor I_8480 (I146117,I146668,I146380);
not I_8481 (I146726,I2514);
DFFARX1 I_8482 (I259088,I2507,I146726,I146752,);
DFFARX1 I_8483 (I146752,I2507,I146726,I146769,);
not I_8484 (I146718,I146769);
not I_8485 (I146791,I146752);
DFFARX1 I_8486 (I259076,I2507,I146726,I146817,);
not I_8487 (I146825,I146817);
and I_8488 (I146842,I146791,I259085);
not I_8489 (I146859,I259082);
nand I_8490 (I146876,I146859,I259085);
not I_8491 (I146893,I259073);
nor I_8492 (I146910,I146893,I259079);
nand I_8493 (I146927,I146910,I259064);
nor I_8494 (I146944,I146927,I146876);
DFFARX1 I_8495 (I146944,I2507,I146726,I146694,);
not I_8496 (I146975,I146927);
not I_8497 (I146992,I259079);
nand I_8498 (I147009,I146992,I259085);
nor I_8499 (I147026,I259079,I259082);
nand I_8500 (I146706,I146842,I147026);
nand I_8501 (I146700,I146791,I259079);
nand I_8502 (I147071,I146893,I259064);
DFFARX1 I_8503 (I147071,I2507,I146726,I146715,);
DFFARX1 I_8504 (I147071,I2507,I146726,I146709,);
not I_8505 (I147116,I259064);
nor I_8506 (I147133,I147116,I259070);
and I_8507 (I147150,I147133,I259067);
or I_8508 (I147167,I147150,I259091);
DFFARX1 I_8509 (I147167,I2507,I146726,I147193,);
nand I_8510 (I147201,I147193,I146859);
nor I_8511 (I146703,I147201,I147009);
nor I_8512 (I146697,I147193,I146825);
DFFARX1 I_8513 (I147193,I2507,I146726,I147255,);
not I_8514 (I147263,I147255);
nor I_8515 (I146712,I147263,I146975);
not I_8516 (I147321,I2514);
DFFARX1 I_8517 (I260720,I2507,I147321,I147347,);
DFFARX1 I_8518 (I147347,I2507,I147321,I147364,);
not I_8519 (I147313,I147364);
not I_8520 (I147386,I147347);
DFFARX1 I_8521 (I260708,I2507,I147321,I147412,);
not I_8522 (I147420,I147412);
and I_8523 (I147437,I147386,I260717);
not I_8524 (I147454,I260714);
nand I_8525 (I147471,I147454,I260717);
not I_8526 (I147488,I260705);
nor I_8527 (I147505,I147488,I260711);
nand I_8528 (I147522,I147505,I260696);
nor I_8529 (I147539,I147522,I147471);
DFFARX1 I_8530 (I147539,I2507,I147321,I147289,);
not I_8531 (I147570,I147522);
not I_8532 (I147587,I260711);
nand I_8533 (I147604,I147587,I260717);
nor I_8534 (I147621,I260711,I260714);
nand I_8535 (I147301,I147437,I147621);
nand I_8536 (I147295,I147386,I260711);
nand I_8537 (I147666,I147488,I260696);
DFFARX1 I_8538 (I147666,I2507,I147321,I147310,);
DFFARX1 I_8539 (I147666,I2507,I147321,I147304,);
not I_8540 (I147711,I260696);
nor I_8541 (I147728,I147711,I260702);
and I_8542 (I147745,I147728,I260699);
or I_8543 (I147762,I147745,I260723);
DFFARX1 I_8544 (I147762,I2507,I147321,I147788,);
nand I_8545 (I147796,I147788,I147454);
nor I_8546 (I147298,I147796,I147604);
nor I_8547 (I147292,I147788,I147420);
DFFARX1 I_8548 (I147788,I2507,I147321,I147850,);
not I_8549 (I147858,I147850);
nor I_8550 (I147307,I147858,I147570);
not I_8551 (I147916,I2514);
DFFARX1 I_8552 (I352457,I2507,I147916,I147942,);
DFFARX1 I_8553 (I147942,I2507,I147916,I147959,);
not I_8554 (I147908,I147959);
not I_8555 (I147981,I147942);
DFFARX1 I_8556 (I352454,I2507,I147916,I148007,);
not I_8557 (I148015,I148007);
and I_8558 (I148032,I147981,I352460);
not I_8559 (I148049,I352445);
nand I_8560 (I148066,I148049,I352460);
not I_8561 (I148083,I352448);
nor I_8562 (I148100,I148083,I352469);
nand I_8563 (I148117,I148100,I352466);
nor I_8564 (I148134,I148117,I148066);
DFFARX1 I_8565 (I148134,I2507,I147916,I147884,);
not I_8566 (I148165,I148117);
not I_8567 (I148182,I352469);
nand I_8568 (I148199,I148182,I352460);
nor I_8569 (I148216,I352469,I352445);
nand I_8570 (I147896,I148032,I148216);
nand I_8571 (I147890,I147981,I352469);
nand I_8572 (I148261,I148083,I352445);
DFFARX1 I_8573 (I148261,I2507,I147916,I147905,);
DFFARX1 I_8574 (I148261,I2507,I147916,I147899,);
not I_8575 (I148306,I352445);
nor I_8576 (I148323,I148306,I352451);
and I_8577 (I148340,I148323,I352463);
or I_8578 (I148357,I148340,I352448);
DFFARX1 I_8579 (I148357,I2507,I147916,I148383,);
nand I_8580 (I148391,I148383,I148049);
nor I_8581 (I147893,I148391,I148199);
nor I_8582 (I147887,I148383,I148015);
DFFARX1 I_8583 (I148383,I2507,I147916,I148445,);
not I_8584 (I148453,I148445);
nor I_8585 (I147902,I148453,I148165);
not I_8586 (I148511,I2514);
DFFARX1 I_8587 (I198527,I2507,I148511,I148537,);
DFFARX1 I_8588 (I148537,I2507,I148511,I148554,);
not I_8589 (I148503,I148554);
not I_8590 (I148576,I148537);
DFFARX1 I_8591 (I198542,I2507,I148511,I148602,);
not I_8592 (I148610,I148602);
and I_8593 (I148627,I148576,I198539);
not I_8594 (I148644,I198527);
nand I_8595 (I148661,I148644,I198539);
not I_8596 (I148678,I198536);
nor I_8597 (I148695,I148678,I198551);
nand I_8598 (I148712,I148695,I198548);
nor I_8599 (I148729,I148712,I148661);
DFFARX1 I_8600 (I148729,I2507,I148511,I148479,);
not I_8601 (I148760,I148712);
not I_8602 (I148777,I198551);
nand I_8603 (I148794,I148777,I198539);
nor I_8604 (I148811,I198551,I198527);
nand I_8605 (I148491,I148627,I148811);
nand I_8606 (I148485,I148576,I198551);
nand I_8607 (I148856,I148678,I198545);
DFFARX1 I_8608 (I148856,I2507,I148511,I148500,);
DFFARX1 I_8609 (I148856,I2507,I148511,I148494,);
not I_8610 (I148901,I198545);
nor I_8611 (I148918,I148901,I198533);
and I_8612 (I148935,I148918,I198554);
or I_8613 (I148952,I148935,I198530);
DFFARX1 I_8614 (I148952,I2507,I148511,I148978,);
nand I_8615 (I148986,I148978,I148644);
nor I_8616 (I148488,I148986,I148794);
nor I_8617 (I148482,I148978,I148610);
DFFARX1 I_8618 (I148978,I2507,I148511,I149040,);
not I_8619 (I149048,I149040);
nor I_8620 (I148497,I149048,I148760);
not I_8621 (I149106,I2514);
DFFARX1 I_8622 (I60445,I2507,I149106,I149132,);
DFFARX1 I_8623 (I149132,I2507,I149106,I149149,);
not I_8624 (I149098,I149149);
not I_8625 (I149171,I149132);
DFFARX1 I_8626 (I60439,I2507,I149106,I149197,);
not I_8627 (I149205,I149197);
and I_8628 (I149222,I149171,I60436);
not I_8629 (I149239,I60457);
nand I_8630 (I149256,I149239,I60436);
not I_8631 (I149273,I60451);
nor I_8632 (I149290,I149273,I60442);
nand I_8633 (I149307,I149290,I60448);
nor I_8634 (I149324,I149307,I149256);
DFFARX1 I_8635 (I149324,I2507,I149106,I149074,);
not I_8636 (I149355,I149307);
not I_8637 (I149372,I60442);
nand I_8638 (I149389,I149372,I60436);
nor I_8639 (I149406,I60442,I60457);
nand I_8640 (I149086,I149222,I149406);
nand I_8641 (I149080,I149171,I60442);
nand I_8642 (I149451,I149273,I60436);
DFFARX1 I_8643 (I149451,I2507,I149106,I149095,);
DFFARX1 I_8644 (I149451,I2507,I149106,I149089,);
not I_8645 (I149496,I60436);
nor I_8646 (I149513,I149496,I60454);
and I_8647 (I149530,I149513,I60460);
or I_8648 (I149547,I149530,I60439);
DFFARX1 I_8649 (I149547,I2507,I149106,I149573,);
nand I_8650 (I149581,I149573,I149239);
nor I_8651 (I149083,I149581,I149389);
nor I_8652 (I149077,I149573,I149205);
DFFARX1 I_8653 (I149573,I2507,I149106,I149635,);
not I_8654 (I149643,I149635);
nor I_8655 (I149092,I149643,I149355);
not I_8656 (I149701,I2514);
DFFARX1 I_8657 (I713869,I2507,I149701,I149727,);
DFFARX1 I_8658 (I149727,I2507,I149701,I149744,);
not I_8659 (I149693,I149744);
not I_8660 (I149766,I149727);
DFFARX1 I_8661 (I713860,I2507,I149701,I149792,);
not I_8662 (I149800,I149792);
and I_8663 (I149817,I149766,I713854);
not I_8664 (I149834,I713848);
nand I_8665 (I149851,I149834,I713854);
not I_8666 (I149868,I713875);
nor I_8667 (I149885,I149868,I713848);
nand I_8668 (I149902,I149885,I713872);
nor I_8669 (I149919,I149902,I149851);
DFFARX1 I_8670 (I149919,I2507,I149701,I149669,);
not I_8671 (I149950,I149902);
not I_8672 (I149967,I713848);
nand I_8673 (I149984,I149967,I713854);
nor I_8674 (I150001,I713848,I713848);
nand I_8675 (I149681,I149817,I150001);
nand I_8676 (I149675,I149766,I713848);
nand I_8677 (I150046,I149868,I713857);
DFFARX1 I_8678 (I150046,I2507,I149701,I149690,);
DFFARX1 I_8679 (I150046,I2507,I149701,I149684,);
not I_8680 (I150091,I713857);
nor I_8681 (I150108,I150091,I713863);
and I_8682 (I150125,I150108,I713866);
or I_8683 (I150142,I150125,I713851);
DFFARX1 I_8684 (I150142,I2507,I149701,I150168,);
nand I_8685 (I150176,I150168,I149834);
nor I_8686 (I149678,I150176,I149984);
nor I_8687 (I149672,I150168,I149800);
DFFARX1 I_8688 (I150168,I2507,I149701,I150230,);
not I_8689 (I150238,I150230);
nor I_8690 (I149687,I150238,I149950);
not I_8691 (I150296,I2514);
DFFARX1 I_8692 (I590751,I2507,I150296,I150322,);
DFFARX1 I_8693 (I150322,I2507,I150296,I150339,);
not I_8694 (I150288,I150339);
not I_8695 (I150361,I150322);
DFFARX1 I_8696 (I590751,I2507,I150296,I150387,);
not I_8697 (I150395,I150387);
and I_8698 (I150412,I150361,I590754);
not I_8699 (I150429,I590766);
nand I_8700 (I150446,I150429,I590754);
not I_8701 (I150463,I590772);
nor I_8702 (I150480,I150463,I590763);
nand I_8703 (I150497,I150480,I590769);
nor I_8704 (I150514,I150497,I150446);
DFFARX1 I_8705 (I150514,I2507,I150296,I150264,);
not I_8706 (I150545,I150497);
not I_8707 (I150562,I590763);
nand I_8708 (I150579,I150562,I590754);
nor I_8709 (I150596,I590763,I590766);
nand I_8710 (I150276,I150412,I150596);
nand I_8711 (I150270,I150361,I590763);
nand I_8712 (I150641,I150463,I590760);
DFFARX1 I_8713 (I150641,I2507,I150296,I150285,);
DFFARX1 I_8714 (I150641,I2507,I150296,I150279,);
not I_8715 (I150686,I590760);
nor I_8716 (I150703,I150686,I590757);
and I_8717 (I150720,I150703,I590775);
or I_8718 (I150737,I150720,I590754);
DFFARX1 I_8719 (I150737,I2507,I150296,I150763,);
nand I_8720 (I150771,I150763,I150429);
nor I_8721 (I150273,I150771,I150579);
nor I_8722 (I150267,I150763,I150395);
DFFARX1 I_8723 (I150763,I2507,I150296,I150825,);
not I_8724 (I150833,I150825);
nor I_8725 (I150282,I150833,I150545);
not I_8726 (I150891,I2514);
DFFARX1 I_8727 (I540791,I2507,I150891,I150917,);
DFFARX1 I_8728 (I150917,I2507,I150891,I150934,);
not I_8729 (I150883,I150934);
not I_8730 (I150956,I150917);
DFFARX1 I_8731 (I540800,I2507,I150891,I150982,);
not I_8732 (I150990,I150982);
and I_8733 (I151007,I150956,I540794);
not I_8734 (I151024,I540788);
nand I_8735 (I151041,I151024,I540794);
not I_8736 (I151058,I540803);
nor I_8737 (I151075,I151058,I540791);
nand I_8738 (I151092,I151075,I540797);
nor I_8739 (I151109,I151092,I151041);
DFFARX1 I_8740 (I151109,I2507,I150891,I150859,);
not I_8741 (I151140,I151092);
not I_8742 (I151157,I540791);
nand I_8743 (I151174,I151157,I540794);
nor I_8744 (I151191,I540791,I540788);
nand I_8745 (I150871,I151007,I151191);
nand I_8746 (I150865,I150956,I540791);
nand I_8747 (I151236,I151058,I540794);
DFFARX1 I_8748 (I151236,I2507,I150891,I150880,);
DFFARX1 I_8749 (I151236,I2507,I150891,I150874,);
not I_8750 (I151281,I540794);
nor I_8751 (I151298,I151281,I540809);
and I_8752 (I151315,I151298,I540806);
or I_8753 (I151332,I151315,I540788);
DFFARX1 I_8754 (I151332,I2507,I150891,I151358,);
nand I_8755 (I151366,I151358,I151024);
nor I_8756 (I150868,I151366,I151174);
nor I_8757 (I150862,I151358,I150990);
DFFARX1 I_8758 (I151358,I2507,I150891,I151420,);
not I_8759 (I151428,I151420);
nor I_8760 (I150877,I151428,I151140);
not I_8761 (I151486,I2514);
DFFARX1 I_8762 (I52540,I2507,I151486,I151512,);
DFFARX1 I_8763 (I151512,I2507,I151486,I151529,);
not I_8764 (I151478,I151529);
not I_8765 (I151551,I151512);
DFFARX1 I_8766 (I52534,I2507,I151486,I151577,);
not I_8767 (I151585,I151577);
and I_8768 (I151602,I151551,I52531);
not I_8769 (I151619,I52552);
nand I_8770 (I151636,I151619,I52531);
not I_8771 (I151653,I52546);
nor I_8772 (I151670,I151653,I52537);
nand I_8773 (I151687,I151670,I52543);
nor I_8774 (I151704,I151687,I151636);
DFFARX1 I_8775 (I151704,I2507,I151486,I151454,);
not I_8776 (I151735,I151687);
not I_8777 (I151752,I52537);
nand I_8778 (I151769,I151752,I52531);
nor I_8779 (I151786,I52537,I52552);
nand I_8780 (I151466,I151602,I151786);
nand I_8781 (I151460,I151551,I52537);
nand I_8782 (I151831,I151653,I52531);
DFFARX1 I_8783 (I151831,I2507,I151486,I151475,);
DFFARX1 I_8784 (I151831,I2507,I151486,I151469,);
not I_8785 (I151876,I52531);
nor I_8786 (I151893,I151876,I52549);
and I_8787 (I151910,I151893,I52555);
or I_8788 (I151927,I151910,I52534);
DFFARX1 I_8789 (I151927,I2507,I151486,I151953,);
nand I_8790 (I151961,I151953,I151619);
nor I_8791 (I151463,I151961,I151769);
nor I_8792 (I151457,I151953,I151585);
DFFARX1 I_8793 (I151953,I2507,I151486,I152015,);
not I_8794 (I152023,I152015);
nor I_8795 (I151472,I152023,I151735);
not I_8796 (I152081,I2514);
DFFARX1 I_8797 (I327606,I2507,I152081,I152107,);
DFFARX1 I_8798 (I152107,I2507,I152081,I152124,);
not I_8799 (I152073,I152124);
not I_8800 (I152146,I152107);
DFFARX1 I_8801 (I327597,I2507,I152081,I152172,);
not I_8802 (I152180,I152172);
and I_8803 (I152197,I152146,I327615);
not I_8804 (I152214,I327612);
nand I_8805 (I152231,I152214,I327615);
not I_8806 (I152248,I327591);
nor I_8807 (I152265,I152248,I327594);
nand I_8808 (I152282,I152265,I327603);
nor I_8809 (I152299,I152282,I152231);
DFFARX1 I_8810 (I152299,I2507,I152081,I152049,);
not I_8811 (I152330,I152282);
not I_8812 (I152347,I327594);
nand I_8813 (I152364,I152347,I327615);
nor I_8814 (I152381,I327594,I327612);
nand I_8815 (I152061,I152197,I152381);
nand I_8816 (I152055,I152146,I327594);
nand I_8817 (I152426,I152248,I327609);
DFFARX1 I_8818 (I152426,I2507,I152081,I152070,);
DFFARX1 I_8819 (I152426,I2507,I152081,I152064,);
not I_8820 (I152471,I327609);
nor I_8821 (I152488,I152471,I327591);
and I_8822 (I152505,I152488,I327600);
or I_8823 (I152522,I152505,I327594);
DFFARX1 I_8824 (I152522,I2507,I152081,I152548,);
nand I_8825 (I152556,I152548,I152214);
nor I_8826 (I152058,I152556,I152364);
nor I_8827 (I152052,I152548,I152180);
DFFARX1 I_8828 (I152548,I2507,I152081,I152610,);
not I_8829 (I152618,I152610);
nor I_8830 (I152067,I152618,I152330);
not I_8831 (I152676,I2514);
DFFARX1 I_8832 (I283760,I2507,I152676,I152702,);
DFFARX1 I_8833 (I152702,I2507,I152676,I152719,);
not I_8834 (I152668,I152719);
not I_8835 (I152741,I152702);
DFFARX1 I_8836 (I283754,I2507,I152676,I152767,);
not I_8837 (I152775,I152767);
and I_8838 (I152792,I152741,I283769);
not I_8839 (I152809,I283766);
nand I_8840 (I152826,I152809,I283769);
not I_8841 (I152843,I283757);
nor I_8842 (I152860,I152843,I283748);
nand I_8843 (I152877,I152860,I283751);
nor I_8844 (I152894,I152877,I152826);
DFFARX1 I_8845 (I152894,I2507,I152676,I152644,);
not I_8846 (I152925,I152877);
not I_8847 (I152942,I283748);
nand I_8848 (I152959,I152942,I283769);
nor I_8849 (I152976,I283748,I283766);
nand I_8850 (I152656,I152792,I152976);
nand I_8851 (I152650,I152741,I283748);
nand I_8852 (I153021,I152843,I283772);
DFFARX1 I_8853 (I153021,I2507,I152676,I152665,);
DFFARX1 I_8854 (I153021,I2507,I152676,I152659,);
not I_8855 (I153066,I283772);
nor I_8856 (I153083,I153066,I283763);
and I_8857 (I153100,I153083,I283748);
or I_8858 (I153117,I153100,I283751);
DFFARX1 I_8859 (I153117,I2507,I152676,I153143,);
nand I_8860 (I153151,I153143,I152809);
nor I_8861 (I152653,I153151,I152959);
nor I_8862 (I152647,I153143,I152775);
DFFARX1 I_8863 (I153143,I2507,I152676,I153205,);
not I_8864 (I153213,I153205);
nor I_8865 (I152662,I153213,I152925);
not I_8866 (I153271,I2514);
DFFARX1 I_8867 (I398697,I2507,I153271,I153297,);
DFFARX1 I_8868 (I153297,I2507,I153271,I153314,);
not I_8869 (I153263,I153314);
not I_8870 (I153336,I153297);
DFFARX1 I_8871 (I398694,I2507,I153271,I153362,);
not I_8872 (I153370,I153362);
and I_8873 (I153387,I153336,I398700);
not I_8874 (I153404,I398685);
nand I_8875 (I153421,I153404,I398700);
not I_8876 (I153438,I398688);
nor I_8877 (I153455,I153438,I398709);
nand I_8878 (I153472,I153455,I398706);
nor I_8879 (I153489,I153472,I153421);
DFFARX1 I_8880 (I153489,I2507,I153271,I153239,);
not I_8881 (I153520,I153472);
not I_8882 (I153537,I398709);
nand I_8883 (I153554,I153537,I398700);
nor I_8884 (I153571,I398709,I398685);
nand I_8885 (I153251,I153387,I153571);
nand I_8886 (I153245,I153336,I398709);
nand I_8887 (I153616,I153438,I398685);
DFFARX1 I_8888 (I153616,I2507,I153271,I153260,);
DFFARX1 I_8889 (I153616,I2507,I153271,I153254,);
not I_8890 (I153661,I398685);
nor I_8891 (I153678,I153661,I398691);
and I_8892 (I153695,I153678,I398703);
or I_8893 (I153712,I153695,I398688);
DFFARX1 I_8894 (I153712,I2507,I153271,I153738,);
nand I_8895 (I153746,I153738,I153404);
nor I_8896 (I153248,I153746,I153554);
nor I_8897 (I153242,I153738,I153370);
DFFARX1 I_8898 (I153738,I2507,I153271,I153800,);
not I_8899 (I153808,I153800);
nor I_8900 (I153257,I153808,I153520);
not I_8901 (I153866,I2514);
DFFARX1 I_8902 (I636413,I2507,I153866,I153892,);
DFFARX1 I_8903 (I153892,I2507,I153866,I153909,);
not I_8904 (I153858,I153909);
not I_8905 (I153931,I153892);
DFFARX1 I_8906 (I636413,I2507,I153866,I153957,);
not I_8907 (I153965,I153957);
and I_8908 (I153982,I153931,I636416);
not I_8909 (I153999,I636428);
nand I_8910 (I154016,I153999,I636416);
not I_8911 (I154033,I636434);
nor I_8912 (I154050,I154033,I636425);
nand I_8913 (I154067,I154050,I636431);
nor I_8914 (I154084,I154067,I154016);
DFFARX1 I_8915 (I154084,I2507,I153866,I153834,);
not I_8916 (I154115,I154067);
not I_8917 (I154132,I636425);
nand I_8918 (I154149,I154132,I636416);
nor I_8919 (I154166,I636425,I636428);
nand I_8920 (I153846,I153982,I154166);
nand I_8921 (I153840,I153931,I636425);
nand I_8922 (I154211,I154033,I636422);
DFFARX1 I_8923 (I154211,I2507,I153866,I153855,);
DFFARX1 I_8924 (I154211,I2507,I153866,I153849,);
not I_8925 (I154256,I636422);
nor I_8926 (I154273,I154256,I636419);
and I_8927 (I154290,I154273,I636437);
or I_8928 (I154307,I154290,I636416);
DFFARX1 I_8929 (I154307,I2507,I153866,I154333,);
nand I_8930 (I154341,I154333,I153999);
nor I_8931 (I153843,I154341,I154149);
nor I_8932 (I153837,I154333,I153965);
DFFARX1 I_8933 (I154333,I2507,I153866,I154395,);
not I_8934 (I154403,I154395);
nor I_8935 (I153852,I154403,I154115);
not I_8936 (I154461,I2514);
DFFARX1 I_8937 (I350145,I2507,I154461,I154487,);
DFFARX1 I_8938 (I154487,I2507,I154461,I154504,);
not I_8939 (I154453,I154504);
not I_8940 (I154526,I154487);
DFFARX1 I_8941 (I350142,I2507,I154461,I154552,);
not I_8942 (I154560,I154552);
and I_8943 (I154577,I154526,I350148);
not I_8944 (I154594,I350133);
nand I_8945 (I154611,I154594,I350148);
not I_8946 (I154628,I350136);
nor I_8947 (I154645,I154628,I350157);
nand I_8948 (I154662,I154645,I350154);
nor I_8949 (I154679,I154662,I154611);
DFFARX1 I_8950 (I154679,I2507,I154461,I154429,);
not I_8951 (I154710,I154662);
not I_8952 (I154727,I350157);
nand I_8953 (I154744,I154727,I350148);
nor I_8954 (I154761,I350157,I350133);
nand I_8955 (I154441,I154577,I154761);
nand I_8956 (I154435,I154526,I350157);
nand I_8957 (I154806,I154628,I350133);
DFFARX1 I_8958 (I154806,I2507,I154461,I154450,);
DFFARX1 I_8959 (I154806,I2507,I154461,I154444,);
not I_8960 (I154851,I350133);
nor I_8961 (I154868,I154851,I350139);
and I_8962 (I154885,I154868,I350151);
or I_8963 (I154902,I154885,I350136);
DFFARX1 I_8964 (I154902,I2507,I154461,I154928,);
nand I_8965 (I154936,I154928,I154594);
nor I_8966 (I154438,I154936,I154744);
nor I_8967 (I154432,I154928,I154560);
DFFARX1 I_8968 (I154928,I2507,I154461,I154990,);
not I_8969 (I154998,I154990);
nor I_8970 (I154447,I154998,I154710);
not I_8971 (I155056,I2514);
DFFARX1 I_8972 (I269968,I2507,I155056,I155082,);
DFFARX1 I_8973 (I155082,I2507,I155056,I155099,);
not I_8974 (I155048,I155099);
not I_8975 (I155121,I155082);
DFFARX1 I_8976 (I269956,I2507,I155056,I155147,);
not I_8977 (I155155,I155147);
and I_8978 (I155172,I155121,I269965);
not I_8979 (I155189,I269962);
nand I_8980 (I155206,I155189,I269965);
not I_8981 (I155223,I269953);
nor I_8982 (I155240,I155223,I269959);
nand I_8983 (I155257,I155240,I269944);
nor I_8984 (I155274,I155257,I155206);
DFFARX1 I_8985 (I155274,I2507,I155056,I155024,);
not I_8986 (I155305,I155257);
not I_8987 (I155322,I269959);
nand I_8988 (I155339,I155322,I269965);
nor I_8989 (I155356,I269959,I269962);
nand I_8990 (I155036,I155172,I155356);
nand I_8991 (I155030,I155121,I269959);
nand I_8992 (I155401,I155223,I269944);
DFFARX1 I_8993 (I155401,I2507,I155056,I155045,);
DFFARX1 I_8994 (I155401,I2507,I155056,I155039,);
not I_8995 (I155446,I269944);
nor I_8996 (I155463,I155446,I269950);
and I_8997 (I155480,I155463,I269947);
or I_8998 (I155497,I155480,I269971);
DFFARX1 I_8999 (I155497,I2507,I155056,I155523,);
nand I_9000 (I155531,I155523,I155189);
nor I_9001 (I155033,I155531,I155339);
nor I_9002 (I155027,I155523,I155155);
DFFARX1 I_9003 (I155523,I2507,I155056,I155585,);
not I_9004 (I155593,I155585);
nor I_9005 (I155042,I155593,I155305);
not I_9006 (I155651,I2514);
DFFARX1 I_9007 (I587283,I2507,I155651,I155677,);
DFFARX1 I_9008 (I155677,I2507,I155651,I155694,);
not I_9009 (I155643,I155694);
not I_9010 (I155716,I155677);
DFFARX1 I_9011 (I587283,I2507,I155651,I155742,);
not I_9012 (I155750,I155742);
and I_9013 (I155767,I155716,I587286);
not I_9014 (I155784,I587298);
nand I_9015 (I155801,I155784,I587286);
not I_9016 (I155818,I587304);
nor I_9017 (I155835,I155818,I587295);
nand I_9018 (I155852,I155835,I587301);
nor I_9019 (I155869,I155852,I155801);
DFFARX1 I_9020 (I155869,I2507,I155651,I155619,);
not I_9021 (I155900,I155852);
not I_9022 (I155917,I587295);
nand I_9023 (I155934,I155917,I587286);
nor I_9024 (I155951,I587295,I587298);
nand I_9025 (I155631,I155767,I155951);
nand I_9026 (I155625,I155716,I587295);
nand I_9027 (I155996,I155818,I587292);
DFFARX1 I_9028 (I155996,I2507,I155651,I155640,);
DFFARX1 I_9029 (I155996,I2507,I155651,I155634,);
not I_9030 (I156041,I587292);
nor I_9031 (I156058,I156041,I587289);
and I_9032 (I156075,I156058,I587307);
or I_9033 (I156092,I156075,I587286);
DFFARX1 I_9034 (I156092,I2507,I155651,I156118,);
nand I_9035 (I156126,I156118,I155784);
nor I_9036 (I155628,I156126,I155934);
nor I_9037 (I155622,I156118,I155750);
DFFARX1 I_9038 (I156118,I2507,I155651,I156180,);
not I_9039 (I156188,I156180);
nor I_9040 (I155637,I156188,I155900);
not I_9041 (I156246,I2514);
DFFARX1 I_9042 (I7760,I2507,I156246,I156272,);
DFFARX1 I_9043 (I156272,I2507,I156246,I156289,);
not I_9044 (I156238,I156289);
not I_9045 (I156311,I156272);
DFFARX1 I_9046 (I7736,I2507,I156246,I156337,);
not I_9047 (I156345,I156337);
and I_9048 (I156362,I156311,I7751);
not I_9049 (I156379,I7739);
nand I_9050 (I156396,I156379,I7751);
not I_9051 (I156413,I7742);
nor I_9052 (I156430,I156413,I7754);
nand I_9053 (I156447,I156430,I7745);
nor I_9054 (I156464,I156447,I156396);
DFFARX1 I_9055 (I156464,I2507,I156246,I156214,);
not I_9056 (I156495,I156447);
not I_9057 (I156512,I7754);
nand I_9058 (I156529,I156512,I7751);
nor I_9059 (I156546,I7754,I7739);
nand I_9060 (I156226,I156362,I156546);
nand I_9061 (I156220,I156311,I7754);
nand I_9062 (I156591,I156413,I7748);
DFFARX1 I_9063 (I156591,I2507,I156246,I156235,);
DFFARX1 I_9064 (I156591,I2507,I156246,I156229,);
not I_9065 (I156636,I7748);
nor I_9066 (I156653,I156636,I7739);
and I_9067 (I156670,I156653,I7736);
or I_9068 (I156687,I156670,I7757);
DFFARX1 I_9069 (I156687,I2507,I156246,I156713,);
nand I_9070 (I156721,I156713,I156379);
nor I_9071 (I156223,I156721,I156529);
nor I_9072 (I156217,I156713,I156345);
DFFARX1 I_9073 (I156713,I2507,I156246,I156775,);
not I_9074 (I156783,I156775);
nor I_9075 (I156232,I156783,I156495);
not I_9076 (I156841,I2514);
DFFARX1 I_9077 (I235152,I2507,I156841,I156867,);
DFFARX1 I_9078 (I156867,I2507,I156841,I156884,);
not I_9079 (I156833,I156884);
not I_9080 (I156906,I156867);
DFFARX1 I_9081 (I235140,I2507,I156841,I156932,);
not I_9082 (I156940,I156932);
and I_9083 (I156957,I156906,I235149);
not I_9084 (I156974,I235146);
nand I_9085 (I156991,I156974,I235149);
not I_9086 (I157008,I235137);
nor I_9087 (I157025,I157008,I235143);
nand I_9088 (I157042,I157025,I235128);
nor I_9089 (I157059,I157042,I156991);
DFFARX1 I_9090 (I157059,I2507,I156841,I156809,);
not I_9091 (I157090,I157042);
not I_9092 (I157107,I235143);
nand I_9093 (I157124,I157107,I235149);
nor I_9094 (I157141,I235143,I235146);
nand I_9095 (I156821,I156957,I157141);
nand I_9096 (I156815,I156906,I235143);
nand I_9097 (I157186,I157008,I235128);
DFFARX1 I_9098 (I157186,I2507,I156841,I156830,);
DFFARX1 I_9099 (I157186,I2507,I156841,I156824,);
not I_9100 (I157231,I235128);
nor I_9101 (I157248,I157231,I235134);
and I_9102 (I157265,I157248,I235131);
or I_9103 (I157282,I157265,I235155);
DFFARX1 I_9104 (I157282,I2507,I156841,I157308,);
nand I_9105 (I157316,I157308,I156974);
nor I_9106 (I156818,I157316,I157124);
nor I_9107 (I156812,I157308,I156940);
DFFARX1 I_9108 (I157308,I2507,I156841,I157370,);
not I_9109 (I157378,I157370);
nor I_9110 (I156827,I157378,I157090);
not I_9111 (I157436,I2514);
DFFARX1 I_9112 (I201689,I2507,I157436,I157462,);
DFFARX1 I_9113 (I157462,I2507,I157436,I157479,);
not I_9114 (I157428,I157479);
not I_9115 (I157501,I157462);
DFFARX1 I_9116 (I201704,I2507,I157436,I157527,);
not I_9117 (I157535,I157527);
and I_9118 (I157552,I157501,I201701);
not I_9119 (I157569,I201689);
nand I_9120 (I157586,I157569,I201701);
not I_9121 (I157603,I201698);
nor I_9122 (I157620,I157603,I201713);
nand I_9123 (I157637,I157620,I201710);
nor I_9124 (I157654,I157637,I157586);
DFFARX1 I_9125 (I157654,I2507,I157436,I157404,);
not I_9126 (I157685,I157637);
not I_9127 (I157702,I201713);
nand I_9128 (I157719,I157702,I201701);
nor I_9129 (I157736,I201713,I201689);
nand I_9130 (I157416,I157552,I157736);
nand I_9131 (I157410,I157501,I201713);
nand I_9132 (I157781,I157603,I201707);
DFFARX1 I_9133 (I157781,I2507,I157436,I157425,);
DFFARX1 I_9134 (I157781,I2507,I157436,I157419,);
not I_9135 (I157826,I201707);
nor I_9136 (I157843,I157826,I201695);
and I_9137 (I157860,I157843,I201716);
or I_9138 (I157877,I157860,I201692);
DFFARX1 I_9139 (I157877,I2507,I157436,I157903,);
nand I_9140 (I157911,I157903,I157569);
nor I_9141 (I157413,I157911,I157719);
nor I_9142 (I157407,I157903,I157535);
DFFARX1 I_9143 (I157903,I2507,I157436,I157965,);
not I_9144 (I157973,I157965);
nor I_9145 (I157422,I157973,I157685);
not I_9146 (I158031,I2514);
DFFARX1 I_9147 (I169542,I2507,I158031,I158057,);
DFFARX1 I_9148 (I158057,I2507,I158031,I158074,);
not I_9149 (I158023,I158074);
not I_9150 (I158096,I158057);
DFFARX1 I_9151 (I169557,I2507,I158031,I158122,);
not I_9152 (I158130,I158122);
and I_9153 (I158147,I158096,I169554);
not I_9154 (I158164,I169542);
nand I_9155 (I158181,I158164,I169554);
not I_9156 (I158198,I169551);
nor I_9157 (I158215,I158198,I169566);
nand I_9158 (I158232,I158215,I169563);
nor I_9159 (I158249,I158232,I158181);
DFFARX1 I_9160 (I158249,I2507,I158031,I157999,);
not I_9161 (I158280,I158232);
not I_9162 (I158297,I169566);
nand I_9163 (I158314,I158297,I169554);
nor I_9164 (I158331,I169566,I169542);
nand I_9165 (I158011,I158147,I158331);
nand I_9166 (I158005,I158096,I169566);
nand I_9167 (I158376,I158198,I169560);
DFFARX1 I_9168 (I158376,I2507,I158031,I158020,);
DFFARX1 I_9169 (I158376,I2507,I158031,I158014,);
not I_9170 (I158421,I169560);
nor I_9171 (I158438,I158421,I169548);
and I_9172 (I158455,I158438,I169569);
or I_9173 (I158472,I158455,I169545);
DFFARX1 I_9174 (I158472,I2507,I158031,I158498,);
nand I_9175 (I158506,I158498,I158164);
nor I_9176 (I158008,I158506,I158314);
nor I_9177 (I158002,I158498,I158130);
DFFARX1 I_9178 (I158498,I2507,I158031,I158560,);
not I_9179 (I158568,I158560);
nor I_9180 (I158017,I158568,I158280);
not I_9181 (I158626,I2514);
DFFARX1 I_9182 (I54121,I2507,I158626,I158652,);
DFFARX1 I_9183 (I158652,I2507,I158626,I158669,);
not I_9184 (I158618,I158669);
not I_9185 (I158691,I158652);
DFFARX1 I_9186 (I54115,I2507,I158626,I158717,);
not I_9187 (I158725,I158717);
and I_9188 (I158742,I158691,I54112);
not I_9189 (I158759,I54133);
nand I_9190 (I158776,I158759,I54112);
not I_9191 (I158793,I54127);
nor I_9192 (I158810,I158793,I54118);
nand I_9193 (I158827,I158810,I54124);
nor I_9194 (I158844,I158827,I158776);
DFFARX1 I_9195 (I158844,I2507,I158626,I158594,);
not I_9196 (I158875,I158827);
not I_9197 (I158892,I54118);
nand I_9198 (I158909,I158892,I54112);
nor I_9199 (I158926,I54118,I54133);
nand I_9200 (I158606,I158742,I158926);
nand I_9201 (I158600,I158691,I54118);
nand I_9202 (I158971,I158793,I54112);
DFFARX1 I_9203 (I158971,I2507,I158626,I158615,);
DFFARX1 I_9204 (I158971,I2507,I158626,I158609,);
not I_9205 (I159016,I54112);
nor I_9206 (I159033,I159016,I54130);
and I_9207 (I159050,I159033,I54136);
or I_9208 (I159067,I159050,I54115);
DFFARX1 I_9209 (I159067,I2507,I158626,I159093,);
nand I_9210 (I159101,I159093,I158759);
nor I_9211 (I158603,I159101,I158909);
nor I_9212 (I158597,I159093,I158725);
DFFARX1 I_9213 (I159093,I2507,I158626,I159155,);
not I_9214 (I159163,I159155);
nor I_9215 (I158612,I159163,I158875);
not I_9216 (I159221,I2514);
DFFARX1 I_9217 (I447090,I2507,I159221,I159247,);
DFFARX1 I_9218 (I159247,I2507,I159221,I159264,);
not I_9219 (I159213,I159264);
not I_9220 (I159286,I159247);
DFFARX1 I_9221 (I447084,I2507,I159221,I159312,);
not I_9222 (I159320,I159312);
and I_9223 (I159337,I159286,I447102);
not I_9224 (I159354,I447090);
nand I_9225 (I159371,I159354,I447102);
not I_9226 (I159388,I447084);
nor I_9227 (I159405,I159388,I447096);
nand I_9228 (I159422,I159405,I447087);
nor I_9229 (I159439,I159422,I159371);
DFFARX1 I_9230 (I159439,I2507,I159221,I159189,);
not I_9231 (I159470,I159422);
not I_9232 (I159487,I447096);
nand I_9233 (I159504,I159487,I447102);
nor I_9234 (I159521,I447096,I447090);
nand I_9235 (I159201,I159337,I159521);
nand I_9236 (I159195,I159286,I447096);
nand I_9237 (I159566,I159388,I447099);
DFFARX1 I_9238 (I159566,I2507,I159221,I159210,);
DFFARX1 I_9239 (I159566,I2507,I159221,I159204,);
not I_9240 (I159611,I447099);
nor I_9241 (I159628,I159611,I447105);
and I_9242 (I159645,I159628,I447087);
or I_9243 (I159662,I159645,I447093);
DFFARX1 I_9244 (I159662,I2507,I159221,I159688,);
nand I_9245 (I159696,I159688,I159354);
nor I_9246 (I159198,I159696,I159504);
nor I_9247 (I159192,I159688,I159320);
DFFARX1 I_9248 (I159688,I2507,I159221,I159750,);
not I_9249 (I159758,I159750);
nor I_9250 (I159207,I159758,I159470);
not I_9251 (I159816,I2514);
DFFARX1 I_9252 (I64661,I2507,I159816,I159842,);
DFFARX1 I_9253 (I159842,I2507,I159816,I159859,);
not I_9254 (I159808,I159859);
not I_9255 (I159881,I159842);
DFFARX1 I_9256 (I64655,I2507,I159816,I159907,);
not I_9257 (I159915,I159907);
and I_9258 (I159932,I159881,I64652);
not I_9259 (I159949,I64673);
nand I_9260 (I159966,I159949,I64652);
not I_9261 (I159983,I64667);
nor I_9262 (I160000,I159983,I64658);
nand I_9263 (I160017,I160000,I64664);
nor I_9264 (I160034,I160017,I159966);
DFFARX1 I_9265 (I160034,I2507,I159816,I159784,);
not I_9266 (I160065,I160017);
not I_9267 (I160082,I64658);
nand I_9268 (I160099,I160082,I64652);
nor I_9269 (I160116,I64658,I64673);
nand I_9270 (I159796,I159932,I160116);
nand I_9271 (I159790,I159881,I64658);
nand I_9272 (I160161,I159983,I64652);
DFFARX1 I_9273 (I160161,I2507,I159816,I159805,);
DFFARX1 I_9274 (I160161,I2507,I159816,I159799,);
not I_9275 (I160206,I64652);
nor I_9276 (I160223,I160206,I64670);
and I_9277 (I160240,I160223,I64676);
or I_9278 (I160257,I160240,I64655);
DFFARX1 I_9279 (I160257,I2507,I159816,I160283,);
nand I_9280 (I160291,I160283,I159949);
nor I_9281 (I159793,I160291,I160099);
nor I_9282 (I159787,I160283,I159915);
DFFARX1 I_9283 (I160283,I2507,I159816,I160345,);
not I_9284 (I160353,I160345);
nor I_9285 (I159802,I160353,I160065);
not I_9286 (I160411,I2514);
DFFARX1 I_9287 (I351879,I2507,I160411,I160437,);
DFFARX1 I_9288 (I160437,I2507,I160411,I160454,);
not I_9289 (I160403,I160454);
not I_9290 (I160476,I160437);
DFFARX1 I_9291 (I351876,I2507,I160411,I160502,);
not I_9292 (I160510,I160502);
and I_9293 (I160527,I160476,I351882);
not I_9294 (I160544,I351867);
nand I_9295 (I160561,I160544,I351882);
not I_9296 (I160578,I351870);
nor I_9297 (I160595,I160578,I351891);
nand I_9298 (I160612,I160595,I351888);
nor I_9299 (I160629,I160612,I160561);
DFFARX1 I_9300 (I160629,I2507,I160411,I160379,);
not I_9301 (I160660,I160612);
not I_9302 (I160677,I351891);
nand I_9303 (I160694,I160677,I351882);
nor I_9304 (I160711,I351891,I351867);
nand I_9305 (I160391,I160527,I160711);
nand I_9306 (I160385,I160476,I351891);
nand I_9307 (I160756,I160578,I351867);
DFFARX1 I_9308 (I160756,I2507,I160411,I160400,);
DFFARX1 I_9309 (I160756,I2507,I160411,I160394,);
not I_9310 (I160801,I351867);
nor I_9311 (I160818,I160801,I351873);
and I_9312 (I160835,I160818,I351885);
or I_9313 (I160852,I160835,I351870);
DFFARX1 I_9314 (I160852,I2507,I160411,I160878,);
nand I_9315 (I160886,I160878,I160544);
nor I_9316 (I160388,I160886,I160694);
nor I_9317 (I160382,I160878,I160510);
DFFARX1 I_9318 (I160878,I2507,I160411,I160940,);
not I_9319 (I160948,I160940);
nor I_9320 (I160397,I160948,I160660);
not I_9321 (I161006,I2514);
DFFARX1 I_9322 (I41473,I2507,I161006,I161032,);
DFFARX1 I_9323 (I161032,I2507,I161006,I161049,);
not I_9324 (I160998,I161049);
not I_9325 (I161071,I161032);
DFFARX1 I_9326 (I41467,I2507,I161006,I161097,);
not I_9327 (I161105,I161097);
and I_9328 (I161122,I161071,I41464);
not I_9329 (I161139,I41485);
nand I_9330 (I161156,I161139,I41464);
not I_9331 (I161173,I41479);
nor I_9332 (I161190,I161173,I41470);
nand I_9333 (I161207,I161190,I41476);
nor I_9334 (I161224,I161207,I161156);
DFFARX1 I_9335 (I161224,I2507,I161006,I160974,);
not I_9336 (I161255,I161207);
not I_9337 (I161272,I41470);
nand I_9338 (I161289,I161272,I41464);
nor I_9339 (I161306,I41470,I41485);
nand I_9340 (I160986,I161122,I161306);
nand I_9341 (I160980,I161071,I41470);
nand I_9342 (I161351,I161173,I41464);
DFFARX1 I_9343 (I161351,I2507,I161006,I160995,);
DFFARX1 I_9344 (I161351,I2507,I161006,I160989,);
not I_9345 (I161396,I41464);
nor I_9346 (I161413,I161396,I41482);
and I_9347 (I161430,I161413,I41488);
or I_9348 (I161447,I161430,I41467);
DFFARX1 I_9349 (I161447,I2507,I161006,I161473,);
nand I_9350 (I161481,I161473,I161139);
nor I_9351 (I160983,I161481,I161289);
nor I_9352 (I160977,I161473,I161105);
DFFARX1 I_9353 (I161473,I2507,I161006,I161535,);
not I_9354 (I161543,I161535);
nor I_9355 (I160992,I161543,I161255);
not I_9356 (I161601,I2514);
DFFARX1 I_9357 (I706729,I2507,I161601,I161627,);
DFFARX1 I_9358 (I161627,I2507,I161601,I161644,);
not I_9359 (I161593,I161644);
not I_9360 (I161666,I161627);
DFFARX1 I_9361 (I706720,I2507,I161601,I161692,);
not I_9362 (I161700,I161692);
and I_9363 (I161717,I161666,I706714);
not I_9364 (I161734,I706708);
nand I_9365 (I161751,I161734,I706714);
not I_9366 (I161768,I706735);
nor I_9367 (I161785,I161768,I706708);
nand I_9368 (I161802,I161785,I706732);
nor I_9369 (I161819,I161802,I161751);
DFFARX1 I_9370 (I161819,I2507,I161601,I161569,);
not I_9371 (I161850,I161802);
not I_9372 (I161867,I706708);
nand I_9373 (I161884,I161867,I706714);
nor I_9374 (I161901,I706708,I706708);
nand I_9375 (I161581,I161717,I161901);
nand I_9376 (I161575,I161666,I706708);
nand I_9377 (I161946,I161768,I706717);
DFFARX1 I_9378 (I161946,I2507,I161601,I161590,);
DFFARX1 I_9379 (I161946,I2507,I161601,I161584,);
not I_9380 (I161991,I706717);
nor I_9381 (I162008,I161991,I706723);
and I_9382 (I162025,I162008,I706726);
or I_9383 (I162042,I162025,I706711);
DFFARX1 I_9384 (I162042,I2507,I161601,I162068,);
nand I_9385 (I162076,I162068,I161734);
nor I_9386 (I161578,I162076,I161884);
nor I_9387 (I161572,I162068,I161700);
DFFARX1 I_9388 (I162068,I2507,I161601,I162130,);
not I_9389 (I162138,I162130);
nor I_9390 (I161587,I162138,I161850);
not I_9391 (I162199,I2514);
DFFARX1 I_9392 (I263428,I2507,I162199,I162225,);
nand I_9393 (I162233,I263440,I263419);
and I_9394 (I162250,I162233,I263443);
DFFARX1 I_9395 (I162250,I2507,I162199,I162276,);
nor I_9396 (I162167,I162276,I162225);
not I_9397 (I162298,I162276);
DFFARX1 I_9398 (I263434,I2507,I162199,I162324,);
nand I_9399 (I162332,I162324,I263416);
not I_9400 (I162349,I162332);
DFFARX1 I_9401 (I162349,I2507,I162199,I162375,);
not I_9402 (I162191,I162375);
nor I_9403 (I162397,I162225,I162332);
nor I_9404 (I162173,I162276,I162397);
DFFARX1 I_9405 (I263431,I2507,I162199,I162437,);
DFFARX1 I_9406 (I162437,I2507,I162199,I162454,);
not I_9407 (I162462,I162454);
not I_9408 (I162479,I162437);
nand I_9409 (I162176,I162479,I162298);
nand I_9410 (I162510,I263416,I263422);
and I_9411 (I162527,I162510,I263425);
DFFARX1 I_9412 (I162527,I2507,I162199,I162553,);
nor I_9413 (I162561,I162553,I162225);
DFFARX1 I_9414 (I162561,I2507,I162199,I162164,);
DFFARX1 I_9415 (I162553,I2507,I162199,I162182,);
nor I_9416 (I162606,I263437,I263422);
not I_9417 (I162623,I162606);
nor I_9418 (I162185,I162462,I162623);
nand I_9419 (I162170,I162479,I162623);
nor I_9420 (I162179,I162225,I162606);
DFFARX1 I_9421 (I162606,I2507,I162199,I162188,);
not I_9422 (I162726,I2514);
DFFARX1 I_9423 (I393495,I2507,I162726,I162752,);
nand I_9424 (I162760,I393486,I393501);
and I_9425 (I162777,I162760,I393507);
DFFARX1 I_9426 (I162777,I2507,I162726,I162803,);
nor I_9427 (I162694,I162803,I162752);
not I_9428 (I162825,I162803);
DFFARX1 I_9429 (I393492,I2507,I162726,I162851,);
nand I_9430 (I162859,I162851,I393486);
not I_9431 (I162876,I162859);
DFFARX1 I_9432 (I162876,I2507,I162726,I162902,);
not I_9433 (I162718,I162902);
nor I_9434 (I162924,I162752,I162859);
nor I_9435 (I162700,I162803,I162924);
DFFARX1 I_9436 (I393489,I2507,I162726,I162964,);
DFFARX1 I_9437 (I162964,I2507,I162726,I162981,);
not I_9438 (I162989,I162981);
not I_9439 (I163006,I162964);
nand I_9440 (I162703,I163006,I162825);
nand I_9441 (I163037,I393483,I393498);
and I_9442 (I163054,I163037,I393483);
DFFARX1 I_9443 (I163054,I2507,I162726,I163080,);
nor I_9444 (I163088,I163080,I162752);
DFFARX1 I_9445 (I163088,I2507,I162726,I162691,);
DFFARX1 I_9446 (I163080,I2507,I162726,I162709,);
nor I_9447 (I163133,I393504,I393498);
not I_9448 (I163150,I163133);
nor I_9449 (I162712,I162989,I163150);
nand I_9450 (I162697,I163006,I163150);
nor I_9451 (I162706,I162752,I163133);
DFFARX1 I_9452 (I163133,I2507,I162726,I162715,);
not I_9453 (I163253,I2514);
DFFARX1 I_9454 (I401587,I2507,I163253,I163279,);
nand I_9455 (I163287,I401578,I401593);
and I_9456 (I163304,I163287,I401599);
DFFARX1 I_9457 (I163304,I2507,I163253,I163330,);
nor I_9458 (I163221,I163330,I163279);
not I_9459 (I163352,I163330);
DFFARX1 I_9460 (I401584,I2507,I163253,I163378,);
nand I_9461 (I163386,I163378,I401578);
not I_9462 (I163403,I163386);
DFFARX1 I_9463 (I163403,I2507,I163253,I163429,);
not I_9464 (I163245,I163429);
nor I_9465 (I163451,I163279,I163386);
nor I_9466 (I163227,I163330,I163451);
DFFARX1 I_9467 (I401581,I2507,I163253,I163491,);
DFFARX1 I_9468 (I163491,I2507,I163253,I163508,);
not I_9469 (I163516,I163508);
not I_9470 (I163533,I163491);
nand I_9471 (I163230,I163533,I163352);
nand I_9472 (I163564,I401575,I401590);
and I_9473 (I163581,I163564,I401575);
DFFARX1 I_9474 (I163581,I2507,I163253,I163607,);
nor I_9475 (I163615,I163607,I163279);
DFFARX1 I_9476 (I163615,I2507,I163253,I163218,);
DFFARX1 I_9477 (I163607,I2507,I163253,I163236,);
nor I_9478 (I163660,I401596,I401590);
not I_9479 (I163677,I163660);
nor I_9480 (I163239,I163516,I163677);
nand I_9481 (I163224,I163533,I163677);
nor I_9482 (I163233,I163279,I163660);
DFFARX1 I_9483 (I163660,I2507,I163253,I163242,);
not I_9484 (I163780,I2514);
DFFARX1 I_9485 (I409101,I2507,I163780,I163806,);
nand I_9486 (I163814,I409092,I409107);
and I_9487 (I163831,I163814,I409113);
DFFARX1 I_9488 (I163831,I2507,I163780,I163857,);
nor I_9489 (I163748,I163857,I163806);
not I_9490 (I163879,I163857);
DFFARX1 I_9491 (I409098,I2507,I163780,I163905,);
nand I_9492 (I163913,I163905,I409092);
not I_9493 (I163930,I163913);
DFFARX1 I_9494 (I163930,I2507,I163780,I163956,);
not I_9495 (I163772,I163956);
nor I_9496 (I163978,I163806,I163913);
nor I_9497 (I163754,I163857,I163978);
DFFARX1 I_9498 (I409095,I2507,I163780,I164018,);
DFFARX1 I_9499 (I164018,I2507,I163780,I164035,);
not I_9500 (I164043,I164035);
not I_9501 (I164060,I164018);
nand I_9502 (I163757,I164060,I163879);
nand I_9503 (I164091,I409089,I409104);
and I_9504 (I164108,I164091,I409089);
DFFARX1 I_9505 (I164108,I2507,I163780,I164134,);
nor I_9506 (I164142,I164134,I163806);
DFFARX1 I_9507 (I164142,I2507,I163780,I163745,);
DFFARX1 I_9508 (I164134,I2507,I163780,I163763,);
nor I_9509 (I164187,I409110,I409104);
not I_9510 (I164204,I164187);
nor I_9511 (I163766,I164043,I164204);
nand I_9512 (I163751,I164060,I164204);
nor I_9513 (I163760,I163806,I164187);
DFFARX1 I_9514 (I164187,I2507,I163780,I163769,);
not I_9515 (I164307,I2514);
DFFARX1 I_9516 (I240036,I2507,I164307,I164333,);
nand I_9517 (I164341,I240048,I240027);
and I_9518 (I164358,I164341,I240051);
DFFARX1 I_9519 (I164358,I2507,I164307,I164384,);
nor I_9520 (I164275,I164384,I164333);
not I_9521 (I164406,I164384);
DFFARX1 I_9522 (I240042,I2507,I164307,I164432,);
nand I_9523 (I164440,I164432,I240024);
not I_9524 (I164457,I164440);
DFFARX1 I_9525 (I164457,I2507,I164307,I164483,);
not I_9526 (I164299,I164483);
nor I_9527 (I164505,I164333,I164440);
nor I_9528 (I164281,I164384,I164505);
DFFARX1 I_9529 (I240039,I2507,I164307,I164545,);
DFFARX1 I_9530 (I164545,I2507,I164307,I164562,);
not I_9531 (I164570,I164562);
not I_9532 (I164587,I164545);
nand I_9533 (I164284,I164587,I164406);
nand I_9534 (I164618,I240024,I240030);
and I_9535 (I164635,I164618,I240033);
DFFARX1 I_9536 (I164635,I2507,I164307,I164661,);
nor I_9537 (I164669,I164661,I164333);
DFFARX1 I_9538 (I164669,I2507,I164307,I164272,);
DFFARX1 I_9539 (I164661,I2507,I164307,I164290,);
nor I_9540 (I164714,I240045,I240030);
not I_9541 (I164731,I164714);
nor I_9542 (I164293,I164570,I164731);
nand I_9543 (I164278,I164587,I164731);
nor I_9544 (I164287,I164333,I164714);
DFFARX1 I_9545 (I164714,I2507,I164307,I164296,);
not I_9546 (I164834,I2514);
DFFARX1 I_9547 (I234052,I2507,I164834,I164860,);
nand I_9548 (I164868,I234064,I234043);
and I_9549 (I164885,I164868,I234067);
DFFARX1 I_9550 (I164885,I2507,I164834,I164911,);
nor I_9551 (I164802,I164911,I164860);
not I_9552 (I164933,I164911);
DFFARX1 I_9553 (I234058,I2507,I164834,I164959,);
nand I_9554 (I164967,I164959,I234040);
not I_9555 (I164984,I164967);
DFFARX1 I_9556 (I164984,I2507,I164834,I165010,);
not I_9557 (I164826,I165010);
nor I_9558 (I165032,I164860,I164967);
nor I_9559 (I164808,I164911,I165032);
DFFARX1 I_9560 (I234055,I2507,I164834,I165072,);
DFFARX1 I_9561 (I165072,I2507,I164834,I165089,);
not I_9562 (I165097,I165089);
not I_9563 (I165114,I165072);
nand I_9564 (I164811,I165114,I164933);
nand I_9565 (I165145,I234040,I234046);
and I_9566 (I165162,I165145,I234049);
DFFARX1 I_9567 (I165162,I2507,I164834,I165188,);
nor I_9568 (I165196,I165188,I164860);
DFFARX1 I_9569 (I165196,I2507,I164834,I164799,);
DFFARX1 I_9570 (I165188,I2507,I164834,I164817,);
nor I_9571 (I165241,I234061,I234046);
not I_9572 (I165258,I165241);
nor I_9573 (I164820,I165097,I165258);
nand I_9574 (I164805,I165114,I165258);
nor I_9575 (I164814,I164860,I165241);
DFFARX1 I_9576 (I165241,I2507,I164834,I164823,);
not I_9577 (I165361,I2514);
DFFARX1 I_9578 (I109209,I2507,I165361,I165387,);
nand I_9579 (I165395,I109209,I109215);
and I_9580 (I165412,I165395,I109233);
DFFARX1 I_9581 (I165412,I2507,I165361,I165438,);
nor I_9582 (I165329,I165438,I165387);
not I_9583 (I165460,I165438);
DFFARX1 I_9584 (I109221,I2507,I165361,I165486,);
nand I_9585 (I165494,I165486,I109218);
not I_9586 (I165511,I165494);
DFFARX1 I_9587 (I165511,I2507,I165361,I165537,);
not I_9588 (I165353,I165537);
nor I_9589 (I165559,I165387,I165494);
nor I_9590 (I165335,I165438,I165559);
DFFARX1 I_9591 (I109227,I2507,I165361,I165599,);
DFFARX1 I_9592 (I165599,I2507,I165361,I165616,);
not I_9593 (I165624,I165616);
not I_9594 (I165641,I165599);
nand I_9595 (I165338,I165641,I165460);
nand I_9596 (I165672,I109212,I109212);
and I_9597 (I165689,I165672,I109224);
DFFARX1 I_9598 (I165689,I2507,I165361,I165715,);
nor I_9599 (I165723,I165715,I165387);
DFFARX1 I_9600 (I165723,I2507,I165361,I165326,);
DFFARX1 I_9601 (I165715,I2507,I165361,I165344,);
nor I_9602 (I165768,I109230,I109212);
not I_9603 (I165785,I165768);
nor I_9604 (I165347,I165624,I165785);
nand I_9605 (I165332,I165641,I165785);
nor I_9606 (I165341,I165387,I165768);
DFFARX1 I_9607 (I165768,I2507,I165361,I165350,);
not I_9608 (I165888,I2514);
DFFARX1 I_9609 (I286131,I2507,I165888,I165914,);
nand I_9610 (I165922,I286131,I286143);
and I_9611 (I165939,I165922,I286128);
DFFARX1 I_9612 (I165939,I2507,I165888,I165965,);
nor I_9613 (I165856,I165965,I165914);
not I_9614 (I165987,I165965);
DFFARX1 I_9615 (I286152,I2507,I165888,I166013,);
nand I_9616 (I166021,I166013,I286149);
not I_9617 (I166038,I166021);
DFFARX1 I_9618 (I166038,I2507,I165888,I166064,);
not I_9619 (I165880,I166064);
nor I_9620 (I166086,I165914,I166021);
nor I_9621 (I165862,I165965,I166086);
DFFARX1 I_9622 (I286140,I2507,I165888,I166126,);
DFFARX1 I_9623 (I166126,I2507,I165888,I166143,);
not I_9624 (I166151,I166143);
not I_9625 (I166168,I166126);
nand I_9626 (I165865,I166168,I165987);
nand I_9627 (I166199,I286128,I286137);
and I_9628 (I166216,I166199,I286146);
DFFARX1 I_9629 (I166216,I2507,I165888,I166242,);
nor I_9630 (I166250,I166242,I165914);
DFFARX1 I_9631 (I166250,I2507,I165888,I165853,);
DFFARX1 I_9632 (I166242,I2507,I165888,I165871,);
nor I_9633 (I166295,I286134,I286137);
not I_9634 (I166312,I166295);
nor I_9635 (I165874,I166151,I166312);
nand I_9636 (I165859,I166168,I166312);
nor I_9637 (I165868,I165914,I166295);
DFFARX1 I_9638 (I166295,I2507,I165888,I165877,);
not I_9639 (I166415,I2514);
DFFARX1 I_9640 (I247108,I2507,I166415,I166441,);
nand I_9641 (I166449,I247120,I247099);
and I_9642 (I166466,I166449,I247123);
DFFARX1 I_9643 (I166466,I2507,I166415,I166492,);
nor I_9644 (I166383,I166492,I166441);
not I_9645 (I166514,I166492);
DFFARX1 I_9646 (I247114,I2507,I166415,I166540,);
nand I_9647 (I166548,I166540,I247096);
not I_9648 (I166565,I166548);
DFFARX1 I_9649 (I166565,I2507,I166415,I166591,);
not I_9650 (I166407,I166591);
nor I_9651 (I166613,I166441,I166548);
nor I_9652 (I166389,I166492,I166613);
DFFARX1 I_9653 (I247111,I2507,I166415,I166653,);
DFFARX1 I_9654 (I166653,I2507,I166415,I166670,);
not I_9655 (I166678,I166670);
not I_9656 (I166695,I166653);
nand I_9657 (I166392,I166695,I166514);
nand I_9658 (I166726,I247096,I247102);
and I_9659 (I166743,I166726,I247105);
DFFARX1 I_9660 (I166743,I2507,I166415,I166769,);
nor I_9661 (I166777,I166769,I166441);
DFFARX1 I_9662 (I166777,I2507,I166415,I166380,);
DFFARX1 I_9663 (I166769,I2507,I166415,I166398,);
nor I_9664 (I166822,I247117,I247102);
not I_9665 (I166839,I166822);
nor I_9666 (I166401,I166678,I166839);
nand I_9667 (I166386,I166695,I166839);
nor I_9668 (I166395,I166441,I166822);
DFFARX1 I_9669 (I166822,I2507,I166415,I166404,);
not I_9670 (I166942,I2514);
DFFARX1 I_9671 (I94929,I2507,I166942,I166968,);
nand I_9672 (I166976,I94929,I94935);
and I_9673 (I166993,I166976,I94953);
DFFARX1 I_9674 (I166993,I2507,I166942,I167019,);
nor I_9675 (I166910,I167019,I166968);
not I_9676 (I167041,I167019);
DFFARX1 I_9677 (I94941,I2507,I166942,I167067,);
nand I_9678 (I167075,I167067,I94938);
not I_9679 (I167092,I167075);
DFFARX1 I_9680 (I167092,I2507,I166942,I167118,);
not I_9681 (I166934,I167118);
nor I_9682 (I167140,I166968,I167075);
nor I_9683 (I166916,I167019,I167140);
DFFARX1 I_9684 (I94947,I2507,I166942,I167180,);
DFFARX1 I_9685 (I167180,I2507,I166942,I167197,);
not I_9686 (I167205,I167197);
not I_9687 (I167222,I167180);
nand I_9688 (I166919,I167222,I167041);
nand I_9689 (I167253,I94932,I94932);
and I_9690 (I167270,I167253,I94944);
DFFARX1 I_9691 (I167270,I2507,I166942,I167296,);
nor I_9692 (I167304,I167296,I166968);
DFFARX1 I_9693 (I167304,I2507,I166942,I166907,);
DFFARX1 I_9694 (I167296,I2507,I166942,I166925,);
nor I_9695 (I167349,I94950,I94932);
not I_9696 (I167366,I167349);
nor I_9697 (I166928,I167205,I167366);
nand I_9698 (I166913,I167222,I167366);
nor I_9699 (I166922,I166968,I167349);
DFFARX1 I_9700 (I167349,I2507,I166942,I166931,);
not I_9701 (I167469,I2514);
DFFARX1 I_9702 (I115159,I2507,I167469,I167495,);
nand I_9703 (I167503,I115159,I115165);
and I_9704 (I167520,I167503,I115183);
DFFARX1 I_9705 (I167520,I2507,I167469,I167546,);
nor I_9706 (I167437,I167546,I167495);
not I_9707 (I167568,I167546);
DFFARX1 I_9708 (I115171,I2507,I167469,I167594,);
nand I_9709 (I167602,I167594,I115168);
not I_9710 (I167619,I167602);
DFFARX1 I_9711 (I167619,I2507,I167469,I167645,);
not I_9712 (I167461,I167645);
nor I_9713 (I167667,I167495,I167602);
nor I_9714 (I167443,I167546,I167667);
DFFARX1 I_9715 (I115177,I2507,I167469,I167707,);
DFFARX1 I_9716 (I167707,I2507,I167469,I167724,);
not I_9717 (I167732,I167724);
not I_9718 (I167749,I167707);
nand I_9719 (I167446,I167749,I167568);
nand I_9720 (I167780,I115162,I115162);
and I_9721 (I167797,I167780,I115174);
DFFARX1 I_9722 (I167797,I2507,I167469,I167823,);
nor I_9723 (I167831,I167823,I167495);
DFFARX1 I_9724 (I167831,I2507,I167469,I167434,);
DFFARX1 I_9725 (I167823,I2507,I167469,I167452,);
nor I_9726 (I167876,I115180,I115162);
not I_9727 (I167893,I167876);
nor I_9728 (I167455,I167732,I167893);
nand I_9729 (I167440,I167749,I167893);
nor I_9730 (I167449,I167495,I167876);
DFFARX1 I_9731 (I167876,I2507,I167469,I167458,);
not I_9732 (I167996,I2514);
DFFARX1 I_9733 (I62547,I2507,I167996,I168022,);
nand I_9734 (I168030,I62559,I62568);
and I_9735 (I168047,I168030,I62547);
DFFARX1 I_9736 (I168047,I2507,I167996,I168073,);
nor I_9737 (I167964,I168073,I168022);
not I_9738 (I168095,I168073);
DFFARX1 I_9739 (I62562,I2507,I167996,I168121,);
nand I_9740 (I168129,I168121,I62550);
not I_9741 (I168146,I168129);
DFFARX1 I_9742 (I168146,I2507,I167996,I168172,);
not I_9743 (I167988,I168172);
nor I_9744 (I168194,I168022,I168129);
nor I_9745 (I167970,I168073,I168194);
DFFARX1 I_9746 (I62553,I2507,I167996,I168234,);
DFFARX1 I_9747 (I168234,I2507,I167996,I168251,);
not I_9748 (I168259,I168251);
not I_9749 (I168276,I168234);
nand I_9750 (I167973,I168276,I168095);
nand I_9751 (I168307,I62544,I62544);
and I_9752 (I168324,I168307,I62556);
DFFARX1 I_9753 (I168324,I2507,I167996,I168350,);
nor I_9754 (I168358,I168350,I168022);
DFFARX1 I_9755 (I168358,I2507,I167996,I167961,);
DFFARX1 I_9756 (I168350,I2507,I167996,I167979,);
nor I_9757 (I168403,I62565,I62544);
not I_9758 (I168420,I168403);
nor I_9759 (I167982,I168259,I168420);
nand I_9760 (I167967,I168276,I168420);
nor I_9761 (I167976,I168022,I168403);
DFFARX1 I_9762 (I168403,I2507,I167996,I167985,);
not I_9763 (I168523,I2514);
DFFARX1 I_9764 (I669408,I2507,I168523,I168549,);
nand I_9765 (I168557,I669405,I669396);
and I_9766 (I168574,I168557,I669393);
DFFARX1 I_9767 (I168574,I2507,I168523,I168600,);
nor I_9768 (I168491,I168600,I168549);
not I_9769 (I168622,I168600);
DFFARX1 I_9770 (I669402,I2507,I168523,I168648,);
nand I_9771 (I168656,I168648,I669411);
not I_9772 (I168673,I168656);
DFFARX1 I_9773 (I168673,I2507,I168523,I168699,);
not I_9774 (I168515,I168699);
nor I_9775 (I168721,I168549,I168656);
nor I_9776 (I168497,I168600,I168721);
DFFARX1 I_9777 (I669414,I2507,I168523,I168761,);
DFFARX1 I_9778 (I168761,I2507,I168523,I168778,);
not I_9779 (I168786,I168778);
not I_9780 (I168803,I168761);
nand I_9781 (I168500,I168803,I168622);
nand I_9782 (I168834,I669393,I669399);
and I_9783 (I168851,I168834,I669417);
DFFARX1 I_9784 (I168851,I2507,I168523,I168877,);
nor I_9785 (I168885,I168877,I168549);
DFFARX1 I_9786 (I168885,I2507,I168523,I168488,);
DFFARX1 I_9787 (I168877,I2507,I168523,I168506,);
nor I_9788 (I168930,I669396,I669399);
not I_9789 (I168947,I168930);
nor I_9790 (I168509,I168786,I168947);
nand I_9791 (I168494,I168803,I168947);
nor I_9792 (I168503,I168549,I168930);
DFFARX1 I_9793 (I168930,I2507,I168523,I168512,);
not I_9794 (I169050,I2514);
DFFARX1 I_9795 (I421817,I2507,I169050,I169076,);
nand I_9796 (I169084,I421808,I421823);
and I_9797 (I169101,I169084,I421829);
DFFARX1 I_9798 (I169101,I2507,I169050,I169127,);
nor I_9799 (I169018,I169127,I169076);
not I_9800 (I169149,I169127);
DFFARX1 I_9801 (I421814,I2507,I169050,I169175,);
nand I_9802 (I169183,I169175,I421808);
not I_9803 (I169200,I169183);
DFFARX1 I_9804 (I169200,I2507,I169050,I169226,);
not I_9805 (I169042,I169226);
nor I_9806 (I169248,I169076,I169183);
nor I_9807 (I169024,I169127,I169248);
DFFARX1 I_9808 (I421811,I2507,I169050,I169288,);
DFFARX1 I_9809 (I169288,I2507,I169050,I169305,);
not I_9810 (I169313,I169305);
not I_9811 (I169330,I169288);
nand I_9812 (I169027,I169330,I169149);
nand I_9813 (I169361,I421805,I421820);
and I_9814 (I169378,I169361,I421805);
DFFARX1 I_9815 (I169378,I2507,I169050,I169404,);
nor I_9816 (I169412,I169404,I169076);
DFFARX1 I_9817 (I169412,I2507,I169050,I169015,);
DFFARX1 I_9818 (I169404,I2507,I169050,I169033,);
nor I_9819 (I169457,I421826,I421820);
not I_9820 (I169474,I169457);
nor I_9821 (I169036,I169313,I169474);
nand I_9822 (I169021,I169330,I169474);
nor I_9823 (I169030,I169076,I169457);
DFFARX1 I_9824 (I169457,I2507,I169050,I169039,);
not I_9825 (I169577,I2514);
DFFARX1 I_9826 (I498971,I2507,I169577,I169603,);
nand I_9827 (I169611,I498968,I498986);
and I_9828 (I169628,I169611,I498977);
DFFARX1 I_9829 (I169628,I2507,I169577,I169654,);
nor I_9830 (I169545,I169654,I169603);
not I_9831 (I169676,I169654);
DFFARX1 I_9832 (I498992,I2507,I169577,I169702,);
nand I_9833 (I169710,I169702,I498974);
not I_9834 (I169727,I169710);
DFFARX1 I_9835 (I169727,I2507,I169577,I169753,);
not I_9836 (I169569,I169753);
nor I_9837 (I169775,I169603,I169710);
nor I_9838 (I169551,I169654,I169775);
DFFARX1 I_9839 (I498980,I2507,I169577,I169815,);
DFFARX1 I_9840 (I169815,I2507,I169577,I169832,);
not I_9841 (I169840,I169832);
not I_9842 (I169857,I169815);
nand I_9843 (I169554,I169857,I169676);
nand I_9844 (I169888,I498968,I498995);
and I_9845 (I169905,I169888,I498983);
DFFARX1 I_9846 (I169905,I2507,I169577,I169931,);
nor I_9847 (I169939,I169931,I169603);
DFFARX1 I_9848 (I169939,I2507,I169577,I169542,);
DFFARX1 I_9849 (I169931,I2507,I169577,I169560,);
nor I_9850 (I169984,I498989,I498995);
not I_9851 (I170001,I169984);
nor I_9852 (I169563,I169840,I170001);
nand I_9853 (I169548,I169857,I170001);
nor I_9854 (I169557,I169603,I169984);
DFFARX1 I_9855 (I169984,I2507,I169577,I169566,);
not I_9856 (I170104,I2514);
DFFARX1 I_9857 (I373843,I2507,I170104,I170130,);
nand I_9858 (I170138,I373834,I373849);
and I_9859 (I170155,I170138,I373855);
DFFARX1 I_9860 (I170155,I2507,I170104,I170181,);
nor I_9861 (I170072,I170181,I170130);
not I_9862 (I170203,I170181);
DFFARX1 I_9863 (I373840,I2507,I170104,I170229,);
nand I_9864 (I170237,I170229,I373834);
not I_9865 (I170254,I170237);
DFFARX1 I_9866 (I170254,I2507,I170104,I170280,);
not I_9867 (I170096,I170280);
nor I_9868 (I170302,I170130,I170237);
nor I_9869 (I170078,I170181,I170302);
DFFARX1 I_9870 (I373837,I2507,I170104,I170342,);
DFFARX1 I_9871 (I170342,I2507,I170104,I170359,);
not I_9872 (I170367,I170359);
not I_9873 (I170384,I170342);
nand I_9874 (I170081,I170384,I170203);
nand I_9875 (I170415,I373831,I373846);
and I_9876 (I170432,I170415,I373831);
DFFARX1 I_9877 (I170432,I2507,I170104,I170458,);
nor I_9878 (I170466,I170458,I170130);
DFFARX1 I_9879 (I170466,I2507,I170104,I170069,);
DFFARX1 I_9880 (I170458,I2507,I170104,I170087,);
nor I_9881 (I170511,I373852,I373846);
not I_9882 (I170528,I170511);
nor I_9883 (I170090,I170367,I170528);
nand I_9884 (I170075,I170384,I170528);
nor I_9885 (I170084,I170130,I170511);
DFFARX1 I_9886 (I170511,I2507,I170104,I170093,);
not I_9887 (I170631,I2514);
DFFARX1 I_9888 (I675188,I2507,I170631,I170657,);
nand I_9889 (I170665,I675185,I675176);
and I_9890 (I170682,I170665,I675173);
DFFARX1 I_9891 (I170682,I2507,I170631,I170708,);
nor I_9892 (I170599,I170708,I170657);
not I_9893 (I170730,I170708);
DFFARX1 I_9894 (I675182,I2507,I170631,I170756,);
nand I_9895 (I170764,I170756,I675191);
not I_9896 (I170781,I170764);
DFFARX1 I_9897 (I170781,I2507,I170631,I170807,);
not I_9898 (I170623,I170807);
nor I_9899 (I170829,I170657,I170764);
nor I_9900 (I170605,I170708,I170829);
DFFARX1 I_9901 (I675194,I2507,I170631,I170869,);
DFFARX1 I_9902 (I170869,I2507,I170631,I170886,);
not I_9903 (I170894,I170886);
not I_9904 (I170911,I170869);
nand I_9905 (I170608,I170911,I170730);
nand I_9906 (I170942,I675173,I675179);
and I_9907 (I170959,I170942,I675197);
DFFARX1 I_9908 (I170959,I2507,I170631,I170985,);
nor I_9909 (I170993,I170985,I170657);
DFFARX1 I_9910 (I170993,I2507,I170631,I170596,);
DFFARX1 I_9911 (I170985,I2507,I170631,I170614,);
nor I_9912 (I171038,I675176,I675179);
not I_9913 (I171055,I171038);
nor I_9914 (I170617,I170894,I171055);
nand I_9915 (I170602,I170911,I171055);
nor I_9916 (I170611,I170657,I171038);
DFFARX1 I_9917 (I171038,I2507,I170631,I170620,);
not I_9918 (I171158,I2514);
DFFARX1 I_9919 (I525457,I2507,I171158,I171184,);
nand I_9920 (I171192,I525454,I525472);
and I_9921 (I171209,I171192,I525463);
DFFARX1 I_9922 (I171209,I2507,I171158,I171235,);
nor I_9923 (I171126,I171235,I171184);
not I_9924 (I171257,I171235);
DFFARX1 I_9925 (I525478,I2507,I171158,I171283,);
nand I_9926 (I171291,I171283,I525460);
not I_9927 (I171308,I171291);
DFFARX1 I_9928 (I171308,I2507,I171158,I171334,);
not I_9929 (I171150,I171334);
nor I_9930 (I171356,I171184,I171291);
nor I_9931 (I171132,I171235,I171356);
DFFARX1 I_9932 (I525466,I2507,I171158,I171396,);
DFFARX1 I_9933 (I171396,I2507,I171158,I171413,);
not I_9934 (I171421,I171413);
not I_9935 (I171438,I171396);
nand I_9936 (I171135,I171438,I171257);
nand I_9937 (I171469,I525454,I525481);
and I_9938 (I171486,I171469,I525469);
DFFARX1 I_9939 (I171486,I2507,I171158,I171512,);
nor I_9940 (I171520,I171512,I171184);
DFFARX1 I_9941 (I171520,I2507,I171158,I171123,);
DFFARX1 I_9942 (I171512,I2507,I171158,I171141,);
nor I_9943 (I171565,I525475,I525481);
not I_9944 (I171582,I171565);
nor I_9945 (I171144,I171421,I171582);
nand I_9946 (I171129,I171438,I171582);
nor I_9947 (I171138,I171184,I171565);
DFFARX1 I_9948 (I171565,I2507,I171158,I171147,);
not I_9949 (I171685,I2514);
DFFARX1 I_9950 (I569963,I2507,I171685,I171711,);
nand I_9951 (I171719,I569960,I569963);
and I_9952 (I171736,I171719,I569972);
DFFARX1 I_9953 (I171736,I2507,I171685,I171762,);
nor I_9954 (I171653,I171762,I171711);
not I_9955 (I171784,I171762);
DFFARX1 I_9956 (I569960,I2507,I171685,I171810,);
nand I_9957 (I171818,I171810,I569978);
not I_9958 (I171835,I171818);
DFFARX1 I_9959 (I171835,I2507,I171685,I171861,);
not I_9960 (I171677,I171861);
nor I_9961 (I171883,I171711,I171818);
nor I_9962 (I171659,I171762,I171883);
DFFARX1 I_9963 (I569966,I2507,I171685,I171923,);
DFFARX1 I_9964 (I171923,I2507,I171685,I171940,);
not I_9965 (I171948,I171940);
not I_9966 (I171965,I171923);
nand I_9967 (I171662,I171965,I171784);
nand I_9968 (I171996,I569975,I569981);
and I_9969 (I172013,I171996,I569966);
DFFARX1 I_9970 (I172013,I2507,I171685,I172039,);
nor I_9971 (I172047,I172039,I171711);
DFFARX1 I_9972 (I172047,I2507,I171685,I171650,);
DFFARX1 I_9973 (I172039,I2507,I171685,I171668,);
nor I_9974 (I172092,I569969,I569981);
not I_9975 (I172109,I172092);
nor I_9976 (I171671,I171948,I172109);
nand I_9977 (I171656,I171965,I172109);
nor I_9978 (I171665,I171711,I172092);
DFFARX1 I_9979 (I172092,I2507,I171685,I171674,);
not I_9980 (I172212,I2514);
DFFARX1 I_9981 (I486051,I2507,I172212,I172238,);
nand I_9982 (I172246,I486048,I486066);
and I_9983 (I172263,I172246,I486057);
DFFARX1 I_9984 (I172263,I2507,I172212,I172289,);
nor I_9985 (I172180,I172289,I172238);
not I_9986 (I172311,I172289);
DFFARX1 I_9987 (I486072,I2507,I172212,I172337,);
nand I_9988 (I172345,I172337,I486054);
not I_9989 (I172362,I172345);
DFFARX1 I_9990 (I172362,I2507,I172212,I172388,);
not I_9991 (I172204,I172388);
nor I_9992 (I172410,I172238,I172345);
nor I_9993 (I172186,I172289,I172410);
DFFARX1 I_9994 (I486060,I2507,I172212,I172450,);
DFFARX1 I_9995 (I172450,I2507,I172212,I172467,);
not I_9996 (I172475,I172467);
not I_9997 (I172492,I172450);
nand I_9998 (I172189,I172492,I172311);
nand I_9999 (I172523,I486048,I486075);
and I_10000 (I172540,I172523,I486063);
DFFARX1 I_10001 (I172540,I2507,I172212,I172566,);
nor I_10002 (I172574,I172566,I172238);
DFFARX1 I_10003 (I172574,I2507,I172212,I172177,);
DFFARX1 I_10004 (I172566,I2507,I172212,I172195,);
nor I_10005 (I172619,I486069,I486075);
not I_10006 (I172636,I172619);
nor I_10007 (I172198,I172475,I172636);
nand I_10008 (I172183,I172492,I172636);
nor I_10009 (I172192,I172238,I172619);
DFFARX1 I_10010 (I172619,I2507,I172212,I172201,);
not I_10011 (I172739,I2514);
DFFARX1 I_10012 (I726959,I2507,I172739,I172765,);
nand I_10013 (I172773,I726938,I726938);
and I_10014 (I172790,I172773,I726965);
DFFARX1 I_10015 (I172790,I2507,I172739,I172816,);
nor I_10016 (I172707,I172816,I172765);
not I_10017 (I172838,I172816);
DFFARX1 I_10018 (I726953,I2507,I172739,I172864,);
nand I_10019 (I172872,I172864,I726956);
not I_10020 (I172889,I172872);
DFFARX1 I_10021 (I172889,I2507,I172739,I172915,);
not I_10022 (I172731,I172915);
nor I_10023 (I172937,I172765,I172872);
nor I_10024 (I172713,I172816,I172937);
DFFARX1 I_10025 (I726947,I2507,I172739,I172977,);
DFFARX1 I_10026 (I172977,I2507,I172739,I172994,);
not I_10027 (I173002,I172994);
not I_10028 (I173019,I172977);
nand I_10029 (I172716,I173019,I172838);
nand I_10030 (I173050,I726944,I726941);
and I_10031 (I173067,I173050,I726962);
DFFARX1 I_10032 (I173067,I2507,I172739,I173093,);
nor I_10033 (I173101,I173093,I172765);
DFFARX1 I_10034 (I173101,I2507,I172739,I172704,);
DFFARX1 I_10035 (I173093,I2507,I172739,I172722,);
nor I_10036 (I173146,I726950,I726941);
not I_10037 (I173163,I173146);
nor I_10038 (I172725,I173002,I173163);
nand I_10039 (I172710,I173019,I173163);
nor I_10040 (I172719,I172765,I173146);
DFFARX1 I_10041 (I173146,I2507,I172739,I172728,);
not I_10042 (I173266,I2514);
DFFARX1 I_10043 (I132414,I2507,I173266,I173292,);
nand I_10044 (I173300,I132414,I132420);
and I_10045 (I173317,I173300,I132438);
DFFARX1 I_10046 (I173317,I2507,I173266,I173343,);
nor I_10047 (I173234,I173343,I173292);
not I_10048 (I173365,I173343);
DFFARX1 I_10049 (I132426,I2507,I173266,I173391,);
nand I_10050 (I173399,I173391,I132423);
not I_10051 (I173416,I173399);
DFFARX1 I_10052 (I173416,I2507,I173266,I173442,);
not I_10053 (I173258,I173442);
nor I_10054 (I173464,I173292,I173399);
nor I_10055 (I173240,I173343,I173464);
DFFARX1 I_10056 (I132432,I2507,I173266,I173504,);
DFFARX1 I_10057 (I173504,I2507,I173266,I173521,);
not I_10058 (I173529,I173521);
not I_10059 (I173546,I173504);
nand I_10060 (I173243,I173546,I173365);
nand I_10061 (I173577,I132417,I132417);
and I_10062 (I173594,I173577,I132429);
DFFARX1 I_10063 (I173594,I2507,I173266,I173620,);
nor I_10064 (I173628,I173620,I173292);
DFFARX1 I_10065 (I173628,I2507,I173266,I173231,);
DFFARX1 I_10066 (I173620,I2507,I173266,I173249,);
nor I_10067 (I173673,I132435,I132417);
not I_10068 (I173690,I173673);
nor I_10069 (I173252,I173529,I173690);
nand I_10070 (I173237,I173546,I173690);
nor I_10071 (I173246,I173292,I173673);
DFFARX1 I_10072 (I173673,I2507,I173266,I173255,);
not I_10073 (I173793,I2514);
DFFARX1 I_10074 (I313734,I2507,I173793,I173819,);
nand I_10075 (I173827,I313719,I313722);
and I_10076 (I173844,I173827,I313737);
DFFARX1 I_10077 (I173844,I2507,I173793,I173870,);
nor I_10078 (I173761,I173870,I173819);
not I_10079 (I173892,I173870);
DFFARX1 I_10080 (I313731,I2507,I173793,I173918,);
nand I_10081 (I173926,I173918,I313722);
not I_10082 (I173943,I173926);
DFFARX1 I_10083 (I173943,I2507,I173793,I173969,);
not I_10084 (I173785,I173969);
nor I_10085 (I173991,I173819,I173926);
nor I_10086 (I173767,I173870,I173991);
DFFARX1 I_10087 (I313728,I2507,I173793,I174031,);
DFFARX1 I_10088 (I174031,I2507,I173793,I174048,);
not I_10089 (I174056,I174048);
not I_10090 (I174073,I174031);
nand I_10091 (I173770,I174073,I173892);
nand I_10092 (I174104,I313743,I313719);
and I_10093 (I174121,I174104,I313740);
DFFARX1 I_10094 (I174121,I2507,I173793,I174147,);
nor I_10095 (I174155,I174147,I173819);
DFFARX1 I_10096 (I174155,I2507,I173793,I173758,);
DFFARX1 I_10097 (I174147,I2507,I173793,I173776,);
nor I_10098 (I174200,I313725,I313719);
not I_10099 (I174217,I174200);
nor I_10100 (I173779,I174056,I174217);
nand I_10101 (I173764,I174073,I174217);
nor I_10102 (I173773,I173819,I174200);
DFFARX1 I_10103 (I174200,I2507,I173793,I173782,);
not I_10104 (I174320,I2514);
DFFARX1 I_10105 (I384825,I2507,I174320,I174346,);
nand I_10106 (I174354,I384816,I384831);
and I_10107 (I174371,I174354,I384837);
DFFARX1 I_10108 (I174371,I2507,I174320,I174397,);
nor I_10109 (I174288,I174397,I174346);
not I_10110 (I174419,I174397);
DFFARX1 I_10111 (I384822,I2507,I174320,I174445,);
nand I_10112 (I174453,I174445,I384816);
not I_10113 (I174470,I174453);
DFFARX1 I_10114 (I174470,I2507,I174320,I174496,);
not I_10115 (I174312,I174496);
nor I_10116 (I174518,I174346,I174453);
nor I_10117 (I174294,I174397,I174518);
DFFARX1 I_10118 (I384819,I2507,I174320,I174558,);
DFFARX1 I_10119 (I174558,I2507,I174320,I174575,);
not I_10120 (I174583,I174575);
not I_10121 (I174600,I174558);
nand I_10122 (I174297,I174600,I174419);
nand I_10123 (I174631,I384813,I384828);
and I_10124 (I174648,I174631,I384813);
DFFARX1 I_10125 (I174648,I2507,I174320,I174674,);
nor I_10126 (I174682,I174674,I174346);
DFFARX1 I_10127 (I174682,I2507,I174320,I174285,);
DFFARX1 I_10128 (I174674,I2507,I174320,I174303,);
nor I_10129 (I174727,I384834,I384828);
not I_10130 (I174744,I174727);
nor I_10131 (I174306,I174583,I174744);
nand I_10132 (I174291,I174600,I174744);
nor I_10133 (I174300,I174346,I174727);
DFFARX1 I_10134 (I174727,I2507,I174320,I174309,);
not I_10135 (I174847,I2514);
DFFARX1 I_10136 (I632945,I2507,I174847,I174873,);
nand I_10137 (I174881,I632960,I632945);
and I_10138 (I174898,I174881,I632963);
DFFARX1 I_10139 (I174898,I2507,I174847,I174924,);
nor I_10140 (I174815,I174924,I174873);
not I_10141 (I174946,I174924);
DFFARX1 I_10142 (I632969,I2507,I174847,I174972,);
nand I_10143 (I174980,I174972,I632951);
not I_10144 (I174997,I174980);
DFFARX1 I_10145 (I174997,I2507,I174847,I175023,);
not I_10146 (I174839,I175023);
nor I_10147 (I175045,I174873,I174980);
nor I_10148 (I174821,I174924,I175045);
DFFARX1 I_10149 (I632948,I2507,I174847,I175085,);
DFFARX1 I_10150 (I175085,I2507,I174847,I175102,);
not I_10151 (I175110,I175102);
not I_10152 (I175127,I175085);
nand I_10153 (I174824,I175127,I174946);
nand I_10154 (I175158,I632948,I632954);
and I_10155 (I175175,I175158,I632966);
DFFARX1 I_10156 (I175175,I2507,I174847,I175201,);
nor I_10157 (I175209,I175201,I174873);
DFFARX1 I_10158 (I175209,I2507,I174847,I174812,);
DFFARX1 I_10159 (I175201,I2507,I174847,I174830,);
nor I_10160 (I175254,I632957,I632954);
not I_10161 (I175271,I175254);
nor I_10162 (I174833,I175110,I175271);
nand I_10163 (I174818,I175127,I175271);
nor I_10164 (I174827,I174873,I175254);
DFFARX1 I_10165 (I175254,I2507,I174847,I174836,);
not I_10166 (I175374,I2514);
DFFARX1 I_10167 (I398119,I2507,I175374,I175400,);
nand I_10168 (I175408,I398110,I398125);
and I_10169 (I175425,I175408,I398131);
DFFARX1 I_10170 (I175425,I2507,I175374,I175451,);
nor I_10171 (I175342,I175451,I175400);
not I_10172 (I175473,I175451);
DFFARX1 I_10173 (I398116,I2507,I175374,I175499,);
nand I_10174 (I175507,I175499,I398110);
not I_10175 (I175524,I175507);
DFFARX1 I_10176 (I175524,I2507,I175374,I175550,);
not I_10177 (I175366,I175550);
nor I_10178 (I175572,I175400,I175507);
nor I_10179 (I175348,I175451,I175572);
DFFARX1 I_10180 (I398113,I2507,I175374,I175612,);
DFFARX1 I_10181 (I175612,I2507,I175374,I175629,);
not I_10182 (I175637,I175629);
not I_10183 (I175654,I175612);
nand I_10184 (I175351,I175654,I175473);
nand I_10185 (I175685,I398107,I398122);
and I_10186 (I175702,I175685,I398107);
DFFARX1 I_10187 (I175702,I2507,I175374,I175728,);
nor I_10188 (I175736,I175728,I175400);
DFFARX1 I_10189 (I175736,I2507,I175374,I175339,);
DFFARX1 I_10190 (I175728,I2507,I175374,I175357,);
nor I_10191 (I175781,I398128,I398122);
not I_10192 (I175798,I175781);
nor I_10193 (I175360,I175637,I175798);
nand I_10194 (I175345,I175654,I175798);
nor I_10195 (I175354,I175400,I175781);
DFFARX1 I_10196 (I175781,I2507,I175374,I175363,);
not I_10197 (I175901,I2514);
DFFARX1 I_10198 (I651255,I2507,I175901,I175927,);
nand I_10199 (I175935,I651237,I651261);
and I_10200 (I175952,I175935,I651252);
DFFARX1 I_10201 (I175952,I2507,I175901,I175978,);
nor I_10202 (I175869,I175978,I175927);
not I_10203 (I176000,I175978);
DFFARX1 I_10204 (I651258,I2507,I175901,I176026,);
nand I_10205 (I176034,I176026,I651246);
not I_10206 (I176051,I176034);
DFFARX1 I_10207 (I176051,I2507,I175901,I176077,);
not I_10208 (I175893,I176077);
nor I_10209 (I176099,I175927,I176034);
nor I_10210 (I175875,I175978,I176099);
DFFARX1 I_10211 (I651237,I2507,I175901,I176139,);
DFFARX1 I_10212 (I176139,I2507,I175901,I176156,);
not I_10213 (I176164,I176156);
not I_10214 (I176181,I176139);
nand I_10215 (I175878,I176181,I176000);
nand I_10216 (I176212,I651243,I651240);
and I_10217 (I176229,I176212,I651249);
DFFARX1 I_10218 (I176229,I2507,I175901,I176255,);
nor I_10219 (I176263,I176255,I175927);
DFFARX1 I_10220 (I176263,I2507,I175901,I175866,);
DFFARX1 I_10221 (I176255,I2507,I175901,I175884,);
nor I_10222 (I176308,I651240,I651240);
not I_10223 (I176325,I176308);
nor I_10224 (I175887,I176164,I176325);
nand I_10225 (I175872,I176181,I176325);
nor I_10226 (I175881,I175927,I176308);
DFFARX1 I_10227 (I176308,I2507,I175901,I175890,);
not I_10228 (I176428,I2514);
DFFARX1 I_10229 (I377311,I2507,I176428,I176454,);
nand I_10230 (I176462,I377302,I377317);
and I_10231 (I176479,I176462,I377323);
DFFARX1 I_10232 (I176479,I2507,I176428,I176505,);
nor I_10233 (I176396,I176505,I176454);
not I_10234 (I176527,I176505);
DFFARX1 I_10235 (I377308,I2507,I176428,I176553,);
nand I_10236 (I176561,I176553,I377302);
not I_10237 (I176578,I176561);
DFFARX1 I_10238 (I176578,I2507,I176428,I176604,);
not I_10239 (I176420,I176604);
nor I_10240 (I176626,I176454,I176561);
nor I_10241 (I176402,I176505,I176626);
DFFARX1 I_10242 (I377305,I2507,I176428,I176666,);
DFFARX1 I_10243 (I176666,I2507,I176428,I176683,);
not I_10244 (I176691,I176683);
not I_10245 (I176708,I176666);
nand I_10246 (I176405,I176708,I176527);
nand I_10247 (I176739,I377299,I377314);
and I_10248 (I176756,I176739,I377299);
DFFARX1 I_10249 (I176756,I2507,I176428,I176782,);
nor I_10250 (I176790,I176782,I176454);
DFFARX1 I_10251 (I176790,I2507,I176428,I176393,);
DFFARX1 I_10252 (I176782,I2507,I176428,I176411,);
nor I_10253 (I176835,I377320,I377314);
not I_10254 (I176852,I176835);
nor I_10255 (I176414,I176691,I176852);
nand I_10256 (I176399,I176708,I176852);
nor I_10257 (I176408,I176454,I176835);
DFFARX1 I_10258 (I176835,I2507,I176428,I176417,);
not I_10259 (I176955,I2514);
DFFARX1 I_10260 (I373265,I2507,I176955,I176981,);
nand I_10261 (I176989,I373256,I373271);
and I_10262 (I177006,I176989,I373277);
DFFARX1 I_10263 (I177006,I2507,I176955,I177032,);
nor I_10264 (I176923,I177032,I176981);
not I_10265 (I177054,I177032);
DFFARX1 I_10266 (I373262,I2507,I176955,I177080,);
nand I_10267 (I177088,I177080,I373256);
not I_10268 (I177105,I177088);
DFFARX1 I_10269 (I177105,I2507,I176955,I177131,);
not I_10270 (I176947,I177131);
nor I_10271 (I177153,I176981,I177088);
nor I_10272 (I176929,I177032,I177153);
DFFARX1 I_10273 (I373259,I2507,I176955,I177193,);
DFFARX1 I_10274 (I177193,I2507,I176955,I177210,);
not I_10275 (I177218,I177210);
not I_10276 (I177235,I177193);
nand I_10277 (I176932,I177235,I177054);
nand I_10278 (I177266,I373253,I373268);
and I_10279 (I177283,I177266,I373253);
DFFARX1 I_10280 (I177283,I2507,I176955,I177309,);
nor I_10281 (I177317,I177309,I176981);
DFFARX1 I_10282 (I177317,I2507,I176955,I176920,);
DFFARX1 I_10283 (I177309,I2507,I176955,I176938,);
nor I_10284 (I177362,I373274,I373268);
not I_10285 (I177379,I177362);
nor I_10286 (I176941,I177218,I177379);
nand I_10287 (I176926,I177235,I177379);
nor I_10288 (I176935,I176981,I177362);
DFFARX1 I_10289 (I177362,I2507,I176955,I176944,);
not I_10290 (I177482,I2514);
DFFARX1 I_10291 (I630055,I2507,I177482,I177508,);
nand I_10292 (I177516,I630070,I630055);
and I_10293 (I177533,I177516,I630073);
DFFARX1 I_10294 (I177533,I2507,I177482,I177559,);
nor I_10295 (I177450,I177559,I177508);
not I_10296 (I177581,I177559);
DFFARX1 I_10297 (I630079,I2507,I177482,I177607,);
nand I_10298 (I177615,I177607,I630061);
not I_10299 (I177632,I177615);
DFFARX1 I_10300 (I177632,I2507,I177482,I177658,);
not I_10301 (I177474,I177658);
nor I_10302 (I177680,I177508,I177615);
nor I_10303 (I177456,I177559,I177680);
DFFARX1 I_10304 (I630058,I2507,I177482,I177720,);
DFFARX1 I_10305 (I177720,I2507,I177482,I177737,);
not I_10306 (I177745,I177737);
not I_10307 (I177762,I177720);
nand I_10308 (I177459,I177762,I177581);
nand I_10309 (I177793,I630058,I630064);
and I_10310 (I177810,I177793,I630076);
DFFARX1 I_10311 (I177810,I2507,I177482,I177836,);
nor I_10312 (I177844,I177836,I177508);
DFFARX1 I_10313 (I177844,I2507,I177482,I177447,);
DFFARX1 I_10314 (I177836,I2507,I177482,I177465,);
nor I_10315 (I177889,I630067,I630064);
not I_10316 (I177906,I177889);
nor I_10317 (I177468,I177745,I177906);
nand I_10318 (I177453,I177762,I177906);
nor I_10319 (I177462,I177508,I177889);
DFFARX1 I_10320 (I177889,I2507,I177482,I177471,);
not I_10321 (I178009,I2514);
DFFARX1 I_10322 (I704349,I2507,I178009,I178035,);
nand I_10323 (I178043,I704328,I704328);
and I_10324 (I178060,I178043,I704355);
DFFARX1 I_10325 (I178060,I2507,I178009,I178086,);
nor I_10326 (I177977,I178086,I178035);
not I_10327 (I178108,I178086);
DFFARX1 I_10328 (I704343,I2507,I178009,I178134,);
nand I_10329 (I178142,I178134,I704346);
not I_10330 (I178159,I178142);
DFFARX1 I_10331 (I178159,I2507,I178009,I178185,);
not I_10332 (I178001,I178185);
nor I_10333 (I178207,I178035,I178142);
nor I_10334 (I177983,I178086,I178207);
DFFARX1 I_10335 (I704337,I2507,I178009,I178247,);
DFFARX1 I_10336 (I178247,I2507,I178009,I178264,);
not I_10337 (I178272,I178264);
not I_10338 (I178289,I178247);
nand I_10339 (I177986,I178289,I178108);
nand I_10340 (I178320,I704334,I704331);
and I_10341 (I178337,I178320,I704352);
DFFARX1 I_10342 (I178337,I2507,I178009,I178363,);
nor I_10343 (I178371,I178363,I178035);
DFFARX1 I_10344 (I178371,I2507,I178009,I177974,);
DFFARX1 I_10345 (I178363,I2507,I178009,I177992,);
nor I_10346 (I178416,I704340,I704331);
not I_10347 (I178433,I178416);
nor I_10348 (I177995,I178272,I178433);
nand I_10349 (I177980,I178289,I178433);
nor I_10350 (I177989,I178035,I178416);
DFFARX1 I_10351 (I178416,I2507,I178009,I177998,);
not I_10352 (I178536,I2514);
DFFARX1 I_10353 (I485405,I2507,I178536,I178562,);
nand I_10354 (I178570,I485402,I485420);
and I_10355 (I178587,I178570,I485411);
DFFARX1 I_10356 (I178587,I2507,I178536,I178613,);
nor I_10357 (I178504,I178613,I178562);
not I_10358 (I178635,I178613);
DFFARX1 I_10359 (I485426,I2507,I178536,I178661,);
nand I_10360 (I178669,I178661,I485408);
not I_10361 (I178686,I178669);
DFFARX1 I_10362 (I178686,I2507,I178536,I178712,);
not I_10363 (I178528,I178712);
nor I_10364 (I178734,I178562,I178669);
nor I_10365 (I178510,I178613,I178734);
DFFARX1 I_10366 (I485414,I2507,I178536,I178774,);
DFFARX1 I_10367 (I178774,I2507,I178536,I178791,);
not I_10368 (I178799,I178791);
not I_10369 (I178816,I178774);
nand I_10370 (I178513,I178816,I178635);
nand I_10371 (I178847,I485402,I485429);
and I_10372 (I178864,I178847,I485417);
DFFARX1 I_10373 (I178864,I2507,I178536,I178890,);
nor I_10374 (I178898,I178890,I178562);
DFFARX1 I_10375 (I178898,I2507,I178536,I178501,);
DFFARX1 I_10376 (I178890,I2507,I178536,I178519,);
nor I_10377 (I178943,I485423,I485429);
not I_10378 (I178960,I178943);
nor I_10379 (I178522,I178799,I178960);
nand I_10380 (I178507,I178816,I178960);
nor I_10381 (I178516,I178562,I178943);
DFFARX1 I_10382 (I178943,I2507,I178536,I178525,);
not I_10383 (I179063,I2514);
DFFARX1 I_10384 (I430750,I2507,I179063,I179089,);
nand I_10385 (I179097,I430753,I430747);
and I_10386 (I179114,I179097,I430759);
DFFARX1 I_10387 (I179114,I2507,I179063,I179140,);
nor I_10388 (I179031,I179140,I179089);
not I_10389 (I179162,I179140);
DFFARX1 I_10390 (I430762,I2507,I179063,I179188,);
nand I_10391 (I179196,I179188,I430753);
not I_10392 (I179213,I179196);
DFFARX1 I_10393 (I179213,I2507,I179063,I179239,);
not I_10394 (I179055,I179239);
nor I_10395 (I179261,I179089,I179196);
nor I_10396 (I179037,I179140,I179261);
DFFARX1 I_10397 (I430765,I2507,I179063,I179301,);
DFFARX1 I_10398 (I179301,I2507,I179063,I179318,);
not I_10399 (I179326,I179318);
not I_10400 (I179343,I179301);
nand I_10401 (I179040,I179343,I179162);
nand I_10402 (I179374,I430747,I430756);
and I_10403 (I179391,I179374,I430750);
DFFARX1 I_10404 (I179391,I2507,I179063,I179417,);
nor I_10405 (I179425,I179417,I179089);
DFFARX1 I_10406 (I179425,I2507,I179063,I179028,);
DFFARX1 I_10407 (I179417,I2507,I179063,I179046,);
nor I_10408 (I179470,I430768,I430756);
not I_10409 (I179487,I179470);
nor I_10410 (I179049,I179326,I179487);
nand I_10411 (I179034,I179343,I179487);
nor I_10412 (I179043,I179089,I179470);
DFFARX1 I_10413 (I179470,I2507,I179063,I179052,);
not I_10414 (I179590,I2514);
DFFARX1 I_10415 (I400431,I2507,I179590,I179616,);
nand I_10416 (I179624,I400422,I400437);
and I_10417 (I179641,I179624,I400443);
DFFARX1 I_10418 (I179641,I2507,I179590,I179667,);
nor I_10419 (I179558,I179667,I179616);
not I_10420 (I179689,I179667);
DFFARX1 I_10421 (I400428,I2507,I179590,I179715,);
nand I_10422 (I179723,I179715,I400422);
not I_10423 (I179740,I179723);
DFFARX1 I_10424 (I179740,I2507,I179590,I179766,);
not I_10425 (I179582,I179766);
nor I_10426 (I179788,I179616,I179723);
nor I_10427 (I179564,I179667,I179788);
DFFARX1 I_10428 (I400425,I2507,I179590,I179828,);
DFFARX1 I_10429 (I179828,I2507,I179590,I179845,);
not I_10430 (I179853,I179845);
not I_10431 (I179870,I179828);
nand I_10432 (I179567,I179870,I179689);
nand I_10433 (I179901,I400419,I400434);
and I_10434 (I179918,I179901,I400419);
DFFARX1 I_10435 (I179918,I2507,I179590,I179944,);
nor I_10436 (I179952,I179944,I179616);
DFFARX1 I_10437 (I179952,I2507,I179590,I179555,);
DFFARX1 I_10438 (I179944,I2507,I179590,I179573,);
nor I_10439 (I179997,I400440,I400434);
not I_10440 (I180014,I179997);
nor I_10441 (I179576,I179853,I180014);
nand I_10442 (I179561,I179870,I180014);
nor I_10443 (I179570,I179616,I179997);
DFFARX1 I_10444 (I179997,I2507,I179590,I179579,);
not I_10445 (I180117,I2514);
DFFARX1 I_10446 (I437074,I2507,I180117,I180143,);
nand I_10447 (I180151,I437077,I437071);
and I_10448 (I180168,I180151,I437083);
DFFARX1 I_10449 (I180168,I2507,I180117,I180194,);
nor I_10450 (I180085,I180194,I180143);
not I_10451 (I180216,I180194);
DFFARX1 I_10452 (I437086,I2507,I180117,I180242,);
nand I_10453 (I180250,I180242,I437077);
not I_10454 (I180267,I180250);
DFFARX1 I_10455 (I180267,I2507,I180117,I180293,);
not I_10456 (I180109,I180293);
nor I_10457 (I180315,I180143,I180250);
nor I_10458 (I180091,I180194,I180315);
DFFARX1 I_10459 (I437089,I2507,I180117,I180355,);
DFFARX1 I_10460 (I180355,I2507,I180117,I180372,);
not I_10461 (I180380,I180372);
not I_10462 (I180397,I180355);
nand I_10463 (I180094,I180397,I180216);
nand I_10464 (I180428,I437071,I437080);
and I_10465 (I180445,I180428,I437074);
DFFARX1 I_10466 (I180445,I2507,I180117,I180471,);
nor I_10467 (I180479,I180471,I180143);
DFFARX1 I_10468 (I180479,I2507,I180117,I180082,);
DFFARX1 I_10469 (I180471,I2507,I180117,I180100,);
nor I_10470 (I180524,I437092,I437080);
not I_10471 (I180541,I180524);
nor I_10472 (I180103,I180380,I180541);
nand I_10473 (I180088,I180397,I180541);
nor I_10474 (I180097,I180143,I180524);
DFFARX1 I_10475 (I180524,I2507,I180117,I180106,);
not I_10476 (I180644,I2514);
DFFARX1 I_10477 (I534501,I2507,I180644,I180670,);
nand I_10478 (I180678,I534498,I534516);
and I_10479 (I180695,I180678,I534507);
DFFARX1 I_10480 (I180695,I2507,I180644,I180721,);
nor I_10481 (I180612,I180721,I180670);
not I_10482 (I180743,I180721);
DFFARX1 I_10483 (I534522,I2507,I180644,I180769,);
nand I_10484 (I180777,I180769,I534504);
not I_10485 (I180794,I180777);
DFFARX1 I_10486 (I180794,I2507,I180644,I180820,);
not I_10487 (I180636,I180820);
nor I_10488 (I180842,I180670,I180777);
nor I_10489 (I180618,I180721,I180842);
DFFARX1 I_10490 (I534510,I2507,I180644,I180882,);
DFFARX1 I_10491 (I180882,I2507,I180644,I180899,);
not I_10492 (I180907,I180899);
not I_10493 (I180924,I180882);
nand I_10494 (I180621,I180924,I180743);
nand I_10495 (I180955,I534498,I534525);
and I_10496 (I180972,I180955,I534513);
DFFARX1 I_10497 (I180972,I2507,I180644,I180998,);
nor I_10498 (I181006,I180998,I180670);
DFFARX1 I_10499 (I181006,I2507,I180644,I180609,);
DFFARX1 I_10500 (I180998,I2507,I180644,I180627,);
nor I_10501 (I181051,I534519,I534525);
not I_10502 (I181068,I181051);
nor I_10503 (I180630,I180907,I181068);
nand I_10504 (I180615,I180924,I181068);
nor I_10505 (I180624,I180670,I181051);
DFFARX1 I_10506 (I181051,I2507,I180644,I180633,);
not I_10507 (I181171,I2514);
DFFARX1 I_10508 (I316046,I2507,I181171,I181197,);
nand I_10509 (I181205,I316031,I316034);
and I_10510 (I181222,I181205,I316049);
DFFARX1 I_10511 (I181222,I2507,I181171,I181248,);
nor I_10512 (I181139,I181248,I181197);
not I_10513 (I181270,I181248);
DFFARX1 I_10514 (I316043,I2507,I181171,I181296,);
nand I_10515 (I181304,I181296,I316034);
not I_10516 (I181321,I181304);
DFFARX1 I_10517 (I181321,I2507,I181171,I181347,);
not I_10518 (I181163,I181347);
nor I_10519 (I181369,I181197,I181304);
nor I_10520 (I181145,I181248,I181369);
DFFARX1 I_10521 (I316040,I2507,I181171,I181409,);
DFFARX1 I_10522 (I181409,I2507,I181171,I181426,);
not I_10523 (I181434,I181426);
not I_10524 (I181451,I181409);
nand I_10525 (I181148,I181451,I181270);
nand I_10526 (I181482,I316055,I316031);
and I_10527 (I181499,I181482,I316052);
DFFARX1 I_10528 (I181499,I2507,I181171,I181525,);
nor I_10529 (I181533,I181525,I181197);
DFFARX1 I_10530 (I181533,I2507,I181171,I181136,);
DFFARX1 I_10531 (I181525,I2507,I181171,I181154,);
nor I_10532 (I181578,I316037,I316031);
not I_10533 (I181595,I181578);
nor I_10534 (I181157,I181434,I181595);
nand I_10535 (I181142,I181451,I181595);
nor I_10536 (I181151,I181197,I181578);
DFFARX1 I_10537 (I181578,I2507,I181171,I181160,);
not I_10538 (I181698,I2514);
DFFARX1 I_10539 (I391761,I2507,I181698,I181724,);
nand I_10540 (I181732,I391752,I391767);
and I_10541 (I181749,I181732,I391773);
DFFARX1 I_10542 (I181749,I2507,I181698,I181775,);
nor I_10543 (I181666,I181775,I181724);
not I_10544 (I181797,I181775);
DFFARX1 I_10545 (I391758,I2507,I181698,I181823,);
nand I_10546 (I181831,I181823,I391752);
not I_10547 (I181848,I181831);
DFFARX1 I_10548 (I181848,I2507,I181698,I181874,);
not I_10549 (I181690,I181874);
nor I_10550 (I181896,I181724,I181831);
nor I_10551 (I181672,I181775,I181896);
DFFARX1 I_10552 (I391755,I2507,I181698,I181936,);
DFFARX1 I_10553 (I181936,I2507,I181698,I181953,);
not I_10554 (I181961,I181953);
not I_10555 (I181978,I181936);
nand I_10556 (I181675,I181978,I181797);
nand I_10557 (I182009,I391749,I391764);
and I_10558 (I182026,I182009,I391749);
DFFARX1 I_10559 (I182026,I2507,I181698,I182052,);
nor I_10560 (I182060,I182052,I181724);
DFFARX1 I_10561 (I182060,I2507,I181698,I181663,);
DFFARX1 I_10562 (I182052,I2507,I181698,I181681,);
nor I_10563 (I182105,I391770,I391764);
not I_10564 (I182122,I182105);
nor I_10565 (I181684,I181961,I182122);
nand I_10566 (I181669,I181978,I182122);
nor I_10567 (I181678,I181724,I182105);
DFFARX1 I_10568 (I182105,I2507,I181698,I181687,);
not I_10569 (I182225,I2514);
DFFARX1 I_10570 (I543596,I2507,I182225,I182251,);
nand I_10571 (I182259,I543593,I543596);
and I_10572 (I182276,I182259,I543605);
DFFARX1 I_10573 (I182276,I2507,I182225,I182302,);
nor I_10574 (I182193,I182302,I182251);
not I_10575 (I182324,I182302);
DFFARX1 I_10576 (I543593,I2507,I182225,I182350,);
nand I_10577 (I182358,I182350,I543611);
not I_10578 (I182375,I182358);
DFFARX1 I_10579 (I182375,I2507,I182225,I182401,);
not I_10580 (I182217,I182401);
nor I_10581 (I182423,I182251,I182358);
nor I_10582 (I182199,I182302,I182423);
DFFARX1 I_10583 (I543599,I2507,I182225,I182463,);
DFFARX1 I_10584 (I182463,I2507,I182225,I182480,);
not I_10585 (I182488,I182480);
not I_10586 (I182505,I182463);
nand I_10587 (I182202,I182505,I182324);
nand I_10588 (I182536,I543608,I543614);
and I_10589 (I182553,I182536,I543599);
DFFARX1 I_10590 (I182553,I2507,I182225,I182579,);
nor I_10591 (I182587,I182579,I182251);
DFFARX1 I_10592 (I182587,I2507,I182225,I182190,);
DFFARX1 I_10593 (I182579,I2507,I182225,I182208,);
nor I_10594 (I182632,I543602,I543614);
not I_10595 (I182649,I182632);
nor I_10596 (I182211,I182488,I182649);
nand I_10597 (I182196,I182505,I182649);
nor I_10598 (I182205,I182251,I182632);
DFFARX1 I_10599 (I182632,I2507,I182225,I182214,);
not I_10600 (I182752,I2514);
DFFARX1 I_10601 (I628321,I2507,I182752,I182778,);
nand I_10602 (I182786,I628336,I628321);
and I_10603 (I182803,I182786,I628339);
DFFARX1 I_10604 (I182803,I2507,I182752,I182829,);
nor I_10605 (I182720,I182829,I182778);
not I_10606 (I182851,I182829);
DFFARX1 I_10607 (I628345,I2507,I182752,I182877,);
nand I_10608 (I182885,I182877,I628327);
not I_10609 (I182902,I182885);
DFFARX1 I_10610 (I182902,I2507,I182752,I182928,);
not I_10611 (I182744,I182928);
nor I_10612 (I182950,I182778,I182885);
nor I_10613 (I182726,I182829,I182950);
DFFARX1 I_10614 (I628324,I2507,I182752,I182990,);
DFFARX1 I_10615 (I182990,I2507,I182752,I183007,);
not I_10616 (I183015,I183007);
not I_10617 (I183032,I182990);
nand I_10618 (I182729,I183032,I182851);
nand I_10619 (I183063,I628324,I628330);
and I_10620 (I183080,I183063,I628342);
DFFARX1 I_10621 (I183080,I2507,I182752,I183106,);
nor I_10622 (I183114,I183106,I182778);
DFFARX1 I_10623 (I183114,I2507,I182752,I182717,);
DFFARX1 I_10624 (I183106,I2507,I182752,I182735,);
nor I_10625 (I183159,I628333,I628330);
not I_10626 (I183176,I183159);
nor I_10627 (I182738,I183015,I183176);
nand I_10628 (I182723,I183032,I183176);
nor I_10629 (I182732,I182778,I183159);
DFFARX1 I_10630 (I183159,I2507,I182752,I182741,);
not I_10631 (I183279,I2514);
DFFARX1 I_10632 (I399275,I2507,I183279,I183305,);
nand I_10633 (I183313,I399266,I399281);
and I_10634 (I183330,I183313,I399287);
DFFARX1 I_10635 (I183330,I2507,I183279,I183356,);
nor I_10636 (I183247,I183356,I183305);
not I_10637 (I183378,I183356);
DFFARX1 I_10638 (I399272,I2507,I183279,I183404,);
nand I_10639 (I183412,I183404,I399266);
not I_10640 (I183429,I183412);
DFFARX1 I_10641 (I183429,I2507,I183279,I183455,);
not I_10642 (I183271,I183455);
nor I_10643 (I183477,I183305,I183412);
nor I_10644 (I183253,I183356,I183477);
DFFARX1 I_10645 (I399269,I2507,I183279,I183517,);
DFFARX1 I_10646 (I183517,I2507,I183279,I183534,);
not I_10647 (I183542,I183534);
not I_10648 (I183559,I183517);
nand I_10649 (I183256,I183559,I183378);
nand I_10650 (I183590,I399263,I399278);
and I_10651 (I183607,I183590,I399263);
DFFARX1 I_10652 (I183607,I2507,I183279,I183633,);
nor I_10653 (I183641,I183633,I183305);
DFFARX1 I_10654 (I183641,I2507,I183279,I183244,);
DFFARX1 I_10655 (I183633,I2507,I183279,I183262,);
nor I_10656 (I183686,I399284,I399278);
not I_10657 (I183703,I183686);
nor I_10658 (I183265,I183542,I183703);
nand I_10659 (I183250,I183559,I183703);
nor I_10660 (I183259,I183305,I183686);
DFFARX1 I_10661 (I183686,I2507,I183279,I183268,);
not I_10662 (I183806,I2514);
DFFARX1 I_10663 (I616183,I2507,I183806,I183832,);
nand I_10664 (I183840,I616198,I616183);
and I_10665 (I183857,I183840,I616201);
DFFARX1 I_10666 (I183857,I2507,I183806,I183883,);
nor I_10667 (I183774,I183883,I183832);
not I_10668 (I183905,I183883);
DFFARX1 I_10669 (I616207,I2507,I183806,I183931,);
nand I_10670 (I183939,I183931,I616189);
not I_10671 (I183956,I183939);
DFFARX1 I_10672 (I183956,I2507,I183806,I183982,);
not I_10673 (I183798,I183982);
nor I_10674 (I184004,I183832,I183939);
nor I_10675 (I183780,I183883,I184004);
DFFARX1 I_10676 (I616186,I2507,I183806,I184044,);
DFFARX1 I_10677 (I184044,I2507,I183806,I184061,);
not I_10678 (I184069,I184061);
not I_10679 (I184086,I184044);
nand I_10680 (I183783,I184086,I183905);
nand I_10681 (I184117,I616186,I616192);
and I_10682 (I184134,I184117,I616204);
DFFARX1 I_10683 (I184134,I2507,I183806,I184160,);
nor I_10684 (I184168,I184160,I183832);
DFFARX1 I_10685 (I184168,I2507,I183806,I183771,);
DFFARX1 I_10686 (I184160,I2507,I183806,I183789,);
nor I_10687 (I184213,I616195,I616192);
not I_10688 (I184230,I184213);
nor I_10689 (I183792,I184069,I184230);
nand I_10690 (I183777,I184086,I184230);
nor I_10691 (I183786,I183832,I184213);
DFFARX1 I_10692 (I184213,I2507,I183806,I183795,);
not I_10693 (I184333,I2514);
DFFARX1 I_10694 (I575723,I2507,I184333,I184359,);
nand I_10695 (I184367,I575738,I575723);
and I_10696 (I184384,I184367,I575741);
DFFARX1 I_10697 (I184384,I2507,I184333,I184410,);
nor I_10698 (I184301,I184410,I184359);
not I_10699 (I184432,I184410);
DFFARX1 I_10700 (I575747,I2507,I184333,I184458,);
nand I_10701 (I184466,I184458,I575729);
not I_10702 (I184483,I184466);
DFFARX1 I_10703 (I184483,I2507,I184333,I184509,);
not I_10704 (I184325,I184509);
nor I_10705 (I184531,I184359,I184466);
nor I_10706 (I184307,I184410,I184531);
DFFARX1 I_10707 (I575726,I2507,I184333,I184571,);
DFFARX1 I_10708 (I184571,I2507,I184333,I184588,);
not I_10709 (I184596,I184588);
not I_10710 (I184613,I184571);
nand I_10711 (I184310,I184613,I184432);
nand I_10712 (I184644,I575726,I575732);
and I_10713 (I184661,I184644,I575744);
DFFARX1 I_10714 (I184661,I2507,I184333,I184687,);
nor I_10715 (I184695,I184687,I184359);
DFFARX1 I_10716 (I184695,I2507,I184333,I184298,);
DFFARX1 I_10717 (I184687,I2507,I184333,I184316,);
nor I_10718 (I184740,I575735,I575732);
not I_10719 (I184757,I184740);
nor I_10720 (I184319,I184596,I184757);
nand I_10721 (I184304,I184613,I184757);
nor I_10722 (I184313,I184359,I184740);
DFFARX1 I_10723 (I184740,I2507,I184333,I184322,);
not I_10724 (I184860,I2514);
DFFARX1 I_10725 (I617339,I2507,I184860,I184886,);
nand I_10726 (I184894,I617354,I617339);
and I_10727 (I184911,I184894,I617357);
DFFARX1 I_10728 (I184911,I2507,I184860,I184937,);
nor I_10729 (I184828,I184937,I184886);
not I_10730 (I184959,I184937);
DFFARX1 I_10731 (I617363,I2507,I184860,I184985,);
nand I_10732 (I184993,I184985,I617345);
not I_10733 (I185010,I184993);
DFFARX1 I_10734 (I185010,I2507,I184860,I185036,);
not I_10735 (I184852,I185036);
nor I_10736 (I185058,I184886,I184993);
nor I_10737 (I184834,I184937,I185058);
DFFARX1 I_10738 (I617342,I2507,I184860,I185098,);
DFFARX1 I_10739 (I185098,I2507,I184860,I185115,);
not I_10740 (I185123,I185115);
not I_10741 (I185140,I185098);
nand I_10742 (I184837,I185140,I184959);
nand I_10743 (I185171,I617342,I617348);
and I_10744 (I185188,I185171,I617360);
DFFARX1 I_10745 (I185188,I2507,I184860,I185214,);
nor I_10746 (I185222,I185214,I184886);
DFFARX1 I_10747 (I185222,I2507,I184860,I184825,);
DFFARX1 I_10748 (I185214,I2507,I184860,I184843,);
nor I_10749 (I185267,I617351,I617348);
not I_10750 (I185284,I185267);
nor I_10751 (I184846,I185123,I185284);
nand I_10752 (I184831,I185140,I185284);
nor I_10753 (I184840,I184886,I185267);
DFFARX1 I_10754 (I185267,I2507,I184860,I184849,);
not I_10755 (I185387,I2514);
DFFARX1 I_10756 (I575145,I2507,I185387,I185413,);
nand I_10757 (I185421,I575160,I575145);
and I_10758 (I185438,I185421,I575163);
DFFARX1 I_10759 (I185438,I2507,I185387,I185464,);
nor I_10760 (I185355,I185464,I185413);
not I_10761 (I185486,I185464);
DFFARX1 I_10762 (I575169,I2507,I185387,I185512,);
nand I_10763 (I185520,I185512,I575151);
not I_10764 (I185537,I185520);
DFFARX1 I_10765 (I185537,I2507,I185387,I185563,);
not I_10766 (I185379,I185563);
nor I_10767 (I185585,I185413,I185520);
nor I_10768 (I185361,I185464,I185585);
DFFARX1 I_10769 (I575148,I2507,I185387,I185625,);
DFFARX1 I_10770 (I185625,I2507,I185387,I185642,);
not I_10771 (I185650,I185642);
not I_10772 (I185667,I185625);
nand I_10773 (I185364,I185667,I185486);
nand I_10774 (I185698,I575148,I575154);
and I_10775 (I185715,I185698,I575166);
DFFARX1 I_10776 (I185715,I2507,I185387,I185741,);
nor I_10777 (I185749,I185741,I185413);
DFFARX1 I_10778 (I185749,I2507,I185387,I185352,);
DFFARX1 I_10779 (I185741,I2507,I185387,I185370,);
nor I_10780 (I185794,I575157,I575154);
not I_10781 (I185811,I185794);
nor I_10782 (I185373,I185650,I185811);
nand I_10783 (I185358,I185667,I185811);
nor I_10784 (I185367,I185413,I185794);
DFFARX1 I_10785 (I185794,I2507,I185387,I185376,);
not I_10786 (I185914,I2514);
DFFARX1 I_10787 (I329340,I2507,I185914,I185940,);
nand I_10788 (I185948,I329325,I329328);
and I_10789 (I185965,I185948,I329343);
DFFARX1 I_10790 (I185965,I2507,I185914,I185991,);
nor I_10791 (I185882,I185991,I185940);
not I_10792 (I186013,I185991);
DFFARX1 I_10793 (I329337,I2507,I185914,I186039,);
nand I_10794 (I186047,I186039,I329328);
not I_10795 (I186064,I186047);
DFFARX1 I_10796 (I186064,I2507,I185914,I186090,);
not I_10797 (I185906,I186090);
nor I_10798 (I186112,I185940,I186047);
nor I_10799 (I185888,I185991,I186112);
DFFARX1 I_10800 (I329334,I2507,I185914,I186152,);
DFFARX1 I_10801 (I186152,I2507,I185914,I186169,);
not I_10802 (I186177,I186169);
not I_10803 (I186194,I186152);
nand I_10804 (I185891,I186194,I186013);
nand I_10805 (I186225,I329349,I329325);
and I_10806 (I186242,I186225,I329346);
DFFARX1 I_10807 (I186242,I2507,I185914,I186268,);
nor I_10808 (I186276,I186268,I185940);
DFFARX1 I_10809 (I186276,I2507,I185914,I185879,);
DFFARX1 I_10810 (I186268,I2507,I185914,I185897,);
nor I_10811 (I186321,I329331,I329325);
not I_10812 (I186338,I186321);
nor I_10813 (I185900,I186177,I186338);
nand I_10814 (I185885,I186194,I186338);
nor I_10815 (I185894,I185940,I186321);
DFFARX1 I_10816 (I186321,I2507,I185914,I185903,);
not I_10817 (I186441,I2514);
DFFARX1 I_10818 (I320670,I2507,I186441,I186467,);
nand I_10819 (I186475,I320655,I320658);
and I_10820 (I186492,I186475,I320673);
DFFARX1 I_10821 (I186492,I2507,I186441,I186518,);
nor I_10822 (I186409,I186518,I186467);
not I_10823 (I186540,I186518);
DFFARX1 I_10824 (I320667,I2507,I186441,I186566,);
nand I_10825 (I186574,I186566,I320658);
not I_10826 (I186591,I186574);
DFFARX1 I_10827 (I186591,I2507,I186441,I186617,);
not I_10828 (I186433,I186617);
nor I_10829 (I186639,I186467,I186574);
nor I_10830 (I186415,I186518,I186639);
DFFARX1 I_10831 (I320664,I2507,I186441,I186679,);
DFFARX1 I_10832 (I186679,I2507,I186441,I186696,);
not I_10833 (I186704,I186696);
not I_10834 (I186721,I186679);
nand I_10835 (I186418,I186721,I186540);
nand I_10836 (I186752,I320679,I320655);
and I_10837 (I186769,I186752,I320676);
DFFARX1 I_10838 (I186769,I2507,I186441,I186795,);
nor I_10839 (I186803,I186795,I186467);
DFFARX1 I_10840 (I186803,I2507,I186441,I186406,);
DFFARX1 I_10841 (I186795,I2507,I186441,I186424,);
nor I_10842 (I186848,I320661,I320655);
not I_10843 (I186865,I186848);
nor I_10844 (I186427,I186704,I186865);
nand I_10845 (I186412,I186721,I186865);
nor I_10846 (I186421,I186467,I186848);
DFFARX1 I_10847 (I186848,I2507,I186441,I186430,);
not I_10848 (I186968,I2514);
DFFARX1 I_10849 (I149669,I2507,I186968,I186994,);
nand I_10850 (I187002,I149669,I149675);
and I_10851 (I187019,I187002,I149693);
DFFARX1 I_10852 (I187019,I2507,I186968,I187045,);
nor I_10853 (I186936,I187045,I186994);
not I_10854 (I187067,I187045);
DFFARX1 I_10855 (I149681,I2507,I186968,I187093,);
nand I_10856 (I187101,I187093,I149678);
not I_10857 (I187118,I187101);
DFFARX1 I_10858 (I187118,I2507,I186968,I187144,);
not I_10859 (I186960,I187144);
nor I_10860 (I187166,I186994,I187101);
nor I_10861 (I186942,I187045,I187166);
DFFARX1 I_10862 (I149687,I2507,I186968,I187206,);
DFFARX1 I_10863 (I187206,I2507,I186968,I187223,);
not I_10864 (I187231,I187223);
not I_10865 (I187248,I187206);
nand I_10866 (I186945,I187248,I187067);
nand I_10867 (I187279,I149672,I149672);
and I_10868 (I187296,I187279,I149684);
DFFARX1 I_10869 (I187296,I2507,I186968,I187322,);
nor I_10870 (I187330,I187322,I186994);
DFFARX1 I_10871 (I187330,I2507,I186968,I186933,);
DFFARX1 I_10872 (I187322,I2507,I186968,I186951,);
nor I_10873 (I187375,I149690,I149672);
not I_10874 (I187392,I187375);
nor I_10875 (I186954,I187231,I187392);
nand I_10876 (I186939,I187248,I187392);
nor I_10877 (I186948,I186994,I187375);
DFFARX1 I_10878 (I187375,I2507,I186968,I186957,);
not I_10879 (I187495,I2514);
DFFARX1 I_10880 (I468167,I2507,I187495,I187521,);
nand I_10881 (I187529,I468170,I468164);
and I_10882 (I187546,I187529,I468176);
DFFARX1 I_10883 (I187546,I2507,I187495,I187572,);
nor I_10884 (I187463,I187572,I187521);
not I_10885 (I187594,I187572);
DFFARX1 I_10886 (I468179,I2507,I187495,I187620,);
nand I_10887 (I187628,I187620,I468170);
not I_10888 (I187645,I187628);
DFFARX1 I_10889 (I187645,I2507,I187495,I187671,);
not I_10890 (I187487,I187671);
nor I_10891 (I187693,I187521,I187628);
nor I_10892 (I187469,I187572,I187693);
DFFARX1 I_10893 (I468182,I2507,I187495,I187733,);
DFFARX1 I_10894 (I187733,I2507,I187495,I187750,);
not I_10895 (I187758,I187750);
not I_10896 (I187775,I187733);
nand I_10897 (I187472,I187775,I187594);
nand I_10898 (I187806,I468164,I468173);
and I_10899 (I187823,I187806,I468167);
DFFARX1 I_10900 (I187823,I2507,I187495,I187849,);
nor I_10901 (I187857,I187849,I187521);
DFFARX1 I_10902 (I187857,I2507,I187495,I187460,);
DFFARX1 I_10903 (I187849,I2507,I187495,I187478,);
nor I_10904 (I187902,I468185,I468173);
not I_10905 (I187919,I187902);
nor I_10906 (I187481,I187758,I187919);
nand I_10907 (I187466,I187775,I187919);
nor I_10908 (I187475,I187521,I187902);
DFFARX1 I_10909 (I187902,I2507,I187495,I187484,);
not I_10910 (I188022,I2514);
DFFARX1 I_10911 (I290296,I2507,I188022,I188048,);
nand I_10912 (I188056,I290296,I290308);
and I_10913 (I188073,I188056,I290293);
DFFARX1 I_10914 (I188073,I2507,I188022,I188099,);
nor I_10915 (I187990,I188099,I188048);
not I_10916 (I188121,I188099);
DFFARX1 I_10917 (I290317,I2507,I188022,I188147,);
nand I_10918 (I188155,I188147,I290314);
not I_10919 (I188172,I188155);
DFFARX1 I_10920 (I188172,I2507,I188022,I188198,);
not I_10921 (I188014,I188198);
nor I_10922 (I188220,I188048,I188155);
nor I_10923 (I187996,I188099,I188220);
DFFARX1 I_10924 (I290305,I2507,I188022,I188260,);
DFFARX1 I_10925 (I188260,I2507,I188022,I188277,);
not I_10926 (I188285,I188277);
not I_10927 (I188302,I188260);
nand I_10928 (I187999,I188302,I188121);
nand I_10929 (I188333,I290293,I290302);
and I_10930 (I188350,I188333,I290311);
DFFARX1 I_10931 (I188350,I2507,I188022,I188376,);
nor I_10932 (I188384,I188376,I188048);
DFFARX1 I_10933 (I188384,I2507,I188022,I187987,);
DFFARX1 I_10934 (I188376,I2507,I188022,I188005,);
nor I_10935 (I188429,I290299,I290302);
not I_10936 (I188446,I188429);
nor I_10937 (I188008,I188285,I188446);
nand I_10938 (I187993,I188302,I188446);
nor I_10939 (I188002,I188048,I188429);
DFFARX1 I_10940 (I188429,I2507,I188022,I188011,);
not I_10941 (I188549,I2514);
DFFARX1 I_10942 (I714464,I2507,I188549,I188575,);
nand I_10943 (I188583,I714443,I714443);
and I_10944 (I188600,I188583,I714470);
DFFARX1 I_10945 (I188600,I2507,I188549,I188626,);
nor I_10946 (I188517,I188626,I188575);
not I_10947 (I188648,I188626);
DFFARX1 I_10948 (I714458,I2507,I188549,I188674,);
nand I_10949 (I188682,I188674,I714461);
not I_10950 (I188699,I188682);
DFFARX1 I_10951 (I188699,I2507,I188549,I188725,);
not I_10952 (I188541,I188725);
nor I_10953 (I188747,I188575,I188682);
nor I_10954 (I188523,I188626,I188747);
DFFARX1 I_10955 (I714452,I2507,I188549,I188787,);
DFFARX1 I_10956 (I188787,I2507,I188549,I188804,);
not I_10957 (I188812,I188804);
not I_10958 (I188829,I188787);
nand I_10959 (I188526,I188829,I188648);
nand I_10960 (I188860,I714449,I714446);
and I_10961 (I188877,I188860,I714467);
DFFARX1 I_10962 (I188877,I2507,I188549,I188903,);
nor I_10963 (I188911,I188903,I188575);
DFFARX1 I_10964 (I188911,I2507,I188549,I188514,);
DFFARX1 I_10965 (I188903,I2507,I188549,I188532,);
nor I_10966 (I188956,I714455,I714446);
not I_10967 (I188973,I188956);
nor I_10968 (I188535,I188812,I188973);
nand I_10969 (I188520,I188829,I188973);
nor I_10970 (I188529,I188575,I188956);
DFFARX1 I_10971 (I188956,I2507,I188549,I188538,);
not I_10972 (I189076,I2514);
DFFARX1 I_10973 (I152049,I2507,I189076,I189102,);
nand I_10974 (I189110,I152049,I152055);
and I_10975 (I189127,I189110,I152073);
DFFARX1 I_10976 (I189127,I2507,I189076,I189153,);
nor I_10977 (I189044,I189153,I189102);
not I_10978 (I189175,I189153);
DFFARX1 I_10979 (I152061,I2507,I189076,I189201,);
nand I_10980 (I189209,I189201,I152058);
not I_10981 (I189226,I189209);
DFFARX1 I_10982 (I189226,I2507,I189076,I189252,);
not I_10983 (I189068,I189252);
nor I_10984 (I189274,I189102,I189209);
nor I_10985 (I189050,I189153,I189274);
DFFARX1 I_10986 (I152067,I2507,I189076,I189314,);
DFFARX1 I_10987 (I189314,I2507,I189076,I189331,);
not I_10988 (I189339,I189331);
not I_10989 (I189356,I189314);
nand I_10990 (I189053,I189356,I189175);
nand I_10991 (I189387,I152052,I152052);
and I_10992 (I189404,I189387,I152064);
DFFARX1 I_10993 (I189404,I2507,I189076,I189430,);
nor I_10994 (I189438,I189430,I189102);
DFFARX1 I_10995 (I189438,I2507,I189076,I189041,);
DFFARX1 I_10996 (I189430,I2507,I189076,I189059,);
nor I_10997 (I189483,I152070,I152052);
not I_10998 (I189500,I189483);
nor I_10999 (I189062,I189339,I189500);
nand I_11000 (I189047,I189356,I189500);
nor I_11001 (I189056,I189102,I189483);
DFFARX1 I_11002 (I189483,I2507,I189076,I189065,);
not I_11003 (I189603,I2514);
DFFARX1 I_11004 (I642007,I2507,I189603,I189629,);
nand I_11005 (I189637,I641989,I642013);
and I_11006 (I189654,I189637,I642004);
DFFARX1 I_11007 (I189654,I2507,I189603,I189680,);
nor I_11008 (I189571,I189680,I189629);
not I_11009 (I189702,I189680);
DFFARX1 I_11010 (I642010,I2507,I189603,I189728,);
nand I_11011 (I189736,I189728,I641998);
not I_11012 (I189753,I189736);
DFFARX1 I_11013 (I189753,I2507,I189603,I189779,);
not I_11014 (I189595,I189779);
nor I_11015 (I189801,I189629,I189736);
nor I_11016 (I189577,I189680,I189801);
DFFARX1 I_11017 (I641989,I2507,I189603,I189841,);
DFFARX1 I_11018 (I189841,I2507,I189603,I189858,);
not I_11019 (I189866,I189858);
not I_11020 (I189883,I189841);
nand I_11021 (I189580,I189883,I189702);
nand I_11022 (I189914,I641995,I641992);
and I_11023 (I189931,I189914,I642001);
DFFARX1 I_11024 (I189931,I2507,I189603,I189957,);
nor I_11025 (I189965,I189957,I189629);
DFFARX1 I_11026 (I189965,I2507,I189603,I189568,);
DFFARX1 I_11027 (I189957,I2507,I189603,I189586,);
nor I_11028 (I190010,I641992,I641992);
not I_11029 (I190027,I190010);
nor I_11030 (I189589,I189866,I190027);
nand I_11031 (I189574,I189883,I190027);
nor I_11032 (I189583,I189629,I190010);
DFFARX1 I_11033 (I190010,I2507,I189603,I189592,);
not I_11034 (I190130,I2514);
DFFARX1 I_11035 (I478945,I2507,I190130,I190156,);
nand I_11036 (I190164,I478942,I478960);
and I_11037 (I190181,I190164,I478951);
DFFARX1 I_11038 (I190181,I2507,I190130,I190207,);
nor I_11039 (I190098,I190207,I190156);
not I_11040 (I190229,I190207);
DFFARX1 I_11041 (I478966,I2507,I190130,I190255,);
nand I_11042 (I190263,I190255,I478948);
not I_11043 (I190280,I190263);
DFFARX1 I_11044 (I190280,I2507,I190130,I190306,);
not I_11045 (I190122,I190306);
nor I_11046 (I190328,I190156,I190263);
nor I_11047 (I190104,I190207,I190328);
DFFARX1 I_11048 (I478954,I2507,I190130,I190368,);
DFFARX1 I_11049 (I190368,I2507,I190130,I190385,);
not I_11050 (I190393,I190385);
not I_11051 (I190410,I190368);
nand I_11052 (I190107,I190410,I190229);
nand I_11053 (I190441,I478942,I478969);
and I_11054 (I190458,I190441,I478957);
DFFARX1 I_11055 (I190458,I2507,I190130,I190484,);
nor I_11056 (I190492,I190484,I190156);
DFFARX1 I_11057 (I190492,I2507,I190130,I190095,);
DFFARX1 I_11058 (I190484,I2507,I190130,I190113,);
nor I_11059 (I190537,I478963,I478969);
not I_11060 (I190554,I190537);
nor I_11061 (I190116,I190393,I190554);
nand I_11062 (I190101,I190410,I190554);
nor I_11063 (I190110,I190156,I190537);
DFFARX1 I_11064 (I190537,I2507,I190130,I190119,);
not I_11065 (I190657,I2514);
DFFARX1 I_11066 (I619073,I2507,I190657,I190683,);
nand I_11067 (I190691,I619088,I619073);
and I_11068 (I190708,I190691,I619091);
DFFARX1 I_11069 (I190708,I2507,I190657,I190734,);
nor I_11070 (I190625,I190734,I190683);
not I_11071 (I190756,I190734);
DFFARX1 I_11072 (I619097,I2507,I190657,I190782,);
nand I_11073 (I190790,I190782,I619079);
not I_11074 (I190807,I190790);
DFFARX1 I_11075 (I190807,I2507,I190657,I190833,);
not I_11076 (I190649,I190833);
nor I_11077 (I190855,I190683,I190790);
nor I_11078 (I190631,I190734,I190855);
DFFARX1 I_11079 (I619076,I2507,I190657,I190895,);
DFFARX1 I_11080 (I190895,I2507,I190657,I190912,);
not I_11081 (I190920,I190912);
not I_11082 (I190937,I190895);
nand I_11083 (I190634,I190937,I190756);
nand I_11084 (I190968,I619076,I619082);
and I_11085 (I190985,I190968,I619094);
DFFARX1 I_11086 (I190985,I2507,I190657,I191011,);
nor I_11087 (I191019,I191011,I190683);
DFFARX1 I_11088 (I191019,I2507,I190657,I190622,);
DFFARX1 I_11089 (I191011,I2507,I190657,I190640,);
nor I_11090 (I191064,I619085,I619082);
not I_11091 (I191081,I191064);
nor I_11092 (I190643,I190920,I191081);
nand I_11093 (I190628,I190937,I191081);
nor I_11094 (I190637,I190683,I191064);
DFFARX1 I_11095 (I191064,I2507,I190657,I190646,);
not I_11096 (I191184,I2514);
DFFARX1 I_11097 (I639831,I2507,I191184,I191210,);
nand I_11098 (I191218,I639813,I639837);
and I_11099 (I191235,I191218,I639828);
DFFARX1 I_11100 (I191235,I2507,I191184,I191261,);
nor I_11101 (I191152,I191261,I191210);
not I_11102 (I191283,I191261);
DFFARX1 I_11103 (I639834,I2507,I191184,I191309,);
nand I_11104 (I191317,I191309,I639822);
not I_11105 (I191334,I191317);
DFFARX1 I_11106 (I191334,I2507,I191184,I191360,);
not I_11107 (I191176,I191360);
nor I_11108 (I191382,I191210,I191317);
nor I_11109 (I191158,I191261,I191382);
DFFARX1 I_11110 (I639813,I2507,I191184,I191422,);
DFFARX1 I_11111 (I191422,I2507,I191184,I191439,);
not I_11112 (I191447,I191439);
not I_11113 (I191464,I191422);
nand I_11114 (I191161,I191464,I191283);
nand I_11115 (I191495,I639819,I639816);
and I_11116 (I191512,I191495,I639825);
DFFARX1 I_11117 (I191512,I2507,I191184,I191538,);
nor I_11118 (I191546,I191538,I191210);
DFFARX1 I_11119 (I191546,I2507,I191184,I191149,);
DFFARX1 I_11120 (I191538,I2507,I191184,I191167,);
nor I_11121 (I191591,I639816,I639816);
not I_11122 (I191608,I191591);
nor I_11123 (I191170,I191447,I191608);
nand I_11124 (I191155,I191464,I191608);
nor I_11125 (I191164,I191210,I191591);
DFFARX1 I_11126 (I191591,I2507,I191184,I191173,);
not I_11127 (I191711,I2514);
DFFARX1 I_11128 (I302174,I2507,I191711,I191737,);
nand I_11129 (I191745,I302159,I302162);
and I_11130 (I191762,I191745,I302177);
DFFARX1 I_11131 (I191762,I2507,I191711,I191788,);
nor I_11132 (I191679,I191788,I191737);
not I_11133 (I191810,I191788);
DFFARX1 I_11134 (I302171,I2507,I191711,I191836,);
nand I_11135 (I191844,I191836,I302162);
not I_11136 (I191861,I191844);
DFFARX1 I_11137 (I191861,I2507,I191711,I191887,);
not I_11138 (I191703,I191887);
nor I_11139 (I191909,I191737,I191844);
nor I_11140 (I191685,I191788,I191909);
DFFARX1 I_11141 (I302168,I2507,I191711,I191949,);
DFFARX1 I_11142 (I191949,I2507,I191711,I191966,);
not I_11143 (I191974,I191966);
not I_11144 (I191991,I191949);
nand I_11145 (I191688,I191991,I191810);
nand I_11146 (I192022,I302183,I302159);
and I_11147 (I192039,I192022,I302180);
DFFARX1 I_11148 (I192039,I2507,I191711,I192065,);
nor I_11149 (I192073,I192065,I191737);
DFFARX1 I_11150 (I192073,I2507,I191711,I191676,);
DFFARX1 I_11151 (I192065,I2507,I191711,I191694,);
nor I_11152 (I192118,I302165,I302159);
not I_11153 (I192135,I192118);
nor I_11154 (I191697,I191974,I192135);
nand I_11155 (I191682,I191991,I192135);
nor I_11156 (I191691,I191737,I192118);
DFFARX1 I_11157 (I192118,I2507,I191711,I191700,);
not I_11158 (I192238,I2514);
DFFARX1 I_11159 (I655607,I2507,I192238,I192264,);
nand I_11160 (I192272,I655589,I655613);
and I_11161 (I192289,I192272,I655604);
DFFARX1 I_11162 (I192289,I2507,I192238,I192315,);
nor I_11163 (I192206,I192315,I192264);
not I_11164 (I192337,I192315);
DFFARX1 I_11165 (I655610,I2507,I192238,I192363,);
nand I_11166 (I192371,I192363,I655598);
not I_11167 (I192388,I192371);
DFFARX1 I_11168 (I192388,I2507,I192238,I192414,);
not I_11169 (I192230,I192414);
nor I_11170 (I192436,I192264,I192371);
nor I_11171 (I192212,I192315,I192436);
DFFARX1 I_11172 (I655589,I2507,I192238,I192476,);
DFFARX1 I_11173 (I192476,I2507,I192238,I192493,);
not I_11174 (I192501,I192493);
not I_11175 (I192518,I192476);
nand I_11176 (I192215,I192518,I192337);
nand I_11177 (I192549,I655595,I655592);
and I_11178 (I192566,I192549,I655601);
DFFARX1 I_11179 (I192566,I2507,I192238,I192592,);
nor I_11180 (I192600,I192592,I192264);
DFFARX1 I_11181 (I192600,I2507,I192238,I192203,);
DFFARX1 I_11182 (I192592,I2507,I192238,I192221,);
nor I_11183 (I192645,I655592,I655592);
not I_11184 (I192662,I192645);
nor I_11185 (I192224,I192501,I192662);
nand I_11186 (I192209,I192518,I192662);
nor I_11187 (I192218,I192264,I192645);
DFFARX1 I_11188 (I192645,I2507,I192238,I192227,);
not I_11189 (I192765,I2514);
DFFARX1 I_11190 (I535147,I2507,I192765,I192791,);
nand I_11191 (I192799,I535144,I535162);
and I_11192 (I192816,I192799,I535153);
DFFARX1 I_11193 (I192816,I2507,I192765,I192842,);
nor I_11194 (I192733,I192842,I192791);
not I_11195 (I192864,I192842);
DFFARX1 I_11196 (I535168,I2507,I192765,I192890,);
nand I_11197 (I192898,I192890,I535150);
not I_11198 (I192915,I192898);
DFFARX1 I_11199 (I192915,I2507,I192765,I192941,);
not I_11200 (I192757,I192941);
nor I_11201 (I192963,I192791,I192898);
nor I_11202 (I192739,I192842,I192963);
DFFARX1 I_11203 (I535156,I2507,I192765,I193003,);
DFFARX1 I_11204 (I193003,I2507,I192765,I193020,);
not I_11205 (I193028,I193020);
not I_11206 (I193045,I193003);
nand I_11207 (I192742,I193045,I192864);
nand I_11208 (I193076,I535144,I535171);
and I_11209 (I193093,I193076,I535159);
DFFARX1 I_11210 (I193093,I2507,I192765,I193119,);
nor I_11211 (I193127,I193119,I192791);
DFFARX1 I_11212 (I193127,I2507,I192765,I192730,);
DFFARX1 I_11213 (I193119,I2507,I192765,I192748,);
nor I_11214 (I193172,I535165,I535171);
not I_11215 (I193189,I193172);
nor I_11216 (I192751,I193028,I193189);
nand I_11217 (I192736,I193045,I193189);
nor I_11218 (I192745,I192791,I193172);
DFFARX1 I_11219 (I193172,I2507,I192765,I192754,);
not I_11220 (I193292,I2514);
DFFARX1 I_11221 (I729934,I2507,I193292,I193318,);
nand I_11222 (I193326,I729913,I729913);
and I_11223 (I193343,I193326,I729940);
DFFARX1 I_11224 (I193343,I2507,I193292,I193369,);
nor I_11225 (I193260,I193369,I193318);
not I_11226 (I193391,I193369);
DFFARX1 I_11227 (I729928,I2507,I193292,I193417,);
nand I_11228 (I193425,I193417,I729931);
not I_11229 (I193442,I193425);
DFFARX1 I_11230 (I193442,I2507,I193292,I193468,);
not I_11231 (I193284,I193468);
nor I_11232 (I193490,I193318,I193425);
nor I_11233 (I193266,I193369,I193490);
DFFARX1 I_11234 (I729922,I2507,I193292,I193530,);
DFFARX1 I_11235 (I193530,I2507,I193292,I193547,);
not I_11236 (I193555,I193547);
not I_11237 (I193572,I193530);
nand I_11238 (I193269,I193572,I193391);
nand I_11239 (I193603,I729919,I729916);
and I_11240 (I193620,I193603,I729937);
DFFARX1 I_11241 (I193620,I2507,I193292,I193646,);
nor I_11242 (I193654,I193646,I193318);
DFFARX1 I_11243 (I193654,I2507,I193292,I193257,);
DFFARX1 I_11244 (I193646,I2507,I193292,I193275,);
nor I_11245 (I193699,I729925,I729916);
not I_11246 (I193716,I193699);
nor I_11247 (I193278,I193555,I193716);
nand I_11248 (I193263,I193572,I193716);
nor I_11249 (I193272,I193318,I193699);
DFFARX1 I_11250 (I193699,I2507,I193292,I193281,);
not I_11251 (I193819,I2514);
DFFARX1 I_11252 (I147884,I2507,I193819,I193845,);
nand I_11253 (I193853,I147884,I147890);
and I_11254 (I193870,I193853,I147908);
DFFARX1 I_11255 (I193870,I2507,I193819,I193896,);
nor I_11256 (I193787,I193896,I193845);
not I_11257 (I193918,I193896);
DFFARX1 I_11258 (I147896,I2507,I193819,I193944,);
nand I_11259 (I193952,I193944,I147893);
not I_11260 (I193969,I193952);
DFFARX1 I_11261 (I193969,I2507,I193819,I193995,);
not I_11262 (I193811,I193995);
nor I_11263 (I194017,I193845,I193952);
nor I_11264 (I193793,I193896,I194017);
DFFARX1 I_11265 (I147902,I2507,I193819,I194057,);
DFFARX1 I_11266 (I194057,I2507,I193819,I194074,);
not I_11267 (I194082,I194074);
not I_11268 (I194099,I194057);
nand I_11269 (I193796,I194099,I193918);
nand I_11270 (I194130,I147887,I147887);
and I_11271 (I194147,I194130,I147899);
DFFARX1 I_11272 (I194147,I2507,I193819,I194173,);
nor I_11273 (I194181,I194173,I193845);
DFFARX1 I_11274 (I194181,I2507,I193819,I193784,);
DFFARX1 I_11275 (I194173,I2507,I193819,I193802,);
nor I_11276 (I194226,I147905,I147887);
not I_11277 (I194243,I194226);
nor I_11278 (I193805,I194082,I194243);
nand I_11279 (I193790,I194099,I194243);
nor I_11280 (I193799,I193845,I194226);
DFFARX1 I_11281 (I194226,I2507,I193819,I193808,);
not I_11282 (I194346,I2514);
DFFARX1 I_11283 (I301596,I2507,I194346,I194372,);
nand I_11284 (I194380,I301581,I301584);
and I_11285 (I194397,I194380,I301599);
DFFARX1 I_11286 (I194397,I2507,I194346,I194423,);
nor I_11287 (I194314,I194423,I194372);
not I_11288 (I194445,I194423);
DFFARX1 I_11289 (I301593,I2507,I194346,I194471,);
nand I_11290 (I194479,I194471,I301584);
not I_11291 (I194496,I194479);
DFFARX1 I_11292 (I194496,I2507,I194346,I194522,);
not I_11293 (I194338,I194522);
nor I_11294 (I194544,I194372,I194479);
nor I_11295 (I194320,I194423,I194544);
DFFARX1 I_11296 (I301590,I2507,I194346,I194584,);
DFFARX1 I_11297 (I194584,I2507,I194346,I194601,);
not I_11298 (I194609,I194601);
not I_11299 (I194626,I194584);
nand I_11300 (I194323,I194626,I194445);
nand I_11301 (I194657,I301605,I301581);
and I_11302 (I194674,I194657,I301602);
DFFARX1 I_11303 (I194674,I2507,I194346,I194700,);
nor I_11304 (I194708,I194700,I194372);
DFFARX1 I_11305 (I194708,I2507,I194346,I194311,);
DFFARX1 I_11306 (I194700,I2507,I194346,I194329,);
nor I_11307 (I194753,I301587,I301581);
not I_11308 (I194770,I194753);
nor I_11309 (I194332,I194609,I194770);
nand I_11310 (I194317,I194626,I194770);
nor I_11311 (I194326,I194372,I194753);
DFFARX1 I_11312 (I194753,I2507,I194346,I194335,);
not I_11313 (I194873,I2514);
DFFARX1 I_11314 (I122894,I2507,I194873,I194899,);
nand I_11315 (I194907,I122894,I122900);
and I_11316 (I194924,I194907,I122918);
DFFARX1 I_11317 (I194924,I2507,I194873,I194950,);
nor I_11318 (I194841,I194950,I194899);
not I_11319 (I194972,I194950);
DFFARX1 I_11320 (I122906,I2507,I194873,I194998,);
nand I_11321 (I195006,I194998,I122903);
not I_11322 (I195023,I195006);
DFFARX1 I_11323 (I195023,I2507,I194873,I195049,);
not I_11324 (I194865,I195049);
nor I_11325 (I195071,I194899,I195006);
nor I_11326 (I194847,I194950,I195071);
DFFARX1 I_11327 (I122912,I2507,I194873,I195111,);
DFFARX1 I_11328 (I195111,I2507,I194873,I195128,);
not I_11329 (I195136,I195128);
not I_11330 (I195153,I195111);
nand I_11331 (I194850,I195153,I194972);
nand I_11332 (I195184,I122897,I122897);
and I_11333 (I195201,I195184,I122909);
DFFARX1 I_11334 (I195201,I2507,I194873,I195227,);
nor I_11335 (I195235,I195227,I194899);
DFFARX1 I_11336 (I195235,I2507,I194873,I194838,);
DFFARX1 I_11337 (I195227,I2507,I194873,I194856,);
nor I_11338 (I195280,I122915,I122897);
not I_11339 (I195297,I195280);
nor I_11340 (I194859,I195136,I195297);
nand I_11341 (I194844,I195153,I195297);
nor I_11342 (I194853,I194899,I195280);
DFFARX1 I_11343 (I195280,I2507,I194873,I194862,);
not I_11344 (I195400,I2514);
DFFARX1 I_11345 (I309688,I2507,I195400,I195426,);
nand I_11346 (I195434,I309673,I309676);
and I_11347 (I195451,I195434,I309691);
DFFARX1 I_11348 (I195451,I2507,I195400,I195477,);
nor I_11349 (I195368,I195477,I195426);
not I_11350 (I195499,I195477);
DFFARX1 I_11351 (I309685,I2507,I195400,I195525,);
nand I_11352 (I195533,I195525,I309676);
not I_11353 (I195550,I195533);
DFFARX1 I_11354 (I195550,I2507,I195400,I195576,);
not I_11355 (I195392,I195576);
nor I_11356 (I195598,I195426,I195533);
nor I_11357 (I195374,I195477,I195598);
DFFARX1 I_11358 (I309682,I2507,I195400,I195638,);
DFFARX1 I_11359 (I195638,I2507,I195400,I195655,);
not I_11360 (I195663,I195655);
not I_11361 (I195680,I195638);
nand I_11362 (I195377,I195680,I195499);
nand I_11363 (I195711,I309697,I309673);
and I_11364 (I195728,I195711,I309694);
DFFARX1 I_11365 (I195728,I2507,I195400,I195754,);
nor I_11366 (I195762,I195754,I195426);
DFFARX1 I_11367 (I195762,I2507,I195400,I195365,);
DFFARX1 I_11368 (I195754,I2507,I195400,I195383,);
nor I_11369 (I195807,I309679,I309673);
not I_11370 (I195824,I195807);
nor I_11371 (I195386,I195663,I195824);
nand I_11372 (I195371,I195680,I195824);
nor I_11373 (I195380,I195426,I195807);
DFFARX1 I_11374 (I195807,I2507,I195400,I195389,);
not I_11375 (I195927,I2514);
DFFARX1 I_11376 (I324138,I2507,I195927,I195953,);
nand I_11377 (I195961,I324123,I324126);
and I_11378 (I195978,I195961,I324141);
DFFARX1 I_11379 (I195978,I2507,I195927,I196004,);
nor I_11380 (I195895,I196004,I195953);
not I_11381 (I196026,I196004);
DFFARX1 I_11382 (I324135,I2507,I195927,I196052,);
nand I_11383 (I196060,I196052,I324126);
not I_11384 (I196077,I196060);
DFFARX1 I_11385 (I196077,I2507,I195927,I196103,);
not I_11386 (I195919,I196103);
nor I_11387 (I196125,I195953,I196060);
nor I_11388 (I195901,I196004,I196125);
DFFARX1 I_11389 (I324132,I2507,I195927,I196165,);
DFFARX1 I_11390 (I196165,I2507,I195927,I196182,);
not I_11391 (I196190,I196182);
not I_11392 (I196207,I196165);
nand I_11393 (I195904,I196207,I196026);
nand I_11394 (I196238,I324147,I324123);
and I_11395 (I196255,I196238,I324144);
DFFARX1 I_11396 (I196255,I2507,I195927,I196281,);
nor I_11397 (I196289,I196281,I195953);
DFFARX1 I_11398 (I196289,I2507,I195927,I195892,);
DFFARX1 I_11399 (I196281,I2507,I195927,I195910,);
nor I_11400 (I196334,I324129,I324123);
not I_11401 (I196351,I196334);
nor I_11402 (I195913,I196190,I196351);
nand I_11403 (I195898,I196207,I196351);
nor I_11404 (I195907,I195953,I196334);
DFFARX1 I_11405 (I196334,I2507,I195927,I195916,);
not I_11406 (I196454,I2514);
DFFARX1 I_11407 (I343212,I2507,I196454,I196480,);
nand I_11408 (I196488,I343197,I343200);
and I_11409 (I196505,I196488,I343215);
DFFARX1 I_11410 (I196505,I2507,I196454,I196531,);
nor I_11411 (I196422,I196531,I196480);
not I_11412 (I196553,I196531);
DFFARX1 I_11413 (I343209,I2507,I196454,I196579,);
nand I_11414 (I196587,I196579,I343200);
not I_11415 (I196604,I196587);
DFFARX1 I_11416 (I196604,I2507,I196454,I196630,);
not I_11417 (I196446,I196630);
nor I_11418 (I196652,I196480,I196587);
nor I_11419 (I196428,I196531,I196652);
DFFARX1 I_11420 (I343206,I2507,I196454,I196692,);
DFFARX1 I_11421 (I196692,I2507,I196454,I196709,);
not I_11422 (I196717,I196709);
not I_11423 (I196734,I196692);
nand I_11424 (I196431,I196734,I196553);
nand I_11425 (I196765,I343221,I343197);
and I_11426 (I196782,I196765,I343218);
DFFARX1 I_11427 (I196782,I2507,I196454,I196808,);
nor I_11428 (I196816,I196808,I196480);
DFFARX1 I_11429 (I196816,I2507,I196454,I196419,);
DFFARX1 I_11430 (I196808,I2507,I196454,I196437,);
nor I_11431 (I196861,I343203,I343197);
not I_11432 (I196878,I196861);
nor I_11433 (I196440,I196717,I196878);
nand I_11434 (I196425,I196734,I196878);
nor I_11435 (I196434,I196480,I196861);
DFFARX1 I_11436 (I196861,I2507,I196454,I196443,);
not I_11437 (I196981,I2514);
DFFARX1 I_11438 (I47264,I2507,I196981,I197007,);
nand I_11439 (I197015,I47276,I47285);
and I_11440 (I197032,I197015,I47264);
DFFARX1 I_11441 (I197032,I2507,I196981,I197058,);
nor I_11442 (I196949,I197058,I197007);
not I_11443 (I197080,I197058);
DFFARX1 I_11444 (I47279,I2507,I196981,I197106,);
nand I_11445 (I197114,I197106,I47267);
not I_11446 (I197131,I197114);
DFFARX1 I_11447 (I197131,I2507,I196981,I197157,);
not I_11448 (I196973,I197157);
nor I_11449 (I197179,I197007,I197114);
nor I_11450 (I196955,I197058,I197179);
DFFARX1 I_11451 (I47270,I2507,I196981,I197219,);
DFFARX1 I_11452 (I197219,I2507,I196981,I197236,);
not I_11453 (I197244,I197236);
not I_11454 (I197261,I197219);
nand I_11455 (I196958,I197261,I197080);
nand I_11456 (I197292,I47261,I47261);
and I_11457 (I197309,I197292,I47273);
DFFARX1 I_11458 (I197309,I2507,I196981,I197335,);
nor I_11459 (I197343,I197335,I197007);
DFFARX1 I_11460 (I197343,I2507,I196981,I196946,);
DFFARX1 I_11461 (I197335,I2507,I196981,I196964,);
nor I_11462 (I197388,I47282,I47261);
not I_11463 (I197405,I197388);
nor I_11464 (I196967,I197244,I197405);
nand I_11465 (I196952,I197261,I197405);
nor I_11466 (I196961,I197007,I197388);
DFFARX1 I_11467 (I197388,I2507,I196981,I196970,);
not I_11468 (I197508,I2514);
DFFARX1 I_11469 (I709704,I2507,I197508,I197534,);
nand I_11470 (I197542,I709683,I709683);
and I_11471 (I197559,I197542,I709710);
DFFARX1 I_11472 (I197559,I2507,I197508,I197585,);
nor I_11473 (I197476,I197585,I197534);
not I_11474 (I197607,I197585);
DFFARX1 I_11475 (I709698,I2507,I197508,I197633,);
nand I_11476 (I197641,I197633,I709701);
not I_11477 (I197658,I197641);
DFFARX1 I_11478 (I197658,I2507,I197508,I197684,);
not I_11479 (I197500,I197684);
nor I_11480 (I197706,I197534,I197641);
nor I_11481 (I197482,I197585,I197706);
DFFARX1 I_11482 (I709692,I2507,I197508,I197746,);
DFFARX1 I_11483 (I197746,I2507,I197508,I197763,);
not I_11484 (I197771,I197763);
not I_11485 (I197788,I197746);
nand I_11486 (I197485,I197788,I197607);
nand I_11487 (I197819,I709689,I709686);
and I_11488 (I197836,I197819,I709707);
DFFARX1 I_11489 (I197836,I2507,I197508,I197862,);
nor I_11490 (I197870,I197862,I197534);
DFFARX1 I_11491 (I197870,I2507,I197508,I197473,);
DFFARX1 I_11492 (I197862,I2507,I197508,I197491,);
nor I_11493 (I197915,I709695,I709686);
not I_11494 (I197932,I197915);
nor I_11495 (I197494,I197771,I197932);
nand I_11496 (I197479,I197788,I197932);
nor I_11497 (I197488,I197534,I197915);
DFFARX1 I_11498 (I197915,I2507,I197508,I197497,);
not I_11499 (I198035,I2514);
DFFARX1 I_11500 (I19330,I2507,I198035,I198061,);
nand I_11501 (I198069,I19354,I19333);
and I_11502 (I198086,I198069,I19330);
DFFARX1 I_11503 (I198086,I2507,I198035,I198112,);
nor I_11504 (I198003,I198112,I198061);
not I_11505 (I198134,I198112);
DFFARX1 I_11506 (I19336,I2507,I198035,I198160,);
nand I_11507 (I198168,I198160,I19345);
not I_11508 (I198185,I198168);
DFFARX1 I_11509 (I198185,I2507,I198035,I198211,);
not I_11510 (I198027,I198211);
nor I_11511 (I198233,I198061,I198168);
nor I_11512 (I198009,I198112,I198233);
DFFARX1 I_11513 (I19339,I2507,I198035,I198273,);
DFFARX1 I_11514 (I198273,I2507,I198035,I198290,);
not I_11515 (I198298,I198290);
not I_11516 (I198315,I198273);
nand I_11517 (I198012,I198315,I198134);
nand I_11518 (I198346,I19351,I19333);
and I_11519 (I198363,I198346,I19342);
DFFARX1 I_11520 (I198363,I2507,I198035,I198389,);
nor I_11521 (I198397,I198389,I198061);
DFFARX1 I_11522 (I198397,I2507,I198035,I198000,);
DFFARX1 I_11523 (I198389,I2507,I198035,I198018,);
nor I_11524 (I198442,I19348,I19333);
not I_11525 (I198459,I198442);
nor I_11526 (I198021,I198298,I198459);
nand I_11527 (I198006,I198315,I198459);
nor I_11528 (I198015,I198061,I198442);
DFFARX1 I_11529 (I198442,I2507,I198035,I198024,);
not I_11530 (I198562,I2514);
DFFARX1 I_11531 (I483467,I2507,I198562,I198588,);
nand I_11532 (I198596,I483464,I483482);
and I_11533 (I198613,I198596,I483473);
DFFARX1 I_11534 (I198613,I2507,I198562,I198639,);
nor I_11535 (I198530,I198639,I198588);
not I_11536 (I198661,I198639);
DFFARX1 I_11537 (I483488,I2507,I198562,I198687,);
nand I_11538 (I198695,I198687,I483470);
not I_11539 (I198712,I198695);
DFFARX1 I_11540 (I198712,I2507,I198562,I198738,);
not I_11541 (I198554,I198738);
nor I_11542 (I198760,I198588,I198695);
nor I_11543 (I198536,I198639,I198760);
DFFARX1 I_11544 (I483476,I2507,I198562,I198800,);
DFFARX1 I_11545 (I198800,I2507,I198562,I198817,);
not I_11546 (I198825,I198817);
not I_11547 (I198842,I198800);
nand I_11548 (I198539,I198842,I198661);
nand I_11549 (I198873,I483464,I483491);
and I_11550 (I198890,I198873,I483479);
DFFARX1 I_11551 (I198890,I2507,I198562,I198916,);
nor I_11552 (I198924,I198916,I198588);
DFFARX1 I_11553 (I198924,I2507,I198562,I198527,);
DFFARX1 I_11554 (I198916,I2507,I198562,I198545,);
nor I_11555 (I198969,I483485,I483491);
not I_11556 (I198986,I198969);
nor I_11557 (I198548,I198825,I198986);
nand I_11558 (I198533,I198842,I198986);
nor I_11559 (I198542,I198588,I198969);
DFFARX1 I_11560 (I198969,I2507,I198562,I198551,);
not I_11561 (I199089,I2514);
DFFARX1 I_11562 (I460789,I2507,I199089,I199115,);
nand I_11563 (I199123,I460792,I460786);
and I_11564 (I199140,I199123,I460798);
DFFARX1 I_11565 (I199140,I2507,I199089,I199166,);
nor I_11566 (I199057,I199166,I199115);
not I_11567 (I199188,I199166);
DFFARX1 I_11568 (I460801,I2507,I199089,I199214,);
nand I_11569 (I199222,I199214,I460792);
not I_11570 (I199239,I199222);
DFFARX1 I_11571 (I199239,I2507,I199089,I199265,);
not I_11572 (I199081,I199265);
nor I_11573 (I199287,I199115,I199222);
nor I_11574 (I199063,I199166,I199287);
DFFARX1 I_11575 (I460804,I2507,I199089,I199327,);
DFFARX1 I_11576 (I199327,I2507,I199089,I199344,);
not I_11577 (I199352,I199344);
not I_11578 (I199369,I199327);
nand I_11579 (I199066,I199369,I199188);
nand I_11580 (I199400,I460786,I460795);
and I_11581 (I199417,I199400,I460789);
DFFARX1 I_11582 (I199417,I2507,I199089,I199443,);
nor I_11583 (I199451,I199443,I199115);
DFFARX1 I_11584 (I199451,I2507,I199089,I199054,);
DFFARX1 I_11585 (I199443,I2507,I199089,I199072,);
nor I_11586 (I199496,I460807,I460795);
not I_11587 (I199513,I199496);
nor I_11588 (I199075,I199352,I199513);
nand I_11589 (I199060,I199369,I199513);
nor I_11590 (I199069,I199115,I199496);
DFFARX1 I_11591 (I199496,I2507,I199089,I199078,);
not I_11592 (I199616,I2514);
DFFARX1 I_11593 (I96119,I2507,I199616,I199642,);
nand I_11594 (I199650,I96119,I96125);
and I_11595 (I199667,I199650,I96143);
DFFARX1 I_11596 (I199667,I2507,I199616,I199693,);
nor I_11597 (I199584,I199693,I199642);
not I_11598 (I199715,I199693);
DFFARX1 I_11599 (I96131,I2507,I199616,I199741,);
nand I_11600 (I199749,I199741,I96128);
not I_11601 (I199766,I199749);
DFFARX1 I_11602 (I199766,I2507,I199616,I199792,);
not I_11603 (I199608,I199792);
nor I_11604 (I199814,I199642,I199749);
nor I_11605 (I199590,I199693,I199814);
DFFARX1 I_11606 (I96137,I2507,I199616,I199854,);
DFFARX1 I_11607 (I199854,I2507,I199616,I199871,);
not I_11608 (I199879,I199871);
not I_11609 (I199896,I199854);
nand I_11610 (I199593,I199896,I199715);
nand I_11611 (I199927,I96122,I96122);
and I_11612 (I199944,I199927,I96134);
DFFARX1 I_11613 (I199944,I2507,I199616,I199970,);
nor I_11614 (I199978,I199970,I199642);
DFFARX1 I_11615 (I199978,I2507,I199616,I199581,);
DFFARX1 I_11616 (I199970,I2507,I199616,I199599,);
nor I_11617 (I200023,I96140,I96122);
not I_11618 (I200040,I200023);
nor I_11619 (I199602,I199879,I200040);
nand I_11620 (I199587,I199896,I200040);
nor I_11621 (I199596,I199642,I200023);
DFFARX1 I_11622 (I200023,I2507,I199616,I199605,);
not I_11623 (I200143,I2514);
DFFARX1 I_11624 (I100284,I2507,I200143,I200169,);
nand I_11625 (I200177,I100284,I100290);
and I_11626 (I200194,I200177,I100308);
DFFARX1 I_11627 (I200194,I2507,I200143,I200220,);
nor I_11628 (I200111,I200220,I200169);
not I_11629 (I200242,I200220);
DFFARX1 I_11630 (I100296,I2507,I200143,I200268,);
nand I_11631 (I200276,I200268,I100293);
not I_11632 (I200293,I200276);
DFFARX1 I_11633 (I200293,I2507,I200143,I200319,);
not I_11634 (I200135,I200319);
nor I_11635 (I200341,I200169,I200276);
nor I_11636 (I200117,I200220,I200341);
DFFARX1 I_11637 (I100302,I2507,I200143,I200381,);
DFFARX1 I_11638 (I200381,I2507,I200143,I200398,);
not I_11639 (I200406,I200398);
not I_11640 (I200423,I200381);
nand I_11641 (I200120,I200423,I200242);
nand I_11642 (I200454,I100287,I100287);
and I_11643 (I200471,I200454,I100299);
DFFARX1 I_11644 (I200471,I2507,I200143,I200497,);
nor I_11645 (I200505,I200497,I200169);
DFFARX1 I_11646 (I200505,I2507,I200143,I200108,);
DFFARX1 I_11647 (I200497,I2507,I200143,I200126,);
nor I_11648 (I200550,I100305,I100287);
not I_11649 (I200567,I200550);
nor I_11650 (I200129,I200406,I200567);
nand I_11651 (I200114,I200423,I200567);
nor I_11652 (I200123,I200169,I200550);
DFFARX1 I_11653 (I200550,I2507,I200143,I200132,);
not I_11654 (I200670,I2514);
DFFARX1 I_11655 (I298031,I2507,I200670,I200696,);
nand I_11656 (I200704,I298031,I298043);
and I_11657 (I200721,I200704,I298028);
DFFARX1 I_11658 (I200721,I2507,I200670,I200747,);
nor I_11659 (I200638,I200747,I200696);
not I_11660 (I200769,I200747);
DFFARX1 I_11661 (I298052,I2507,I200670,I200795,);
nand I_11662 (I200803,I200795,I298049);
not I_11663 (I200820,I200803);
DFFARX1 I_11664 (I200820,I2507,I200670,I200846,);
not I_11665 (I200662,I200846);
nor I_11666 (I200868,I200696,I200803);
nor I_11667 (I200644,I200747,I200868);
DFFARX1 I_11668 (I298040,I2507,I200670,I200908,);
DFFARX1 I_11669 (I200908,I2507,I200670,I200925,);
not I_11670 (I200933,I200925);
not I_11671 (I200950,I200908);
nand I_11672 (I200647,I200950,I200769);
nand I_11673 (I200981,I298028,I298037);
and I_11674 (I200998,I200981,I298046);
DFFARX1 I_11675 (I200998,I2507,I200670,I201024,);
nor I_11676 (I201032,I201024,I200696);
DFFARX1 I_11677 (I201032,I2507,I200670,I200635,);
DFFARX1 I_11678 (I201024,I2507,I200670,I200653,);
nor I_11679 (I201077,I298034,I298037);
not I_11680 (I201094,I201077);
nor I_11681 (I200656,I200933,I201094);
nand I_11682 (I200641,I200950,I201094);
nor I_11683 (I200650,I200696,I201077);
DFFARX1 I_11684 (I201077,I2507,I200670,I200659,);
not I_11685 (I201197,I2514);
DFFARX1 I_11686 (I420083,I2507,I201197,I201223,);
nand I_11687 (I201231,I420074,I420089);
and I_11688 (I201248,I201231,I420095);
DFFARX1 I_11689 (I201248,I2507,I201197,I201274,);
nor I_11690 (I201165,I201274,I201223);
not I_11691 (I201296,I201274);
DFFARX1 I_11692 (I420080,I2507,I201197,I201322,);
nand I_11693 (I201330,I201322,I420074);
not I_11694 (I201347,I201330);
DFFARX1 I_11695 (I201347,I2507,I201197,I201373,);
not I_11696 (I201189,I201373);
nor I_11697 (I201395,I201223,I201330);
nor I_11698 (I201171,I201274,I201395);
DFFARX1 I_11699 (I420077,I2507,I201197,I201435,);
DFFARX1 I_11700 (I201435,I2507,I201197,I201452,);
not I_11701 (I201460,I201452);
not I_11702 (I201477,I201435);
nand I_11703 (I201174,I201477,I201296);
nand I_11704 (I201508,I420071,I420086);
and I_11705 (I201525,I201508,I420071);
DFFARX1 I_11706 (I201525,I2507,I201197,I201551,);
nor I_11707 (I201559,I201551,I201223);
DFFARX1 I_11708 (I201559,I2507,I201197,I201162,);
DFFARX1 I_11709 (I201551,I2507,I201197,I201180,);
nor I_11710 (I201604,I420092,I420086);
not I_11711 (I201621,I201604);
nor I_11712 (I201183,I201460,I201621);
nand I_11713 (I201168,I201477,I201621);
nor I_11714 (I201177,I201223,I201604);
DFFARX1 I_11715 (I201604,I2507,I201197,I201186,);
not I_11716 (I201724,I2514);
DFFARX1 I_11717 (I608669,I2507,I201724,I201750,);
nand I_11718 (I201758,I608684,I608669);
and I_11719 (I201775,I201758,I608687);
DFFARX1 I_11720 (I201775,I2507,I201724,I201801,);
nor I_11721 (I201692,I201801,I201750);
not I_11722 (I201823,I201801);
DFFARX1 I_11723 (I608693,I2507,I201724,I201849,);
nand I_11724 (I201857,I201849,I608675);
not I_11725 (I201874,I201857);
DFFARX1 I_11726 (I201874,I2507,I201724,I201900,);
not I_11727 (I201716,I201900);
nor I_11728 (I201922,I201750,I201857);
nor I_11729 (I201698,I201801,I201922);
DFFARX1 I_11730 (I608672,I2507,I201724,I201962,);
DFFARX1 I_11731 (I201962,I2507,I201724,I201979,);
not I_11732 (I201987,I201979);
not I_11733 (I202004,I201962);
nand I_11734 (I201701,I202004,I201823);
nand I_11735 (I202035,I608672,I608678);
and I_11736 (I202052,I202035,I608690);
DFFARX1 I_11737 (I202052,I2507,I201724,I202078,);
nor I_11738 (I202086,I202078,I201750);
DFFARX1 I_11739 (I202086,I2507,I201724,I201689,);
DFFARX1 I_11740 (I202078,I2507,I201724,I201707,);
nor I_11741 (I202131,I608681,I608678);
not I_11742 (I202148,I202131);
nor I_11743 (I201710,I201987,I202148);
nand I_11744 (I201695,I202004,I202148);
nor I_11745 (I201704,I201750,I202131);
DFFARX1 I_11746 (I202131,I2507,I201724,I201713,);
not I_11747 (I202251,I2514);
DFFARX1 I_11748 (I470275,I2507,I202251,I202277,);
nand I_11749 (I202285,I470278,I470272);
and I_11750 (I202302,I202285,I470284);
DFFARX1 I_11751 (I202302,I2507,I202251,I202328,);
nor I_11752 (I202219,I202328,I202277);
not I_11753 (I202350,I202328);
DFFARX1 I_11754 (I470287,I2507,I202251,I202376,);
nand I_11755 (I202384,I202376,I470278);
not I_11756 (I202401,I202384);
DFFARX1 I_11757 (I202401,I2507,I202251,I202427,);
not I_11758 (I202243,I202427);
nor I_11759 (I202449,I202277,I202384);
nor I_11760 (I202225,I202328,I202449);
DFFARX1 I_11761 (I470290,I2507,I202251,I202489,);
DFFARX1 I_11762 (I202489,I2507,I202251,I202506,);
not I_11763 (I202514,I202506);
not I_11764 (I202531,I202489);
nand I_11765 (I202228,I202531,I202350);
nand I_11766 (I202562,I470272,I470281);
and I_11767 (I202579,I202562,I470275);
DFFARX1 I_11768 (I202579,I2507,I202251,I202605,);
nor I_11769 (I202613,I202605,I202277);
DFFARX1 I_11770 (I202613,I2507,I202251,I202216,);
DFFARX1 I_11771 (I202605,I2507,I202251,I202234,);
nor I_11772 (I202658,I470293,I470281);
not I_11773 (I202675,I202658);
nor I_11774 (I202237,I202514,I202675);
nand I_11775 (I202222,I202531,I202675);
nor I_11776 (I202231,I202277,I202658);
DFFARX1 I_11777 (I202658,I2507,I202251,I202240,);
not I_11778 (I202778,I2514);
DFFARX1 I_11779 (I677500,I2507,I202778,I202804,);
nand I_11780 (I202812,I677497,I677488);
and I_11781 (I202829,I202812,I677485);
DFFARX1 I_11782 (I202829,I2507,I202778,I202855,);
nor I_11783 (I202746,I202855,I202804);
not I_11784 (I202877,I202855);
DFFARX1 I_11785 (I677494,I2507,I202778,I202903,);
nand I_11786 (I202911,I202903,I677503);
not I_11787 (I202928,I202911);
DFFARX1 I_11788 (I202928,I2507,I202778,I202954,);
not I_11789 (I202770,I202954);
nor I_11790 (I202976,I202804,I202911);
nor I_11791 (I202752,I202855,I202976);
DFFARX1 I_11792 (I677506,I2507,I202778,I203016,);
DFFARX1 I_11793 (I203016,I2507,I202778,I203033,);
not I_11794 (I203041,I203033);
not I_11795 (I203058,I203016);
nand I_11796 (I202755,I203058,I202877);
nand I_11797 (I203089,I677485,I677491);
and I_11798 (I203106,I203089,I677509);
DFFARX1 I_11799 (I203106,I2507,I202778,I203132,);
nor I_11800 (I203140,I203132,I202804);
DFFARX1 I_11801 (I203140,I2507,I202778,I202743,);
DFFARX1 I_11802 (I203132,I2507,I202778,I202761,);
nor I_11803 (I203185,I677488,I677491);
not I_11804 (I203202,I203185);
nor I_11805 (I202764,I203041,I203202);
nand I_11806 (I202749,I203058,I203202);
nor I_11807 (I202758,I202804,I203185);
DFFARX1 I_11808 (I203185,I2507,I202778,I202767,);
not I_11809 (I203305,I2514);
DFFARX1 I_11810 (I323560,I2507,I203305,I203331,);
nand I_11811 (I203339,I323545,I323548);
and I_11812 (I203356,I203339,I323563);
DFFARX1 I_11813 (I203356,I2507,I203305,I203382,);
nor I_11814 (I203273,I203382,I203331);
not I_11815 (I203404,I203382);
DFFARX1 I_11816 (I323557,I2507,I203305,I203430,);
nand I_11817 (I203438,I203430,I323548);
not I_11818 (I203455,I203438);
DFFARX1 I_11819 (I203455,I2507,I203305,I203481,);
not I_11820 (I203297,I203481);
nor I_11821 (I203503,I203331,I203438);
nor I_11822 (I203279,I203382,I203503);
DFFARX1 I_11823 (I323554,I2507,I203305,I203543,);
DFFARX1 I_11824 (I203543,I2507,I203305,I203560,);
not I_11825 (I203568,I203560);
not I_11826 (I203585,I203543);
nand I_11827 (I203282,I203585,I203404);
nand I_11828 (I203616,I323569,I323545);
and I_11829 (I203633,I203616,I323566);
DFFARX1 I_11830 (I203633,I2507,I203305,I203659,);
nor I_11831 (I203667,I203659,I203331);
DFFARX1 I_11832 (I203667,I2507,I203305,I203270,);
DFFARX1 I_11833 (I203659,I2507,I203305,I203288,);
nor I_11834 (I203712,I323551,I323545);
not I_11835 (I203729,I203712);
nor I_11836 (I203291,I203568,I203729);
nand I_11837 (I203276,I203585,I203729);
nor I_11838 (I203285,I203331,I203712);
DFFARX1 I_11839 (I203712,I2507,I203305,I203294,);
not I_11840 (I203832,I2514);
DFFARX1 I_11841 (I396963,I2507,I203832,I203858,);
nand I_11842 (I203866,I396954,I396969);
and I_11843 (I203883,I203866,I396975);
DFFARX1 I_11844 (I203883,I2507,I203832,I203909,);
nor I_11845 (I203800,I203909,I203858);
not I_11846 (I203931,I203909);
DFFARX1 I_11847 (I396960,I2507,I203832,I203957,);
nand I_11848 (I203965,I203957,I396954);
not I_11849 (I203982,I203965);
DFFARX1 I_11850 (I203982,I2507,I203832,I204008,);
not I_11851 (I203824,I204008);
nor I_11852 (I204030,I203858,I203965);
nor I_11853 (I203806,I203909,I204030);
DFFARX1 I_11854 (I396957,I2507,I203832,I204070,);
DFFARX1 I_11855 (I204070,I2507,I203832,I204087,);
not I_11856 (I204095,I204087);
not I_11857 (I204112,I204070);
nand I_11858 (I203809,I204112,I203931);
nand I_11859 (I204143,I396951,I396966);
and I_11860 (I204160,I204143,I396951);
DFFARX1 I_11861 (I204160,I2507,I203832,I204186,);
nor I_11862 (I204194,I204186,I203858);
DFFARX1 I_11863 (I204194,I2507,I203832,I203797,);
DFFARX1 I_11864 (I204186,I2507,I203832,I203815,);
nor I_11865 (I204239,I396972,I396966);
not I_11866 (I204256,I204239);
nor I_11867 (I203818,I204095,I204256);
nand I_11868 (I203803,I204112,I204256);
nor I_11869 (I203812,I203858,I204239);
DFFARX1 I_11870 (I204239,I2507,I203832,I203821,);
not I_11871 (I204359,I2514);
DFFARX1 I_11872 (I81519,I2507,I204359,I204385,);
nand I_11873 (I204393,I81531,I81540);
and I_11874 (I204410,I204393,I81519);
DFFARX1 I_11875 (I204410,I2507,I204359,I204436,);
nor I_11876 (I204327,I204436,I204385);
not I_11877 (I204458,I204436);
DFFARX1 I_11878 (I81534,I2507,I204359,I204484,);
nand I_11879 (I204492,I204484,I81522);
not I_11880 (I204509,I204492);
DFFARX1 I_11881 (I204509,I2507,I204359,I204535,);
not I_11882 (I204351,I204535);
nor I_11883 (I204557,I204385,I204492);
nor I_11884 (I204333,I204436,I204557);
DFFARX1 I_11885 (I81525,I2507,I204359,I204597,);
DFFARX1 I_11886 (I204597,I2507,I204359,I204614,);
not I_11887 (I204622,I204614);
not I_11888 (I204639,I204597);
nand I_11889 (I204336,I204639,I204458);
nand I_11890 (I204670,I81516,I81516);
and I_11891 (I204687,I204670,I81528);
DFFARX1 I_11892 (I204687,I2507,I204359,I204713,);
nor I_11893 (I204721,I204713,I204385);
DFFARX1 I_11894 (I204721,I2507,I204359,I204324,);
DFFARX1 I_11895 (I204713,I2507,I204359,I204342,);
nor I_11896 (I204766,I81537,I81516);
not I_11897 (I204783,I204766);
nor I_11898 (I204345,I204622,I204783);
nand I_11899 (I204330,I204639,I204783);
nor I_11900 (I204339,I204385,I204766);
DFFARX1 I_11901 (I204766,I2507,I204359,I204348,);
not I_11902 (I204886,I2514);
DFFARX1 I_11903 (I131224,I2507,I204886,I204912,);
nand I_11904 (I204920,I131224,I131230);
and I_11905 (I204937,I204920,I131248);
DFFARX1 I_11906 (I204937,I2507,I204886,I204963,);
nor I_11907 (I204854,I204963,I204912);
not I_11908 (I204985,I204963);
DFFARX1 I_11909 (I131236,I2507,I204886,I205011,);
nand I_11910 (I205019,I205011,I131233);
not I_11911 (I205036,I205019);
DFFARX1 I_11912 (I205036,I2507,I204886,I205062,);
not I_11913 (I204878,I205062);
nor I_11914 (I205084,I204912,I205019);
nor I_11915 (I204860,I204963,I205084);
DFFARX1 I_11916 (I131242,I2507,I204886,I205124,);
DFFARX1 I_11917 (I205124,I2507,I204886,I205141,);
not I_11918 (I205149,I205141);
not I_11919 (I205166,I205124);
nand I_11920 (I204863,I205166,I204985);
nand I_11921 (I205197,I131227,I131227);
and I_11922 (I205214,I205197,I131239);
DFFARX1 I_11923 (I205214,I2507,I204886,I205240,);
nor I_11924 (I205248,I205240,I204912);
DFFARX1 I_11925 (I205248,I2507,I204886,I204851,);
DFFARX1 I_11926 (I205240,I2507,I204886,I204869,);
nor I_11927 (I205293,I131245,I131227);
not I_11928 (I205310,I205293);
nor I_11929 (I204872,I205149,I205310);
nand I_11930 (I204857,I205166,I205310);
nor I_11931 (I204866,I204912,I205293);
DFFARX1 I_11932 (I205293,I2507,I204886,I204875,);
not I_11933 (I205413,I2514);
DFFARX1 I_11934 (I379623,I2507,I205413,I205439,);
nand I_11935 (I205447,I379614,I379629);
and I_11936 (I205464,I205447,I379635);
DFFARX1 I_11937 (I205464,I2507,I205413,I205490,);
nor I_11938 (I205381,I205490,I205439);
not I_11939 (I205512,I205490);
DFFARX1 I_11940 (I379620,I2507,I205413,I205538,);
nand I_11941 (I205546,I205538,I379614);
not I_11942 (I205563,I205546);
DFFARX1 I_11943 (I205563,I2507,I205413,I205589,);
not I_11944 (I205405,I205589);
nor I_11945 (I205611,I205439,I205546);
nor I_11946 (I205387,I205490,I205611);
DFFARX1 I_11947 (I379617,I2507,I205413,I205651,);
DFFARX1 I_11948 (I205651,I2507,I205413,I205668,);
not I_11949 (I205676,I205668);
not I_11950 (I205693,I205651);
nand I_11951 (I205390,I205693,I205512);
nand I_11952 (I205724,I379611,I379626);
and I_11953 (I205741,I205724,I379611);
DFFARX1 I_11954 (I205741,I2507,I205413,I205767,);
nor I_11955 (I205775,I205767,I205439);
DFFARX1 I_11956 (I205775,I2507,I205413,I205378,);
DFFARX1 I_11957 (I205767,I2507,I205413,I205396,);
nor I_11958 (I205820,I379632,I379626);
not I_11959 (I205837,I205820);
nor I_11960 (I205399,I205676,I205837);
nand I_11961 (I205384,I205693,I205837);
nor I_11962 (I205393,I205439,I205820);
DFFARX1 I_11963 (I205820,I2507,I205413,I205402,);
not I_11964 (I205940,I2514);
DFFARX1 I_11965 (I450776,I2507,I205940,I205966,);
nand I_11966 (I205974,I450779,I450773);
and I_11967 (I205991,I205974,I450785);
DFFARX1 I_11968 (I205991,I2507,I205940,I206017,);
nor I_11969 (I205908,I206017,I205966);
not I_11970 (I206039,I206017);
DFFARX1 I_11971 (I450788,I2507,I205940,I206065,);
nand I_11972 (I206073,I206065,I450779);
not I_11973 (I206090,I206073);
DFFARX1 I_11974 (I206090,I2507,I205940,I206116,);
not I_11975 (I205932,I206116);
nor I_11976 (I206138,I205966,I206073);
nor I_11977 (I205914,I206017,I206138);
DFFARX1 I_11978 (I450791,I2507,I205940,I206178,);
DFFARX1 I_11979 (I206178,I2507,I205940,I206195,);
not I_11980 (I206203,I206195);
not I_11981 (I206220,I206178);
nand I_11982 (I205917,I206220,I206039);
nand I_11983 (I206251,I450773,I450782);
and I_11984 (I206268,I206251,I450776);
DFFARX1 I_11985 (I206268,I2507,I205940,I206294,);
nor I_11986 (I206302,I206294,I205966);
DFFARX1 I_11987 (I206302,I2507,I205940,I205905,);
DFFARX1 I_11988 (I206294,I2507,I205940,I205923,);
nor I_11989 (I206347,I450794,I450782);
not I_11990 (I206364,I206347);
nor I_11991 (I205926,I206203,I206364);
nand I_11992 (I205911,I206220,I206364);
nor I_11993 (I205920,I205966,I206347);
DFFARX1 I_11994 (I206347,I2507,I205940,I205929,);
not I_11995 (I206467,I2514);
DFFARX1 I_11996 (I604623,I2507,I206467,I206493,);
nand I_11997 (I206501,I604638,I604623);
and I_11998 (I206518,I206501,I604641);
DFFARX1 I_11999 (I206518,I2507,I206467,I206544,);
nor I_12000 (I206435,I206544,I206493);
not I_12001 (I206566,I206544);
DFFARX1 I_12002 (I604647,I2507,I206467,I206592,);
nand I_12003 (I206600,I206592,I604629);
not I_12004 (I206617,I206600);
DFFARX1 I_12005 (I206617,I2507,I206467,I206643,);
not I_12006 (I206459,I206643);
nor I_12007 (I206665,I206493,I206600);
nor I_12008 (I206441,I206544,I206665);
DFFARX1 I_12009 (I604626,I2507,I206467,I206705,);
DFFARX1 I_12010 (I206705,I2507,I206467,I206722,);
not I_12011 (I206730,I206722);
not I_12012 (I206747,I206705);
nand I_12013 (I206444,I206747,I206566);
nand I_12014 (I206778,I604626,I604632);
and I_12015 (I206795,I206778,I604644);
DFFARX1 I_12016 (I206795,I2507,I206467,I206821,);
nor I_12017 (I206829,I206821,I206493);
DFFARX1 I_12018 (I206829,I2507,I206467,I206432,);
DFFARX1 I_12019 (I206821,I2507,I206467,I206450,);
nor I_12020 (I206874,I604635,I604632);
not I_12021 (I206891,I206874);
nor I_12022 (I206453,I206730,I206891);
nand I_12023 (I206438,I206747,I206891);
nor I_12024 (I206447,I206493,I206874);
DFFARX1 I_12025 (I206874,I2507,I206467,I206456,);
not I_12026 (I206994,I2514);
DFFARX1 I_12027 (I465005,I2507,I206994,I207020,);
nand I_12028 (I207028,I465008,I465002);
and I_12029 (I207045,I207028,I465014);
DFFARX1 I_12030 (I207045,I2507,I206994,I207071,);
nor I_12031 (I206962,I207071,I207020);
not I_12032 (I207093,I207071);
DFFARX1 I_12033 (I465017,I2507,I206994,I207119,);
nand I_12034 (I207127,I207119,I465008);
not I_12035 (I207144,I207127);
DFFARX1 I_12036 (I207144,I2507,I206994,I207170,);
not I_12037 (I206986,I207170);
nor I_12038 (I207192,I207020,I207127);
nor I_12039 (I206968,I207071,I207192);
DFFARX1 I_12040 (I465020,I2507,I206994,I207232,);
DFFARX1 I_12041 (I207232,I2507,I206994,I207249,);
not I_12042 (I207257,I207249);
not I_12043 (I207274,I207232);
nand I_12044 (I206971,I207274,I207093);
nand I_12045 (I207305,I465002,I465011);
and I_12046 (I207322,I207305,I465005);
DFFARX1 I_12047 (I207322,I2507,I206994,I207348,);
nor I_12048 (I207356,I207348,I207020);
DFFARX1 I_12049 (I207356,I2507,I206994,I206959,);
DFFARX1 I_12050 (I207348,I2507,I206994,I206977,);
nor I_12051 (I207401,I465023,I465011);
not I_12052 (I207418,I207401);
nor I_12053 (I206980,I207257,I207418);
nand I_12054 (I206965,I207274,I207418);
nor I_12055 (I206974,I207020,I207401);
DFFARX1 I_12056 (I207401,I2507,I206994,I206983,);
not I_12057 (I207521,I2514);
DFFARX1 I_12058 (I439182,I2507,I207521,I207547,);
nand I_12059 (I207555,I439185,I439179);
and I_12060 (I207572,I207555,I439191);
DFFARX1 I_12061 (I207572,I2507,I207521,I207598,);
nor I_12062 (I207489,I207598,I207547);
not I_12063 (I207620,I207598);
DFFARX1 I_12064 (I439194,I2507,I207521,I207646,);
nand I_12065 (I207654,I207646,I439185);
not I_12066 (I207671,I207654);
DFFARX1 I_12067 (I207671,I2507,I207521,I207697,);
not I_12068 (I207513,I207697);
nor I_12069 (I207719,I207547,I207654);
nor I_12070 (I207495,I207598,I207719);
DFFARX1 I_12071 (I439197,I2507,I207521,I207759,);
DFFARX1 I_12072 (I207759,I2507,I207521,I207776,);
not I_12073 (I207784,I207776);
not I_12074 (I207801,I207759);
nand I_12075 (I207498,I207801,I207620);
nand I_12076 (I207832,I439179,I439188);
and I_12077 (I207849,I207832,I439182);
DFFARX1 I_12078 (I207849,I2507,I207521,I207875,);
nor I_12079 (I207883,I207875,I207547);
DFFARX1 I_12080 (I207883,I2507,I207521,I207486,);
DFFARX1 I_12081 (I207875,I2507,I207521,I207504,);
nor I_12082 (I207928,I439200,I439188);
not I_12083 (I207945,I207928);
nor I_12084 (I207507,I207784,I207945);
nand I_12085 (I207492,I207801,I207945);
nor I_12086 (I207501,I207547,I207928);
DFFARX1 I_12087 (I207928,I2507,I207521,I207510,);
not I_12088 (I208048,I2514);
DFFARX1 I_12089 (I436020,I2507,I208048,I208074,);
nand I_12090 (I208082,I436023,I436017);
and I_12091 (I208099,I208082,I436029);
DFFARX1 I_12092 (I208099,I2507,I208048,I208125,);
nor I_12093 (I208016,I208125,I208074);
not I_12094 (I208147,I208125);
DFFARX1 I_12095 (I436032,I2507,I208048,I208173,);
nand I_12096 (I208181,I208173,I436023);
not I_12097 (I208198,I208181);
DFFARX1 I_12098 (I208198,I2507,I208048,I208224,);
not I_12099 (I208040,I208224);
nor I_12100 (I208246,I208074,I208181);
nor I_12101 (I208022,I208125,I208246);
DFFARX1 I_12102 (I436035,I2507,I208048,I208286,);
DFFARX1 I_12103 (I208286,I2507,I208048,I208303,);
not I_12104 (I208311,I208303);
not I_12105 (I208328,I208286);
nand I_12106 (I208025,I208328,I208147);
nand I_12107 (I208359,I436017,I436026);
and I_12108 (I208376,I208359,I436020);
DFFARX1 I_12109 (I208376,I2507,I208048,I208402,);
nor I_12110 (I208410,I208402,I208074);
DFFARX1 I_12111 (I208410,I2507,I208048,I208013,);
DFFARX1 I_12112 (I208402,I2507,I208048,I208031,);
nor I_12113 (I208455,I436038,I436026);
not I_12114 (I208472,I208455);
nor I_12115 (I208034,I208311,I208472);
nand I_12116 (I208019,I208328,I208472);
nor I_12117 (I208028,I208074,I208455);
DFFARX1 I_12118 (I208455,I2507,I208048,I208037,);
not I_12119 (I208575,I2514);
DFFARX1 I_12120 (I569402,I2507,I208575,I208601,);
nand I_12121 (I208609,I569399,I569402);
and I_12122 (I208626,I208609,I569411);
DFFARX1 I_12123 (I208626,I2507,I208575,I208652,);
nor I_12124 (I208543,I208652,I208601);
not I_12125 (I208674,I208652);
DFFARX1 I_12126 (I569399,I2507,I208575,I208700,);
nand I_12127 (I208708,I208700,I569417);
not I_12128 (I208725,I208708);
DFFARX1 I_12129 (I208725,I2507,I208575,I208751,);
not I_12130 (I208567,I208751);
nor I_12131 (I208773,I208601,I208708);
nor I_12132 (I208549,I208652,I208773);
DFFARX1 I_12133 (I569405,I2507,I208575,I208813,);
DFFARX1 I_12134 (I208813,I2507,I208575,I208830,);
not I_12135 (I208838,I208830);
not I_12136 (I208855,I208813);
nand I_12137 (I208552,I208855,I208674);
nand I_12138 (I208886,I569414,I569420);
and I_12139 (I208903,I208886,I569405);
DFFARX1 I_12140 (I208903,I2507,I208575,I208929,);
nor I_12141 (I208937,I208929,I208601);
DFFARX1 I_12142 (I208937,I2507,I208575,I208540,);
DFFARX1 I_12143 (I208929,I2507,I208575,I208558,);
nor I_12144 (I208982,I569408,I569420);
not I_12145 (I208999,I208982);
nor I_12146 (I208561,I208838,I208999);
nand I_12147 (I208546,I208855,I208999);
nor I_12148 (I208555,I208601,I208982);
DFFARX1 I_12149 (I208982,I2507,I208575,I208564,);
not I_12150 (I209102,I2514);
DFFARX1 I_12151 (I368063,I2507,I209102,I209128,);
nand I_12152 (I209136,I368054,I368069);
and I_12153 (I209153,I209136,I368075);
DFFARX1 I_12154 (I209153,I2507,I209102,I209179,);
nor I_12155 (I209070,I209179,I209128);
not I_12156 (I209201,I209179);
DFFARX1 I_12157 (I368060,I2507,I209102,I209227,);
nand I_12158 (I209235,I209227,I368054);
not I_12159 (I209252,I209235);
DFFARX1 I_12160 (I209252,I2507,I209102,I209278,);
not I_12161 (I209094,I209278);
nor I_12162 (I209300,I209128,I209235);
nor I_12163 (I209076,I209179,I209300);
DFFARX1 I_12164 (I368057,I2507,I209102,I209340,);
DFFARX1 I_12165 (I209340,I2507,I209102,I209357,);
not I_12166 (I209365,I209357);
not I_12167 (I209382,I209340);
nand I_12168 (I209079,I209382,I209201);
nand I_12169 (I209413,I368051,I368066);
and I_12170 (I209430,I209413,I368051);
DFFARX1 I_12171 (I209430,I2507,I209102,I209456,);
nor I_12172 (I209464,I209456,I209128);
DFFARX1 I_12173 (I209464,I2507,I209102,I209067,);
DFFARX1 I_12174 (I209456,I2507,I209102,I209085,);
nor I_12175 (I209509,I368072,I368066);
not I_12176 (I209526,I209509);
nor I_12177 (I209088,I209365,I209526);
nand I_12178 (I209073,I209382,I209526);
nor I_12179 (I209082,I209128,I209509);
DFFARX1 I_12180 (I209509,I2507,I209102,I209091,);
not I_12181 (I209629,I2514);
DFFARX1 I_12182 (I429696,I2507,I209629,I209655,);
nand I_12183 (I209663,I429699,I429693);
and I_12184 (I209680,I209663,I429705);
DFFARX1 I_12185 (I209680,I2507,I209629,I209706,);
nor I_12186 (I209597,I209706,I209655);
not I_12187 (I209728,I209706);
DFFARX1 I_12188 (I429708,I2507,I209629,I209754,);
nand I_12189 (I209762,I209754,I429699);
not I_12190 (I209779,I209762);
DFFARX1 I_12191 (I209779,I2507,I209629,I209805,);
not I_12192 (I209621,I209805);
nor I_12193 (I209827,I209655,I209762);
nor I_12194 (I209603,I209706,I209827);
DFFARX1 I_12195 (I429711,I2507,I209629,I209867,);
DFFARX1 I_12196 (I209867,I2507,I209629,I209884,);
not I_12197 (I209892,I209884);
not I_12198 (I209909,I209867);
nand I_12199 (I209606,I209909,I209728);
nand I_12200 (I209940,I429693,I429702);
and I_12201 (I209957,I209940,I429696);
DFFARX1 I_12202 (I209957,I2507,I209629,I209983,);
nor I_12203 (I209991,I209983,I209655);
DFFARX1 I_12204 (I209991,I2507,I209629,I209594,);
DFFARX1 I_12205 (I209983,I2507,I209629,I209612,);
nor I_12206 (I210036,I429714,I429702);
not I_12207 (I210053,I210036);
nor I_12208 (I209615,I209892,I210053);
nand I_12209 (I209600,I209909,I210053);
nor I_12210 (I209609,I209655,I210036);
DFFARX1 I_12211 (I210036,I2507,I209629,I209618,);
not I_12212 (I210156,I2514);
DFFARX1 I_12213 (I606357,I2507,I210156,I210182,);
nand I_12214 (I210190,I606372,I606357);
and I_12215 (I210207,I210190,I606375);
DFFARX1 I_12216 (I210207,I2507,I210156,I210233,);
nor I_12217 (I210124,I210233,I210182);
not I_12218 (I210255,I210233);
DFFARX1 I_12219 (I606381,I2507,I210156,I210281,);
nand I_12220 (I210289,I210281,I606363);
not I_12221 (I210306,I210289);
DFFARX1 I_12222 (I210306,I2507,I210156,I210332,);
not I_12223 (I210148,I210332);
nor I_12224 (I210354,I210182,I210289);
nor I_12225 (I210130,I210233,I210354);
DFFARX1 I_12226 (I606360,I2507,I210156,I210394,);
DFFARX1 I_12227 (I210394,I2507,I210156,I210411,);
not I_12228 (I210419,I210411);
not I_12229 (I210436,I210394);
nand I_12230 (I210133,I210436,I210255);
nand I_12231 (I210467,I606360,I606366);
and I_12232 (I210484,I210467,I606378);
DFFARX1 I_12233 (I210484,I2507,I210156,I210510,);
nor I_12234 (I210518,I210510,I210182);
DFFARX1 I_12235 (I210518,I2507,I210156,I210121,);
DFFARX1 I_12236 (I210510,I2507,I210156,I210139,);
nor I_12237 (I210563,I606369,I606366);
not I_12238 (I210580,I210563);
nor I_12239 (I210142,I210419,I210580);
nand I_12240 (I210127,I210436,I210580);
nor I_12241 (I210136,I210182,I210563);
DFFARX1 I_12242 (I210563,I2507,I210156,I210145,);
not I_12243 (I210683,I2514);
DFFARX1 I_12244 (I653975,I2507,I210683,I210709,);
nand I_12245 (I210717,I653957,I653981);
and I_12246 (I210734,I210717,I653972);
DFFARX1 I_12247 (I210734,I2507,I210683,I210760,);
nor I_12248 (I210651,I210760,I210709);
not I_12249 (I210782,I210760);
DFFARX1 I_12250 (I653978,I2507,I210683,I210808,);
nand I_12251 (I210816,I210808,I653966);
not I_12252 (I210833,I210816);
DFFARX1 I_12253 (I210833,I2507,I210683,I210859,);
not I_12254 (I210675,I210859);
nor I_12255 (I210881,I210709,I210816);
nor I_12256 (I210657,I210760,I210881);
DFFARX1 I_12257 (I653957,I2507,I210683,I210921,);
DFFARX1 I_12258 (I210921,I2507,I210683,I210938,);
not I_12259 (I210946,I210938);
not I_12260 (I210963,I210921);
nand I_12261 (I210660,I210963,I210782);
nand I_12262 (I210994,I653963,I653960);
and I_12263 (I211011,I210994,I653969);
DFFARX1 I_12264 (I211011,I2507,I210683,I211037,);
nor I_12265 (I211045,I211037,I210709);
DFFARX1 I_12266 (I211045,I2507,I210683,I210648,);
DFFARX1 I_12267 (I211037,I2507,I210683,I210666,);
nor I_12268 (I211090,I653960,I653960);
not I_12269 (I211107,I211090);
nor I_12270 (I210669,I210946,I211107);
nand I_12271 (I210654,I210963,I211107);
nor I_12272 (I210663,I210709,I211090);
DFFARX1 I_12273 (I211090,I2507,I210683,I210672,);
not I_12274 (I211210,I2514);
DFFARX1 I_12275 (I282561,I2507,I211210,I211236,);
nand I_12276 (I211244,I282561,I282573);
and I_12277 (I211261,I211244,I282558);
DFFARX1 I_12278 (I211261,I2507,I211210,I211287,);
nor I_12279 (I211178,I211287,I211236);
not I_12280 (I211309,I211287);
DFFARX1 I_12281 (I282582,I2507,I211210,I211335,);
nand I_12282 (I211343,I211335,I282579);
not I_12283 (I211360,I211343);
DFFARX1 I_12284 (I211360,I2507,I211210,I211386,);
not I_12285 (I211202,I211386);
nor I_12286 (I211408,I211236,I211343);
nor I_12287 (I211184,I211287,I211408);
DFFARX1 I_12288 (I282570,I2507,I211210,I211448,);
DFFARX1 I_12289 (I211448,I2507,I211210,I211465,);
not I_12290 (I211473,I211465);
not I_12291 (I211490,I211448);
nand I_12292 (I211187,I211490,I211309);
nand I_12293 (I211521,I282558,I282567);
and I_12294 (I211538,I211521,I282576);
DFFARX1 I_12295 (I211538,I2507,I211210,I211564,);
nor I_12296 (I211572,I211564,I211236);
DFFARX1 I_12297 (I211572,I2507,I211210,I211175,);
DFFARX1 I_12298 (I211564,I2507,I211210,I211193,);
nor I_12299 (I211617,I282564,I282567);
not I_12300 (I211634,I211617);
nor I_12301 (I211196,I211473,I211634);
nand I_12302 (I211181,I211490,I211634);
nor I_12303 (I211190,I211236,I211617);
DFFARX1 I_12304 (I211617,I2507,I211210,I211199,);
not I_12305 (I211737,I2514);
DFFARX1 I_12306 (I545279,I2507,I211737,I211763,);
nand I_12307 (I211771,I545276,I545279);
and I_12308 (I211788,I211771,I545288);
DFFARX1 I_12309 (I211788,I2507,I211737,I211814,);
nor I_12310 (I211705,I211814,I211763);
not I_12311 (I211836,I211814);
DFFARX1 I_12312 (I545276,I2507,I211737,I211862,);
nand I_12313 (I211870,I211862,I545294);
not I_12314 (I211887,I211870);
DFFARX1 I_12315 (I211887,I2507,I211737,I211913,);
not I_12316 (I211729,I211913);
nor I_12317 (I211935,I211763,I211870);
nor I_12318 (I211711,I211814,I211935);
DFFARX1 I_12319 (I545282,I2507,I211737,I211975,);
DFFARX1 I_12320 (I211975,I2507,I211737,I211992,);
not I_12321 (I212000,I211992);
not I_12322 (I212017,I211975);
nand I_12323 (I211714,I212017,I211836);
nand I_12324 (I212048,I545291,I545297);
and I_12325 (I212065,I212048,I545282);
DFFARX1 I_12326 (I212065,I2507,I211737,I212091,);
nor I_12327 (I212099,I212091,I211763);
DFFARX1 I_12328 (I212099,I2507,I211737,I211702,);
DFFARX1 I_12329 (I212091,I2507,I211737,I211720,);
nor I_12330 (I212144,I545285,I545297);
not I_12331 (I212161,I212144);
nor I_12332 (I211723,I212000,I212161);
nand I_12333 (I211708,I212017,I212161);
nor I_12334 (I211717,I211763,I212144);
DFFARX1 I_12335 (I212144,I2507,I211737,I211726,);
not I_12336 (I212264,I2514);
DFFARX1 I_12337 (I291486,I2507,I212264,I212290,);
nand I_12338 (I212298,I291486,I291498);
and I_12339 (I212315,I212298,I291483);
DFFARX1 I_12340 (I212315,I2507,I212264,I212341,);
nor I_12341 (I212232,I212341,I212290);
not I_12342 (I212363,I212341);
DFFARX1 I_12343 (I291507,I2507,I212264,I212389,);
nand I_12344 (I212397,I212389,I291504);
not I_12345 (I212414,I212397);
DFFARX1 I_12346 (I212414,I2507,I212264,I212440,);
not I_12347 (I212256,I212440);
nor I_12348 (I212462,I212290,I212397);
nor I_12349 (I212238,I212341,I212462);
DFFARX1 I_12350 (I291495,I2507,I212264,I212502,);
DFFARX1 I_12351 (I212502,I2507,I212264,I212519,);
not I_12352 (I212527,I212519);
not I_12353 (I212544,I212502);
nand I_12354 (I212241,I212544,I212363);
nand I_12355 (I212575,I291483,I291492);
and I_12356 (I212592,I212575,I291501);
DFFARX1 I_12357 (I212592,I2507,I212264,I212618,);
nor I_12358 (I212626,I212618,I212290);
DFFARX1 I_12359 (I212626,I2507,I212264,I212229,);
DFFARX1 I_12360 (I212618,I2507,I212264,I212247,);
nor I_12361 (I212671,I291489,I291492);
not I_12362 (I212688,I212671);
nor I_12363 (I212250,I212527,I212688);
nand I_12364 (I212235,I212544,I212688);
nor I_12365 (I212244,I212290,I212671);
DFFARX1 I_12366 (I212671,I2507,I212264,I212253,);
not I_12367 (I212791,I2514);
DFFARX1 I_12368 (I346677,I2507,I212791,I212817,);
nand I_12369 (I212825,I346668,I346683);
and I_12370 (I212842,I212825,I346689);
DFFARX1 I_12371 (I212842,I2507,I212791,I212868,);
nor I_12372 (I212759,I212868,I212817);
not I_12373 (I212890,I212868);
DFFARX1 I_12374 (I346674,I2507,I212791,I212916,);
nand I_12375 (I212924,I212916,I346668);
not I_12376 (I212941,I212924);
DFFARX1 I_12377 (I212941,I2507,I212791,I212967,);
not I_12378 (I212783,I212967);
nor I_12379 (I212989,I212817,I212924);
nor I_12380 (I212765,I212868,I212989);
DFFARX1 I_12381 (I346671,I2507,I212791,I213029,);
DFFARX1 I_12382 (I213029,I2507,I212791,I213046,);
not I_12383 (I213054,I213046);
not I_12384 (I213071,I213029);
nand I_12385 (I212768,I213071,I212890);
nand I_12386 (I213102,I346665,I346680);
and I_12387 (I213119,I213102,I346665);
DFFARX1 I_12388 (I213119,I2507,I212791,I213145,);
nor I_12389 (I213153,I213145,I212817);
DFFARX1 I_12390 (I213153,I2507,I212791,I212756,);
DFFARX1 I_12391 (I213145,I2507,I212791,I212774,);
nor I_12392 (I213198,I346686,I346680);
not I_12393 (I213215,I213198);
nor I_12394 (I212777,I213054,I213215);
nand I_12395 (I212762,I213071,I213215);
nor I_12396 (I212771,I212817,I213198);
DFFARX1 I_12397 (I213198,I2507,I212791,I212780,);
not I_12398 (I213318,I2514);
DFFARX1 I_12399 (I338588,I2507,I213318,I213344,);
nand I_12400 (I213352,I338573,I338576);
and I_12401 (I213369,I213352,I338591);
DFFARX1 I_12402 (I213369,I2507,I213318,I213395,);
nor I_12403 (I213286,I213395,I213344);
not I_12404 (I213417,I213395);
DFFARX1 I_12405 (I338585,I2507,I213318,I213443,);
nand I_12406 (I213451,I213443,I338576);
not I_12407 (I213468,I213451);
DFFARX1 I_12408 (I213468,I2507,I213318,I213494,);
not I_12409 (I213310,I213494);
nor I_12410 (I213516,I213344,I213451);
nor I_12411 (I213292,I213395,I213516);
DFFARX1 I_12412 (I338582,I2507,I213318,I213556,);
DFFARX1 I_12413 (I213556,I2507,I213318,I213573,);
not I_12414 (I213581,I213573);
not I_12415 (I213598,I213556);
nand I_12416 (I213295,I213598,I213417);
nand I_12417 (I213629,I338597,I338573);
and I_12418 (I213646,I213629,I338594);
DFFARX1 I_12419 (I213646,I2507,I213318,I213672,);
nor I_12420 (I213680,I213672,I213344);
DFFARX1 I_12421 (I213680,I2507,I213318,I213283,);
DFFARX1 I_12422 (I213672,I2507,I213318,I213301,);
nor I_12423 (I213725,I338579,I338573);
not I_12424 (I213742,I213725);
nor I_12425 (I213304,I213581,I213742);
nand I_12426 (I213289,I213598,I213742);
nor I_12427 (I213298,I213344,I213725);
DFFARX1 I_12428 (I213725,I2507,I213318,I213307,);
not I_12429 (I213845,I2514);
DFFARX1 I_12430 (I294461,I2507,I213845,I213871,);
nand I_12431 (I213879,I294461,I294473);
and I_12432 (I213896,I213879,I294458);
DFFARX1 I_12433 (I213896,I2507,I213845,I213922,);
nor I_12434 (I213813,I213922,I213871);
not I_12435 (I213944,I213922);
DFFARX1 I_12436 (I294482,I2507,I213845,I213970,);
nand I_12437 (I213978,I213970,I294479);
not I_12438 (I213995,I213978);
DFFARX1 I_12439 (I213995,I2507,I213845,I214021,);
not I_12440 (I213837,I214021);
nor I_12441 (I214043,I213871,I213978);
nor I_12442 (I213819,I213922,I214043);
DFFARX1 I_12443 (I294470,I2507,I213845,I214083,);
DFFARX1 I_12444 (I214083,I2507,I213845,I214100,);
not I_12445 (I214108,I214100);
not I_12446 (I214125,I214083);
nand I_12447 (I213822,I214125,I213944);
nand I_12448 (I214156,I294458,I294467);
and I_12449 (I214173,I214156,I294476);
DFFARX1 I_12450 (I214173,I2507,I213845,I214199,);
nor I_12451 (I214207,I214199,I213871);
DFFARX1 I_12452 (I214207,I2507,I213845,I213810,);
DFFARX1 I_12453 (I214199,I2507,I213845,I213828,);
nor I_12454 (I214252,I294464,I294467);
not I_12455 (I214269,I214252);
nor I_12456 (I213831,I214108,I214269);
nand I_12457 (I213816,I214125,I214269);
nor I_12458 (I213825,I213871,I214252);
DFFARX1 I_12459 (I214252,I2507,I213845,I213834,);
not I_12460 (I214372,I2514);
DFFARX1 I_12461 (I333964,I2507,I214372,I214398,);
nand I_12462 (I214406,I333949,I333952);
and I_12463 (I214423,I214406,I333967);
DFFARX1 I_12464 (I214423,I2507,I214372,I214449,);
nor I_12465 (I214340,I214449,I214398);
not I_12466 (I214471,I214449);
DFFARX1 I_12467 (I333961,I2507,I214372,I214497,);
nand I_12468 (I214505,I214497,I333952);
not I_12469 (I214522,I214505);
DFFARX1 I_12470 (I214522,I2507,I214372,I214548,);
not I_12471 (I214364,I214548);
nor I_12472 (I214570,I214398,I214505);
nor I_12473 (I214346,I214449,I214570);
DFFARX1 I_12474 (I333958,I2507,I214372,I214610,);
DFFARX1 I_12475 (I214610,I2507,I214372,I214627,);
not I_12476 (I214635,I214627);
not I_12477 (I214652,I214610);
nand I_12478 (I214349,I214652,I214471);
nand I_12479 (I214683,I333973,I333949);
and I_12480 (I214700,I214683,I333970);
DFFARX1 I_12481 (I214700,I2507,I214372,I214726,);
nor I_12482 (I214734,I214726,I214398);
DFFARX1 I_12483 (I214734,I2507,I214372,I214337,);
DFFARX1 I_12484 (I214726,I2507,I214372,I214355,);
nor I_12485 (I214779,I333955,I333949);
not I_12486 (I214796,I214779);
nor I_12487 (I214358,I214635,I214796);
nand I_12488 (I214343,I214652,I214796);
nor I_12489 (I214352,I214398,I214779);
DFFARX1 I_12490 (I214779,I2507,I214372,I214361,);
not I_12491 (I214899,I2514);
DFFARX1 I_12492 (I1396,I2507,I214899,I214925,);
nand I_12493 (I214933,I2484,I1836);
and I_12494 (I214950,I214933,I1532);
DFFARX1 I_12495 (I214950,I2507,I214899,I214976,);
nor I_12496 (I214867,I214976,I214925);
not I_12497 (I214998,I214976);
DFFARX1 I_12498 (I2068,I2507,I214899,I215024,);
nand I_12499 (I215032,I215024,I1468);
not I_12500 (I215049,I215032);
DFFARX1 I_12501 (I215049,I2507,I214899,I215075,);
not I_12502 (I214891,I215075);
nor I_12503 (I215097,I214925,I215032);
nor I_12504 (I214873,I214976,I215097);
DFFARX1 I_12505 (I2156,I2507,I214899,I215137,);
DFFARX1 I_12506 (I215137,I2507,I214899,I215154,);
not I_12507 (I215162,I215154);
not I_12508 (I215179,I215137);
nand I_12509 (I214876,I215179,I214998);
nand I_12510 (I215210,I2076,I2420);
and I_12511 (I215227,I215210,I2300);
DFFARX1 I_12512 (I215227,I2507,I214899,I215253,);
nor I_12513 (I215261,I215253,I214925);
DFFARX1 I_12514 (I215261,I2507,I214899,I214864,);
DFFARX1 I_12515 (I215253,I2507,I214899,I214882,);
nor I_12516 (I215306,I2316,I2420);
not I_12517 (I215323,I215306);
nor I_12518 (I214885,I215162,I215323);
nand I_12519 (I214870,I215179,I215323);
nor I_12520 (I214879,I214925,I215306);
DFFARX1 I_12521 (I215306,I2507,I214899,I214888,);
not I_12522 (I215426,I2514);
DFFARX1 I_12523 (I35670,I2507,I215426,I215452,);
nand I_12524 (I215460,I35682,I35691);
and I_12525 (I215477,I215460,I35670);
DFFARX1 I_12526 (I215477,I2507,I215426,I215503,);
nor I_12527 (I215394,I215503,I215452);
not I_12528 (I215525,I215503);
DFFARX1 I_12529 (I35685,I2507,I215426,I215551,);
nand I_12530 (I215559,I215551,I35673);
not I_12531 (I215576,I215559);
DFFARX1 I_12532 (I215576,I2507,I215426,I215602,);
not I_12533 (I215418,I215602);
nor I_12534 (I215624,I215452,I215559);
nor I_12535 (I215400,I215503,I215624);
DFFARX1 I_12536 (I35676,I2507,I215426,I215664,);
DFFARX1 I_12537 (I215664,I2507,I215426,I215681,);
not I_12538 (I215689,I215681);
not I_12539 (I215706,I215664);
nand I_12540 (I215403,I215706,I215525);
nand I_12541 (I215737,I35667,I35667);
and I_12542 (I215754,I215737,I35679);
DFFARX1 I_12543 (I215754,I2507,I215426,I215780,);
nor I_12544 (I215788,I215780,I215452);
DFFARX1 I_12545 (I215788,I2507,I215426,I215391,);
DFFARX1 I_12546 (I215780,I2507,I215426,I215409,);
nor I_12547 (I215833,I35688,I35667);
not I_12548 (I215850,I215833);
nor I_12549 (I215412,I215689,I215850);
nand I_12550 (I215397,I215706,I215850);
nor I_12551 (I215406,I215452,I215833);
DFFARX1 I_12552 (I215833,I2507,I215426,I215415,);
not I_12553 (I215953,I2514);
DFFARX1 I_12554 (I464478,I2507,I215953,I215979,);
nand I_12555 (I215987,I464481,I464475);
and I_12556 (I216004,I215987,I464487);
DFFARX1 I_12557 (I216004,I2507,I215953,I216030,);
nor I_12558 (I215921,I216030,I215979);
not I_12559 (I216052,I216030);
DFFARX1 I_12560 (I464490,I2507,I215953,I216078,);
nand I_12561 (I216086,I216078,I464481);
not I_12562 (I216103,I216086);
DFFARX1 I_12563 (I216103,I2507,I215953,I216129,);
not I_12564 (I215945,I216129);
nor I_12565 (I216151,I215979,I216086);
nor I_12566 (I215927,I216030,I216151);
DFFARX1 I_12567 (I464493,I2507,I215953,I216191,);
DFFARX1 I_12568 (I216191,I2507,I215953,I216208,);
not I_12569 (I216216,I216208);
not I_12570 (I216233,I216191);
nand I_12571 (I215930,I216233,I216052);
nand I_12572 (I216264,I464475,I464484);
and I_12573 (I216281,I216264,I464478);
DFFARX1 I_12574 (I216281,I2507,I215953,I216307,);
nor I_12575 (I216315,I216307,I215979);
DFFARX1 I_12576 (I216315,I2507,I215953,I215918,);
DFFARX1 I_12577 (I216307,I2507,I215953,I215936,);
nor I_12578 (I216360,I464496,I464484);
not I_12579 (I216377,I216360);
nor I_12580 (I215939,I216216,I216377);
nand I_12581 (I215924,I216233,I216377);
nor I_12582 (I215933,I215979,I216360);
DFFARX1 I_12583 (I216360,I2507,I215953,I215942,);
not I_12584 (I216480,I2514);
DFFARX1 I_12585 (I44629,I2507,I216480,I216506,);
nand I_12586 (I216514,I44641,I44650);
and I_12587 (I216531,I216514,I44629);
DFFARX1 I_12588 (I216531,I2507,I216480,I216557,);
nor I_12589 (I216448,I216557,I216506);
not I_12590 (I216579,I216557);
DFFARX1 I_12591 (I44644,I2507,I216480,I216605,);
nand I_12592 (I216613,I216605,I44632);
not I_12593 (I216630,I216613);
DFFARX1 I_12594 (I216630,I2507,I216480,I216656,);
not I_12595 (I216472,I216656);
nor I_12596 (I216678,I216506,I216613);
nor I_12597 (I216454,I216557,I216678);
DFFARX1 I_12598 (I44635,I2507,I216480,I216718,);
DFFARX1 I_12599 (I216718,I2507,I216480,I216735,);
not I_12600 (I216743,I216735);
not I_12601 (I216760,I216718);
nand I_12602 (I216457,I216760,I216579);
nand I_12603 (I216791,I44626,I44626);
and I_12604 (I216808,I216791,I44638);
DFFARX1 I_12605 (I216808,I2507,I216480,I216834,);
nor I_12606 (I216842,I216834,I216506);
DFFARX1 I_12607 (I216842,I2507,I216480,I216445,);
DFFARX1 I_12608 (I216834,I2507,I216480,I216463,);
nor I_12609 (I216887,I44647,I44626);
not I_12610 (I216904,I216887);
nor I_12611 (I216466,I216743,I216904);
nand I_12612 (I216451,I216760,I216904);
nor I_12613 (I216460,I216506,I216887);
DFFARX1 I_12614 (I216887,I2507,I216480,I216469,);
not I_12615 (I217007,I2514);
DFFARX1 I_12616 (I700184,I2507,I217007,I217033,);
nand I_12617 (I217041,I700163,I700163);
and I_12618 (I217058,I217041,I700190);
DFFARX1 I_12619 (I217058,I2507,I217007,I217084,);
nor I_12620 (I216975,I217084,I217033);
not I_12621 (I217106,I217084);
DFFARX1 I_12622 (I700178,I2507,I217007,I217132,);
nand I_12623 (I217140,I217132,I700181);
not I_12624 (I217157,I217140);
DFFARX1 I_12625 (I217157,I2507,I217007,I217183,);
not I_12626 (I216999,I217183);
nor I_12627 (I217205,I217033,I217140);
nor I_12628 (I216981,I217084,I217205);
DFFARX1 I_12629 (I700172,I2507,I217007,I217245,);
DFFARX1 I_12630 (I217245,I2507,I217007,I217262,);
not I_12631 (I217270,I217262);
not I_12632 (I217287,I217245);
nand I_12633 (I216984,I217287,I217106);
nand I_12634 (I217318,I700169,I700166);
and I_12635 (I217335,I217318,I700187);
DFFARX1 I_12636 (I217335,I2507,I217007,I217361,);
nor I_12637 (I217369,I217361,I217033);
DFFARX1 I_12638 (I217369,I2507,I217007,I216972,);
DFFARX1 I_12639 (I217361,I2507,I217007,I216990,);
nor I_12640 (I217414,I700175,I700166);
not I_12641 (I217431,I217414);
nor I_12642 (I216993,I217270,I217431);
nand I_12643 (I216978,I217287,I217431);
nor I_12644 (I216987,I217033,I217414);
DFFARX1 I_12645 (I217414,I2507,I217007,I216996,);
not I_12646 (I217534,I2514);
DFFARX1 I_12647 (I1932,I2507,I217534,I217560,);
nand I_12648 (I217568,I1700,I1612);
and I_12649 (I217585,I217568,I2052);
DFFARX1 I_12650 (I217585,I2507,I217534,I217611,);
nor I_12651 (I217502,I217611,I217560);
not I_12652 (I217633,I217611);
DFFARX1 I_12653 (I1740,I2507,I217534,I217659,);
nand I_12654 (I217667,I217659,I1980);
not I_12655 (I217684,I217667);
DFFARX1 I_12656 (I217684,I2507,I217534,I217710,);
not I_12657 (I217526,I217710);
nor I_12658 (I217732,I217560,I217667);
nor I_12659 (I217508,I217611,I217732);
DFFARX1 I_12660 (I2196,I2507,I217534,I217772,);
DFFARX1 I_12661 (I217772,I2507,I217534,I217789,);
not I_12662 (I217797,I217789);
not I_12663 (I217814,I217772);
nand I_12664 (I217511,I217814,I217633);
nand I_12665 (I217845,I2340,I1508);
and I_12666 (I217862,I217845,I1404);
DFFARX1 I_12667 (I217862,I2507,I217534,I217888,);
nor I_12668 (I217896,I217888,I217560);
DFFARX1 I_12669 (I217896,I2507,I217534,I217499,);
DFFARX1 I_12670 (I217888,I2507,I217534,I217517,);
nor I_12671 (I217941,I1972,I1508);
not I_12672 (I217958,I217941);
nor I_12673 (I217520,I217797,I217958);
nand I_12674 (I217505,I217814,I217958);
nor I_12675 (I217514,I217560,I217941);
DFFARX1 I_12676 (I217941,I2507,I217534,I217523,);
not I_12677 (I218061,I2514);
DFFARX1 I_12678 (I13006,I2507,I218061,I218087,);
nand I_12679 (I218095,I13030,I13009);
and I_12680 (I218112,I218095,I13006);
DFFARX1 I_12681 (I218112,I2507,I218061,I218138,);
nor I_12682 (I218029,I218138,I218087);
not I_12683 (I218160,I218138);
DFFARX1 I_12684 (I13012,I2507,I218061,I218186,);
nand I_12685 (I218194,I218186,I13021);
not I_12686 (I218211,I218194);
DFFARX1 I_12687 (I218211,I2507,I218061,I218237,);
not I_12688 (I218053,I218237);
nor I_12689 (I218259,I218087,I218194);
nor I_12690 (I218035,I218138,I218259);
DFFARX1 I_12691 (I13015,I2507,I218061,I218299,);
DFFARX1 I_12692 (I218299,I2507,I218061,I218316,);
not I_12693 (I218324,I218316);
not I_12694 (I218341,I218299);
nand I_12695 (I218038,I218341,I218160);
nand I_12696 (I218372,I13027,I13009);
and I_12697 (I218389,I218372,I13018);
DFFARX1 I_12698 (I218389,I2507,I218061,I218415,);
nor I_12699 (I218423,I218415,I218087);
DFFARX1 I_12700 (I218423,I2507,I218061,I218026,);
DFFARX1 I_12701 (I218415,I2507,I218061,I218044,);
nor I_12702 (I218468,I13024,I13009);
not I_12703 (I218485,I218468);
nor I_12704 (I218047,I218324,I218485);
nand I_12705 (I218032,I218341,I218485);
nor I_12706 (I218041,I218087,I218468);
DFFARX1 I_12707 (I218468,I2507,I218061,I218050,);
not I_12708 (I218588,I2514);
DFFARX1 I_12709 (I709109,I2507,I218588,I218614,);
nand I_12710 (I218622,I709088,I709088);
and I_12711 (I218639,I218622,I709115);
DFFARX1 I_12712 (I218639,I2507,I218588,I218665,);
nor I_12713 (I218556,I218665,I218614);
not I_12714 (I218687,I218665);
DFFARX1 I_12715 (I709103,I2507,I218588,I218713,);
nand I_12716 (I218721,I218713,I709106);
not I_12717 (I218738,I218721);
DFFARX1 I_12718 (I218738,I2507,I218588,I218764,);
not I_12719 (I218580,I218764);
nor I_12720 (I218786,I218614,I218721);
nor I_12721 (I218562,I218665,I218786);
DFFARX1 I_12722 (I709097,I2507,I218588,I218826,);
DFFARX1 I_12723 (I218826,I2507,I218588,I218843,);
not I_12724 (I218851,I218843);
not I_12725 (I218868,I218826);
nand I_12726 (I218565,I218868,I218687);
nand I_12727 (I218899,I709094,I709091);
and I_12728 (I218916,I218899,I709112);
DFFARX1 I_12729 (I218916,I2507,I218588,I218942,);
nor I_12730 (I218950,I218942,I218614);
DFFARX1 I_12731 (I218950,I2507,I218588,I218553,);
DFFARX1 I_12732 (I218942,I2507,I218588,I218571,);
nor I_12733 (I218995,I709100,I709091);
not I_12734 (I219012,I218995);
nor I_12735 (I218574,I218851,I219012);
nand I_12736 (I218559,I218868,I219012);
nor I_12737 (I218568,I218614,I218995);
DFFARX1 I_12738 (I218995,I2507,I218588,I218577,);
not I_12739 (I219115,I2514);
DFFARX1 I_12740 (I380201,I2507,I219115,I219141,);
nand I_12741 (I219149,I380192,I380207);
and I_12742 (I219166,I219149,I380213);
DFFARX1 I_12743 (I219166,I2507,I219115,I219192,);
nor I_12744 (I219083,I219192,I219141);
not I_12745 (I219214,I219192);
DFFARX1 I_12746 (I380198,I2507,I219115,I219240,);
nand I_12747 (I219248,I219240,I380192);
not I_12748 (I219265,I219248);
DFFARX1 I_12749 (I219265,I2507,I219115,I219291,);
not I_12750 (I219107,I219291);
nor I_12751 (I219313,I219141,I219248);
nor I_12752 (I219089,I219192,I219313);
DFFARX1 I_12753 (I380195,I2507,I219115,I219353,);
DFFARX1 I_12754 (I219353,I2507,I219115,I219370,);
not I_12755 (I219378,I219370);
not I_12756 (I219395,I219353);
nand I_12757 (I219092,I219395,I219214);
nand I_12758 (I219426,I380189,I380204);
and I_12759 (I219443,I219426,I380189);
DFFARX1 I_12760 (I219443,I2507,I219115,I219469,);
nor I_12761 (I219477,I219469,I219141);
DFFARX1 I_12762 (I219477,I2507,I219115,I219080,);
DFFARX1 I_12763 (I219469,I2507,I219115,I219098,);
nor I_12764 (I219522,I380210,I380204);
not I_12765 (I219539,I219522);
nor I_12766 (I219101,I219378,I219539);
nand I_12767 (I219086,I219395,I219539);
nor I_12768 (I219095,I219141,I219522);
DFFARX1 I_12769 (I219522,I2507,I219115,I219104,);
not I_12770 (I219642,I2514);
DFFARX1 I_12771 (I643639,I2507,I219642,I219668,);
nand I_12772 (I219676,I643621,I643645);
and I_12773 (I219693,I219676,I643636);
DFFARX1 I_12774 (I219693,I2507,I219642,I219719,);
nor I_12775 (I219610,I219719,I219668);
not I_12776 (I219741,I219719);
DFFARX1 I_12777 (I643642,I2507,I219642,I219767,);
nand I_12778 (I219775,I219767,I643630);
not I_12779 (I219792,I219775);
DFFARX1 I_12780 (I219792,I2507,I219642,I219818,);
not I_12781 (I219634,I219818);
nor I_12782 (I219840,I219668,I219775);
nor I_12783 (I219616,I219719,I219840);
DFFARX1 I_12784 (I643621,I2507,I219642,I219880,);
DFFARX1 I_12785 (I219880,I2507,I219642,I219897,);
not I_12786 (I219905,I219897);
not I_12787 (I219922,I219880);
nand I_12788 (I219619,I219922,I219741);
nand I_12789 (I219953,I643627,I643624);
and I_12790 (I219970,I219953,I643633);
DFFARX1 I_12791 (I219970,I2507,I219642,I219996,);
nor I_12792 (I220004,I219996,I219668);
DFFARX1 I_12793 (I220004,I2507,I219642,I219607,);
DFFARX1 I_12794 (I219996,I2507,I219642,I219625,);
nor I_12795 (I220049,I643624,I643624);
not I_12796 (I220066,I220049);
nor I_12797 (I219628,I219905,I220066);
nand I_12798 (I219613,I219922,I220066);
nor I_12799 (I219622,I219668,I220049);
DFFARX1 I_12800 (I220049,I2507,I219642,I219631,);
not I_12801 (I220169,I2514);
DFFARX1 I_12802 (I667674,I2507,I220169,I220195,);
nand I_12803 (I220203,I667671,I667662);
and I_12804 (I220220,I220203,I667659);
DFFARX1 I_12805 (I220220,I2507,I220169,I220246,);
nor I_12806 (I220137,I220246,I220195);
not I_12807 (I220268,I220246);
DFFARX1 I_12808 (I667668,I2507,I220169,I220294,);
nand I_12809 (I220302,I220294,I667677);
not I_12810 (I220319,I220302);
DFFARX1 I_12811 (I220319,I2507,I220169,I220345,);
not I_12812 (I220161,I220345);
nor I_12813 (I220367,I220195,I220302);
nor I_12814 (I220143,I220246,I220367);
DFFARX1 I_12815 (I667680,I2507,I220169,I220407,);
DFFARX1 I_12816 (I220407,I2507,I220169,I220424,);
not I_12817 (I220432,I220424);
not I_12818 (I220449,I220407);
nand I_12819 (I220146,I220449,I220268);
nand I_12820 (I220480,I667659,I667665);
and I_12821 (I220497,I220480,I667683);
DFFARX1 I_12822 (I220497,I2507,I220169,I220523,);
nor I_12823 (I220531,I220523,I220195);
DFFARX1 I_12824 (I220531,I2507,I220169,I220134,);
DFFARX1 I_12825 (I220523,I2507,I220169,I220152,);
nor I_12826 (I220576,I667662,I667665);
not I_12827 (I220593,I220576);
nor I_12828 (I220155,I220432,I220593);
nand I_12829 (I220140,I220449,I220593);
nor I_12830 (I220149,I220195,I220576);
DFFARX1 I_12831 (I220576,I2507,I220169,I220158,);
not I_12832 (I220696,I2514);
DFFARX1 I_12833 (I237860,I2507,I220696,I220722,);
nand I_12834 (I220730,I237872,I237851);
and I_12835 (I220747,I220730,I237875);
DFFARX1 I_12836 (I220747,I2507,I220696,I220773,);
nor I_12837 (I220664,I220773,I220722);
not I_12838 (I220795,I220773);
DFFARX1 I_12839 (I237866,I2507,I220696,I220821,);
nand I_12840 (I220829,I220821,I237848);
not I_12841 (I220846,I220829);
DFFARX1 I_12842 (I220846,I2507,I220696,I220872,);
not I_12843 (I220688,I220872);
nor I_12844 (I220894,I220722,I220829);
nor I_12845 (I220670,I220773,I220894);
DFFARX1 I_12846 (I237863,I2507,I220696,I220934,);
DFFARX1 I_12847 (I220934,I2507,I220696,I220951,);
not I_12848 (I220959,I220951);
not I_12849 (I220976,I220934);
nand I_12850 (I220673,I220976,I220795);
nand I_12851 (I221007,I237848,I237854);
and I_12852 (I221024,I221007,I237857);
DFFARX1 I_12853 (I221024,I2507,I220696,I221050,);
nor I_12854 (I221058,I221050,I220722);
DFFARX1 I_12855 (I221058,I2507,I220696,I220661,);
DFFARX1 I_12856 (I221050,I2507,I220696,I220679,);
nor I_12857 (I221103,I237869,I237854);
not I_12858 (I221120,I221103);
nor I_12859 (I220682,I220959,I221120);
nand I_12860 (I220667,I220976,I221120);
nor I_12861 (I220676,I220722,I221103);
DFFARX1 I_12862 (I221103,I2507,I220696,I220685,);
not I_12863 (I221223,I2514);
DFFARX1 I_12864 (I138959,I2507,I221223,I221249,);
nand I_12865 (I221257,I138959,I138965);
and I_12866 (I221274,I221257,I138983);
DFFARX1 I_12867 (I221274,I2507,I221223,I221300,);
nor I_12868 (I221191,I221300,I221249);
not I_12869 (I221322,I221300);
DFFARX1 I_12870 (I138971,I2507,I221223,I221348,);
nand I_12871 (I221356,I221348,I138968);
not I_12872 (I221373,I221356);
DFFARX1 I_12873 (I221373,I2507,I221223,I221399,);
not I_12874 (I221215,I221399);
nor I_12875 (I221421,I221249,I221356);
nor I_12876 (I221197,I221300,I221421);
DFFARX1 I_12877 (I138977,I2507,I221223,I221461,);
DFFARX1 I_12878 (I221461,I2507,I221223,I221478,);
not I_12879 (I221486,I221478);
not I_12880 (I221503,I221461);
nand I_12881 (I221200,I221503,I221322);
nand I_12882 (I221534,I138962,I138962);
and I_12883 (I221551,I221534,I138974);
DFFARX1 I_12884 (I221551,I2507,I221223,I221577,);
nor I_12885 (I221585,I221577,I221249);
DFFARX1 I_12886 (I221585,I2507,I221223,I221188,);
DFFARX1 I_12887 (I221577,I2507,I221223,I221206,);
nor I_12888 (I221630,I138980,I138962);
not I_12889 (I221647,I221630);
nor I_12890 (I221209,I221486,I221647);
nand I_12891 (I221194,I221503,I221647);
nor I_12892 (I221203,I221249,I221630);
DFFARX1 I_12893 (I221630,I2507,I221223,I221212,);
not I_12894 (I221750,I2514);
DFFARX1 I_12895 (I266692,I2507,I221750,I221776,);
nand I_12896 (I221784,I266704,I266683);
and I_12897 (I221801,I221784,I266707);
DFFARX1 I_12898 (I221801,I2507,I221750,I221827,);
nor I_12899 (I221718,I221827,I221776);
not I_12900 (I221849,I221827);
DFFARX1 I_12901 (I266698,I2507,I221750,I221875,);
nand I_12902 (I221883,I221875,I266680);
not I_12903 (I221900,I221883);
DFFARX1 I_12904 (I221900,I2507,I221750,I221926,);
not I_12905 (I221742,I221926);
nor I_12906 (I221948,I221776,I221883);
nor I_12907 (I221724,I221827,I221948);
DFFARX1 I_12908 (I266695,I2507,I221750,I221988,);
DFFARX1 I_12909 (I221988,I2507,I221750,I222005,);
not I_12910 (I222013,I222005);
not I_12911 (I222030,I221988);
nand I_12912 (I221727,I222030,I221849);
nand I_12913 (I222061,I266680,I266686);
and I_12914 (I222078,I222061,I266689);
DFFARX1 I_12915 (I222078,I2507,I221750,I222104,);
nor I_12916 (I222112,I222104,I221776);
DFFARX1 I_12917 (I222112,I2507,I221750,I221715,);
DFFARX1 I_12918 (I222104,I2507,I221750,I221733,);
nor I_12919 (I222157,I266701,I266686);
not I_12920 (I222174,I222157);
nor I_12921 (I221736,I222013,I222174);
nand I_12922 (I221721,I222030,I222174);
nor I_12923 (I221730,I221776,I222157);
DFFARX1 I_12924 (I222157,I2507,I221750,I221739,);
not I_12925 (I222277,I2514);
DFFARX1 I_12926 (I406789,I2507,I222277,I222303,);
nand I_12927 (I222311,I406780,I406795);
and I_12928 (I222328,I222311,I406801);
DFFARX1 I_12929 (I222328,I2507,I222277,I222354,);
nor I_12930 (I222245,I222354,I222303);
not I_12931 (I222376,I222354);
DFFARX1 I_12932 (I406786,I2507,I222277,I222402,);
nand I_12933 (I222410,I222402,I406780);
not I_12934 (I222427,I222410);
DFFARX1 I_12935 (I222427,I2507,I222277,I222453,);
not I_12936 (I222269,I222453);
nor I_12937 (I222475,I222303,I222410);
nor I_12938 (I222251,I222354,I222475);
DFFARX1 I_12939 (I406783,I2507,I222277,I222515,);
DFFARX1 I_12940 (I222515,I2507,I222277,I222532,);
not I_12941 (I222540,I222532);
not I_12942 (I222557,I222515);
nand I_12943 (I222254,I222557,I222376);
nand I_12944 (I222588,I406777,I406792);
and I_12945 (I222605,I222588,I406777);
DFFARX1 I_12946 (I222605,I2507,I222277,I222631,);
nor I_12947 (I222639,I222631,I222303);
DFFARX1 I_12948 (I222639,I2507,I222277,I222242,);
DFFARX1 I_12949 (I222631,I2507,I222277,I222260,);
nor I_12950 (I222684,I406798,I406792);
not I_12951 (I222701,I222684);
nor I_12952 (I222263,I222540,I222701);
nand I_12953 (I222248,I222557,I222701);
nor I_12954 (I222257,I222303,I222684);
DFFARX1 I_12955 (I222684,I2507,I222277,I222266,);
not I_12956 (I222804,I2514);
DFFARX1 I_12957 (I626587,I2507,I222804,I222830,);
nand I_12958 (I222838,I626602,I626587);
and I_12959 (I222855,I222838,I626605);
DFFARX1 I_12960 (I222855,I2507,I222804,I222881,);
nor I_12961 (I222772,I222881,I222830);
not I_12962 (I222903,I222881);
DFFARX1 I_12963 (I626611,I2507,I222804,I222929,);
nand I_12964 (I222937,I222929,I626593);
not I_12965 (I222954,I222937);
DFFARX1 I_12966 (I222954,I2507,I222804,I222980,);
not I_12967 (I222796,I222980);
nor I_12968 (I223002,I222830,I222937);
nor I_12969 (I222778,I222881,I223002);
DFFARX1 I_12970 (I626590,I2507,I222804,I223042,);
DFFARX1 I_12971 (I223042,I2507,I222804,I223059,);
not I_12972 (I223067,I223059);
not I_12973 (I223084,I223042);
nand I_12974 (I222781,I223084,I222903);
nand I_12975 (I223115,I626590,I626596);
and I_12976 (I223132,I223115,I626608);
DFFARX1 I_12977 (I223132,I2507,I222804,I223158,);
nor I_12978 (I223166,I223158,I222830);
DFFARX1 I_12979 (I223166,I2507,I222804,I222769,);
DFFARX1 I_12980 (I223158,I2507,I222804,I222787,);
nor I_12981 (I223211,I626599,I626596);
not I_12982 (I223228,I223211);
nor I_12983 (I222790,I223067,I223228);
nand I_12984 (I222775,I223084,I223228);
nor I_12985 (I222784,I222830,I223211);
DFFARX1 I_12986 (I223211,I2507,I222804,I222793,);
not I_12987 (I223331,I2514);
DFFARX1 I_12988 (I73614,I2507,I223331,I223357,);
nand I_12989 (I223365,I73626,I73635);
and I_12990 (I223382,I223365,I73614);
DFFARX1 I_12991 (I223382,I2507,I223331,I223408,);
nor I_12992 (I223299,I223408,I223357);
not I_12993 (I223430,I223408);
DFFARX1 I_12994 (I73629,I2507,I223331,I223456,);
nand I_12995 (I223464,I223456,I73617);
not I_12996 (I223481,I223464);
DFFARX1 I_12997 (I223481,I2507,I223331,I223507,);
not I_12998 (I223323,I223507);
nor I_12999 (I223529,I223357,I223464);
nor I_13000 (I223305,I223408,I223529);
DFFARX1 I_13001 (I73620,I2507,I223331,I223569,);
DFFARX1 I_13002 (I223569,I2507,I223331,I223586,);
not I_13003 (I223594,I223586);
not I_13004 (I223611,I223569);
nand I_13005 (I223308,I223611,I223430);
nand I_13006 (I223642,I73611,I73611);
and I_13007 (I223659,I223642,I73623);
DFFARX1 I_13008 (I223659,I2507,I223331,I223685,);
nor I_13009 (I223693,I223685,I223357);
DFFARX1 I_13010 (I223693,I2507,I223331,I223296,);
DFFARX1 I_13011 (I223685,I2507,I223331,I223314,);
nor I_13012 (I223738,I73632,I73611);
not I_13013 (I223755,I223738);
nor I_13014 (I223317,I223594,I223755);
nand I_13015 (I223302,I223611,I223755);
nor I_13016 (I223311,I223357,I223738);
DFFARX1 I_13017 (I223738,I2507,I223331,I223320,);
not I_13018 (I223858,I2514);
DFFARX1 I_13019 (I76249,I2507,I223858,I223884,);
nand I_13020 (I223892,I76261,I76270);
and I_13021 (I223909,I223892,I76249);
DFFARX1 I_13022 (I223909,I2507,I223858,I223935,);
nor I_13023 (I223826,I223935,I223884);
not I_13024 (I223957,I223935);
DFFARX1 I_13025 (I76264,I2507,I223858,I223983,);
nand I_13026 (I223991,I223983,I76252);
not I_13027 (I224008,I223991);
DFFARX1 I_13028 (I224008,I2507,I223858,I224034,);
not I_13029 (I223850,I224034);
nor I_13030 (I224056,I223884,I223991);
nor I_13031 (I223832,I223935,I224056);
DFFARX1 I_13032 (I76255,I2507,I223858,I224096,);
DFFARX1 I_13033 (I224096,I2507,I223858,I224113,);
not I_13034 (I224121,I224113);
not I_13035 (I224138,I224096);
nand I_13036 (I223835,I224138,I223957);
nand I_13037 (I224169,I76246,I76246);
and I_13038 (I224186,I224169,I76258);
DFFARX1 I_13039 (I224186,I2507,I223858,I224212,);
nor I_13040 (I224220,I224212,I223884);
DFFARX1 I_13041 (I224220,I2507,I223858,I223823,);
DFFARX1 I_13042 (I224212,I2507,I223858,I223841,);
nor I_13043 (I224265,I76267,I76246);
not I_13044 (I224282,I224265);
nor I_13045 (I223844,I224121,I224282);
nand I_13046 (I223829,I224138,I224282);
nor I_13047 (I223838,I223884,I224265);
DFFARX1 I_13048 (I224265,I2507,I223858,I223847,);
not I_13049 (I224385,I2514);
DFFARX1 I_13050 (I259620,I2507,I224385,I224411,);
nand I_13051 (I224419,I259632,I259611);
and I_13052 (I224436,I224419,I259635);
DFFARX1 I_13053 (I224436,I2507,I224385,I224462,);
nor I_13054 (I224353,I224462,I224411);
not I_13055 (I224484,I224462);
DFFARX1 I_13056 (I259626,I2507,I224385,I224510,);
nand I_13057 (I224518,I224510,I259608);
not I_13058 (I224535,I224518);
DFFARX1 I_13059 (I224535,I2507,I224385,I224561,);
not I_13060 (I224377,I224561);
nor I_13061 (I224583,I224411,I224518);
nor I_13062 (I224359,I224462,I224583);
DFFARX1 I_13063 (I259623,I2507,I224385,I224623,);
DFFARX1 I_13064 (I224623,I2507,I224385,I224640,);
not I_13065 (I224648,I224640);
not I_13066 (I224665,I224623);
nand I_13067 (I224362,I224665,I224484);
nand I_13068 (I224696,I259608,I259614);
and I_13069 (I224713,I224696,I259617);
DFFARX1 I_13070 (I224713,I2507,I224385,I224739,);
nor I_13071 (I224747,I224739,I224411);
DFFARX1 I_13072 (I224747,I2507,I224385,I224350,);
DFFARX1 I_13073 (I224739,I2507,I224385,I224368,);
nor I_13074 (I224792,I259629,I259614);
not I_13075 (I224809,I224792);
nor I_13076 (I224371,I224648,I224809);
nand I_13077 (I224356,I224665,I224809);
nor I_13078 (I224365,I224411,I224792);
DFFARX1 I_13079 (I224792,I2507,I224385,I224374,);
not I_13080 (I224912,I2514);
DFFARX1 I_13081 (I271588,I2507,I224912,I224938,);
nand I_13082 (I224946,I271600,I271579);
and I_13083 (I224963,I224946,I271603);
DFFARX1 I_13084 (I224963,I2507,I224912,I224989,);
nor I_13085 (I224880,I224989,I224938);
not I_13086 (I225011,I224989);
DFFARX1 I_13087 (I271594,I2507,I224912,I225037,);
nand I_13088 (I225045,I225037,I271576);
not I_13089 (I225062,I225045);
DFFARX1 I_13090 (I225062,I2507,I224912,I225088,);
not I_13091 (I224904,I225088);
nor I_13092 (I225110,I224938,I225045);
nor I_13093 (I224886,I224989,I225110);
DFFARX1 I_13094 (I271591,I2507,I224912,I225150,);
DFFARX1 I_13095 (I225150,I2507,I224912,I225167,);
not I_13096 (I225175,I225167);
not I_13097 (I225192,I225150);
nand I_13098 (I224889,I225192,I225011);
nand I_13099 (I225223,I271576,I271582);
and I_13100 (I225240,I225223,I271585);
DFFARX1 I_13101 (I225240,I2507,I224912,I225266,);
nor I_13102 (I225274,I225266,I224938);
DFFARX1 I_13103 (I225274,I2507,I224912,I224877,);
DFFARX1 I_13104 (I225266,I2507,I224912,I224895,);
nor I_13105 (I225319,I271597,I271582);
not I_13106 (I225336,I225319);
nor I_13107 (I224898,I225175,I225336);
nand I_13108 (I224883,I225192,I225336);
nor I_13109 (I224892,I224938,I225319);
DFFARX1 I_13110 (I225319,I2507,I224912,I224901,);
not I_13111 (I225439,I2514);
DFFARX1 I_13112 (I586127,I2507,I225439,I225465,);
nand I_13113 (I225473,I586142,I586127);
and I_13114 (I225490,I225473,I586145);
DFFARX1 I_13115 (I225490,I2507,I225439,I225516,);
nor I_13116 (I225407,I225516,I225465);
not I_13117 (I225538,I225516);
DFFARX1 I_13118 (I586151,I2507,I225439,I225564,);
nand I_13119 (I225572,I225564,I586133);
not I_13120 (I225589,I225572);
DFFARX1 I_13121 (I225589,I2507,I225439,I225615,);
not I_13122 (I225431,I225615);
nor I_13123 (I225637,I225465,I225572);
nor I_13124 (I225413,I225516,I225637);
DFFARX1 I_13125 (I586130,I2507,I225439,I225677,);
DFFARX1 I_13126 (I225677,I2507,I225439,I225694,);
not I_13127 (I225702,I225694);
not I_13128 (I225719,I225677);
nand I_13129 (I225416,I225719,I225538);
nand I_13130 (I225750,I586130,I586136);
and I_13131 (I225767,I225750,I586148);
DFFARX1 I_13132 (I225767,I2507,I225439,I225793,);
nor I_13133 (I225801,I225793,I225465);
DFFARX1 I_13134 (I225801,I2507,I225439,I225404,);
DFFARX1 I_13135 (I225793,I2507,I225439,I225422,);
nor I_13136 (I225846,I586139,I586136);
not I_13137 (I225863,I225846);
nor I_13138 (I225425,I225702,I225863);
nand I_13139 (I225410,I225719,I225863);
nor I_13140 (I225419,I225465,I225846);
DFFARX1 I_13141 (I225846,I2507,I225439,I225428,);
not I_13142 (I225966,I2514);
DFFARX1 I_13143 (I564914,I2507,I225966,I225992,);
nand I_13144 (I226000,I564911,I564914);
and I_13145 (I226017,I226000,I564923);
DFFARX1 I_13146 (I226017,I2507,I225966,I226043,);
nor I_13147 (I225934,I226043,I225992);
not I_13148 (I226065,I226043);
DFFARX1 I_13149 (I564911,I2507,I225966,I226091,);
nand I_13150 (I226099,I226091,I564929);
not I_13151 (I226116,I226099);
DFFARX1 I_13152 (I226116,I2507,I225966,I226142,);
not I_13153 (I225958,I226142);
nor I_13154 (I226164,I225992,I226099);
nor I_13155 (I225940,I226043,I226164);
DFFARX1 I_13156 (I564917,I2507,I225966,I226204,);
DFFARX1 I_13157 (I226204,I2507,I225966,I226221,);
not I_13158 (I226229,I226221);
not I_13159 (I226246,I226204);
nand I_13160 (I225943,I226246,I226065);
nand I_13161 (I226277,I564926,I564932);
and I_13162 (I226294,I226277,I564917);
DFFARX1 I_13163 (I226294,I2507,I225966,I226320,);
nor I_13164 (I226328,I226320,I225992);
DFFARX1 I_13165 (I226328,I2507,I225966,I225931,);
DFFARX1 I_13166 (I226320,I2507,I225966,I225949,);
nor I_13167 (I226373,I564920,I564932);
not I_13168 (I226390,I226373);
nor I_13169 (I225952,I226229,I226390);
nand I_13170 (I225937,I226246,I226390);
nor I_13171 (I225946,I225992,I226373);
DFFARX1 I_13172 (I226373,I2507,I225966,I225955,);
not I_13173 (I226493,I2514);
DFFARX1 I_13174 (I275396,I2507,I226493,I226519,);
nand I_13175 (I226527,I275408,I275387);
and I_13176 (I226544,I226527,I275411);
DFFARX1 I_13177 (I226544,I2507,I226493,I226570,);
nor I_13178 (I226461,I226570,I226519);
not I_13179 (I226592,I226570);
DFFARX1 I_13180 (I275402,I2507,I226493,I226618,);
nand I_13181 (I226626,I226618,I275384);
not I_13182 (I226643,I226626);
DFFARX1 I_13183 (I226643,I2507,I226493,I226669,);
not I_13184 (I226485,I226669);
nor I_13185 (I226691,I226519,I226626);
nor I_13186 (I226467,I226570,I226691);
DFFARX1 I_13187 (I275399,I2507,I226493,I226731,);
DFFARX1 I_13188 (I226731,I2507,I226493,I226748,);
not I_13189 (I226756,I226748);
not I_13190 (I226773,I226731);
nand I_13191 (I226470,I226773,I226592);
nand I_13192 (I226804,I275384,I275390);
and I_13193 (I226821,I226804,I275393);
DFFARX1 I_13194 (I226821,I2507,I226493,I226847,);
nor I_13195 (I226855,I226847,I226519);
DFFARX1 I_13196 (I226855,I2507,I226493,I226458,);
DFFARX1 I_13197 (I226847,I2507,I226493,I226476,);
nor I_13198 (I226900,I275405,I275390);
not I_13199 (I226917,I226900);
nor I_13200 (I226479,I226756,I226917);
nand I_13201 (I226464,I226773,I226917);
nor I_13202 (I226473,I226519,I226900);
DFFARX1 I_13203 (I226900,I2507,I226493,I226482,);
not I_13204 (I227020,I2514);
DFFARX1 I_13205 (I156214,I2507,I227020,I227046,);
nand I_13206 (I227054,I156214,I156220);
and I_13207 (I227071,I227054,I156238);
DFFARX1 I_13208 (I227071,I2507,I227020,I227097,);
nor I_13209 (I226988,I227097,I227046);
not I_13210 (I227119,I227097);
DFFARX1 I_13211 (I156226,I2507,I227020,I227145,);
nand I_13212 (I227153,I227145,I156223);
not I_13213 (I227170,I227153);
DFFARX1 I_13214 (I227170,I2507,I227020,I227196,);
not I_13215 (I227012,I227196);
nor I_13216 (I227218,I227046,I227153);
nor I_13217 (I226994,I227097,I227218);
DFFARX1 I_13218 (I156232,I2507,I227020,I227258,);
DFFARX1 I_13219 (I227258,I2507,I227020,I227275,);
not I_13220 (I227283,I227275);
not I_13221 (I227300,I227258);
nand I_13222 (I226997,I227300,I227119);
nand I_13223 (I227331,I156217,I156217);
and I_13224 (I227348,I227331,I156229);
DFFARX1 I_13225 (I227348,I2507,I227020,I227374,);
nor I_13226 (I227382,I227374,I227046);
DFFARX1 I_13227 (I227382,I2507,I227020,I226985,);
DFFARX1 I_13228 (I227374,I2507,I227020,I227003,);
nor I_13229 (I227427,I156235,I156217);
not I_13230 (I227444,I227427);
nor I_13231 (I227006,I227283,I227444);
nand I_13232 (I226991,I227300,I227444);
nor I_13233 (I227000,I227046,I227427);
DFFARX1 I_13234 (I227427,I2507,I227020,I227009,);
not I_13235 (I227547,I2514);
DFFARX1 I_13236 (I650696,I2507,I227547,I227573,);
DFFARX1 I_13237 (I227573,I2507,I227547,I227590,);
not I_13238 (I227539,I227590);
not I_13239 (I227612,I227573);
nand I_13240 (I227629,I650708,I650711);
and I_13241 (I227646,I227629,I650714);
DFFARX1 I_13242 (I227646,I2507,I227547,I227672,);
not I_13243 (I227680,I227672);
DFFARX1 I_13244 (I650699,I2507,I227547,I227706,);
and I_13245 (I227714,I227706,I650705);
nand I_13246 (I227731,I227706,I650705);
nand I_13247 (I227518,I227680,I227731);
DFFARX1 I_13248 (I650693,I2507,I227547,I227771,);
nor I_13249 (I227779,I227771,I227714);
DFFARX1 I_13250 (I227779,I2507,I227547,I227512,);
nor I_13251 (I227527,I227771,I227672);
nand I_13252 (I227824,I650696,I650717);
and I_13253 (I227841,I227824,I650702);
DFFARX1 I_13254 (I227841,I2507,I227547,I227867,);
nor I_13255 (I227515,I227867,I227771);
not I_13256 (I227889,I227867);
nor I_13257 (I227906,I227889,I227680);
nor I_13258 (I227923,I227612,I227906);
DFFARX1 I_13259 (I227923,I2507,I227547,I227530,);
nor I_13260 (I227954,I227889,I227771);
nor I_13261 (I227971,I650693,I650717);
nor I_13262 (I227521,I227971,I227954);
not I_13263 (I228002,I227971);
nand I_13264 (I227524,I227731,I228002);
DFFARX1 I_13265 (I227971,I2507,I227547,I227536,);
DFFARX1 I_13266 (I227971,I2507,I227547,I227533,);
not I_13267 (I228091,I2514);
DFFARX1 I_13268 (I578038,I2507,I228091,I228117,);
DFFARX1 I_13269 (I228117,I2507,I228091,I228134,);
not I_13270 (I228083,I228134);
not I_13271 (I228156,I228117);
nand I_13272 (I228173,I578050,I578038);
and I_13273 (I228190,I228173,I578041);
DFFARX1 I_13274 (I228190,I2507,I228091,I228216,);
not I_13275 (I228224,I228216);
DFFARX1 I_13276 (I578059,I2507,I228091,I228250,);
and I_13277 (I228258,I228250,I578035);
nand I_13278 (I228275,I228250,I578035);
nand I_13279 (I228062,I228224,I228275);
DFFARX1 I_13280 (I578053,I2507,I228091,I228315,);
nor I_13281 (I228323,I228315,I228258);
DFFARX1 I_13282 (I228323,I2507,I228091,I228056,);
nor I_13283 (I228071,I228315,I228216);
nand I_13284 (I228368,I578047,I578044);
and I_13285 (I228385,I228368,I578056);
DFFARX1 I_13286 (I228385,I2507,I228091,I228411,);
nor I_13287 (I228059,I228411,I228315);
not I_13288 (I228433,I228411);
nor I_13289 (I228450,I228433,I228224);
nor I_13290 (I228467,I228156,I228450);
DFFARX1 I_13291 (I228467,I2507,I228091,I228074,);
nor I_13292 (I228498,I228433,I228315);
nor I_13293 (I228515,I578035,I578044);
nor I_13294 (I228065,I228515,I228498);
not I_13295 (I228546,I228515);
nand I_13296 (I228068,I228275,I228546);
DFFARX1 I_13297 (I228515,I2507,I228091,I228080,);
DFFARX1 I_13298 (I228515,I2507,I228091,I228077,);
not I_13299 (I228635,I2514);
DFFARX1 I_13300 (I351292,I2507,I228635,I228661,);
DFFARX1 I_13301 (I228661,I2507,I228635,I228678,);
not I_13302 (I228627,I228678);
not I_13303 (I228700,I228661);
nand I_13304 (I228717,I351313,I351304);
and I_13305 (I228734,I228717,I351292);
DFFARX1 I_13306 (I228734,I2507,I228635,I228760,);
not I_13307 (I228768,I228760);
DFFARX1 I_13308 (I351298,I2507,I228635,I228794,);
and I_13309 (I228802,I228794,I351295);
nand I_13310 (I228819,I228794,I351295);
nand I_13311 (I228606,I228768,I228819);
DFFARX1 I_13312 (I351289,I2507,I228635,I228859,);
nor I_13313 (I228867,I228859,I228802);
DFFARX1 I_13314 (I228867,I2507,I228635,I228600,);
nor I_13315 (I228615,I228859,I228760);
nand I_13316 (I228912,I351289,I351301);
and I_13317 (I228929,I228912,I351310);
DFFARX1 I_13318 (I228929,I2507,I228635,I228955,);
nor I_13319 (I228603,I228955,I228859);
not I_13320 (I228977,I228955);
nor I_13321 (I228994,I228977,I228768);
nor I_13322 (I229011,I228700,I228994);
DFFARX1 I_13323 (I229011,I2507,I228635,I228618,);
nor I_13324 (I229042,I228977,I228859);
nor I_13325 (I229059,I351307,I351301);
nor I_13326 (I228609,I229059,I229042);
not I_13327 (I229090,I229059);
nand I_13328 (I228612,I228819,I229090);
DFFARX1 I_13329 (I229059,I2507,I228635,I228624,);
DFFARX1 I_13330 (I229059,I2507,I228635,I228621,);
not I_13331 (I229179,I2514);
DFFARX1 I_13332 (I128258,I2507,I229179,I229205,);
DFFARX1 I_13333 (I229205,I2507,I229179,I229222,);
not I_13334 (I229171,I229222);
not I_13335 (I229244,I229205);
nand I_13336 (I229261,I128270,I128249);
and I_13337 (I229278,I229261,I128252);
DFFARX1 I_13338 (I229278,I2507,I229179,I229304,);
not I_13339 (I229312,I229304);
DFFARX1 I_13340 (I128261,I2507,I229179,I229338,);
and I_13341 (I229346,I229338,I128273);
nand I_13342 (I229363,I229338,I128273);
nand I_13343 (I229150,I229312,I229363);
DFFARX1 I_13344 (I128267,I2507,I229179,I229403,);
nor I_13345 (I229411,I229403,I229346);
DFFARX1 I_13346 (I229411,I2507,I229179,I229144,);
nor I_13347 (I229159,I229403,I229304);
nand I_13348 (I229456,I128255,I128252);
and I_13349 (I229473,I229456,I128264);
DFFARX1 I_13350 (I229473,I2507,I229179,I229499,);
nor I_13351 (I229147,I229499,I229403);
not I_13352 (I229521,I229499);
nor I_13353 (I229538,I229521,I229312);
nor I_13354 (I229555,I229244,I229538);
DFFARX1 I_13355 (I229555,I2507,I229179,I229162,);
nor I_13356 (I229586,I229521,I229403);
nor I_13357 (I229603,I128249,I128252);
nor I_13358 (I229153,I229603,I229586);
not I_13359 (I229634,I229603);
nand I_13360 (I229156,I229363,I229634);
DFFARX1 I_13361 (I229603,I2507,I229179,I229168,);
DFFARX1 I_13362 (I229603,I2507,I229179,I229165,);
not I_13363 (I229723,I2514);
DFFARX1 I_13364 (I390596,I2507,I229723,I229749,);
DFFARX1 I_13365 (I229749,I2507,I229723,I229766,);
not I_13366 (I229715,I229766);
not I_13367 (I229788,I229749);
nand I_13368 (I229805,I390617,I390608);
and I_13369 (I229822,I229805,I390596);
DFFARX1 I_13370 (I229822,I2507,I229723,I229848,);
not I_13371 (I229856,I229848);
DFFARX1 I_13372 (I390602,I2507,I229723,I229882,);
and I_13373 (I229890,I229882,I390599);
nand I_13374 (I229907,I229882,I390599);
nand I_13375 (I229694,I229856,I229907);
DFFARX1 I_13376 (I390593,I2507,I229723,I229947,);
nor I_13377 (I229955,I229947,I229890);
DFFARX1 I_13378 (I229955,I2507,I229723,I229688,);
nor I_13379 (I229703,I229947,I229848);
nand I_13380 (I230000,I390593,I390605);
and I_13381 (I230017,I230000,I390614);
DFFARX1 I_13382 (I230017,I2507,I229723,I230043,);
nor I_13383 (I229691,I230043,I229947);
not I_13384 (I230065,I230043);
nor I_13385 (I230082,I230065,I229856);
nor I_13386 (I230099,I229788,I230082);
DFFARX1 I_13387 (I230099,I2507,I229723,I229706,);
nor I_13388 (I230130,I230065,I229947);
nor I_13389 (I230147,I390611,I390605);
nor I_13390 (I229697,I230147,I230130);
not I_13391 (I230178,I230147);
nand I_13392 (I229700,I229907,I230178);
DFFARX1 I_13393 (I230147,I2507,I229723,I229712,);
DFFARX1 I_13394 (I230147,I2507,I229723,I229709,);
not I_13395 (I230267,I2514);
DFFARX1 I_13396 (I432340,I2507,I230267,I230293,);
DFFARX1 I_13397 (I230293,I2507,I230267,I230310,);
not I_13398 (I230259,I230310);
not I_13399 (I230332,I230293);
nand I_13400 (I230349,I432334,I432331);
and I_13401 (I230366,I230349,I432346);
DFFARX1 I_13402 (I230366,I2507,I230267,I230392,);
not I_13403 (I230400,I230392);
DFFARX1 I_13404 (I432334,I2507,I230267,I230426,);
and I_13405 (I230434,I230426,I432328);
nand I_13406 (I230451,I230426,I432328);
nand I_13407 (I230238,I230400,I230451);
DFFARX1 I_13408 (I432328,I2507,I230267,I230491,);
nor I_13409 (I230499,I230491,I230434);
DFFARX1 I_13410 (I230499,I2507,I230267,I230232,);
nor I_13411 (I230247,I230491,I230392);
nand I_13412 (I230544,I432343,I432337);
and I_13413 (I230561,I230544,I432331);
DFFARX1 I_13414 (I230561,I2507,I230267,I230587,);
nor I_13415 (I230235,I230587,I230491);
not I_13416 (I230609,I230587);
nor I_13417 (I230626,I230609,I230400);
nor I_13418 (I230643,I230332,I230626);
DFFARX1 I_13419 (I230643,I2507,I230267,I230250,);
nor I_13420 (I230674,I230609,I230491);
nor I_13421 (I230691,I432349,I432337);
nor I_13422 (I230241,I230691,I230674);
not I_13423 (I230722,I230691);
nand I_13424 (I230244,I230451,I230722);
DFFARX1 I_13425 (I230691,I2507,I230267,I230256,);
DFFARX1 I_13426 (I230691,I2507,I230267,I230253,);
not I_13427 (I230811,I2514);
DFFARX1 I_13428 (I59915,I2507,I230811,I230837,);
DFFARX1 I_13429 (I230837,I2507,I230811,I230854,);
not I_13430 (I230803,I230854);
not I_13431 (I230876,I230837);
nand I_13432 (I230893,I59930,I59909);
and I_13433 (I230910,I230893,I59912);
DFFARX1 I_13434 (I230910,I2507,I230811,I230936,);
not I_13435 (I230944,I230936);
DFFARX1 I_13436 (I59918,I2507,I230811,I230970,);
and I_13437 (I230978,I230970,I59912);
nand I_13438 (I230995,I230970,I59912);
nand I_13439 (I230782,I230944,I230995);
DFFARX1 I_13440 (I59927,I2507,I230811,I231035,);
nor I_13441 (I231043,I231035,I230978);
DFFARX1 I_13442 (I231043,I2507,I230811,I230776,);
nor I_13443 (I230791,I231035,I230936);
nand I_13444 (I231088,I59909,I59924);
and I_13445 (I231105,I231088,I59921);
DFFARX1 I_13446 (I231105,I2507,I230811,I231131,);
nor I_13447 (I230779,I231131,I231035);
not I_13448 (I231153,I231131);
nor I_13449 (I231170,I231153,I230944);
nor I_13450 (I231187,I230876,I231170);
DFFARX1 I_13451 (I231187,I2507,I230811,I230794,);
nor I_13452 (I231218,I231153,I231035);
nor I_13453 (I231235,I59933,I59924);
nor I_13454 (I230785,I231235,I231218);
not I_13455 (I231266,I231235);
nand I_13456 (I230788,I230995,I231266);
DFFARX1 I_13457 (I231235,I2507,I230811,I230800,);
DFFARX1 I_13458 (I231235,I2507,I230811,I230797,);
not I_13459 (I231355,I2514);
DFFARX1 I_13460 (I165347,I2507,I231355,I231381,);
DFFARX1 I_13461 (I231381,I2507,I231355,I231398,);
not I_13462 (I231347,I231398);
not I_13463 (I231420,I231381);
nand I_13464 (I231437,I165326,I165350);
and I_13465 (I231454,I231437,I165353);
DFFARX1 I_13466 (I231454,I2507,I231355,I231480,);
not I_13467 (I231488,I231480);
DFFARX1 I_13468 (I165335,I2507,I231355,I231514,);
and I_13469 (I231522,I231514,I165341);
nand I_13470 (I231539,I231514,I165341);
nand I_13471 (I231326,I231488,I231539);
DFFARX1 I_13472 (I165329,I2507,I231355,I231579,);
nor I_13473 (I231587,I231579,I231522);
DFFARX1 I_13474 (I231587,I2507,I231355,I231320,);
nor I_13475 (I231335,I231579,I231480);
nand I_13476 (I231632,I165338,I165326);
and I_13477 (I231649,I231632,I165332);
DFFARX1 I_13478 (I231649,I2507,I231355,I231675,);
nor I_13479 (I231323,I231675,I231579);
not I_13480 (I231697,I231675);
nor I_13481 (I231714,I231697,I231488);
nor I_13482 (I231731,I231420,I231714);
DFFARX1 I_13483 (I231731,I2507,I231355,I231338,);
nor I_13484 (I231762,I231697,I231579);
nor I_13485 (I231779,I165344,I165326);
nor I_13486 (I231329,I231779,I231762);
not I_13487 (I231810,I231779);
nand I_13488 (I231332,I231539,I231810);
DFFARX1 I_13489 (I231779,I2507,I231355,I231344,);
DFFARX1 I_13490 (I231779,I2507,I231355,I231341,);
not I_13491 (I231899,I2514);
DFFARX1 I_13492 (I546398,I2507,I231899,I231925,);
DFFARX1 I_13493 (I231925,I2507,I231899,I231942,);
not I_13494 (I231891,I231942);
not I_13495 (I231964,I231925);
nand I_13496 (I231981,I546398,I546416);
and I_13497 (I231998,I231981,I546410);
DFFARX1 I_13498 (I231998,I2507,I231899,I232024,);
not I_13499 (I232032,I232024);
DFFARX1 I_13500 (I546404,I2507,I231899,I232058,);
and I_13501 (I232066,I232058,I546413);
nand I_13502 (I232083,I232058,I546413);
nand I_13503 (I231870,I232032,I232083);
DFFARX1 I_13504 (I546401,I2507,I231899,I232123,);
nor I_13505 (I232131,I232123,I232066);
DFFARX1 I_13506 (I232131,I2507,I231899,I231864,);
nor I_13507 (I231879,I232123,I232024);
nand I_13508 (I232176,I546401,I546419);
and I_13509 (I232193,I232176,I546404);
DFFARX1 I_13510 (I232193,I2507,I231899,I232219,);
nor I_13511 (I231867,I232219,I232123);
not I_13512 (I232241,I232219);
nor I_13513 (I232258,I232241,I232032);
nor I_13514 (I232275,I231964,I232258);
DFFARX1 I_13515 (I232275,I2507,I231899,I231882,);
nor I_13516 (I232306,I232241,I232123);
nor I_13517 (I232323,I546407,I546419);
nor I_13518 (I231873,I232323,I232306);
not I_13519 (I232354,I232323);
nand I_13520 (I231876,I232083,I232354);
DFFARX1 I_13521 (I232323,I2507,I231899,I231888,);
DFFARX1 I_13522 (I232323,I2507,I231899,I231885,);
not I_13523 (I232443,I2514);
DFFARX1 I_13524 (I186954,I2507,I232443,I232469,);
DFFARX1 I_13525 (I232469,I2507,I232443,I232486,);
not I_13526 (I232435,I232486);
not I_13527 (I232508,I232469);
nand I_13528 (I232525,I186933,I186957);
and I_13529 (I232542,I232525,I186960);
DFFARX1 I_13530 (I232542,I2507,I232443,I232568,);
not I_13531 (I232576,I232568);
DFFARX1 I_13532 (I186942,I2507,I232443,I232602,);
and I_13533 (I232610,I232602,I186948);
nand I_13534 (I232627,I232602,I186948);
nand I_13535 (I232414,I232576,I232627);
DFFARX1 I_13536 (I186936,I2507,I232443,I232667,);
nor I_13537 (I232675,I232667,I232610);
DFFARX1 I_13538 (I232675,I2507,I232443,I232408,);
nor I_13539 (I232423,I232667,I232568);
nand I_13540 (I232720,I186945,I186933);
and I_13541 (I232737,I232720,I186939);
DFFARX1 I_13542 (I232737,I2507,I232443,I232763,);
nor I_13543 (I232411,I232763,I232667);
not I_13544 (I232785,I232763);
nor I_13545 (I232802,I232785,I232576);
nor I_13546 (I232819,I232508,I232802);
DFFARX1 I_13547 (I232819,I2507,I232443,I232426,);
nor I_13548 (I232850,I232785,I232667);
nor I_13549 (I232867,I186951,I186933);
nor I_13550 (I232417,I232867,I232850);
not I_13551 (I232898,I232867);
nand I_13552 (I232420,I232627,I232898);
DFFARX1 I_13553 (I232867,I2507,I232443,I232432,);
DFFARX1 I_13554 (I232867,I2507,I232443,I232429,);
not I_13555 (I232987,I2514);
DFFARX1 I_13556 (I427010,I2507,I232987,I233013,);
DFFARX1 I_13557 (I233013,I2507,I232987,I233030,);
not I_13558 (I232979,I233030);
not I_13559 (I233052,I233013);
nand I_13560 (I233069,I427031,I427022);
and I_13561 (I233086,I233069,I427010);
DFFARX1 I_13562 (I233086,I2507,I232987,I233112,);
not I_13563 (I233120,I233112);
DFFARX1 I_13564 (I427016,I2507,I232987,I233146,);
and I_13565 (I233154,I233146,I427013);
nand I_13566 (I233171,I233146,I427013);
nand I_13567 (I232958,I233120,I233171);
DFFARX1 I_13568 (I427007,I2507,I232987,I233211,);
nor I_13569 (I233219,I233211,I233154);
DFFARX1 I_13570 (I233219,I2507,I232987,I232952,);
nor I_13571 (I232967,I233211,I233112);
nand I_13572 (I233264,I427007,I427019);
and I_13573 (I233281,I233264,I427028);
DFFARX1 I_13574 (I233281,I2507,I232987,I233307,);
nor I_13575 (I232955,I233307,I233211);
not I_13576 (I233329,I233307);
nor I_13577 (I233346,I233329,I233120);
nor I_13578 (I233363,I233052,I233346);
DFFARX1 I_13579 (I233363,I2507,I232987,I232970,);
nor I_13580 (I233394,I233329,I233211);
nor I_13581 (I233411,I427025,I427019);
nor I_13582 (I232961,I233411,I233394);
not I_13583 (I233442,I233411);
nand I_13584 (I232964,I233171,I233442);
DFFARX1 I_13585 (I233411,I2507,I232987,I232976,);
DFFARX1 I_13586 (I233411,I2507,I232987,I232973,);
not I_13587 (I233531,I2514);
DFFARX1 I_13588 (I163239,I2507,I233531,I233557,);
DFFARX1 I_13589 (I233557,I2507,I233531,I233574,);
not I_13590 (I233523,I233574);
not I_13591 (I233596,I233557);
nand I_13592 (I233613,I163218,I163242);
and I_13593 (I233630,I233613,I163245);
DFFARX1 I_13594 (I233630,I2507,I233531,I233656,);
not I_13595 (I233664,I233656);
DFFARX1 I_13596 (I163227,I2507,I233531,I233690,);
and I_13597 (I233698,I233690,I163233);
nand I_13598 (I233715,I233690,I163233);
nand I_13599 (I233502,I233664,I233715);
DFFARX1 I_13600 (I163221,I2507,I233531,I233755,);
nor I_13601 (I233763,I233755,I233698);
DFFARX1 I_13602 (I233763,I2507,I233531,I233496,);
nor I_13603 (I233511,I233755,I233656);
nand I_13604 (I233808,I163230,I163218);
and I_13605 (I233825,I233808,I163224);
DFFARX1 I_13606 (I233825,I2507,I233531,I233851,);
nor I_13607 (I233499,I233851,I233755);
not I_13608 (I233873,I233851);
nor I_13609 (I233890,I233873,I233664);
nor I_13610 (I233907,I233596,I233890);
DFFARX1 I_13611 (I233907,I2507,I233531,I233514,);
nor I_13612 (I233938,I233873,I233755);
nor I_13613 (I233955,I163236,I163218);
nor I_13614 (I233505,I233955,I233938);
not I_13615 (I233986,I233955);
nand I_13616 (I233508,I233715,I233986);
DFFARX1 I_13617 (I233955,I2507,I233531,I233520,);
DFFARX1 I_13618 (I233955,I2507,I233531,I233517,);
not I_13619 (I234075,I2514);
DFFARX1 I_13620 (I716850,I2507,I234075,I234101,);
DFFARX1 I_13621 (I234101,I2507,I234075,I234118,);
not I_13622 (I234067,I234118);
not I_13623 (I234140,I234101);
nand I_13624 (I234157,I716826,I716847);
and I_13625 (I234174,I234157,I716844);
DFFARX1 I_13626 (I234174,I2507,I234075,I234200,);
not I_13627 (I234208,I234200);
DFFARX1 I_13628 (I716823,I2507,I234075,I234234,);
and I_13629 (I234242,I234234,I716835);
nand I_13630 (I234259,I234234,I716835);
nand I_13631 (I234046,I234208,I234259);
DFFARX1 I_13632 (I716838,I2507,I234075,I234299,);
nor I_13633 (I234307,I234299,I234242);
DFFARX1 I_13634 (I234307,I2507,I234075,I234040,);
nor I_13635 (I234055,I234299,I234200);
nand I_13636 (I234352,I716841,I716829);
and I_13637 (I234369,I234352,I716832);
DFFARX1 I_13638 (I234369,I2507,I234075,I234395,);
nor I_13639 (I234043,I234395,I234299);
not I_13640 (I234417,I234395);
nor I_13641 (I234434,I234417,I234208);
nor I_13642 (I234451,I234140,I234434);
DFFARX1 I_13643 (I234451,I2507,I234075,I234058,);
nor I_13644 (I234482,I234417,I234299);
nor I_13645 (I234499,I716823,I716829);
nor I_13646 (I234049,I234499,I234482);
not I_13647 (I234530,I234499);
nand I_13648 (I234052,I234259,I234530);
DFFARX1 I_13649 (I234499,I2507,I234075,I234064,);
DFFARX1 I_13650 (I234499,I2507,I234075,I234061,);
not I_13651 (I234619,I2514);
DFFARX1 I_13652 (I333374,I2507,I234619,I234645,);
DFFARX1 I_13653 (I234645,I2507,I234619,I234662,);
not I_13654 (I234611,I234662);
not I_13655 (I234684,I234645);
nand I_13656 (I234701,I333371,I333392);
and I_13657 (I234718,I234701,I333395);
DFFARX1 I_13658 (I234718,I2507,I234619,I234744,);
not I_13659 (I234752,I234744);
DFFARX1 I_13660 (I333380,I2507,I234619,I234778,);
and I_13661 (I234786,I234778,I333383);
nand I_13662 (I234803,I234778,I333383);
nand I_13663 (I234590,I234752,I234803);
DFFARX1 I_13664 (I333386,I2507,I234619,I234843,);
nor I_13665 (I234851,I234843,I234786);
DFFARX1 I_13666 (I234851,I2507,I234619,I234584,);
nor I_13667 (I234599,I234843,I234744);
nand I_13668 (I234896,I333371,I333377);
and I_13669 (I234913,I234896,I333389);
DFFARX1 I_13670 (I234913,I2507,I234619,I234939,);
nor I_13671 (I234587,I234939,I234843);
not I_13672 (I234961,I234939);
nor I_13673 (I234978,I234961,I234752);
nor I_13674 (I234995,I234684,I234978);
DFFARX1 I_13675 (I234995,I2507,I234619,I234602,);
nor I_13676 (I235026,I234961,I234843);
nor I_13677 (I235043,I333374,I333377);
nor I_13678 (I234593,I235043,I235026);
not I_13679 (I235074,I235043);
nand I_13680 (I234596,I234803,I235074);
DFFARX1 I_13681 (I235043,I2507,I234619,I234608,);
DFFARX1 I_13682 (I235043,I2507,I234619,I234605,);
not I_13683 (I235163,I2514);
DFFARX1 I_13684 (I63077,I2507,I235163,I235189,);
DFFARX1 I_13685 (I235189,I2507,I235163,I235206,);
not I_13686 (I235155,I235206);
not I_13687 (I235228,I235189);
nand I_13688 (I235245,I63092,I63071);
and I_13689 (I235262,I235245,I63074);
DFFARX1 I_13690 (I235262,I2507,I235163,I235288,);
not I_13691 (I235296,I235288);
DFFARX1 I_13692 (I63080,I2507,I235163,I235322,);
and I_13693 (I235330,I235322,I63074);
nand I_13694 (I235347,I235322,I63074);
nand I_13695 (I235134,I235296,I235347);
DFFARX1 I_13696 (I63089,I2507,I235163,I235387,);
nor I_13697 (I235395,I235387,I235330);
DFFARX1 I_13698 (I235395,I2507,I235163,I235128,);
nor I_13699 (I235143,I235387,I235288);
nand I_13700 (I235440,I63071,I63086);
and I_13701 (I235457,I235440,I63083);
DFFARX1 I_13702 (I235457,I2507,I235163,I235483,);
nor I_13703 (I235131,I235483,I235387);
not I_13704 (I235505,I235483);
nor I_13705 (I235522,I235505,I235296);
nor I_13706 (I235539,I235228,I235522);
DFFARX1 I_13707 (I235539,I2507,I235163,I235146,);
nor I_13708 (I235570,I235505,I235387);
nor I_13709 (I235587,I63095,I63086);
nor I_13710 (I235137,I235587,I235570);
not I_13711 (I235618,I235587);
nand I_13712 (I235140,I235347,I235618);
DFFARX1 I_13713 (I235587,I2507,I235163,I235152,);
DFFARX1 I_13714 (I235587,I2507,I235163,I235149,);
not I_13715 (I235707,I2514);
DFFARX1 I_13716 (I668833,I2507,I235707,I235733,);
DFFARX1 I_13717 (I235733,I2507,I235707,I235750,);
not I_13718 (I235699,I235750);
not I_13719 (I235772,I235733);
nand I_13720 (I235789,I668830,I668827);
and I_13721 (I235806,I235789,I668815);
DFFARX1 I_13722 (I235806,I2507,I235707,I235832,);
not I_13723 (I235840,I235832);
DFFARX1 I_13724 (I668839,I2507,I235707,I235866,);
and I_13725 (I235874,I235866,I668824);
nand I_13726 (I235891,I235866,I668824);
nand I_13727 (I235678,I235840,I235891);
DFFARX1 I_13728 (I668818,I2507,I235707,I235931,);
nor I_13729 (I235939,I235931,I235874);
DFFARX1 I_13730 (I235939,I2507,I235707,I235672,);
nor I_13731 (I235687,I235931,I235832);
nand I_13732 (I235984,I668815,I668821);
and I_13733 (I236001,I235984,I668836);
DFFARX1 I_13734 (I236001,I2507,I235707,I236027,);
nor I_13735 (I235675,I236027,I235931);
not I_13736 (I236049,I236027);
nor I_13737 (I236066,I236049,I235840);
nor I_13738 (I236083,I235772,I236066);
DFFARX1 I_13739 (I236083,I2507,I235707,I235690,);
nor I_13740 (I236114,I236049,I235931);
nor I_13741 (I236131,I668818,I668821);
nor I_13742 (I235681,I236131,I236114);
not I_13743 (I236162,I236131);
nand I_13744 (I235684,I235891,I236162);
DFFARX1 I_13745 (I236131,I2507,I235707,I235696,);
DFFARX1 I_13746 (I236131,I2507,I235707,I235693,);
not I_13747 (I236251,I2514);
DFFARX1 I_13748 (I25666,I2507,I236251,I236277,);
DFFARX1 I_13749 (I236277,I2507,I236251,I236294,);
not I_13750 (I236243,I236294);
not I_13751 (I236316,I236277);
nand I_13752 (I236333,I25654,I25669);
and I_13753 (I236350,I236333,I25657);
DFFARX1 I_13754 (I236350,I2507,I236251,I236376,);
not I_13755 (I236384,I236376);
DFFARX1 I_13756 (I25678,I2507,I236251,I236410,);
and I_13757 (I236418,I236410,I25672);
nand I_13758 (I236435,I236410,I25672);
nand I_13759 (I236222,I236384,I236435);
DFFARX1 I_13760 (I25675,I2507,I236251,I236475,);
nor I_13761 (I236483,I236475,I236418);
DFFARX1 I_13762 (I236483,I2507,I236251,I236216,);
nor I_13763 (I236231,I236475,I236376);
nand I_13764 (I236528,I25654,I25657);
and I_13765 (I236545,I236528,I25660);
DFFARX1 I_13766 (I236545,I2507,I236251,I236571,);
nor I_13767 (I236219,I236571,I236475);
not I_13768 (I236593,I236571);
nor I_13769 (I236610,I236593,I236384);
nor I_13770 (I236627,I236316,I236610);
DFFARX1 I_13771 (I236627,I2507,I236251,I236234,);
nor I_13772 (I236658,I236593,I236475);
nor I_13773 (I236675,I25663,I25657);
nor I_13774 (I236225,I236675,I236658);
not I_13775 (I236706,I236675);
nand I_13776 (I236228,I236435,I236706);
DFFARX1 I_13777 (I236675,I2507,I236251,I236240,);
DFFARX1 I_13778 (I236675,I2507,I236251,I236237,);
not I_13779 (I236795,I2514);
DFFARX1 I_13780 (I104458,I2507,I236795,I236821,);
DFFARX1 I_13781 (I236821,I2507,I236795,I236838,);
not I_13782 (I236787,I236838);
not I_13783 (I236860,I236821);
nand I_13784 (I236877,I104470,I104449);
and I_13785 (I236894,I236877,I104452);
DFFARX1 I_13786 (I236894,I2507,I236795,I236920,);
not I_13787 (I236928,I236920);
DFFARX1 I_13788 (I104461,I2507,I236795,I236954,);
and I_13789 (I236962,I236954,I104473);
nand I_13790 (I236979,I236954,I104473);
nand I_13791 (I236766,I236928,I236979);
DFFARX1 I_13792 (I104467,I2507,I236795,I237019,);
nor I_13793 (I237027,I237019,I236962);
DFFARX1 I_13794 (I237027,I2507,I236795,I236760,);
nor I_13795 (I236775,I237019,I236920);
nand I_13796 (I237072,I104455,I104452);
and I_13797 (I237089,I237072,I104464);
DFFARX1 I_13798 (I237089,I2507,I236795,I237115,);
nor I_13799 (I236763,I237115,I237019);
not I_13800 (I237137,I237115);
nor I_13801 (I237154,I237137,I236928);
nor I_13802 (I237171,I236860,I237154);
DFFARX1 I_13803 (I237171,I2507,I236795,I236778,);
nor I_13804 (I237202,I237137,I237019);
nor I_13805 (I237219,I104449,I104452);
nor I_13806 (I236769,I237219,I237202);
not I_13807 (I237250,I237219);
nand I_13808 (I236772,I236979,I237250);
DFFARX1 I_13809 (I237219,I2507,I236795,I236784,);
DFFARX1 I_13810 (I237219,I2507,I236795,I236781,);
not I_13811 (I237339,I2514);
DFFARX1 I_13812 (I206980,I2507,I237339,I237365,);
DFFARX1 I_13813 (I237365,I2507,I237339,I237382,);
not I_13814 (I237331,I237382);
not I_13815 (I237404,I237365);
nand I_13816 (I237421,I206959,I206983);
and I_13817 (I237438,I237421,I206986);
DFFARX1 I_13818 (I237438,I2507,I237339,I237464,);
not I_13819 (I237472,I237464);
DFFARX1 I_13820 (I206968,I2507,I237339,I237498,);
and I_13821 (I237506,I237498,I206974);
nand I_13822 (I237523,I237498,I206974);
nand I_13823 (I237310,I237472,I237523);
DFFARX1 I_13824 (I206962,I2507,I237339,I237563,);
nor I_13825 (I237571,I237563,I237506);
DFFARX1 I_13826 (I237571,I2507,I237339,I237304,);
nor I_13827 (I237319,I237563,I237464);
nand I_13828 (I237616,I206971,I206959);
and I_13829 (I237633,I237616,I206965);
DFFARX1 I_13830 (I237633,I2507,I237339,I237659,);
nor I_13831 (I237307,I237659,I237563);
not I_13832 (I237681,I237659);
nor I_13833 (I237698,I237681,I237472);
nor I_13834 (I237715,I237404,I237698);
DFFARX1 I_13835 (I237715,I2507,I237339,I237322,);
nor I_13836 (I237746,I237681,I237563);
nor I_13837 (I237763,I206977,I206959);
nor I_13838 (I237313,I237763,I237746);
not I_13839 (I237794,I237763);
nand I_13840 (I237316,I237523,I237794);
DFFARX1 I_13841 (I237763,I2507,I237339,I237328,);
DFFARX1 I_13842 (I237763,I2507,I237339,I237325,);
not I_13843 (I237883,I2514);
DFFARX1 I_13844 (I153843,I2507,I237883,I237909,);
DFFARX1 I_13845 (I237909,I2507,I237883,I237926,);
not I_13846 (I237875,I237926);
not I_13847 (I237948,I237909);
nand I_13848 (I237965,I153855,I153834);
and I_13849 (I237982,I237965,I153837);
DFFARX1 I_13850 (I237982,I2507,I237883,I238008,);
not I_13851 (I238016,I238008);
DFFARX1 I_13852 (I153846,I2507,I237883,I238042,);
and I_13853 (I238050,I238042,I153858);
nand I_13854 (I238067,I238042,I153858);
nand I_13855 (I237854,I238016,I238067);
DFFARX1 I_13856 (I153852,I2507,I237883,I238107,);
nor I_13857 (I238115,I238107,I238050);
DFFARX1 I_13858 (I238115,I2507,I237883,I237848,);
nor I_13859 (I237863,I238107,I238008);
nand I_13860 (I238160,I153840,I153837);
and I_13861 (I238177,I238160,I153849);
DFFARX1 I_13862 (I238177,I2507,I237883,I238203,);
nor I_13863 (I237851,I238203,I238107);
not I_13864 (I238225,I238203);
nor I_13865 (I238242,I238225,I238016);
nor I_13866 (I238259,I237948,I238242);
DFFARX1 I_13867 (I238259,I2507,I237883,I237866,);
nor I_13868 (I238290,I238225,I238107);
nor I_13869 (I238307,I153834,I153837);
nor I_13870 (I237857,I238307,I238290);
not I_13871 (I238338,I238307);
nand I_13872 (I237860,I238067,I238338);
DFFARX1 I_13873 (I238307,I2507,I237883,I237872,);
DFFARX1 I_13874 (I238307,I2507,I237883,I237869,);
not I_13875 (I238427,I2514);
DFFARX1 I_13876 (I719825,I2507,I238427,I238453,);
DFFARX1 I_13877 (I238453,I2507,I238427,I238470,);
not I_13878 (I238419,I238470);
not I_13879 (I238492,I238453);
nand I_13880 (I238509,I719801,I719822);
and I_13881 (I238526,I238509,I719819);
DFFARX1 I_13882 (I238526,I2507,I238427,I238552,);
not I_13883 (I238560,I238552);
DFFARX1 I_13884 (I719798,I2507,I238427,I238586,);
and I_13885 (I238594,I238586,I719810);
nand I_13886 (I238611,I238586,I719810);
nand I_13887 (I238398,I238560,I238611);
DFFARX1 I_13888 (I719813,I2507,I238427,I238651,);
nor I_13889 (I238659,I238651,I238594);
DFFARX1 I_13890 (I238659,I2507,I238427,I238392,);
nor I_13891 (I238407,I238651,I238552);
nand I_13892 (I238704,I719816,I719804);
and I_13893 (I238721,I238704,I719807);
DFFARX1 I_13894 (I238721,I2507,I238427,I238747,);
nor I_13895 (I238395,I238747,I238651);
not I_13896 (I238769,I238747);
nor I_13897 (I238786,I238769,I238560);
nor I_13898 (I238803,I238492,I238786);
DFFARX1 I_13899 (I238803,I2507,I238427,I238410,);
nor I_13900 (I238834,I238769,I238651);
nor I_13901 (I238851,I719798,I719804);
nor I_13902 (I238401,I238851,I238834);
not I_13903 (I238882,I238851);
nand I_13904 (I238404,I238611,I238882);
DFFARX1 I_13905 (I238851,I2507,I238427,I238416,);
DFFARX1 I_13906 (I238851,I2507,I238427,I238413,);
not I_13907 (I238971,I2514);
DFFARX1 I_13908 (I82049,I2507,I238971,I238997,);
DFFARX1 I_13909 (I238997,I2507,I238971,I239014,);
not I_13910 (I238963,I239014);
not I_13911 (I239036,I238997);
nand I_13912 (I239053,I82064,I82043);
and I_13913 (I239070,I239053,I82046);
DFFARX1 I_13914 (I239070,I2507,I238971,I239096,);
not I_13915 (I239104,I239096);
DFFARX1 I_13916 (I82052,I2507,I238971,I239130,);
and I_13917 (I239138,I239130,I82046);
nand I_13918 (I239155,I239130,I82046);
nand I_13919 (I238942,I239104,I239155);
DFFARX1 I_13920 (I82061,I2507,I238971,I239195,);
nor I_13921 (I239203,I239195,I239138);
DFFARX1 I_13922 (I239203,I2507,I238971,I238936,);
nor I_13923 (I238951,I239195,I239096);
nand I_13924 (I239248,I82043,I82058);
and I_13925 (I239265,I239248,I82055);
DFFARX1 I_13926 (I239265,I2507,I238971,I239291,);
nor I_13927 (I238939,I239291,I239195);
not I_13928 (I239313,I239291);
nor I_13929 (I239330,I239313,I239104);
nor I_13930 (I239347,I239036,I239330);
DFFARX1 I_13931 (I239347,I2507,I238971,I238954,);
nor I_13932 (I239378,I239313,I239195);
nor I_13933 (I239395,I82067,I82058);
nor I_13934 (I238945,I239395,I239378);
not I_13935 (I239426,I239395);
nand I_13936 (I238948,I239155,I239426);
DFFARX1 I_13937 (I239395,I2507,I238971,I238960,);
DFFARX1 I_13938 (I239395,I2507,I238971,I238957,);
not I_13939 (I239515,I2514);
DFFARX1 I_13940 (I679237,I2507,I239515,I239541,);
DFFARX1 I_13941 (I239541,I2507,I239515,I239558,);
not I_13942 (I239507,I239558);
not I_13943 (I239580,I239541);
nand I_13944 (I239597,I679234,I679231);
and I_13945 (I239614,I239597,I679219);
DFFARX1 I_13946 (I239614,I2507,I239515,I239640,);
not I_13947 (I239648,I239640);
DFFARX1 I_13948 (I679243,I2507,I239515,I239674,);
and I_13949 (I239682,I239674,I679228);
nand I_13950 (I239699,I239674,I679228);
nand I_13951 (I239486,I239648,I239699);
DFFARX1 I_13952 (I679222,I2507,I239515,I239739,);
nor I_13953 (I239747,I239739,I239682);
DFFARX1 I_13954 (I239747,I2507,I239515,I239480,);
nor I_13955 (I239495,I239739,I239640);
nand I_13956 (I239792,I679219,I679225);
and I_13957 (I239809,I239792,I679240);
DFFARX1 I_13958 (I239809,I2507,I239515,I239835,);
nor I_13959 (I239483,I239835,I239739);
not I_13960 (I239857,I239835);
nor I_13961 (I239874,I239857,I239648);
nor I_13962 (I239891,I239580,I239874);
DFFARX1 I_13963 (I239891,I2507,I239515,I239498,);
nor I_13964 (I239922,I239857,I239739);
nor I_13965 (I239939,I679222,I679225);
nor I_13966 (I239489,I239939,I239922);
not I_13967 (I239970,I239939);
nand I_13968 (I239492,I239699,I239970);
DFFARX1 I_13969 (I239939,I2507,I239515,I239504,);
DFFARX1 I_13970 (I239939,I2507,I239515,I239501,);
not I_13971 (I240059,I2514);
DFFARX1 I_13972 (I507372,I2507,I240059,I240085,);
DFFARX1 I_13973 (I240085,I2507,I240059,I240102,);
not I_13974 (I240051,I240102);
not I_13975 (I240124,I240085);
nand I_13976 (I240141,I507387,I507375);
and I_13977 (I240158,I240141,I507366);
DFFARX1 I_13978 (I240158,I2507,I240059,I240184,);
not I_13979 (I240192,I240184);
DFFARX1 I_13980 (I507378,I2507,I240059,I240218,);
and I_13981 (I240226,I240218,I507369);
nand I_13982 (I240243,I240218,I507369);
nand I_13983 (I240030,I240192,I240243);
DFFARX1 I_13984 (I507384,I2507,I240059,I240283,);
nor I_13985 (I240291,I240283,I240226);
DFFARX1 I_13986 (I240291,I2507,I240059,I240024,);
nor I_13987 (I240039,I240283,I240184);
nand I_13988 (I240336,I507393,I507381);
and I_13989 (I240353,I240336,I507390);
DFFARX1 I_13990 (I240353,I2507,I240059,I240379,);
nor I_13991 (I240027,I240379,I240283);
not I_13992 (I240401,I240379);
nor I_13993 (I240418,I240401,I240192);
nor I_13994 (I240435,I240124,I240418);
DFFARX1 I_13995 (I240435,I2507,I240059,I240042,);
nor I_13996 (I240466,I240401,I240283);
nor I_13997 (I240483,I507366,I507381);
nor I_13998 (I240033,I240483,I240466);
not I_13999 (I240514,I240483);
nand I_14000 (I240036,I240243,I240514);
DFFARX1 I_14001 (I240483,I2507,I240059,I240048,);
DFFARX1 I_14002 (I240483,I2507,I240059,I240045,);
not I_14003 (I240603,I2514);
DFFARX1 I_14004 (I204345,I2507,I240603,I240629,);
DFFARX1 I_14005 (I240629,I2507,I240603,I240646,);
not I_14006 (I240595,I240646);
not I_14007 (I240668,I240629);
nand I_14008 (I240685,I204324,I204348);
and I_14009 (I240702,I240685,I204351);
DFFARX1 I_14010 (I240702,I2507,I240603,I240728,);
not I_14011 (I240736,I240728);
DFFARX1 I_14012 (I204333,I2507,I240603,I240762,);
and I_14013 (I240770,I240762,I204339);
nand I_14014 (I240787,I240762,I204339);
nand I_14015 (I240574,I240736,I240787);
DFFARX1 I_14016 (I204327,I2507,I240603,I240827,);
nor I_14017 (I240835,I240827,I240770);
DFFARX1 I_14018 (I240835,I2507,I240603,I240568,);
nor I_14019 (I240583,I240827,I240728);
nand I_14020 (I240880,I204336,I204324);
and I_14021 (I240897,I240880,I204330);
DFFARX1 I_14022 (I240897,I2507,I240603,I240923,);
nor I_14023 (I240571,I240923,I240827);
not I_14024 (I240945,I240923);
nor I_14025 (I240962,I240945,I240736);
nor I_14026 (I240979,I240668,I240962);
DFFARX1 I_14027 (I240979,I2507,I240603,I240586,);
nor I_14028 (I241010,I240945,I240827);
nor I_14029 (I241027,I204342,I204324);
nor I_14030 (I240577,I241027,I241010);
not I_14031 (I241058,I241027);
nand I_14032 (I240580,I240787,I241058);
DFFARX1 I_14033 (I241027,I2507,I240603,I240592,);
DFFARX1 I_14034 (I241027,I2507,I240603,I240589,);
not I_14035 (I241147,I2514);
DFFARX1 I_14036 (I517708,I2507,I241147,I241173,);
DFFARX1 I_14037 (I241173,I2507,I241147,I241190,);
not I_14038 (I241139,I241190);
not I_14039 (I241212,I241173);
nand I_14040 (I241229,I517723,I517711);
and I_14041 (I241246,I241229,I517702);
DFFARX1 I_14042 (I241246,I2507,I241147,I241272,);
not I_14043 (I241280,I241272);
DFFARX1 I_14044 (I517714,I2507,I241147,I241306,);
and I_14045 (I241314,I241306,I517705);
nand I_14046 (I241331,I241306,I517705);
nand I_14047 (I241118,I241280,I241331);
DFFARX1 I_14048 (I517720,I2507,I241147,I241371,);
nor I_14049 (I241379,I241371,I241314);
DFFARX1 I_14050 (I241379,I2507,I241147,I241112,);
nor I_14051 (I241127,I241371,I241272);
nand I_14052 (I241424,I517729,I517717);
and I_14053 (I241441,I241424,I517726);
DFFARX1 I_14054 (I241441,I2507,I241147,I241467,);
nor I_14055 (I241115,I241467,I241371);
not I_14056 (I241489,I241467);
nor I_14057 (I241506,I241489,I241280);
nor I_14058 (I241523,I241212,I241506);
DFFARX1 I_14059 (I241523,I2507,I241147,I241130,);
nor I_14060 (I241554,I241489,I241371);
nor I_14061 (I241571,I517702,I517717);
nor I_14062 (I241121,I241571,I241554);
not I_14063 (I241602,I241571);
nand I_14064 (I241124,I241331,I241602);
DFFARX1 I_14065 (I241571,I2507,I241147,I241136,);
DFFARX1 I_14066 (I241571,I2507,I241147,I241133,);
not I_14067 (I241691,I2514);
DFFARX1 I_14068 (I361696,I2507,I241691,I241717,);
DFFARX1 I_14069 (I241717,I2507,I241691,I241734,);
not I_14070 (I241683,I241734);
not I_14071 (I241756,I241717);
nand I_14072 (I241773,I361717,I361708);
and I_14073 (I241790,I241773,I361696);
DFFARX1 I_14074 (I241790,I2507,I241691,I241816,);
not I_14075 (I241824,I241816);
DFFARX1 I_14076 (I361702,I2507,I241691,I241850,);
and I_14077 (I241858,I241850,I361699);
nand I_14078 (I241875,I241850,I361699);
nand I_14079 (I241662,I241824,I241875);
DFFARX1 I_14080 (I361693,I2507,I241691,I241915,);
nor I_14081 (I241923,I241915,I241858);
DFFARX1 I_14082 (I241923,I2507,I241691,I241656,);
nor I_14083 (I241671,I241915,I241816);
nand I_14084 (I241968,I361693,I361705);
and I_14085 (I241985,I241968,I361714);
DFFARX1 I_14086 (I241985,I2507,I241691,I242011,);
nor I_14087 (I241659,I242011,I241915);
not I_14088 (I242033,I242011);
nor I_14089 (I242050,I242033,I241824);
nor I_14090 (I242067,I241756,I242050);
DFFARX1 I_14091 (I242067,I2507,I241691,I241674,);
nor I_14092 (I242098,I242033,I241915);
nor I_14093 (I242115,I361711,I361705);
nor I_14094 (I241665,I242115,I242098);
not I_14095 (I242146,I242115);
nand I_14096 (I241668,I241875,I242146);
DFFARX1 I_14097 (I242115,I2507,I241691,I241680,);
DFFARX1 I_14098 (I242115,I2507,I241691,I241677,);
not I_14099 (I242235,I2514);
DFFARX1 I_14100 (I143728,I2507,I242235,I242261,);
DFFARX1 I_14101 (I242261,I2507,I242235,I242278,);
not I_14102 (I242227,I242278);
not I_14103 (I242300,I242261);
nand I_14104 (I242317,I143740,I143719);
and I_14105 (I242334,I242317,I143722);
DFFARX1 I_14106 (I242334,I2507,I242235,I242360,);
not I_14107 (I242368,I242360);
DFFARX1 I_14108 (I143731,I2507,I242235,I242394,);
and I_14109 (I242402,I242394,I143743);
nand I_14110 (I242419,I242394,I143743);
nand I_14111 (I242206,I242368,I242419);
DFFARX1 I_14112 (I143737,I2507,I242235,I242459,);
nor I_14113 (I242467,I242459,I242402);
DFFARX1 I_14114 (I242467,I2507,I242235,I242200,);
nor I_14115 (I242215,I242459,I242360);
nand I_14116 (I242512,I143725,I143722);
and I_14117 (I242529,I242512,I143734);
DFFARX1 I_14118 (I242529,I2507,I242235,I242555,);
nor I_14119 (I242203,I242555,I242459);
not I_14120 (I242577,I242555);
nor I_14121 (I242594,I242577,I242368);
nor I_14122 (I242611,I242300,I242594);
DFFARX1 I_14123 (I242611,I2507,I242235,I242218,);
nor I_14124 (I242642,I242577,I242459);
nor I_14125 (I242659,I143719,I143722);
nor I_14126 (I242209,I242659,I242642);
not I_14127 (I242690,I242659);
nand I_14128 (I242212,I242419,I242690);
DFFARX1 I_14129 (I242659,I2507,I242235,I242224,);
DFFARX1 I_14130 (I242659,I2507,I242235,I242221,);
not I_14131 (I242779,I2514);
DFFARX1 I_14132 (I412560,I2507,I242779,I242805,);
DFFARX1 I_14133 (I242805,I2507,I242779,I242822,);
not I_14134 (I242771,I242822);
not I_14135 (I242844,I242805);
nand I_14136 (I242861,I412581,I412572);
and I_14137 (I242878,I242861,I412560);
DFFARX1 I_14138 (I242878,I2507,I242779,I242904,);
not I_14139 (I242912,I242904);
DFFARX1 I_14140 (I412566,I2507,I242779,I242938,);
and I_14141 (I242946,I242938,I412563);
nand I_14142 (I242963,I242938,I412563);
nand I_14143 (I242750,I242912,I242963);
DFFARX1 I_14144 (I412557,I2507,I242779,I243003,);
nor I_14145 (I243011,I243003,I242946);
DFFARX1 I_14146 (I243011,I2507,I242779,I242744,);
nor I_14147 (I242759,I243003,I242904);
nand I_14148 (I243056,I412557,I412569);
and I_14149 (I243073,I243056,I412578);
DFFARX1 I_14150 (I243073,I2507,I242779,I243099,);
nor I_14151 (I242747,I243099,I243003);
not I_14152 (I243121,I243099);
nor I_14153 (I243138,I243121,I242912);
nor I_14154 (I243155,I242844,I243138);
DFFARX1 I_14155 (I243155,I2507,I242779,I242762,);
nor I_14156 (I243186,I243121,I243003);
nor I_14157 (I243203,I412575,I412569);
nor I_14158 (I242753,I243203,I243186);
not I_14159 (I243234,I243203);
nand I_14160 (I242756,I242963,I243234);
DFFARX1 I_14161 (I243203,I2507,I242779,I242768,);
DFFARX1 I_14162 (I243203,I2507,I242779,I242765,);
not I_14163 (I243323,I2514);
DFFARX1 I_14164 (I28301,I2507,I243323,I243349,);
DFFARX1 I_14165 (I243349,I2507,I243323,I243366,);
not I_14166 (I243315,I243366);
not I_14167 (I243388,I243349);
nand I_14168 (I243405,I28289,I28304);
and I_14169 (I243422,I243405,I28292);
DFFARX1 I_14170 (I243422,I2507,I243323,I243448,);
not I_14171 (I243456,I243448);
DFFARX1 I_14172 (I28313,I2507,I243323,I243482,);
and I_14173 (I243490,I243482,I28307);
nand I_14174 (I243507,I243482,I28307);
nand I_14175 (I243294,I243456,I243507);
DFFARX1 I_14176 (I28310,I2507,I243323,I243547,);
nor I_14177 (I243555,I243547,I243490);
DFFARX1 I_14178 (I243555,I2507,I243323,I243288,);
nor I_14179 (I243303,I243547,I243448);
nand I_14180 (I243600,I28289,I28292);
and I_14181 (I243617,I243600,I28295);
DFFARX1 I_14182 (I243617,I2507,I243323,I243643,);
nor I_14183 (I243291,I243643,I243547);
not I_14184 (I243665,I243643);
nor I_14185 (I243682,I243665,I243456);
nor I_14186 (I243699,I243388,I243682);
DFFARX1 I_14187 (I243699,I2507,I243323,I243306,);
nor I_14188 (I243730,I243665,I243547);
nor I_14189 (I243747,I28298,I28292);
nor I_14190 (I243297,I243747,I243730);
not I_14191 (I243778,I243747);
nand I_14192 (I243300,I243507,I243778);
DFFARX1 I_14193 (I243747,I2507,I243323,I243312,);
DFFARX1 I_14194 (I243747,I2507,I243323,I243309,);
not I_14195 (I243867,I2514);
DFFARX1 I_14196 (I423542,I2507,I243867,I243893,);
DFFARX1 I_14197 (I243893,I2507,I243867,I243910,);
not I_14198 (I243859,I243910);
not I_14199 (I243932,I243893);
nand I_14200 (I243949,I423563,I423554);
and I_14201 (I243966,I243949,I423542);
DFFARX1 I_14202 (I243966,I2507,I243867,I243992,);
not I_14203 (I244000,I243992);
DFFARX1 I_14204 (I423548,I2507,I243867,I244026,);
and I_14205 (I244034,I244026,I423545);
nand I_14206 (I244051,I244026,I423545);
nand I_14207 (I243838,I244000,I244051);
DFFARX1 I_14208 (I423539,I2507,I243867,I244091,);
nor I_14209 (I244099,I244091,I244034);
DFFARX1 I_14210 (I244099,I2507,I243867,I243832,);
nor I_14211 (I243847,I244091,I243992);
nand I_14212 (I244144,I423539,I423551);
and I_14213 (I244161,I244144,I423560);
DFFARX1 I_14214 (I244161,I2507,I243867,I244187,);
nor I_14215 (I243835,I244187,I244091);
not I_14216 (I244209,I244187);
nor I_14217 (I244226,I244209,I244000);
nor I_14218 (I244243,I243932,I244226);
DFFARX1 I_14219 (I244243,I2507,I243867,I243850,);
nor I_14220 (I244274,I244209,I244091);
nor I_14221 (I244291,I423557,I423551);
nor I_14222 (I243841,I244291,I244274);
not I_14223 (I244322,I244291);
nand I_14224 (I243844,I244051,I244322);
DFFARX1 I_14225 (I244291,I2507,I243867,I243856,);
DFFARX1 I_14226 (I244291,I2507,I243867,I243853,);
not I_14227 (I244411,I2514);
DFFARX1 I_14228 (I179576,I2507,I244411,I244437,);
DFFARX1 I_14229 (I244437,I2507,I244411,I244454,);
not I_14230 (I244403,I244454);
not I_14231 (I244476,I244437);
nand I_14232 (I244493,I179555,I179579);
and I_14233 (I244510,I244493,I179582);
DFFARX1 I_14234 (I244510,I2507,I244411,I244536,);
not I_14235 (I244544,I244536);
DFFARX1 I_14236 (I179564,I2507,I244411,I244570,);
and I_14237 (I244578,I244570,I179570);
nand I_14238 (I244595,I244570,I179570);
nand I_14239 (I244382,I244544,I244595);
DFFARX1 I_14240 (I179558,I2507,I244411,I244635,);
nor I_14241 (I244643,I244635,I244578);
DFFARX1 I_14242 (I244643,I2507,I244411,I244376,);
nor I_14243 (I244391,I244635,I244536);
nand I_14244 (I244688,I179567,I179555);
and I_14245 (I244705,I244688,I179561);
DFFARX1 I_14246 (I244705,I2507,I244411,I244731,);
nor I_14247 (I244379,I244731,I244635);
not I_14248 (I244753,I244731);
nor I_14249 (I244770,I244753,I244544);
nor I_14250 (I244787,I244476,I244770);
DFFARX1 I_14251 (I244787,I2507,I244411,I244394,);
nor I_14252 (I244818,I244753,I244635);
nor I_14253 (I244835,I179573,I179555);
nor I_14254 (I244385,I244835,I244818);
not I_14255 (I244866,I244835);
nand I_14256 (I244388,I244595,I244866);
DFFARX1 I_14257 (I244835,I2507,I244411,I244400,);
DFFARX1 I_14258 (I244835,I2507,I244411,I244397,);
not I_14259 (I244955,I2514);
DFFARX1 I_14260 (I573992,I2507,I244955,I244981,);
DFFARX1 I_14261 (I244981,I2507,I244955,I244998,);
not I_14262 (I244947,I244998);
not I_14263 (I245020,I244981);
nand I_14264 (I245037,I574004,I573992);
and I_14265 (I245054,I245037,I573995);
DFFARX1 I_14266 (I245054,I2507,I244955,I245080,);
not I_14267 (I245088,I245080);
DFFARX1 I_14268 (I574013,I2507,I244955,I245114,);
and I_14269 (I245122,I245114,I573989);
nand I_14270 (I245139,I245114,I573989);
nand I_14271 (I244926,I245088,I245139);
DFFARX1 I_14272 (I574007,I2507,I244955,I245179,);
nor I_14273 (I245187,I245179,I245122);
DFFARX1 I_14274 (I245187,I2507,I244955,I244920,);
nor I_14275 (I244935,I245179,I245080);
nand I_14276 (I245232,I574001,I573998);
and I_14277 (I245249,I245232,I574010);
DFFARX1 I_14278 (I245249,I2507,I244955,I245275,);
nor I_14279 (I244923,I245275,I245179);
not I_14280 (I245297,I245275);
nor I_14281 (I245314,I245297,I245088);
nor I_14282 (I245331,I245020,I245314);
DFFARX1 I_14283 (I245331,I2507,I244955,I244938,);
nor I_14284 (I245362,I245297,I245179);
nor I_14285 (I245379,I573989,I573998);
nor I_14286 (I244929,I245379,I245362);
not I_14287 (I245410,I245379);
nand I_14288 (I244932,I245139,I245410);
DFFARX1 I_14289 (I245379,I2507,I244955,I244944,);
DFFARX1 I_14290 (I245379,I2507,I244955,I244941,);
not I_14291 (I245499,I2514);
DFFARX1 I_14292 (I111003,I2507,I245499,I245525,);
DFFARX1 I_14293 (I245525,I2507,I245499,I245542,);
not I_14294 (I245491,I245542);
not I_14295 (I245564,I245525);
nand I_14296 (I245581,I111015,I110994);
and I_14297 (I245598,I245581,I110997);
DFFARX1 I_14298 (I245598,I2507,I245499,I245624,);
not I_14299 (I245632,I245624);
DFFARX1 I_14300 (I111006,I2507,I245499,I245658,);
and I_14301 (I245666,I245658,I111018);
nand I_14302 (I245683,I245658,I111018);
nand I_14303 (I245470,I245632,I245683);
DFFARX1 I_14304 (I111012,I2507,I245499,I245723,);
nor I_14305 (I245731,I245723,I245666);
DFFARX1 I_14306 (I245731,I2507,I245499,I245464,);
nor I_14307 (I245479,I245723,I245624);
nand I_14308 (I245776,I111000,I110997);
and I_14309 (I245793,I245776,I111009);
DFFARX1 I_14310 (I245793,I2507,I245499,I245819,);
nor I_14311 (I245467,I245819,I245723);
not I_14312 (I245841,I245819);
nor I_14313 (I245858,I245841,I245632);
nor I_14314 (I245875,I245564,I245858);
DFFARX1 I_14315 (I245875,I2507,I245499,I245482,);
nor I_14316 (I245906,I245841,I245723);
nor I_14317 (I245923,I110994,I110997);
nor I_14318 (I245473,I245923,I245906);
not I_14319 (I245954,I245923);
nand I_14320 (I245476,I245683,I245954);
DFFARX1 I_14321 (I245923,I2507,I245499,I245488,);
DFFARX1 I_14322 (I245923,I2507,I245499,I245485,);
not I_14323 (I246043,I2514);
DFFARX1 I_14324 (I136588,I2507,I246043,I246069,);
DFFARX1 I_14325 (I246069,I2507,I246043,I246086,);
not I_14326 (I246035,I246086);
not I_14327 (I246108,I246069);
nand I_14328 (I246125,I136600,I136579);
and I_14329 (I246142,I246125,I136582);
DFFARX1 I_14330 (I246142,I2507,I246043,I246168,);
not I_14331 (I246176,I246168);
DFFARX1 I_14332 (I136591,I2507,I246043,I246202,);
and I_14333 (I246210,I246202,I136603);
nand I_14334 (I246227,I246202,I136603);
nand I_14335 (I246014,I246176,I246227);
DFFARX1 I_14336 (I136597,I2507,I246043,I246267,);
nor I_14337 (I246275,I246267,I246210);
DFFARX1 I_14338 (I246275,I2507,I246043,I246008,);
nor I_14339 (I246023,I246267,I246168);
nand I_14340 (I246320,I136585,I136582);
and I_14341 (I246337,I246320,I136594);
DFFARX1 I_14342 (I246337,I2507,I246043,I246363,);
nor I_14343 (I246011,I246363,I246267);
not I_14344 (I246385,I246363);
nor I_14345 (I246402,I246385,I246176);
nor I_14346 (I246419,I246108,I246402);
DFFARX1 I_14347 (I246419,I2507,I246043,I246026,);
nor I_14348 (I246450,I246385,I246267);
nor I_14349 (I246467,I136579,I136582);
nor I_14350 (I246017,I246467,I246450);
not I_14351 (I246498,I246467);
nand I_14352 (I246020,I246227,I246498);
DFFARX1 I_14353 (I246467,I2507,I246043,I246032,);
DFFARX1 I_14354 (I246467,I2507,I246043,I246029,);
not I_14355 (I246587,I2514);
DFFARX1 I_14356 (I690670,I2507,I246587,I246613,);
DFFARX1 I_14357 (I246613,I2507,I246587,I246630,);
not I_14358 (I246579,I246630);
not I_14359 (I246652,I246613);
nand I_14360 (I246669,I690646,I690667);
and I_14361 (I246686,I246669,I690664);
DFFARX1 I_14362 (I246686,I2507,I246587,I246712,);
not I_14363 (I246720,I246712);
DFFARX1 I_14364 (I690643,I2507,I246587,I246746,);
and I_14365 (I246754,I246746,I690655);
nand I_14366 (I246771,I246746,I690655);
nand I_14367 (I246558,I246720,I246771);
DFFARX1 I_14368 (I690658,I2507,I246587,I246811,);
nor I_14369 (I246819,I246811,I246754);
DFFARX1 I_14370 (I246819,I2507,I246587,I246552,);
nor I_14371 (I246567,I246811,I246712);
nand I_14372 (I246864,I690661,I690649);
and I_14373 (I246881,I246864,I690652);
DFFARX1 I_14374 (I246881,I2507,I246587,I246907,);
nor I_14375 (I246555,I246907,I246811);
not I_14376 (I246929,I246907);
nor I_14377 (I246946,I246929,I246720);
nor I_14378 (I246963,I246652,I246946);
DFFARX1 I_14379 (I246963,I2507,I246587,I246570,);
nor I_14380 (I246994,I246929,I246811);
nor I_14381 (I247011,I690643,I690649);
nor I_14382 (I246561,I247011,I246994);
not I_14383 (I247042,I247011);
nand I_14384 (I246564,I246771,I247042);
DFFARX1 I_14385 (I247011,I2507,I246587,I246576,);
DFFARX1 I_14386 (I247011,I2507,I246587,I246573,);
not I_14387 (I247131,I2514);
DFFARX1 I_14388 (I126473,I2507,I247131,I247157,);
DFFARX1 I_14389 (I247157,I2507,I247131,I247174,);
not I_14390 (I247123,I247174);
not I_14391 (I247196,I247157);
nand I_14392 (I247213,I126485,I126464);
and I_14393 (I247230,I247213,I126467);
DFFARX1 I_14394 (I247230,I2507,I247131,I247256,);
not I_14395 (I247264,I247256);
DFFARX1 I_14396 (I126476,I2507,I247131,I247290,);
and I_14397 (I247298,I247290,I126488);
nand I_14398 (I247315,I247290,I126488);
nand I_14399 (I247102,I247264,I247315);
DFFARX1 I_14400 (I126482,I2507,I247131,I247355,);
nor I_14401 (I247363,I247355,I247298);
DFFARX1 I_14402 (I247363,I2507,I247131,I247096,);
nor I_14403 (I247111,I247355,I247256);
nand I_14404 (I247408,I126470,I126467);
and I_14405 (I247425,I247408,I126479);
DFFARX1 I_14406 (I247425,I2507,I247131,I247451,);
nor I_14407 (I247099,I247451,I247355);
not I_14408 (I247473,I247451);
nor I_14409 (I247490,I247473,I247264);
nor I_14410 (I247507,I247196,I247490);
DFFARX1 I_14411 (I247507,I2507,I247131,I247114,);
nor I_14412 (I247538,I247473,I247355);
nor I_14413 (I247555,I126464,I126467);
nor I_14414 (I247105,I247555,I247538);
not I_14415 (I247586,I247555);
nand I_14416 (I247108,I247315,I247586);
DFFARX1 I_14417 (I247555,I2507,I247131,I247120,);
DFFARX1 I_14418 (I247555,I2507,I247131,I247117,);
not I_14419 (I247675,I2514);
DFFARX1 I_14420 (I86016,I2507,I247675,I247701,);
DFFARX1 I_14421 (I247701,I2507,I247675,I247718,);
not I_14422 (I247667,I247718);
not I_14423 (I247740,I247701);
nand I_14424 (I247757,I86025,I86028);
and I_14425 (I247774,I247757,I86007);
DFFARX1 I_14426 (I247774,I2507,I247675,I247800,);
not I_14427 (I247808,I247800);
DFFARX1 I_14428 (I86022,I2507,I247675,I247834,);
and I_14429 (I247842,I247834,I86010);
nand I_14430 (I247859,I247834,I86010);
nand I_14431 (I247646,I247808,I247859);
DFFARX1 I_14432 (I86004,I2507,I247675,I247899,);
nor I_14433 (I247907,I247899,I247842);
DFFARX1 I_14434 (I247907,I2507,I247675,I247640,);
nor I_14435 (I247655,I247899,I247800);
nand I_14436 (I247952,I86019,I86013);
and I_14437 (I247969,I247952,I86004);
DFFARX1 I_14438 (I247969,I2507,I247675,I247995,);
nor I_14439 (I247643,I247995,I247899);
not I_14440 (I248017,I247995);
nor I_14441 (I248034,I248017,I247808);
nor I_14442 (I248051,I247740,I248034);
DFFARX1 I_14443 (I248051,I2507,I247675,I247658,);
nor I_14444 (I248082,I248017,I247899);
nor I_14445 (I248099,I86031,I86013);
nor I_14446 (I247649,I248099,I248082);
not I_14447 (I248130,I248099);
nand I_14448 (I247652,I247859,I248130);
DFFARX1 I_14449 (I248099,I2507,I247675,I247664,);
DFFARX1 I_14450 (I248099,I2507,I247675,I247661,);
not I_14451 (I248219,I2514);
DFFARX1 I_14452 (I97318,I2507,I248219,I248245,);
DFFARX1 I_14453 (I248245,I2507,I248219,I248262,);
not I_14454 (I248211,I248262);
not I_14455 (I248284,I248245);
nand I_14456 (I248301,I97330,I97309);
and I_14457 (I248318,I248301,I97312);
DFFARX1 I_14458 (I248318,I2507,I248219,I248344,);
not I_14459 (I248352,I248344);
DFFARX1 I_14460 (I97321,I2507,I248219,I248378,);
and I_14461 (I248386,I248378,I97333);
nand I_14462 (I248403,I248378,I97333);
nand I_14463 (I248190,I248352,I248403);
DFFARX1 I_14464 (I97327,I2507,I248219,I248443,);
nor I_14465 (I248451,I248443,I248386);
DFFARX1 I_14466 (I248451,I2507,I248219,I248184,);
nor I_14467 (I248199,I248443,I248344);
nand I_14468 (I248496,I97315,I97312);
and I_14469 (I248513,I248496,I97324);
DFFARX1 I_14470 (I248513,I2507,I248219,I248539,);
nor I_14471 (I248187,I248539,I248443);
not I_14472 (I248561,I248539);
nor I_14473 (I248578,I248561,I248352);
nor I_14474 (I248595,I248284,I248578);
DFFARX1 I_14475 (I248595,I2507,I248219,I248202,);
nor I_14476 (I248626,I248561,I248443);
nor I_14477 (I248643,I97309,I97312);
nor I_14478 (I248193,I248643,I248626);
not I_14479 (I248674,I248643);
nand I_14480 (I248196,I248403,I248674);
DFFARX1 I_14481 (I248643,I2507,I248219,I248208,);
DFFARX1 I_14482 (I248643,I2507,I248219,I248205,);
not I_14483 (I248763,I2514);
DFFARX1 I_14484 (I146108,I2507,I248763,I248789,);
DFFARX1 I_14485 (I248789,I2507,I248763,I248806,);
not I_14486 (I248755,I248806);
not I_14487 (I248828,I248789);
nand I_14488 (I248845,I146120,I146099);
and I_14489 (I248862,I248845,I146102);
DFFARX1 I_14490 (I248862,I2507,I248763,I248888,);
not I_14491 (I248896,I248888);
DFFARX1 I_14492 (I146111,I2507,I248763,I248922,);
and I_14493 (I248930,I248922,I146123);
nand I_14494 (I248947,I248922,I146123);
nand I_14495 (I248734,I248896,I248947);
DFFARX1 I_14496 (I146117,I2507,I248763,I248987,);
nor I_14497 (I248995,I248987,I248930);
DFFARX1 I_14498 (I248995,I2507,I248763,I248728,);
nor I_14499 (I248743,I248987,I248888);
nand I_14500 (I249040,I146105,I146102);
and I_14501 (I249057,I249040,I146114);
DFFARX1 I_14502 (I249057,I2507,I248763,I249083,);
nor I_14503 (I248731,I249083,I248987);
not I_14504 (I249105,I249083);
nor I_14505 (I249122,I249105,I248896);
nor I_14506 (I249139,I248828,I249122);
DFFARX1 I_14507 (I249139,I2507,I248763,I248746,);
nor I_14508 (I249170,I249105,I248987);
nor I_14509 (I249187,I146099,I146102);
nor I_14510 (I248737,I249187,I249170);
not I_14511 (I249218,I249187);
nand I_14512 (I248740,I248947,I249218);
DFFARX1 I_14513 (I249187,I2507,I248763,I248752,);
DFFARX1 I_14514 (I249187,I2507,I248763,I248749,);
not I_14515 (I249307,I2514);
DFFARX1 I_14516 (I117548,I2507,I249307,I249333,);
DFFARX1 I_14517 (I249333,I2507,I249307,I249350,);
not I_14518 (I249299,I249350);
not I_14519 (I249372,I249333);
nand I_14520 (I249389,I117560,I117539);
and I_14521 (I249406,I249389,I117542);
DFFARX1 I_14522 (I249406,I2507,I249307,I249432,);
not I_14523 (I249440,I249432);
DFFARX1 I_14524 (I117551,I2507,I249307,I249466,);
and I_14525 (I249474,I249466,I117563);
nand I_14526 (I249491,I249466,I117563);
nand I_14527 (I249278,I249440,I249491);
DFFARX1 I_14528 (I117557,I2507,I249307,I249531,);
nor I_14529 (I249539,I249531,I249474);
DFFARX1 I_14530 (I249539,I2507,I249307,I249272,);
nor I_14531 (I249287,I249531,I249432);
nand I_14532 (I249584,I117545,I117542);
and I_14533 (I249601,I249584,I117554);
DFFARX1 I_14534 (I249601,I2507,I249307,I249627,);
nor I_14535 (I249275,I249627,I249531);
not I_14536 (I249649,I249627);
nor I_14537 (I249666,I249649,I249440);
nor I_14538 (I249683,I249372,I249666);
DFFARX1 I_14539 (I249683,I2507,I249307,I249290,);
nor I_14540 (I249714,I249649,I249531);
nor I_14541 (I249731,I117539,I117542);
nor I_14542 (I249281,I249731,I249714);
not I_14543 (I249762,I249731);
nand I_14544 (I249284,I249491,I249762);
DFFARX1 I_14545 (I249731,I2507,I249307,I249296,);
DFFARX1 I_14546 (I249731,I2507,I249307,I249293,);
not I_14547 (I249851,I2514);
DFFARX1 I_14548 (I205399,I2507,I249851,I249877,);
DFFARX1 I_14549 (I249877,I2507,I249851,I249894,);
not I_14550 (I249843,I249894);
not I_14551 (I249916,I249877);
nand I_14552 (I249933,I205378,I205402);
and I_14553 (I249950,I249933,I205405);
DFFARX1 I_14554 (I249950,I2507,I249851,I249976,);
not I_14555 (I249984,I249976);
DFFARX1 I_14556 (I205387,I2507,I249851,I250010,);
and I_14557 (I250018,I250010,I205393);
nand I_14558 (I250035,I250010,I205393);
nand I_14559 (I249822,I249984,I250035);
DFFARX1 I_14560 (I205381,I2507,I249851,I250075,);
nor I_14561 (I250083,I250075,I250018);
DFFARX1 I_14562 (I250083,I2507,I249851,I249816,);
nor I_14563 (I249831,I250075,I249976);
nand I_14564 (I250128,I205390,I205378);
and I_14565 (I250145,I250128,I205384);
DFFARX1 I_14566 (I250145,I2507,I249851,I250171,);
nor I_14567 (I249819,I250171,I250075);
not I_14568 (I250193,I250171);
nor I_14569 (I250210,I250193,I249984);
nor I_14570 (I250227,I249916,I250210);
DFFARX1 I_14571 (I250227,I2507,I249851,I249834,);
nor I_14572 (I250258,I250193,I250075);
nor I_14573 (I250275,I205396,I205378);
nor I_14574 (I249825,I250275,I250258);
not I_14575 (I250306,I250275);
nand I_14576 (I249828,I250035,I250306);
DFFARX1 I_14577 (I250275,I2507,I249851,I249840,);
DFFARX1 I_14578 (I250275,I2507,I249851,I249837,);
not I_14579 (I250395,I2514);
DFFARX1 I_14580 (I159793,I2507,I250395,I250421,);
DFFARX1 I_14581 (I250421,I2507,I250395,I250438,);
not I_14582 (I250387,I250438);
not I_14583 (I250460,I250421);
nand I_14584 (I250477,I159805,I159784);
and I_14585 (I250494,I250477,I159787);
DFFARX1 I_14586 (I250494,I2507,I250395,I250520,);
not I_14587 (I250528,I250520);
DFFARX1 I_14588 (I159796,I2507,I250395,I250554,);
and I_14589 (I250562,I250554,I159808);
nand I_14590 (I250579,I250554,I159808);
nand I_14591 (I250366,I250528,I250579);
DFFARX1 I_14592 (I159802,I2507,I250395,I250619,);
nor I_14593 (I250627,I250619,I250562);
DFFARX1 I_14594 (I250627,I2507,I250395,I250360,);
nor I_14595 (I250375,I250619,I250520);
nand I_14596 (I250672,I159790,I159787);
and I_14597 (I250689,I250672,I159799);
DFFARX1 I_14598 (I250689,I2507,I250395,I250715,);
nor I_14599 (I250363,I250715,I250619);
not I_14600 (I250737,I250715);
nor I_14601 (I250754,I250737,I250528);
nor I_14602 (I250771,I250460,I250754);
DFFARX1 I_14603 (I250771,I2507,I250395,I250378,);
nor I_14604 (I250802,I250737,I250619);
nor I_14605 (I250819,I159784,I159787);
nor I_14606 (I250369,I250819,I250802);
not I_14607 (I250850,I250819);
nand I_14608 (I250372,I250579,I250850);
DFFARX1 I_14609 (I250819,I2507,I250395,I250384,);
DFFARX1 I_14610 (I250819,I2507,I250395,I250381,);
not I_14611 (I250939,I2514);
DFFARX1 I_14612 (I676347,I2507,I250939,I250965,);
DFFARX1 I_14613 (I250965,I2507,I250939,I250982,);
not I_14614 (I250931,I250982);
not I_14615 (I251004,I250965);
nand I_14616 (I251021,I676344,I676341);
and I_14617 (I251038,I251021,I676329);
DFFARX1 I_14618 (I251038,I2507,I250939,I251064,);
not I_14619 (I251072,I251064);
DFFARX1 I_14620 (I676353,I2507,I250939,I251098,);
and I_14621 (I251106,I251098,I676338);
nand I_14622 (I251123,I251098,I676338);
nand I_14623 (I250910,I251072,I251123);
DFFARX1 I_14624 (I676332,I2507,I250939,I251163,);
nor I_14625 (I251171,I251163,I251106);
DFFARX1 I_14626 (I251171,I2507,I250939,I250904,);
nor I_14627 (I250919,I251163,I251064);
nand I_14628 (I251216,I676329,I676335);
and I_14629 (I251233,I251216,I676350);
DFFARX1 I_14630 (I251233,I2507,I250939,I251259,);
nor I_14631 (I250907,I251259,I251163);
not I_14632 (I251281,I251259);
nor I_14633 (I251298,I251281,I251072);
nor I_14634 (I251315,I251004,I251298);
DFFARX1 I_14635 (I251315,I2507,I250939,I250922,);
nor I_14636 (I251346,I251281,I251163);
nor I_14637 (I251363,I676332,I676335);
nor I_14638 (I250913,I251363,I251346);
not I_14639 (I251394,I251363);
nand I_14640 (I250916,I251123,I251394);
DFFARX1 I_14641 (I251363,I2507,I250939,I250928,);
DFFARX1 I_14642 (I251363,I2507,I250939,I250925,);
not I_14643 (I251483,I2514);
DFFARX1 I_14644 (I63604,I2507,I251483,I251509,);
DFFARX1 I_14645 (I251509,I2507,I251483,I251526,);
not I_14646 (I251475,I251526);
not I_14647 (I251548,I251509);
nand I_14648 (I251565,I63619,I63598);
and I_14649 (I251582,I251565,I63601);
DFFARX1 I_14650 (I251582,I2507,I251483,I251608,);
not I_14651 (I251616,I251608);
DFFARX1 I_14652 (I63607,I2507,I251483,I251642,);
and I_14653 (I251650,I251642,I63601);
nand I_14654 (I251667,I251642,I63601);
nand I_14655 (I251454,I251616,I251667);
DFFARX1 I_14656 (I63616,I2507,I251483,I251707,);
nor I_14657 (I251715,I251707,I251650);
DFFARX1 I_14658 (I251715,I2507,I251483,I251448,);
nor I_14659 (I251463,I251707,I251608);
nand I_14660 (I251760,I63598,I63613);
and I_14661 (I251777,I251760,I63610);
DFFARX1 I_14662 (I251777,I2507,I251483,I251803,);
nor I_14663 (I251451,I251803,I251707);
not I_14664 (I251825,I251803);
nor I_14665 (I251842,I251825,I251616);
nor I_14666 (I251859,I251548,I251842);
DFFARX1 I_14667 (I251859,I2507,I251483,I251466,);
nor I_14668 (I251890,I251825,I251707);
nor I_14669 (I251907,I63622,I63613);
nor I_14670 (I251457,I251907,I251890);
not I_14671 (I251938,I251907);
nand I_14672 (I251460,I251667,I251938);
DFFARX1 I_14673 (I251907,I2507,I251483,I251472,);
DFFARX1 I_14674 (I251907,I2507,I251483,I251469,);
not I_14675 (I252027,I2514);
DFFARX1 I_14676 (I289701,I2507,I252027,I252053,);
DFFARX1 I_14677 (I252053,I2507,I252027,I252070,);
not I_14678 (I252019,I252070);
not I_14679 (I252092,I252053);
nand I_14680 (I252109,I289704,I289722);
and I_14681 (I252126,I252109,I289710);
DFFARX1 I_14682 (I252126,I2507,I252027,I252152,);
not I_14683 (I252160,I252152);
DFFARX1 I_14684 (I289701,I2507,I252027,I252186,);
and I_14685 (I252194,I252186,I289719);
nand I_14686 (I252211,I252186,I289719);
nand I_14687 (I251998,I252160,I252211);
DFFARX1 I_14688 (I289713,I2507,I252027,I252251,);
nor I_14689 (I252259,I252251,I252194);
DFFARX1 I_14690 (I252259,I2507,I252027,I251992,);
nor I_14691 (I252007,I252251,I252152);
nand I_14692 (I252304,I289716,I289698);
and I_14693 (I252321,I252304,I289707);
DFFARX1 I_14694 (I252321,I2507,I252027,I252347,);
nor I_14695 (I251995,I252347,I252251);
not I_14696 (I252369,I252347);
nor I_14697 (I252386,I252369,I252160);
nor I_14698 (I252403,I252092,I252386);
DFFARX1 I_14699 (I252403,I2507,I252027,I252010,);
nor I_14700 (I252434,I252369,I252251);
nor I_14701 (I252451,I289698,I289698);
nor I_14702 (I252001,I252451,I252434);
not I_14703 (I252482,I252451);
nand I_14704 (I252004,I252211,I252482);
DFFARX1 I_14705 (I252451,I2507,I252027,I252016,);
DFFARX1 I_14706 (I252451,I2507,I252027,I252013,);
not I_14707 (I252571,I2514);
DFFARX1 I_14708 (I670567,I2507,I252571,I252597,);
DFFARX1 I_14709 (I252597,I2507,I252571,I252614,);
not I_14710 (I252563,I252614);
not I_14711 (I252636,I252597);
nand I_14712 (I252653,I670564,I670561);
and I_14713 (I252670,I252653,I670549);
DFFARX1 I_14714 (I252670,I2507,I252571,I252696,);
not I_14715 (I252704,I252696);
DFFARX1 I_14716 (I670573,I2507,I252571,I252730,);
and I_14717 (I252738,I252730,I670558);
nand I_14718 (I252755,I252730,I670558);
nand I_14719 (I252542,I252704,I252755);
DFFARX1 I_14720 (I670552,I2507,I252571,I252795,);
nor I_14721 (I252803,I252795,I252738);
DFFARX1 I_14722 (I252803,I2507,I252571,I252536,);
nor I_14723 (I252551,I252795,I252696);
nand I_14724 (I252848,I670549,I670555);
and I_14725 (I252865,I252848,I670570);
DFFARX1 I_14726 (I252865,I2507,I252571,I252891,);
nor I_14727 (I252539,I252891,I252795);
not I_14728 (I252913,I252891);
nor I_14729 (I252930,I252913,I252704);
nor I_14730 (I252947,I252636,I252930);
DFFARX1 I_14731 (I252947,I2507,I252571,I252554,);
nor I_14732 (I252978,I252913,I252795);
nor I_14733 (I252995,I670552,I670555);
nor I_14734 (I252545,I252995,I252978);
not I_14735 (I253026,I252995);
nand I_14736 (I252548,I252755,I253026);
DFFARX1 I_14737 (I252995,I2507,I252571,I252560,);
DFFARX1 I_14738 (I252995,I2507,I252571,I252557,);
not I_14739 (I253115,I2514);
DFFARX1 I_14740 (I89583,I2507,I253115,I253141,);
DFFARX1 I_14741 (I253141,I2507,I253115,I253158,);
not I_14742 (I253107,I253158);
not I_14743 (I253180,I253141);
nand I_14744 (I253197,I89595,I89574);
and I_14745 (I253214,I253197,I89577);
DFFARX1 I_14746 (I253214,I2507,I253115,I253240,);
not I_14747 (I253248,I253240);
DFFARX1 I_14748 (I89586,I2507,I253115,I253274,);
and I_14749 (I253282,I253274,I89598);
nand I_14750 (I253299,I253274,I89598);
nand I_14751 (I253086,I253248,I253299);
DFFARX1 I_14752 (I89592,I2507,I253115,I253339,);
nor I_14753 (I253347,I253339,I253282);
DFFARX1 I_14754 (I253347,I2507,I253115,I253080,);
nor I_14755 (I253095,I253339,I253240);
nand I_14756 (I253392,I89580,I89577);
and I_14757 (I253409,I253392,I89589);
DFFARX1 I_14758 (I253409,I2507,I253115,I253435,);
nor I_14759 (I253083,I253435,I253339);
not I_14760 (I253457,I253435);
nor I_14761 (I253474,I253457,I253248);
nor I_14762 (I253491,I253180,I253474);
DFFARX1 I_14763 (I253491,I2507,I253115,I253098,);
nor I_14764 (I253522,I253457,I253339);
nor I_14765 (I253539,I89574,I89577);
nor I_14766 (I253089,I253539,I253522);
not I_14767 (I253570,I253539);
nand I_14768 (I253092,I253299,I253570);
DFFARX1 I_14769 (I253539,I2507,I253115,I253104,);
DFFARX1 I_14770 (I253539,I2507,I253115,I253101,);
not I_14771 (I253659,I2514);
DFFARX1 I_14772 (I347824,I2507,I253659,I253685,);
DFFARX1 I_14773 (I253685,I2507,I253659,I253702,);
not I_14774 (I253651,I253702);
not I_14775 (I253724,I253685);
nand I_14776 (I253741,I347845,I347836);
and I_14777 (I253758,I253741,I347824);
DFFARX1 I_14778 (I253758,I2507,I253659,I253784,);
not I_14779 (I253792,I253784);
DFFARX1 I_14780 (I347830,I2507,I253659,I253818,);
and I_14781 (I253826,I253818,I347827);
nand I_14782 (I253843,I253818,I347827);
nand I_14783 (I253630,I253792,I253843);
DFFARX1 I_14784 (I347821,I2507,I253659,I253883,);
nor I_14785 (I253891,I253883,I253826);
DFFARX1 I_14786 (I253891,I2507,I253659,I253624,);
nor I_14787 (I253639,I253883,I253784);
nand I_14788 (I253936,I347821,I347833);
and I_14789 (I253953,I253936,I347842);
DFFARX1 I_14790 (I253953,I2507,I253659,I253979,);
nor I_14791 (I253627,I253979,I253883);
not I_14792 (I254001,I253979);
nor I_14793 (I254018,I254001,I253792);
nor I_14794 (I254035,I253724,I254018);
DFFARX1 I_14795 (I254035,I2507,I253659,I253642,);
nor I_14796 (I254066,I254001,I253883);
nor I_14797 (I254083,I347839,I347833);
nor I_14798 (I253633,I254083,I254066);
not I_14799 (I254114,I254083);
nand I_14800 (I253636,I253843,I254114);
DFFARX1 I_14801 (I254083,I2507,I253659,I253648,);
DFFARX1 I_14802 (I254083,I2507,I253659,I253645,);
not I_14803 (I254203,I2514);
DFFARX1 I_14804 (I225952,I2507,I254203,I254229,);
DFFARX1 I_14805 (I254229,I2507,I254203,I254246,);
not I_14806 (I254195,I254246);
not I_14807 (I254268,I254229);
nand I_14808 (I254285,I225931,I225955);
and I_14809 (I254302,I254285,I225958);
DFFARX1 I_14810 (I254302,I2507,I254203,I254328,);
not I_14811 (I254336,I254328);
DFFARX1 I_14812 (I225940,I2507,I254203,I254362,);
and I_14813 (I254370,I254362,I225946);
nand I_14814 (I254387,I254362,I225946);
nand I_14815 (I254174,I254336,I254387);
DFFARX1 I_14816 (I225934,I2507,I254203,I254427,);
nor I_14817 (I254435,I254427,I254370);
DFFARX1 I_14818 (I254435,I2507,I254203,I254168,);
nor I_14819 (I254183,I254427,I254328);
nand I_14820 (I254480,I225943,I225931);
and I_14821 (I254497,I254480,I225937);
DFFARX1 I_14822 (I254497,I2507,I254203,I254523,);
nor I_14823 (I254171,I254523,I254427);
not I_14824 (I254545,I254523);
nor I_14825 (I254562,I254545,I254336);
nor I_14826 (I254579,I254268,I254562);
DFFARX1 I_14827 (I254579,I2507,I254203,I254186,);
nor I_14828 (I254610,I254545,I254427);
nor I_14829 (I254627,I225949,I225931);
nor I_14830 (I254177,I254627,I254610);
not I_14831 (I254658,I254627);
nand I_14832 (I254180,I254387,I254658);
DFFARX1 I_14833 (I254627,I2507,I254203,I254192,);
DFFARX1 I_14834 (I254627,I2507,I254203,I254189,);
not I_14835 (I254747,I2514);
DFFARX1 I_14836 (I659400,I2507,I254747,I254773,);
DFFARX1 I_14837 (I254773,I2507,I254747,I254790,);
not I_14838 (I254739,I254790);
not I_14839 (I254812,I254773);
nand I_14840 (I254829,I659412,I659415);
and I_14841 (I254846,I254829,I659418);
DFFARX1 I_14842 (I254846,I2507,I254747,I254872,);
not I_14843 (I254880,I254872);
DFFARX1 I_14844 (I659403,I2507,I254747,I254906,);
and I_14845 (I254914,I254906,I659409);
nand I_14846 (I254931,I254906,I659409);
nand I_14847 (I254718,I254880,I254931);
DFFARX1 I_14848 (I659397,I2507,I254747,I254971,);
nor I_14849 (I254979,I254971,I254914);
DFFARX1 I_14850 (I254979,I2507,I254747,I254712,);
nor I_14851 (I254727,I254971,I254872);
nand I_14852 (I255024,I659400,I659421);
and I_14853 (I255041,I255024,I659406);
DFFARX1 I_14854 (I255041,I2507,I254747,I255067,);
nor I_14855 (I254715,I255067,I254971);
not I_14856 (I255089,I255067);
nor I_14857 (I255106,I255089,I254880);
nor I_14858 (I255123,I254812,I255106);
DFFARX1 I_14859 (I255123,I2507,I254747,I254730,);
nor I_14860 (I255154,I255089,I254971);
nor I_14861 (I255171,I659397,I659421);
nor I_14862 (I254721,I255171,I255154);
not I_14863 (I255202,I255171);
nand I_14864 (I254724,I254931,I255202);
DFFARX1 I_14865 (I255171,I2507,I254747,I254736,);
DFFARX1 I_14866 (I255171,I2507,I254747,I254733,);
not I_14867 (I255291,I2514);
DFFARX1 I_14868 (I710900,I2507,I255291,I255317,);
DFFARX1 I_14869 (I255317,I2507,I255291,I255334,);
not I_14870 (I255283,I255334);
not I_14871 (I255356,I255317);
nand I_14872 (I255373,I710876,I710897);
and I_14873 (I255390,I255373,I710894);
DFFARX1 I_14874 (I255390,I2507,I255291,I255416,);
not I_14875 (I255424,I255416);
DFFARX1 I_14876 (I710873,I2507,I255291,I255450,);
and I_14877 (I255458,I255450,I710885);
nand I_14878 (I255475,I255450,I710885);
nand I_14879 (I255262,I255424,I255475);
DFFARX1 I_14880 (I710888,I2507,I255291,I255515,);
nor I_14881 (I255523,I255515,I255458);
DFFARX1 I_14882 (I255523,I2507,I255291,I255256,);
nor I_14883 (I255271,I255515,I255416);
nand I_14884 (I255568,I710891,I710879);
and I_14885 (I255585,I255568,I710882);
DFFARX1 I_14886 (I255585,I2507,I255291,I255611,);
nor I_14887 (I255259,I255611,I255515);
not I_14888 (I255633,I255611);
nor I_14889 (I255650,I255633,I255424);
nor I_14890 (I255667,I255356,I255650);
DFFARX1 I_14891 (I255667,I2507,I255291,I255274,);
nor I_14892 (I255698,I255633,I255515);
nor I_14893 (I255715,I710873,I710879);
nor I_14894 (I255265,I255715,I255698);
not I_14895 (I255746,I255715);
nand I_14896 (I255268,I255475,I255746);
DFFARX1 I_14897 (I255715,I2507,I255291,I255280,);
DFFARX1 I_14898 (I255715,I2507,I255291,I255277,);
not I_14899 (I255835,I2514);
DFFARX1 I_14900 (I23031,I2507,I255835,I255861,);
DFFARX1 I_14901 (I255861,I2507,I255835,I255878,);
not I_14902 (I255827,I255878);
not I_14903 (I255900,I255861);
nand I_14904 (I255917,I23019,I23034);
and I_14905 (I255934,I255917,I23022);
DFFARX1 I_14906 (I255934,I2507,I255835,I255960,);
not I_14907 (I255968,I255960);
DFFARX1 I_14908 (I23043,I2507,I255835,I255994,);
and I_14909 (I256002,I255994,I23037);
nand I_14910 (I256019,I255994,I23037);
nand I_14911 (I255806,I255968,I256019);
DFFARX1 I_14912 (I23040,I2507,I255835,I256059,);
nor I_14913 (I256067,I256059,I256002);
DFFARX1 I_14914 (I256067,I2507,I255835,I255800,);
nor I_14915 (I255815,I256059,I255960);
nand I_14916 (I256112,I23019,I23022);
and I_14917 (I256129,I256112,I23025);
DFFARX1 I_14918 (I256129,I2507,I255835,I256155,);
nor I_14919 (I255803,I256155,I256059);
not I_14920 (I256177,I256155);
nor I_14921 (I256194,I256177,I255968);
nor I_14922 (I256211,I255900,I256194);
DFFARX1 I_14923 (I256211,I2507,I255835,I255818,);
nor I_14924 (I256242,I256177,I256059);
nor I_14925 (I256259,I23028,I23022);
nor I_14926 (I255809,I256259,I256242);
not I_14927 (I256290,I256259);
nand I_14928 (I255812,I256019,I256290);
DFFARX1 I_14929 (I256259,I2507,I255835,I255824,);
DFFARX1 I_14930 (I256259,I2507,I255835,I255821,);
not I_14931 (I256379,I2514);
DFFARX1 I_14932 (I188535,I2507,I256379,I256405,);
DFFARX1 I_14933 (I256405,I2507,I256379,I256422,);
not I_14934 (I256371,I256422);
not I_14935 (I256444,I256405);
nand I_14936 (I256461,I188514,I188538);
and I_14937 (I256478,I256461,I188541);
DFFARX1 I_14938 (I256478,I2507,I256379,I256504,);
not I_14939 (I256512,I256504);
DFFARX1 I_14940 (I188523,I2507,I256379,I256538,);
and I_14941 (I256546,I256538,I188529);
nand I_14942 (I256563,I256538,I188529);
nand I_14943 (I256350,I256512,I256563);
DFFARX1 I_14944 (I188517,I2507,I256379,I256603,);
nor I_14945 (I256611,I256603,I256546);
DFFARX1 I_14946 (I256611,I2507,I256379,I256344,);
nor I_14947 (I256359,I256603,I256504);
nand I_14948 (I256656,I188526,I188514);
and I_14949 (I256673,I256656,I188520);
DFFARX1 I_14950 (I256673,I2507,I256379,I256699,);
nor I_14951 (I256347,I256699,I256603);
not I_14952 (I256721,I256699);
nor I_14953 (I256738,I256721,I256512);
nor I_14954 (I256755,I256444,I256738);
DFFARX1 I_14955 (I256755,I2507,I256379,I256362,);
nor I_14956 (I256786,I256721,I256603);
nor I_14957 (I256803,I188532,I188514);
nor I_14958 (I256353,I256803,I256786);
not I_14959 (I256834,I256803);
nand I_14960 (I256356,I256563,I256834);
DFFARX1 I_14961 (I256803,I2507,I256379,I256368,);
DFFARX1 I_14962 (I256803,I2507,I256379,I256365,);
not I_14963 (I256923,I2514);
DFFARX1 I_14964 (I565472,I2507,I256923,I256949,);
DFFARX1 I_14965 (I256949,I2507,I256923,I256966,);
not I_14966 (I256915,I256966);
not I_14967 (I256988,I256949);
nand I_14968 (I257005,I565472,I565490);
and I_14969 (I257022,I257005,I565484);
DFFARX1 I_14970 (I257022,I2507,I256923,I257048,);
not I_14971 (I257056,I257048);
DFFARX1 I_14972 (I565478,I2507,I256923,I257082,);
and I_14973 (I257090,I257082,I565487);
nand I_14974 (I257107,I257082,I565487);
nand I_14975 (I256894,I257056,I257107);
DFFARX1 I_14976 (I565475,I2507,I256923,I257147,);
nor I_14977 (I257155,I257147,I257090);
DFFARX1 I_14978 (I257155,I2507,I256923,I256888,);
nor I_14979 (I256903,I257147,I257048);
nand I_14980 (I257200,I565475,I565493);
and I_14981 (I257217,I257200,I565478);
DFFARX1 I_14982 (I257217,I2507,I256923,I257243,);
nor I_14983 (I256891,I257243,I257147);
not I_14984 (I257265,I257243);
nor I_14985 (I257282,I257265,I257056);
nor I_14986 (I257299,I256988,I257282);
DFFARX1 I_14987 (I257299,I2507,I256923,I256906,);
nor I_14988 (I257330,I257265,I257147);
nor I_14989 (I257347,I565481,I565493);
nor I_14990 (I256897,I257347,I257330);
not I_14991 (I257378,I257347);
nand I_14992 (I256900,I257107,I257378);
DFFARX1 I_14993 (I257347,I2507,I256923,I256912,);
DFFARX1 I_14994 (I257347,I2507,I256923,I256909,);
not I_14995 (I257467,I2514);
DFFARX1 I_14996 (I211723,I2507,I257467,I257493,);
DFFARX1 I_14997 (I257493,I2507,I257467,I257510,);
not I_14998 (I257459,I257510);
not I_14999 (I257532,I257493);
nand I_15000 (I257549,I211702,I211726);
and I_15001 (I257566,I257549,I211729);
DFFARX1 I_15002 (I257566,I2507,I257467,I257592,);
not I_15003 (I257600,I257592);
DFFARX1 I_15004 (I211711,I2507,I257467,I257626,);
and I_15005 (I257634,I257626,I211717);
nand I_15006 (I257651,I257626,I211717);
nand I_15007 (I257438,I257600,I257651);
DFFARX1 I_15008 (I211705,I2507,I257467,I257691,);
nor I_15009 (I257699,I257691,I257634);
DFFARX1 I_15010 (I257699,I2507,I257467,I257432,);
nor I_15011 (I257447,I257691,I257592);
nand I_15012 (I257744,I211714,I211702);
and I_15013 (I257761,I257744,I211708);
DFFARX1 I_15014 (I257761,I2507,I257467,I257787,);
nor I_15015 (I257435,I257787,I257691);
not I_15016 (I257809,I257787);
nor I_15017 (I257826,I257809,I257600);
nor I_15018 (I257843,I257532,I257826);
DFFARX1 I_15019 (I257843,I2507,I257467,I257450,);
nor I_15020 (I257874,I257809,I257691);
nor I_15021 (I257891,I211720,I211702);
nor I_15022 (I257441,I257891,I257874);
not I_15023 (I257922,I257891);
nand I_15024 (I257444,I257651,I257922);
DFFARX1 I_15025 (I257891,I2507,I257467,I257456,);
DFFARX1 I_15026 (I257891,I2507,I257467,I257453,);
not I_15027 (I258011,I2514);
DFFARX1 I_15028 (I218047,I2507,I258011,I258037,);
DFFARX1 I_15029 (I258037,I2507,I258011,I258054,);
not I_15030 (I258003,I258054);
not I_15031 (I258076,I258037);
nand I_15032 (I258093,I218026,I218050);
and I_15033 (I258110,I258093,I218053);
DFFARX1 I_15034 (I258110,I2507,I258011,I258136,);
not I_15035 (I258144,I258136);
DFFARX1 I_15036 (I218035,I2507,I258011,I258170,);
and I_15037 (I258178,I258170,I218041);
nand I_15038 (I258195,I258170,I218041);
nand I_15039 (I257982,I258144,I258195);
DFFARX1 I_15040 (I218029,I2507,I258011,I258235,);
nor I_15041 (I258243,I258235,I258178);
DFFARX1 I_15042 (I258243,I2507,I258011,I257976,);
nor I_15043 (I257991,I258235,I258136);
nand I_15044 (I258288,I218038,I218026);
and I_15045 (I258305,I258288,I218032);
DFFARX1 I_15046 (I258305,I2507,I258011,I258331,);
nor I_15047 (I257979,I258331,I258235);
not I_15048 (I258353,I258331);
nor I_15049 (I258370,I258353,I258144);
nor I_15050 (I258387,I258076,I258370);
DFFARX1 I_15051 (I258387,I2507,I258011,I257994,);
nor I_15052 (I258418,I258353,I258235);
nor I_15053 (I258435,I218044,I218026);
nor I_15054 (I257985,I258435,I258418);
not I_15055 (I258466,I258435);
nand I_15056 (I257988,I258195,I258466);
DFFARX1 I_15057 (I258435,I2507,I258011,I258000,);
DFFARX1 I_15058 (I258435,I2507,I258011,I257997,);
not I_15059 (I258555,I2514);
DFFARX1 I_15060 (I339154,I2507,I258555,I258581,);
DFFARX1 I_15061 (I258581,I2507,I258555,I258598,);
not I_15062 (I258547,I258598);
not I_15063 (I258620,I258581);
nand I_15064 (I258637,I339151,I339172);
and I_15065 (I258654,I258637,I339175);
DFFARX1 I_15066 (I258654,I2507,I258555,I258680,);
not I_15067 (I258688,I258680);
DFFARX1 I_15068 (I339160,I2507,I258555,I258714,);
and I_15069 (I258722,I258714,I339163);
nand I_15070 (I258739,I258714,I339163);
nand I_15071 (I258526,I258688,I258739);
DFFARX1 I_15072 (I339166,I2507,I258555,I258779,);
nor I_15073 (I258787,I258779,I258722);
DFFARX1 I_15074 (I258787,I2507,I258555,I258520,);
nor I_15075 (I258535,I258779,I258680);
nand I_15076 (I258832,I339151,I339157);
and I_15077 (I258849,I258832,I339169);
DFFARX1 I_15078 (I258849,I2507,I258555,I258875,);
nor I_15079 (I258523,I258875,I258779);
not I_15080 (I258897,I258875);
nor I_15081 (I258914,I258897,I258688);
nor I_15082 (I258931,I258620,I258914);
DFFARX1 I_15083 (I258931,I2507,I258555,I258538,);
nor I_15084 (I258962,I258897,I258779);
nor I_15085 (I258979,I339154,I339157);
nor I_15086 (I258529,I258979,I258962);
not I_15087 (I259010,I258979);
nand I_15088 (I258532,I258739,I259010);
DFFARX1 I_15089 (I258979,I2507,I258555,I258544,);
DFFARX1 I_15090 (I258979,I2507,I258555,I258541,);
not I_15091 (I259099,I2514);
DFFARX1 I_15092 (I708520,I2507,I259099,I259125,);
DFFARX1 I_15093 (I259125,I2507,I259099,I259142,);
not I_15094 (I259091,I259142);
not I_15095 (I259164,I259125);
nand I_15096 (I259181,I708496,I708517);
and I_15097 (I259198,I259181,I708514);
DFFARX1 I_15098 (I259198,I2507,I259099,I259224,);
not I_15099 (I259232,I259224);
DFFARX1 I_15100 (I708493,I2507,I259099,I259258,);
and I_15101 (I259266,I259258,I708505);
nand I_15102 (I259283,I259258,I708505);
nand I_15103 (I259070,I259232,I259283);
DFFARX1 I_15104 (I708508,I2507,I259099,I259323,);
nor I_15105 (I259331,I259323,I259266);
DFFARX1 I_15106 (I259331,I2507,I259099,I259064,);
nor I_15107 (I259079,I259323,I259224);
nand I_15108 (I259376,I708511,I708499);
and I_15109 (I259393,I259376,I708502);
DFFARX1 I_15110 (I259393,I2507,I259099,I259419,);
nor I_15111 (I259067,I259419,I259323);
not I_15112 (I259441,I259419);
nor I_15113 (I259458,I259441,I259232);
nor I_15114 (I259475,I259164,I259458);
DFFARX1 I_15115 (I259475,I2507,I259099,I259082,);
nor I_15116 (I259506,I259441,I259323);
nor I_15117 (I259523,I708493,I708499);
nor I_15118 (I259073,I259523,I259506);
not I_15119 (I259554,I259523);
nand I_15120 (I259076,I259283,I259554);
DFFARX1 I_15121 (I259523,I2507,I259099,I259088,);
DFFARX1 I_15122 (I259523,I2507,I259099,I259085,);
not I_15123 (I259643,I2514);
DFFARX1 I_15124 (I103863,I2507,I259643,I259669,);
DFFARX1 I_15125 (I259669,I2507,I259643,I259686,);
not I_15126 (I259635,I259686);
not I_15127 (I259708,I259669);
nand I_15128 (I259725,I103875,I103854);
and I_15129 (I259742,I259725,I103857);
DFFARX1 I_15130 (I259742,I2507,I259643,I259768,);
not I_15131 (I259776,I259768);
DFFARX1 I_15132 (I103866,I2507,I259643,I259802,);
and I_15133 (I259810,I259802,I103878);
nand I_15134 (I259827,I259802,I103878);
nand I_15135 (I259614,I259776,I259827);
DFFARX1 I_15136 (I103872,I2507,I259643,I259867,);
nor I_15137 (I259875,I259867,I259810);
DFFARX1 I_15138 (I259875,I2507,I259643,I259608,);
nor I_15139 (I259623,I259867,I259768);
nand I_15140 (I259920,I103860,I103857);
and I_15141 (I259937,I259920,I103869);
DFFARX1 I_15142 (I259937,I2507,I259643,I259963,);
nor I_15143 (I259611,I259963,I259867);
not I_15144 (I259985,I259963);
nor I_15145 (I260002,I259985,I259776);
nor I_15146 (I260019,I259708,I260002);
DFFARX1 I_15147 (I260019,I2507,I259643,I259626,);
nor I_15148 (I260050,I259985,I259867);
nor I_15149 (I260067,I103854,I103857);
nor I_15150 (I259617,I260067,I260050);
not I_15151 (I260098,I260067);
nand I_15152 (I259620,I259827,I260098);
DFFARX1 I_15153 (I260067,I2507,I259643,I259632,);
DFFARX1 I_15154 (I260067,I2507,I259643,I259629,);
not I_15155 (I260187,I2514);
DFFARX1 I_15156 (I306208,I2507,I260187,I260213,);
DFFARX1 I_15157 (I260213,I2507,I260187,I260230,);
not I_15158 (I260179,I260230);
not I_15159 (I260252,I260213);
nand I_15160 (I260269,I306205,I306226);
and I_15161 (I260286,I260269,I306229);
DFFARX1 I_15162 (I260286,I2507,I260187,I260312,);
not I_15163 (I260320,I260312);
DFFARX1 I_15164 (I306214,I2507,I260187,I260346,);
and I_15165 (I260354,I260346,I306217);
nand I_15166 (I260371,I260346,I306217);
nand I_15167 (I260158,I260320,I260371);
DFFARX1 I_15168 (I306220,I2507,I260187,I260411,);
nor I_15169 (I260419,I260411,I260354);
DFFARX1 I_15170 (I260419,I2507,I260187,I260152,);
nor I_15171 (I260167,I260411,I260312);
nand I_15172 (I260464,I306205,I306211);
and I_15173 (I260481,I260464,I306223);
DFFARX1 I_15174 (I260481,I2507,I260187,I260507,);
nor I_15175 (I260155,I260507,I260411);
not I_15176 (I260529,I260507);
nor I_15177 (I260546,I260529,I260320);
nor I_15178 (I260563,I260252,I260546);
DFFARX1 I_15179 (I260563,I2507,I260187,I260170,);
nor I_15180 (I260594,I260529,I260411);
nor I_15181 (I260611,I306208,I306211);
nor I_15182 (I260161,I260611,I260594);
not I_15183 (I260642,I260611);
nand I_15184 (I260164,I260371,I260642);
DFFARX1 I_15185 (I260611,I2507,I260187,I260176,);
DFFARX1 I_15186 (I260611,I2507,I260187,I260173,);
not I_15187 (I260731,I2514);
DFFARX1 I_15188 (I721610,I2507,I260731,I260757,);
DFFARX1 I_15189 (I260757,I2507,I260731,I260774,);
not I_15190 (I260723,I260774);
not I_15191 (I260796,I260757);
nand I_15192 (I260813,I721586,I721607);
and I_15193 (I260830,I260813,I721604);
DFFARX1 I_15194 (I260830,I2507,I260731,I260856,);
not I_15195 (I260864,I260856);
DFFARX1 I_15196 (I721583,I2507,I260731,I260890,);
and I_15197 (I260898,I260890,I721595);
nand I_15198 (I260915,I260890,I721595);
nand I_15199 (I260702,I260864,I260915);
DFFARX1 I_15200 (I721598,I2507,I260731,I260955,);
nor I_15201 (I260963,I260955,I260898);
DFFARX1 I_15202 (I260963,I2507,I260731,I260696,);
nor I_15203 (I260711,I260955,I260856);
nand I_15204 (I261008,I721601,I721589);
and I_15205 (I261025,I261008,I721592);
DFFARX1 I_15206 (I261025,I2507,I260731,I261051,);
nor I_15207 (I260699,I261051,I260955);
not I_15208 (I261073,I261051);
nor I_15209 (I261090,I261073,I260864);
nor I_15210 (I261107,I260796,I261090);
DFFARX1 I_15211 (I261107,I2507,I260731,I260714,);
nor I_15212 (I261138,I261073,I260955);
nor I_15213 (I261155,I721583,I721589);
nor I_15214 (I260705,I261155,I261138);
not I_15215 (I261186,I261155);
nand I_15216 (I260708,I260915,I261186);
DFFARX1 I_15217 (I261155,I2507,I260731,I260720,);
DFFARX1 I_15218 (I261155,I2507,I260731,I260717,);
not I_15219 (I261275,I2514);
DFFARX1 I_15220 (I558179,I2507,I261275,I261301,);
DFFARX1 I_15221 (I261301,I2507,I261275,I261318,);
not I_15222 (I261267,I261318);
not I_15223 (I261340,I261301);
nand I_15224 (I261357,I558179,I558197);
and I_15225 (I261374,I261357,I558191);
DFFARX1 I_15226 (I261374,I2507,I261275,I261400,);
not I_15227 (I261408,I261400);
DFFARX1 I_15228 (I558185,I2507,I261275,I261434,);
and I_15229 (I261442,I261434,I558194);
nand I_15230 (I261459,I261434,I558194);
nand I_15231 (I261246,I261408,I261459);
DFFARX1 I_15232 (I558182,I2507,I261275,I261499,);
nor I_15233 (I261507,I261499,I261442);
DFFARX1 I_15234 (I261507,I2507,I261275,I261240,);
nor I_15235 (I261255,I261499,I261400);
nand I_15236 (I261552,I558182,I558200);
and I_15237 (I261569,I261552,I558185);
DFFARX1 I_15238 (I261569,I2507,I261275,I261595,);
nor I_15239 (I261243,I261595,I261499);
not I_15240 (I261617,I261595);
nor I_15241 (I261634,I261617,I261408);
nor I_15242 (I261651,I261340,I261634);
DFFARX1 I_15243 (I261651,I2507,I261275,I261258,);
nor I_15244 (I261682,I261617,I261499);
nor I_15245 (I261699,I558188,I558200);
nor I_15246 (I261249,I261699,I261682);
not I_15247 (I261730,I261699);
nand I_15248 (I261252,I261459,I261730);
DFFARX1 I_15249 (I261699,I2507,I261275,I261264,);
DFFARX1 I_15250 (I261699,I2507,I261275,I261261,);
not I_15251 (I261819,I2514);
DFFARX1 I_15252 (I532566,I2507,I261819,I261845,);
DFFARX1 I_15253 (I261845,I2507,I261819,I261862,);
not I_15254 (I261811,I261862);
not I_15255 (I261884,I261845);
nand I_15256 (I261901,I532581,I532569);
and I_15257 (I261918,I261901,I532560);
DFFARX1 I_15258 (I261918,I2507,I261819,I261944,);
not I_15259 (I261952,I261944);
DFFARX1 I_15260 (I532572,I2507,I261819,I261978,);
and I_15261 (I261986,I261978,I532563);
nand I_15262 (I262003,I261978,I532563);
nand I_15263 (I261790,I261952,I262003);
DFFARX1 I_15264 (I532578,I2507,I261819,I262043,);
nor I_15265 (I262051,I262043,I261986);
DFFARX1 I_15266 (I262051,I2507,I261819,I261784,);
nor I_15267 (I261799,I262043,I261944);
nand I_15268 (I262096,I532587,I532575);
and I_15269 (I262113,I262096,I532584);
DFFARX1 I_15270 (I262113,I2507,I261819,I262139,);
nor I_15271 (I261787,I262139,I262043);
not I_15272 (I262161,I262139);
nor I_15273 (I262178,I262161,I261952);
nor I_15274 (I262195,I261884,I262178);
DFFARX1 I_15275 (I262195,I2507,I261819,I261802,);
nor I_15276 (I262226,I262161,I262043);
nor I_15277 (I262243,I532560,I532575);
nor I_15278 (I261793,I262243,I262226);
not I_15279 (I262274,I262243);
nand I_15280 (I261796,I262003,I262274);
DFFARX1 I_15281 (I262243,I2507,I261819,I261808,);
DFFARX1 I_15282 (I262243,I2507,I261819,I261805,);
not I_15283 (I262363,I2514);
DFFARX1 I_15284 (I19869,I2507,I262363,I262389,);
DFFARX1 I_15285 (I262389,I2507,I262363,I262406,);
not I_15286 (I262355,I262406);
not I_15287 (I262428,I262389);
nand I_15288 (I262445,I19857,I19872);
and I_15289 (I262462,I262445,I19860);
DFFARX1 I_15290 (I262462,I2507,I262363,I262488,);
not I_15291 (I262496,I262488);
DFFARX1 I_15292 (I19881,I2507,I262363,I262522,);
and I_15293 (I262530,I262522,I19875);
nand I_15294 (I262547,I262522,I19875);
nand I_15295 (I262334,I262496,I262547);
DFFARX1 I_15296 (I19878,I2507,I262363,I262587,);
nor I_15297 (I262595,I262587,I262530);
DFFARX1 I_15298 (I262595,I2507,I262363,I262328,);
nor I_15299 (I262343,I262587,I262488);
nand I_15300 (I262640,I19857,I19860);
and I_15301 (I262657,I262640,I19863);
DFFARX1 I_15302 (I262657,I2507,I262363,I262683,);
nor I_15303 (I262331,I262683,I262587);
not I_15304 (I262705,I262683);
nor I_15305 (I262722,I262705,I262496);
nor I_15306 (I262739,I262428,I262722);
DFFARX1 I_15307 (I262739,I2507,I262363,I262346,);
nor I_15308 (I262770,I262705,I262587);
nor I_15309 (I262787,I19866,I19860);
nor I_15310 (I262337,I262787,I262770);
not I_15311 (I262818,I262787);
nand I_15312 (I262340,I262547,I262818);
DFFARX1 I_15313 (I262787,I2507,I262363,I262352,);
DFFARX1 I_15314 (I262787,I2507,I262363,I262349,);
not I_15315 (I262907,I2514);
DFFARX1 I_15316 (I311988,I2507,I262907,I262933,);
DFFARX1 I_15317 (I262933,I2507,I262907,I262950,);
not I_15318 (I262899,I262950);
not I_15319 (I262972,I262933);
nand I_15320 (I262989,I311985,I312006);
and I_15321 (I263006,I262989,I312009);
DFFARX1 I_15322 (I263006,I2507,I262907,I263032,);
not I_15323 (I263040,I263032);
DFFARX1 I_15324 (I311994,I2507,I262907,I263066,);
and I_15325 (I263074,I263066,I311997);
nand I_15326 (I263091,I263066,I311997);
nand I_15327 (I262878,I263040,I263091);
DFFARX1 I_15328 (I312000,I2507,I262907,I263131,);
nor I_15329 (I263139,I263131,I263074);
DFFARX1 I_15330 (I263139,I2507,I262907,I262872,);
nor I_15331 (I262887,I263131,I263032);
nand I_15332 (I263184,I311985,I311991);
and I_15333 (I263201,I263184,I312003);
DFFARX1 I_15334 (I263201,I2507,I262907,I263227,);
nor I_15335 (I262875,I263227,I263131);
not I_15336 (I263249,I263227);
nor I_15337 (I263266,I263249,I263040);
nor I_15338 (I263283,I262972,I263266);
DFFARX1 I_15339 (I263283,I2507,I262907,I262890,);
nor I_15340 (I263314,I263249,I263131);
nor I_15341 (I263331,I311988,I311991);
nor I_15342 (I262881,I263331,I263314);
not I_15343 (I263362,I263331);
nand I_15344 (I262884,I263091,I263362);
DFFARX1 I_15345 (I263331,I2507,I262907,I262896,);
DFFARX1 I_15346 (I263331,I2507,I262907,I262893,);
not I_15347 (I263451,I2514);
DFFARX1 I_15348 (I66766,I2507,I263451,I263477,);
DFFARX1 I_15349 (I263477,I2507,I263451,I263494,);
not I_15350 (I263443,I263494);
not I_15351 (I263516,I263477);
nand I_15352 (I263533,I66781,I66760);
and I_15353 (I263550,I263533,I66763);
DFFARX1 I_15354 (I263550,I2507,I263451,I263576,);
not I_15355 (I263584,I263576);
DFFARX1 I_15356 (I66769,I2507,I263451,I263610,);
and I_15357 (I263618,I263610,I66763);
nand I_15358 (I263635,I263610,I66763);
nand I_15359 (I263422,I263584,I263635);
DFFARX1 I_15360 (I66778,I2507,I263451,I263675,);
nor I_15361 (I263683,I263675,I263618);
DFFARX1 I_15362 (I263683,I2507,I263451,I263416,);
nor I_15363 (I263431,I263675,I263576);
nand I_15364 (I263728,I66760,I66775);
and I_15365 (I263745,I263728,I66772);
DFFARX1 I_15366 (I263745,I2507,I263451,I263771,);
nor I_15367 (I263419,I263771,I263675);
not I_15368 (I263793,I263771);
nor I_15369 (I263810,I263793,I263584);
nor I_15370 (I263827,I263516,I263810);
DFFARX1 I_15371 (I263827,I2507,I263451,I263434,);
nor I_15372 (I263858,I263793,I263675);
nor I_15373 (I263875,I66784,I66775);
nor I_15374 (I263425,I263875,I263858);
not I_15375 (I263906,I263875);
nand I_15376 (I263428,I263635,I263906);
DFFARX1 I_15377 (I263875,I2507,I263451,I263440,);
DFFARX1 I_15378 (I263875,I2507,I263451,I263437,);
not I_15379 (I263995,I2514);
DFFARX1 I_15380 (I157413,I2507,I263995,I264021,);
DFFARX1 I_15381 (I264021,I2507,I263995,I264038,);
not I_15382 (I263987,I264038);
not I_15383 (I264060,I264021);
nand I_15384 (I264077,I157425,I157404);
and I_15385 (I264094,I264077,I157407);
DFFARX1 I_15386 (I264094,I2507,I263995,I264120,);
not I_15387 (I264128,I264120);
DFFARX1 I_15388 (I157416,I2507,I263995,I264154,);
and I_15389 (I264162,I264154,I157428);
nand I_15390 (I264179,I264154,I157428);
nand I_15391 (I263966,I264128,I264179);
DFFARX1 I_15392 (I157422,I2507,I263995,I264219,);
nor I_15393 (I264227,I264219,I264162);
DFFARX1 I_15394 (I264227,I2507,I263995,I263960,);
nor I_15395 (I263975,I264219,I264120);
nand I_15396 (I264272,I157410,I157407);
and I_15397 (I264289,I264272,I157419);
DFFARX1 I_15398 (I264289,I2507,I263995,I264315,);
nor I_15399 (I263963,I264315,I264219);
not I_15400 (I264337,I264315);
nor I_15401 (I264354,I264337,I264128);
nor I_15402 (I264371,I264060,I264354);
DFFARX1 I_15403 (I264371,I2507,I263995,I263978,);
nor I_15404 (I264402,I264337,I264219);
nor I_15405 (I264419,I157404,I157407);
nor I_15406 (I263969,I264419,I264402);
not I_15407 (I264450,I264419);
nand I_15408 (I263972,I264179,I264450);
DFFARX1 I_15409 (I264419,I2507,I263995,I263984,);
DFFARX1 I_15410 (I264419,I2507,I263995,I263981,);
not I_15411 (I264539,I2514);
DFFARX1 I_15412 (I54645,I2507,I264539,I264565,);
DFFARX1 I_15413 (I264565,I2507,I264539,I264582,);
not I_15414 (I264531,I264582);
not I_15415 (I264604,I264565);
nand I_15416 (I264621,I54660,I54639);
and I_15417 (I264638,I264621,I54642);
DFFARX1 I_15418 (I264638,I2507,I264539,I264664,);
not I_15419 (I264672,I264664);
DFFARX1 I_15420 (I54648,I2507,I264539,I264698,);
and I_15421 (I264706,I264698,I54642);
nand I_15422 (I264723,I264698,I54642);
nand I_15423 (I264510,I264672,I264723);
DFFARX1 I_15424 (I54657,I2507,I264539,I264763,);
nor I_15425 (I264771,I264763,I264706);
DFFARX1 I_15426 (I264771,I2507,I264539,I264504,);
nor I_15427 (I264519,I264763,I264664);
nand I_15428 (I264816,I54639,I54654);
and I_15429 (I264833,I264816,I54651);
DFFARX1 I_15430 (I264833,I2507,I264539,I264859,);
nor I_15431 (I264507,I264859,I264763);
not I_15432 (I264881,I264859);
nor I_15433 (I264898,I264881,I264672);
nor I_15434 (I264915,I264604,I264898);
DFFARX1 I_15435 (I264915,I2507,I264539,I264522,);
nor I_15436 (I264946,I264881,I264763);
nor I_15437 (I264963,I54663,I54654);
nor I_15438 (I264513,I264963,I264946);
not I_15439 (I264994,I264963);
nand I_15440 (I264516,I264723,I264994);
DFFARX1 I_15441 (I264963,I2507,I264539,I264528,);
DFFARX1 I_15442 (I264963,I2507,I264539,I264525,);
not I_15443 (I265083,I2514);
DFFARX1 I_15444 (I678659,I2507,I265083,I265109,);
DFFARX1 I_15445 (I265109,I2507,I265083,I265126,);
not I_15446 (I265075,I265126);
not I_15447 (I265148,I265109);
nand I_15448 (I265165,I678656,I678653);
and I_15449 (I265182,I265165,I678641);
DFFARX1 I_15450 (I265182,I2507,I265083,I265208,);
not I_15451 (I265216,I265208);
DFFARX1 I_15452 (I678665,I2507,I265083,I265242,);
and I_15453 (I265250,I265242,I678650);
nand I_15454 (I265267,I265242,I678650);
nand I_15455 (I265054,I265216,I265267);
DFFARX1 I_15456 (I678644,I2507,I265083,I265307,);
nor I_15457 (I265315,I265307,I265250);
DFFARX1 I_15458 (I265315,I2507,I265083,I265048,);
nor I_15459 (I265063,I265307,I265208);
nand I_15460 (I265360,I678641,I678647);
and I_15461 (I265377,I265360,I678662);
DFFARX1 I_15462 (I265377,I2507,I265083,I265403,);
nor I_15463 (I265051,I265403,I265307);
not I_15464 (I265425,I265403);
nor I_15465 (I265442,I265425,I265216);
nor I_15466 (I265459,I265148,I265442);
DFFARX1 I_15467 (I265459,I2507,I265083,I265066,);
nor I_15468 (I265490,I265425,I265307);
nor I_15469 (I265507,I678644,I678647);
nor I_15470 (I265057,I265507,I265490);
not I_15471 (I265538,I265507);
nand I_15472 (I265060,I265267,I265538);
DFFARX1 I_15473 (I265507,I2507,I265083,I265072,);
DFFARX1 I_15474 (I265507,I2507,I265083,I265069,);
not I_15475 (I265627,I2514);
DFFARX1 I_15476 (I281966,I2507,I265627,I265653,);
DFFARX1 I_15477 (I265653,I2507,I265627,I265670,);
not I_15478 (I265619,I265670);
not I_15479 (I265692,I265653);
nand I_15480 (I265709,I281969,I281987);
and I_15481 (I265726,I265709,I281975);
DFFARX1 I_15482 (I265726,I2507,I265627,I265752,);
not I_15483 (I265760,I265752);
DFFARX1 I_15484 (I281966,I2507,I265627,I265786,);
and I_15485 (I265794,I265786,I281984);
nand I_15486 (I265811,I265786,I281984);
nand I_15487 (I265598,I265760,I265811);
DFFARX1 I_15488 (I281978,I2507,I265627,I265851,);
nor I_15489 (I265859,I265851,I265794);
DFFARX1 I_15490 (I265859,I2507,I265627,I265592,);
nor I_15491 (I265607,I265851,I265752);
nand I_15492 (I265904,I281981,I281963);
and I_15493 (I265921,I265904,I281972);
DFFARX1 I_15494 (I265921,I2507,I265627,I265947,);
nor I_15495 (I265595,I265947,I265851);
not I_15496 (I265969,I265947);
nor I_15497 (I265986,I265969,I265760);
nor I_15498 (I266003,I265692,I265986);
DFFARX1 I_15499 (I266003,I2507,I265627,I265610,);
nor I_15500 (I266034,I265969,I265851);
nor I_15501 (I266051,I281963,I281963);
nor I_15502 (I265601,I266051,I266034);
not I_15503 (I266082,I266051);
nand I_15504 (I265604,I265811,I266082);
DFFARX1 I_15505 (I266051,I2507,I265627,I265616,);
DFFARX1 I_15506 (I266051,I2507,I265627,I265613,);
not I_15507 (I266171,I2514);
DFFARX1 I_15508 (I321236,I2507,I266171,I266197,);
DFFARX1 I_15509 (I266197,I2507,I266171,I266214,);
not I_15510 (I266163,I266214);
not I_15511 (I266236,I266197);
nand I_15512 (I266253,I321233,I321254);
and I_15513 (I266270,I266253,I321257);
DFFARX1 I_15514 (I266270,I2507,I266171,I266296,);
not I_15515 (I266304,I266296);
DFFARX1 I_15516 (I321242,I2507,I266171,I266330,);
and I_15517 (I266338,I266330,I321245);
nand I_15518 (I266355,I266330,I321245);
nand I_15519 (I266142,I266304,I266355);
DFFARX1 I_15520 (I321248,I2507,I266171,I266395,);
nor I_15521 (I266403,I266395,I266338);
DFFARX1 I_15522 (I266403,I2507,I266171,I266136,);
nor I_15523 (I266151,I266395,I266296);
nand I_15524 (I266448,I321233,I321239);
and I_15525 (I266465,I266448,I321251);
DFFARX1 I_15526 (I266465,I2507,I266171,I266491,);
nor I_15527 (I266139,I266491,I266395);
not I_15528 (I266513,I266491);
nor I_15529 (I266530,I266513,I266304);
nor I_15530 (I266547,I266236,I266530);
DFFARX1 I_15531 (I266547,I2507,I266171,I266154,);
nor I_15532 (I266578,I266513,I266395);
nor I_15533 (I266595,I321236,I321239);
nor I_15534 (I266145,I266595,I266578);
not I_15535 (I266626,I266595);
nand I_15536 (I266148,I266355,I266626);
DFFARX1 I_15537 (I266595,I2507,I266171,I266160,);
DFFARX1 I_15538 (I266595,I2507,I266171,I266157,);
not I_15539 (I266715,I2514);
DFFARX1 I_15540 (I353026,I2507,I266715,I266741,);
DFFARX1 I_15541 (I266741,I2507,I266715,I266758,);
not I_15542 (I266707,I266758);
not I_15543 (I266780,I266741);
nand I_15544 (I266797,I353047,I353038);
and I_15545 (I266814,I266797,I353026);
DFFARX1 I_15546 (I266814,I2507,I266715,I266840,);
not I_15547 (I266848,I266840);
DFFARX1 I_15548 (I353032,I2507,I266715,I266874,);
and I_15549 (I266882,I266874,I353029);
nand I_15550 (I266899,I266874,I353029);
nand I_15551 (I266686,I266848,I266899);
DFFARX1 I_15552 (I353023,I2507,I266715,I266939,);
nor I_15553 (I266947,I266939,I266882);
DFFARX1 I_15554 (I266947,I2507,I266715,I266680,);
nor I_15555 (I266695,I266939,I266840);
nand I_15556 (I266992,I353023,I353035);
and I_15557 (I267009,I266992,I353044);
DFFARX1 I_15558 (I267009,I2507,I266715,I267035,);
nor I_15559 (I266683,I267035,I266939);
not I_15560 (I267057,I267035);
nor I_15561 (I267074,I267057,I266848);
nor I_15562 (I267091,I266780,I267074);
DFFARX1 I_15563 (I267091,I2507,I266715,I266698,);
nor I_15564 (I267122,I267057,I266939);
nor I_15565 (I267139,I353041,I353035);
nor I_15566 (I266689,I267139,I267122);
not I_15567 (I267170,I267139);
nand I_15568 (I266692,I266899,I267170);
DFFARX1 I_15569 (I267139,I2507,I266715,I266704,);
DFFARX1 I_15570 (I267139,I2507,I266715,I266701,);
not I_15571 (I267259,I2514);
DFFARX1 I_15572 (I458690,I2507,I267259,I267285,);
DFFARX1 I_15573 (I267285,I2507,I267259,I267302,);
not I_15574 (I267251,I267302);
not I_15575 (I267324,I267285);
nand I_15576 (I267341,I458684,I458681);
and I_15577 (I267358,I267341,I458696);
DFFARX1 I_15578 (I267358,I2507,I267259,I267384,);
not I_15579 (I267392,I267384);
DFFARX1 I_15580 (I458684,I2507,I267259,I267418,);
and I_15581 (I267426,I267418,I458678);
nand I_15582 (I267443,I267418,I458678);
nand I_15583 (I267230,I267392,I267443);
DFFARX1 I_15584 (I458678,I2507,I267259,I267483,);
nor I_15585 (I267491,I267483,I267426);
DFFARX1 I_15586 (I267491,I2507,I267259,I267224,);
nor I_15587 (I267239,I267483,I267384);
nand I_15588 (I267536,I458693,I458687);
and I_15589 (I267553,I267536,I458681);
DFFARX1 I_15590 (I267553,I2507,I267259,I267579,);
nor I_15591 (I267227,I267579,I267483);
not I_15592 (I267601,I267579);
nor I_15593 (I267618,I267601,I267392);
nor I_15594 (I267635,I267324,I267618);
DFFARX1 I_15595 (I267635,I2507,I267259,I267242,);
nor I_15596 (I267666,I267601,I267483);
nor I_15597 (I267683,I458699,I458687);
nor I_15598 (I267233,I267683,I267666);
not I_15599 (I267714,I267683);
nand I_15600 (I267236,I267443,I267714);
DFFARX1 I_15601 (I267683,I2507,I267259,I267248,);
DFFARX1 I_15602 (I267683,I2507,I267259,I267245,);
not I_15603 (I267803,I2514);
DFFARX1 I_15604 (I576304,I2507,I267803,I267829,);
DFFARX1 I_15605 (I267829,I2507,I267803,I267846,);
not I_15606 (I267795,I267846);
not I_15607 (I267868,I267829);
nand I_15608 (I267885,I576316,I576304);
and I_15609 (I267902,I267885,I576307);
DFFARX1 I_15610 (I267902,I2507,I267803,I267928,);
not I_15611 (I267936,I267928);
DFFARX1 I_15612 (I576325,I2507,I267803,I267962,);
and I_15613 (I267970,I267962,I576301);
nand I_15614 (I267987,I267962,I576301);
nand I_15615 (I267774,I267936,I267987);
DFFARX1 I_15616 (I576319,I2507,I267803,I268027,);
nor I_15617 (I268035,I268027,I267970);
DFFARX1 I_15618 (I268035,I2507,I267803,I267768,);
nor I_15619 (I267783,I268027,I267928);
nand I_15620 (I268080,I576313,I576310);
and I_15621 (I268097,I268080,I576322);
DFFARX1 I_15622 (I268097,I2507,I267803,I268123,);
nor I_15623 (I267771,I268123,I268027);
not I_15624 (I268145,I268123);
nor I_15625 (I268162,I268145,I267936);
nor I_15626 (I268179,I267868,I268162);
DFFARX1 I_15627 (I268179,I2507,I267803,I267786,);
nor I_15628 (I268210,I268145,I268027);
nor I_15629 (I268227,I576301,I576310);
nor I_15630 (I267777,I268227,I268210);
not I_15631 (I268258,I268227);
nand I_15632 (I267780,I267987,I268258);
DFFARX1 I_15633 (I268227,I2507,I267803,I267792,);
DFFARX1 I_15634 (I268227,I2507,I267803,I267789,);
not I_15635 (I268347,I2514);
DFFARX1 I_15636 (I46213,I2507,I268347,I268373,);
DFFARX1 I_15637 (I268373,I2507,I268347,I268390,);
not I_15638 (I268339,I268390);
not I_15639 (I268412,I268373);
nand I_15640 (I268429,I46228,I46207);
and I_15641 (I268446,I268429,I46210);
DFFARX1 I_15642 (I268446,I2507,I268347,I268472,);
not I_15643 (I268480,I268472);
DFFARX1 I_15644 (I46216,I2507,I268347,I268506,);
and I_15645 (I268514,I268506,I46210);
nand I_15646 (I268531,I268506,I46210);
nand I_15647 (I268318,I268480,I268531);
DFFARX1 I_15648 (I46225,I2507,I268347,I268571,);
nor I_15649 (I268579,I268571,I268514);
DFFARX1 I_15650 (I268579,I2507,I268347,I268312,);
nor I_15651 (I268327,I268571,I268472);
nand I_15652 (I268624,I46207,I46222);
and I_15653 (I268641,I268624,I46219);
DFFARX1 I_15654 (I268641,I2507,I268347,I268667,);
nor I_15655 (I268315,I268667,I268571);
not I_15656 (I268689,I268667);
nor I_15657 (I268706,I268689,I268480);
nor I_15658 (I268723,I268412,I268706);
DFFARX1 I_15659 (I268723,I2507,I268347,I268330,);
nor I_15660 (I268754,I268689,I268571);
nor I_15661 (I268771,I46231,I46222);
nor I_15662 (I268321,I268771,I268754);
not I_15663 (I268802,I268771);
nand I_15664 (I268324,I268531,I268802);
DFFARX1 I_15665 (I268771,I2507,I268347,I268336,);
DFFARX1 I_15666 (I268771,I2507,I268347,I268333,);
not I_15667 (I268891,I2514);
DFFARX1 I_15668 (I520938,I2507,I268891,I268917,);
DFFARX1 I_15669 (I268917,I2507,I268891,I268934,);
not I_15670 (I268883,I268934);
not I_15671 (I268956,I268917);
nand I_15672 (I268973,I520953,I520941);
and I_15673 (I268990,I268973,I520932);
DFFARX1 I_15674 (I268990,I2507,I268891,I269016,);
not I_15675 (I269024,I269016);
DFFARX1 I_15676 (I520944,I2507,I268891,I269050,);
and I_15677 (I269058,I269050,I520935);
nand I_15678 (I269075,I269050,I520935);
nand I_15679 (I268862,I269024,I269075);
DFFARX1 I_15680 (I520950,I2507,I268891,I269115,);
nor I_15681 (I269123,I269115,I269058);
DFFARX1 I_15682 (I269123,I2507,I268891,I268856,);
nor I_15683 (I268871,I269115,I269016);
nand I_15684 (I269168,I520959,I520947);
and I_15685 (I269185,I269168,I520956);
DFFARX1 I_15686 (I269185,I2507,I268891,I269211,);
nor I_15687 (I268859,I269211,I269115);
not I_15688 (I269233,I269211);
nor I_15689 (I269250,I269233,I269024);
nor I_15690 (I269267,I268956,I269250);
DFFARX1 I_15691 (I269267,I2507,I268891,I268874,);
nor I_15692 (I269298,I269233,I269115);
nor I_15693 (I269315,I520932,I520947);
nor I_15694 (I268865,I269315,I269298);
not I_15695 (I269346,I269315);
nand I_15696 (I268868,I269075,I269346);
DFFARX1 I_15697 (I269315,I2507,I268891,I268880,);
DFFARX1 I_15698 (I269315,I2507,I268891,I268877,);
not I_15699 (I269435,I2514);
DFFARX1 I_15700 (I207507,I2507,I269435,I269461,);
DFFARX1 I_15701 (I269461,I2507,I269435,I269478,);
not I_15702 (I269427,I269478);
not I_15703 (I269500,I269461);
nand I_15704 (I269517,I207486,I207510);
and I_15705 (I269534,I269517,I207513);
DFFARX1 I_15706 (I269534,I2507,I269435,I269560,);
not I_15707 (I269568,I269560);
DFFARX1 I_15708 (I207495,I2507,I269435,I269594,);
and I_15709 (I269602,I269594,I207501);
nand I_15710 (I269619,I269594,I207501);
nand I_15711 (I269406,I269568,I269619);
DFFARX1 I_15712 (I207489,I2507,I269435,I269659,);
nor I_15713 (I269667,I269659,I269602);
DFFARX1 I_15714 (I269667,I2507,I269435,I269400,);
nor I_15715 (I269415,I269659,I269560);
nand I_15716 (I269712,I207498,I207486);
and I_15717 (I269729,I269712,I207492);
DFFARX1 I_15718 (I269729,I2507,I269435,I269755,);
nor I_15719 (I269403,I269755,I269659);
not I_15720 (I269777,I269755);
nor I_15721 (I269794,I269777,I269568);
nor I_15722 (I269811,I269500,I269794);
DFFARX1 I_15723 (I269811,I2507,I269435,I269418,);
nor I_15724 (I269842,I269777,I269659);
nor I_15725 (I269859,I207504,I207486);
nor I_15726 (I269409,I269859,I269842);
not I_15727 (I269890,I269859);
nand I_15728 (I269412,I269619,I269890);
DFFARX1 I_15729 (I269859,I2507,I269435,I269424,);
DFFARX1 I_15730 (I269859,I2507,I269435,I269421,);
not I_15731 (I269979,I2514);
DFFARX1 I_15732 (I521584,I2507,I269979,I270005,);
DFFARX1 I_15733 (I270005,I2507,I269979,I270022,);
not I_15734 (I269971,I270022);
not I_15735 (I270044,I270005);
nand I_15736 (I270061,I521599,I521587);
and I_15737 (I270078,I270061,I521578);
DFFARX1 I_15738 (I270078,I2507,I269979,I270104,);
not I_15739 (I270112,I270104);
DFFARX1 I_15740 (I521590,I2507,I269979,I270138,);
and I_15741 (I270146,I270138,I521581);
nand I_15742 (I270163,I270138,I521581);
nand I_15743 (I269950,I270112,I270163);
DFFARX1 I_15744 (I521596,I2507,I269979,I270203,);
nor I_15745 (I270211,I270203,I270146);
DFFARX1 I_15746 (I270211,I2507,I269979,I269944,);
nor I_15747 (I269959,I270203,I270104);
nand I_15748 (I270256,I521605,I521593);
and I_15749 (I270273,I270256,I521602);
DFFARX1 I_15750 (I270273,I2507,I269979,I270299,);
nor I_15751 (I269947,I270299,I270203);
not I_15752 (I270321,I270299);
nor I_15753 (I270338,I270321,I270112);
nor I_15754 (I270355,I270044,I270338);
DFFARX1 I_15755 (I270355,I2507,I269979,I269962,);
nor I_15756 (I270386,I270321,I270203);
nor I_15757 (I270403,I521578,I521593);
nor I_15758 (I269953,I270403,I270386);
not I_15759 (I270434,I270403);
nand I_15760 (I269956,I270163,I270434);
DFFARX1 I_15761 (I270403,I2507,I269979,I269968,);
DFFARX1 I_15762 (I270403,I2507,I269979,I269965,);
not I_15763 (I270523,I2514);
DFFARX1 I_15764 (I428651,I2507,I270523,I270549,);
DFFARX1 I_15765 (I270549,I2507,I270523,I270566,);
not I_15766 (I270515,I270566);
not I_15767 (I270588,I270549);
nand I_15768 (I270605,I428645,I428642);
and I_15769 (I270622,I270605,I428657);
DFFARX1 I_15770 (I270622,I2507,I270523,I270648,);
not I_15771 (I270656,I270648);
DFFARX1 I_15772 (I428645,I2507,I270523,I270682,);
and I_15773 (I270690,I270682,I428639);
nand I_15774 (I270707,I270682,I428639);
nand I_15775 (I270494,I270656,I270707);
DFFARX1 I_15776 (I428639,I2507,I270523,I270747,);
nor I_15777 (I270755,I270747,I270690);
DFFARX1 I_15778 (I270755,I2507,I270523,I270488,);
nor I_15779 (I270503,I270747,I270648);
nand I_15780 (I270800,I428654,I428648);
and I_15781 (I270817,I270800,I428642);
DFFARX1 I_15782 (I270817,I2507,I270523,I270843,);
nor I_15783 (I270491,I270843,I270747);
not I_15784 (I270865,I270843);
nor I_15785 (I270882,I270865,I270656);
nor I_15786 (I270899,I270588,I270882);
DFFARX1 I_15787 (I270899,I2507,I270523,I270506,);
nor I_15788 (I270930,I270865,I270747);
nor I_15789 (I270947,I428660,I428648);
nor I_15790 (I270497,I270947,I270930);
not I_15791 (I270978,I270947);
nand I_15792 (I270500,I270707,I270978);
DFFARX1 I_15793 (I270947,I2507,I270523,I270512,);
DFFARX1 I_15794 (I270947,I2507,I270523,I270509,);
not I_15795 (I271067,I2514);
DFFARX1 I_15796 (I437610,I2507,I271067,I271093,);
DFFARX1 I_15797 (I271093,I2507,I271067,I271110,);
not I_15798 (I271059,I271110);
not I_15799 (I271132,I271093);
nand I_15800 (I271149,I437604,I437601);
and I_15801 (I271166,I271149,I437616);
DFFARX1 I_15802 (I271166,I2507,I271067,I271192,);
not I_15803 (I271200,I271192);
DFFARX1 I_15804 (I437604,I2507,I271067,I271226,);
and I_15805 (I271234,I271226,I437598);
nand I_15806 (I271251,I271226,I437598);
nand I_15807 (I271038,I271200,I271251);
DFFARX1 I_15808 (I437598,I2507,I271067,I271291,);
nor I_15809 (I271299,I271291,I271234);
DFFARX1 I_15810 (I271299,I2507,I271067,I271032,);
nor I_15811 (I271047,I271291,I271192);
nand I_15812 (I271344,I437613,I437607);
and I_15813 (I271361,I271344,I437601);
DFFARX1 I_15814 (I271361,I2507,I271067,I271387,);
nor I_15815 (I271035,I271387,I271291);
not I_15816 (I271409,I271387);
nor I_15817 (I271426,I271409,I271200);
nor I_15818 (I271443,I271132,I271426);
DFFARX1 I_15819 (I271443,I2507,I271067,I271050,);
nor I_15820 (I271474,I271409,I271291);
nor I_15821 (I271491,I437619,I437607);
nor I_15822 (I271041,I271491,I271474);
not I_15823 (I271522,I271491);
nand I_15824 (I271044,I271251,I271522);
DFFARX1 I_15825 (I271491,I2507,I271067,I271056,);
DFFARX1 I_15826 (I271491,I2507,I271067,I271053,);
not I_15827 (I271611,I2514);
DFFARX1 I_15828 (I362274,I2507,I271611,I271637,);
DFFARX1 I_15829 (I271637,I2507,I271611,I271654,);
not I_15830 (I271603,I271654);
not I_15831 (I271676,I271637);
nand I_15832 (I271693,I362295,I362286);
and I_15833 (I271710,I271693,I362274);
DFFARX1 I_15834 (I271710,I2507,I271611,I271736,);
not I_15835 (I271744,I271736);
DFFARX1 I_15836 (I362280,I2507,I271611,I271770,);
and I_15837 (I271778,I271770,I362277);
nand I_15838 (I271795,I271770,I362277);
nand I_15839 (I271582,I271744,I271795);
DFFARX1 I_15840 (I362271,I2507,I271611,I271835,);
nor I_15841 (I271843,I271835,I271778);
DFFARX1 I_15842 (I271843,I2507,I271611,I271576,);
nor I_15843 (I271591,I271835,I271736);
nand I_15844 (I271888,I362271,I362283);
and I_15845 (I271905,I271888,I362292);
DFFARX1 I_15846 (I271905,I2507,I271611,I271931,);
nor I_15847 (I271579,I271931,I271835);
not I_15848 (I271953,I271931);
nor I_15849 (I271970,I271953,I271744);
nor I_15850 (I271987,I271676,I271970);
DFFARX1 I_15851 (I271987,I2507,I271611,I271594,);
nor I_15852 (I272018,I271953,I271835);
nor I_15853 (I272035,I362289,I362283);
nor I_15854 (I271585,I272035,I272018);
not I_15855 (I272066,I272035);
nand I_15856 (I271588,I271795,I272066);
DFFARX1 I_15857 (I272035,I2507,I271611,I271600,);
DFFARX1 I_15858 (I272035,I2507,I271611,I271597,);
not I_15859 (I272155,I2514);
DFFARX1 I_15860 (I74144,I2507,I272155,I272181,);
DFFARX1 I_15861 (I272181,I2507,I272155,I272198,);
not I_15862 (I272147,I272198);
not I_15863 (I272220,I272181);
nand I_15864 (I272237,I74159,I74138);
and I_15865 (I272254,I272237,I74141);
DFFARX1 I_15866 (I272254,I2507,I272155,I272280,);
not I_15867 (I272288,I272280);
DFFARX1 I_15868 (I74147,I2507,I272155,I272314,);
and I_15869 (I272322,I272314,I74141);
nand I_15870 (I272339,I272314,I74141);
nand I_15871 (I272126,I272288,I272339);
DFFARX1 I_15872 (I74156,I2507,I272155,I272379,);
nor I_15873 (I272387,I272379,I272322);
DFFARX1 I_15874 (I272387,I2507,I272155,I272120,);
nor I_15875 (I272135,I272379,I272280);
nand I_15876 (I272432,I74138,I74153);
and I_15877 (I272449,I272432,I74150);
DFFARX1 I_15878 (I272449,I2507,I272155,I272475,);
nor I_15879 (I272123,I272475,I272379);
not I_15880 (I272497,I272475);
nor I_15881 (I272514,I272497,I272288);
nor I_15882 (I272531,I272220,I272514);
DFFARX1 I_15883 (I272531,I2507,I272155,I272138,);
nor I_15884 (I272562,I272497,I272379);
nor I_15885 (I272579,I74162,I74153);
nor I_15886 (I272129,I272579,I272562);
not I_15887 (I272610,I272579);
nand I_15888 (I272132,I272339,I272610);
DFFARX1 I_15889 (I272579,I2507,I272155,I272144,);
DFFARX1 I_15890 (I272579,I2507,I272155,I272141,);
not I_15891 (I272699,I2514);
DFFARX1 I_15892 (I163766,I2507,I272699,I272725,);
DFFARX1 I_15893 (I272725,I2507,I272699,I272742,);
not I_15894 (I272691,I272742);
not I_15895 (I272764,I272725);
nand I_15896 (I272781,I163745,I163769);
and I_15897 (I272798,I272781,I163772);
DFFARX1 I_15898 (I272798,I2507,I272699,I272824,);
not I_15899 (I272832,I272824);
DFFARX1 I_15900 (I163754,I2507,I272699,I272858,);
and I_15901 (I272866,I272858,I163760);
nand I_15902 (I272883,I272858,I163760);
nand I_15903 (I272670,I272832,I272883);
DFFARX1 I_15904 (I163748,I2507,I272699,I272923,);
nor I_15905 (I272931,I272923,I272866);
DFFARX1 I_15906 (I272931,I2507,I272699,I272664,);
nor I_15907 (I272679,I272923,I272824);
nand I_15908 (I272976,I163757,I163745);
and I_15909 (I272993,I272976,I163751);
DFFARX1 I_15910 (I272993,I2507,I272699,I273019,);
nor I_15911 (I272667,I273019,I272923);
not I_15912 (I273041,I273019);
nor I_15913 (I273058,I273041,I272832);
nor I_15914 (I273075,I272764,I273058);
DFFARX1 I_15915 (I273075,I2507,I272699,I272682,);
nor I_15916 (I273106,I273041,I272923);
nor I_15917 (I273123,I163763,I163745);
nor I_15918 (I272673,I273123,I273106);
not I_15919 (I273154,I273123);
nand I_15920 (I272676,I272883,I273154);
DFFARX1 I_15921 (I273123,I2507,I272699,I272688,);
DFFARX1 I_15922 (I273123,I2507,I272699,I272685,);
not I_15923 (I273243,I2514);
DFFARX1 I_15924 (I609828,I2507,I273243,I273269,);
DFFARX1 I_15925 (I273269,I2507,I273243,I273286,);
not I_15926 (I273235,I273286);
not I_15927 (I273308,I273269);
nand I_15928 (I273325,I609840,I609828);
and I_15929 (I273342,I273325,I609831);
DFFARX1 I_15930 (I273342,I2507,I273243,I273368,);
not I_15931 (I273376,I273368);
DFFARX1 I_15932 (I609849,I2507,I273243,I273402,);
and I_15933 (I273410,I273402,I609825);
nand I_15934 (I273427,I273402,I609825);
nand I_15935 (I273214,I273376,I273427);
DFFARX1 I_15936 (I609843,I2507,I273243,I273467,);
nor I_15937 (I273475,I273467,I273410);
DFFARX1 I_15938 (I273475,I2507,I273243,I273208,);
nor I_15939 (I273223,I273467,I273368);
nand I_15940 (I273520,I609837,I609834);
and I_15941 (I273537,I273520,I609846);
DFFARX1 I_15942 (I273537,I2507,I273243,I273563,);
nor I_15943 (I273211,I273563,I273467);
not I_15944 (I273585,I273563);
nor I_15945 (I273602,I273585,I273376);
nor I_15946 (I273619,I273308,I273602);
DFFARX1 I_15947 (I273619,I2507,I273243,I273226,);
nor I_15948 (I273650,I273585,I273467);
nor I_15949 (I273667,I609825,I609834);
nor I_15950 (I273217,I273667,I273650);
not I_15951 (I273698,I273667);
nand I_15952 (I273220,I273427,I273698);
DFFARX1 I_15953 (I273667,I2507,I273243,I273232,);
DFFARX1 I_15954 (I273667,I2507,I273243,I273229,);
not I_15955 (I273787,I2514);
DFFARX1 I_15956 (I344356,I2507,I273787,I273813,);
DFFARX1 I_15957 (I273813,I2507,I273787,I273830,);
not I_15958 (I273779,I273830);
not I_15959 (I273852,I273813);
nand I_15960 (I273869,I344353,I344374);
and I_15961 (I273886,I273869,I344377);
DFFARX1 I_15962 (I273886,I2507,I273787,I273912,);
not I_15963 (I273920,I273912);
DFFARX1 I_15964 (I344362,I2507,I273787,I273946,);
and I_15965 (I273954,I273946,I344365);
nand I_15966 (I273971,I273946,I344365);
nand I_15967 (I273758,I273920,I273971);
DFFARX1 I_15968 (I344368,I2507,I273787,I274011,);
nor I_15969 (I274019,I274011,I273954);
DFFARX1 I_15970 (I274019,I2507,I273787,I273752,);
nor I_15971 (I273767,I274011,I273912);
nand I_15972 (I274064,I344353,I344359);
and I_15973 (I274081,I274064,I344371);
DFFARX1 I_15974 (I274081,I2507,I273787,I274107,);
nor I_15975 (I273755,I274107,I274011);
not I_15976 (I274129,I274107);
nor I_15977 (I274146,I274129,I273920);
nor I_15978 (I274163,I273852,I274146);
DFFARX1 I_15979 (I274163,I2507,I273787,I273770,);
nor I_15980 (I274194,I274129,I274011);
nor I_15981 (I274211,I344356,I344359);
nor I_15982 (I273761,I274211,I274194);
not I_15983 (I274242,I274211);
nand I_15984 (I273764,I273971,I274242);
DFFARX1 I_15985 (I274211,I2507,I273787,I273776,);
DFFARX1 I_15986 (I274211,I2507,I273787,I273773,);
not I_15987 (I274331,I2514);
DFFARX1 I_15988 (I129448,I2507,I274331,I274357,);
DFFARX1 I_15989 (I274357,I2507,I274331,I274374,);
not I_15990 (I274323,I274374);
not I_15991 (I274396,I274357);
nand I_15992 (I274413,I129460,I129439);
and I_15993 (I274430,I274413,I129442);
DFFARX1 I_15994 (I274430,I2507,I274331,I274456,);
not I_15995 (I274464,I274456);
DFFARX1 I_15996 (I129451,I2507,I274331,I274490,);
and I_15997 (I274498,I274490,I129463);
nand I_15998 (I274515,I274490,I129463);
nand I_15999 (I274302,I274464,I274515);
DFFARX1 I_16000 (I129457,I2507,I274331,I274555,);
nor I_16001 (I274563,I274555,I274498);
DFFARX1 I_16002 (I274563,I2507,I274331,I274296,);
nor I_16003 (I274311,I274555,I274456);
nand I_16004 (I274608,I129445,I129442);
and I_16005 (I274625,I274608,I129454);
DFFARX1 I_16006 (I274625,I2507,I274331,I274651,);
nor I_16007 (I274299,I274651,I274555);
not I_16008 (I274673,I274651);
nor I_16009 (I274690,I274673,I274464);
nor I_16010 (I274707,I274396,I274690);
DFFARX1 I_16011 (I274707,I2507,I274331,I274314,);
nor I_16012 (I274738,I274673,I274555);
nor I_16013 (I274755,I129439,I129442);
nor I_16014 (I274305,I274755,I274738);
not I_16015 (I274786,I274755);
nand I_16016 (I274308,I274515,I274786);
DFFARX1 I_16017 (I274755,I2507,I274331,I274320,);
DFFARX1 I_16018 (I274755,I2507,I274331,I274317,);
not I_16019 (I274875,I2514);
DFFARX1 I_16020 (I590176,I2507,I274875,I274901,);
DFFARX1 I_16021 (I274901,I2507,I274875,I274918,);
not I_16022 (I274867,I274918);
not I_16023 (I274940,I274901);
nand I_16024 (I274957,I590188,I590176);
and I_16025 (I274974,I274957,I590179);
DFFARX1 I_16026 (I274974,I2507,I274875,I275000,);
not I_16027 (I275008,I275000);
DFFARX1 I_16028 (I590197,I2507,I274875,I275034,);
and I_16029 (I275042,I275034,I590173);
nand I_16030 (I275059,I275034,I590173);
nand I_16031 (I274846,I275008,I275059);
DFFARX1 I_16032 (I590191,I2507,I274875,I275099,);
nor I_16033 (I275107,I275099,I275042);
DFFARX1 I_16034 (I275107,I2507,I274875,I274840,);
nor I_16035 (I274855,I275099,I275000);
nand I_16036 (I275152,I590185,I590182);
and I_16037 (I275169,I275152,I590194);
DFFARX1 I_16038 (I275169,I2507,I274875,I275195,);
nor I_16039 (I274843,I275195,I275099);
not I_16040 (I275217,I275195);
nor I_16041 (I275234,I275217,I275008);
nor I_16042 (I275251,I274940,I275234);
DFFARX1 I_16043 (I275251,I2507,I274875,I274858,);
nor I_16044 (I275282,I275217,I275099);
nor I_16045 (I275299,I590173,I590182);
nor I_16046 (I274849,I275299,I275282);
not I_16047 (I275330,I275299);
nand I_16048 (I274852,I275059,I275330);
DFFARX1 I_16049 (I275299,I2507,I274875,I274864,);
DFFARX1 I_16050 (I275299,I2507,I274875,I274861,);
not I_16051 (I275419,I2514);
DFFARX1 I_16052 (I215939,I2507,I275419,I275445,);
DFFARX1 I_16053 (I275445,I2507,I275419,I275462,);
not I_16054 (I275411,I275462);
not I_16055 (I275484,I275445);
nand I_16056 (I275501,I215918,I215942);
and I_16057 (I275518,I275501,I215945);
DFFARX1 I_16058 (I275518,I2507,I275419,I275544,);
not I_16059 (I275552,I275544);
DFFARX1 I_16060 (I215927,I2507,I275419,I275578,);
and I_16061 (I275586,I275578,I215933);
nand I_16062 (I275603,I275578,I215933);
nand I_16063 (I275390,I275552,I275603);
DFFARX1 I_16064 (I215921,I2507,I275419,I275643,);
nor I_16065 (I275651,I275643,I275586);
DFFARX1 I_16066 (I275651,I2507,I275419,I275384,);
nor I_16067 (I275399,I275643,I275544);
nand I_16068 (I275696,I215930,I215918);
and I_16069 (I275713,I275696,I215924);
DFFARX1 I_16070 (I275713,I2507,I275419,I275739,);
nor I_16071 (I275387,I275739,I275643);
not I_16072 (I275761,I275739);
nor I_16073 (I275778,I275761,I275552);
nor I_16074 (I275795,I275484,I275778);
DFFARX1 I_16075 (I275795,I2507,I275419,I275402,);
nor I_16076 (I275826,I275761,I275643);
nor I_16077 (I275843,I215936,I215918);
nor I_16078 (I275393,I275843,I275826);
not I_16079 (I275874,I275843);
nand I_16080 (I275396,I275603,I275874);
DFFARX1 I_16081 (I275843,I2507,I275419,I275408,);
DFFARX1 I_16082 (I275843,I2507,I275419,I275405,);
not I_16083 (I275963,I2514);
DFFARX1 I_16084 (I557057,I2507,I275963,I275989,);
DFFARX1 I_16085 (I275989,I2507,I275963,I276006,);
not I_16086 (I275955,I276006);
not I_16087 (I276028,I275989);
nand I_16088 (I276045,I557057,I557075);
and I_16089 (I276062,I276045,I557069);
DFFARX1 I_16090 (I276062,I2507,I275963,I276088,);
not I_16091 (I276096,I276088);
DFFARX1 I_16092 (I557063,I2507,I275963,I276122,);
and I_16093 (I276130,I276122,I557072);
nand I_16094 (I276147,I276122,I557072);
nand I_16095 (I275934,I276096,I276147);
DFFARX1 I_16096 (I557060,I2507,I275963,I276187,);
nor I_16097 (I276195,I276187,I276130);
DFFARX1 I_16098 (I276195,I2507,I275963,I275928,);
nor I_16099 (I275943,I276187,I276088);
nand I_16100 (I276240,I557060,I557078);
and I_16101 (I276257,I276240,I557063);
DFFARX1 I_16102 (I276257,I2507,I275963,I276283,);
nor I_16103 (I275931,I276283,I276187);
not I_16104 (I276305,I276283);
nor I_16105 (I276322,I276305,I276096);
nor I_16106 (I276339,I276028,I276322);
DFFARX1 I_16107 (I276339,I2507,I275963,I275946,);
nor I_16108 (I276370,I276305,I276187);
nor I_16109 (I276387,I557066,I557078);
nor I_16110 (I275937,I276387,I276370);
not I_16111 (I276418,I276387);
nand I_16112 (I275940,I276147,I276418);
DFFARX1 I_16113 (I276387,I2507,I275963,I275952,);
DFFARX1 I_16114 (I276387,I2507,I275963,I275949,);
not I_16115 (I276507,I2514);
DFFARX1 I_16116 (I363430,I2507,I276507,I276533,);
DFFARX1 I_16117 (I276533,I2507,I276507,I276550,);
not I_16118 (I276499,I276550);
not I_16119 (I276572,I276533);
nand I_16120 (I276589,I363451,I363442);
and I_16121 (I276606,I276589,I363430);
DFFARX1 I_16122 (I276606,I2507,I276507,I276632,);
not I_16123 (I276640,I276632);
DFFARX1 I_16124 (I363436,I2507,I276507,I276666,);
and I_16125 (I276674,I276666,I363433);
nand I_16126 (I276691,I276666,I363433);
nand I_16127 (I276478,I276640,I276691);
DFFARX1 I_16128 (I363427,I2507,I276507,I276731,);
nor I_16129 (I276739,I276731,I276674);
DFFARX1 I_16130 (I276739,I2507,I276507,I276472,);
nor I_16131 (I276487,I276731,I276632);
nand I_16132 (I276784,I363427,I363439);
and I_16133 (I276801,I276784,I363448);
DFFARX1 I_16134 (I276801,I2507,I276507,I276827,);
nor I_16135 (I276475,I276827,I276731);
not I_16136 (I276849,I276827);
nor I_16137 (I276866,I276849,I276640);
nor I_16138 (I276883,I276572,I276866);
DFFARX1 I_16139 (I276883,I2507,I276507,I276490,);
nor I_16140 (I276914,I276849,I276731);
nor I_16141 (I276931,I363445,I363439);
nor I_16142 (I276481,I276931,I276914);
not I_16143 (I276962,I276931);
nand I_16144 (I276484,I276691,I276962);
DFFARX1 I_16145 (I276931,I2507,I276507,I276496,);
DFFARX1 I_16146 (I276931,I2507,I276507,I276493,);
not I_16147 (I277051,I2514);
DFFARX1 I_16148 (I648520,I2507,I277051,I277077,);
DFFARX1 I_16149 (I277077,I2507,I277051,I277094,);
not I_16150 (I277043,I277094);
not I_16151 (I277116,I277077);
nand I_16152 (I277133,I648532,I648535);
and I_16153 (I277150,I277133,I648538);
DFFARX1 I_16154 (I277150,I2507,I277051,I277176,);
not I_16155 (I277184,I277176);
DFFARX1 I_16156 (I648523,I2507,I277051,I277210,);
and I_16157 (I277218,I277210,I648529);
nand I_16158 (I277235,I277210,I648529);
nand I_16159 (I277022,I277184,I277235);
DFFARX1 I_16160 (I648517,I2507,I277051,I277275,);
nor I_16161 (I277283,I277275,I277218);
DFFARX1 I_16162 (I277283,I2507,I277051,I277016,);
nor I_16163 (I277031,I277275,I277176);
nand I_16164 (I277328,I648520,I648541);
and I_16165 (I277345,I277328,I648526);
DFFARX1 I_16166 (I277345,I2507,I277051,I277371,);
nor I_16167 (I277019,I277371,I277275);
not I_16168 (I277393,I277371);
nor I_16169 (I277410,I277393,I277184);
nor I_16170 (I277427,I277116,I277410);
DFFARX1 I_16171 (I277427,I2507,I277051,I277034,);
nor I_16172 (I277458,I277393,I277275);
nor I_16173 (I277475,I648517,I648541);
nor I_16174 (I277025,I277475,I277458);
not I_16175 (I277506,I277475);
nand I_16176 (I277028,I277235,I277506);
DFFARX1 I_16177 (I277475,I2507,I277051,I277040,);
DFFARX1 I_16178 (I277475,I2507,I277051,I277037,);
not I_16179 (I277595,I2514);
DFFARX1 I_16180 (I391174,I2507,I277595,I277621,);
DFFARX1 I_16181 (I277621,I2507,I277595,I277638,);
not I_16182 (I277587,I277638);
not I_16183 (I277660,I277621);
nand I_16184 (I277677,I391195,I391186);
and I_16185 (I277694,I277677,I391174);
DFFARX1 I_16186 (I277694,I2507,I277595,I277720,);
not I_16187 (I277728,I277720);
DFFARX1 I_16188 (I391180,I2507,I277595,I277754,);
and I_16189 (I277762,I277754,I391177);
nand I_16190 (I277779,I277754,I391177);
nand I_16191 (I277566,I277728,I277779);
DFFARX1 I_16192 (I391171,I2507,I277595,I277819,);
nor I_16193 (I277827,I277819,I277762);
DFFARX1 I_16194 (I277827,I2507,I277595,I277560,);
nor I_16195 (I277575,I277819,I277720);
nand I_16196 (I277872,I391171,I391183);
and I_16197 (I277889,I277872,I391192);
DFFARX1 I_16198 (I277889,I2507,I277595,I277915,);
nor I_16199 (I277563,I277915,I277819);
not I_16200 (I277937,I277915);
nor I_16201 (I277954,I277937,I277728);
nor I_16202 (I277971,I277660,I277954);
DFFARX1 I_16203 (I277971,I2507,I277595,I277578,);
nor I_16204 (I278002,I277937,I277819);
nor I_16205 (I278019,I391189,I391183);
nor I_16206 (I277569,I278019,I278002);
not I_16207 (I278050,I278019);
nand I_16208 (I277572,I277779,I278050);
DFFARX1 I_16209 (I278019,I2507,I277595,I277584,);
DFFARX1 I_16210 (I278019,I2507,I277595,I277581,);
not I_16211 (I278139,I2514);
DFFARX1 I_16212 (I55699,I2507,I278139,I278165,);
DFFARX1 I_16213 (I278165,I2507,I278139,I278182,);
not I_16214 (I278131,I278182);
not I_16215 (I278204,I278165);
nand I_16216 (I278221,I55714,I55693);
and I_16217 (I278238,I278221,I55696);
DFFARX1 I_16218 (I278238,I2507,I278139,I278264,);
not I_16219 (I278272,I278264);
DFFARX1 I_16220 (I55702,I2507,I278139,I278298,);
and I_16221 (I278306,I278298,I55696);
nand I_16222 (I278323,I278298,I55696);
nand I_16223 (I278110,I278272,I278323);
DFFARX1 I_16224 (I55711,I2507,I278139,I278363,);
nor I_16225 (I278371,I278363,I278306);
DFFARX1 I_16226 (I278371,I2507,I278139,I278104,);
nor I_16227 (I278119,I278363,I278264);
nand I_16228 (I278416,I55693,I55708);
and I_16229 (I278433,I278416,I55705);
DFFARX1 I_16230 (I278433,I2507,I278139,I278459,);
nor I_16231 (I278107,I278459,I278363);
not I_16232 (I278481,I278459);
nor I_16233 (I278498,I278481,I278272);
nor I_16234 (I278515,I278204,I278498);
DFFARX1 I_16235 (I278515,I2507,I278139,I278122,);
nor I_16236 (I278546,I278481,I278363);
nor I_16237 (I278563,I55717,I55708);
nor I_16238 (I278113,I278563,I278546);
not I_16239 (I278594,I278563);
nand I_16240 (I278116,I278323,I278594);
DFFARX1 I_16241 (I278563,I2507,I278139,I278128,);
DFFARX1 I_16242 (I278563,I2507,I278139,I278125,);
not I_16243 (I278683,I2514);
DFFARX1 I_16244 (I2535,I2507,I278683,I278709,);
DFFARX1 I_16245 (I278709,I2507,I278683,I278726,);
not I_16246 (I278675,I278726);
not I_16247 (I278748,I278709);
nand I_16248 (I278765,I2538,I2526);
and I_16249 (I278782,I278765,I2532);
DFFARX1 I_16250 (I278782,I2507,I278683,I278808,);
not I_16251 (I278816,I278808);
DFFARX1 I_16252 (I2520,I2507,I278683,I278842,);
and I_16253 (I278850,I278842,I2517);
nand I_16254 (I278867,I278842,I2517);
nand I_16255 (I278654,I278816,I278867);
DFFARX1 I_16256 (I2523,I2507,I278683,I278907,);
nor I_16257 (I278915,I278907,I278850);
DFFARX1 I_16258 (I278915,I2507,I278683,I278648,);
nor I_16259 (I278663,I278907,I278808);
nand I_16260 (I278960,I2523,I2520);
and I_16261 (I278977,I278960,I2517);
DFFARX1 I_16262 (I278977,I2507,I278683,I279003,);
nor I_16263 (I278651,I279003,I278907);
not I_16264 (I279025,I279003);
nor I_16265 (I279042,I279025,I278816);
nor I_16266 (I279059,I278748,I279042);
DFFARX1 I_16267 (I279059,I2507,I278683,I278666,);
nor I_16268 (I279090,I279025,I278907);
nor I_16269 (I279107,I2529,I2520);
nor I_16270 (I278657,I279107,I279090);
not I_16271 (I279138,I279107);
nand I_16272 (I278660,I278867,I279138);
DFFARX1 I_16273 (I279107,I2507,I278683,I278672,);
DFFARX1 I_16274 (I279107,I2507,I278683,I278669,);
not I_16275 (I279227,I2514);
DFFARX1 I_16276 (I329906,I2507,I279227,I279253,);
DFFARX1 I_16277 (I279253,I2507,I279227,I279270,);
not I_16278 (I279219,I279270);
not I_16279 (I279292,I279253);
nand I_16280 (I279309,I329903,I329924);
and I_16281 (I279326,I279309,I329927);
DFFARX1 I_16282 (I279326,I2507,I279227,I279352,);
not I_16283 (I279360,I279352);
DFFARX1 I_16284 (I329912,I2507,I279227,I279386,);
and I_16285 (I279394,I279386,I329915);
nand I_16286 (I279411,I279386,I329915);
nand I_16287 (I279198,I279360,I279411);
DFFARX1 I_16288 (I329918,I2507,I279227,I279451,);
nor I_16289 (I279459,I279451,I279394);
DFFARX1 I_16290 (I279459,I2507,I279227,I279192,);
nor I_16291 (I279207,I279451,I279352);
nand I_16292 (I279504,I329903,I329909);
and I_16293 (I279521,I279504,I329921);
DFFARX1 I_16294 (I279521,I2507,I279227,I279547,);
nor I_16295 (I279195,I279547,I279451);
not I_16296 (I279569,I279547);
nor I_16297 (I279586,I279569,I279360);
nor I_16298 (I279603,I279292,I279586);
DFFARX1 I_16299 (I279603,I2507,I279227,I279210,);
nor I_16300 (I279634,I279569,I279451);
nor I_16301 (I279651,I329906,I329909);
nor I_16302 (I279201,I279651,I279634);
not I_16303 (I279682,I279651);
nand I_16304 (I279204,I279411,I279682);
DFFARX1 I_16305 (I279651,I2507,I279227,I279216,);
DFFARX1 I_16306 (I279651,I2507,I279227,I279213,);
not I_16307 (I279771,I2514);
DFFARX1 I_16308 (I305052,I2507,I279771,I279797,);
DFFARX1 I_16309 (I279797,I2507,I279771,I279814,);
not I_16310 (I279763,I279814);
not I_16311 (I279836,I279797);
nand I_16312 (I279853,I305049,I305070);
and I_16313 (I279870,I279853,I305073);
DFFARX1 I_16314 (I279870,I2507,I279771,I279896,);
not I_16315 (I279904,I279896);
DFFARX1 I_16316 (I305058,I2507,I279771,I279930,);
and I_16317 (I279938,I279930,I305061);
nand I_16318 (I279955,I279930,I305061);
nand I_16319 (I279742,I279904,I279955);
DFFARX1 I_16320 (I305064,I2507,I279771,I279995,);
nor I_16321 (I280003,I279995,I279938);
DFFARX1 I_16322 (I280003,I2507,I279771,I279736,);
nor I_16323 (I279751,I279995,I279896);
nand I_16324 (I280048,I305049,I305055);
and I_16325 (I280065,I280048,I305067);
DFFARX1 I_16326 (I280065,I2507,I279771,I280091,);
nor I_16327 (I279739,I280091,I279995);
not I_16328 (I280113,I280091);
nor I_16329 (I280130,I280113,I279904);
nor I_16330 (I280147,I279836,I280130);
DFFARX1 I_16331 (I280147,I2507,I279771,I279754,);
nor I_16332 (I280178,I280113,I279995);
nor I_16333 (I280195,I305052,I305055);
nor I_16334 (I279745,I280195,I280178);
not I_16335 (I280226,I280195);
nand I_16336 (I279748,I279955,I280226);
DFFARX1 I_16337 (I280195,I2507,I279771,I279760,);
DFFARX1 I_16338 (I280195,I2507,I279771,I279757,);
not I_16339 (I280315,I2514);
DFFARX1 I_16340 (I526106,I2507,I280315,I280341,);
DFFARX1 I_16341 (I280341,I2507,I280315,I280358,);
not I_16342 (I280307,I280358);
not I_16343 (I280380,I280341);
nand I_16344 (I280397,I526121,I526109);
and I_16345 (I280414,I280397,I526100);
DFFARX1 I_16346 (I280414,I2507,I280315,I280440,);
not I_16347 (I280448,I280440);
DFFARX1 I_16348 (I526112,I2507,I280315,I280474,);
and I_16349 (I280482,I280474,I526103);
nand I_16350 (I280499,I280474,I526103);
nand I_16351 (I280286,I280448,I280499);
DFFARX1 I_16352 (I526118,I2507,I280315,I280539,);
nor I_16353 (I280547,I280539,I280482);
DFFARX1 I_16354 (I280547,I2507,I280315,I280280,);
nor I_16355 (I280295,I280539,I280440);
nand I_16356 (I280592,I526127,I526115);
and I_16357 (I280609,I280592,I526124);
DFFARX1 I_16358 (I280609,I2507,I280315,I280635,);
nor I_16359 (I280283,I280635,I280539);
not I_16360 (I280657,I280635);
nor I_16361 (I280674,I280657,I280448);
nor I_16362 (I280691,I280380,I280674);
DFFARX1 I_16363 (I280691,I2507,I280315,I280298,);
nor I_16364 (I280722,I280657,I280539);
nor I_16365 (I280739,I526100,I526115);
nor I_16366 (I280289,I280739,I280722);
not I_16367 (I280770,I280739);
nand I_16368 (I280292,I280499,I280770);
DFFARX1 I_16369 (I280739,I2507,I280315,I280304,);
DFFARX1 I_16370 (I280739,I2507,I280315,I280301,);
not I_16371 (I280859,I2514);
DFFARX1 I_16372 (I608094,I2507,I280859,I280885,);
DFFARX1 I_16373 (I280885,I2507,I280859,I280902,);
not I_16374 (I280851,I280902);
not I_16375 (I280924,I280885);
nand I_16376 (I280941,I608106,I608094);
and I_16377 (I280958,I280941,I608097);
DFFARX1 I_16378 (I280958,I2507,I280859,I280984,);
not I_16379 (I280992,I280984);
DFFARX1 I_16380 (I608115,I2507,I280859,I281018,);
and I_16381 (I281026,I281018,I608091);
nand I_16382 (I281043,I281018,I608091);
nand I_16383 (I280830,I280992,I281043);
DFFARX1 I_16384 (I608109,I2507,I280859,I281083,);
nor I_16385 (I281091,I281083,I281026);
DFFARX1 I_16386 (I281091,I2507,I280859,I280824,);
nor I_16387 (I280839,I281083,I280984);
nand I_16388 (I281136,I608103,I608100);
and I_16389 (I281153,I281136,I608112);
DFFARX1 I_16390 (I281153,I2507,I280859,I281179,);
nor I_16391 (I280827,I281179,I281083);
not I_16392 (I281201,I281179);
nor I_16393 (I281218,I281201,I280992);
nor I_16394 (I281235,I280924,I281218);
DFFARX1 I_16395 (I281235,I2507,I280859,I280842,);
nor I_16396 (I281266,I281201,I281083);
nor I_16397 (I281283,I608091,I608100);
nor I_16398 (I280833,I281283,I281266);
not I_16399 (I281314,I281283);
nand I_16400 (I280836,I281043,I281314);
DFFARX1 I_16401 (I281283,I2507,I280859,I280848,);
DFFARX1 I_16402 (I281283,I2507,I280859,I280845,);
not I_16403 (I281400,I2514);
DFFARX1 I_16404 (I202758,I2507,I281400,I281426,);
DFFARX1 I_16405 (I281426,I2507,I281400,I281443,);
not I_16406 (I281392,I281443);
DFFARX1 I_16407 (I202746,I2507,I281400,I281474,);
not I_16408 (I281482,I202749);
nor I_16409 (I281499,I281426,I281482);
not I_16410 (I281516,I202752);
not I_16411 (I281533,I202764);
nand I_16412 (I281550,I281533,I202752);
nor I_16413 (I281567,I281482,I281550);
nor I_16414 (I281584,I281474,I281567);
DFFARX1 I_16415 (I281533,I2507,I281400,I281389,);
nor I_16416 (I281615,I202764,I202755);
nand I_16417 (I281632,I281615,I202743);
nor I_16418 (I281649,I281632,I281516);
nand I_16419 (I281374,I281649,I202749);
DFFARX1 I_16420 (I281632,I2507,I281400,I281386,);
nand I_16421 (I281694,I281516,I202764);
nor I_16422 (I281711,I281516,I202764);
nand I_16423 (I281380,I281499,I281711);
not I_16424 (I281742,I202761);
nor I_16425 (I281759,I281742,I281694);
DFFARX1 I_16426 (I281759,I2507,I281400,I281368,);
nor I_16427 (I281790,I281742,I202767);
and I_16428 (I281807,I281790,I202770);
or I_16429 (I281824,I281807,I202743);
DFFARX1 I_16430 (I281824,I2507,I281400,I281850,);
nor I_16431 (I281858,I281850,I281474);
nor I_16432 (I281377,I281426,I281858);
not I_16433 (I281889,I281850);
nor I_16434 (I281906,I281889,I281584);
DFFARX1 I_16435 (I281906,I2507,I281400,I281383,);
nand I_16436 (I281937,I281889,I281516);
nor I_16437 (I281371,I281742,I281937);
not I_16438 (I281995,I2514);
DFFARX1 I_16439 (I96714,I2507,I281995,I282021,);
DFFARX1 I_16440 (I282021,I2507,I281995,I282038,);
not I_16441 (I281987,I282038);
DFFARX1 I_16442 (I96738,I2507,I281995,I282069,);
not I_16443 (I282077,I96732);
nor I_16444 (I282094,I282021,I282077);
not I_16445 (I282111,I96726);
not I_16446 (I282128,I96723);
nand I_16447 (I282145,I282128,I96726);
nor I_16448 (I282162,I282077,I282145);
nor I_16449 (I282179,I282069,I282162);
DFFARX1 I_16450 (I282128,I2507,I281995,I281984,);
nor I_16451 (I282210,I96723,I96717);
nand I_16452 (I282227,I282210,I96735);
nor I_16453 (I282244,I282227,I282111);
nand I_16454 (I281969,I282244,I96732);
DFFARX1 I_16455 (I282227,I2507,I281995,I281981,);
nand I_16456 (I282289,I282111,I96723);
nor I_16457 (I282306,I282111,I96723);
nand I_16458 (I281975,I282094,I282306);
not I_16459 (I282337,I96729);
nor I_16460 (I282354,I282337,I282289);
DFFARX1 I_16461 (I282354,I2507,I281995,I281963,);
nor I_16462 (I282385,I282337,I96714);
and I_16463 (I282402,I282385,I96720);
or I_16464 (I282419,I282402,I96717);
DFFARX1 I_16465 (I282419,I2507,I281995,I282445,);
nor I_16466 (I282453,I282445,I282069);
nor I_16467 (I281972,I282021,I282453);
not I_16468 (I282484,I282445);
nor I_16469 (I282501,I282484,I282179);
DFFARX1 I_16470 (I282501,I2507,I281995,I281978,);
nand I_16471 (I282532,I282484,I282111);
nor I_16472 (I281966,I282337,I282532);
not I_16473 (I282590,I2514);
DFFARX1 I_16474 (I450255,I2507,I282590,I282616,);
DFFARX1 I_16475 (I282616,I2507,I282590,I282633,);
not I_16476 (I282582,I282633);
DFFARX1 I_16477 (I450252,I2507,I282590,I282664,);
not I_16478 (I282672,I450252);
nor I_16479 (I282689,I282616,I282672);
not I_16480 (I282706,I450249);
not I_16481 (I282723,I450264);
nand I_16482 (I282740,I282723,I450249);
nor I_16483 (I282757,I282672,I282740);
nor I_16484 (I282774,I282664,I282757);
DFFARX1 I_16485 (I282723,I2507,I282590,I282579,);
nor I_16486 (I282805,I450264,I450258);
nand I_16487 (I282822,I282805,I450246);
nor I_16488 (I282839,I282822,I282706);
nand I_16489 (I282564,I282839,I450252);
DFFARX1 I_16490 (I282822,I2507,I282590,I282576,);
nand I_16491 (I282884,I282706,I450264);
nor I_16492 (I282901,I282706,I450264);
nand I_16493 (I282570,I282689,I282901);
not I_16494 (I282932,I450267);
nor I_16495 (I282949,I282932,I282884);
DFFARX1 I_16496 (I282949,I2507,I282590,I282558,);
nor I_16497 (I282980,I282932,I450246);
and I_16498 (I282997,I282980,I450261);
or I_16499 (I283014,I282997,I450249);
DFFARX1 I_16500 (I283014,I2507,I282590,I283040,);
nor I_16501 (I283048,I283040,I282664);
nor I_16502 (I282567,I282616,I283048);
not I_16503 (I283079,I283040);
nor I_16504 (I283096,I283079,I282774);
DFFARX1 I_16505 (I283096,I2507,I282590,I282573,);
nand I_16506 (I283127,I283079,I282706);
nor I_16507 (I282561,I282932,I283127);
not I_16508 (I283185,I2514);
DFFARX1 I_16509 (I25127,I2507,I283185,I283211,);
DFFARX1 I_16510 (I283211,I2507,I283185,I283228,);
not I_16511 (I283177,I283228);
DFFARX1 I_16512 (I25127,I2507,I283185,I283259,);
not I_16513 (I283267,I25142);
nor I_16514 (I283284,I283211,I283267);
not I_16515 (I283301,I25145);
not I_16516 (I283318,I25136);
nand I_16517 (I283335,I283318,I25145);
nor I_16518 (I283352,I283267,I283335);
nor I_16519 (I283369,I283259,I283352);
DFFARX1 I_16520 (I283318,I2507,I283185,I283174,);
nor I_16521 (I283400,I25136,I25148);
nand I_16522 (I283417,I283400,I25130);
nor I_16523 (I283434,I283417,I283301);
nand I_16524 (I283159,I283434,I25142);
DFFARX1 I_16525 (I283417,I2507,I283185,I283171,);
nand I_16526 (I283479,I283301,I25136);
nor I_16527 (I283496,I283301,I25136);
nand I_16528 (I283165,I283284,I283496);
not I_16529 (I283527,I25130);
nor I_16530 (I283544,I283527,I283479);
DFFARX1 I_16531 (I283544,I2507,I283185,I283153,);
nor I_16532 (I283575,I283527,I25139);
and I_16533 (I283592,I283575,I25133);
or I_16534 (I283609,I283592,I25151);
DFFARX1 I_16535 (I283609,I2507,I283185,I283635,);
nor I_16536 (I283643,I283635,I283259);
nor I_16537 (I283162,I283211,I283643);
not I_16538 (I283674,I283635);
nor I_16539 (I283691,I283674,I283369);
DFFARX1 I_16540 (I283691,I2507,I283185,I283168,);
nand I_16541 (I283722,I283674,I283301);
nor I_16542 (I283156,I283527,I283722);
not I_16543 (I283780,I2514);
DFFARX1 I_16544 (I460268,I2507,I283780,I283806,);
DFFARX1 I_16545 (I283806,I2507,I283780,I283823,);
not I_16546 (I283772,I283823);
DFFARX1 I_16547 (I460265,I2507,I283780,I283854,);
not I_16548 (I283862,I460265);
nor I_16549 (I283879,I283806,I283862);
not I_16550 (I283896,I460262);
not I_16551 (I283913,I460277);
nand I_16552 (I283930,I283913,I460262);
nor I_16553 (I283947,I283862,I283930);
nor I_16554 (I283964,I283854,I283947);
DFFARX1 I_16555 (I283913,I2507,I283780,I283769,);
nor I_16556 (I283995,I460277,I460271);
nand I_16557 (I284012,I283995,I460259);
nor I_16558 (I284029,I284012,I283896);
nand I_16559 (I283754,I284029,I460265);
DFFARX1 I_16560 (I284012,I2507,I283780,I283766,);
nand I_16561 (I284074,I283896,I460277);
nor I_16562 (I284091,I283896,I460277);
nand I_16563 (I283760,I283879,I284091);
not I_16564 (I284122,I460280);
nor I_16565 (I284139,I284122,I284074);
DFFARX1 I_16566 (I284139,I2507,I283780,I283748,);
nor I_16567 (I284170,I284122,I460259);
and I_16568 (I284187,I284170,I460274);
or I_16569 (I284204,I284187,I460262);
DFFARX1 I_16570 (I284204,I2507,I283780,I284230,);
nor I_16571 (I284238,I284230,I283854);
nor I_16572 (I283757,I283806,I284238);
not I_16573 (I284269,I284230);
nor I_16574 (I284286,I284269,I283964);
DFFARX1 I_16575 (I284286,I2507,I283780,I283763,);
nand I_16576 (I284317,I284269,I283896);
nor I_16577 (I283751,I284122,I284317);
not I_16578 (I284375,I2514);
DFFARX1 I_16579 (I357656,I2507,I284375,I284401,);
DFFARX1 I_16580 (I284401,I2507,I284375,I284418,);
not I_16581 (I284367,I284418);
DFFARX1 I_16582 (I357650,I2507,I284375,I284449,);
not I_16583 (I284457,I357647);
nor I_16584 (I284474,I284401,I284457);
not I_16585 (I284491,I357659);
not I_16586 (I284508,I357662);
nand I_16587 (I284525,I284508,I357659);
nor I_16588 (I284542,I284457,I284525);
nor I_16589 (I284559,I284449,I284542);
DFFARX1 I_16590 (I284508,I2507,I284375,I284364,);
nor I_16591 (I284590,I357662,I357671);
nand I_16592 (I284607,I284590,I357665);
nor I_16593 (I284624,I284607,I284491);
nand I_16594 (I284349,I284624,I357647);
DFFARX1 I_16595 (I284607,I2507,I284375,I284361,);
nand I_16596 (I284669,I284491,I357662);
nor I_16597 (I284686,I284491,I357662);
nand I_16598 (I284355,I284474,I284686);
not I_16599 (I284717,I357653);
nor I_16600 (I284734,I284717,I284669);
DFFARX1 I_16601 (I284734,I2507,I284375,I284343,);
nor I_16602 (I284765,I284717,I357668);
and I_16603 (I284782,I284765,I357647);
or I_16604 (I284799,I284782,I357650);
DFFARX1 I_16605 (I284799,I2507,I284375,I284825,);
nor I_16606 (I284833,I284825,I284449);
nor I_16607 (I284352,I284401,I284833);
not I_16608 (I284864,I284825);
nor I_16609 (I284881,I284864,I284559);
DFFARX1 I_16610 (I284881,I2507,I284375,I284358,);
nand I_16611 (I284912,I284864,I284491);
nor I_16612 (I284346,I284717,I284912);
not I_16613 (I284970,I2514);
DFFARX1 I_16614 (I656677,I2507,I284970,I284996,);
DFFARX1 I_16615 (I284996,I2507,I284970,I285013,);
not I_16616 (I284962,I285013);
DFFARX1 I_16617 (I656692,I2507,I284970,I285044,);
not I_16618 (I285052,I656701);
nor I_16619 (I285069,I284996,I285052);
not I_16620 (I285086,I656680);
not I_16621 (I285103,I656686);
nand I_16622 (I285120,I285103,I656680);
nor I_16623 (I285137,I285052,I285120);
nor I_16624 (I285154,I285044,I285137);
DFFARX1 I_16625 (I285103,I2507,I284970,I284959,);
nor I_16626 (I285185,I656686,I656698);
nand I_16627 (I285202,I285185,I656695);
nor I_16628 (I285219,I285202,I285086);
nand I_16629 (I284944,I285219,I656701);
DFFARX1 I_16630 (I285202,I2507,I284970,I284956,);
nand I_16631 (I285264,I285086,I656686);
nor I_16632 (I285281,I285086,I656686);
nand I_16633 (I284950,I285069,I285281);
not I_16634 (I285312,I656677);
nor I_16635 (I285329,I285312,I285264);
DFFARX1 I_16636 (I285329,I2507,I284970,I284938,);
nor I_16637 (I285360,I285312,I656689);
and I_16638 (I285377,I285360,I656683);
or I_16639 (I285394,I285377,I656680);
DFFARX1 I_16640 (I285394,I2507,I284970,I285420,);
nor I_16641 (I285428,I285420,I285044);
nor I_16642 (I284947,I284996,I285428);
not I_16643 (I285459,I285420);
nor I_16644 (I285476,I285459,I285154);
DFFARX1 I_16645 (I285476,I2507,I284970,I284953,);
nand I_16646 (I285507,I285459,I285086);
nor I_16647 (I284941,I285312,I285507);
not I_16648 (I285565,I2514);
DFFARX1 I_16649 (I730508,I2507,I285565,I285591,);
DFFARX1 I_16650 (I285591,I2507,I285565,I285608,);
not I_16651 (I285557,I285608);
DFFARX1 I_16652 (I730514,I2507,I285565,I285639,);
not I_16653 (I285647,I730529);
nor I_16654 (I285664,I285591,I285647);
not I_16655 (I285681,I730520);
not I_16656 (I285698,I730517);
nand I_16657 (I285715,I285698,I730520);
nor I_16658 (I285732,I285647,I285715);
nor I_16659 (I285749,I285639,I285732);
DFFARX1 I_16660 (I285698,I2507,I285565,I285554,);
nor I_16661 (I285780,I730517,I730508);
nand I_16662 (I285797,I285780,I730532);
nor I_16663 (I285814,I285797,I285681);
nand I_16664 (I285539,I285814,I730529);
DFFARX1 I_16665 (I285797,I2507,I285565,I285551,);
nand I_16666 (I285859,I285681,I730517);
nor I_16667 (I285876,I285681,I730517);
nand I_16668 (I285545,I285664,I285876);
not I_16669 (I285907,I730526);
nor I_16670 (I285924,I285907,I285859);
DFFARX1 I_16671 (I285924,I2507,I285565,I285533,);
nor I_16672 (I285955,I285907,I730511);
and I_16673 (I285972,I285955,I730523);
or I_16674 (I285989,I285972,I730535);
DFFARX1 I_16675 (I285989,I2507,I285565,I286015,);
nor I_16676 (I286023,I286015,I285639);
nor I_16677 (I285542,I285591,I286023);
not I_16678 (I286054,I286015);
nor I_16679 (I286071,I286054,I285749);
DFFARX1 I_16680 (I286071,I2507,I285565,I285548,);
nand I_16681 (I286102,I286054,I285681);
nor I_16682 (I285536,I285907,I286102);
not I_16683 (I286160,I2514);
DFFARX1 I_16684 (I380776,I2507,I286160,I286186,);
DFFARX1 I_16685 (I286186,I2507,I286160,I286203,);
not I_16686 (I286152,I286203);
DFFARX1 I_16687 (I380770,I2507,I286160,I286234,);
not I_16688 (I286242,I380767);
nor I_16689 (I286259,I286186,I286242);
not I_16690 (I286276,I380779);
not I_16691 (I286293,I380782);
nand I_16692 (I286310,I286293,I380779);
nor I_16693 (I286327,I286242,I286310);
nor I_16694 (I286344,I286234,I286327);
DFFARX1 I_16695 (I286293,I2507,I286160,I286149,);
nor I_16696 (I286375,I380782,I380791);
nand I_16697 (I286392,I286375,I380785);
nor I_16698 (I286409,I286392,I286276);
nand I_16699 (I286134,I286409,I380767);
DFFARX1 I_16700 (I286392,I2507,I286160,I286146,);
nand I_16701 (I286454,I286276,I380782);
nor I_16702 (I286471,I286276,I380782);
nand I_16703 (I286140,I286259,I286471);
not I_16704 (I286502,I380773);
nor I_16705 (I286519,I286502,I286454);
DFFARX1 I_16706 (I286519,I2507,I286160,I286128,);
nor I_16707 (I286550,I286502,I380788);
and I_16708 (I286567,I286550,I380767);
or I_16709 (I286584,I286567,I380770);
DFFARX1 I_16710 (I286584,I2507,I286160,I286610,);
nor I_16711 (I286618,I286610,I286234);
nor I_16712 (I286137,I286186,I286618);
not I_16713 (I286649,I286610);
nor I_16714 (I286666,I286649,I286344);
DFFARX1 I_16715 (I286666,I2507,I286160,I286143,);
nand I_16716 (I286697,I286649,I286276);
nor I_16717 (I286131,I286502,I286697);
not I_16718 (I286755,I2514);
DFFARX1 I_16719 (I336264,I2507,I286755,I286781,);
DFFARX1 I_16720 (I286781,I2507,I286755,I286798,);
not I_16721 (I286747,I286798);
DFFARX1 I_16722 (I336276,I2507,I286755,I286829,);
not I_16723 (I286837,I336261);
nor I_16724 (I286854,I286781,I286837);
not I_16725 (I286871,I336279);
not I_16726 (I286888,I336270);
nand I_16727 (I286905,I286888,I336279);
nor I_16728 (I286922,I286837,I286905);
nor I_16729 (I286939,I286829,I286922);
DFFARX1 I_16730 (I286888,I2507,I286755,I286744,);
nor I_16731 (I286970,I336270,I336282);
nand I_16732 (I286987,I286970,I336285);
nor I_16733 (I287004,I286987,I286871);
nand I_16734 (I286729,I287004,I336261);
DFFARX1 I_16735 (I286987,I2507,I286755,I286741,);
nand I_16736 (I287049,I286871,I336270);
nor I_16737 (I287066,I286871,I336270);
nand I_16738 (I286735,I286854,I287066);
not I_16739 (I287097,I336261);
nor I_16740 (I287114,I287097,I287049);
DFFARX1 I_16741 (I287114,I2507,I286755,I286723,);
nor I_16742 (I287145,I287097,I336273);
and I_16743 (I287162,I287145,I336267);
or I_16744 (I287179,I287162,I336264);
DFFARX1 I_16745 (I287179,I2507,I286755,I287205,);
nor I_16746 (I287213,I287205,I286829);
nor I_16747 (I286732,I286781,I287213);
not I_16748 (I287244,I287205);
nor I_16749 (I287261,I287244,I286939);
DFFARX1 I_16750 (I287261,I2507,I286755,I286738,);
nand I_16751 (I287292,I287244,I286871);
nor I_16752 (I286726,I287097,I287292);
not I_16753 (I287350,I2514);
DFFARX1 I_16754 (I238392,I2507,I287350,I287376,);
DFFARX1 I_16755 (I287376,I2507,I287350,I287393,);
not I_16756 (I287342,I287393);
DFFARX1 I_16757 (I238416,I2507,I287350,I287424,);
not I_16758 (I287432,I238395);
nor I_16759 (I287449,I287376,I287432);
not I_16760 (I287466,I238401);
not I_16761 (I287483,I238407);
nand I_16762 (I287500,I287483,I238401);
nor I_16763 (I287517,I287432,I287500);
nor I_16764 (I287534,I287424,I287517);
DFFARX1 I_16765 (I287483,I2507,I287350,I287339,);
nor I_16766 (I287565,I238407,I238419);
nand I_16767 (I287582,I287565,I238413);
nor I_16768 (I287599,I287582,I287466);
nand I_16769 (I287324,I287599,I238395);
DFFARX1 I_16770 (I287582,I2507,I287350,I287336,);
nand I_16771 (I287644,I287466,I238407);
nor I_16772 (I287661,I287466,I238407);
nand I_16773 (I287330,I287449,I287661);
not I_16774 (I287692,I238398);
nor I_16775 (I287709,I287692,I287644);
DFFARX1 I_16776 (I287709,I2507,I287350,I287318,);
nor I_16777 (I287740,I287692,I238392);
and I_16778 (I287757,I287740,I238410);
or I_16779 (I287774,I287757,I238404);
DFFARX1 I_16780 (I287774,I2507,I287350,I287800,);
nor I_16781 (I287808,I287800,I287424);
nor I_16782 (I287327,I287376,I287808);
not I_16783 (I287839,I287800);
nor I_16784 (I287856,I287839,I287534);
DFFARX1 I_16785 (I287856,I2507,I287350,I287333,);
nand I_16786 (I287887,I287839,I287466);
nor I_16787 (I287321,I287692,I287887);
not I_16788 (I287945,I2514);
DFFARX1 I_16789 (I473443,I2507,I287945,I287971,);
DFFARX1 I_16790 (I287971,I2507,I287945,I287988,);
not I_16791 (I287937,I287988);
DFFARX1 I_16792 (I473440,I2507,I287945,I288019,);
not I_16793 (I288027,I473440);
nor I_16794 (I288044,I287971,I288027);
not I_16795 (I288061,I473437);
not I_16796 (I288078,I473452);
nand I_16797 (I288095,I288078,I473437);
nor I_16798 (I288112,I288027,I288095);
nor I_16799 (I288129,I288019,I288112);
DFFARX1 I_16800 (I288078,I2507,I287945,I287934,);
nor I_16801 (I288160,I473452,I473446);
nand I_16802 (I288177,I288160,I473434);
nor I_16803 (I288194,I288177,I288061);
nand I_16804 (I287919,I288194,I473440);
DFFARX1 I_16805 (I288177,I2507,I287945,I287931,);
nand I_16806 (I288239,I288061,I473452);
nor I_16807 (I288256,I288061,I473452);
nand I_16808 (I287925,I288044,I288256);
not I_16809 (I288287,I473455);
nor I_16810 (I288304,I288287,I288239);
DFFARX1 I_16811 (I288304,I2507,I287945,I287913,);
nor I_16812 (I288335,I288287,I473434);
and I_16813 (I288352,I288335,I473449);
or I_16814 (I288369,I288352,I473437);
DFFARX1 I_16815 (I288369,I2507,I287945,I288395,);
nor I_16816 (I288403,I288395,I288019);
nor I_16817 (I287922,I287971,I288403);
not I_16818 (I288434,I288395);
nor I_16819 (I288451,I288434,I288129);
DFFARX1 I_16820 (I288451,I2507,I287945,I287928,);
nand I_16821 (I288482,I288434,I288061);
nor I_16822 (I287916,I288287,I288482);
not I_16823 (I288540,I2514);
DFFARX1 I_16824 (I242200,I2507,I288540,I288566,);
DFFARX1 I_16825 (I288566,I2507,I288540,I288583,);
not I_16826 (I288532,I288583);
DFFARX1 I_16827 (I242224,I2507,I288540,I288614,);
not I_16828 (I288622,I242203);
nor I_16829 (I288639,I288566,I288622);
not I_16830 (I288656,I242209);
not I_16831 (I288673,I242215);
nand I_16832 (I288690,I288673,I242209);
nor I_16833 (I288707,I288622,I288690);
nor I_16834 (I288724,I288614,I288707);
DFFARX1 I_16835 (I288673,I2507,I288540,I288529,);
nor I_16836 (I288755,I242215,I242227);
nand I_16837 (I288772,I288755,I242221);
nor I_16838 (I288789,I288772,I288656);
nand I_16839 (I288514,I288789,I242203);
DFFARX1 I_16840 (I288772,I2507,I288540,I288526,);
nand I_16841 (I288834,I288656,I242215);
nor I_16842 (I288851,I288656,I242215);
nand I_16843 (I288520,I288639,I288851);
not I_16844 (I288882,I242206);
nor I_16845 (I288899,I288882,I288834);
DFFARX1 I_16846 (I288899,I2507,I288540,I288508,);
nor I_16847 (I288930,I288882,I242200);
and I_16848 (I288947,I288930,I242218);
or I_16849 (I288964,I288947,I242212);
DFFARX1 I_16850 (I288964,I2507,I288540,I288990,);
nor I_16851 (I288998,I288990,I288614);
nor I_16852 (I288517,I288566,I288998);
not I_16853 (I289029,I288990);
nor I_16854 (I289046,I289029,I288724);
DFFARX1 I_16855 (I289046,I2507,I288540,I288523,);
nand I_16856 (I289077,I289029,I288656);
nor I_16857 (I288511,I288882,I289077);
not I_16858 (I289135,I2514);
DFFARX1 I_16859 (I664837,I2507,I289135,I289161,);
DFFARX1 I_16860 (I289161,I2507,I289135,I289178,);
not I_16861 (I289127,I289178);
DFFARX1 I_16862 (I664852,I2507,I289135,I289209,);
not I_16863 (I289217,I664861);
nor I_16864 (I289234,I289161,I289217);
not I_16865 (I289251,I664840);
not I_16866 (I289268,I664846);
nand I_16867 (I289285,I289268,I664840);
nor I_16868 (I289302,I289217,I289285);
nor I_16869 (I289319,I289209,I289302);
DFFARX1 I_16870 (I289268,I2507,I289135,I289124,);
nor I_16871 (I289350,I664846,I664858);
nand I_16872 (I289367,I289350,I664855);
nor I_16873 (I289384,I289367,I289251);
nand I_16874 (I289109,I289384,I664861);
DFFARX1 I_16875 (I289367,I2507,I289135,I289121,);
nand I_16876 (I289429,I289251,I664846);
nor I_16877 (I289446,I289251,I664846);
nand I_16878 (I289115,I289234,I289446);
not I_16879 (I289477,I664837);
nor I_16880 (I289494,I289477,I289429);
DFFARX1 I_16881 (I289494,I2507,I289135,I289103,);
nor I_16882 (I289525,I289477,I664849);
and I_16883 (I289542,I289525,I664843);
or I_16884 (I289559,I289542,I664840);
DFFARX1 I_16885 (I289559,I2507,I289135,I289585,);
nor I_16886 (I289593,I289585,I289209);
nor I_16887 (I289112,I289161,I289593);
not I_16888 (I289624,I289585);
nor I_16889 (I289641,I289624,I289319);
DFFARX1 I_16890 (I289641,I2507,I289135,I289118,);
nand I_16891 (I289672,I289624,I289251);
nor I_16892 (I289106,I289477,I289672);
not I_16893 (I289730,I2514);
DFFARX1 I_16894 (I56229,I2507,I289730,I289756,);
DFFARX1 I_16895 (I289756,I2507,I289730,I289773,);
not I_16896 (I289722,I289773);
DFFARX1 I_16897 (I56241,I2507,I289730,I289804,);
not I_16898 (I289812,I56232);
nor I_16899 (I289829,I289756,I289812);
not I_16900 (I289846,I56223);
not I_16901 (I289863,I56220);
nand I_16902 (I289880,I289863,I56223);
nor I_16903 (I289897,I289812,I289880);
nor I_16904 (I289914,I289804,I289897);
DFFARX1 I_16905 (I289863,I2507,I289730,I289719,);
nor I_16906 (I289945,I56220,I56220);
nand I_16907 (I289962,I289945,I56238);
nor I_16908 (I289979,I289962,I289846);
nand I_16909 (I289704,I289979,I56232);
DFFARX1 I_16910 (I289962,I2507,I289730,I289716,);
nand I_16911 (I290024,I289846,I56220);
nor I_16912 (I290041,I289846,I56220);
nand I_16913 (I289710,I289829,I290041);
not I_16914 (I290072,I56244);
nor I_16915 (I290089,I290072,I290024);
DFFARX1 I_16916 (I290089,I2507,I289730,I289698,);
nor I_16917 (I290120,I290072,I56223);
and I_16918 (I290137,I290120,I56226);
or I_16919 (I290154,I290137,I56235);
DFFARX1 I_16920 (I290154,I2507,I289730,I290180,);
nor I_16921 (I290188,I290180,I289804);
nor I_16922 (I289707,I289756,I290188);
not I_16923 (I290219,I290180);
nor I_16924 (I290236,I290219,I289914);
DFFARX1 I_16925 (I290236,I2507,I289730,I289713,);
nand I_16926 (I290267,I290219,I289846);
nor I_16927 (I289701,I290072,I290267);
not I_16928 (I290325,I2514);
DFFARX1 I_16929 (I418346,I2507,I290325,I290351,);
DFFARX1 I_16930 (I290351,I2507,I290325,I290368,);
not I_16931 (I290317,I290368);
DFFARX1 I_16932 (I418340,I2507,I290325,I290399,);
not I_16933 (I290407,I418337);
nor I_16934 (I290424,I290351,I290407);
not I_16935 (I290441,I418349);
not I_16936 (I290458,I418352);
nand I_16937 (I290475,I290458,I418349);
nor I_16938 (I290492,I290407,I290475);
nor I_16939 (I290509,I290399,I290492);
DFFARX1 I_16940 (I290458,I2507,I290325,I290314,);
nor I_16941 (I290540,I418352,I418361);
nand I_16942 (I290557,I290540,I418355);
nor I_16943 (I290574,I290557,I290441);
nand I_16944 (I290299,I290574,I418337);
DFFARX1 I_16945 (I290557,I2507,I290325,I290311,);
nand I_16946 (I290619,I290441,I418352);
nor I_16947 (I290636,I290441,I418352);
nand I_16948 (I290305,I290424,I290636);
not I_16949 (I290667,I418343);
nor I_16950 (I290684,I290667,I290619);
DFFARX1 I_16951 (I290684,I2507,I290325,I290293,);
nor I_16952 (I290715,I290667,I418358);
and I_16953 (I290732,I290715,I418337);
or I_16954 (I290749,I290732,I418340);
DFFARX1 I_16955 (I290749,I2507,I290325,I290775,);
nor I_16956 (I290783,I290775,I290399);
nor I_16957 (I290302,I290351,I290783);
not I_16958 (I290814,I290775);
nor I_16959 (I290831,I290814,I290509);
DFFARX1 I_16960 (I290831,I2507,I290325,I290308,);
nand I_16961 (I290862,I290814,I290441);
nor I_16962 (I290296,I290667,I290862);
not I_16963 (I290920,I2514);
DFFARX1 I_16964 (I668246,I2507,I290920,I290946,);
DFFARX1 I_16965 (I290946,I2507,I290920,I290963,);
not I_16966 (I290912,I290963);
DFFARX1 I_16967 (I668252,I2507,I290920,I290994,);
not I_16968 (I291002,I668240);
nor I_16969 (I291019,I290946,I291002);
not I_16970 (I291036,I668243);
not I_16971 (I291053,I668249);
nand I_16972 (I291070,I291053,I668243);
nor I_16973 (I291087,I291002,I291070);
nor I_16974 (I291104,I290994,I291087);
DFFARX1 I_16975 (I291053,I2507,I290920,I290909,);
nor I_16976 (I291135,I668249,I668240);
nand I_16977 (I291152,I291135,I668258);
nor I_16978 (I291169,I291152,I291036);
nand I_16979 (I290894,I291169,I668240);
DFFARX1 I_16980 (I291152,I2507,I290920,I290906,);
nand I_16981 (I291214,I291036,I668249);
nor I_16982 (I291231,I291036,I668249);
nand I_16983 (I290900,I291019,I291231);
not I_16984 (I291262,I668237);
nor I_16985 (I291279,I291262,I291214);
DFFARX1 I_16986 (I291279,I2507,I290920,I290888,);
nor I_16987 (I291310,I291262,I668261);
and I_16988 (I291327,I291310,I668237);
or I_16989 (I291344,I291327,I668255);
DFFARX1 I_16990 (I291344,I2507,I290920,I291370,);
nor I_16991 (I291378,I291370,I290994);
nor I_16992 (I290897,I290946,I291378);
not I_16993 (I291409,I291370);
nor I_16994 (I291426,I291409,I291104);
DFFARX1 I_16995 (I291426,I2507,I290920,I290903,);
nand I_16996 (I291457,I291409,I291036);
nor I_16997 (I290891,I291262,I291457);
not I_16998 (I291515,I2514);
DFFARX1 I_16999 (I491877,I2507,I291515,I291541,);
DFFARX1 I_17000 (I291541,I2507,I291515,I291558,);
not I_17001 (I291507,I291558);
DFFARX1 I_17002 (I491865,I2507,I291515,I291589,);
not I_17003 (I291597,I491862);
nor I_17004 (I291614,I291541,I291597);
not I_17005 (I291631,I491874);
not I_17006 (I291648,I491871);
nand I_17007 (I291665,I291648,I491874);
nor I_17008 (I291682,I291597,I291665);
nor I_17009 (I291699,I291589,I291682);
DFFARX1 I_17010 (I291648,I2507,I291515,I291504,);
nor I_17011 (I291730,I491871,I491880);
nand I_17012 (I291747,I291730,I491883);
nor I_17013 (I291764,I291747,I291631);
nand I_17014 (I291489,I291764,I491862);
DFFARX1 I_17015 (I291747,I2507,I291515,I291501,);
nand I_17016 (I291809,I291631,I491871);
nor I_17017 (I291826,I291631,I491871);
nand I_17018 (I291495,I291614,I291826);
not I_17019 (I291857,I491886);
nor I_17020 (I291874,I291857,I291809);
DFFARX1 I_17021 (I291874,I2507,I291515,I291483,);
nor I_17022 (I291905,I291857,I491889);
and I_17023 (I291922,I291905,I491868);
or I_17024 (I291939,I291922,I491862);
DFFARX1 I_17025 (I291939,I2507,I291515,I291965,);
nor I_17026 (I291973,I291965,I291589);
nor I_17027 (I291492,I291541,I291973);
not I_17028 (I292004,I291965);
nor I_17029 (I292021,I292004,I291699);
DFFARX1 I_17030 (I292021,I2507,I291515,I291498,);
nand I_17031 (I292052,I292004,I291631);
nor I_17032 (I291486,I291857,I292052);
not I_17033 (I292110,I2514);
DFFARX1 I_17034 (I273752,I2507,I292110,I292136,);
DFFARX1 I_17035 (I292136,I2507,I292110,I292153,);
not I_17036 (I292102,I292153);
DFFARX1 I_17037 (I273776,I2507,I292110,I292184,);
not I_17038 (I292192,I273755);
nor I_17039 (I292209,I292136,I292192);
not I_17040 (I292226,I273761);
not I_17041 (I292243,I273767);
nand I_17042 (I292260,I292243,I273761);
nor I_17043 (I292277,I292192,I292260);
nor I_17044 (I292294,I292184,I292277);
DFFARX1 I_17045 (I292243,I2507,I292110,I292099,);
nor I_17046 (I292325,I273767,I273779);
nand I_17047 (I292342,I292325,I273773);
nor I_17048 (I292359,I292342,I292226);
nand I_17049 (I292084,I292359,I273755);
DFFARX1 I_17050 (I292342,I2507,I292110,I292096,);
nand I_17051 (I292404,I292226,I273767);
nor I_17052 (I292421,I292226,I273767);
nand I_17053 (I292090,I292209,I292421);
not I_17054 (I292452,I273758);
nor I_17055 (I292469,I292452,I292404);
DFFARX1 I_17056 (I292469,I2507,I292110,I292078,);
nor I_17057 (I292500,I292452,I273752);
and I_17058 (I292517,I292500,I273770);
or I_17059 (I292534,I292517,I273764);
DFFARX1 I_17060 (I292534,I2507,I292110,I292560,);
nor I_17061 (I292568,I292560,I292184);
nor I_17062 (I292087,I292136,I292568);
not I_17063 (I292599,I292560);
nor I_17064 (I292616,I292599,I292294);
DFFARX1 I_17065 (I292616,I2507,I292110,I292093,);
nand I_17066 (I292647,I292599,I292226);
nor I_17067 (I292081,I292452,I292647);
not I_17068 (I292705,I2514);
DFFARX1 I_17069 (I133604,I2507,I292705,I292731,);
DFFARX1 I_17070 (I292731,I2507,I292705,I292748,);
not I_17071 (I292697,I292748);
DFFARX1 I_17072 (I133628,I2507,I292705,I292779,);
not I_17073 (I292787,I133622);
nor I_17074 (I292804,I292731,I292787);
not I_17075 (I292821,I133616);
not I_17076 (I292838,I133613);
nand I_17077 (I292855,I292838,I133616);
nor I_17078 (I292872,I292787,I292855);
nor I_17079 (I292889,I292779,I292872);
DFFARX1 I_17080 (I292838,I2507,I292705,I292694,);
nor I_17081 (I292920,I133613,I133607);
nand I_17082 (I292937,I292920,I133625);
nor I_17083 (I292954,I292937,I292821);
nand I_17084 (I292679,I292954,I133622);
DFFARX1 I_17085 (I292937,I2507,I292705,I292691,);
nand I_17086 (I292999,I292821,I133613);
nor I_17087 (I293016,I292821,I133613);
nand I_17088 (I292685,I292804,I293016);
not I_17089 (I293047,I133619);
nor I_17090 (I293064,I293047,I292999);
DFFARX1 I_17091 (I293064,I2507,I292705,I292673,);
nor I_17092 (I293095,I293047,I133604);
and I_17093 (I293112,I293095,I133610);
or I_17094 (I293129,I293112,I133607);
DFFARX1 I_17095 (I293129,I2507,I292705,I293155,);
nor I_17096 (I293163,I293155,I292779);
nor I_17097 (I292682,I292731,I293163);
not I_17098 (I293194,I293155);
nor I_17099 (I293211,I293194,I292889);
DFFARX1 I_17100 (I293211,I2507,I292705,I292688,);
nand I_17101 (I293242,I293194,I292821);
nor I_17102 (I292676,I293047,I293242);
not I_17103 (I293300,I2514);
DFFARX1 I_17104 (I150859,I2507,I293300,I293326,);
DFFARX1 I_17105 (I293326,I2507,I293300,I293343,);
not I_17106 (I293292,I293343);
DFFARX1 I_17107 (I150883,I2507,I293300,I293374,);
not I_17108 (I293382,I150877);
nor I_17109 (I293399,I293326,I293382);
not I_17110 (I293416,I150871);
not I_17111 (I293433,I150868);
nand I_17112 (I293450,I293433,I150871);
nor I_17113 (I293467,I293382,I293450);
nor I_17114 (I293484,I293374,I293467);
DFFARX1 I_17115 (I293433,I2507,I293300,I293289,);
nor I_17116 (I293515,I150868,I150862);
nand I_17117 (I293532,I293515,I150880);
nor I_17118 (I293549,I293532,I293416);
nand I_17119 (I293274,I293549,I150877);
DFFARX1 I_17120 (I293532,I2507,I293300,I293286,);
nand I_17121 (I293594,I293416,I150868);
nor I_17122 (I293611,I293416,I150868);
nand I_17123 (I293280,I293399,I293611);
not I_17124 (I293642,I150874);
nor I_17125 (I293659,I293642,I293594);
DFFARX1 I_17126 (I293659,I2507,I293300,I293268,);
nor I_17127 (I293690,I293642,I150859);
and I_17128 (I293707,I293690,I150865);
or I_17129 (I293724,I293707,I150862);
DFFARX1 I_17130 (I293724,I2507,I293300,I293750,);
nor I_17131 (I293758,I293750,I293374);
nor I_17132 (I293277,I293326,I293758);
not I_17133 (I293789,I293750);
nor I_17134 (I293806,I293789,I293484);
DFFARX1 I_17135 (I293806,I2507,I293300,I293283,);
nand I_17136 (I293837,I293789,I293416);
nor I_17137 (I293271,I293642,I293837);
not I_17138 (I293895,I2514);
DFFARX1 I_17139 (I607531,I2507,I293895,I293921,);
DFFARX1 I_17140 (I293921,I2507,I293895,I293938,);
not I_17141 (I293887,I293938);
DFFARX1 I_17142 (I607513,I2507,I293895,I293969,);
not I_17143 (I293977,I607519);
nor I_17144 (I293994,I293921,I293977);
not I_17145 (I294011,I607534);
not I_17146 (I294028,I607525);
nand I_17147 (I294045,I294028,I607534);
nor I_17148 (I294062,I293977,I294045);
nor I_17149 (I294079,I293969,I294062);
DFFARX1 I_17150 (I294028,I2507,I293895,I293884,);
nor I_17151 (I294110,I607525,I607537);
nand I_17152 (I294127,I294110,I607516);
nor I_17153 (I294144,I294127,I294011);
nand I_17154 (I293869,I294144,I607519);
DFFARX1 I_17155 (I294127,I2507,I293895,I293881,);
nand I_17156 (I294189,I294011,I607525);
nor I_17157 (I294206,I294011,I607525);
nand I_17158 (I293875,I293994,I294206);
not I_17159 (I294237,I607522);
nor I_17160 (I294254,I294237,I294189);
DFFARX1 I_17161 (I294254,I2507,I293895,I293863,);
nor I_17162 (I294285,I294237,I607528);
and I_17163 (I294302,I294285,I607513);
or I_17164 (I294319,I294302,I607516);
DFFARX1 I_17165 (I294319,I2507,I293895,I294345,);
nor I_17166 (I294353,I294345,I293969);
nor I_17167 (I293872,I293921,I294353);
not I_17168 (I294384,I294345);
nor I_17169 (I294401,I294384,I294079);
DFFARX1 I_17170 (I294401,I2507,I293895,I293878,);
nand I_17171 (I294432,I294384,I294011);
nor I_17172 (I293866,I294237,I294432);
not I_17173 (I294490,I2514);
DFFARX1 I_17174 (I612155,I2507,I294490,I294516,);
DFFARX1 I_17175 (I294516,I2507,I294490,I294533,);
not I_17176 (I294482,I294533);
DFFARX1 I_17177 (I612137,I2507,I294490,I294564,);
not I_17178 (I294572,I612143);
nor I_17179 (I294589,I294516,I294572);
not I_17180 (I294606,I612158);
not I_17181 (I294623,I612149);
nand I_17182 (I294640,I294623,I612158);
nor I_17183 (I294657,I294572,I294640);
nor I_17184 (I294674,I294564,I294657);
DFFARX1 I_17185 (I294623,I2507,I294490,I294479,);
nor I_17186 (I294705,I612149,I612161);
nand I_17187 (I294722,I294705,I612140);
nor I_17188 (I294739,I294722,I294606);
nand I_17189 (I294464,I294739,I612143);
DFFARX1 I_17190 (I294722,I2507,I294490,I294476,);
nand I_17191 (I294784,I294606,I612149);
nor I_17192 (I294801,I294606,I612149);
nand I_17193 (I294470,I294589,I294801);
not I_17194 (I294832,I612146);
nor I_17195 (I294849,I294832,I294784);
DFFARX1 I_17196 (I294849,I2507,I294490,I294458,);
nor I_17197 (I294880,I294832,I612152);
and I_17198 (I294897,I294880,I612137);
or I_17199 (I294914,I294897,I612140);
DFFARX1 I_17200 (I294914,I2507,I294490,I294940,);
nor I_17201 (I294948,I294940,I294564);
nor I_17202 (I294467,I294516,I294948);
not I_17203 (I294979,I294940);
nor I_17204 (I294996,I294979,I294674);
DFFARX1 I_17205 (I294996,I2507,I294490,I294473,);
nand I_17206 (I295027,I294979,I294606);
nor I_17207 (I294461,I294832,I295027);
not I_17208 (I295085,I2514);
DFFARX1 I_17209 (I657221,I2507,I295085,I295111,);
DFFARX1 I_17210 (I295111,I2507,I295085,I295128,);
not I_17211 (I295077,I295128);
DFFARX1 I_17212 (I657236,I2507,I295085,I295159,);
not I_17213 (I295167,I657245);
nor I_17214 (I295184,I295111,I295167);
not I_17215 (I295201,I657224);
not I_17216 (I295218,I657230);
nand I_17217 (I295235,I295218,I657224);
nor I_17218 (I295252,I295167,I295235);
nor I_17219 (I295269,I295159,I295252);
DFFARX1 I_17220 (I295218,I2507,I295085,I295074,);
nor I_17221 (I295300,I657230,I657242);
nand I_17222 (I295317,I295300,I657239);
nor I_17223 (I295334,I295317,I295201);
nand I_17224 (I295059,I295334,I657245);
DFFARX1 I_17225 (I295317,I2507,I295085,I295071,);
nand I_17226 (I295379,I295201,I657230);
nor I_17227 (I295396,I295201,I657230);
nand I_17228 (I295065,I295184,I295396);
not I_17229 (I295427,I657221);
nor I_17230 (I295444,I295427,I295379);
DFFARX1 I_17231 (I295444,I2507,I295085,I295053,);
nor I_17232 (I295475,I295427,I657233);
and I_17233 (I295492,I295475,I657227);
or I_17234 (I295509,I295492,I657224);
DFFARX1 I_17235 (I295509,I2507,I295085,I295535,);
nor I_17236 (I295543,I295535,I295159);
nor I_17237 (I295062,I295111,I295543);
not I_17238 (I295574,I295535);
nor I_17239 (I295591,I295574,I295269);
DFFARX1 I_17240 (I295591,I2507,I295085,I295068,);
nand I_17241 (I295622,I295574,I295201);
nor I_17242 (I295056,I295427,I295622);
not I_17243 (I295680,I2514);
DFFARX1 I_17244 (I536451,I2507,I295680,I295706,);
DFFARX1 I_17245 (I295706,I2507,I295680,I295723,);
not I_17246 (I295672,I295723);
DFFARX1 I_17247 (I536439,I2507,I295680,I295754,);
not I_17248 (I295762,I536436);
nor I_17249 (I295779,I295706,I295762);
not I_17250 (I295796,I536448);
not I_17251 (I295813,I536445);
nand I_17252 (I295830,I295813,I536448);
nor I_17253 (I295847,I295762,I295830);
nor I_17254 (I295864,I295754,I295847);
DFFARX1 I_17255 (I295813,I2507,I295680,I295669,);
nor I_17256 (I295895,I536445,I536454);
nand I_17257 (I295912,I295895,I536457);
nor I_17258 (I295929,I295912,I295796);
nand I_17259 (I295654,I295929,I536436);
DFFARX1 I_17260 (I295912,I2507,I295680,I295666,);
nand I_17261 (I295974,I295796,I536445);
nor I_17262 (I295991,I295796,I536445);
nand I_17263 (I295660,I295779,I295991);
not I_17264 (I296022,I536460);
nor I_17265 (I296039,I296022,I295974);
DFFARX1 I_17266 (I296039,I2507,I295680,I295648,);
nor I_17267 (I296070,I296022,I536463);
and I_17268 (I296087,I296070,I536442);
or I_17269 (I296104,I296087,I536436);
DFFARX1 I_17270 (I296104,I2507,I295680,I296130,);
nor I_17271 (I296138,I296130,I295754);
nor I_17272 (I295657,I295706,I296138);
not I_17273 (I296169,I296130);
nor I_17274 (I296186,I296169,I295864);
DFFARX1 I_17275 (I296186,I2507,I295680,I295663,);
nand I_17276 (I296217,I296169,I295796);
nor I_17277 (I295651,I296022,I296217);
not I_17278 (I296275,I2514);
DFFARX1 I_17279 (I57283,I2507,I296275,I296301,);
DFFARX1 I_17280 (I296301,I2507,I296275,I296318,);
not I_17281 (I296267,I296318);
DFFARX1 I_17282 (I57295,I2507,I296275,I296349,);
not I_17283 (I296357,I57286);
nor I_17284 (I296374,I296301,I296357);
not I_17285 (I296391,I57277);
not I_17286 (I296408,I57274);
nand I_17287 (I296425,I296408,I57277);
nor I_17288 (I296442,I296357,I296425);
nor I_17289 (I296459,I296349,I296442);
DFFARX1 I_17290 (I296408,I2507,I296275,I296264,);
nor I_17291 (I296490,I57274,I57274);
nand I_17292 (I296507,I296490,I57292);
nor I_17293 (I296524,I296507,I296391);
nand I_17294 (I296249,I296524,I57286);
DFFARX1 I_17295 (I296507,I2507,I296275,I296261,);
nand I_17296 (I296569,I296391,I57274);
nor I_17297 (I296586,I296391,I57274);
nand I_17298 (I296255,I296374,I296586);
not I_17299 (I296617,I57298);
nor I_17300 (I296634,I296617,I296569);
DFFARX1 I_17301 (I296634,I2507,I296275,I296243,);
nor I_17302 (I296665,I296617,I57277);
and I_17303 (I296682,I296665,I57280);
or I_17304 (I296699,I296682,I57289);
DFFARX1 I_17305 (I296699,I2507,I296275,I296725,);
nor I_17306 (I296733,I296725,I296349);
nor I_17307 (I296252,I296301,I296733);
not I_17308 (I296764,I296725);
nor I_17309 (I296781,I296764,I296459);
DFFARX1 I_17310 (I296781,I2507,I296275,I296258,);
nand I_17311 (I296812,I296764,I296391);
nor I_17312 (I296246,I296617,I296812);
not I_17313 (I296870,I2514);
DFFARX1 I_17314 (I718013,I2507,I296870,I296896,);
DFFARX1 I_17315 (I296896,I2507,I296870,I296913,);
not I_17316 (I296862,I296913);
DFFARX1 I_17317 (I718019,I2507,I296870,I296944,);
not I_17318 (I296952,I718034);
nor I_17319 (I296969,I296896,I296952);
not I_17320 (I296986,I718025);
not I_17321 (I297003,I718022);
nand I_17322 (I297020,I297003,I718025);
nor I_17323 (I297037,I296952,I297020);
nor I_17324 (I297054,I296944,I297037);
DFFARX1 I_17325 (I297003,I2507,I296870,I296859,);
nor I_17326 (I297085,I718022,I718013);
nand I_17327 (I297102,I297085,I718037);
nor I_17328 (I297119,I297102,I296986);
nand I_17329 (I296844,I297119,I718034);
DFFARX1 I_17330 (I297102,I2507,I296870,I296856,);
nand I_17331 (I297164,I296986,I718022);
nor I_17332 (I297181,I296986,I718022);
nand I_17333 (I296850,I296969,I297181);
not I_17334 (I297212,I718031);
nor I_17335 (I297229,I297212,I297164);
DFFARX1 I_17336 (I297229,I2507,I296870,I296838,);
nor I_17337 (I297260,I297212,I718016);
and I_17338 (I297277,I297260,I718028);
or I_17339 (I297294,I297277,I718040);
DFFARX1 I_17340 (I297294,I2507,I296870,I297320,);
nor I_17341 (I297328,I297320,I296944);
nor I_17342 (I296847,I296896,I297328);
not I_17343 (I297359,I297320);
nor I_17344 (I297376,I297359,I297054);
DFFARX1 I_17345 (I297376,I2507,I296870,I296853,);
nand I_17346 (I297407,I297359,I296986);
nor I_17347 (I296841,I297212,I297407);
not I_17348 (I297465,I2514);
DFFARX1 I_17349 (I435499,I2507,I297465,I297491,);
DFFARX1 I_17350 (I297491,I2507,I297465,I297508,);
not I_17351 (I297457,I297508);
DFFARX1 I_17352 (I435496,I2507,I297465,I297539,);
not I_17353 (I297547,I435496);
nor I_17354 (I297564,I297491,I297547);
not I_17355 (I297581,I435493);
not I_17356 (I297598,I435508);
nand I_17357 (I297615,I297598,I435493);
nor I_17358 (I297632,I297547,I297615);
nor I_17359 (I297649,I297539,I297632);
DFFARX1 I_17360 (I297598,I2507,I297465,I297454,);
nor I_17361 (I297680,I435508,I435502);
nand I_17362 (I297697,I297680,I435490);
nor I_17363 (I297714,I297697,I297581);
nand I_17364 (I297439,I297714,I435496);
DFFARX1 I_17365 (I297697,I2507,I297465,I297451,);
nand I_17366 (I297759,I297581,I435508);
nor I_17367 (I297776,I297581,I435508);
nand I_17368 (I297445,I297564,I297776);
not I_17369 (I297807,I435511);
nor I_17370 (I297824,I297807,I297759);
DFFARX1 I_17371 (I297824,I2507,I297465,I297433,);
nor I_17372 (I297855,I297807,I435490);
and I_17373 (I297872,I297855,I435505);
or I_17374 (I297889,I297872,I435493);
DFFARX1 I_17375 (I297889,I2507,I297465,I297915,);
nor I_17376 (I297923,I297915,I297539);
nor I_17377 (I297442,I297491,I297923);
not I_17378 (I297954,I297915);
nor I_17379 (I297971,I297954,I297649);
DFFARX1 I_17380 (I297971,I2507,I297465,I297448,);
nand I_17381 (I298002,I297954,I297581);
nor I_17382 (I297436,I297807,I298002);
not I_17383 (I298060,I2514);
DFFARX1 I_17384 (I99689,I2507,I298060,I298086,);
DFFARX1 I_17385 (I298086,I2507,I298060,I298103,);
not I_17386 (I298052,I298103);
DFFARX1 I_17387 (I99713,I2507,I298060,I298134,);
not I_17388 (I298142,I99707);
nor I_17389 (I298159,I298086,I298142);
not I_17390 (I298176,I99701);
not I_17391 (I298193,I99698);
nand I_17392 (I298210,I298193,I99701);
nor I_17393 (I298227,I298142,I298210);
nor I_17394 (I298244,I298134,I298227);
DFFARX1 I_17395 (I298193,I2507,I298060,I298049,);
nor I_17396 (I298275,I99698,I99692);
nand I_17397 (I298292,I298275,I99710);
nor I_17398 (I298309,I298292,I298176);
nand I_17399 (I298034,I298309,I99707);
DFFARX1 I_17400 (I298292,I2507,I298060,I298046,);
nand I_17401 (I298354,I298176,I99698);
nor I_17402 (I298371,I298176,I99698);
nand I_17403 (I298040,I298159,I298371);
not I_17404 (I298402,I99704);
nor I_17405 (I298419,I298402,I298354);
DFFARX1 I_17406 (I298419,I2507,I298060,I298028,);
nor I_17407 (I298450,I298402,I99689);
and I_17408 (I298467,I298450,I99695);
or I_17409 (I298484,I298467,I99692);
DFFARX1 I_17410 (I298484,I2507,I298060,I298510,);
nor I_17411 (I298518,I298510,I298134);
nor I_17412 (I298037,I298086,I298518);
not I_17413 (I298549,I298510);
nor I_17414 (I298566,I298549,I298244);
DFFARX1 I_17415 (I298566,I2507,I298060,I298043,);
nand I_17416 (I298597,I298549,I298176);
nor I_17417 (I298031,I298402,I298597);
not I_17418 (I298655,I2514);
DFFARX1 I_17419 (I623137,I2507,I298655,I298681,);
DFFARX1 I_17420 (I298681,I2507,I298655,I298698,);
not I_17421 (I298647,I298698);
DFFARX1 I_17422 (I623119,I2507,I298655,I298729,);
not I_17423 (I298737,I623125);
nor I_17424 (I298754,I298681,I298737);
not I_17425 (I298771,I623140);
not I_17426 (I298788,I623131);
nand I_17427 (I298805,I298788,I623140);
nor I_17428 (I298822,I298737,I298805);
nor I_17429 (I298839,I298729,I298822);
DFFARX1 I_17430 (I298788,I2507,I298655,I298644,);
nor I_17431 (I298870,I623131,I623143);
nand I_17432 (I298887,I298870,I623122);
nor I_17433 (I298904,I298887,I298771);
nand I_17434 (I298629,I298904,I623125);
DFFARX1 I_17435 (I298887,I2507,I298655,I298641,);
nand I_17436 (I298949,I298771,I623131);
nor I_17437 (I298966,I298771,I623131);
nand I_17438 (I298635,I298754,I298966);
not I_17439 (I298997,I623128);
nor I_17440 (I299014,I298997,I298949);
DFFARX1 I_17441 (I299014,I2507,I298655,I298623,);
nor I_17442 (I299045,I298997,I623134);
and I_17443 (I299062,I299045,I623119);
or I_17444 (I299079,I299062,I623122);
DFFARX1 I_17445 (I299079,I2507,I298655,I299105,);
nor I_17446 (I299113,I299105,I298729);
nor I_17447 (I298632,I298681,I299113);
not I_17448 (I299144,I299105);
nor I_17449 (I299161,I299144,I298839);
DFFARX1 I_17450 (I299161,I2507,I298655,I298638,);
nand I_17451 (I299192,I299144,I298771);
nor I_17452 (I298626,I298997,I299192);
not I_17453 (I299250,I2514);
DFFARX1 I_17454 (I462376,I2507,I299250,I299276,);
DFFARX1 I_17455 (I299276,I2507,I299250,I299293,);
not I_17456 (I299242,I299293);
DFFARX1 I_17457 (I462373,I2507,I299250,I299324,);
not I_17458 (I299332,I462373);
nor I_17459 (I299349,I299276,I299332);
not I_17460 (I299366,I462370);
not I_17461 (I299383,I462385);
nand I_17462 (I299400,I299383,I462370);
nor I_17463 (I299417,I299332,I299400);
nor I_17464 (I299434,I299324,I299417);
DFFARX1 I_17465 (I299383,I2507,I299250,I299239,);
nor I_17466 (I299465,I462385,I462379);
nand I_17467 (I299482,I299465,I462367);
nor I_17468 (I299499,I299482,I299366);
nand I_17469 (I299224,I299499,I462373);
DFFARX1 I_17470 (I299482,I2507,I299250,I299236,);
nand I_17471 (I299544,I299366,I462385);
nor I_17472 (I299561,I299366,I462385);
nand I_17473 (I299230,I299349,I299561);
not I_17474 (I299592,I462388);
nor I_17475 (I299609,I299592,I299544);
DFFARX1 I_17476 (I299609,I2507,I299250,I299218,);
nor I_17477 (I299640,I299592,I462367);
and I_17478 (I299657,I299640,I462382);
or I_17479 (I299674,I299657,I462370);
DFFARX1 I_17480 (I299674,I2507,I299250,I299700,);
nor I_17481 (I299708,I299700,I299324);
nor I_17482 (I299227,I299276,I299708);
not I_17483 (I299739,I299700);
nor I_17484 (I299756,I299739,I299434);
DFFARX1 I_17485 (I299756,I2507,I299250,I299233,);
nand I_17486 (I299787,I299739,I299366);
nor I_17487 (I299221,I299592,I299787);
not I_17488 (I299845,I2514);
DFFARX1 I_17489 (I444985,I2507,I299845,I299871,);
DFFARX1 I_17490 (I299871,I2507,I299845,I299888,);
not I_17491 (I299837,I299888);
DFFARX1 I_17492 (I444982,I2507,I299845,I299919,);
not I_17493 (I299927,I444982);
nor I_17494 (I299944,I299871,I299927);
not I_17495 (I299961,I444979);
not I_17496 (I299978,I444994);
nand I_17497 (I299995,I299978,I444979);
nor I_17498 (I300012,I299927,I299995);
nor I_17499 (I300029,I299919,I300012);
DFFARX1 I_17500 (I299978,I2507,I299845,I299834,);
nor I_17501 (I300060,I444994,I444988);
nand I_17502 (I300077,I300060,I444976);
nor I_17503 (I300094,I300077,I299961);
nand I_17504 (I299819,I300094,I444982);
DFFARX1 I_17505 (I300077,I2507,I299845,I299831,);
nand I_17506 (I300139,I299961,I444994);
nor I_17507 (I300156,I299961,I444994);
nand I_17508 (I299825,I299944,I300156);
not I_17509 (I300187,I444997);
nor I_17510 (I300204,I300187,I300139);
DFFARX1 I_17511 (I300204,I2507,I299845,I299813,);
nor I_17512 (I300235,I300187,I444976);
and I_17513 (I300252,I300235,I444991);
or I_17514 (I300269,I300252,I444979);
DFFARX1 I_17515 (I300269,I2507,I299845,I300295,);
nor I_17516 (I300303,I300295,I299919);
nor I_17517 (I299822,I299871,I300303);
not I_17518 (I300334,I300295);
nor I_17519 (I300351,I300334,I300029);
DFFARX1 I_17520 (I300351,I2507,I299845,I299828,);
nand I_17521 (I300382,I300334,I299961);
nor I_17522 (I299816,I300187,I300382);
not I_17523 (I300440,I2514);
DFFARX1 I_17524 (I166922,I2507,I300440,I300466,);
DFFARX1 I_17525 (I300466,I2507,I300440,I300483,);
not I_17526 (I300432,I300483);
DFFARX1 I_17527 (I166910,I2507,I300440,I300514,);
not I_17528 (I300522,I166913);
nor I_17529 (I300539,I300466,I300522);
not I_17530 (I300556,I166916);
not I_17531 (I300573,I166928);
nand I_17532 (I300590,I300573,I166916);
nor I_17533 (I300607,I300522,I300590);
nor I_17534 (I300624,I300514,I300607);
DFFARX1 I_17535 (I300573,I2507,I300440,I300429,);
nor I_17536 (I300655,I166928,I166919);
nand I_17537 (I300672,I300655,I166907);
nor I_17538 (I300689,I300672,I300556);
nand I_17539 (I300414,I300689,I166913);
DFFARX1 I_17540 (I300672,I2507,I300440,I300426,);
nand I_17541 (I300734,I300556,I166928);
nor I_17542 (I300751,I300556,I166928);
nand I_17543 (I300420,I300539,I300751);
not I_17544 (I300782,I166925);
nor I_17545 (I300799,I300782,I300734);
DFFARX1 I_17546 (I300799,I2507,I300440,I300408,);
nor I_17547 (I300830,I300782,I166931);
and I_17548 (I300847,I300830,I166934);
or I_17549 (I300864,I300847,I166907);
DFFARX1 I_17550 (I300864,I2507,I300440,I300890,);
nor I_17551 (I300898,I300890,I300514);
nor I_17552 (I300417,I300466,I300898);
not I_17553 (I300929,I300890);
nor I_17554 (I300946,I300929,I300624);
DFFARX1 I_17555 (I300946,I2507,I300440,I300423,);
nand I_17556 (I300977,I300929,I300556);
nor I_17557 (I300411,I300782,I300977);
not I_17558 (I301035,I2514);
DFFARX1 I_17559 (I45177,I2507,I301035,I301061,);
not I_17560 (I301069,I301061);
DFFARX1 I_17561 (I45156,I2507,I301035,I301095,);
not I_17562 (I301103,I45153);
nand I_17563 (I301120,I301103,I45168);
not I_17564 (I301137,I301120);
nor I_17565 (I301154,I301137,I45156);
nor I_17566 (I301171,I301069,I301154);
DFFARX1 I_17567 (I301171,I2507,I301035,I301021,);
not I_17568 (I301202,I45156);
nand I_17569 (I301219,I301202,I301137);
and I_17570 (I301236,I301202,I45159);
nand I_17571 (I301253,I301236,I45174);
nor I_17572 (I301018,I301253,I301202);
and I_17573 (I301009,I301095,I301253);
not I_17574 (I301298,I301253);
nand I_17575 (I301012,I301095,I301298);
nor I_17576 (I301006,I301061,I301253);
not I_17577 (I301343,I45165);
nor I_17578 (I301360,I301343,I45159);
nand I_17579 (I301377,I301360,I301202);
nor I_17580 (I301015,I301120,I301377);
nor I_17581 (I301408,I301343,I45153);
and I_17582 (I301425,I301408,I45162);
or I_17583 (I301442,I301425,I45171);
DFFARX1 I_17584 (I301442,I2507,I301035,I301468,);
nor I_17585 (I301476,I301468,I301219);
DFFARX1 I_17586 (I301476,I2507,I301035,I301003,);
DFFARX1 I_17587 (I301468,I2507,I301035,I301027,);
not I_17588 (I301521,I301468);
nor I_17589 (I301538,I301521,I301095);
nor I_17590 (I301555,I301360,I301538);
DFFARX1 I_17591 (I301555,I2507,I301035,I301024,);
not I_17592 (I301613,I2514);
DFFARX1 I_17593 (I428118,I2507,I301613,I301639,);
not I_17594 (I301647,I301639);
DFFARX1 I_17595 (I428118,I2507,I301613,I301673,);
not I_17596 (I301681,I428115);
nand I_17597 (I301698,I301681,I428130);
not I_17598 (I301715,I301698);
nor I_17599 (I301732,I301715,I428124);
nor I_17600 (I301749,I301647,I301732);
DFFARX1 I_17601 (I301749,I2507,I301613,I301599,);
not I_17602 (I301780,I428124);
nand I_17603 (I301797,I301780,I301715);
and I_17604 (I301814,I301780,I428121);
nand I_17605 (I301831,I301814,I428112);
nor I_17606 (I301596,I301831,I301780);
and I_17607 (I301587,I301673,I301831);
not I_17608 (I301876,I301831);
nand I_17609 (I301590,I301673,I301876);
nor I_17610 (I301584,I301639,I301831);
not I_17611 (I301921,I428133);
nor I_17612 (I301938,I301921,I428121);
nand I_17613 (I301955,I301938,I301780);
nor I_17614 (I301593,I301698,I301955);
nor I_17615 (I301986,I301921,I428112);
and I_17616 (I302003,I301986,I428115);
or I_17617 (I302020,I302003,I428127);
DFFARX1 I_17618 (I302020,I2507,I301613,I302046,);
nor I_17619 (I302054,I302046,I301797);
DFFARX1 I_17620 (I302054,I2507,I301613,I301581,);
DFFARX1 I_17621 (I302046,I2507,I301613,I301605,);
not I_17622 (I302099,I302046);
nor I_17623 (I302116,I302099,I301673);
nor I_17624 (I302133,I301938,I302116);
DFFARX1 I_17625 (I302133,I2507,I301613,I301602,);
not I_17626 (I302191,I2514);
DFFARX1 I_17627 (I376721,I2507,I302191,I302217,);
not I_17628 (I302225,I302217);
DFFARX1 I_17629 (I376733,I2507,I302191,I302251,);
not I_17630 (I302259,I376724);
nand I_17631 (I302276,I302259,I376727);
not I_17632 (I302293,I302276);
nor I_17633 (I302310,I302293,I376730);
nor I_17634 (I302327,I302225,I302310);
DFFARX1 I_17635 (I302327,I2507,I302191,I302177,);
not I_17636 (I302358,I376730);
nand I_17637 (I302375,I302358,I302293);
and I_17638 (I302392,I302358,I376724);
nand I_17639 (I302409,I302392,I376736);
nor I_17640 (I302174,I302409,I302358);
and I_17641 (I302165,I302251,I302409);
not I_17642 (I302454,I302409);
nand I_17643 (I302168,I302251,I302454);
nor I_17644 (I302162,I302217,I302409);
not I_17645 (I302499,I376742);
nor I_17646 (I302516,I302499,I376724);
nand I_17647 (I302533,I302516,I302358);
nor I_17648 (I302171,I302276,I302533);
nor I_17649 (I302564,I302499,I376721);
and I_17650 (I302581,I302564,I376739);
or I_17651 (I302598,I302581,I376745);
DFFARX1 I_17652 (I302598,I2507,I302191,I302624,);
nor I_17653 (I302632,I302624,I302375);
DFFARX1 I_17654 (I302632,I2507,I302191,I302159,);
DFFARX1 I_17655 (I302624,I2507,I302191,I302183,);
not I_17656 (I302677,I302624);
nor I_17657 (I302694,I302677,I302251);
nor I_17658 (I302711,I302516,I302694);
DFFARX1 I_17659 (I302711,I2507,I302191,I302180,);
not I_17660 (I302769,I2514);
DFFARX1 I_17661 (I1628,I2507,I302769,I302795,);
not I_17662 (I302803,I302795);
DFFARX1 I_17663 (I1684,I2507,I302769,I302829,);
not I_17664 (I302837,I1412);
nand I_17665 (I302854,I302837,I2444);
not I_17666 (I302871,I302854);
nor I_17667 (I302888,I302871,I1540);
nor I_17668 (I302905,I302803,I302888);
DFFARX1 I_17669 (I302905,I2507,I302769,I302755,);
not I_17670 (I302936,I1540);
nand I_17671 (I302953,I302936,I302871);
and I_17672 (I302970,I302936,I1852);
nand I_17673 (I302987,I302970,I2348);
nor I_17674 (I302752,I302987,I302936);
and I_17675 (I302743,I302829,I302987);
not I_17676 (I303032,I302987);
nand I_17677 (I302746,I302829,I303032);
nor I_17678 (I302740,I302795,I302987);
not I_17679 (I303077,I1660);
nor I_17680 (I303094,I303077,I1852);
nand I_17681 (I303111,I303094,I302936);
nor I_17682 (I302749,I302854,I303111);
nor I_17683 (I303142,I303077,I2044);
and I_17684 (I303159,I303142,I1364);
or I_17685 (I303176,I303159,I2292);
DFFARX1 I_17686 (I303176,I2507,I302769,I303202,);
nor I_17687 (I303210,I303202,I302953);
DFFARX1 I_17688 (I303210,I2507,I302769,I302737,);
DFFARX1 I_17689 (I303202,I2507,I302769,I302761,);
not I_17690 (I303255,I303202);
nor I_17691 (I303272,I303255,I302829);
nor I_17692 (I303289,I303094,I303272);
DFFARX1 I_17693 (I303289,I2507,I302769,I302758,);
not I_17694 (I303347,I2514);
DFFARX1 I_17695 (I283156,I2507,I303347,I303373,);
not I_17696 (I303381,I303373);
DFFARX1 I_17697 (I283168,I2507,I303347,I303407,);
not I_17698 (I303415,I283174);
nand I_17699 (I303432,I303415,I283165);
not I_17700 (I303449,I303432);
nor I_17701 (I303466,I303449,I283171);
nor I_17702 (I303483,I303381,I303466);
DFFARX1 I_17703 (I303483,I2507,I303347,I303333,);
not I_17704 (I303514,I283171);
nand I_17705 (I303531,I303514,I303449);
and I_17706 (I303548,I303514,I283162);
nand I_17707 (I303565,I303548,I283153);
nor I_17708 (I303330,I303565,I303514);
and I_17709 (I303321,I303407,I303565);
not I_17710 (I303610,I303565);
nand I_17711 (I303324,I303407,I303610);
nor I_17712 (I303318,I303373,I303565);
not I_17713 (I303655,I283159);
nor I_17714 (I303672,I303655,I283162);
nand I_17715 (I303689,I303672,I303514);
nor I_17716 (I303327,I303432,I303689);
nor I_17717 (I303720,I303655,I283156);
and I_17718 (I303737,I303720,I283153);
or I_17719 (I303754,I303737,I283177);
DFFARX1 I_17720 (I303754,I2507,I303347,I303780,);
nor I_17721 (I303788,I303780,I303531);
DFFARX1 I_17722 (I303788,I2507,I303347,I303315,);
DFFARX1 I_17723 (I303780,I2507,I303347,I303339,);
not I_17724 (I303833,I303780);
nor I_17725 (I303850,I303833,I303407);
nor I_17726 (I303867,I303672,I303850);
DFFARX1 I_17727 (I303867,I2507,I303347,I303336,);
not I_17728 (I303925,I2514);
DFFARX1 I_17729 (I614449,I2507,I303925,I303951,);
not I_17730 (I303959,I303951);
DFFARX1 I_17731 (I614455,I2507,I303925,I303985,);
not I_17732 (I303993,I614449);
nand I_17733 (I304010,I303993,I614452);
not I_17734 (I304027,I304010);
nor I_17735 (I304044,I304027,I614470);
nor I_17736 (I304061,I303959,I304044);
DFFARX1 I_17737 (I304061,I2507,I303925,I303911,);
not I_17738 (I304092,I614470);
nand I_17739 (I304109,I304092,I304027);
and I_17740 (I304126,I304092,I614473);
nand I_17741 (I304143,I304126,I614452);
nor I_17742 (I303908,I304143,I304092);
and I_17743 (I303899,I303985,I304143);
not I_17744 (I304188,I304143);
nand I_17745 (I303902,I303985,I304188);
nor I_17746 (I303896,I303951,I304143);
not I_17747 (I304233,I614458);
nor I_17748 (I304250,I304233,I614473);
nand I_17749 (I304267,I304250,I304092);
nor I_17750 (I303905,I304010,I304267);
nor I_17751 (I304298,I304233,I614464);
and I_17752 (I304315,I304298,I614461);
or I_17753 (I304332,I304315,I614467);
DFFARX1 I_17754 (I304332,I2507,I303925,I304358,);
nor I_17755 (I304366,I304358,I304109);
DFFARX1 I_17756 (I304366,I2507,I303925,I303893,);
DFFARX1 I_17757 (I304358,I2507,I303925,I303917,);
not I_17758 (I304411,I304358);
nor I_17759 (I304428,I304411,I303985);
nor I_17760 (I304445,I304250,I304428);
DFFARX1 I_17761 (I304445,I2507,I303925,I303914,);
not I_17762 (I304503,I2514);
DFFARX1 I_17763 (I206438,I2507,I304503,I304529,);
not I_17764 (I304537,I304529);
DFFARX1 I_17765 (I206453,I2507,I304503,I304563,);
not I_17766 (I304571,I206456);
nand I_17767 (I304588,I304571,I206435);
not I_17768 (I304605,I304588);
nor I_17769 (I304622,I304605,I206459);
nor I_17770 (I304639,I304537,I304622);
DFFARX1 I_17771 (I304639,I2507,I304503,I304489,);
not I_17772 (I304670,I206459);
nand I_17773 (I304687,I304670,I304605);
and I_17774 (I304704,I304670,I206441);
nand I_17775 (I304721,I304704,I206432);
nor I_17776 (I304486,I304721,I304670);
and I_17777 (I304477,I304563,I304721);
not I_17778 (I304766,I304721);
nand I_17779 (I304480,I304563,I304766);
nor I_17780 (I304474,I304529,I304721);
not I_17781 (I304811,I206432);
nor I_17782 (I304828,I304811,I206441);
nand I_17783 (I304845,I304828,I304670);
nor I_17784 (I304483,I304588,I304845);
nor I_17785 (I304876,I304811,I206447);
and I_17786 (I304893,I304876,I206450);
or I_17787 (I304910,I304893,I206444);
DFFARX1 I_17788 (I304910,I2507,I304503,I304936,);
nor I_17789 (I304944,I304936,I304687);
DFFARX1 I_17790 (I304944,I2507,I304503,I304471,);
DFFARX1 I_17791 (I304936,I2507,I304503,I304495,);
not I_17792 (I304989,I304936);
nor I_17793 (I305006,I304989,I304563);
nor I_17794 (I305023,I304828,I305006);
DFFARX1 I_17795 (I305023,I2507,I304503,I304492,);
not I_17796 (I305081,I2514);
DFFARX1 I_17797 (I499620,I2507,I305081,I305107,);
not I_17798 (I305115,I305107);
DFFARX1 I_17799 (I499617,I2507,I305081,I305141,);
not I_17800 (I305149,I499614);
nand I_17801 (I305166,I305149,I499641);
not I_17802 (I305183,I305166);
nor I_17803 (I305200,I305183,I499629);
nor I_17804 (I305217,I305115,I305200);
DFFARX1 I_17805 (I305217,I2507,I305081,I305067,);
not I_17806 (I305248,I499629);
nand I_17807 (I305265,I305248,I305183);
and I_17808 (I305282,I305248,I499635);
nand I_17809 (I305299,I305282,I499626);
nor I_17810 (I305064,I305299,I305248);
and I_17811 (I305055,I305141,I305299);
not I_17812 (I305344,I305299);
nand I_17813 (I305058,I305141,I305344);
nor I_17814 (I305052,I305107,I305299);
not I_17815 (I305389,I499623);
nor I_17816 (I305406,I305389,I499635);
nand I_17817 (I305423,I305406,I305248);
nor I_17818 (I305061,I305166,I305423);
nor I_17819 (I305454,I305389,I499638);
and I_17820 (I305471,I305454,I499632);
or I_17821 (I305488,I305471,I499614);
DFFARX1 I_17822 (I305488,I2507,I305081,I305514,);
nor I_17823 (I305522,I305514,I305265);
DFFARX1 I_17824 (I305522,I2507,I305081,I305049,);
DFFARX1 I_17825 (I305514,I2507,I305081,I305073,);
not I_17826 (I305567,I305514);
nor I_17827 (I305584,I305567,I305141);
nor I_17828 (I305601,I305406,I305584);
DFFARX1 I_17829 (I305601,I2507,I305081,I305070,);
not I_17830 (I305659,I2514);
DFFARX1 I_17831 (I547541,I2507,I305659,I305685,);
not I_17832 (I305693,I305685);
DFFARX1 I_17833 (I547532,I2507,I305659,I305719,);
not I_17834 (I305727,I547526);
nand I_17835 (I305744,I305727,I547538);
not I_17836 (I305761,I305744);
nor I_17837 (I305778,I305761,I547529);
nor I_17838 (I305795,I305693,I305778);
DFFARX1 I_17839 (I305795,I2507,I305659,I305645,);
not I_17840 (I305826,I547529);
nand I_17841 (I305843,I305826,I305761);
and I_17842 (I305860,I305826,I547535);
nand I_17843 (I305877,I305860,I547520);
nor I_17844 (I305642,I305877,I305826);
and I_17845 (I305633,I305719,I305877);
not I_17846 (I305922,I305877);
nand I_17847 (I305636,I305719,I305922);
nor I_17848 (I305630,I305685,I305877);
not I_17849 (I305967,I547520);
nor I_17850 (I305984,I305967,I547535);
nand I_17851 (I306001,I305984,I305826);
nor I_17852 (I305639,I305744,I306001);
nor I_17853 (I306032,I305967,I547523);
and I_17854 (I306049,I306032,I547526);
or I_17855 (I306066,I306049,I547523);
DFFARX1 I_17856 (I306066,I2507,I305659,I306092,);
nor I_17857 (I306100,I306092,I305843);
DFFARX1 I_17858 (I306100,I2507,I305659,I305627,);
DFFARX1 I_17859 (I306092,I2507,I305659,I305651,);
not I_17860 (I306145,I306092);
nor I_17861 (I306162,I306145,I305719);
nor I_17862 (I306179,I305984,I306162);
DFFARX1 I_17863 (I306179,I2507,I305659,I305648,);
not I_17864 (I306237,I2514);
DFFARX1 I_17865 (I515124,I2507,I306237,I306263,);
not I_17866 (I306271,I306263);
DFFARX1 I_17867 (I515121,I2507,I306237,I306297,);
not I_17868 (I306305,I515118);
nand I_17869 (I306322,I306305,I515145);
not I_17870 (I306339,I306322);
nor I_17871 (I306356,I306339,I515133);
nor I_17872 (I306373,I306271,I306356);
DFFARX1 I_17873 (I306373,I2507,I306237,I306223,);
not I_17874 (I306404,I515133);
nand I_17875 (I306421,I306404,I306339);
and I_17876 (I306438,I306404,I515139);
nand I_17877 (I306455,I306438,I515130);
nor I_17878 (I306220,I306455,I306404);
and I_17879 (I306211,I306297,I306455);
not I_17880 (I306500,I306455);
nand I_17881 (I306214,I306297,I306500);
nor I_17882 (I306208,I306263,I306455);
not I_17883 (I306545,I515127);
nor I_17884 (I306562,I306545,I515139);
nand I_17885 (I306579,I306562,I306404);
nor I_17886 (I306217,I306322,I306579);
nor I_17887 (I306610,I306545,I515142);
and I_17888 (I306627,I306610,I515136);
or I_17889 (I306644,I306627,I515118);
DFFARX1 I_17890 (I306644,I2507,I306237,I306670,);
nor I_17891 (I306678,I306670,I306421);
DFFARX1 I_17892 (I306678,I2507,I306237,I306205,);
DFFARX1 I_17893 (I306670,I2507,I306237,I306229,);
not I_17894 (I306723,I306670);
nor I_17895 (I306740,I306723,I306297);
nor I_17896 (I306757,I306562,I306740);
DFFARX1 I_17897 (I306757,I2507,I306237,I306226,);
not I_17898 (I306815,I2514);
DFFARX1 I_17899 (I538380,I2507,I306815,I306841,);
not I_17900 (I306849,I306841);
DFFARX1 I_17901 (I538377,I2507,I306815,I306875,);
not I_17902 (I306883,I538374);
nand I_17903 (I306900,I306883,I538401);
not I_17904 (I306917,I306900);
nor I_17905 (I306934,I306917,I538389);
nor I_17906 (I306951,I306849,I306934);
DFFARX1 I_17907 (I306951,I2507,I306815,I306801,);
not I_17908 (I306982,I538389);
nand I_17909 (I306999,I306982,I306917);
and I_17910 (I307016,I306982,I538395);
nand I_17911 (I307033,I307016,I538386);
nor I_17912 (I306798,I307033,I306982);
and I_17913 (I306789,I306875,I307033);
not I_17914 (I307078,I307033);
nand I_17915 (I306792,I306875,I307078);
nor I_17916 (I306786,I306841,I307033);
not I_17917 (I307123,I538383);
nor I_17918 (I307140,I307123,I538395);
nand I_17919 (I307157,I307140,I306982);
nor I_17920 (I306795,I306900,I307157);
nor I_17921 (I307188,I307123,I538398);
and I_17922 (I307205,I307188,I538392);
or I_17923 (I307222,I307205,I538374);
DFFARX1 I_17924 (I307222,I2507,I306815,I307248,);
nor I_17925 (I307256,I307248,I306999);
DFFARX1 I_17926 (I307256,I2507,I306815,I306783,);
DFFARX1 I_17927 (I307248,I2507,I306815,I306807,);
not I_17928 (I307301,I307248);
nor I_17929 (I307318,I307301,I306875);
nor I_17930 (I307335,I307140,I307318);
DFFARX1 I_17931 (I307335,I2507,I306815,I306804,);
not I_17932 (I307393,I2514);
DFFARX1 I_17933 (I106249,I2507,I307393,I307419,);
not I_17934 (I307427,I307419);
DFFARX1 I_17935 (I106234,I2507,I307393,I307453,);
not I_17936 (I307461,I106252);
nand I_17937 (I307478,I307461,I106237);
not I_17938 (I307495,I307478);
nor I_17939 (I307512,I307495,I106234);
nor I_17940 (I307529,I307427,I307512);
DFFARX1 I_17941 (I307529,I2507,I307393,I307379,);
not I_17942 (I307560,I106234);
nand I_17943 (I307577,I307560,I307495);
and I_17944 (I307594,I307560,I106237);
nand I_17945 (I307611,I307594,I106258);
nor I_17946 (I307376,I307611,I307560);
and I_17947 (I307367,I307453,I307611);
not I_17948 (I307656,I307611);
nand I_17949 (I307370,I307453,I307656);
nor I_17950 (I307364,I307419,I307611);
not I_17951 (I307701,I106246);
nor I_17952 (I307718,I307701,I106237);
nand I_17953 (I307735,I307718,I307560);
nor I_17954 (I307373,I307478,I307735);
nor I_17955 (I307766,I307701,I106240);
and I_17956 (I307783,I307766,I106255);
or I_17957 (I307800,I307783,I106243);
DFFARX1 I_17958 (I307800,I2507,I307393,I307826,);
nor I_17959 (I307834,I307826,I307577);
DFFARX1 I_17960 (I307834,I2507,I307393,I307361,);
DFFARX1 I_17961 (I307826,I2507,I307393,I307385,);
not I_17962 (I307879,I307826);
nor I_17963 (I307896,I307879,I307453);
nor I_17964 (I307913,I307718,I307896);
DFFARX1 I_17965 (I307913,I2507,I307393,I307382,);
not I_17966 (I307971,I2514);
DFFARX1 I_17967 (I71527,I2507,I307971,I307997,);
not I_17968 (I308005,I307997);
DFFARX1 I_17969 (I71506,I2507,I307971,I308031,);
not I_17970 (I308039,I71503);
nand I_17971 (I308056,I308039,I71518);
not I_17972 (I308073,I308056);
nor I_17973 (I308090,I308073,I71506);
nor I_17974 (I308107,I308005,I308090);
DFFARX1 I_17975 (I308107,I2507,I307971,I307957,);
not I_17976 (I308138,I71506);
nand I_17977 (I308155,I308138,I308073);
and I_17978 (I308172,I308138,I71509);
nand I_17979 (I308189,I308172,I71524);
nor I_17980 (I307954,I308189,I308138);
and I_17981 (I307945,I308031,I308189);
not I_17982 (I308234,I308189);
nand I_17983 (I307948,I308031,I308234);
nor I_17984 (I307942,I307997,I308189);
not I_17985 (I308279,I71515);
nor I_17986 (I308296,I308279,I71509);
nand I_17987 (I308313,I308296,I308138);
nor I_17988 (I307951,I308056,I308313);
nor I_17989 (I308344,I308279,I71503);
and I_17990 (I308361,I308344,I71512);
or I_17991 (I308378,I308361,I71521);
DFFARX1 I_17992 (I308378,I2507,I307971,I308404,);
nor I_17993 (I308412,I308404,I308155);
DFFARX1 I_17994 (I308412,I2507,I307971,I307939,);
DFFARX1 I_17995 (I308404,I2507,I307971,I307963,);
not I_17996 (I308457,I308404);
nor I_17997 (I308474,I308457,I308031);
nor I_17998 (I308491,I308296,I308474);
DFFARX1 I_17999 (I308491,I2507,I307971,I307960,);
not I_18000 (I308549,I2514);
DFFARX1 I_18001 (I636991,I2507,I308549,I308575,);
not I_18002 (I308583,I308575);
DFFARX1 I_18003 (I636997,I2507,I308549,I308609,);
not I_18004 (I308617,I636991);
nand I_18005 (I308634,I308617,I636994);
not I_18006 (I308651,I308634);
nor I_18007 (I308668,I308651,I637012);
nor I_18008 (I308685,I308583,I308668);
DFFARX1 I_18009 (I308685,I2507,I308549,I308535,);
not I_18010 (I308716,I637012);
nand I_18011 (I308733,I308716,I308651);
and I_18012 (I308750,I308716,I637015);
nand I_18013 (I308767,I308750,I636994);
nor I_18014 (I308532,I308767,I308716);
and I_18015 (I308523,I308609,I308767);
not I_18016 (I308812,I308767);
nand I_18017 (I308526,I308609,I308812);
nor I_18018 (I308520,I308575,I308767);
not I_18019 (I308857,I637000);
nor I_18020 (I308874,I308857,I637015);
nand I_18021 (I308891,I308874,I308716);
nor I_18022 (I308529,I308634,I308891);
nor I_18023 (I308922,I308857,I637006);
and I_18024 (I308939,I308922,I637003);
or I_18025 (I308956,I308939,I637009);
DFFARX1 I_18026 (I308956,I2507,I308549,I308982,);
nor I_18027 (I308990,I308982,I308733);
DFFARX1 I_18028 (I308990,I2507,I308549,I308517,);
DFFARX1 I_18029 (I308982,I2507,I308549,I308541,);
not I_18030 (I309035,I308982);
nor I_18031 (I309052,I309035,I308609);
nor I_18032 (I309069,I308874,I309052);
DFFARX1 I_18033 (I309069,I2507,I308549,I308538,);
not I_18034 (I309127,I2514);
DFFARX1 I_18035 (I33583,I2507,I309127,I309153,);
not I_18036 (I309161,I309153);
DFFARX1 I_18037 (I33562,I2507,I309127,I309187,);
not I_18038 (I309195,I33559);
nand I_18039 (I309212,I309195,I33574);
not I_18040 (I309229,I309212);
nor I_18041 (I309246,I309229,I33562);
nor I_18042 (I309263,I309161,I309246);
DFFARX1 I_18043 (I309263,I2507,I309127,I309113,);
not I_18044 (I309294,I33562);
nand I_18045 (I309311,I309294,I309229);
and I_18046 (I309328,I309294,I33565);
nand I_18047 (I309345,I309328,I33580);
nor I_18048 (I309110,I309345,I309294);
and I_18049 (I309101,I309187,I309345);
not I_18050 (I309390,I309345);
nand I_18051 (I309104,I309187,I309390);
nor I_18052 (I309098,I309153,I309345);
not I_18053 (I309435,I33571);
nor I_18054 (I309452,I309435,I33565);
nand I_18055 (I309469,I309452,I309294);
nor I_18056 (I309107,I309212,I309469);
nor I_18057 (I309500,I309435,I33559);
and I_18058 (I309517,I309500,I33568);
or I_18059 (I309534,I309517,I33577);
DFFARX1 I_18060 (I309534,I2507,I309127,I309560,);
nor I_18061 (I309568,I309560,I309311);
DFFARX1 I_18062 (I309568,I2507,I309127,I309095,);
DFFARX1 I_18063 (I309560,I2507,I309127,I309119,);
not I_18064 (I309613,I309560);
nor I_18065 (I309630,I309613,I309187);
nor I_18066 (I309647,I309452,I309630);
DFFARX1 I_18067 (I309647,I2507,I309127,I309116,);
not I_18068 (I309705,I2514);
DFFARX1 I_18069 (I465535,I2507,I309705,I309731,);
not I_18070 (I309739,I309731);
DFFARX1 I_18071 (I465535,I2507,I309705,I309765,);
not I_18072 (I309773,I465532);
nand I_18073 (I309790,I309773,I465547);
not I_18074 (I309807,I309790);
nor I_18075 (I309824,I309807,I465541);
nor I_18076 (I309841,I309739,I309824);
DFFARX1 I_18077 (I309841,I2507,I309705,I309691,);
not I_18078 (I309872,I465541);
nand I_18079 (I309889,I309872,I309807);
and I_18080 (I309906,I309872,I465538);
nand I_18081 (I309923,I309906,I465529);
nor I_18082 (I309688,I309923,I309872);
and I_18083 (I309679,I309765,I309923);
not I_18084 (I309968,I309923);
nand I_18085 (I309682,I309765,I309968);
nor I_18086 (I309676,I309731,I309923);
not I_18087 (I310013,I465550);
nor I_18088 (I310030,I310013,I465538);
nand I_18089 (I310047,I310030,I309872);
nor I_18090 (I309685,I309790,I310047);
nor I_18091 (I310078,I310013,I465529);
and I_18092 (I310095,I310078,I465532);
or I_18093 (I310112,I310095,I465544);
DFFARX1 I_18094 (I310112,I2507,I309705,I310138,);
nor I_18095 (I310146,I310138,I309889);
DFFARX1 I_18096 (I310146,I2507,I309705,I309673,);
DFFARX1 I_18097 (I310138,I2507,I309705,I309697,);
not I_18098 (I310191,I310138);
nor I_18099 (I310208,I310191,I309765);
nor I_18100 (I310225,I310030,I310208);
DFFARX1 I_18101 (I310225,I2507,I309705,I309694,);
not I_18102 (I310283,I2514);
DFFARX1 I_18103 (I257988,I2507,I310283,I310309,);
not I_18104 (I310317,I310309);
DFFARX1 I_18105 (I258000,I2507,I310283,I310343,);
not I_18106 (I310351,I257976);
nand I_18107 (I310368,I310351,I258003);
not I_18108 (I310385,I310368);
nor I_18109 (I310402,I310385,I257991);
nor I_18110 (I310419,I310317,I310402);
DFFARX1 I_18111 (I310419,I2507,I310283,I310269,);
not I_18112 (I310450,I257991);
nand I_18113 (I310467,I310450,I310385);
and I_18114 (I310484,I310450,I257976);
nand I_18115 (I310501,I310484,I257979);
nor I_18116 (I310266,I310501,I310450);
and I_18117 (I310257,I310343,I310501);
not I_18118 (I310546,I310501);
nand I_18119 (I310260,I310343,I310546);
nor I_18120 (I310254,I310309,I310501);
not I_18121 (I310591,I257985);
nor I_18122 (I310608,I310591,I257976);
nand I_18123 (I310625,I310608,I310450);
nor I_18124 (I310263,I310368,I310625);
nor I_18125 (I310656,I310591,I257994);
and I_18126 (I310673,I310656,I257982);
or I_18127 (I310690,I310673,I257997);
DFFARX1 I_18128 (I310690,I2507,I310283,I310716,);
nor I_18129 (I310724,I310716,I310467);
DFFARX1 I_18130 (I310724,I2507,I310283,I310251,);
DFFARX1 I_18131 (I310716,I2507,I310283,I310275,);
not I_18132 (I310769,I310716);
nor I_18133 (I310786,I310769,I310343);
nor I_18134 (I310803,I310608,I310786);
DFFARX1 I_18135 (I310803,I2507,I310283,I310272,);
not I_18136 (I310861,I2514);
DFFARX1 I_18137 (I680965,I2507,I310861,I310887,);
not I_18138 (I310895,I310887);
DFFARX1 I_18139 (I680977,I2507,I310861,I310921,);
not I_18140 (I310929,I680968);
nand I_18141 (I310946,I310929,I680956);
not I_18142 (I310963,I310946);
nor I_18143 (I310980,I310963,I680953);
nor I_18144 (I310997,I310895,I310980);
DFFARX1 I_18145 (I310997,I2507,I310861,I310847,);
not I_18146 (I311028,I680953);
nand I_18147 (I311045,I311028,I310963);
and I_18148 (I311062,I311028,I680959);
nand I_18149 (I311079,I311062,I680956);
nor I_18150 (I310844,I311079,I311028);
and I_18151 (I310835,I310921,I311079);
not I_18152 (I311124,I311079);
nand I_18153 (I310838,I310921,I311124);
nor I_18154 (I310832,I310887,I311079);
not I_18155 (I311169,I680974);
nor I_18156 (I311186,I311169,I680959);
nand I_18157 (I311203,I311186,I311028);
nor I_18158 (I310841,I310946,I311203);
nor I_18159 (I311234,I311169,I680962);
and I_18160 (I311251,I311234,I680953);
or I_18161 (I311268,I311251,I680971);
DFFARX1 I_18162 (I311268,I2507,I310861,I311294,);
nor I_18163 (I311302,I311294,I311045);
DFFARX1 I_18164 (I311302,I2507,I310861,I310829,);
DFFARX1 I_18165 (I311294,I2507,I310861,I310853,);
not I_18166 (I311347,I311294);
nor I_18167 (I311364,I311347,I310921);
nor I_18168 (I311381,I311186,I311364);
DFFARX1 I_18169 (I311381,I2507,I310861,I310850,);
not I_18170 (I311439,I2514);
DFFARX1 I_18171 (I425273,I2507,I311439,I311465,);
not I_18172 (I311473,I311465);
DFFARX1 I_18173 (I425285,I2507,I311439,I311499,);
not I_18174 (I311507,I425276);
nand I_18175 (I311524,I311507,I425279);
not I_18176 (I311541,I311524);
nor I_18177 (I311558,I311541,I425282);
nor I_18178 (I311575,I311473,I311558);
DFFARX1 I_18179 (I311575,I2507,I311439,I311425,);
not I_18180 (I311606,I425282);
nand I_18181 (I311623,I311606,I311541);
and I_18182 (I311640,I311606,I425276);
nand I_18183 (I311657,I311640,I425288);
nor I_18184 (I311422,I311657,I311606);
and I_18185 (I311413,I311499,I311657);
not I_18186 (I311702,I311657);
nand I_18187 (I311416,I311499,I311702);
nor I_18188 (I311410,I311465,I311657);
not I_18189 (I311747,I425294);
nor I_18190 (I311764,I311747,I425276);
nand I_18191 (I311781,I311764,I311606);
nor I_18192 (I311419,I311524,I311781);
nor I_18193 (I311812,I311747,I425273);
and I_18194 (I311829,I311812,I425291);
or I_18195 (I311846,I311829,I425297);
DFFARX1 I_18196 (I311846,I2507,I311439,I311872,);
nor I_18197 (I311880,I311872,I311623);
DFFARX1 I_18198 (I311880,I2507,I311439,I311407,);
DFFARX1 I_18199 (I311872,I2507,I311439,I311431,);
not I_18200 (I311925,I311872);
nor I_18201 (I311942,I311925,I311499);
nor I_18202 (I311959,I311764,I311942);
DFFARX1 I_18203 (I311959,I2507,I311439,I311428,);
not I_18204 (I312017,I2514);
DFFARX1 I_18205 (I61514,I2507,I312017,I312043,);
not I_18206 (I312051,I312043);
DFFARX1 I_18207 (I61493,I2507,I312017,I312077,);
not I_18208 (I312085,I61490);
nand I_18209 (I312102,I312085,I61505);
not I_18210 (I312119,I312102);
nor I_18211 (I312136,I312119,I61493);
nor I_18212 (I312153,I312051,I312136);
DFFARX1 I_18213 (I312153,I2507,I312017,I312003,);
not I_18214 (I312184,I61493);
nand I_18215 (I312201,I312184,I312119);
and I_18216 (I312218,I312184,I61496);
nand I_18217 (I312235,I312218,I61511);
nor I_18218 (I312000,I312235,I312184);
and I_18219 (I311991,I312077,I312235);
not I_18220 (I312280,I312235);
nand I_18221 (I311994,I312077,I312280);
nor I_18222 (I311988,I312043,I312235);
not I_18223 (I312325,I61502);
nor I_18224 (I312342,I312325,I61496);
nand I_18225 (I312359,I312342,I312184);
nor I_18226 (I311997,I312102,I312359);
nor I_18227 (I312390,I312325,I61490);
and I_18228 (I312407,I312390,I61499);
or I_18229 (I312424,I312407,I61508);
DFFARX1 I_18230 (I312424,I2507,I312017,I312450,);
nor I_18231 (I312458,I312450,I312201);
DFFARX1 I_18232 (I312458,I2507,I312017,I311985,);
DFFARX1 I_18233 (I312450,I2507,I312017,I312009,);
not I_18234 (I312503,I312450);
nor I_18235 (I312520,I312503,I312077);
nor I_18236 (I312537,I312342,I312520);
DFFARX1 I_18237 (I312537,I2507,I312017,I312006,);
not I_18238 (I312595,I2514);
DFFARX1 I_18239 (I51501,I2507,I312595,I312621,);
not I_18240 (I312629,I312621);
DFFARX1 I_18241 (I51480,I2507,I312595,I312655,);
not I_18242 (I312663,I51477);
nand I_18243 (I312680,I312663,I51492);
not I_18244 (I312697,I312680);
nor I_18245 (I312714,I312697,I51480);
nor I_18246 (I312731,I312629,I312714);
DFFARX1 I_18247 (I312731,I2507,I312595,I312581,);
not I_18248 (I312762,I51480);
nand I_18249 (I312779,I312762,I312697);
and I_18250 (I312796,I312762,I51483);
nand I_18251 (I312813,I312796,I51498);
nor I_18252 (I312578,I312813,I312762);
and I_18253 (I312569,I312655,I312813);
not I_18254 (I312858,I312813);
nand I_18255 (I312572,I312655,I312858);
nor I_18256 (I312566,I312621,I312813);
not I_18257 (I312903,I51489);
nor I_18258 (I312920,I312903,I51483);
nand I_18259 (I312937,I312920,I312762);
nor I_18260 (I312575,I312680,I312937);
nor I_18261 (I312968,I312903,I51477);
and I_18262 (I312985,I312968,I51486);
or I_18263 (I313002,I312985,I51495);
DFFARX1 I_18264 (I313002,I2507,I312595,I313028,);
nor I_18265 (I313036,I313028,I312779);
DFFARX1 I_18266 (I313036,I2507,I312595,I312563,);
DFFARX1 I_18267 (I313028,I2507,I312595,I312587,);
not I_18268 (I313081,I313028);
nor I_18269 (I313098,I313081,I312655);
nor I_18270 (I313115,I312920,I313098);
DFFARX1 I_18271 (I313115,I2507,I312595,I312584,);
not I_18272 (I313173,I2514);
DFFARX1 I_18273 (I296841,I2507,I313173,I313199,);
not I_18274 (I313207,I313199);
DFFARX1 I_18275 (I296853,I2507,I313173,I313233,);
not I_18276 (I313241,I296859);
nand I_18277 (I313258,I313241,I296850);
not I_18278 (I313275,I313258);
nor I_18279 (I313292,I313275,I296856);
nor I_18280 (I313309,I313207,I313292);
DFFARX1 I_18281 (I313309,I2507,I313173,I313159,);
not I_18282 (I313340,I296856);
nand I_18283 (I313357,I313340,I313275);
and I_18284 (I313374,I313340,I296847);
nand I_18285 (I313391,I313374,I296838);
nor I_18286 (I313156,I313391,I313340);
and I_18287 (I313147,I313233,I313391);
not I_18288 (I313436,I313391);
nand I_18289 (I313150,I313233,I313436);
nor I_18290 (I313144,I313199,I313391);
not I_18291 (I313481,I296844);
nor I_18292 (I313498,I313481,I296847);
nand I_18293 (I313515,I313498,I313340);
nor I_18294 (I313153,I313258,I313515);
nor I_18295 (I313546,I313481,I296841);
and I_18296 (I313563,I313546,I296838);
or I_18297 (I313580,I313563,I296862);
DFFARX1 I_18298 (I313580,I2507,I313173,I313606,);
nor I_18299 (I313614,I313606,I313357);
DFFARX1 I_18300 (I313614,I2507,I313173,I313141,);
DFFARX1 I_18301 (I313606,I2507,I313173,I313165,);
not I_18302 (I313659,I313606);
nor I_18303 (I313676,I313659,I313233);
nor I_18304 (I313693,I313498,I313676);
DFFARX1 I_18305 (I313693,I2507,I313173,I313162,);
not I_18306 (I313751,I2514);
DFFARX1 I_18307 (I647447,I2507,I313751,I313777,);
not I_18308 (I313785,I313777);
DFFARX1 I_18309 (I647441,I2507,I313751,I313811,);
not I_18310 (I313819,I647450);
nand I_18311 (I313836,I313819,I647429);
not I_18312 (I313853,I313836);
nor I_18313 (I313870,I313853,I647438);
nor I_18314 (I313887,I313785,I313870);
DFFARX1 I_18315 (I313887,I2507,I313751,I313737,);
not I_18316 (I313918,I647438);
nand I_18317 (I313935,I313918,I313853);
and I_18318 (I313952,I313918,I647453);
nand I_18319 (I313969,I313952,I647432);
nor I_18320 (I313734,I313969,I313918);
and I_18321 (I313725,I313811,I313969);
not I_18322 (I314014,I313969);
nand I_18323 (I313728,I313811,I314014);
nor I_18324 (I313722,I313777,I313969);
not I_18325 (I314059,I647435);
nor I_18326 (I314076,I314059,I647453);
nand I_18327 (I314093,I314076,I313918);
nor I_18328 (I313731,I313836,I314093);
nor I_18329 (I314124,I314059,I647444);
and I_18330 (I314141,I314124,I647432);
or I_18331 (I314158,I314141,I647429);
DFFARX1 I_18332 (I314158,I2507,I313751,I314184,);
nor I_18333 (I314192,I314184,I313935);
DFFARX1 I_18334 (I314192,I2507,I313751,I313719,);
DFFARX1 I_18335 (I314184,I2507,I313751,I313743,);
not I_18336 (I314237,I314184);
nor I_18337 (I314254,I314237,I313811);
nor I_18338 (I314271,I314076,I314254);
DFFARX1 I_18339 (I314271,I2507,I313751,I313740,);
not I_18340 (I314329,I2514);
DFFARX1 I_18341 (I213289,I2507,I314329,I314355,);
not I_18342 (I314363,I314355);
DFFARX1 I_18343 (I213304,I2507,I314329,I314389,);
not I_18344 (I314397,I213307);
nand I_18345 (I314414,I314397,I213286);
not I_18346 (I314431,I314414);
nor I_18347 (I314448,I314431,I213310);
nor I_18348 (I314465,I314363,I314448);
DFFARX1 I_18349 (I314465,I2507,I314329,I314315,);
not I_18350 (I314496,I213310);
nand I_18351 (I314513,I314496,I314431);
and I_18352 (I314530,I314496,I213292);
nand I_18353 (I314547,I314530,I213283);
nor I_18354 (I314312,I314547,I314496);
and I_18355 (I314303,I314389,I314547);
not I_18356 (I314592,I314547);
nand I_18357 (I314306,I314389,I314592);
nor I_18358 (I314300,I314355,I314547);
not I_18359 (I314637,I213283);
nor I_18360 (I314654,I314637,I213292);
nand I_18361 (I314671,I314654,I314496);
nor I_18362 (I314309,I314414,I314671);
nor I_18363 (I314702,I314637,I213298);
and I_18364 (I314719,I314702,I213301);
or I_18365 (I314736,I314719,I213295);
DFFARX1 I_18366 (I314736,I2507,I314329,I314762,);
nor I_18367 (I314770,I314762,I314513);
DFFARX1 I_18368 (I314770,I2507,I314329,I314297,);
DFFARX1 I_18369 (I314762,I2507,I314329,I314321,);
not I_18370 (I314815,I314762);
nor I_18371 (I314832,I314815,I314389);
nor I_18372 (I314849,I314654,I314832);
DFFARX1 I_18373 (I314849,I2507,I314329,I314318,);
not I_18374 (I314907,I2514);
DFFARX1 I_18375 (I500912,I2507,I314907,I314933,);
not I_18376 (I314941,I314933);
DFFARX1 I_18377 (I500909,I2507,I314907,I314967,);
not I_18378 (I314975,I500906);
nand I_18379 (I314992,I314975,I500933);
not I_18380 (I315009,I314992);
nor I_18381 (I315026,I315009,I500921);
nor I_18382 (I315043,I314941,I315026);
DFFARX1 I_18383 (I315043,I2507,I314907,I314893,);
not I_18384 (I315074,I500921);
nand I_18385 (I315091,I315074,I315009);
and I_18386 (I315108,I315074,I500927);
nand I_18387 (I315125,I315108,I500918);
nor I_18388 (I314890,I315125,I315074);
and I_18389 (I314881,I314967,I315125);
not I_18390 (I315170,I315125);
nand I_18391 (I314884,I314967,I315170);
nor I_18392 (I314878,I314933,I315125);
not I_18393 (I315215,I500915);
nor I_18394 (I315232,I315215,I500927);
nand I_18395 (I315249,I315232,I315074);
nor I_18396 (I314887,I314992,I315249);
nor I_18397 (I315280,I315215,I500930);
and I_18398 (I315297,I315280,I500924);
or I_18399 (I315314,I315297,I500906);
DFFARX1 I_18400 (I315314,I2507,I314907,I315340,);
nor I_18401 (I315348,I315340,I315091);
DFFARX1 I_18402 (I315348,I2507,I314907,I314875,);
DFFARX1 I_18403 (I315340,I2507,I314907,I314899,);
not I_18404 (I315393,I315340);
nor I_18405 (I315410,I315393,I314967);
nor I_18406 (I315427,I315232,I315410);
DFFARX1 I_18407 (I315427,I2507,I314907,I314896,);
not I_18408 (I315485,I2514);
DFFARX1 I_18409 (I446563,I2507,I315485,I315511,);
not I_18410 (I315519,I315511);
DFFARX1 I_18411 (I446563,I2507,I315485,I315545,);
not I_18412 (I315553,I446560);
nand I_18413 (I315570,I315553,I446575);
not I_18414 (I315587,I315570);
nor I_18415 (I315604,I315587,I446569);
nor I_18416 (I315621,I315519,I315604);
DFFARX1 I_18417 (I315621,I2507,I315485,I315471,);
not I_18418 (I315652,I446569);
nand I_18419 (I315669,I315652,I315587);
and I_18420 (I315686,I315652,I446566);
nand I_18421 (I315703,I315686,I446557);
nor I_18422 (I315468,I315703,I315652);
and I_18423 (I315459,I315545,I315703);
not I_18424 (I315748,I315703);
nand I_18425 (I315462,I315545,I315748);
nor I_18426 (I315456,I315511,I315703);
not I_18427 (I315793,I446578);
nor I_18428 (I315810,I315793,I446566);
nand I_18429 (I315827,I315810,I315652);
nor I_18430 (I315465,I315570,I315827);
nor I_18431 (I315858,I315793,I446557);
and I_18432 (I315875,I315858,I446560);
or I_18433 (I315892,I315875,I446572);
DFFARX1 I_18434 (I315892,I2507,I315485,I315918,);
nor I_18435 (I315926,I315918,I315669);
DFFARX1 I_18436 (I315926,I2507,I315485,I315453,);
DFFARX1 I_18437 (I315918,I2507,I315485,I315477,);
not I_18438 (I315971,I315918);
nor I_18439 (I315988,I315971,I315545);
nor I_18440 (I316005,I315810,I315988);
DFFARX1 I_18441 (I316005,I2507,I315485,I315474,);
not I_18442 (I316063,I2514);
DFFARX1 I_18443 (I222775,I2507,I316063,I316089,);
not I_18444 (I316097,I316089);
DFFARX1 I_18445 (I222790,I2507,I316063,I316123,);
not I_18446 (I316131,I222793);
nand I_18447 (I316148,I316131,I222772);
not I_18448 (I316165,I316148);
nor I_18449 (I316182,I316165,I222796);
nor I_18450 (I316199,I316097,I316182);
DFFARX1 I_18451 (I316199,I2507,I316063,I316049,);
not I_18452 (I316230,I222796);
nand I_18453 (I316247,I316230,I316165);
and I_18454 (I316264,I316230,I222778);
nand I_18455 (I316281,I316264,I222769);
nor I_18456 (I316046,I316281,I316230);
and I_18457 (I316037,I316123,I316281);
not I_18458 (I316326,I316281);
nand I_18459 (I316040,I316123,I316326);
nor I_18460 (I316034,I316089,I316281);
not I_18461 (I316371,I222769);
nor I_18462 (I316388,I316371,I222778);
nand I_18463 (I316405,I316388,I316230);
nor I_18464 (I316043,I316148,I316405);
nor I_18465 (I316436,I316371,I222784);
and I_18466 (I316453,I316436,I222787);
or I_18467 (I316470,I316453,I222781);
DFFARX1 I_18468 (I316470,I2507,I316063,I316496,);
nor I_18469 (I316504,I316496,I316247);
DFFARX1 I_18470 (I316504,I2507,I316063,I316031,);
DFFARX1 I_18471 (I316496,I2507,I316063,I316055,);
not I_18472 (I316549,I316496);
nor I_18473 (I316566,I316549,I316123);
nor I_18474 (I316583,I316388,I316566);
DFFARX1 I_18475 (I316583,I2507,I316063,I316052,);
not I_18476 (I316641,I2514);
DFFARX1 I_18477 (I125289,I2507,I316641,I316667,);
not I_18478 (I316675,I316667);
DFFARX1 I_18479 (I125274,I2507,I316641,I316701,);
not I_18480 (I316709,I125292);
nand I_18481 (I316726,I316709,I125277);
not I_18482 (I316743,I316726);
nor I_18483 (I316760,I316743,I125274);
nor I_18484 (I316777,I316675,I316760);
DFFARX1 I_18485 (I316777,I2507,I316641,I316627,);
not I_18486 (I316808,I125274);
nand I_18487 (I316825,I316808,I316743);
and I_18488 (I316842,I316808,I125277);
nand I_18489 (I316859,I316842,I125298);
nor I_18490 (I316624,I316859,I316808);
and I_18491 (I316615,I316701,I316859);
not I_18492 (I316904,I316859);
nand I_18493 (I316618,I316701,I316904);
nor I_18494 (I316612,I316667,I316859);
not I_18495 (I316949,I125286);
nor I_18496 (I316966,I316949,I125277);
nand I_18497 (I316983,I316966,I316808);
nor I_18498 (I316621,I316726,I316983);
nor I_18499 (I317014,I316949,I125280);
and I_18500 (I317031,I317014,I125295);
or I_18501 (I317048,I317031,I125283);
DFFARX1 I_18502 (I317048,I2507,I316641,I317074,);
nor I_18503 (I317082,I317074,I316825);
DFFARX1 I_18504 (I317082,I2507,I316641,I316609,);
DFFARX1 I_18505 (I317074,I2507,I316641,I316633,);
not I_18506 (I317127,I317074);
nor I_18507 (I317144,I317127,I316701);
nor I_18508 (I317161,I316966,I317144);
DFFARX1 I_18509 (I317161,I2507,I316641,I316630,);
not I_18510 (I317219,I2514);
DFFARX1 I_18511 (I239492,I2507,I317219,I317245,);
not I_18512 (I317253,I317245);
DFFARX1 I_18513 (I239504,I2507,I317219,I317279,);
not I_18514 (I317287,I239480);
nand I_18515 (I317304,I317287,I239507);
not I_18516 (I317321,I317304);
nor I_18517 (I317338,I317321,I239495);
nor I_18518 (I317355,I317253,I317338);
DFFARX1 I_18519 (I317355,I2507,I317219,I317205,);
not I_18520 (I317386,I239495);
nand I_18521 (I317403,I317386,I317321);
and I_18522 (I317420,I317386,I239480);
nand I_18523 (I317437,I317420,I239483);
nor I_18524 (I317202,I317437,I317386);
and I_18525 (I317193,I317279,I317437);
not I_18526 (I317482,I317437);
nand I_18527 (I317196,I317279,I317482);
nor I_18528 (I317190,I317245,I317437);
not I_18529 (I317527,I239489);
nor I_18530 (I317544,I317527,I239480);
nand I_18531 (I317561,I317544,I317386);
nor I_18532 (I317199,I317304,I317561);
nor I_18533 (I317592,I317527,I239498);
and I_18534 (I317609,I317592,I239486);
or I_18535 (I317626,I317609,I239501);
DFFARX1 I_18536 (I317626,I2507,I317219,I317652,);
nor I_18537 (I317660,I317652,I317403);
DFFARX1 I_18538 (I317660,I2507,I317219,I317187,);
DFFARX1 I_18539 (I317652,I2507,I317219,I317211,);
not I_18540 (I317705,I317652);
nor I_18541 (I317722,I317705,I317279);
nor I_18542 (I317739,I317544,I317722);
DFFARX1 I_18543 (I317739,I2507,I317219,I317208,);
not I_18544 (I317797,I2514);
DFFARX1 I_18545 (I573411,I2507,I317797,I317823,);
not I_18546 (I317831,I317823);
DFFARX1 I_18547 (I573417,I2507,I317797,I317857,);
not I_18548 (I317865,I573411);
nand I_18549 (I317882,I317865,I573414);
not I_18550 (I317899,I317882);
nor I_18551 (I317916,I317899,I573432);
nor I_18552 (I317933,I317831,I317916);
DFFARX1 I_18553 (I317933,I2507,I317797,I317783,);
not I_18554 (I317964,I573432);
nand I_18555 (I317981,I317964,I317899);
and I_18556 (I317998,I317964,I573435);
nand I_18557 (I318015,I317998,I573414);
nor I_18558 (I317780,I318015,I317964);
and I_18559 (I317771,I317857,I318015);
not I_18560 (I318060,I318015);
nand I_18561 (I317774,I317857,I318060);
nor I_18562 (I317768,I317823,I318015);
not I_18563 (I318105,I573420);
nor I_18564 (I318122,I318105,I573435);
nand I_18565 (I318139,I318122,I317964);
nor I_18566 (I317777,I317882,I318139);
nor I_18567 (I318170,I318105,I573426);
and I_18568 (I318187,I318170,I573423);
or I_18569 (I318204,I318187,I573429);
DFFARX1 I_18570 (I318204,I2507,I317797,I318230,);
nor I_18571 (I318238,I318230,I317981);
DFFARX1 I_18572 (I318238,I2507,I317797,I317765,);
DFFARX1 I_18573 (I318230,I2507,I317797,I317789,);
not I_18574 (I318283,I318230);
nor I_18575 (I318300,I318283,I317857);
nor I_18576 (I318317,I318122,I318300);
DFFARX1 I_18577 (I318317,I2507,I317797,I317786,);
not I_18578 (I318375,I2514);
DFFARX1 I_18579 (I555956,I2507,I318375,I318401,);
not I_18580 (I318409,I318401);
DFFARX1 I_18581 (I555947,I2507,I318375,I318435,);
not I_18582 (I318443,I555941);
nand I_18583 (I318460,I318443,I555953);
not I_18584 (I318477,I318460);
nor I_18585 (I318494,I318477,I555944);
nor I_18586 (I318511,I318409,I318494);
DFFARX1 I_18587 (I318511,I2507,I318375,I318361,);
not I_18588 (I318542,I555944);
nand I_18589 (I318559,I318542,I318477);
and I_18590 (I318576,I318542,I555950);
nand I_18591 (I318593,I318576,I555935);
nor I_18592 (I318358,I318593,I318542);
and I_18593 (I318349,I318435,I318593);
not I_18594 (I318638,I318593);
nand I_18595 (I318352,I318435,I318638);
nor I_18596 (I318346,I318401,I318593);
not I_18597 (I318683,I555935);
nor I_18598 (I318700,I318683,I555950);
nand I_18599 (I318717,I318700,I318542);
nor I_18600 (I318355,I318460,I318717);
nor I_18601 (I318748,I318683,I555938);
and I_18602 (I318765,I318748,I555941);
or I_18603 (I318782,I318765,I555938);
DFFARX1 I_18604 (I318782,I2507,I318375,I318808,);
nor I_18605 (I318816,I318808,I318559);
DFFARX1 I_18606 (I318816,I2507,I318375,I318343,);
DFFARX1 I_18607 (I318808,I2507,I318375,I318367,);
not I_18608 (I318861,I318808);
nor I_18609 (I318878,I318861,I318435);
nor I_18610 (I318895,I318700,I318878);
DFFARX1 I_18611 (I318895,I2507,I318375,I318364,);
not I_18612 (I318953,I2514);
DFFARX1 I_18613 (I649623,I2507,I318953,I318979,);
not I_18614 (I318987,I318979);
DFFARX1 I_18615 (I649617,I2507,I318953,I319013,);
not I_18616 (I319021,I649626);
nand I_18617 (I319038,I319021,I649605);
not I_18618 (I319055,I319038);
nor I_18619 (I319072,I319055,I649614);
nor I_18620 (I319089,I318987,I319072);
DFFARX1 I_18621 (I319089,I2507,I318953,I318939,);
not I_18622 (I319120,I649614);
nand I_18623 (I319137,I319120,I319055);
and I_18624 (I319154,I319120,I649629);
nand I_18625 (I319171,I319154,I649608);
nor I_18626 (I318936,I319171,I319120);
and I_18627 (I318927,I319013,I319171);
not I_18628 (I319216,I319171);
nand I_18629 (I318930,I319013,I319216);
nor I_18630 (I318924,I318979,I319171);
not I_18631 (I319261,I649611);
nor I_18632 (I319278,I319261,I649629);
nand I_18633 (I319295,I319278,I319120);
nor I_18634 (I318933,I319038,I319295);
nor I_18635 (I319326,I319261,I649620);
and I_18636 (I319343,I319326,I649608);
or I_18637 (I319360,I319343,I649605);
DFFARX1 I_18638 (I319360,I2507,I318953,I319386,);
nor I_18639 (I319394,I319386,I319137);
DFFARX1 I_18640 (I319394,I2507,I318953,I318921,);
DFFARX1 I_18641 (I319386,I2507,I318953,I318945,);
not I_18642 (I319439,I319386);
nor I_18643 (I319456,I319439,I319013);
nor I_18644 (I319473,I319278,I319456);
DFFARX1 I_18645 (I319473,I2507,I318953,I318942,);
not I_18646 (I319531,I2514);
DFFARX1 I_18647 (I552590,I2507,I319531,I319557,);
not I_18648 (I319565,I319557);
DFFARX1 I_18649 (I552581,I2507,I319531,I319591,);
not I_18650 (I319599,I552575);
nand I_18651 (I319616,I319599,I552587);
not I_18652 (I319633,I319616);
nor I_18653 (I319650,I319633,I552578);
nor I_18654 (I319667,I319565,I319650);
DFFARX1 I_18655 (I319667,I2507,I319531,I319517,);
not I_18656 (I319698,I552578);
nand I_18657 (I319715,I319698,I319633);
and I_18658 (I319732,I319698,I552584);
nand I_18659 (I319749,I319732,I552569);
nor I_18660 (I319514,I319749,I319698);
and I_18661 (I319505,I319591,I319749);
not I_18662 (I319794,I319749);
nand I_18663 (I319508,I319591,I319794);
nor I_18664 (I319502,I319557,I319749);
not I_18665 (I319839,I552569);
nor I_18666 (I319856,I319839,I552584);
nand I_18667 (I319873,I319856,I319698);
nor I_18668 (I319511,I319616,I319873);
nor I_18669 (I319904,I319839,I552572);
and I_18670 (I319921,I319904,I552575);
or I_18671 (I319938,I319921,I552572);
DFFARX1 I_18672 (I319938,I2507,I319531,I319964,);
nor I_18673 (I319972,I319964,I319715);
DFFARX1 I_18674 (I319972,I2507,I319531,I319499,);
DFFARX1 I_18675 (I319964,I2507,I319531,I319523,);
not I_18676 (I320017,I319964);
nor I_18677 (I320034,I320017,I319591);
nor I_18678 (I320051,I319856,I320034);
DFFARX1 I_18679 (I320051,I2507,I319531,I319520,);
not I_18680 (I320109,I2514);
DFFARX1 I_18681 (I421227,I2507,I320109,I320135,);
not I_18682 (I320143,I320135);
DFFARX1 I_18683 (I421239,I2507,I320109,I320169,);
not I_18684 (I320177,I421230);
nand I_18685 (I320194,I320177,I421233);
not I_18686 (I320211,I320194);
nor I_18687 (I320228,I320211,I421236);
nor I_18688 (I320245,I320143,I320228);
DFFARX1 I_18689 (I320245,I2507,I320109,I320095,);
not I_18690 (I320276,I421236);
nand I_18691 (I320293,I320276,I320211);
and I_18692 (I320310,I320276,I421230);
nand I_18693 (I320327,I320310,I421242);
nor I_18694 (I320092,I320327,I320276);
and I_18695 (I320083,I320169,I320327);
not I_18696 (I320372,I320327);
nand I_18697 (I320086,I320169,I320372);
nor I_18698 (I320080,I320135,I320327);
not I_18699 (I320417,I421248);
nor I_18700 (I320434,I320417,I421230);
nand I_18701 (I320451,I320434,I320276);
nor I_18702 (I320089,I320194,I320451);
nor I_18703 (I320482,I320417,I421227);
and I_18704 (I320499,I320482,I421245);
or I_18705 (I320516,I320499,I421251);
DFFARX1 I_18706 (I320516,I2507,I320109,I320542,);
nor I_18707 (I320550,I320542,I320293);
DFFARX1 I_18708 (I320550,I2507,I320109,I320077,);
DFFARX1 I_18709 (I320542,I2507,I320109,I320101,);
not I_18710 (I320595,I320542);
nor I_18711 (I320612,I320595,I320169);
nor I_18712 (I320629,I320434,I320612);
DFFARX1 I_18713 (I320629,I2507,I320109,I320098,);
not I_18714 (I320687,I2514);
DFFARX1 I_18715 (I137189,I2507,I320687,I320713,);
not I_18716 (I320721,I320713);
DFFARX1 I_18717 (I137174,I2507,I320687,I320747,);
not I_18718 (I320755,I137192);
nand I_18719 (I320772,I320755,I137177);
not I_18720 (I320789,I320772);
nor I_18721 (I320806,I320789,I137174);
nor I_18722 (I320823,I320721,I320806);
DFFARX1 I_18723 (I320823,I2507,I320687,I320673,);
not I_18724 (I320854,I137174);
nand I_18725 (I320871,I320854,I320789);
and I_18726 (I320888,I320854,I137177);
nand I_18727 (I320905,I320888,I137198);
nor I_18728 (I320670,I320905,I320854);
and I_18729 (I320661,I320747,I320905);
not I_18730 (I320950,I320905);
nand I_18731 (I320664,I320747,I320950);
nor I_18732 (I320658,I320713,I320905);
not I_18733 (I320995,I137186);
nor I_18734 (I321012,I320995,I137177);
nand I_18735 (I321029,I321012,I320854);
nor I_18736 (I320667,I320772,I321029);
nor I_18737 (I321060,I320995,I137180);
and I_18738 (I321077,I321060,I137195);
or I_18739 (I321094,I321077,I137183);
DFFARX1 I_18740 (I321094,I2507,I320687,I321120,);
nor I_18741 (I321128,I321120,I320871);
DFFARX1 I_18742 (I321128,I2507,I320687,I320655,);
DFFARX1 I_18743 (I321120,I2507,I320687,I320679,);
not I_18744 (I321173,I321120);
nor I_18745 (I321190,I321173,I320747);
nor I_18746 (I321207,I321012,I321190);
DFFARX1 I_18747 (I321207,I2507,I320687,I320676,);
not I_18748 (I321265,I2514);
DFFARX1 I_18749 (I539687,I2507,I321265,I321291,);
not I_18750 (I321299,I321291);
DFFARX1 I_18751 (I539678,I2507,I321265,I321325,);
not I_18752 (I321333,I539672);
nand I_18753 (I321350,I321333,I539684);
not I_18754 (I321367,I321350);
nor I_18755 (I321384,I321367,I539675);
nor I_18756 (I321401,I321299,I321384);
DFFARX1 I_18757 (I321401,I2507,I321265,I321251,);
not I_18758 (I321432,I539675);
nand I_18759 (I321449,I321432,I321367);
and I_18760 (I321466,I321432,I539681);
nand I_18761 (I321483,I321466,I539666);
nor I_18762 (I321248,I321483,I321432);
and I_18763 (I321239,I321325,I321483);
not I_18764 (I321528,I321483);
nand I_18765 (I321242,I321325,I321528);
nor I_18766 (I321236,I321291,I321483);
not I_18767 (I321573,I539666);
nor I_18768 (I321590,I321573,I539681);
nand I_18769 (I321607,I321590,I321432);
nor I_18770 (I321245,I321350,I321607);
nor I_18771 (I321638,I321573,I539669);
and I_18772 (I321655,I321638,I539672);
or I_18773 (I321672,I321655,I539669);
DFFARX1 I_18774 (I321672,I2507,I321265,I321698,);
nor I_18775 (I321706,I321698,I321449);
DFFARX1 I_18776 (I321706,I2507,I321265,I321233,);
DFFARX1 I_18777 (I321698,I2507,I321265,I321257,);
not I_18778 (I321751,I321698);
nor I_18779 (I321768,I321751,I321325);
nor I_18780 (I321785,I321590,I321768);
DFFARX1 I_18781 (I321785,I2507,I321265,I321254,);
not I_18782 (I321843,I2514);
DFFARX1 I_18783 (I496390,I2507,I321843,I321869,);
not I_18784 (I321877,I321869);
DFFARX1 I_18785 (I496387,I2507,I321843,I321903,);
not I_18786 (I321911,I496384);
nand I_18787 (I321928,I321911,I496411);
not I_18788 (I321945,I321928);
nor I_18789 (I321962,I321945,I496399);
nor I_18790 (I321979,I321877,I321962);
DFFARX1 I_18791 (I321979,I2507,I321843,I321829,);
not I_18792 (I322010,I496399);
nand I_18793 (I322027,I322010,I321945);
and I_18794 (I322044,I322010,I496405);
nand I_18795 (I322061,I322044,I496396);
nor I_18796 (I321826,I322061,I322010);
and I_18797 (I321817,I321903,I322061);
not I_18798 (I322106,I322061);
nand I_18799 (I321820,I321903,I322106);
nor I_18800 (I321814,I321869,I322061);
not I_18801 (I322151,I496393);
nor I_18802 (I322168,I322151,I496405);
nand I_18803 (I322185,I322168,I322010);
nor I_18804 (I321823,I321928,I322185);
nor I_18805 (I322216,I322151,I496408);
and I_18806 (I322233,I322216,I496402);
or I_18807 (I322250,I322233,I496384);
DFFARX1 I_18808 (I322250,I2507,I321843,I322276,);
nor I_18809 (I322284,I322276,I322027);
DFFARX1 I_18810 (I322284,I2507,I321843,I321811,);
DFFARX1 I_18811 (I322276,I2507,I321843,I321835,);
not I_18812 (I322329,I322276);
nor I_18813 (I322346,I322329,I321903);
nor I_18814 (I322363,I322168,I322346);
DFFARX1 I_18815 (I322363,I2507,I321843,I321832,);
not I_18816 (I322421,I2514);
DFFARX1 I_18817 (I619651,I2507,I322421,I322447,);
not I_18818 (I322455,I322447);
DFFARX1 I_18819 (I619657,I2507,I322421,I322481,);
not I_18820 (I322489,I619651);
nand I_18821 (I322506,I322489,I619654);
not I_18822 (I322523,I322506);
nor I_18823 (I322540,I322523,I619672);
nor I_18824 (I322557,I322455,I322540);
DFFARX1 I_18825 (I322557,I2507,I322421,I322407,);
not I_18826 (I322588,I619672);
nand I_18827 (I322605,I322588,I322523);
and I_18828 (I322622,I322588,I619675);
nand I_18829 (I322639,I322622,I619654);
nor I_18830 (I322404,I322639,I322588);
and I_18831 (I322395,I322481,I322639);
not I_18832 (I322684,I322639);
nand I_18833 (I322398,I322481,I322684);
nor I_18834 (I322392,I322447,I322639);
not I_18835 (I322729,I619660);
nor I_18836 (I322746,I322729,I619675);
nand I_18837 (I322763,I322746,I322588);
nor I_18838 (I322401,I322506,I322763);
nor I_18839 (I322794,I322729,I619666);
and I_18840 (I322811,I322794,I619663);
or I_18841 (I322828,I322811,I619669);
DFFARX1 I_18842 (I322828,I2507,I322421,I322854,);
nor I_18843 (I322862,I322854,I322605);
DFFARX1 I_18844 (I322862,I2507,I322421,I322389,);
DFFARX1 I_18845 (I322854,I2507,I322421,I322413,);
not I_18846 (I322907,I322854);
nor I_18847 (I322924,I322907,I322481);
nor I_18848 (I322941,I322746,I322924);
DFFARX1 I_18849 (I322941,I2507,I322421,I322410,);
not I_18850 (I322999,I2514);
DFFARX1 I_18851 (I147304,I2507,I322999,I323025,);
not I_18852 (I323033,I323025);
DFFARX1 I_18853 (I147289,I2507,I322999,I323059,);
not I_18854 (I323067,I147307);
nand I_18855 (I323084,I323067,I147292);
not I_18856 (I323101,I323084);
nor I_18857 (I323118,I323101,I147289);
nor I_18858 (I323135,I323033,I323118);
DFFARX1 I_18859 (I323135,I2507,I322999,I322985,);
not I_18860 (I323166,I147289);
nand I_18861 (I323183,I323166,I323101);
and I_18862 (I323200,I323166,I147292);
nand I_18863 (I323217,I323200,I147313);
nor I_18864 (I322982,I323217,I323166);
and I_18865 (I322973,I323059,I323217);
not I_18866 (I323262,I323217);
nand I_18867 (I322976,I323059,I323262);
nor I_18868 (I322970,I323025,I323217);
not I_18869 (I323307,I147301);
nor I_18870 (I323324,I323307,I147292);
nand I_18871 (I323341,I323324,I323166);
nor I_18872 (I322979,I323084,I323341);
nor I_18873 (I323372,I323307,I147295);
and I_18874 (I323389,I323372,I147310);
or I_18875 (I323406,I323389,I147298);
DFFARX1 I_18876 (I323406,I2507,I322999,I323432,);
nor I_18877 (I323440,I323432,I323183);
DFFARX1 I_18878 (I323440,I2507,I322999,I322967,);
DFFARX1 I_18879 (I323432,I2507,I322999,I322991,);
not I_18880 (I323485,I323432);
nor I_18881 (I323502,I323485,I323059);
nor I_18882 (I323519,I323324,I323502);
DFFARX1 I_18883 (I323519,I2507,I322999,I322988,);
not I_18884 (I323577,I2514);
DFFARX1 I_18885 (I273220,I2507,I323577,I323603,);
not I_18886 (I323611,I323603);
DFFARX1 I_18887 (I273232,I2507,I323577,I323637,);
not I_18888 (I323645,I273208);
nand I_18889 (I323662,I323645,I273235);
not I_18890 (I323679,I323662);
nor I_18891 (I323696,I323679,I273223);
nor I_18892 (I323713,I323611,I323696);
DFFARX1 I_18893 (I323713,I2507,I323577,I323563,);
not I_18894 (I323744,I273223);
nand I_18895 (I323761,I323744,I323679);
and I_18896 (I323778,I323744,I273208);
nand I_18897 (I323795,I323778,I273211);
nor I_18898 (I323560,I323795,I323744);
and I_18899 (I323551,I323637,I323795);
not I_18900 (I323840,I323795);
nand I_18901 (I323554,I323637,I323840);
nor I_18902 (I323548,I323603,I323795);
not I_18903 (I323885,I273217);
nor I_18904 (I323902,I323885,I273208);
nand I_18905 (I323919,I323902,I323744);
nor I_18906 (I323557,I323662,I323919);
nor I_18907 (I323950,I323885,I273226);
and I_18908 (I323967,I323950,I273214);
or I_18909 (I323984,I323967,I273229);
DFFARX1 I_18910 (I323984,I2507,I323577,I324010,);
nor I_18911 (I324018,I324010,I323761);
DFFARX1 I_18912 (I324018,I2507,I323577,I323545,);
DFFARX1 I_18913 (I324010,I2507,I323577,I323569,);
not I_18914 (I324063,I324010);
nor I_18915 (I324080,I324063,I323637);
nor I_18916 (I324097,I323902,I324080);
DFFARX1 I_18917 (I324097,I2507,I323577,I323566,);
not I_18918 (I324155,I2514);
DFFARX1 I_18919 (I427591,I2507,I324155,I324181,);
not I_18920 (I324189,I324181);
DFFARX1 I_18921 (I427591,I2507,I324155,I324215,);
not I_18922 (I324223,I427588);
nand I_18923 (I324240,I324223,I427603);
not I_18924 (I324257,I324240);
nor I_18925 (I324274,I324257,I427597);
nor I_18926 (I324291,I324189,I324274);
DFFARX1 I_18927 (I324291,I2507,I324155,I324141,);
not I_18928 (I324322,I427597);
nand I_18929 (I324339,I324322,I324257);
and I_18930 (I324356,I324322,I427594);
nand I_18931 (I324373,I324356,I427585);
nor I_18932 (I324138,I324373,I324322);
and I_18933 (I324129,I324215,I324373);
not I_18934 (I324418,I324373);
nand I_18935 (I324132,I324215,I324418);
nor I_18936 (I324126,I324181,I324373);
not I_18937 (I324463,I427606);
nor I_18938 (I324480,I324463,I427594);
nand I_18939 (I324497,I324480,I324322);
nor I_18940 (I324135,I324240,I324497);
nor I_18941 (I324528,I324463,I427585);
and I_18942 (I324545,I324528,I427588);
or I_18943 (I324562,I324545,I427600);
DFFARX1 I_18944 (I324562,I2507,I324155,I324588,);
nor I_18945 (I324596,I324588,I324339);
DFFARX1 I_18946 (I324596,I2507,I324155,I324123,);
DFFARX1 I_18947 (I324588,I2507,I324155,I324147,);
not I_18948 (I324641,I324588);
nor I_18949 (I324658,I324641,I324215);
nor I_18950 (I324675,I324480,I324658);
DFFARX1 I_18951 (I324675,I2507,I324155,I324144,);
not I_18952 (I324733,I2514);
DFFARX1 I_18953 (I375565,I2507,I324733,I324759,);
not I_18954 (I324767,I324759);
DFFARX1 I_18955 (I375577,I2507,I324733,I324793,);
not I_18956 (I324801,I375568);
nand I_18957 (I324818,I324801,I375571);
not I_18958 (I324835,I324818);
nor I_18959 (I324852,I324835,I375574);
nor I_18960 (I324869,I324767,I324852);
DFFARX1 I_18961 (I324869,I2507,I324733,I324719,);
not I_18962 (I324900,I375574);
nand I_18963 (I324917,I324900,I324835);
and I_18964 (I324934,I324900,I375568);
nand I_18965 (I324951,I324934,I375580);
nor I_18966 (I324716,I324951,I324900);
and I_18967 (I324707,I324793,I324951);
not I_18968 (I324996,I324951);
nand I_18969 (I324710,I324793,I324996);
nor I_18970 (I324704,I324759,I324951);
not I_18971 (I325041,I375586);
nor I_18972 (I325058,I325041,I375568);
nand I_18973 (I325075,I325058,I324900);
nor I_18974 (I324713,I324818,I325075);
nor I_18975 (I325106,I325041,I375565);
and I_18976 (I325123,I325106,I375583);
or I_18977 (I325140,I325123,I375589);
DFFARX1 I_18978 (I325140,I2507,I324733,I325166,);
nor I_18979 (I325174,I325166,I324917);
DFFARX1 I_18980 (I325174,I2507,I324733,I324701,);
DFFARX1 I_18981 (I325166,I2507,I324733,I324725,);
not I_18982 (I325219,I325166);
nor I_18983 (I325236,I325219,I324793);
nor I_18984 (I325253,I325058,I325236);
DFFARX1 I_18985 (I325253,I2507,I324733,I324722,);
not I_18986 (I325311,I2514);
DFFARX1 I_18987 (I93159,I2507,I325311,I325337,);
not I_18988 (I325345,I325337);
DFFARX1 I_18989 (I93144,I2507,I325311,I325371,);
not I_18990 (I325379,I93162);
nand I_18991 (I325396,I325379,I93147);
not I_18992 (I325413,I325396);
nor I_18993 (I325430,I325413,I93144);
nor I_18994 (I325447,I325345,I325430);
DFFARX1 I_18995 (I325447,I2507,I325311,I325297,);
not I_18996 (I325478,I93144);
nand I_18997 (I325495,I325478,I325413);
and I_18998 (I325512,I325478,I93147);
nand I_18999 (I325529,I325512,I93168);
nor I_19000 (I325294,I325529,I325478);
and I_19001 (I325285,I325371,I325529);
not I_19002 (I325574,I325529);
nand I_19003 (I325288,I325371,I325574);
nor I_19004 (I325282,I325337,I325529);
not I_19005 (I325619,I93156);
nor I_19006 (I325636,I325619,I93147);
nand I_19007 (I325653,I325636,I325478);
nor I_19008 (I325291,I325396,I325653);
nor I_19009 (I325684,I325619,I93150);
and I_19010 (I325701,I325684,I93165);
or I_19011 (I325718,I325701,I93153);
DFFARX1 I_19012 (I325718,I2507,I325311,I325744,);
nor I_19013 (I325752,I325744,I325495);
DFFARX1 I_19014 (I325752,I2507,I325311,I325279,);
DFFARX1 I_19015 (I325744,I2507,I325311,I325303,);
not I_19016 (I325797,I325744);
nor I_19017 (I325814,I325797,I325371);
nor I_19018 (I325831,I325636,I325814);
DFFARX1 I_19019 (I325831,I2507,I325311,I325300,);
not I_19020 (I325889,I2514);
DFFARX1 I_19021 (I541931,I2507,I325889,I325915,);
not I_19022 (I325923,I325915);
DFFARX1 I_19023 (I541922,I2507,I325889,I325949,);
not I_19024 (I325957,I541916);
nand I_19025 (I325974,I325957,I541928);
not I_19026 (I325991,I325974);
nor I_19027 (I326008,I325991,I541919);
nor I_19028 (I326025,I325923,I326008);
DFFARX1 I_19029 (I326025,I2507,I325889,I325875,);
not I_19030 (I326056,I541919);
nand I_19031 (I326073,I326056,I325991);
and I_19032 (I326090,I326056,I541925);
nand I_19033 (I326107,I326090,I541910);
nor I_19034 (I325872,I326107,I326056);
and I_19035 (I325863,I325949,I326107);
not I_19036 (I326152,I326107);
nand I_19037 (I325866,I325949,I326152);
nor I_19038 (I325860,I325915,I326107);
not I_19039 (I326197,I541910);
nor I_19040 (I326214,I326197,I541925);
nand I_19041 (I326231,I326214,I326056);
nor I_19042 (I325869,I325974,I326231);
nor I_19043 (I326262,I326197,I541913);
and I_19044 (I326279,I326262,I541916);
or I_19045 (I326296,I326279,I541913);
DFFARX1 I_19046 (I326296,I2507,I325889,I326322,);
nor I_19047 (I326330,I326322,I326073);
DFFARX1 I_19048 (I326330,I2507,I325889,I325857,);
DFFARX1 I_19049 (I326322,I2507,I325889,I325881,);
not I_19050 (I326375,I326322);
nor I_19051 (I326392,I326375,I325949);
nor I_19052 (I326409,I326214,I326392);
DFFARX1 I_19053 (I326409,I2507,I325889,I325878,);
not I_19054 (I326467,I2514);
DFFARX1 I_19055 (I6685,I2507,I326467,I326493,);
not I_19056 (I326501,I326493);
DFFARX1 I_19057 (I6688,I2507,I326467,I326527,);
not I_19058 (I326535,I6682);
nand I_19059 (I326552,I326535,I6706);
not I_19060 (I326569,I326552);
nor I_19061 (I326586,I326569,I6685);
nor I_19062 (I326603,I326501,I326586);
DFFARX1 I_19063 (I326603,I2507,I326467,I326453,);
not I_19064 (I326634,I6685);
nand I_19065 (I326651,I326634,I326569);
and I_19066 (I326668,I326634,I6700);
nand I_19067 (I326685,I326668,I6694);
nor I_19068 (I326450,I326685,I326634);
and I_19069 (I326441,I326527,I326685);
not I_19070 (I326730,I326685);
nand I_19071 (I326444,I326527,I326730);
nor I_19072 (I326438,I326493,I326685);
not I_19073 (I326775,I6703);
nor I_19074 (I326792,I326775,I6700);
nand I_19075 (I326809,I326792,I326634);
nor I_19076 (I326447,I326552,I326809);
nor I_19077 (I326840,I326775,I6682);
and I_19078 (I326857,I326840,I6691);
or I_19079 (I326874,I326857,I6697);
DFFARX1 I_19080 (I326874,I2507,I326467,I326900,);
nor I_19081 (I326908,I326900,I326651);
DFFARX1 I_19082 (I326908,I2507,I326467,I326435,);
DFFARX1 I_19083 (I326900,I2507,I326467,I326459,);
not I_19084 (I326953,I326900);
nor I_19085 (I326970,I326953,I326527);
nor I_19086 (I326987,I326792,I326970);
DFFARX1 I_19087 (I326987,I2507,I326467,I326456,);
not I_19088 (I327045,I2514);
DFFARX1 I_19089 (I187466,I2507,I327045,I327071,);
not I_19090 (I327079,I327071);
DFFARX1 I_19091 (I187481,I2507,I327045,I327105,);
not I_19092 (I327113,I187484);
nand I_19093 (I327130,I327113,I187463);
not I_19094 (I327147,I327130);
nor I_19095 (I327164,I327147,I187487);
nor I_19096 (I327181,I327079,I327164);
DFFARX1 I_19097 (I327181,I2507,I327045,I327031,);
not I_19098 (I327212,I187487);
nand I_19099 (I327229,I327212,I327147);
and I_19100 (I327246,I327212,I187469);
nand I_19101 (I327263,I327246,I187460);
nor I_19102 (I327028,I327263,I327212);
and I_19103 (I327019,I327105,I327263);
not I_19104 (I327308,I327263);
nand I_19105 (I327022,I327105,I327308);
nor I_19106 (I327016,I327071,I327263);
not I_19107 (I327353,I187460);
nor I_19108 (I327370,I327353,I187469);
nand I_19109 (I327387,I327370,I327212);
nor I_19110 (I327025,I327130,I327387);
nor I_19111 (I327418,I327353,I187475);
and I_19112 (I327435,I327418,I187478);
or I_19113 (I327452,I327435,I187472);
DFFARX1 I_19114 (I327452,I2507,I327045,I327478,);
nor I_19115 (I327486,I327478,I327229);
DFFARX1 I_19116 (I327486,I2507,I327045,I327013,);
DFFARX1 I_19117 (I327478,I2507,I327045,I327037,);
not I_19118 (I327531,I327478);
nor I_19119 (I327548,I327531,I327105);
nor I_19120 (I327565,I327370,I327548);
DFFARX1 I_19121 (I327565,I2507,I327045,I327034,);
not I_19122 (I327623,I2514);
DFFARX1 I_19123 (I160394,I2507,I327623,I327649,);
not I_19124 (I327657,I327649);
DFFARX1 I_19125 (I160379,I2507,I327623,I327683,);
not I_19126 (I327691,I160397);
nand I_19127 (I327708,I327691,I160382);
not I_19128 (I327725,I327708);
nor I_19129 (I327742,I327725,I160379);
nor I_19130 (I327759,I327657,I327742);
DFFARX1 I_19131 (I327759,I2507,I327623,I327609,);
not I_19132 (I327790,I160379);
nand I_19133 (I327807,I327790,I327725);
and I_19134 (I327824,I327790,I160382);
nand I_19135 (I327841,I327824,I160403);
nor I_19136 (I327606,I327841,I327790);
and I_19137 (I327597,I327683,I327841);
not I_19138 (I327886,I327841);
nand I_19139 (I327600,I327683,I327886);
nor I_19140 (I327594,I327649,I327841);
not I_19141 (I327931,I160391);
nor I_19142 (I327948,I327931,I160382);
nand I_19143 (I327965,I327948,I327790);
nor I_19144 (I327603,I327708,I327965);
nor I_19145 (I327996,I327931,I160385);
and I_19146 (I328013,I327996,I160400);
or I_19147 (I328030,I328013,I160388);
DFFARX1 I_19148 (I328030,I2507,I327623,I328056,);
nor I_19149 (I328064,I328056,I327807);
DFFARX1 I_19150 (I328064,I2507,I327623,I327591,);
DFFARX1 I_19151 (I328056,I2507,I327623,I327615,);
not I_19152 (I328109,I328056);
nor I_19153 (I328126,I328109,I327683);
nor I_19154 (I328143,I327948,I328126);
DFFARX1 I_19155 (I328143,I2507,I327623,I327612,);
not I_19156 (I328201,I2514);
DFFARX1 I_19157 (I698973,I2507,I328201,I328227,);
not I_19158 (I328235,I328227);
DFFARX1 I_19159 (I698973,I2507,I328201,I328261,);
not I_19160 (I328269,I698997);
nand I_19161 (I328286,I328269,I698979);
not I_19162 (I328303,I328286);
nor I_19163 (I328320,I328303,I698994);
nor I_19164 (I328337,I328235,I328320);
DFFARX1 I_19165 (I328337,I2507,I328201,I328187,);
not I_19166 (I328368,I698994);
nand I_19167 (I328385,I328368,I328303);
and I_19168 (I328402,I328368,I698976);
nand I_19169 (I328419,I328402,I698985);
nor I_19170 (I328184,I328419,I328368);
and I_19171 (I328175,I328261,I328419);
not I_19172 (I328464,I328419);
nand I_19173 (I328178,I328261,I328464);
nor I_19174 (I328172,I328227,I328419);
not I_19175 (I328509,I698982);
nor I_19176 (I328526,I328509,I698976);
nand I_19177 (I328543,I328526,I328368);
nor I_19178 (I328181,I328286,I328543);
nor I_19179 (I328574,I328509,I698991);
and I_19180 (I328591,I328574,I699000);
or I_19181 (I328608,I328591,I698988);
DFFARX1 I_19182 (I328608,I2507,I328201,I328634,);
nor I_19183 (I328642,I328634,I328385);
DFFARX1 I_19184 (I328642,I2507,I328201,I328169,);
DFFARX1 I_19185 (I328634,I2507,I328201,I328193,);
not I_19186 (I328687,I328634);
nor I_19187 (I328704,I328687,I328261);
nor I_19188 (I328721,I328526,I328704);
DFFARX1 I_19189 (I328721,I2507,I328201,I328190,);
not I_19190 (I328779,I2514);
DFFARX1 I_19191 (I544736,I2507,I328779,I328805,);
not I_19192 (I328813,I328805);
DFFARX1 I_19193 (I544727,I2507,I328779,I328839,);
not I_19194 (I328847,I544721);
nand I_19195 (I328864,I328847,I544733);
not I_19196 (I328881,I328864);
nor I_19197 (I328898,I328881,I544724);
nor I_19198 (I328915,I328813,I328898);
DFFARX1 I_19199 (I328915,I2507,I328779,I328765,);
not I_19200 (I328946,I544724);
nand I_19201 (I328963,I328946,I328881);
and I_19202 (I328980,I328946,I544730);
nand I_19203 (I328997,I328980,I544715);
nor I_19204 (I328762,I328997,I328946);
and I_19205 (I328753,I328839,I328997);
not I_19206 (I329042,I328997);
nand I_19207 (I328756,I328839,I329042);
nor I_19208 (I328750,I328805,I328997);
not I_19209 (I329087,I544715);
nor I_19210 (I329104,I329087,I544730);
nand I_19211 (I329121,I329104,I328946);
nor I_19212 (I328759,I328864,I329121);
nor I_19213 (I329152,I329087,I544718);
and I_19214 (I329169,I329152,I544721);
or I_19215 (I329186,I329169,I544718);
DFFARX1 I_19216 (I329186,I2507,I328779,I329212,);
nor I_19217 (I329220,I329212,I328963);
DFFARX1 I_19218 (I329220,I2507,I328779,I328747,);
DFFARX1 I_19219 (I329212,I2507,I328779,I328771,);
not I_19220 (I329265,I329212);
nor I_19221 (I329282,I329265,I328839);
nor I_19222 (I329299,I329104,I329282);
DFFARX1 I_19223 (I329299,I2507,I328779,I328768,);
not I_19224 (I329357,I2514);
DFFARX1 I_19225 (I671139,I2507,I329357,I329383,);
not I_19226 (I329391,I329383);
DFFARX1 I_19227 (I671151,I2507,I329357,I329417,);
not I_19228 (I329425,I671142);
nand I_19229 (I329442,I329425,I671130);
not I_19230 (I329459,I329442);
nor I_19231 (I329476,I329459,I671127);
nor I_19232 (I329493,I329391,I329476);
DFFARX1 I_19233 (I329493,I2507,I329357,I329343,);
not I_19234 (I329524,I671127);
nand I_19235 (I329541,I329524,I329459);
and I_19236 (I329558,I329524,I671133);
nand I_19237 (I329575,I329558,I671130);
nor I_19238 (I329340,I329575,I329524);
and I_19239 (I329331,I329417,I329575);
not I_19240 (I329620,I329575);
nand I_19241 (I329334,I329417,I329620);
nor I_19242 (I329328,I329383,I329575);
not I_19243 (I329665,I671148);
nor I_19244 (I329682,I329665,I671133);
nand I_19245 (I329699,I329682,I329524);
nor I_19246 (I329337,I329442,I329699);
nor I_19247 (I329730,I329665,I671136);
and I_19248 (I329747,I329730,I671127);
or I_19249 (I329764,I329747,I671145);
DFFARX1 I_19250 (I329764,I2507,I329357,I329790,);
nor I_19251 (I329798,I329790,I329541);
DFFARX1 I_19252 (I329798,I2507,I329357,I329325,);
DFFARX1 I_19253 (I329790,I2507,I329357,I329349,);
not I_19254 (I329843,I329790);
nor I_19255 (I329860,I329843,I329417);
nor I_19256 (I329877,I329682,I329860);
DFFARX1 I_19257 (I329877,I2507,I329357,I329346,);
not I_19258 (I329935,I2514);
DFFARX1 I_19259 (I357069,I2507,I329935,I329961,);
not I_19260 (I329969,I329961);
DFFARX1 I_19261 (I357081,I2507,I329935,I329995,);
not I_19262 (I330003,I357072);
nand I_19263 (I330020,I330003,I357075);
not I_19264 (I330037,I330020);
nor I_19265 (I330054,I330037,I357078);
nor I_19266 (I330071,I329969,I330054);
DFFARX1 I_19267 (I330071,I2507,I329935,I329921,);
not I_19268 (I330102,I357078);
nand I_19269 (I330119,I330102,I330037);
and I_19270 (I330136,I330102,I357072);
nand I_19271 (I330153,I330136,I357084);
nor I_19272 (I329918,I330153,I330102);
and I_19273 (I329909,I329995,I330153);
not I_19274 (I330198,I330153);
nand I_19275 (I329912,I329995,I330198);
nor I_19276 (I329906,I329961,I330153);
not I_19277 (I330243,I357090);
nor I_19278 (I330260,I330243,I357072);
nand I_19279 (I330277,I330260,I330102);
nor I_19280 (I329915,I330020,I330277);
nor I_19281 (I330308,I330243,I357069);
and I_19282 (I330325,I330308,I357087);
or I_19283 (I330342,I330325,I357093);
DFFARX1 I_19284 (I330342,I2507,I329935,I330368,);
nor I_19285 (I330376,I330368,I330119);
DFFARX1 I_19286 (I330376,I2507,I329935,I329903,);
DFFARX1 I_19287 (I330368,I2507,I329935,I329927,);
not I_19288 (I330421,I330368);
nor I_19289 (I330438,I330421,I329995);
nor I_19290 (I330455,I330260,I330438);
DFFARX1 I_19291 (I330455,I2507,I329935,I329924,);
not I_19292 (I330513,I2514);
DFFARX1 I_19293 (I193263,I2507,I330513,I330539,);
not I_19294 (I330547,I330539);
DFFARX1 I_19295 (I193278,I2507,I330513,I330573,);
not I_19296 (I330581,I193281);
nand I_19297 (I330598,I330581,I193260);
not I_19298 (I330615,I330598);
nor I_19299 (I330632,I330615,I193284);
nor I_19300 (I330649,I330547,I330632);
DFFARX1 I_19301 (I330649,I2507,I330513,I330499,);
not I_19302 (I330680,I193284);
nand I_19303 (I330697,I330680,I330615);
and I_19304 (I330714,I330680,I193266);
nand I_19305 (I330731,I330714,I193257);
nor I_19306 (I330496,I330731,I330680);
and I_19307 (I330487,I330573,I330731);
not I_19308 (I330776,I330731);
nand I_19309 (I330490,I330573,I330776);
nor I_19310 (I330484,I330539,I330731);
not I_19311 (I330821,I193257);
nor I_19312 (I330838,I330821,I193266);
nand I_19313 (I330855,I330838,I330680);
nor I_19314 (I330493,I330598,I330855);
nor I_19315 (I330886,I330821,I193272);
and I_19316 (I330903,I330886,I193275);
or I_19317 (I330920,I330903,I193269);
DFFARX1 I_19318 (I330920,I2507,I330513,I330946,);
nor I_19319 (I330954,I330946,I330697);
DFFARX1 I_19320 (I330954,I2507,I330513,I330481,);
DFFARX1 I_19321 (I330946,I2507,I330513,I330505,);
not I_19322 (I330999,I330946);
nor I_19323 (I331016,I330999,I330573);
nor I_19324 (I331033,I330838,I331016);
DFFARX1 I_19325 (I331033,I2507,I330513,I330502,);
not I_19326 (I331091,I2514);
DFFARX1 I_19327 (I235684,I2507,I331091,I331117,);
not I_19328 (I331125,I331117);
DFFARX1 I_19329 (I235696,I2507,I331091,I331151,);
not I_19330 (I331159,I235672);
nand I_19331 (I331176,I331159,I235699);
not I_19332 (I331193,I331176);
nor I_19333 (I331210,I331193,I235687);
nor I_19334 (I331227,I331125,I331210);
DFFARX1 I_19335 (I331227,I2507,I331091,I331077,);
not I_19336 (I331258,I235687);
nand I_19337 (I331275,I331258,I331193);
and I_19338 (I331292,I331258,I235672);
nand I_19339 (I331309,I331292,I235675);
nor I_19340 (I331074,I331309,I331258);
and I_19341 (I331065,I331151,I331309);
not I_19342 (I331354,I331309);
nand I_19343 (I331068,I331151,I331354);
nor I_19344 (I331062,I331117,I331309);
not I_19345 (I331399,I235681);
nor I_19346 (I331416,I331399,I235672);
nand I_19347 (I331433,I331416,I331258);
nor I_19348 (I331071,I331176,I331433);
nor I_19349 (I331464,I331399,I235690);
and I_19350 (I331481,I331464,I235678);
or I_19351 (I331498,I331481,I235693);
DFFARX1 I_19352 (I331498,I2507,I331091,I331524,);
nor I_19353 (I331532,I331524,I331275);
DFFARX1 I_19354 (I331532,I2507,I331091,I331059,);
DFFARX1 I_19355 (I331524,I2507,I331091,I331083,);
not I_19356 (I331577,I331524);
nor I_19357 (I331594,I331577,I331151);
nor I_19358 (I331611,I331416,I331594);
DFFARX1 I_19359 (I331611,I2507,I331091,I331080,);
not I_19360 (I331669,I2514);
DFFARX1 I_19361 (I502204,I2507,I331669,I331695,);
not I_19362 (I331703,I331695);
DFFARX1 I_19363 (I502201,I2507,I331669,I331729,);
not I_19364 (I331737,I502198);
nand I_19365 (I331754,I331737,I502225);
not I_19366 (I331771,I331754);
nor I_19367 (I331788,I331771,I502213);
nor I_19368 (I331805,I331703,I331788);
DFFARX1 I_19369 (I331805,I2507,I331669,I331655,);
not I_19370 (I331836,I502213);
nand I_19371 (I331853,I331836,I331771);
and I_19372 (I331870,I331836,I502219);
nand I_19373 (I331887,I331870,I502210);
nor I_19374 (I331652,I331887,I331836);
and I_19375 (I331643,I331729,I331887);
not I_19376 (I331932,I331887);
nand I_19377 (I331646,I331729,I331932);
nor I_19378 (I331640,I331695,I331887);
not I_19379 (I331977,I502207);
nor I_19380 (I331994,I331977,I502219);
nand I_19381 (I332011,I331994,I331836);
nor I_19382 (I331649,I331754,I332011);
nor I_19383 (I332042,I331977,I502222);
and I_19384 (I332059,I332042,I502216);
or I_19385 (I332076,I332059,I502198);
DFFARX1 I_19386 (I332076,I2507,I331669,I332102,);
nor I_19387 (I332110,I332102,I331853);
DFFARX1 I_19388 (I332110,I2507,I331669,I331637,);
DFFARX1 I_19389 (I332102,I2507,I331669,I331661,);
not I_19390 (I332155,I332102);
nor I_19391 (I332172,I332155,I331729);
nor I_19392 (I332189,I331994,I332172);
DFFARX1 I_19393 (I332189,I2507,I331669,I331658,);
not I_19394 (I332247,I2514);
DFFARX1 I_19395 (I447617,I2507,I332247,I332273,);
not I_19396 (I332281,I332273);
DFFARX1 I_19397 (I447617,I2507,I332247,I332307,);
not I_19398 (I332315,I447614);
nand I_19399 (I332332,I332315,I447629);
not I_19400 (I332349,I332332);
nor I_19401 (I332366,I332349,I447623);
nor I_19402 (I332383,I332281,I332366);
DFFARX1 I_19403 (I332383,I2507,I332247,I332233,);
not I_19404 (I332414,I447623);
nand I_19405 (I332431,I332414,I332349);
and I_19406 (I332448,I332414,I447620);
nand I_19407 (I332465,I332448,I447611);
nor I_19408 (I332230,I332465,I332414);
and I_19409 (I332221,I332307,I332465);
not I_19410 (I332510,I332465);
nand I_19411 (I332224,I332307,I332510);
nor I_19412 (I332218,I332273,I332465);
not I_19413 (I332555,I447632);
nor I_19414 (I332572,I332555,I447620);
nand I_19415 (I332589,I332572,I332414);
nor I_19416 (I332227,I332332,I332589);
nor I_19417 (I332620,I332555,I447611);
and I_19418 (I332637,I332620,I447614);
or I_19419 (I332654,I332637,I447626);
DFFARX1 I_19420 (I332654,I2507,I332247,I332680,);
nor I_19421 (I332688,I332680,I332431);
DFFARX1 I_19422 (I332688,I2507,I332247,I332215,);
DFFARX1 I_19423 (I332680,I2507,I332247,I332239,);
not I_19424 (I332733,I332680);
nor I_19425 (I332750,I332733,I332307);
nor I_19426 (I332767,I332572,I332750);
DFFARX1 I_19427 (I332767,I2507,I332247,I332236,);
not I_19428 (I332825,I2514);
DFFARX1 I_19429 (I574567,I2507,I332825,I332851,);
not I_19430 (I332859,I332851);
DFFARX1 I_19431 (I574573,I2507,I332825,I332885,);
not I_19432 (I332893,I574567);
nand I_19433 (I332910,I332893,I574570);
not I_19434 (I332927,I332910);
nor I_19435 (I332944,I332927,I574588);
nor I_19436 (I332961,I332859,I332944);
DFFARX1 I_19437 (I332961,I2507,I332825,I332811,);
not I_19438 (I332992,I574588);
nand I_19439 (I333009,I332992,I332927);
and I_19440 (I333026,I332992,I574591);
nand I_19441 (I333043,I333026,I574570);
nor I_19442 (I332808,I333043,I332992);
and I_19443 (I332799,I332885,I333043);
not I_19444 (I333088,I333043);
nand I_19445 (I332802,I332885,I333088);
nor I_19446 (I332796,I332851,I333043);
not I_19447 (I333133,I574576);
nor I_19448 (I333150,I333133,I574591);
nand I_19449 (I333167,I333150,I332992);
nor I_19450 (I332805,I332910,I333167);
nor I_19451 (I333198,I333133,I574582);
and I_19452 (I333215,I333198,I574579);
or I_19453 (I333232,I333215,I574585);
DFFARX1 I_19454 (I333232,I2507,I332825,I333258,);
nor I_19455 (I333266,I333258,I333009);
DFFARX1 I_19456 (I333266,I2507,I332825,I332793,);
DFFARX1 I_19457 (I333258,I2507,I332825,I332817,);
not I_19458 (I333311,I333258);
nor I_19459 (I333328,I333311,I332885);
nor I_19460 (I333345,I333150,I333328);
DFFARX1 I_19461 (I333345,I2507,I332825,I332814,);
not I_19462 (I333403,I2514);
DFFARX1 I_19463 (I430226,I2507,I333403,I333429,);
not I_19464 (I333437,I333429);
DFFARX1 I_19465 (I430226,I2507,I333403,I333463,);
not I_19466 (I333471,I430223);
nand I_19467 (I333488,I333471,I430238);
not I_19468 (I333505,I333488);
nor I_19469 (I333522,I333505,I430232);
nor I_19470 (I333539,I333437,I333522);
DFFARX1 I_19471 (I333539,I2507,I333403,I333389,);
not I_19472 (I333570,I430232);
nand I_19473 (I333587,I333570,I333505);
and I_19474 (I333604,I333570,I430229);
nand I_19475 (I333621,I333604,I430220);
nor I_19476 (I333386,I333621,I333570);
and I_19477 (I333377,I333463,I333621);
not I_19478 (I333666,I333621);
nand I_19479 (I333380,I333463,I333666);
nor I_19480 (I333374,I333429,I333621);
not I_19481 (I333711,I430241);
nor I_19482 (I333728,I333711,I430229);
nand I_19483 (I333745,I333728,I333570);
nor I_19484 (I333383,I333488,I333745);
nor I_19485 (I333776,I333711,I430220);
and I_19486 (I333793,I333776,I430223);
or I_19487 (I333810,I333793,I430235);
DFFARX1 I_19488 (I333810,I2507,I333403,I333836,);
nor I_19489 (I333844,I333836,I333587);
DFFARX1 I_19490 (I333844,I2507,I333403,I333371,);
DFFARX1 I_19491 (I333836,I2507,I333403,I333395,);
not I_19492 (I333889,I333836);
nor I_19493 (I333906,I333889,I333463);
nor I_19494 (I333923,I333728,I333906);
DFFARX1 I_19495 (I333923,I2507,I333403,I333392,);
not I_19496 (I333981,I2514);
DFFARX1 I_19497 (I203803,I2507,I333981,I334007,);
not I_19498 (I334015,I334007);
DFFARX1 I_19499 (I203818,I2507,I333981,I334041,);
not I_19500 (I334049,I203821);
nand I_19501 (I334066,I334049,I203800);
not I_19502 (I334083,I334066);
nor I_19503 (I334100,I334083,I203824);
nor I_19504 (I334117,I334015,I334100);
DFFARX1 I_19505 (I334117,I2507,I333981,I333967,);
not I_19506 (I334148,I203824);
nand I_19507 (I334165,I334148,I334083);
and I_19508 (I334182,I334148,I203806);
nand I_19509 (I334199,I334182,I203797);
nor I_19510 (I333964,I334199,I334148);
and I_19511 (I333955,I334041,I334199);
not I_19512 (I334244,I334199);
nand I_19513 (I333958,I334041,I334244);
nor I_19514 (I333952,I334007,I334199);
not I_19515 (I334289,I203797);
nor I_19516 (I334306,I334289,I203806);
nand I_19517 (I334323,I334306,I334148);
nor I_19518 (I333961,I334066,I334323);
nor I_19519 (I334354,I334289,I203812);
and I_19520 (I334371,I334354,I203815);
or I_19521 (I334388,I334371,I203809);
DFFARX1 I_19522 (I334388,I2507,I333981,I334414,);
nor I_19523 (I334422,I334414,I334165);
DFFARX1 I_19524 (I334422,I2507,I333981,I333949,);
DFFARX1 I_19525 (I334414,I2507,I333981,I333973,);
not I_19526 (I334467,I334414);
nor I_19527 (I334484,I334467,I334041);
nor I_19528 (I334501,I334306,I334484);
DFFARX1 I_19529 (I334501,I2507,I333981,I333970,);
not I_19530 (I334559,I2514);
DFFARX1 I_19531 (I79959,I2507,I334559,I334585,);
not I_19532 (I334593,I334585);
DFFARX1 I_19533 (I79938,I2507,I334559,I334619,);
not I_19534 (I334627,I79935);
nand I_19535 (I334644,I334627,I79950);
not I_19536 (I334661,I334644);
nor I_19537 (I334678,I334661,I79938);
nor I_19538 (I334695,I334593,I334678);
DFFARX1 I_19539 (I334695,I2507,I334559,I334545,);
not I_19540 (I334726,I79938);
nand I_19541 (I334743,I334726,I334661);
and I_19542 (I334760,I334726,I79941);
nand I_19543 (I334777,I334760,I79956);
nor I_19544 (I334542,I334777,I334726);
and I_19545 (I334533,I334619,I334777);
not I_19546 (I334822,I334777);
nand I_19547 (I334536,I334619,I334822);
nor I_19548 (I334530,I334585,I334777);
not I_19549 (I334867,I79947);
nor I_19550 (I334884,I334867,I79941);
nand I_19551 (I334901,I334884,I334726);
nor I_19552 (I334539,I334644,I334901);
nor I_19553 (I334932,I334867,I79935);
and I_19554 (I334949,I334932,I79944);
or I_19555 (I334966,I334949,I79953);
DFFARX1 I_19556 (I334966,I2507,I334559,I334992,);
nor I_19557 (I335000,I334992,I334743);
DFFARX1 I_19558 (I335000,I2507,I334559,I334527,);
DFFARX1 I_19559 (I334992,I2507,I334559,I334551,);
not I_19560 (I335045,I334992);
nor I_19561 (I335062,I335045,I334619);
nor I_19562 (I335079,I334884,I335062);
DFFARX1 I_19563 (I335079,I2507,I334559,I334548,);
not I_19564 (I335137,I2514);
DFFARX1 I_19565 (I387703,I2507,I335137,I335163,);
not I_19566 (I335171,I335163);
DFFARX1 I_19567 (I387715,I2507,I335137,I335197,);
not I_19568 (I335205,I387706);
nand I_19569 (I335222,I335205,I387709);
not I_19570 (I335239,I335222);
nor I_19571 (I335256,I335239,I387712);
nor I_19572 (I335273,I335171,I335256);
DFFARX1 I_19573 (I335273,I2507,I335137,I335123,);
not I_19574 (I335304,I387712);
nand I_19575 (I335321,I335304,I335239);
and I_19576 (I335338,I335304,I387706);
nand I_19577 (I335355,I335338,I387718);
nor I_19578 (I335120,I335355,I335304);
and I_19579 (I335111,I335197,I335355);
not I_19580 (I335400,I335355);
nand I_19581 (I335114,I335197,I335400);
nor I_19582 (I335108,I335163,I335355);
not I_19583 (I335445,I387724);
nor I_19584 (I335462,I335445,I387706);
nand I_19585 (I335479,I335462,I335304);
nor I_19586 (I335117,I335222,I335479);
nor I_19587 (I335510,I335445,I387703);
and I_19588 (I335527,I335510,I387721);
or I_19589 (I335544,I335527,I387727);
DFFARX1 I_19590 (I335544,I2507,I335137,I335570,);
nor I_19591 (I335578,I335570,I335321);
DFFARX1 I_19592 (I335578,I2507,I335137,I335105,);
DFFARX1 I_19593 (I335570,I2507,I335137,I335129,);
not I_19594 (I335623,I335570);
nor I_19595 (I335640,I335623,I335197);
nor I_19596 (I335657,I335462,I335640);
DFFARX1 I_19597 (I335657,I2507,I335137,I335126,);
not I_19598 (I335715,I2514);
DFFARX1 I_19599 (I131834,I2507,I335715,I335741,);
not I_19600 (I335749,I335741);
DFFARX1 I_19601 (I131819,I2507,I335715,I335775,);
not I_19602 (I335783,I131837);
nand I_19603 (I335800,I335783,I131822);
not I_19604 (I335817,I335800);
nor I_19605 (I335834,I335817,I131819);
nor I_19606 (I335851,I335749,I335834);
DFFARX1 I_19607 (I335851,I2507,I335715,I335701,);
not I_19608 (I335882,I131819);
nand I_19609 (I335899,I335882,I335817);
and I_19610 (I335916,I335882,I131822);
nand I_19611 (I335933,I335916,I131843);
nor I_19612 (I335698,I335933,I335882);
and I_19613 (I335689,I335775,I335933);
not I_19614 (I335978,I335933);
nand I_19615 (I335692,I335775,I335978);
nor I_19616 (I335686,I335741,I335933);
not I_19617 (I336023,I131831);
nor I_19618 (I336040,I336023,I131822);
nand I_19619 (I336057,I336040,I335882);
nor I_19620 (I335695,I335800,I336057);
nor I_19621 (I336088,I336023,I131825);
and I_19622 (I336105,I336088,I131840);
or I_19623 (I336122,I336105,I131828);
DFFARX1 I_19624 (I336122,I2507,I335715,I336148,);
nor I_19625 (I336156,I336148,I335899);
DFFARX1 I_19626 (I336156,I2507,I335715,I335683,);
DFFARX1 I_19627 (I336148,I2507,I335715,I335707,);
not I_19628 (I336201,I336148);
nor I_19629 (I336218,I336201,I335775);
nor I_19630 (I336235,I336040,I336218);
DFFARX1 I_19631 (I336235,I2507,I335715,I335704,);
not I_19632 (I336293,I2514);
DFFARX1 I_19633 (I199587,I2507,I336293,I336319,);
not I_19634 (I336327,I336319);
DFFARX1 I_19635 (I199602,I2507,I336293,I336353,);
not I_19636 (I336361,I199605);
nand I_19637 (I336378,I336361,I199584);
not I_19638 (I336395,I336378);
nor I_19639 (I336412,I336395,I199608);
nor I_19640 (I336429,I336327,I336412);
DFFARX1 I_19641 (I336429,I2507,I336293,I336279,);
not I_19642 (I336460,I199608);
nand I_19643 (I336477,I336460,I336395);
and I_19644 (I336494,I336460,I199590);
nand I_19645 (I336511,I336494,I199581);
nor I_19646 (I336276,I336511,I336460);
and I_19647 (I336267,I336353,I336511);
not I_19648 (I336556,I336511);
nand I_19649 (I336270,I336353,I336556);
nor I_19650 (I336264,I336319,I336511);
not I_19651 (I336601,I199581);
nor I_19652 (I336618,I336601,I199590);
nand I_19653 (I336635,I336618,I336460);
nor I_19654 (I336273,I336378,I336635);
nor I_19655 (I336666,I336601,I199596);
and I_19656 (I336683,I336666,I199599);
or I_19657 (I336700,I336683,I199593);
DFFARX1 I_19658 (I336700,I2507,I336293,I336726,);
nor I_19659 (I336734,I336726,I336477);
DFFARX1 I_19660 (I336734,I2507,I336293,I336261,);
DFFARX1 I_19661 (I336726,I2507,I336293,I336285,);
not I_19662 (I336779,I336726);
nor I_19663 (I336796,I336779,I336353);
nor I_19664 (I336813,I336618,I336796);
DFFARX1 I_19665 (I336813,I2507,I336293,I336282,);
not I_19666 (I336871,I2514);
DFFARX1 I_19667 (I425851,I2507,I336871,I336897,);
not I_19668 (I336905,I336897);
DFFARX1 I_19669 (I425863,I2507,I336871,I336931,);
not I_19670 (I336939,I425854);
nand I_19671 (I336956,I336939,I425857);
not I_19672 (I336973,I336956);
nor I_19673 (I336990,I336973,I425860);
nor I_19674 (I337007,I336905,I336990);
DFFARX1 I_19675 (I337007,I2507,I336871,I336857,);
not I_19676 (I337038,I425860);
nand I_19677 (I337055,I337038,I336973);
and I_19678 (I337072,I337038,I425854);
nand I_19679 (I337089,I337072,I425866);
nor I_19680 (I336854,I337089,I337038);
and I_19681 (I336845,I336931,I337089);
not I_19682 (I337134,I337089);
nand I_19683 (I336848,I336931,I337134);
nor I_19684 (I336842,I336897,I337089);
not I_19685 (I337179,I425872);
nor I_19686 (I337196,I337179,I425854);
nand I_19687 (I337213,I337196,I337038);
nor I_19688 (I336851,I336956,I337213);
nor I_19689 (I337244,I337179,I425851);
and I_19690 (I337261,I337244,I425869);
or I_19691 (I337278,I337261,I425875);
DFFARX1 I_19692 (I337278,I2507,I336871,I337304,);
nor I_19693 (I337312,I337304,I337055);
DFFARX1 I_19694 (I337312,I2507,I336871,I336839,);
DFFARX1 I_19695 (I337304,I2507,I336871,I336863,);
not I_19696 (I337357,I337304);
nor I_19697 (I337374,I337357,I336931);
nor I_19698 (I337391,I337196,I337374);
DFFARX1 I_19699 (I337391,I2507,I336871,I336860,);
not I_19700 (I337449,I2514);
DFFARX1 I_19701 (I130644,I2507,I337449,I337475,);
not I_19702 (I337483,I337475);
DFFARX1 I_19703 (I130629,I2507,I337449,I337509,);
not I_19704 (I337517,I130647);
nand I_19705 (I337534,I337517,I130632);
not I_19706 (I337551,I337534);
nor I_19707 (I337568,I337551,I130629);
nor I_19708 (I337585,I337483,I337568);
DFFARX1 I_19709 (I337585,I2507,I337449,I337435,);
not I_19710 (I337616,I130629);
nand I_19711 (I337633,I337616,I337551);
and I_19712 (I337650,I337616,I130632);
nand I_19713 (I337667,I337650,I130653);
nor I_19714 (I337432,I337667,I337616);
and I_19715 (I337423,I337509,I337667);
not I_19716 (I337712,I337667);
nand I_19717 (I337426,I337509,I337712);
nor I_19718 (I337420,I337475,I337667);
not I_19719 (I337757,I130641);
nor I_19720 (I337774,I337757,I130632);
nand I_19721 (I337791,I337774,I337616);
nor I_19722 (I337429,I337534,I337791);
nor I_19723 (I337822,I337757,I130635);
and I_19724 (I337839,I337822,I130650);
or I_19725 (I337856,I337839,I130638);
DFFARX1 I_19726 (I337856,I2507,I337449,I337882,);
nor I_19727 (I337890,I337882,I337633);
DFFARX1 I_19728 (I337890,I2507,I337449,I337417,);
DFFARX1 I_19729 (I337882,I2507,I337449,I337441,);
not I_19730 (I337935,I337882);
nor I_19731 (I337952,I337935,I337509);
nor I_19732 (I337969,I337774,I337952);
DFFARX1 I_19733 (I337969,I2507,I337449,I337438,);
not I_19734 (I338027,I2514);
DFFARX1 I_19735 (I234596,I2507,I338027,I338053,);
not I_19736 (I338061,I338053);
DFFARX1 I_19737 (I234608,I2507,I338027,I338087,);
not I_19738 (I338095,I234584);
nand I_19739 (I338112,I338095,I234611);
not I_19740 (I338129,I338112);
nor I_19741 (I338146,I338129,I234599);
nor I_19742 (I338163,I338061,I338146);
DFFARX1 I_19743 (I338163,I2507,I338027,I338013,);
not I_19744 (I338194,I234599);
nand I_19745 (I338211,I338194,I338129);
and I_19746 (I338228,I338194,I234584);
nand I_19747 (I338245,I338228,I234587);
nor I_19748 (I338010,I338245,I338194);
and I_19749 (I338001,I338087,I338245);
not I_19750 (I338290,I338245);
nand I_19751 (I338004,I338087,I338290);
nor I_19752 (I337998,I338053,I338245);
not I_19753 (I338335,I234593);
nor I_19754 (I338352,I338335,I234584);
nand I_19755 (I338369,I338352,I338194);
nor I_19756 (I338007,I338112,I338369);
nor I_19757 (I338400,I338335,I234602);
and I_19758 (I338417,I338400,I234590);
or I_19759 (I338434,I338417,I234605);
DFFARX1 I_19760 (I338434,I2507,I338027,I338460,);
nor I_19761 (I338468,I338460,I338211);
DFFARX1 I_19762 (I338468,I2507,I338027,I337995,);
DFFARX1 I_19763 (I338460,I2507,I338027,I338019,);
not I_19764 (I338513,I338460);
nor I_19765 (I338530,I338513,I338087);
nor I_19766 (I338547,I338352,I338530);
DFFARX1 I_19767 (I338547,I2507,I338027,I338016,);
not I_19768 (I338605,I2514);
DFFARX1 I_19769 (I49393,I2507,I338605,I338631,);
not I_19770 (I338639,I338631);
DFFARX1 I_19771 (I49372,I2507,I338605,I338665,);
not I_19772 (I338673,I49369);
nand I_19773 (I338690,I338673,I49384);
not I_19774 (I338707,I338690);
nor I_19775 (I338724,I338707,I49372);
nor I_19776 (I338741,I338639,I338724);
DFFARX1 I_19777 (I338741,I2507,I338605,I338591,);
not I_19778 (I338772,I49372);
nand I_19779 (I338789,I338772,I338707);
and I_19780 (I338806,I338772,I49375);
nand I_19781 (I338823,I338806,I49390);
nor I_19782 (I338588,I338823,I338772);
and I_19783 (I338579,I338665,I338823);
not I_19784 (I338868,I338823);
nand I_19785 (I338582,I338665,I338868);
nor I_19786 (I338576,I338631,I338823);
not I_19787 (I338913,I49381);
nor I_19788 (I338930,I338913,I49375);
nand I_19789 (I338947,I338930,I338772);
nor I_19790 (I338585,I338690,I338947);
nor I_19791 (I338978,I338913,I49369);
and I_19792 (I338995,I338978,I49378);
or I_19793 (I339012,I338995,I49387);
DFFARX1 I_19794 (I339012,I2507,I338605,I339038,);
nor I_19795 (I339046,I339038,I338789);
DFFARX1 I_19796 (I339046,I2507,I338605,I338573,);
DFFARX1 I_19797 (I339038,I2507,I338605,I338597,);
not I_19798 (I339091,I339038);
nor I_19799 (I339108,I339091,I338665);
nor I_19800 (I339125,I338930,I339108);
DFFARX1 I_19801 (I339125,I2507,I338605,I338594,);
not I_19802 (I339183,I2514);
DFFARX1 I_19803 (I466589,I2507,I339183,I339209,);
not I_19804 (I339217,I339209);
DFFARX1 I_19805 (I466589,I2507,I339183,I339243,);
not I_19806 (I339251,I466586);
nand I_19807 (I339268,I339251,I466601);
not I_19808 (I339285,I339268);
nor I_19809 (I339302,I339285,I466595);
nor I_19810 (I339319,I339217,I339302);
DFFARX1 I_19811 (I339319,I2507,I339183,I339169,);
not I_19812 (I339350,I466595);
nand I_19813 (I339367,I339350,I339285);
and I_19814 (I339384,I339350,I466592);
nand I_19815 (I339401,I339384,I466583);
nor I_19816 (I339166,I339401,I339350);
and I_19817 (I339157,I339243,I339401);
not I_19818 (I339446,I339401);
nand I_19819 (I339160,I339243,I339446);
nor I_19820 (I339154,I339209,I339401);
not I_19821 (I339491,I466604);
nor I_19822 (I339508,I339491,I466592);
nand I_19823 (I339525,I339508,I339350);
nor I_19824 (I339163,I339268,I339525);
nor I_19825 (I339556,I339491,I466583);
and I_19826 (I339573,I339556,I466586);
or I_19827 (I339590,I339573,I466598);
DFFARX1 I_19828 (I339590,I2507,I339183,I339616,);
nor I_19829 (I339624,I339616,I339367);
DFFARX1 I_19830 (I339624,I2507,I339183,I339151,);
DFFARX1 I_19831 (I339616,I2507,I339183,I339175,);
not I_19832 (I339669,I339616);
nor I_19833 (I339686,I339669,I339243);
nor I_19834 (I339703,I339508,I339686);
DFFARX1 I_19835 (I339703,I2507,I339183,I339172,);
not I_19836 (I339761,I2514);
DFFARX1 I_19837 (I537734,I2507,I339761,I339787,);
not I_19838 (I339795,I339787);
DFFARX1 I_19839 (I537731,I2507,I339761,I339821,);
not I_19840 (I339829,I537728);
nand I_19841 (I339846,I339829,I537755);
not I_19842 (I339863,I339846);
nor I_19843 (I339880,I339863,I537743);
nor I_19844 (I339897,I339795,I339880);
DFFARX1 I_19845 (I339897,I2507,I339761,I339747,);
not I_19846 (I339928,I537743);
nand I_19847 (I339945,I339928,I339863);
and I_19848 (I339962,I339928,I537749);
nand I_19849 (I339979,I339962,I537740);
nor I_19850 (I339744,I339979,I339928);
and I_19851 (I339735,I339821,I339979);
not I_19852 (I340024,I339979);
nand I_19853 (I339738,I339821,I340024);
nor I_19854 (I339732,I339787,I339979);
not I_19855 (I340069,I537737);
nor I_19856 (I340086,I340069,I537749);
nand I_19857 (I340103,I340086,I339928);
nor I_19858 (I339741,I339846,I340103);
nor I_19859 (I340134,I340069,I537752);
and I_19860 (I340151,I340134,I537746);
or I_19861 (I340168,I340151,I537728);
DFFARX1 I_19862 (I340168,I2507,I339761,I340194,);
nor I_19863 (I340202,I340194,I339945);
DFFARX1 I_19864 (I340202,I2507,I339761,I339729,);
DFFARX1 I_19865 (I340194,I2507,I339761,I339753,);
not I_19866 (I340247,I340194);
nor I_19867 (I340264,I340247,I339821);
nor I_19868 (I340281,I340086,I340264);
DFFARX1 I_19869 (I340281,I2507,I339761,I339750,);
not I_19870 (I340339,I2514);
DFFARX1 I_19871 (I707303,I2507,I340339,I340365,);
not I_19872 (I340373,I340365);
DFFARX1 I_19873 (I707303,I2507,I340339,I340399,);
not I_19874 (I340407,I707327);
nand I_19875 (I340424,I340407,I707309);
not I_19876 (I340441,I340424);
nor I_19877 (I340458,I340441,I707324);
nor I_19878 (I340475,I340373,I340458);
DFFARX1 I_19879 (I340475,I2507,I340339,I340325,);
not I_19880 (I340506,I707324);
nand I_19881 (I340523,I340506,I340441);
and I_19882 (I340540,I340506,I707306);
nand I_19883 (I340557,I340540,I707315);
nor I_19884 (I340322,I340557,I340506);
and I_19885 (I340313,I340399,I340557);
not I_19886 (I340602,I340557);
nand I_19887 (I340316,I340399,I340602);
nor I_19888 (I340310,I340365,I340557);
not I_19889 (I340647,I707312);
nor I_19890 (I340664,I340647,I707306);
nand I_19891 (I340681,I340664,I340506);
nor I_19892 (I340319,I340424,I340681);
nor I_19893 (I340712,I340647,I707321);
and I_19894 (I340729,I340712,I707330);
or I_19895 (I340746,I340729,I707318);
DFFARX1 I_19896 (I340746,I2507,I340339,I340772,);
nor I_19897 (I340780,I340772,I340523);
DFFARX1 I_19898 (I340780,I2507,I340339,I340307,);
DFFARX1 I_19899 (I340772,I2507,I340339,I340331,);
not I_19900 (I340825,I340772);
nor I_19901 (I340842,I340825,I340399);
nor I_19902 (I340859,I340664,I340842);
DFFARX1 I_19903 (I340859,I2507,I340339,I340328,);
not I_19904 (I340917,I2514);
DFFARX1 I_19905 (I484116,I2507,I340917,I340943,);
not I_19906 (I340951,I340943);
DFFARX1 I_19907 (I484113,I2507,I340917,I340977,);
not I_19908 (I340985,I484110);
nand I_19909 (I341002,I340985,I484137);
not I_19910 (I341019,I341002);
nor I_19911 (I341036,I341019,I484125);
nor I_19912 (I341053,I340951,I341036);
DFFARX1 I_19913 (I341053,I2507,I340917,I340903,);
not I_19914 (I341084,I484125);
nand I_19915 (I341101,I341084,I341019);
and I_19916 (I341118,I341084,I484131);
nand I_19917 (I341135,I341118,I484122);
nor I_19918 (I340900,I341135,I341084);
and I_19919 (I340891,I340977,I341135);
not I_19920 (I341180,I341135);
nand I_19921 (I340894,I340977,I341180);
nor I_19922 (I340888,I340943,I341135);
not I_19923 (I341225,I484119);
nor I_19924 (I341242,I341225,I484131);
nand I_19925 (I341259,I341242,I341084);
nor I_19926 (I340897,I341002,I341259);
nor I_19927 (I341290,I341225,I484134);
and I_19928 (I341307,I341290,I484128);
or I_19929 (I341324,I341307,I484110);
DFFARX1 I_19930 (I341324,I2507,I340917,I341350,);
nor I_19931 (I341358,I341350,I341101);
DFFARX1 I_19932 (I341358,I2507,I340917,I340885,);
DFFARX1 I_19933 (I341350,I2507,I340917,I340909,);
not I_19934 (I341403,I341350);
nor I_19935 (I341420,I341403,I340977);
nor I_19936 (I341437,I341242,I341420);
DFFARX1 I_19937 (I341437,I2507,I340917,I340906,);
not I_19938 (I341495,I2514);
DFFARX1 I_19939 (I3719,I2507,I341495,I341521,);
not I_19940 (I341529,I341521);
DFFARX1 I_19941 (I3707,I2507,I341495,I341555,);
not I_19942 (I341563,I3716);
nand I_19943 (I341580,I341563,I3713);
not I_19944 (I341597,I341580);
nor I_19945 (I341614,I341597,I3722);
nor I_19946 (I341631,I341529,I341614);
DFFARX1 I_19947 (I341631,I2507,I341495,I341481,);
not I_19948 (I341662,I3722);
nand I_19949 (I341679,I341662,I341597);
and I_19950 (I341696,I341662,I3710);
nand I_19951 (I341713,I341696,I3713);
nor I_19952 (I341478,I341713,I341662);
and I_19953 (I341469,I341555,I341713);
not I_19954 (I341758,I341713);
nand I_19955 (I341472,I341555,I341758);
nor I_19956 (I341466,I341521,I341713);
not I_19957 (I341803,I3728);
nor I_19958 (I341820,I341803,I3710);
nand I_19959 (I341837,I341820,I341662);
nor I_19960 (I341475,I341580,I341837);
nor I_19961 (I341868,I341803,I3710);
and I_19962 (I341885,I341868,I3725);
or I_19963 (I341902,I341885,I3707);
DFFARX1 I_19964 (I341902,I2507,I341495,I341928,);
nor I_19965 (I341936,I341928,I341679);
DFFARX1 I_19966 (I341936,I2507,I341495,I341463,);
DFFARX1 I_19967 (I341928,I2507,I341495,I341487,);
not I_19968 (I341981,I341928);
nor I_19969 (I341998,I341981,I341555);
nor I_19970 (I342015,I341820,I341998);
DFFARX1 I_19971 (I342015,I2507,I341495,I341484,);
not I_19972 (I342073,I2514);
DFFARX1 I_19973 (I472386,I2507,I342073,I342099,);
not I_19974 (I342107,I342099);
DFFARX1 I_19975 (I472386,I2507,I342073,I342133,);
not I_19976 (I342141,I472383);
nand I_19977 (I342158,I342141,I472398);
not I_19978 (I342175,I342158);
nor I_19979 (I342192,I342175,I472392);
nor I_19980 (I342209,I342107,I342192);
DFFARX1 I_19981 (I342209,I2507,I342073,I342059,);
not I_19982 (I342240,I472392);
nand I_19983 (I342257,I342240,I342175);
and I_19984 (I342274,I342240,I472389);
nand I_19985 (I342291,I342274,I472380);
nor I_19986 (I342056,I342291,I342240);
and I_19987 (I342047,I342133,I342291);
not I_19988 (I342336,I342291);
nand I_19989 (I342050,I342133,I342336);
nor I_19990 (I342044,I342099,I342291);
not I_19991 (I342381,I472401);
nor I_19992 (I342398,I342381,I472389);
nand I_19993 (I342415,I342398,I342240);
nor I_19994 (I342053,I342158,I342415);
nor I_19995 (I342446,I342381,I472380);
and I_19996 (I342463,I342446,I472383);
or I_19997 (I342480,I342463,I472395);
DFFARX1 I_19998 (I342480,I2507,I342073,I342506,);
nor I_19999 (I342514,I342506,I342257);
DFFARX1 I_20000 (I342514,I2507,I342073,I342041,);
DFFARX1 I_20001 (I342506,I2507,I342073,I342065,);
not I_20002 (I342559,I342506);
nor I_20003 (I342576,I342559,I342133);
nor I_20004 (I342593,I342398,I342576);
DFFARX1 I_20005 (I342593,I2507,I342073,I342062,);
not I_20006 (I342651,I2514);
DFFARX1 I_20007 (I95539,I2507,I342651,I342677,);
not I_20008 (I342685,I342677);
DFFARX1 I_20009 (I95524,I2507,I342651,I342711,);
not I_20010 (I342719,I95542);
nand I_20011 (I342736,I342719,I95527);
not I_20012 (I342753,I342736);
nor I_20013 (I342770,I342753,I95524);
nor I_20014 (I342787,I342685,I342770);
DFFARX1 I_20015 (I342787,I2507,I342651,I342637,);
not I_20016 (I342818,I95524);
nand I_20017 (I342835,I342818,I342753);
and I_20018 (I342852,I342818,I95527);
nand I_20019 (I342869,I342852,I95548);
nor I_20020 (I342634,I342869,I342818);
and I_20021 (I342625,I342711,I342869);
not I_20022 (I342914,I342869);
nand I_20023 (I342628,I342711,I342914);
nor I_20024 (I342622,I342677,I342869);
not I_20025 (I342959,I95536);
nor I_20026 (I342976,I342959,I95527);
nand I_20027 (I342993,I342976,I342818);
nor I_20028 (I342631,I342736,I342993);
nor I_20029 (I343024,I342959,I95530);
and I_20030 (I343041,I343024,I95545);
or I_20031 (I343058,I343041,I95533);
DFFARX1 I_20032 (I343058,I2507,I342651,I343084,);
nor I_20033 (I343092,I343084,I342835);
DFFARX1 I_20034 (I343092,I2507,I342651,I342619,);
DFFARX1 I_20035 (I343084,I2507,I342651,I342643,);
not I_20036 (I343137,I343084);
nor I_20037 (I343154,I343137,I342711);
nor I_20038 (I343171,I342976,I343154);
DFFARX1 I_20039 (I343171,I2507,I342651,I342640,);
not I_20040 (I343229,I2514);
DFFARX1 I_20041 (I275940,I2507,I343229,I343255,);
not I_20042 (I343263,I343255);
DFFARX1 I_20043 (I275952,I2507,I343229,I343289,);
not I_20044 (I343297,I275928);
nand I_20045 (I343314,I343297,I275955);
not I_20046 (I343331,I343314);
nor I_20047 (I343348,I343331,I275943);
nor I_20048 (I343365,I343263,I343348);
DFFARX1 I_20049 (I343365,I2507,I343229,I343215,);
not I_20050 (I343396,I275943);
nand I_20051 (I343413,I343396,I343331);
and I_20052 (I343430,I343396,I275928);
nand I_20053 (I343447,I343430,I275931);
nor I_20054 (I343212,I343447,I343396);
and I_20055 (I343203,I343289,I343447);
not I_20056 (I343492,I343447);
nand I_20057 (I343206,I343289,I343492);
nor I_20058 (I343200,I343255,I343447);
not I_20059 (I343537,I275937);
nor I_20060 (I343554,I343537,I275928);
nand I_20061 (I343571,I343554,I343396);
nor I_20062 (I343209,I343314,I343571);
nor I_20063 (I343602,I343537,I275946);
and I_20064 (I343619,I343602,I275934);
or I_20065 (I343636,I343619,I275949);
DFFARX1 I_20066 (I343636,I2507,I343229,I343662,);
nor I_20067 (I343670,I343662,I343413);
DFFARX1 I_20068 (I343670,I2507,I343229,I343197,);
DFFARX1 I_20069 (I343662,I2507,I343229,I343221,);
not I_20070 (I343715,I343662);
nor I_20071 (I343732,I343715,I343289);
nor I_20072 (I343749,I343554,I343732);
DFFARX1 I_20073 (I343749,I2507,I343229,I343218,);
not I_20074 (I343807,I2514);
DFFARX1 I_20075 (I299816,I2507,I343807,I343833,);
not I_20076 (I343841,I343833);
DFFARX1 I_20077 (I299828,I2507,I343807,I343867,);
not I_20078 (I343875,I299834);
nand I_20079 (I343892,I343875,I299825);
not I_20080 (I343909,I343892);
nor I_20081 (I343926,I343909,I299831);
nor I_20082 (I343943,I343841,I343926);
DFFARX1 I_20083 (I343943,I2507,I343807,I343793,);
not I_20084 (I343974,I299831);
nand I_20085 (I343991,I343974,I343909);
and I_20086 (I344008,I343974,I299822);
nand I_20087 (I344025,I344008,I299813);
nor I_20088 (I343790,I344025,I343974);
and I_20089 (I343781,I343867,I344025);
not I_20090 (I344070,I344025);
nand I_20091 (I343784,I343867,I344070);
nor I_20092 (I343778,I343833,I344025);
not I_20093 (I344115,I299819);
nor I_20094 (I344132,I344115,I299822);
nand I_20095 (I344149,I344132,I343974);
nor I_20096 (I343787,I343892,I344149);
nor I_20097 (I344180,I344115,I299816);
and I_20098 (I344197,I344180,I299813);
or I_20099 (I344214,I344197,I299837);
DFFARX1 I_20100 (I344214,I2507,I343807,I344240,);
nor I_20101 (I344248,I344240,I343991);
DFFARX1 I_20102 (I344248,I2507,I343807,I343775,);
DFFARX1 I_20103 (I344240,I2507,I343807,I343799,);
not I_20104 (I344293,I344240);
nor I_20105 (I344310,I344293,I343867);
nor I_20106 (I344327,I344132,I344310);
DFFARX1 I_20107 (I344327,I2507,I343807,I343796,);
not I_20108 (I344385,I2514);
DFFARX1 I_20109 (I560444,I2507,I344385,I344411,);
not I_20110 (I344419,I344411);
DFFARX1 I_20111 (I560435,I2507,I344385,I344445,);
not I_20112 (I344453,I560429);
nand I_20113 (I344470,I344453,I560441);
not I_20114 (I344487,I344470);
nor I_20115 (I344504,I344487,I560432);
nor I_20116 (I344521,I344419,I344504);
DFFARX1 I_20117 (I344521,I2507,I344385,I344371,);
not I_20118 (I344552,I560432);
nand I_20119 (I344569,I344552,I344487);
and I_20120 (I344586,I344552,I560438);
nand I_20121 (I344603,I344586,I560423);
nor I_20122 (I344368,I344603,I344552);
and I_20123 (I344359,I344445,I344603);
not I_20124 (I344648,I344603);
nand I_20125 (I344362,I344445,I344648);
nor I_20126 (I344356,I344411,I344603);
not I_20127 (I344693,I560423);
nor I_20128 (I344710,I344693,I560438);
nand I_20129 (I344727,I344710,I344552);
nor I_20130 (I344365,I344470,I344727);
nor I_20131 (I344758,I344693,I560426);
and I_20132 (I344775,I344758,I560429);
or I_20133 (I344792,I344775,I560426);
DFFARX1 I_20134 (I344792,I2507,I344385,I344818,);
nor I_20135 (I344826,I344818,I344569);
DFFARX1 I_20136 (I344826,I2507,I344385,I344353,);
DFFARX1 I_20137 (I344818,I2507,I344385,I344377,);
not I_20138 (I344871,I344818);
nor I_20139 (I344888,I344871,I344445);
nor I_20140 (I344905,I344710,I344888);
DFFARX1 I_20141 (I344905,I2507,I344385,I344374,);
not I_20142 (I344963,I2514);
DFFARX1 I_20143 (I369785,I2507,I344963,I344989,);
not I_20144 (I344997,I344989);
DFFARX1 I_20145 (I369797,I2507,I344963,I345023,);
not I_20146 (I345031,I369788);
nand I_20147 (I345048,I345031,I369791);
not I_20148 (I345065,I345048);
nor I_20149 (I345082,I345065,I369794);
nor I_20150 (I345099,I344997,I345082);
DFFARX1 I_20151 (I345099,I2507,I344963,I344949,);
not I_20152 (I345130,I369794);
nand I_20153 (I345147,I345130,I345065);
and I_20154 (I345164,I345130,I369788);
nand I_20155 (I345181,I345164,I369800);
nor I_20156 (I344946,I345181,I345130);
and I_20157 (I344937,I345023,I345181);
not I_20158 (I345226,I345181);
nand I_20159 (I344940,I345023,I345226);
nor I_20160 (I344934,I344989,I345181);
not I_20161 (I345271,I369806);
nor I_20162 (I345288,I345271,I369788);
nand I_20163 (I345305,I345288,I345130);
nor I_20164 (I344943,I345048,I345305);
nor I_20165 (I345336,I345271,I369785);
and I_20166 (I345353,I345336,I369803);
or I_20167 (I345370,I345353,I369809);
DFFARX1 I_20168 (I345370,I2507,I344963,I345396,);
nor I_20169 (I345404,I345396,I345147);
DFFARX1 I_20170 (I345404,I2507,I344963,I344931,);
DFFARX1 I_20171 (I345396,I2507,I344963,I344955,);
not I_20172 (I345449,I345396);
nor I_20173 (I345466,I345449,I345023);
nor I_20174 (I345483,I345288,I345466);
DFFARX1 I_20175 (I345483,I2507,I344963,I344952,);
not I_20176 (I345541,I2514);
DFFARX1 I_20177 (I469224,I2507,I345541,I345567,);
not I_20178 (I345575,I345567);
DFFARX1 I_20179 (I469224,I2507,I345541,I345601,);
not I_20180 (I345609,I469221);
nand I_20181 (I345626,I345609,I469236);
not I_20182 (I345643,I345626);
nor I_20183 (I345660,I345643,I469230);
nor I_20184 (I345677,I345575,I345660);
DFFARX1 I_20185 (I345677,I2507,I345541,I345527,);
not I_20186 (I345708,I469230);
nand I_20187 (I345725,I345708,I345643);
and I_20188 (I345742,I345708,I469227);
nand I_20189 (I345759,I345742,I469218);
nor I_20190 (I345524,I345759,I345708);
and I_20191 (I345515,I345601,I345759);
not I_20192 (I345804,I345759);
nand I_20193 (I345518,I345601,I345804);
nor I_20194 (I345512,I345567,I345759);
not I_20195 (I345849,I469239);
nor I_20196 (I345866,I345849,I469227);
nand I_20197 (I345883,I345866,I345708);
nor I_20198 (I345521,I345626,I345883);
nor I_20199 (I345914,I345849,I469218);
and I_20200 (I345931,I345914,I469221);
or I_20201 (I345948,I345931,I469233);
DFFARX1 I_20202 (I345948,I2507,I345541,I345974,);
nor I_20203 (I345982,I345974,I345725);
DFFARX1 I_20204 (I345982,I2507,I345541,I345509,);
DFFARX1 I_20205 (I345974,I2507,I345541,I345533,);
not I_20206 (I346027,I345974);
nor I_20207 (I346044,I346027,I345601);
nor I_20208 (I346061,I345866,I346044);
DFFARX1 I_20209 (I346061,I2507,I345541,I345530,);
not I_20210 (I346119,I2514);
DFFARX1 I_20211 (I671717,I2507,I346119,I346145,);
not I_20212 (I346153,I346145);
DFFARX1 I_20213 (I671729,I2507,I346119,I346179,);
not I_20214 (I346187,I671720);
nand I_20215 (I346204,I346187,I671708);
not I_20216 (I346221,I346204);
nor I_20217 (I346238,I346221,I671705);
nor I_20218 (I346255,I346153,I346238);
DFFARX1 I_20219 (I346255,I2507,I346119,I346105,);
not I_20220 (I346286,I671705);
nand I_20221 (I346303,I346286,I346221);
and I_20222 (I346320,I346286,I671711);
nand I_20223 (I346337,I346320,I671708);
nor I_20224 (I346102,I346337,I346286);
and I_20225 (I346093,I346179,I346337);
not I_20226 (I346382,I346337);
nand I_20227 (I346096,I346179,I346382);
nor I_20228 (I346090,I346145,I346337);
not I_20229 (I346427,I671726);
nor I_20230 (I346444,I346427,I671711);
nand I_20231 (I346461,I346444,I346286);
nor I_20232 (I346099,I346204,I346461);
nor I_20233 (I346492,I346427,I671714);
and I_20234 (I346509,I346492,I671705);
or I_20235 (I346526,I346509,I671723);
DFFARX1 I_20236 (I346526,I2507,I346119,I346552,);
nor I_20237 (I346560,I346552,I346303);
DFFARX1 I_20238 (I346560,I2507,I346119,I346087,);
DFFARX1 I_20239 (I346552,I2507,I346119,I346111,);
not I_20240 (I346605,I346552);
nor I_20241 (I346622,I346605,I346179);
nor I_20242 (I346639,I346444,I346622);
DFFARX1 I_20243 (I346639,I2507,I346119,I346108,);
not I_20244 (I346697,I2514);
DFFARX1 I_20245 (I278657,I2507,I346697,I346723,);
not I_20246 (I346731,I346723);
nand I_20247 (I346748,I278648,I278666);
and I_20248 (I346765,I346748,I278669);
DFFARX1 I_20249 (I346765,I2507,I346697,I346791,);
not I_20250 (I346799,I278663);
DFFARX1 I_20251 (I278651,I2507,I346697,I346825,);
not I_20252 (I346833,I346825);
nor I_20253 (I346850,I346833,I346731);
and I_20254 (I346867,I346850,I278663);
nor I_20255 (I346884,I346833,I346799);
nor I_20256 (I346680,I346791,I346884);
DFFARX1 I_20257 (I278660,I2507,I346697,I346924,);
nor I_20258 (I346932,I346924,I346791);
not I_20259 (I346949,I346932);
not I_20260 (I346966,I346924);
nor I_20261 (I346983,I346966,I346867);
DFFARX1 I_20262 (I346983,I2507,I346697,I346683,);
nand I_20263 (I347014,I278675,I278672);
and I_20264 (I347031,I347014,I278654);
DFFARX1 I_20265 (I347031,I2507,I346697,I347057,);
nor I_20266 (I347065,I347057,I346924);
DFFARX1 I_20267 (I347065,I2507,I346697,I346665,);
nand I_20268 (I347096,I347057,I346966);
nand I_20269 (I346674,I346949,I347096);
not I_20270 (I347127,I347057);
nor I_20271 (I347144,I347127,I346867);
DFFARX1 I_20272 (I347144,I2507,I346697,I346686,);
nor I_20273 (I347175,I278648,I278672);
or I_20274 (I346677,I346924,I347175);
nor I_20275 (I346668,I347057,I347175);
or I_20276 (I346671,I346791,I347175);
DFFARX1 I_20277 (I347175,I2507,I346697,I346689,);
not I_20278 (I347275,I2514);
DFFARX1 I_20279 (I541355,I2507,I347275,I347301,);
not I_20280 (I347309,I347301);
nand I_20281 (I347326,I541352,I541370);
and I_20282 (I347343,I347326,I541367);
DFFARX1 I_20283 (I347343,I2507,I347275,I347369,);
not I_20284 (I347377,I541349);
DFFARX1 I_20285 (I541352,I2507,I347275,I347403,);
not I_20286 (I347411,I347403);
nor I_20287 (I347428,I347411,I347309);
and I_20288 (I347445,I347428,I541349);
nor I_20289 (I347462,I347411,I347377);
nor I_20290 (I347258,I347369,I347462);
DFFARX1 I_20291 (I541361,I2507,I347275,I347502,);
nor I_20292 (I347510,I347502,I347369);
not I_20293 (I347527,I347510);
not I_20294 (I347544,I347502);
nor I_20295 (I347561,I347544,I347445);
DFFARX1 I_20296 (I347561,I2507,I347275,I347261,);
nand I_20297 (I347592,I541364,I541349);
and I_20298 (I347609,I347592,I541355);
DFFARX1 I_20299 (I347609,I2507,I347275,I347635,);
nor I_20300 (I347643,I347635,I347502);
DFFARX1 I_20301 (I347643,I2507,I347275,I347243,);
nand I_20302 (I347674,I347635,I347544);
nand I_20303 (I347252,I347527,I347674);
not I_20304 (I347705,I347635);
nor I_20305 (I347722,I347705,I347445);
DFFARX1 I_20306 (I347722,I2507,I347275,I347264,);
nor I_20307 (I347753,I541358,I541349);
or I_20308 (I347255,I347502,I347753);
nor I_20309 (I347246,I347635,I347753);
or I_20310 (I347249,I347369,I347753);
DFFARX1 I_20311 (I347753,I2507,I347275,I347267,);
not I_20312 (I347853,I2514);
DFFARX1 I_20313 (I13545,I2507,I347853,I347879,);
not I_20314 (I347887,I347879);
nand I_20315 (I347904,I13542,I13533);
and I_20316 (I347921,I347904,I13533);
DFFARX1 I_20317 (I347921,I2507,I347853,I347947,);
not I_20318 (I347955,I13536);
DFFARX1 I_20319 (I13551,I2507,I347853,I347981,);
not I_20320 (I347989,I347981);
nor I_20321 (I348006,I347989,I347887);
and I_20322 (I348023,I348006,I13536);
nor I_20323 (I348040,I347989,I347955);
nor I_20324 (I347836,I347947,I348040);
DFFARX1 I_20325 (I13536,I2507,I347853,I348080,);
nor I_20326 (I348088,I348080,I347947);
not I_20327 (I348105,I348088);
not I_20328 (I348122,I348080);
nor I_20329 (I348139,I348122,I348023);
DFFARX1 I_20330 (I348139,I2507,I347853,I347839,);
nand I_20331 (I348170,I13554,I13539);
and I_20332 (I348187,I348170,I13557);
DFFARX1 I_20333 (I348187,I2507,I347853,I348213,);
nor I_20334 (I348221,I348213,I348080);
DFFARX1 I_20335 (I348221,I2507,I347853,I347821,);
nand I_20336 (I348252,I348213,I348122);
nand I_20337 (I347830,I348105,I348252);
not I_20338 (I348283,I348213);
nor I_20339 (I348300,I348283,I348023);
DFFARX1 I_20340 (I348300,I2507,I347853,I347842,);
nor I_20341 (I348331,I13548,I13539);
or I_20342 (I347833,I348080,I348331);
nor I_20343 (I347824,I348213,I348331);
or I_20344 (I347827,I347947,I348331);
DFFARX1 I_20345 (I348331,I2507,I347853,I347845,);
not I_20346 (I348431,I2514);
DFFARX1 I_20347 (I122299,I2507,I348431,I348457,);
not I_20348 (I348465,I348457);
nand I_20349 (I348482,I122302,I122323);
and I_20350 (I348499,I348482,I122311);
DFFARX1 I_20351 (I348499,I2507,I348431,I348525,);
not I_20352 (I348533,I122308);
DFFARX1 I_20353 (I122299,I2507,I348431,I348559,);
not I_20354 (I348567,I348559);
nor I_20355 (I348584,I348567,I348465);
and I_20356 (I348601,I348584,I122308);
nor I_20357 (I348618,I348567,I348533);
nor I_20358 (I348414,I348525,I348618);
DFFARX1 I_20359 (I122317,I2507,I348431,I348658,);
nor I_20360 (I348666,I348658,I348525);
not I_20361 (I348683,I348666);
not I_20362 (I348700,I348658);
nor I_20363 (I348717,I348700,I348601);
DFFARX1 I_20364 (I348717,I2507,I348431,I348417,);
nand I_20365 (I348748,I122302,I122305);
and I_20366 (I348765,I348748,I122314);
DFFARX1 I_20367 (I348765,I2507,I348431,I348791,);
nor I_20368 (I348799,I348791,I348658);
DFFARX1 I_20369 (I348799,I2507,I348431,I348399,);
nand I_20370 (I348830,I348791,I348700);
nand I_20371 (I348408,I348683,I348830);
not I_20372 (I348861,I348791);
nor I_20373 (I348878,I348861,I348601);
DFFARX1 I_20374 (I348878,I2507,I348431,I348420,);
nor I_20375 (I348909,I122320,I122305);
or I_20376 (I348411,I348658,I348909);
nor I_20377 (I348402,I348791,I348909);
or I_20378 (I348405,I348525,I348909);
DFFARX1 I_20379 (I348909,I2507,I348431,I348423,);
not I_20380 (I349009,I2514);
DFFARX1 I_20381 (I183795,I2507,I349009,I349035,);
not I_20382 (I349043,I349035);
nand I_20383 (I349060,I183798,I183774);
and I_20384 (I349077,I349060,I183771);
DFFARX1 I_20385 (I349077,I2507,I349009,I349103,);
not I_20386 (I349111,I183777);
DFFARX1 I_20387 (I183771,I2507,I349009,I349137,);
not I_20388 (I349145,I349137);
nor I_20389 (I349162,I349145,I349043);
and I_20390 (I349179,I349162,I183777);
nor I_20391 (I349196,I349145,I349111);
nor I_20392 (I348992,I349103,I349196);
DFFARX1 I_20393 (I183780,I2507,I349009,I349236,);
nor I_20394 (I349244,I349236,I349103);
not I_20395 (I349261,I349244);
not I_20396 (I349278,I349236);
nor I_20397 (I349295,I349278,I349179);
DFFARX1 I_20398 (I349295,I2507,I349009,I348995,);
nand I_20399 (I349326,I183783,I183792);
and I_20400 (I349343,I349326,I183789);
DFFARX1 I_20401 (I349343,I2507,I349009,I349369,);
nor I_20402 (I349377,I349369,I349236);
DFFARX1 I_20403 (I349377,I2507,I349009,I348977,);
nand I_20404 (I349408,I349369,I349278);
nand I_20405 (I348986,I349261,I349408);
not I_20406 (I349439,I349369);
nor I_20407 (I349456,I349439,I349179);
DFFARX1 I_20408 (I349456,I2507,I349009,I348998,);
nor I_20409 (I349487,I183786,I183792);
or I_20410 (I348989,I349236,I349487);
nor I_20411 (I348980,I349369,I349487);
or I_20412 (I348983,I349103,I349487);
DFFARX1 I_20413 (I349487,I2507,I349009,I349001,);
not I_20414 (I349587,I2514);
DFFARX1 I_20415 (I191173,I2507,I349587,I349613,);
not I_20416 (I349621,I349613);
nand I_20417 (I349638,I191176,I191152);
and I_20418 (I349655,I349638,I191149);
DFFARX1 I_20419 (I349655,I2507,I349587,I349681,);
not I_20420 (I349689,I191155);
DFFARX1 I_20421 (I191149,I2507,I349587,I349715,);
not I_20422 (I349723,I349715);
nor I_20423 (I349740,I349723,I349621);
and I_20424 (I349757,I349740,I191155);
nor I_20425 (I349774,I349723,I349689);
nor I_20426 (I349570,I349681,I349774);
DFFARX1 I_20427 (I191158,I2507,I349587,I349814,);
nor I_20428 (I349822,I349814,I349681);
not I_20429 (I349839,I349822);
not I_20430 (I349856,I349814);
nor I_20431 (I349873,I349856,I349757);
DFFARX1 I_20432 (I349873,I2507,I349587,I349573,);
nand I_20433 (I349904,I191161,I191170);
and I_20434 (I349921,I349904,I191167);
DFFARX1 I_20435 (I349921,I2507,I349587,I349947,);
nor I_20436 (I349955,I349947,I349814);
DFFARX1 I_20437 (I349955,I2507,I349587,I349555,);
nand I_20438 (I349986,I349947,I349856);
nand I_20439 (I349564,I349839,I349986);
not I_20440 (I350017,I349947);
nor I_20441 (I350034,I350017,I349757);
DFFARX1 I_20442 (I350034,I2507,I349587,I349576,);
nor I_20443 (I350065,I191164,I191170);
or I_20444 (I349567,I349814,I350065);
nor I_20445 (I349558,I349947,I350065);
or I_20446 (I349561,I349681,I350065);
DFFARX1 I_20447 (I350065,I2507,I349587,I349579,);
not I_20448 (I350165,I2514);
DFFARX1 I_20449 (I200659,I2507,I350165,I350191,);
not I_20450 (I350199,I350191);
nand I_20451 (I350216,I200662,I200638);
and I_20452 (I350233,I350216,I200635);
DFFARX1 I_20453 (I350233,I2507,I350165,I350259,);
not I_20454 (I350267,I200641);
DFFARX1 I_20455 (I200635,I2507,I350165,I350293,);
not I_20456 (I350301,I350293);
nor I_20457 (I350318,I350301,I350199);
and I_20458 (I350335,I350318,I200641);
nor I_20459 (I350352,I350301,I350267);
nor I_20460 (I350148,I350259,I350352);
DFFARX1 I_20461 (I200644,I2507,I350165,I350392,);
nor I_20462 (I350400,I350392,I350259);
not I_20463 (I350417,I350400);
not I_20464 (I350434,I350392);
nor I_20465 (I350451,I350434,I350335);
DFFARX1 I_20466 (I350451,I2507,I350165,I350151,);
nand I_20467 (I350482,I200647,I200656);
and I_20468 (I350499,I350482,I200653);
DFFARX1 I_20469 (I350499,I2507,I350165,I350525,);
nor I_20470 (I350533,I350525,I350392);
DFFARX1 I_20471 (I350533,I2507,I350165,I350133,);
nand I_20472 (I350564,I350525,I350434);
nand I_20473 (I350142,I350417,I350564);
not I_20474 (I350595,I350525);
nor I_20475 (I350612,I350595,I350335);
DFFARX1 I_20476 (I350612,I2507,I350165,I350154,);
nor I_20477 (I350643,I200650,I200656);
or I_20478 (I350145,I350392,I350643);
nor I_20479 (I350136,I350525,I350643);
or I_20480 (I350139,I350259,I350643);
DFFARX1 I_20481 (I350643,I2507,I350165,I350157,);
not I_20482 (I350743,I2514);
DFFARX1 I_20483 (I500284,I2507,I350743,I350769,);
not I_20484 (I350777,I350769);
nand I_20485 (I350794,I500260,I500275);
and I_20486 (I350811,I350794,I500287);
DFFARX1 I_20487 (I350811,I2507,I350743,I350837,);
not I_20488 (I350845,I500272);
DFFARX1 I_20489 (I500263,I2507,I350743,I350871,);
not I_20490 (I350879,I350871);
nor I_20491 (I350896,I350879,I350777);
and I_20492 (I350913,I350896,I500272);
nor I_20493 (I350930,I350879,I350845);
nor I_20494 (I350726,I350837,I350930);
DFFARX1 I_20495 (I500260,I2507,I350743,I350970,);
nor I_20496 (I350978,I350970,I350837);
not I_20497 (I350995,I350978);
not I_20498 (I351012,I350970);
nor I_20499 (I351029,I351012,I350913);
DFFARX1 I_20500 (I351029,I2507,I350743,I350729,);
nand I_20501 (I351060,I500278,I500269);
and I_20502 (I351077,I351060,I500281);
DFFARX1 I_20503 (I351077,I2507,I350743,I351103,);
nor I_20504 (I351111,I351103,I350970);
DFFARX1 I_20505 (I351111,I2507,I350743,I350711,);
nand I_20506 (I351142,I351103,I351012);
nand I_20507 (I350720,I350995,I351142);
not I_20508 (I351173,I351103);
nor I_20509 (I351190,I351173,I350913);
DFFARX1 I_20510 (I351190,I2507,I350743,I350732,);
nor I_20511 (I351221,I500266,I500269);
or I_20512 (I350723,I350970,I351221);
nor I_20513 (I350714,I351103,I351221);
or I_20514 (I350717,I350837,I351221);
DFFARX1 I_20515 (I351221,I2507,I350743,I350735,);
not I_20516 (I351321,I2514);
DFFARX1 I_20517 (I146694,I2507,I351321,I351347,);
not I_20518 (I351355,I351347);
nand I_20519 (I351372,I146697,I146718);
and I_20520 (I351389,I351372,I146706);
DFFARX1 I_20521 (I351389,I2507,I351321,I351415,);
not I_20522 (I351423,I146703);
DFFARX1 I_20523 (I146694,I2507,I351321,I351449,);
not I_20524 (I351457,I351449);
nor I_20525 (I351474,I351457,I351355);
and I_20526 (I351491,I351474,I146703);
nor I_20527 (I351508,I351457,I351423);
nor I_20528 (I351304,I351415,I351508);
DFFARX1 I_20529 (I146712,I2507,I351321,I351548,);
nor I_20530 (I351556,I351548,I351415);
not I_20531 (I351573,I351556);
not I_20532 (I351590,I351548);
nor I_20533 (I351607,I351590,I351491);
DFFARX1 I_20534 (I351607,I2507,I351321,I351307,);
nand I_20535 (I351638,I146697,I146700);
and I_20536 (I351655,I351638,I146709);
DFFARX1 I_20537 (I351655,I2507,I351321,I351681,);
nor I_20538 (I351689,I351681,I351548);
DFFARX1 I_20539 (I351689,I2507,I351321,I351289,);
nand I_20540 (I351720,I351681,I351590);
nand I_20541 (I351298,I351573,I351720);
not I_20542 (I351751,I351681);
nor I_20543 (I351768,I351751,I351491);
DFFARX1 I_20544 (I351768,I2507,I351321,I351310,);
nor I_20545 (I351799,I146715,I146700);
or I_20546 (I351301,I351548,I351799);
nor I_20547 (I351292,I351681,I351799);
or I_20548 (I351295,I351415,I351799);
DFFARX1 I_20549 (I351799,I2507,I351321,I351313,);
not I_20550 (I351899,I2514);
DFFARX1 I_20551 (I214361,I2507,I351899,I351925,);
not I_20552 (I351933,I351925);
nand I_20553 (I351950,I214364,I214340);
and I_20554 (I351967,I351950,I214337);
DFFARX1 I_20555 (I351967,I2507,I351899,I351993,);
not I_20556 (I352001,I214343);
DFFARX1 I_20557 (I214337,I2507,I351899,I352027,);
not I_20558 (I352035,I352027);
nor I_20559 (I352052,I352035,I351933);
and I_20560 (I352069,I352052,I214343);
nor I_20561 (I352086,I352035,I352001);
nor I_20562 (I351882,I351993,I352086);
DFFARX1 I_20563 (I214346,I2507,I351899,I352126,);
nor I_20564 (I352134,I352126,I351993);
not I_20565 (I352151,I352134);
not I_20566 (I352168,I352126);
nor I_20567 (I352185,I352168,I352069);
DFFARX1 I_20568 (I352185,I2507,I351899,I351885,);
nand I_20569 (I352216,I214349,I214358);
and I_20570 (I352233,I352216,I214355);
DFFARX1 I_20571 (I352233,I2507,I351899,I352259,);
nor I_20572 (I352267,I352259,I352126);
DFFARX1 I_20573 (I352267,I2507,I351899,I351867,);
nand I_20574 (I352298,I352259,I352168);
nand I_20575 (I351876,I352151,I352298);
not I_20576 (I352329,I352259);
nor I_20577 (I352346,I352329,I352069);
DFFARX1 I_20578 (I352346,I2507,I351899,I351888,);
nor I_20579 (I352377,I214352,I214358);
or I_20580 (I351879,I352126,I352377);
nor I_20581 (I351870,I352259,I352377);
or I_20582 (I351873,I351993,I352377);
DFFARX1 I_20583 (I352377,I2507,I351899,I351891,);
not I_20584 (I352477,I2514);
DFFARX1 I_20585 (I65182,I2507,I352477,I352503,);
not I_20586 (I352511,I352503);
nand I_20587 (I352528,I65191,I65200);
and I_20588 (I352545,I352528,I65179);
DFFARX1 I_20589 (I352545,I2507,I352477,I352571,);
not I_20590 (I352579,I65182);
DFFARX1 I_20591 (I65197,I2507,I352477,I352605,);
not I_20592 (I352613,I352605);
nor I_20593 (I352630,I352613,I352511);
and I_20594 (I352647,I352630,I65182);
nor I_20595 (I352664,I352613,I352579);
nor I_20596 (I352460,I352571,I352664);
DFFARX1 I_20597 (I65188,I2507,I352477,I352704,);
nor I_20598 (I352712,I352704,I352571);
not I_20599 (I352729,I352712);
not I_20600 (I352746,I352704);
nor I_20601 (I352763,I352746,I352647);
DFFARX1 I_20602 (I352763,I2507,I352477,I352463,);
nand I_20603 (I352794,I65203,I65179);
and I_20604 (I352811,I352794,I65185);
DFFARX1 I_20605 (I352811,I2507,I352477,I352837,);
nor I_20606 (I352845,I352837,I352704);
DFFARX1 I_20607 (I352845,I2507,I352477,I352445,);
nand I_20608 (I352876,I352837,I352746);
nand I_20609 (I352454,I352729,I352876);
not I_20610 (I352907,I352837);
nor I_20611 (I352924,I352907,I352647);
DFFARX1 I_20612 (I352924,I2507,I352477,I352466,);
nor I_20613 (I352955,I65194,I65179);
or I_20614 (I352457,I352704,I352955);
nor I_20615 (I352448,I352837,I352955);
or I_20616 (I352451,I352571,I352955);
DFFARX1 I_20617 (I352955,I2507,I352477,I352469,);
not I_20618 (I353055,I2514);
DFFARX1 I_20619 (I712685,I2507,I353055,I353081,);
not I_20620 (I353089,I353081);
nand I_20621 (I353106,I712670,I712658);
and I_20622 (I353123,I353106,I712673);
DFFARX1 I_20623 (I353123,I2507,I353055,I353149,);
not I_20624 (I353157,I712658);
DFFARX1 I_20625 (I712676,I2507,I353055,I353183,);
not I_20626 (I353191,I353183);
nor I_20627 (I353208,I353191,I353089);
and I_20628 (I353225,I353208,I712658);
nor I_20629 (I353242,I353191,I353157);
nor I_20630 (I353038,I353149,I353242);
DFFARX1 I_20631 (I712664,I2507,I353055,I353282,);
nor I_20632 (I353290,I353282,I353149);
not I_20633 (I353307,I353290);
not I_20634 (I353324,I353282);
nor I_20635 (I353341,I353324,I353225);
DFFARX1 I_20636 (I353341,I2507,I353055,I353041,);
nand I_20637 (I353372,I712661,I712667);
and I_20638 (I353389,I353372,I712682);
DFFARX1 I_20639 (I353389,I2507,I353055,I353415,);
nor I_20640 (I353423,I353415,I353282);
DFFARX1 I_20641 (I353423,I2507,I353055,I353023,);
nand I_20642 (I353454,I353415,I353324);
nand I_20643 (I353032,I353307,I353454);
not I_20644 (I353485,I353415);
nor I_20645 (I353502,I353485,I353225);
DFFARX1 I_20646 (I353502,I2507,I353055,I353044,);
nor I_20647 (I353533,I712679,I712667);
or I_20648 (I353035,I353282,I353533);
nor I_20649 (I353026,I353415,I353533);
or I_20650 (I353029,I353149,I353533);
DFFARX1 I_20651 (I353533,I2507,I353055,I353047,);
not I_20652 (I353633,I2514);
DFFARX1 I_20653 (I583833,I2507,I353633,I353659,);
not I_20654 (I353667,I353659);
nand I_20655 (I353684,I583815,I583827);
and I_20656 (I353701,I353684,I583830);
DFFARX1 I_20657 (I353701,I2507,I353633,I353727,);
not I_20658 (I353735,I583824);
DFFARX1 I_20659 (I583821,I2507,I353633,I353761,);
not I_20660 (I353769,I353761);
nor I_20661 (I353786,I353769,I353667);
and I_20662 (I353803,I353786,I583824);
nor I_20663 (I353820,I353769,I353735);
nor I_20664 (I353616,I353727,I353820);
DFFARX1 I_20665 (I583839,I2507,I353633,I353860,);
nor I_20666 (I353868,I353860,I353727);
not I_20667 (I353885,I353868);
not I_20668 (I353902,I353860);
nor I_20669 (I353919,I353902,I353803);
DFFARX1 I_20670 (I353919,I2507,I353633,I353619,);
nand I_20671 (I353950,I583818,I583818);
and I_20672 (I353967,I353950,I583815);
DFFARX1 I_20673 (I353967,I2507,I353633,I353993,);
nor I_20674 (I354001,I353993,I353860);
DFFARX1 I_20675 (I354001,I2507,I353633,I353601,);
nand I_20676 (I354032,I353993,I353902);
nand I_20677 (I353610,I353885,I354032);
not I_20678 (I354063,I353993);
nor I_20679 (I354080,I354063,I353803);
DFFARX1 I_20680 (I354080,I2507,I353633,I353622,);
nor I_20681 (I354111,I583836,I583818);
or I_20682 (I353613,I353860,I354111);
nor I_20683 (I353604,I353993,I354111);
or I_20684 (I353607,I353727,I354111);
DFFARX1 I_20685 (I354111,I2507,I353633,I353625,);
not I_20686 (I354211,I2514);
DFFARX1 I_20687 (I230241,I2507,I354211,I354237,);
not I_20688 (I354245,I354237);
nand I_20689 (I354262,I230232,I230250);
and I_20690 (I354279,I354262,I230253);
DFFARX1 I_20691 (I354279,I2507,I354211,I354305,);
not I_20692 (I354313,I230247);
DFFARX1 I_20693 (I230235,I2507,I354211,I354339,);
not I_20694 (I354347,I354339);
nor I_20695 (I354364,I354347,I354245);
and I_20696 (I354381,I354364,I230247);
nor I_20697 (I354398,I354347,I354313);
nor I_20698 (I354194,I354305,I354398);
DFFARX1 I_20699 (I230244,I2507,I354211,I354438,);
nor I_20700 (I354446,I354438,I354305);
not I_20701 (I354463,I354446);
not I_20702 (I354480,I354438);
nor I_20703 (I354497,I354480,I354381);
DFFARX1 I_20704 (I354497,I2507,I354211,I354197,);
nand I_20705 (I354528,I230259,I230256);
and I_20706 (I354545,I354528,I230238);
DFFARX1 I_20707 (I354545,I2507,I354211,I354571,);
nor I_20708 (I354579,I354571,I354438);
DFFARX1 I_20709 (I354579,I2507,I354211,I354179,);
nand I_20710 (I354610,I354571,I354480);
nand I_20711 (I354188,I354463,I354610);
not I_20712 (I354641,I354571);
nor I_20713 (I354658,I354641,I354381);
DFFARX1 I_20714 (I354658,I2507,I354211,I354200,);
nor I_20715 (I354689,I230232,I230256);
or I_20716 (I354191,I354438,I354689);
nor I_20717 (I354182,I354571,I354689);
or I_20718 (I354185,I354305,I354689);
DFFARX1 I_20719 (I354689,I2507,I354211,I354203,);
not I_20720 (I354789,I2514);
DFFARX1 I_20721 (I47791,I2507,I354789,I354815,);
not I_20722 (I354823,I354815);
nand I_20723 (I354840,I47800,I47809);
and I_20724 (I354857,I354840,I47788);
DFFARX1 I_20725 (I354857,I2507,I354789,I354883,);
not I_20726 (I354891,I47791);
DFFARX1 I_20727 (I47806,I2507,I354789,I354917,);
not I_20728 (I354925,I354917);
nor I_20729 (I354942,I354925,I354823);
and I_20730 (I354959,I354942,I47791);
nor I_20731 (I354976,I354925,I354891);
nor I_20732 (I354772,I354883,I354976);
DFFARX1 I_20733 (I47797,I2507,I354789,I355016,);
nor I_20734 (I355024,I355016,I354883);
not I_20735 (I355041,I355024);
not I_20736 (I355058,I355016);
nor I_20737 (I355075,I355058,I354959);
DFFARX1 I_20738 (I355075,I2507,I354789,I354775,);
nand I_20739 (I355106,I47812,I47788);
and I_20740 (I355123,I355106,I47794);
DFFARX1 I_20741 (I355123,I2507,I354789,I355149,);
nor I_20742 (I355157,I355149,I355016);
DFFARX1 I_20743 (I355157,I2507,I354789,I354757,);
nand I_20744 (I355188,I355149,I355058);
nand I_20745 (I354766,I355041,I355188);
not I_20746 (I355219,I355149);
nor I_20747 (I355236,I355219,I354959);
DFFARX1 I_20748 (I355236,I2507,I354789,I354778,);
nor I_20749 (I355267,I47803,I47788);
or I_20750 (I354769,I355016,I355267);
nor I_20751 (I354760,I355149,I355267);
or I_20752 (I354763,I354883,I355267);
DFFARX1 I_20753 (I355267,I2507,I354789,I354781,);
not I_20754 (I355367,I2514);
DFFARX1 I_20755 (I84231,I2507,I355367,I355393,);
not I_20756 (I355401,I355393);
nand I_20757 (I355418,I84246,I84219);
and I_20758 (I355435,I355418,I84234);
DFFARX1 I_20759 (I355435,I2507,I355367,I355461,);
not I_20760 (I355469,I84237);
DFFARX1 I_20761 (I84222,I2507,I355367,I355495,);
not I_20762 (I355503,I355495);
nor I_20763 (I355520,I355503,I355401);
and I_20764 (I355537,I355520,I84237);
nor I_20765 (I355554,I355503,I355469);
nor I_20766 (I355350,I355461,I355554);
DFFARX1 I_20767 (I84228,I2507,I355367,I355594,);
nor I_20768 (I355602,I355594,I355461);
not I_20769 (I355619,I355602);
not I_20770 (I355636,I355594);
nor I_20771 (I355653,I355636,I355537);
DFFARX1 I_20772 (I355653,I2507,I355367,I355353,);
nand I_20773 (I355684,I84243,I84225);
and I_20774 (I355701,I355684,I84240);
DFFARX1 I_20775 (I355701,I2507,I355367,I355727,);
nor I_20776 (I355735,I355727,I355594);
DFFARX1 I_20777 (I355735,I2507,I355367,I355335,);
nand I_20778 (I355766,I355727,I355636);
nand I_20779 (I355344,I355619,I355766);
not I_20780 (I355797,I355727);
nor I_20781 (I355814,I355797,I355537);
DFFARX1 I_20782 (I355814,I2507,I355367,I355356,);
nor I_20783 (I355845,I84219,I84225);
or I_20784 (I355347,I355594,I355845);
nor I_20785 (I355338,I355727,I355845);
or I_20786 (I355341,I355461,I355845);
DFFARX1 I_20787 (I355845,I2507,I355367,I355359,);
not I_20788 (I355945,I2514);
DFFARX1 I_20789 (I127059,I2507,I355945,I355971,);
not I_20790 (I355979,I355971);
nand I_20791 (I355996,I127062,I127083);
and I_20792 (I356013,I355996,I127071);
DFFARX1 I_20793 (I356013,I2507,I355945,I356039,);
not I_20794 (I356047,I127068);
DFFARX1 I_20795 (I127059,I2507,I355945,I356073,);
not I_20796 (I356081,I356073);
nor I_20797 (I356098,I356081,I355979);
and I_20798 (I356115,I356098,I127068);
nor I_20799 (I356132,I356081,I356047);
nor I_20800 (I355928,I356039,I356132);
DFFARX1 I_20801 (I127077,I2507,I355945,I356172,);
nor I_20802 (I356180,I356172,I356039);
not I_20803 (I356197,I356180);
not I_20804 (I356214,I356172);
nor I_20805 (I356231,I356214,I356115);
DFFARX1 I_20806 (I356231,I2507,I355945,I355931,);
nand I_20807 (I356262,I127062,I127065);
and I_20808 (I356279,I356262,I127074);
DFFARX1 I_20809 (I356279,I2507,I355945,I356305,);
nor I_20810 (I356313,I356305,I356172);
DFFARX1 I_20811 (I356313,I2507,I355945,I355913,);
nand I_20812 (I356344,I356305,I356214);
nand I_20813 (I355922,I356197,I356344);
not I_20814 (I356375,I356305);
nor I_20815 (I356392,I356375,I356115);
DFFARX1 I_20816 (I356392,I2507,I355945,I355934,);
nor I_20817 (I356423,I127080,I127065);
or I_20818 (I355925,I356172,I356423);
nor I_20819 (I355916,I356305,I356423);
or I_20820 (I355919,I356039,I356423);
DFFARX1 I_20821 (I356423,I2507,I355945,I355937,);
not I_20822 (I356523,I2514);
DFFARX1 I_20823 (I253633,I2507,I356523,I356549,);
not I_20824 (I356557,I356549);
nand I_20825 (I356574,I253624,I253642);
and I_20826 (I356591,I356574,I253645);
DFFARX1 I_20827 (I356591,I2507,I356523,I356617,);
not I_20828 (I356625,I253639);
DFFARX1 I_20829 (I253627,I2507,I356523,I356651,);
not I_20830 (I356659,I356651);
nor I_20831 (I356676,I356659,I356557);
and I_20832 (I356693,I356676,I253639);
nor I_20833 (I356710,I356659,I356625);
nor I_20834 (I356506,I356617,I356710);
DFFARX1 I_20835 (I253636,I2507,I356523,I356750,);
nor I_20836 (I356758,I356750,I356617);
not I_20837 (I356775,I356758);
not I_20838 (I356792,I356750);
nor I_20839 (I356809,I356792,I356693);
DFFARX1 I_20840 (I356809,I2507,I356523,I356509,);
nand I_20841 (I356840,I253651,I253648);
and I_20842 (I356857,I356840,I253630);
DFFARX1 I_20843 (I356857,I2507,I356523,I356883,);
nor I_20844 (I356891,I356883,I356750);
DFFARX1 I_20845 (I356891,I2507,I356523,I356491,);
nand I_20846 (I356922,I356883,I356792);
nand I_20847 (I356500,I356775,I356922);
not I_20848 (I356953,I356883);
nor I_20849 (I356970,I356953,I356693);
DFFARX1 I_20850 (I356970,I2507,I356523,I356512,);
nor I_20851 (I357001,I253624,I253648);
or I_20852 (I356503,I356750,I357001);
nor I_20853 (I356494,I356883,I357001);
or I_20854 (I356497,I356617,I357001);
DFFARX1 I_20855 (I357001,I2507,I356523,I356515,);
not I_20856 (I357101,I2514);
DFFARX1 I_20857 (I24612,I2507,I357101,I357127,);
not I_20858 (I357135,I357127);
nand I_20859 (I357152,I24609,I24600);
and I_20860 (I357169,I357152,I24600);
DFFARX1 I_20861 (I357169,I2507,I357101,I357195,);
not I_20862 (I357203,I24603);
DFFARX1 I_20863 (I24618,I2507,I357101,I357229,);
not I_20864 (I357237,I357229);
nor I_20865 (I357254,I357237,I357135);
and I_20866 (I357271,I357254,I24603);
nor I_20867 (I357288,I357237,I357203);
nor I_20868 (I357084,I357195,I357288);
DFFARX1 I_20869 (I24603,I2507,I357101,I357328,);
nor I_20870 (I357336,I357328,I357195);
not I_20871 (I357353,I357336);
not I_20872 (I357370,I357328);
nor I_20873 (I357387,I357370,I357271);
DFFARX1 I_20874 (I357387,I2507,I357101,I357087,);
nand I_20875 (I357418,I24621,I24606);
and I_20876 (I357435,I357418,I24624);
DFFARX1 I_20877 (I357435,I2507,I357101,I357461,);
nor I_20878 (I357469,I357461,I357328);
DFFARX1 I_20879 (I357469,I2507,I357101,I357069,);
nand I_20880 (I357500,I357461,I357370);
nand I_20881 (I357078,I357353,I357500);
not I_20882 (I357531,I357461);
nor I_20883 (I357548,I357531,I357271);
DFFARX1 I_20884 (I357548,I2507,I357101,I357090,);
nor I_20885 (I357579,I24615,I24606);
or I_20886 (I357081,I357328,I357579);
nor I_20887 (I357072,I357461,I357579);
or I_20888 (I357075,I357195,I357579);
DFFARX1 I_20889 (I357579,I2507,I357101,I357093,);
not I_20890 (I357679,I2514);
DFFARX1 I_20891 (I686663,I2507,I357679,I357705,);
not I_20892 (I357713,I357705);
nand I_20893 (I357730,I686651,I686669);
and I_20894 (I357747,I357730,I686660);
DFFARX1 I_20895 (I357747,I2507,I357679,I357773,);
not I_20896 (I357781,I686675);
DFFARX1 I_20897 (I686672,I2507,I357679,I357807,);
not I_20898 (I357815,I357807);
nor I_20899 (I357832,I357815,I357713);
and I_20900 (I357849,I357832,I686675);
nor I_20901 (I357866,I357815,I357781);
nor I_20902 (I357662,I357773,I357866);
DFFARX1 I_20903 (I686654,I2507,I357679,I357906,);
nor I_20904 (I357914,I357906,I357773);
not I_20905 (I357931,I357914);
not I_20906 (I357948,I357906);
nor I_20907 (I357965,I357948,I357849);
DFFARX1 I_20908 (I357965,I2507,I357679,I357665,);
nand I_20909 (I357996,I686648,I686648);
and I_20910 (I358013,I357996,I686657);
DFFARX1 I_20911 (I358013,I2507,I357679,I358039,);
nor I_20912 (I358047,I358039,I357906);
DFFARX1 I_20913 (I358047,I2507,I357679,I357647,);
nand I_20914 (I358078,I358039,I357948);
nand I_20915 (I357656,I357931,I358078);
not I_20916 (I358109,I358039);
nor I_20917 (I358126,I358109,I357849);
DFFARX1 I_20918 (I358126,I2507,I357679,I357668,);
nor I_20919 (I358157,I686666,I686648);
or I_20920 (I357659,I357906,I358157);
nor I_20921 (I357650,I358039,I358157);
or I_20922 (I357653,I357773,I358157);
DFFARX1 I_20923 (I358157,I2507,I357679,I357671,);
not I_20924 (I358257,I2514);
DFFARX1 I_20925 (I168512,I2507,I358257,I358283,);
not I_20926 (I358291,I358283);
nand I_20927 (I358308,I168515,I168491);
and I_20928 (I358325,I358308,I168488);
DFFARX1 I_20929 (I358325,I2507,I358257,I358351,);
not I_20930 (I358359,I168494);
DFFARX1 I_20931 (I168488,I2507,I358257,I358385,);
not I_20932 (I358393,I358385);
nor I_20933 (I358410,I358393,I358291);
and I_20934 (I358427,I358410,I168494);
nor I_20935 (I358444,I358393,I358359);
nor I_20936 (I358240,I358351,I358444);
DFFARX1 I_20937 (I168497,I2507,I358257,I358484,);
nor I_20938 (I358492,I358484,I358351);
not I_20939 (I358509,I358492);
not I_20940 (I358526,I358484);
nor I_20941 (I358543,I358526,I358427);
DFFARX1 I_20942 (I358543,I2507,I358257,I358243,);
nand I_20943 (I358574,I168500,I168509);
and I_20944 (I358591,I358574,I168506);
DFFARX1 I_20945 (I358591,I2507,I358257,I358617,);
nor I_20946 (I358625,I358617,I358484);
DFFARX1 I_20947 (I358625,I2507,I358257,I358225,);
nand I_20948 (I358656,I358617,I358526);
nand I_20949 (I358234,I358509,I358656);
not I_20950 (I358687,I358617);
nor I_20951 (I358704,I358687,I358427);
DFFARX1 I_20952 (I358704,I2507,I358257,I358246,);
nor I_20953 (I358735,I168503,I168509);
or I_20954 (I358237,I358484,I358735);
nor I_20955 (I358228,I358617,I358735);
or I_20956 (I358231,I358351,I358735);
DFFARX1 I_20957 (I358735,I2507,I358257,I358249,);
not I_20958 (I358835,I2514);
DFFARX1 I_20959 (I728750,I2507,I358835,I358861,);
not I_20960 (I358869,I358861);
nand I_20961 (I358886,I728735,I728723);
and I_20962 (I358903,I358886,I728738);
DFFARX1 I_20963 (I358903,I2507,I358835,I358929,);
not I_20964 (I358937,I728723);
DFFARX1 I_20965 (I728741,I2507,I358835,I358963,);
not I_20966 (I358971,I358963);
nor I_20967 (I358988,I358971,I358869);
and I_20968 (I359005,I358988,I728723);
nor I_20969 (I359022,I358971,I358937);
nor I_20970 (I358818,I358929,I359022);
DFFARX1 I_20971 (I728729,I2507,I358835,I359062,);
nor I_20972 (I359070,I359062,I358929);
not I_20973 (I359087,I359070);
not I_20974 (I359104,I359062);
nor I_20975 (I359121,I359104,I359005);
DFFARX1 I_20976 (I359121,I2507,I358835,I358821,);
nand I_20977 (I359152,I728726,I728732);
and I_20978 (I359169,I359152,I728747);
DFFARX1 I_20979 (I359169,I2507,I358835,I359195,);
nor I_20980 (I359203,I359195,I359062);
DFFARX1 I_20981 (I359203,I2507,I358835,I358803,);
nand I_20982 (I359234,I359195,I359104);
nand I_20983 (I358812,I359087,I359234);
not I_20984 (I359265,I359195);
nor I_20985 (I359282,I359265,I359005);
DFFARX1 I_20986 (I359282,I2507,I358835,I358824,);
nor I_20987 (I359313,I728744,I728732);
or I_20988 (I358815,I359062,I359313);
nor I_20989 (I358806,I359195,I359313);
or I_20990 (I358809,I358929,I359313);
DFFARX1 I_20991 (I359313,I2507,I358835,I358827,);
not I_20992 (I359413,I2514);
DFFARX1 I_20993 (I624293,I2507,I359413,I359439,);
not I_20994 (I359447,I359439);
nand I_20995 (I359464,I624275,I624287);
and I_20996 (I359481,I359464,I624290);
DFFARX1 I_20997 (I359481,I2507,I359413,I359507,);
not I_20998 (I359515,I624284);
DFFARX1 I_20999 (I624281,I2507,I359413,I359541,);
not I_21000 (I359549,I359541);
nor I_21001 (I359566,I359549,I359447);
and I_21002 (I359583,I359566,I624284);
nor I_21003 (I359600,I359549,I359515);
nor I_21004 (I359396,I359507,I359600);
DFFARX1 I_21005 (I624299,I2507,I359413,I359640,);
nor I_21006 (I359648,I359640,I359507);
not I_21007 (I359665,I359648);
not I_21008 (I359682,I359640);
nor I_21009 (I359699,I359682,I359583);
DFFARX1 I_21010 (I359699,I2507,I359413,I359399,);
nand I_21011 (I359730,I624278,I624278);
and I_21012 (I359747,I359730,I624275);
DFFARX1 I_21013 (I359747,I2507,I359413,I359773,);
nor I_21014 (I359781,I359773,I359640);
DFFARX1 I_21015 (I359781,I2507,I359413,I359381,);
nand I_21016 (I359812,I359773,I359682);
nand I_21017 (I359390,I359665,I359812);
not I_21018 (I359843,I359773);
nor I_21019 (I359860,I359843,I359583);
DFFARX1 I_21020 (I359860,I2507,I359413,I359402,);
nor I_21021 (I359891,I624296,I624278);
or I_21022 (I359393,I359640,I359891);
nor I_21023 (I359384,I359773,I359891);
or I_21024 (I359387,I359507,I359891);
DFFARX1 I_21025 (I359891,I2507,I359413,I359405,);
not I_21026 (I359991,I2514);
DFFARX1 I_21027 (I141339,I2507,I359991,I360017,);
not I_21028 (I360025,I360017);
nand I_21029 (I360042,I141342,I141363);
and I_21030 (I360059,I360042,I141351);
DFFARX1 I_21031 (I360059,I2507,I359991,I360085,);
not I_21032 (I360093,I141348);
DFFARX1 I_21033 (I141339,I2507,I359991,I360119,);
not I_21034 (I360127,I360119);
nor I_21035 (I360144,I360127,I360025);
and I_21036 (I360161,I360144,I141348);
nor I_21037 (I360178,I360127,I360093);
nor I_21038 (I359974,I360085,I360178);
DFFARX1 I_21039 (I141357,I2507,I359991,I360218,);
nor I_21040 (I360226,I360218,I360085);
not I_21041 (I360243,I360226);
not I_21042 (I360260,I360218);
nor I_21043 (I360277,I360260,I360161);
DFFARX1 I_21044 (I360277,I2507,I359991,I359977,);
nand I_21045 (I360308,I141342,I141345);
and I_21046 (I360325,I360308,I141354);
DFFARX1 I_21047 (I360325,I2507,I359991,I360351,);
nor I_21048 (I360359,I360351,I360218);
DFFARX1 I_21049 (I360359,I2507,I359991,I359959,);
nand I_21050 (I360390,I360351,I360260);
nand I_21051 (I359968,I360243,I360390);
not I_21052 (I360421,I360351);
nor I_21053 (I360438,I360421,I360161);
DFFARX1 I_21054 (I360438,I2507,I359991,I359980,);
nor I_21055 (I360469,I141360,I141345);
or I_21056 (I359971,I360218,I360469);
nor I_21057 (I359962,I360351,I360469);
or I_21058 (I359965,I360085,I360469);
DFFARX1 I_21059 (I360469,I2507,I359991,I359983,);
not I_21060 (I360569,I2514);
DFFARX1 I_21061 (I249281,I2507,I360569,I360595,);
not I_21062 (I360603,I360595);
nand I_21063 (I360620,I249272,I249290);
and I_21064 (I360637,I360620,I249293);
DFFARX1 I_21065 (I360637,I2507,I360569,I360663,);
not I_21066 (I360671,I249287);
DFFARX1 I_21067 (I249275,I2507,I360569,I360697,);
not I_21068 (I360705,I360697);
nor I_21069 (I360722,I360705,I360603);
and I_21070 (I360739,I360722,I249287);
nor I_21071 (I360756,I360705,I360671);
nor I_21072 (I360552,I360663,I360756);
DFFARX1 I_21073 (I249284,I2507,I360569,I360796,);
nor I_21074 (I360804,I360796,I360663);
not I_21075 (I360821,I360804);
not I_21076 (I360838,I360796);
nor I_21077 (I360855,I360838,I360739);
DFFARX1 I_21078 (I360855,I2507,I360569,I360555,);
nand I_21079 (I360886,I249299,I249296);
and I_21080 (I360903,I360886,I249278);
DFFARX1 I_21081 (I360903,I2507,I360569,I360929,);
nor I_21082 (I360937,I360929,I360796);
DFFARX1 I_21083 (I360937,I2507,I360569,I360537,);
nand I_21084 (I360968,I360929,I360838);
nand I_21085 (I360546,I360821,I360968);
not I_21086 (I360999,I360929);
nor I_21087 (I361016,I360999,I360739);
DFFARX1 I_21088 (I361016,I2507,I360569,I360558,);
nor I_21089 (I361047,I249272,I249296);
or I_21090 (I360549,I360796,I361047);
nor I_21091 (I360540,I360929,I361047);
or I_21092 (I360543,I360663,I361047);
DFFARX1 I_21093 (I361047,I2507,I360569,I360561,);
not I_21094 (I361147,I2514);
DFFARX1 I_21095 (I46737,I2507,I361147,I361173,);
not I_21096 (I361181,I361173);
nand I_21097 (I361198,I46746,I46755);
and I_21098 (I361215,I361198,I46734);
DFFARX1 I_21099 (I361215,I2507,I361147,I361241,);
not I_21100 (I361249,I46737);
DFFARX1 I_21101 (I46752,I2507,I361147,I361275,);
not I_21102 (I361283,I361275);
nor I_21103 (I361300,I361283,I361181);
and I_21104 (I361317,I361300,I46737);
nor I_21105 (I361334,I361283,I361249);
nor I_21106 (I361130,I361241,I361334);
DFFARX1 I_21107 (I46743,I2507,I361147,I361374,);
nor I_21108 (I361382,I361374,I361241);
not I_21109 (I361399,I361382);
not I_21110 (I361416,I361374);
nor I_21111 (I361433,I361416,I361317);
DFFARX1 I_21112 (I361433,I2507,I361147,I361133,);
nand I_21113 (I361464,I46758,I46734);
and I_21114 (I361481,I361464,I46740);
DFFARX1 I_21115 (I361481,I2507,I361147,I361507,);
nor I_21116 (I361515,I361507,I361374);
DFFARX1 I_21117 (I361515,I2507,I361147,I361115,);
nand I_21118 (I361546,I361507,I361416);
nand I_21119 (I361124,I361399,I361546);
not I_21120 (I361577,I361507);
nor I_21121 (I361594,I361577,I361317);
DFFARX1 I_21122 (I361594,I2507,I361147,I361136,);
nor I_21123 (I361625,I46749,I46734);
or I_21124 (I361127,I361374,I361625);
nor I_21125 (I361118,I361507,I361625);
or I_21126 (I361121,I361241,I361625);
DFFARX1 I_21127 (I361625,I2507,I361147,I361139,);
not I_21128 (I361725,I2514);
DFFARX1 I_21129 (I592503,I2507,I361725,I361751,);
not I_21130 (I361759,I361751);
nand I_21131 (I361776,I592485,I592497);
and I_21132 (I361793,I361776,I592500);
DFFARX1 I_21133 (I361793,I2507,I361725,I361819,);
not I_21134 (I361827,I592494);
DFFARX1 I_21135 (I592491,I2507,I361725,I361853,);
not I_21136 (I361861,I361853);
nor I_21137 (I361878,I361861,I361759);
and I_21138 (I361895,I361878,I592494);
nor I_21139 (I361912,I361861,I361827);
nor I_21140 (I361708,I361819,I361912);
DFFARX1 I_21141 (I592509,I2507,I361725,I361952,);
nor I_21142 (I361960,I361952,I361819);
not I_21143 (I361977,I361960);
not I_21144 (I361994,I361952);
nor I_21145 (I362011,I361994,I361895);
DFFARX1 I_21146 (I362011,I2507,I361725,I361711,);
nand I_21147 (I362042,I592488,I592488);
and I_21148 (I362059,I362042,I592485);
DFFARX1 I_21149 (I362059,I2507,I361725,I362085,);
nor I_21150 (I362093,I362085,I361952);
DFFARX1 I_21151 (I362093,I2507,I361725,I361693,);
nand I_21152 (I362124,I362085,I361994);
nand I_21153 (I361702,I361977,I362124);
not I_21154 (I362155,I362085);
nor I_21155 (I362172,I362155,I361895);
DFFARX1 I_21156 (I362172,I2507,I361725,I361714,);
nor I_21157 (I362203,I592506,I592488);
or I_21158 (I361705,I361952,I362203);
nor I_21159 (I361696,I362085,I362203);
or I_21160 (I361699,I361819,I362203);
DFFARX1 I_21161 (I362203,I2507,I361725,I361717,);
not I_21162 (I362303,I2514);
DFFARX1 I_21163 (I138364,I2507,I362303,I362329,);
not I_21164 (I362337,I362329);
nand I_21165 (I362354,I138367,I138388);
and I_21166 (I362371,I362354,I138376);
DFFARX1 I_21167 (I362371,I2507,I362303,I362397,);
not I_21168 (I362405,I138373);
DFFARX1 I_21169 (I138364,I2507,I362303,I362431,);
not I_21170 (I362439,I362431);
nor I_21171 (I362456,I362439,I362337);
and I_21172 (I362473,I362456,I138373);
nor I_21173 (I362490,I362439,I362405);
nor I_21174 (I362286,I362397,I362490);
DFFARX1 I_21175 (I138382,I2507,I362303,I362530,);
nor I_21176 (I362538,I362530,I362397);
not I_21177 (I362555,I362538);
not I_21178 (I362572,I362530);
nor I_21179 (I362589,I362572,I362473);
DFFARX1 I_21180 (I362589,I2507,I362303,I362289,);
nand I_21181 (I362620,I138367,I138370);
and I_21182 (I362637,I362620,I138379);
DFFARX1 I_21183 (I362637,I2507,I362303,I362663,);
nor I_21184 (I362671,I362663,I362530);
DFFARX1 I_21185 (I362671,I2507,I362303,I362271,);
nand I_21186 (I362702,I362663,I362572);
nand I_21187 (I362280,I362555,I362702);
not I_21188 (I362733,I362663);
nor I_21189 (I362750,I362733,I362473);
DFFARX1 I_21190 (I362750,I2507,I362303,I362292,);
nor I_21191 (I362781,I138385,I138370);
or I_21192 (I362283,I362530,I362781);
nor I_21193 (I362274,I362663,I362781);
or I_21194 (I362277,I362397,I362781);
DFFARX1 I_21195 (I362781,I2507,I362303,I362295,);
not I_21196 (I362881,I2514);
DFFARX1 I_21197 (I48845,I2507,I362881,I362907,);
not I_21198 (I362915,I362907);
nand I_21199 (I362932,I48854,I48863);
and I_21200 (I362949,I362932,I48842);
DFFARX1 I_21201 (I362949,I2507,I362881,I362975,);
not I_21202 (I362983,I48845);
DFFARX1 I_21203 (I48860,I2507,I362881,I363009,);
not I_21204 (I363017,I363009);
nor I_21205 (I363034,I363017,I362915);
and I_21206 (I363051,I363034,I48845);
nor I_21207 (I363068,I363017,I362983);
nor I_21208 (I362864,I362975,I363068);
DFFARX1 I_21209 (I48851,I2507,I362881,I363108,);
nor I_21210 (I363116,I363108,I362975);
not I_21211 (I363133,I363116);
not I_21212 (I363150,I363108);
nor I_21213 (I363167,I363150,I363051);
DFFARX1 I_21214 (I363167,I2507,I362881,I362867,);
nand I_21215 (I363198,I48866,I48842);
and I_21216 (I363215,I363198,I48848);
DFFARX1 I_21217 (I363215,I2507,I362881,I363241,);
nor I_21218 (I363249,I363241,I363108);
DFFARX1 I_21219 (I363249,I2507,I362881,I362849,);
nand I_21220 (I363280,I363241,I363150);
nand I_21221 (I362858,I363133,I363280);
not I_21222 (I363311,I363241);
nor I_21223 (I363328,I363311,I363051);
DFFARX1 I_21224 (I363328,I2507,I362881,I362870,);
nor I_21225 (I363359,I48857,I48842);
or I_21226 (I362861,I363108,I363359);
nor I_21227 (I362852,I363241,I363359);
or I_21228 (I362855,I362975,I363359);
DFFARX1 I_21229 (I363359,I2507,I362881,I362873,);
not I_21230 (I363459,I2514);
DFFARX1 I_21231 (I346087,I2507,I363459,I363485,);
not I_21232 (I363493,I363485);
nand I_21233 (I363510,I346096,I346105);
and I_21234 (I363527,I363510,I346111);
DFFARX1 I_21235 (I363527,I2507,I363459,I363553,);
not I_21236 (I363561,I346108);
DFFARX1 I_21237 (I346093,I2507,I363459,I363587,);
not I_21238 (I363595,I363587);
nor I_21239 (I363612,I363595,I363493);
and I_21240 (I363629,I363612,I346108);
nor I_21241 (I363646,I363595,I363561);
nor I_21242 (I363442,I363553,I363646);
DFFARX1 I_21243 (I346102,I2507,I363459,I363686,);
nor I_21244 (I363694,I363686,I363553);
not I_21245 (I363711,I363694);
not I_21246 (I363728,I363686);
nor I_21247 (I363745,I363728,I363629);
DFFARX1 I_21248 (I363745,I2507,I363459,I363445,);
nand I_21249 (I363776,I346099,I346090);
and I_21250 (I363793,I363776,I346087);
DFFARX1 I_21251 (I363793,I2507,I363459,I363819,);
nor I_21252 (I363827,I363819,I363686);
DFFARX1 I_21253 (I363827,I2507,I363459,I363427,);
nand I_21254 (I363858,I363819,I363728);
nand I_21255 (I363436,I363711,I363858);
not I_21256 (I363889,I363819);
nor I_21257 (I363906,I363889,I363629);
DFFARX1 I_21258 (I363906,I2507,I363459,I363448,);
nor I_21259 (I363937,I346090,I346090);
or I_21260 (I363439,I363686,I363937);
nor I_21261 (I363430,I363819,I363937);
or I_21262 (I363433,I363553,I363937);
DFFARX1 I_21263 (I363937,I2507,I363459,I363451,);
not I_21264 (I364037,I2514);
DFFARX1 I_21265 (I36724,I2507,I364037,I364063,);
not I_21266 (I364071,I364063);
nand I_21267 (I364088,I36733,I36742);
and I_21268 (I364105,I364088,I36721);
DFFARX1 I_21269 (I364105,I2507,I364037,I364131,);
not I_21270 (I364139,I36724);
DFFARX1 I_21271 (I36739,I2507,I364037,I364165,);
not I_21272 (I364173,I364165);
nor I_21273 (I364190,I364173,I364071);
and I_21274 (I364207,I364190,I36724);
nor I_21275 (I364224,I364173,I364139);
nor I_21276 (I364020,I364131,I364224);
DFFARX1 I_21277 (I36730,I2507,I364037,I364264,);
nor I_21278 (I364272,I364264,I364131);
not I_21279 (I364289,I364272);
not I_21280 (I364306,I364264);
nor I_21281 (I364323,I364306,I364207);
DFFARX1 I_21282 (I364323,I2507,I364037,I364023,);
nand I_21283 (I364354,I36745,I36721);
and I_21284 (I364371,I364354,I36727);
DFFARX1 I_21285 (I364371,I2507,I364037,I364397,);
nor I_21286 (I364405,I364397,I364264);
DFFARX1 I_21287 (I364405,I2507,I364037,I364005,);
nand I_21288 (I364436,I364397,I364306);
nand I_21289 (I364014,I364289,I364436);
not I_21290 (I364467,I364397);
nor I_21291 (I364484,I364467,I364207);
DFFARX1 I_21292 (I364484,I2507,I364037,I364026,);
nor I_21293 (I364515,I36736,I36721);
or I_21294 (I364017,I364264,I364515);
nor I_21295 (I364008,I364397,I364515);
or I_21296 (I364011,I364131,I364515);
DFFARX1 I_21297 (I364515,I2507,I364037,I364029,);
not I_21298 (I364615,I2514);
DFFARX1 I_21299 (I32517,I2507,I364615,I364641,);
not I_21300 (I364649,I364641);
nand I_21301 (I364666,I32514,I32505);
and I_21302 (I364683,I364666,I32505);
DFFARX1 I_21303 (I364683,I2507,I364615,I364709,);
not I_21304 (I364717,I32508);
DFFARX1 I_21305 (I32523,I2507,I364615,I364743,);
not I_21306 (I364751,I364743);
nor I_21307 (I364768,I364751,I364649);
and I_21308 (I364785,I364768,I32508);
nor I_21309 (I364802,I364751,I364717);
nor I_21310 (I364598,I364709,I364802);
DFFARX1 I_21311 (I32508,I2507,I364615,I364842,);
nor I_21312 (I364850,I364842,I364709);
not I_21313 (I364867,I364850);
not I_21314 (I364884,I364842);
nor I_21315 (I364901,I364884,I364785);
DFFARX1 I_21316 (I364901,I2507,I364615,I364601,);
nand I_21317 (I364932,I32526,I32511);
and I_21318 (I364949,I364932,I32529);
DFFARX1 I_21319 (I364949,I2507,I364615,I364975,);
nor I_21320 (I364983,I364975,I364842);
DFFARX1 I_21321 (I364983,I2507,I364615,I364583,);
nand I_21322 (I365014,I364975,I364884);
nand I_21323 (I364592,I364867,I365014);
not I_21324 (I365045,I364975);
nor I_21325 (I365062,I365045,I364785);
DFFARX1 I_21326 (I365062,I2507,I364615,I364604,);
nor I_21327 (I365093,I32520,I32511);
or I_21328 (I364595,I364842,I365093);
nor I_21329 (I364586,I364975,I365093);
or I_21330 (I364589,I364709,I365093);
DFFARX1 I_21331 (I365093,I2507,I364615,I364607,);
not I_21332 (I365193,I2514);
DFFARX1 I_21333 (I252545,I2507,I365193,I365219,);
not I_21334 (I365227,I365219);
nand I_21335 (I365244,I252536,I252554);
and I_21336 (I365261,I365244,I252557);
DFFARX1 I_21337 (I365261,I2507,I365193,I365287,);
not I_21338 (I365295,I252551);
DFFARX1 I_21339 (I252539,I2507,I365193,I365321,);
not I_21340 (I365329,I365321);
nor I_21341 (I365346,I365329,I365227);
and I_21342 (I365363,I365346,I252551);
nor I_21343 (I365380,I365329,I365295);
nor I_21344 (I365176,I365287,I365380);
DFFARX1 I_21345 (I252548,I2507,I365193,I365420,);
nor I_21346 (I365428,I365420,I365287);
not I_21347 (I365445,I365428);
not I_21348 (I365462,I365420);
nor I_21349 (I365479,I365462,I365363);
DFFARX1 I_21350 (I365479,I2507,I365193,I365179,);
nand I_21351 (I365510,I252563,I252560);
and I_21352 (I365527,I365510,I252542);
DFFARX1 I_21353 (I365527,I2507,I365193,I365553,);
nor I_21354 (I365561,I365553,I365420);
DFFARX1 I_21355 (I365561,I2507,I365193,I365161,);
nand I_21356 (I365592,I365553,I365462);
nand I_21357 (I365170,I365445,I365592);
not I_21358 (I365623,I365553);
nor I_21359 (I365640,I365623,I365363);
DFFARX1 I_21360 (I365640,I2507,I365193,I365182,);
nor I_21361 (I365671,I252536,I252560);
or I_21362 (I365173,I365420,I365671);
nor I_21363 (I365164,I365553,I365671);
or I_21364 (I365167,I365287,I365671);
DFFARX1 I_21365 (I365671,I2507,I365193,I365185,);
not I_21366 (I365771,I2514);
DFFARX1 I_21367 (I277569,I2507,I365771,I365797,);
not I_21368 (I365805,I365797);
nand I_21369 (I365822,I277560,I277578);
and I_21370 (I365839,I365822,I277581);
DFFARX1 I_21371 (I365839,I2507,I365771,I365865,);
not I_21372 (I365873,I277575);
DFFARX1 I_21373 (I277563,I2507,I365771,I365899,);
not I_21374 (I365907,I365899);
nor I_21375 (I365924,I365907,I365805);
and I_21376 (I365941,I365924,I277575);
nor I_21377 (I365958,I365907,I365873);
nor I_21378 (I365754,I365865,I365958);
DFFARX1 I_21379 (I277572,I2507,I365771,I365998,);
nor I_21380 (I366006,I365998,I365865);
not I_21381 (I366023,I366006);
not I_21382 (I366040,I365998);
nor I_21383 (I366057,I366040,I365941);
DFFARX1 I_21384 (I366057,I2507,I365771,I365757,);
nand I_21385 (I366088,I277587,I277584);
and I_21386 (I366105,I366088,I277566);
DFFARX1 I_21387 (I366105,I2507,I365771,I366131,);
nor I_21388 (I366139,I366131,I365998);
DFFARX1 I_21389 (I366139,I2507,I365771,I365739,);
nand I_21390 (I366170,I366131,I366040);
nand I_21391 (I365748,I366023,I366170);
not I_21392 (I366201,I366131);
nor I_21393 (I366218,I366201,I365941);
DFFARX1 I_21394 (I366218,I2507,I365771,I365760,);
nor I_21395 (I366249,I277560,I277584);
or I_21396 (I365751,I365998,I366249);
nor I_21397 (I365742,I366131,I366249);
or I_21398 (I365745,I365865,I366249);
DFFARX1 I_21399 (I366249,I2507,I365771,I365763,);
not I_21400 (I366349,I2514);
DFFARX1 I_21401 (I658309,I2507,I366349,I366375,);
not I_21402 (I366383,I366375);
nand I_21403 (I366400,I658312,I658321);
and I_21404 (I366417,I366400,I658324);
DFFARX1 I_21405 (I366417,I2507,I366349,I366443,);
not I_21406 (I366451,I658333);
DFFARX1 I_21407 (I658315,I2507,I366349,I366477,);
not I_21408 (I366485,I366477);
nor I_21409 (I366502,I366485,I366383);
and I_21410 (I366519,I366502,I658333);
nor I_21411 (I366536,I366485,I366451);
nor I_21412 (I366332,I366443,I366536);
DFFARX1 I_21413 (I658312,I2507,I366349,I366576,);
nor I_21414 (I366584,I366576,I366443);
not I_21415 (I366601,I366584);
not I_21416 (I366618,I366576);
nor I_21417 (I366635,I366618,I366519);
DFFARX1 I_21418 (I366635,I2507,I366349,I366335,);
nand I_21419 (I366666,I658330,I658309);
and I_21420 (I366683,I366666,I658327);
DFFARX1 I_21421 (I366683,I2507,I366349,I366709,);
nor I_21422 (I366717,I366709,I366576);
DFFARX1 I_21423 (I366717,I2507,I366349,I366317,);
nand I_21424 (I366748,I366709,I366618);
nand I_21425 (I366326,I366601,I366748);
not I_21426 (I366779,I366709);
nor I_21427 (I366796,I366779,I366519);
DFFARX1 I_21428 (I366796,I2507,I366349,I366338,);
nor I_21429 (I366827,I658318,I658309);
or I_21430 (I366329,I366576,I366827);
nor I_21431 (I366320,I366709,I366827);
or I_21432 (I366323,I366443,I366827);
DFFARX1 I_21433 (I366827,I2507,I366349,I366341,);
not I_21434 (I366927,I2514);
DFFARX1 I_21435 (I702570,I2507,I366927,I366953,);
not I_21436 (I366961,I366953);
nand I_21437 (I366978,I702555,I702543);
and I_21438 (I366995,I366978,I702558);
DFFARX1 I_21439 (I366995,I2507,I366927,I367021,);
not I_21440 (I367029,I702543);
DFFARX1 I_21441 (I702561,I2507,I366927,I367055,);
not I_21442 (I367063,I367055);
nor I_21443 (I367080,I367063,I366961);
and I_21444 (I367097,I367080,I702543);
nor I_21445 (I367114,I367063,I367029);
nor I_21446 (I366910,I367021,I367114);
DFFARX1 I_21447 (I702549,I2507,I366927,I367154,);
nor I_21448 (I367162,I367154,I367021);
not I_21449 (I367179,I367162);
not I_21450 (I367196,I367154);
nor I_21451 (I367213,I367196,I367097);
DFFARX1 I_21452 (I367213,I2507,I366927,I366913,);
nand I_21453 (I367244,I702546,I702552);
and I_21454 (I367261,I367244,I702567);
DFFARX1 I_21455 (I367261,I2507,I366927,I367287,);
nor I_21456 (I367295,I367287,I367154);
DFFARX1 I_21457 (I367295,I2507,I366927,I366895,);
nand I_21458 (I367326,I367287,I367196);
nand I_21459 (I366904,I367179,I367326);
not I_21460 (I367357,I367287);
nor I_21461 (I367374,I367357,I367097);
DFFARX1 I_21462 (I367374,I2507,I366927,I366916,);
nor I_21463 (I367405,I702564,I702552);
or I_21464 (I366907,I367154,I367405);
nor I_21465 (I366898,I367287,I367405);
or I_21466 (I366901,I367021,I367405);
DFFARX1 I_21467 (I367405,I2507,I366927,I366919,);
not I_21468 (I367505,I2514);
DFFARX1 I_21469 (I549770,I2507,I367505,I367531,);
not I_21470 (I367539,I367531);
nand I_21471 (I367556,I549767,I549785);
and I_21472 (I367573,I367556,I549782);
DFFARX1 I_21473 (I367573,I2507,I367505,I367599,);
not I_21474 (I367607,I549764);
DFFARX1 I_21475 (I549767,I2507,I367505,I367633,);
not I_21476 (I367641,I367633);
nor I_21477 (I367658,I367641,I367539);
and I_21478 (I367675,I367658,I549764);
nor I_21479 (I367692,I367641,I367607);
nor I_21480 (I367488,I367599,I367692);
DFFARX1 I_21481 (I549776,I2507,I367505,I367732,);
nor I_21482 (I367740,I367732,I367599);
not I_21483 (I367757,I367740);
not I_21484 (I367774,I367732);
nor I_21485 (I367791,I367774,I367675);
DFFARX1 I_21486 (I367791,I2507,I367505,I367491,);
nand I_21487 (I367822,I549779,I549764);
and I_21488 (I367839,I367822,I549770);
DFFARX1 I_21489 (I367839,I2507,I367505,I367865,);
nor I_21490 (I367873,I367865,I367732);
DFFARX1 I_21491 (I367873,I2507,I367505,I367473,);
nand I_21492 (I367904,I367865,I367774);
nand I_21493 (I367482,I367757,I367904);
not I_21494 (I367935,I367865);
nor I_21495 (I367952,I367935,I367675);
DFFARX1 I_21496 (I367952,I2507,I367505,I367494,);
nor I_21497 (I367983,I549773,I549764);
or I_21498 (I367485,I367732,I367983);
nor I_21499 (I367476,I367865,I367983);
or I_21500 (I367479,I367599,I367983);
DFFARX1 I_21501 (I367983,I2507,I367505,I367497,);
not I_21502 (I368083,I2514);
DFFARX1 I_21503 (I307361,I2507,I368083,I368109,);
not I_21504 (I368117,I368109);
nand I_21505 (I368134,I307370,I307379);
and I_21506 (I368151,I368134,I307385);
DFFARX1 I_21507 (I368151,I2507,I368083,I368177,);
not I_21508 (I368185,I307382);
DFFARX1 I_21509 (I307367,I2507,I368083,I368211,);
not I_21510 (I368219,I368211);
nor I_21511 (I368236,I368219,I368117);
and I_21512 (I368253,I368236,I307382);
nor I_21513 (I368270,I368219,I368185);
nor I_21514 (I368066,I368177,I368270);
DFFARX1 I_21515 (I307376,I2507,I368083,I368310,);
nor I_21516 (I368318,I368310,I368177);
not I_21517 (I368335,I368318);
not I_21518 (I368352,I368310);
nor I_21519 (I368369,I368352,I368253);
DFFARX1 I_21520 (I368369,I2507,I368083,I368069,);
nand I_21521 (I368400,I307373,I307364);
and I_21522 (I368417,I368400,I307361);
DFFARX1 I_21523 (I368417,I2507,I368083,I368443,);
nor I_21524 (I368451,I368443,I368310);
DFFARX1 I_21525 (I368451,I2507,I368083,I368051,);
nand I_21526 (I368482,I368443,I368352);
nand I_21527 (I368060,I368335,I368482);
not I_21528 (I368513,I368443);
nor I_21529 (I368530,I368513,I368253);
DFFARX1 I_21530 (I368530,I2507,I368083,I368072,);
nor I_21531 (I368561,I307364,I307364);
or I_21532 (I368063,I368310,I368561);
nor I_21533 (I368054,I368443,I368561);
or I_21534 (I368057,I368177,I368561);
DFFARX1 I_21535 (I368561,I2507,I368083,I368075,);
not I_21536 (I368661,I2514);
DFFARX1 I_21537 (I492532,I2507,I368661,I368687,);
not I_21538 (I368695,I368687);
nand I_21539 (I368712,I492508,I492523);
and I_21540 (I368729,I368712,I492535);
DFFARX1 I_21541 (I368729,I2507,I368661,I368755,);
not I_21542 (I368763,I492520);
DFFARX1 I_21543 (I492511,I2507,I368661,I368789,);
not I_21544 (I368797,I368789);
nor I_21545 (I368814,I368797,I368695);
and I_21546 (I368831,I368814,I492520);
nor I_21547 (I368848,I368797,I368763);
nor I_21548 (I368644,I368755,I368848);
DFFARX1 I_21549 (I492508,I2507,I368661,I368888,);
nor I_21550 (I368896,I368888,I368755);
not I_21551 (I368913,I368896);
not I_21552 (I368930,I368888);
nor I_21553 (I368947,I368930,I368831);
DFFARX1 I_21554 (I368947,I2507,I368661,I368647,);
nand I_21555 (I368978,I492526,I492517);
and I_21556 (I368995,I368978,I492529);
DFFARX1 I_21557 (I368995,I2507,I368661,I369021,);
nor I_21558 (I369029,I369021,I368888);
DFFARX1 I_21559 (I369029,I2507,I368661,I368629,);
nand I_21560 (I369060,I369021,I368930);
nand I_21561 (I368638,I368913,I369060);
not I_21562 (I369091,I369021);
nor I_21563 (I369108,I369091,I368831);
DFFARX1 I_21564 (I369108,I2507,I368661,I368650,);
nor I_21565 (I369139,I492514,I492517);
or I_21566 (I368641,I368888,I369139);
nor I_21567 (I368632,I369021,I369139);
or I_21568 (I368635,I368755,I369139);
DFFARX1 I_21569 (I369139,I2507,I368661,I368653,);
not I_21570 (I369239,I2514);
DFFARX1 I_21571 (I328169,I2507,I369239,I369265,);
not I_21572 (I369273,I369265);
nand I_21573 (I369290,I328178,I328187);
and I_21574 (I369307,I369290,I328193);
DFFARX1 I_21575 (I369307,I2507,I369239,I369333,);
not I_21576 (I369341,I328190);
DFFARX1 I_21577 (I328175,I2507,I369239,I369367,);
not I_21578 (I369375,I369367);
nor I_21579 (I369392,I369375,I369273);
and I_21580 (I369409,I369392,I328190);
nor I_21581 (I369426,I369375,I369341);
nor I_21582 (I369222,I369333,I369426);
DFFARX1 I_21583 (I328184,I2507,I369239,I369466,);
nor I_21584 (I369474,I369466,I369333);
not I_21585 (I369491,I369474);
not I_21586 (I369508,I369466);
nor I_21587 (I369525,I369508,I369409);
DFFARX1 I_21588 (I369525,I2507,I369239,I369225,);
nand I_21589 (I369556,I328181,I328172);
and I_21590 (I369573,I369556,I328169);
DFFARX1 I_21591 (I369573,I2507,I369239,I369599,);
nor I_21592 (I369607,I369599,I369466);
DFFARX1 I_21593 (I369607,I2507,I369239,I369207,);
nand I_21594 (I369638,I369599,I369508);
nand I_21595 (I369216,I369491,I369638);
not I_21596 (I369669,I369599);
nor I_21597 (I369686,I369669,I369409);
DFFARX1 I_21598 (I369686,I2507,I369239,I369228,);
nor I_21599 (I369717,I328172,I328172);
or I_21600 (I369219,I369466,I369717);
nor I_21601 (I369210,I369599,I369717);
or I_21602 (I369213,I369333,I369717);
DFFARX1 I_21603 (I369717,I2507,I369239,I369231,);
not I_21604 (I369817,I2514);
DFFARX1 I_21605 (I245473,I2507,I369817,I369843,);
not I_21606 (I369851,I369843);
nand I_21607 (I369868,I245464,I245482);
and I_21608 (I369885,I369868,I245485);
DFFARX1 I_21609 (I369885,I2507,I369817,I369911,);
not I_21610 (I369919,I245479);
DFFARX1 I_21611 (I245467,I2507,I369817,I369945,);
not I_21612 (I369953,I369945);
nor I_21613 (I369970,I369953,I369851);
and I_21614 (I369987,I369970,I245479);
nor I_21615 (I370004,I369953,I369919);
nor I_21616 (I369800,I369911,I370004);
DFFARX1 I_21617 (I245476,I2507,I369817,I370044,);
nor I_21618 (I370052,I370044,I369911);
not I_21619 (I370069,I370052);
not I_21620 (I370086,I370044);
nor I_21621 (I370103,I370086,I369987);
DFFARX1 I_21622 (I370103,I2507,I369817,I369803,);
nand I_21623 (I370134,I245491,I245488);
and I_21624 (I370151,I370134,I245470);
DFFARX1 I_21625 (I370151,I2507,I369817,I370177,);
nor I_21626 (I370185,I370177,I370044);
DFFARX1 I_21627 (I370185,I2507,I369817,I369785,);
nand I_21628 (I370216,I370177,I370086);
nand I_21629 (I369794,I370069,I370216);
not I_21630 (I370247,I370177);
nor I_21631 (I370264,I370247,I369987);
DFFARX1 I_21632 (I370264,I2507,I369817,I369806,);
nor I_21633 (I370295,I245464,I245488);
or I_21634 (I369797,I370044,I370295);
nor I_21635 (I369788,I370177,I370295);
or I_21636 (I369791,I369911,I370295);
DFFARX1 I_21637 (I370295,I2507,I369817,I369809,);
not I_21638 (I370395,I2514);
DFFARX1 I_21639 (I580365,I2507,I370395,I370421,);
not I_21640 (I370429,I370421);
nand I_21641 (I370446,I580347,I580359);
and I_21642 (I370463,I370446,I580362);
DFFARX1 I_21643 (I370463,I2507,I370395,I370489,);
not I_21644 (I370497,I580356);
DFFARX1 I_21645 (I580353,I2507,I370395,I370523,);
not I_21646 (I370531,I370523);
nor I_21647 (I370548,I370531,I370429);
and I_21648 (I370565,I370548,I580356);
nor I_21649 (I370582,I370531,I370497);
nor I_21650 (I370378,I370489,I370582);
DFFARX1 I_21651 (I580371,I2507,I370395,I370622,);
nor I_21652 (I370630,I370622,I370489);
not I_21653 (I370647,I370630);
not I_21654 (I370664,I370622);
nor I_21655 (I370681,I370664,I370565);
DFFARX1 I_21656 (I370681,I2507,I370395,I370381,);
nand I_21657 (I370712,I580350,I580350);
and I_21658 (I370729,I370712,I580347);
DFFARX1 I_21659 (I370729,I2507,I370395,I370755,);
nor I_21660 (I370763,I370755,I370622);
DFFARX1 I_21661 (I370763,I2507,I370395,I370363,);
nand I_21662 (I370794,I370755,I370664);
nand I_21663 (I370372,I370647,I370794);
not I_21664 (I370825,I370755);
nor I_21665 (I370842,I370825,I370565);
DFFARX1 I_21666 (I370842,I2507,I370395,I370384,);
nor I_21667 (I370873,I580368,I580350);
or I_21668 (I370375,I370622,I370873);
nor I_21669 (I370366,I370755,I370873);
or I_21670 (I370369,I370489,I370873);
DFFARX1 I_21671 (I370873,I2507,I370395,I370387,);
not I_21672 (I370973,I2514);
DFFARX1 I_21673 (I23558,I2507,I370973,I370999,);
not I_21674 (I371007,I370999);
nand I_21675 (I371024,I23555,I23546);
and I_21676 (I371041,I371024,I23546);
DFFARX1 I_21677 (I371041,I2507,I370973,I371067,);
not I_21678 (I371075,I23549);
DFFARX1 I_21679 (I23564,I2507,I370973,I371101,);
not I_21680 (I371109,I371101);
nor I_21681 (I371126,I371109,I371007);
and I_21682 (I371143,I371126,I23549);
nor I_21683 (I371160,I371109,I371075);
nor I_21684 (I370956,I371067,I371160);
DFFARX1 I_21685 (I23549,I2507,I370973,I371200,);
nor I_21686 (I371208,I371200,I371067);
not I_21687 (I371225,I371208);
not I_21688 (I371242,I371200);
nor I_21689 (I371259,I371242,I371143);
DFFARX1 I_21690 (I371259,I2507,I370973,I370959,);
nand I_21691 (I371290,I23567,I23552);
and I_21692 (I371307,I371290,I23570);
DFFARX1 I_21693 (I371307,I2507,I370973,I371333,);
nor I_21694 (I371341,I371333,I371200);
DFFARX1 I_21695 (I371341,I2507,I370973,I370941,);
nand I_21696 (I371372,I371333,I371242);
nand I_21697 (I370950,I371225,I371372);
not I_21698 (I371403,I371333);
nor I_21699 (I371420,I371403,I371143);
DFFARX1 I_21700 (I371420,I2507,I370973,I370962,);
nor I_21701 (I371451,I23561,I23552);
or I_21702 (I370953,I371200,I371451);
nor I_21703 (I370944,I371333,I371451);
or I_21704 (I370947,I371067,I371451);
DFFARX1 I_21705 (I371451,I2507,I370973,I370965,);
not I_21706 (I371551,I2514);
DFFARX1 I_21707 (I488010,I2507,I371551,I371577,);
not I_21708 (I371585,I371577);
nand I_21709 (I371602,I487986,I488001);
and I_21710 (I371619,I371602,I488013);
DFFARX1 I_21711 (I371619,I2507,I371551,I371645,);
not I_21712 (I371653,I487998);
DFFARX1 I_21713 (I487989,I2507,I371551,I371679,);
not I_21714 (I371687,I371679);
nor I_21715 (I371704,I371687,I371585);
and I_21716 (I371721,I371704,I487998);
nor I_21717 (I371738,I371687,I371653);
nor I_21718 (I371534,I371645,I371738);
DFFARX1 I_21719 (I487986,I2507,I371551,I371778,);
nor I_21720 (I371786,I371778,I371645);
not I_21721 (I371803,I371786);
not I_21722 (I371820,I371778);
nor I_21723 (I371837,I371820,I371721);
DFFARX1 I_21724 (I371837,I2507,I371551,I371537,);
nand I_21725 (I371868,I488004,I487995);
and I_21726 (I371885,I371868,I488007);
DFFARX1 I_21727 (I371885,I2507,I371551,I371911,);
nor I_21728 (I371919,I371911,I371778);
DFFARX1 I_21729 (I371919,I2507,I371551,I371519,);
nand I_21730 (I371950,I371911,I371820);
nand I_21731 (I371528,I371803,I371950);
not I_21732 (I371981,I371911);
nor I_21733 (I371998,I371981,I371721);
DFFARX1 I_21734 (I371998,I2507,I371551,I371540,);
nor I_21735 (I372029,I487992,I487995);
or I_21736 (I371531,I371778,I372029);
nor I_21737 (I371522,I371911,I372029);
or I_21738 (I371525,I371645,I372029);
DFFARX1 I_21739 (I372029,I2507,I371551,I371543,);
not I_21740 (I372129,I2514);
DFFARX1 I_21741 (I476084,I2507,I372129,I372155,);
not I_21742 (I372163,I372155);
nand I_21743 (I372180,I476072,I476090);
and I_21744 (I372197,I372180,I476087);
DFFARX1 I_21745 (I372197,I2507,I372129,I372223,);
not I_21746 (I372231,I476078);
DFFARX1 I_21747 (I476075,I2507,I372129,I372257,);
not I_21748 (I372265,I372257);
nor I_21749 (I372282,I372265,I372163);
and I_21750 (I372299,I372282,I476078);
nor I_21751 (I372316,I372265,I372231);
nor I_21752 (I372112,I372223,I372316);
DFFARX1 I_21753 (I476069,I2507,I372129,I372356,);
nor I_21754 (I372364,I372356,I372223);
not I_21755 (I372381,I372364);
not I_21756 (I372398,I372356);
nor I_21757 (I372415,I372398,I372299);
DFFARX1 I_21758 (I372415,I2507,I372129,I372115,);
nand I_21759 (I372446,I476069,I476072);
and I_21760 (I372463,I372446,I476075);
DFFARX1 I_21761 (I372463,I2507,I372129,I372489,);
nor I_21762 (I372497,I372489,I372356);
DFFARX1 I_21763 (I372497,I2507,I372129,I372097,);
nand I_21764 (I372528,I372489,I372398);
nand I_21765 (I372106,I372381,I372528);
not I_21766 (I372559,I372489);
nor I_21767 (I372576,I372559,I372299);
DFFARX1 I_21768 (I372576,I2507,I372129,I372118,);
nor I_21769 (I372607,I476081,I476072);
or I_21770 (I372109,I372356,I372607);
nor I_21771 (I372100,I372489,I372607);
or I_21772 (I372103,I372223,I372607);
DFFARX1 I_21773 (I372607,I2507,I372129,I372121,);
not I_21774 (I372707,I2514);
DFFARX1 I_21775 (I188011,I2507,I372707,I372733,);
not I_21776 (I372741,I372733);
nand I_21777 (I372758,I188014,I187990);
and I_21778 (I372775,I372758,I187987);
DFFARX1 I_21779 (I372775,I2507,I372707,I372801,);
not I_21780 (I372809,I187993);
DFFARX1 I_21781 (I187987,I2507,I372707,I372835,);
not I_21782 (I372843,I372835);
nor I_21783 (I372860,I372843,I372741);
and I_21784 (I372877,I372860,I187993);
nor I_21785 (I372894,I372843,I372809);
nor I_21786 (I372690,I372801,I372894);
DFFARX1 I_21787 (I187996,I2507,I372707,I372934,);
nor I_21788 (I372942,I372934,I372801);
not I_21789 (I372959,I372942);
not I_21790 (I372976,I372934);
nor I_21791 (I372993,I372976,I372877);
DFFARX1 I_21792 (I372993,I2507,I372707,I372693,);
nand I_21793 (I373024,I187999,I188008);
and I_21794 (I373041,I373024,I188005);
DFFARX1 I_21795 (I373041,I2507,I372707,I373067,);
nor I_21796 (I373075,I373067,I372934);
DFFARX1 I_21797 (I373075,I2507,I372707,I372675,);
nand I_21798 (I373106,I373067,I372976);
nand I_21799 (I372684,I372959,I373106);
not I_21800 (I373137,I373067);
nor I_21801 (I373154,I373137,I372877);
DFFARX1 I_21802 (I373154,I2507,I372707,I372696,);
nor I_21803 (I373185,I188002,I188008);
or I_21804 (I372687,I372934,I373185);
nor I_21805 (I372678,I373067,I373185);
or I_21806 (I372681,I372801,I373185);
DFFARX1 I_21807 (I373185,I2507,I372707,I372699,);
not I_21808 (I373285,I2514);
DFFARX1 I_21809 (I38832,I2507,I373285,I373311,);
not I_21810 (I373319,I373311);
nand I_21811 (I373336,I38841,I38850);
and I_21812 (I373353,I373336,I38829);
DFFARX1 I_21813 (I373353,I2507,I373285,I373379,);
not I_21814 (I373387,I38832);
DFFARX1 I_21815 (I38847,I2507,I373285,I373413,);
not I_21816 (I373421,I373413);
nor I_21817 (I373438,I373421,I373319);
and I_21818 (I373455,I373438,I38832);
nor I_21819 (I373472,I373421,I373387);
nor I_21820 (I373268,I373379,I373472);
DFFARX1 I_21821 (I38838,I2507,I373285,I373512,);
nor I_21822 (I373520,I373512,I373379);
not I_21823 (I373537,I373520);
not I_21824 (I373554,I373512);
nor I_21825 (I373571,I373554,I373455);
DFFARX1 I_21826 (I373571,I2507,I373285,I373271,);
nand I_21827 (I373602,I38853,I38829);
and I_21828 (I373619,I373602,I38835);
DFFARX1 I_21829 (I373619,I2507,I373285,I373645,);
nor I_21830 (I373653,I373645,I373512);
DFFARX1 I_21831 (I373653,I2507,I373285,I373253,);
nand I_21832 (I373684,I373645,I373554);
nand I_21833 (I373262,I373537,I373684);
not I_21834 (I373715,I373645);
nor I_21835 (I373732,I373715,I373455);
DFFARX1 I_21836 (I373732,I2507,I373285,I373274,);
nor I_21837 (I373763,I38844,I38829);
or I_21838 (I373265,I373512,I373763);
nor I_21839 (I373256,I373645,I373763);
or I_21840 (I373259,I373379,I373763);
DFFARX1 I_21841 (I373763,I2507,I373285,I373277,);
not I_21842 (I373863,I2514);
DFFARX1 I_21843 (I331637,I2507,I373863,I373889,);
not I_21844 (I373897,I373889);
nand I_21845 (I373914,I331646,I331655);
and I_21846 (I373931,I373914,I331661);
DFFARX1 I_21847 (I373931,I2507,I373863,I373957,);
not I_21848 (I373965,I331658);
DFFARX1 I_21849 (I331643,I2507,I373863,I373991,);
not I_21850 (I373999,I373991);
nor I_21851 (I374016,I373999,I373897);
and I_21852 (I374033,I374016,I331658);
nor I_21853 (I374050,I373999,I373965);
nor I_21854 (I373846,I373957,I374050);
DFFARX1 I_21855 (I331652,I2507,I373863,I374090,);
nor I_21856 (I374098,I374090,I373957);
not I_21857 (I374115,I374098);
not I_21858 (I374132,I374090);
nor I_21859 (I374149,I374132,I374033);
DFFARX1 I_21860 (I374149,I2507,I373863,I373849,);
nand I_21861 (I374180,I331649,I331640);
and I_21862 (I374197,I374180,I331637);
DFFARX1 I_21863 (I374197,I2507,I373863,I374223,);
nor I_21864 (I374231,I374223,I374090);
DFFARX1 I_21865 (I374231,I2507,I373863,I373831,);
nand I_21866 (I374262,I374223,I374132);
nand I_21867 (I373840,I374115,I374262);
not I_21868 (I374293,I374223);
nor I_21869 (I374310,I374293,I374033);
DFFARX1 I_21870 (I374310,I2507,I373863,I373852,);
nor I_21871 (I374341,I331640,I331640);
or I_21872 (I373843,I374090,I374341);
nor I_21873 (I373834,I374223,I374341);
or I_21874 (I373837,I373957,I374341);
DFFARX1 I_21875 (I374341,I2507,I373863,I373855,);
not I_21876 (I374441,I2514);
DFFARX1 I_21877 (I43048,I2507,I374441,I374467,);
not I_21878 (I374475,I374467);
nand I_21879 (I374492,I43057,I43066);
and I_21880 (I374509,I374492,I43045);
DFFARX1 I_21881 (I374509,I2507,I374441,I374535,);
not I_21882 (I374543,I43048);
DFFARX1 I_21883 (I43063,I2507,I374441,I374569,);
not I_21884 (I374577,I374569);
nor I_21885 (I374594,I374577,I374475);
and I_21886 (I374611,I374594,I43048);
nor I_21887 (I374628,I374577,I374543);
nor I_21888 (I374424,I374535,I374628);
DFFARX1 I_21889 (I43054,I2507,I374441,I374668,);
nor I_21890 (I374676,I374668,I374535);
not I_21891 (I374693,I374676);
not I_21892 (I374710,I374668);
nor I_21893 (I374727,I374710,I374611);
DFFARX1 I_21894 (I374727,I2507,I374441,I374427,);
nand I_21895 (I374758,I43069,I43045);
and I_21896 (I374775,I374758,I43051);
DFFARX1 I_21897 (I374775,I2507,I374441,I374801,);
nor I_21898 (I374809,I374801,I374668);
DFFARX1 I_21899 (I374809,I2507,I374441,I374409,);
nand I_21900 (I374840,I374801,I374710);
nand I_21901 (I374418,I374693,I374840);
not I_21902 (I374871,I374801);
nor I_21903 (I374888,I374871,I374611);
DFFARX1 I_21904 (I374888,I2507,I374441,I374430,);
nor I_21905 (I374919,I43060,I43045);
or I_21906 (I374421,I374668,I374919);
nor I_21907 (I374412,I374801,I374919);
or I_21908 (I374415,I374535,I374919);
DFFARX1 I_21909 (I374919,I2507,I374441,I374433,);
not I_21910 (I375019,I2514);
DFFARX1 I_21911 (I171147,I2507,I375019,I375045,);
not I_21912 (I375053,I375045);
nand I_21913 (I375070,I171150,I171126);
and I_21914 (I375087,I375070,I171123);
DFFARX1 I_21915 (I375087,I2507,I375019,I375113,);
not I_21916 (I375121,I171129);
DFFARX1 I_21917 (I171123,I2507,I375019,I375147,);
not I_21918 (I375155,I375147);
nor I_21919 (I375172,I375155,I375053);
and I_21920 (I375189,I375172,I171129);
nor I_21921 (I375206,I375155,I375121);
nor I_21922 (I375002,I375113,I375206);
DFFARX1 I_21923 (I171132,I2507,I375019,I375246,);
nor I_21924 (I375254,I375246,I375113);
not I_21925 (I375271,I375254);
not I_21926 (I375288,I375246);
nor I_21927 (I375305,I375288,I375189);
DFFARX1 I_21928 (I375305,I2507,I375019,I375005,);
nand I_21929 (I375336,I171135,I171144);
and I_21930 (I375353,I375336,I171141);
DFFARX1 I_21931 (I375353,I2507,I375019,I375379,);
nor I_21932 (I375387,I375379,I375246);
DFFARX1 I_21933 (I375387,I2507,I375019,I374987,);
nand I_21934 (I375418,I375379,I375288);
nand I_21935 (I374996,I375271,I375418);
not I_21936 (I375449,I375379);
nor I_21937 (I375466,I375449,I375189);
DFFARX1 I_21938 (I375466,I2507,I375019,I375008,);
nor I_21939 (I375497,I171138,I171144);
or I_21940 (I374999,I375246,I375497);
nor I_21941 (I374990,I375379,I375497);
or I_21942 (I374993,I375113,I375497);
DFFARX1 I_21943 (I375497,I2507,I375019,I375011,);
not I_21944 (I375597,I2514);
DFFARX1 I_21945 (I681531,I2507,I375597,I375623,);
not I_21946 (I375631,I375623);
nand I_21947 (I375648,I681555,I681537);
and I_21948 (I375665,I375648,I681543);
DFFARX1 I_21949 (I375665,I2507,I375597,I375691,);
not I_21950 (I375699,I681549);
DFFARX1 I_21951 (I681534,I2507,I375597,I375725,);
not I_21952 (I375733,I375725);
nor I_21953 (I375750,I375733,I375631);
and I_21954 (I375767,I375750,I681549);
nor I_21955 (I375784,I375733,I375699);
nor I_21956 (I375580,I375691,I375784);
DFFARX1 I_21957 (I681546,I2507,I375597,I375824,);
nor I_21958 (I375832,I375824,I375691);
not I_21959 (I375849,I375832);
not I_21960 (I375866,I375824);
nor I_21961 (I375883,I375866,I375767);
DFFARX1 I_21962 (I375883,I2507,I375597,I375583,);
nand I_21963 (I375914,I681552,I681540);
and I_21964 (I375931,I375914,I681534);
DFFARX1 I_21965 (I375931,I2507,I375597,I375957,);
nor I_21966 (I375965,I375957,I375824);
DFFARX1 I_21967 (I375965,I2507,I375597,I375565,);
nand I_21968 (I375996,I375957,I375866);
nand I_21969 (I375574,I375849,I375996);
not I_21970 (I376027,I375957);
nor I_21971 (I376044,I376027,I375767);
DFFARX1 I_21972 (I376044,I2507,I375597,I375586,);
nor I_21973 (I376075,I681531,I681540);
or I_21974 (I375577,I375824,I376075);
nor I_21975 (I375568,I375957,I376075);
or I_21976 (I375571,I375691,I376075);
DFFARX1 I_21977 (I376075,I2507,I375597,I375589,);
not I_21978 (I376175,I2514);
DFFARX1 I_21979 (I77303,I2507,I376175,I376201,);
not I_21980 (I376209,I376201);
nand I_21981 (I376226,I77312,I77321);
and I_21982 (I376243,I376226,I77300);
DFFARX1 I_21983 (I376243,I2507,I376175,I376269,);
not I_21984 (I376277,I77303);
DFFARX1 I_21985 (I77318,I2507,I376175,I376303,);
not I_21986 (I376311,I376303);
nor I_21987 (I376328,I376311,I376209);
and I_21988 (I376345,I376328,I77303);
nor I_21989 (I376362,I376311,I376277);
nor I_21990 (I376158,I376269,I376362);
DFFARX1 I_21991 (I77309,I2507,I376175,I376402,);
nor I_21992 (I376410,I376402,I376269);
not I_21993 (I376427,I376410);
not I_21994 (I376444,I376402);
nor I_21995 (I376461,I376444,I376345);
DFFARX1 I_21996 (I376461,I2507,I376175,I376161,);
nand I_21997 (I376492,I77324,I77300);
and I_21998 (I376509,I376492,I77306);
DFFARX1 I_21999 (I376509,I2507,I376175,I376535,);
nor I_22000 (I376543,I376535,I376402);
DFFARX1 I_22001 (I376543,I2507,I376175,I376143,);
nand I_22002 (I376574,I376535,I376444);
nand I_22003 (I376152,I376427,I376574);
not I_22004 (I376605,I376535);
nor I_22005 (I376622,I376605,I376345);
DFFARX1 I_22006 (I376622,I2507,I376175,I376164,);
nor I_22007 (I376653,I77315,I77300);
or I_22008 (I376155,I376402,I376653);
nor I_22009 (I376146,I376535,I376653);
or I_22010 (I376149,I376269,I376653);
DFFARX1 I_22011 (I376653,I2507,I376175,I376167,);
not I_22012 (I376753,I2514);
DFFARX1 I_22013 (I563795,I2507,I376753,I376779,);
not I_22014 (I376787,I376779);
nand I_22015 (I376804,I563792,I563810);
and I_22016 (I376821,I376804,I563807);
DFFARX1 I_22017 (I376821,I2507,I376753,I376847,);
not I_22018 (I376855,I563789);
DFFARX1 I_22019 (I563792,I2507,I376753,I376881,);
not I_22020 (I376889,I376881);
nor I_22021 (I376906,I376889,I376787);
and I_22022 (I376923,I376906,I563789);
nor I_22023 (I376940,I376889,I376855);
nor I_22024 (I376736,I376847,I376940);
DFFARX1 I_22025 (I563801,I2507,I376753,I376980,);
nor I_22026 (I376988,I376980,I376847);
not I_22027 (I377005,I376988);
not I_22028 (I377022,I376980);
nor I_22029 (I377039,I377022,I376923);
DFFARX1 I_22030 (I377039,I2507,I376753,I376739,);
nand I_22031 (I377070,I563804,I563789);
and I_22032 (I377087,I377070,I563795);
DFFARX1 I_22033 (I377087,I2507,I376753,I377113,);
nor I_22034 (I377121,I377113,I376980);
DFFARX1 I_22035 (I377121,I2507,I376753,I376721,);
nand I_22036 (I377152,I377113,I377022);
nand I_22037 (I376730,I377005,I377152);
not I_22038 (I377183,I377113);
nor I_22039 (I377200,I377183,I376923);
DFFARX1 I_22040 (I377200,I2507,I376753,I376742,);
nor I_22041 (I377231,I563798,I563789);
or I_22042 (I376733,I376980,I377231);
nor I_22043 (I376724,I377113,I377231);
or I_22044 (I376727,I376847,I377231);
DFFARX1 I_22045 (I377231,I2507,I376753,I376745,);
not I_22046 (I377331,I2514);
DFFARX1 I_22047 (I724585,I2507,I377331,I377357,);
not I_22048 (I377365,I377357);
nand I_22049 (I377382,I724570,I724558);
and I_22050 (I377399,I377382,I724573);
DFFARX1 I_22051 (I377399,I2507,I377331,I377425,);
not I_22052 (I377433,I724558);
DFFARX1 I_22053 (I724576,I2507,I377331,I377459,);
not I_22054 (I377467,I377459);
nor I_22055 (I377484,I377467,I377365);
and I_22056 (I377501,I377484,I724558);
nor I_22057 (I377518,I377467,I377433);
nor I_22058 (I377314,I377425,I377518);
DFFARX1 I_22059 (I724564,I2507,I377331,I377558,);
nor I_22060 (I377566,I377558,I377425);
not I_22061 (I377583,I377566);
not I_22062 (I377600,I377558);
nor I_22063 (I377617,I377600,I377501);
DFFARX1 I_22064 (I377617,I2507,I377331,I377317,);
nand I_22065 (I377648,I724561,I724567);
and I_22066 (I377665,I377648,I724582);
DFFARX1 I_22067 (I377665,I2507,I377331,I377691,);
nor I_22068 (I377699,I377691,I377558);
DFFARX1 I_22069 (I377699,I2507,I377331,I377299,);
nand I_22070 (I377730,I377691,I377600);
nand I_22071 (I377308,I377583,I377730);
not I_22072 (I377761,I377691);
nor I_22073 (I377778,I377761,I377501);
DFFARX1 I_22074 (I377778,I2507,I377331,I377320,);
nor I_22075 (I377809,I724579,I724567);
or I_22076 (I377311,I377558,I377809);
nor I_22077 (I377302,I377691,I377809);
or I_22078 (I377305,I377425,I377809);
DFFARX1 I_22079 (I377809,I2507,I377331,I377323,);
not I_22080 (I377909,I2514);
DFFARX1 I_22081 (I213834,I2507,I377909,I377935,);
not I_22082 (I377943,I377935);
nand I_22083 (I377960,I213837,I213813);
and I_22084 (I377977,I377960,I213810);
DFFARX1 I_22085 (I377977,I2507,I377909,I378003,);
not I_22086 (I378011,I213816);
DFFARX1 I_22087 (I213810,I2507,I377909,I378037,);
not I_22088 (I378045,I378037);
nor I_22089 (I378062,I378045,I377943);
and I_22090 (I378079,I378062,I213816);
nor I_22091 (I378096,I378045,I378011);
nor I_22092 (I377892,I378003,I378096);
DFFARX1 I_22093 (I213819,I2507,I377909,I378136,);
nor I_22094 (I378144,I378136,I378003);
not I_22095 (I378161,I378144);
not I_22096 (I378178,I378136);
nor I_22097 (I378195,I378178,I378079);
DFFARX1 I_22098 (I378195,I2507,I377909,I377895,);
nand I_22099 (I378226,I213822,I213831);
and I_22100 (I378243,I378226,I213828);
DFFARX1 I_22101 (I378243,I2507,I377909,I378269,);
nor I_22102 (I378277,I378269,I378136);
DFFARX1 I_22103 (I378277,I2507,I377909,I377877,);
nand I_22104 (I378308,I378269,I378178);
nand I_22105 (I377886,I378161,I378308);
not I_22106 (I378339,I378269);
nor I_22107 (I378356,I378339,I378079);
DFFARX1 I_22108 (I378356,I2507,I377909,I377898,);
nor I_22109 (I378387,I213825,I213831);
or I_22110 (I377889,I378136,I378387);
nor I_22111 (I377880,I378269,I378387);
or I_22112 (I377883,I378003,I378387);
DFFARX1 I_22113 (I378387,I2507,I377909,I377901,);
not I_22114 (I378487,I2514);
DFFARX1 I_22115 (I663205,I2507,I378487,I378513,);
not I_22116 (I378521,I378513);
nand I_22117 (I378538,I663208,I663217);
and I_22118 (I378555,I378538,I663220);
DFFARX1 I_22119 (I378555,I2507,I378487,I378581,);
not I_22120 (I378589,I663229);
DFFARX1 I_22121 (I663211,I2507,I378487,I378615,);
not I_22122 (I378623,I378615);
nor I_22123 (I378640,I378623,I378521);
and I_22124 (I378657,I378640,I663229);
nor I_22125 (I378674,I378623,I378589);
nor I_22126 (I378470,I378581,I378674);
DFFARX1 I_22127 (I663208,I2507,I378487,I378714,);
nor I_22128 (I378722,I378714,I378581);
not I_22129 (I378739,I378722);
not I_22130 (I378756,I378714);
nor I_22131 (I378773,I378756,I378657);
DFFARX1 I_22132 (I378773,I2507,I378487,I378473,);
nand I_22133 (I378804,I663226,I663205);
and I_22134 (I378821,I378804,I663223);
DFFARX1 I_22135 (I378821,I2507,I378487,I378847,);
nor I_22136 (I378855,I378847,I378714);
DFFARX1 I_22137 (I378855,I2507,I378487,I378455,);
nand I_22138 (I378886,I378847,I378756);
nand I_22139 (I378464,I378739,I378886);
not I_22140 (I378917,I378847);
nor I_22141 (I378934,I378917,I378657);
DFFARX1 I_22142 (I378934,I2507,I378487,I378476,);
nor I_22143 (I378965,I663214,I663205);
or I_22144 (I378467,I378714,I378965);
nor I_22145 (I378458,I378847,I378965);
or I_22146 (I378461,I378581,I378965);
DFFARX1 I_22147 (I378965,I2507,I378487,I378479,);
not I_22148 (I379065,I2514);
DFFARX1 I_22149 (I693050,I2507,I379065,I379091,);
not I_22150 (I379099,I379091);
nand I_22151 (I379116,I693035,I693023);
and I_22152 (I379133,I379116,I693038);
DFFARX1 I_22153 (I379133,I2507,I379065,I379159,);
not I_22154 (I379167,I693023);
DFFARX1 I_22155 (I693041,I2507,I379065,I379193,);
not I_22156 (I379201,I379193);
nor I_22157 (I379218,I379201,I379099);
and I_22158 (I379235,I379218,I693023);
nor I_22159 (I379252,I379201,I379167);
nor I_22160 (I379048,I379159,I379252);
DFFARX1 I_22161 (I693029,I2507,I379065,I379292,);
nor I_22162 (I379300,I379292,I379159);
not I_22163 (I379317,I379300);
not I_22164 (I379334,I379292);
nor I_22165 (I379351,I379334,I379235);
DFFARX1 I_22166 (I379351,I2507,I379065,I379051,);
nand I_22167 (I379382,I693026,I693032);
and I_22168 (I379399,I379382,I693047);
DFFARX1 I_22169 (I379399,I2507,I379065,I379425,);
nor I_22170 (I379433,I379425,I379292);
DFFARX1 I_22171 (I379433,I2507,I379065,I379033,);
nand I_22172 (I379464,I379425,I379334);
nand I_22173 (I379042,I379317,I379464);
not I_22174 (I379495,I379425);
nor I_22175 (I379512,I379495,I379235);
DFFARX1 I_22176 (I379512,I2507,I379065,I379054,);
nor I_22177 (I379543,I693044,I693032);
or I_22178 (I379045,I379292,I379543);
nor I_22179 (I379036,I379425,I379543);
or I_22180 (I379039,I379159,I379543);
DFFARX1 I_22181 (I379543,I2507,I379065,I379057,);
not I_22182 (I379643,I2514);
DFFARX1 I_22183 (I497054,I2507,I379643,I379669,);
not I_22184 (I379677,I379669);
nand I_22185 (I379694,I497030,I497045);
and I_22186 (I379711,I379694,I497057);
DFFARX1 I_22187 (I379711,I2507,I379643,I379737,);
not I_22188 (I379745,I497042);
DFFARX1 I_22189 (I497033,I2507,I379643,I379771,);
not I_22190 (I379779,I379771);
nor I_22191 (I379796,I379779,I379677);
and I_22192 (I379813,I379796,I497042);
nor I_22193 (I379830,I379779,I379745);
nor I_22194 (I379626,I379737,I379830);
DFFARX1 I_22195 (I497030,I2507,I379643,I379870,);
nor I_22196 (I379878,I379870,I379737);
not I_22197 (I379895,I379878);
not I_22198 (I379912,I379870);
nor I_22199 (I379929,I379912,I379813);
DFFARX1 I_22200 (I379929,I2507,I379643,I379629,);
nand I_22201 (I379960,I497048,I497039);
and I_22202 (I379977,I379960,I497051);
DFFARX1 I_22203 (I379977,I2507,I379643,I380003,);
nor I_22204 (I380011,I380003,I379870);
DFFARX1 I_22205 (I380011,I2507,I379643,I379611,);
nand I_22206 (I380042,I380003,I379912);
nand I_22207 (I379620,I379895,I380042);
not I_22208 (I380073,I380003);
nor I_22209 (I380090,I380073,I379813);
DFFARX1 I_22210 (I380090,I2507,I379643,I379632,);
nor I_22211 (I380121,I497036,I497039);
or I_22212 (I379623,I379870,I380121);
nor I_22213 (I379614,I380003,I380121);
or I_22214 (I379617,I379737,I380121);
DFFARX1 I_22215 (I380121,I2507,I379643,I379635,);
not I_22216 (I380221,I2514);
DFFARX1 I_22217 (I572851,I2507,I380221,I380247,);
not I_22218 (I380255,I380247);
nand I_22219 (I380272,I572833,I572845);
and I_22220 (I380289,I380272,I572848);
DFFARX1 I_22221 (I380289,I2507,I380221,I380315,);
not I_22222 (I380323,I572842);
DFFARX1 I_22223 (I572839,I2507,I380221,I380349,);
not I_22224 (I380357,I380349);
nor I_22225 (I380374,I380357,I380255);
and I_22226 (I380391,I380374,I572842);
nor I_22227 (I380408,I380357,I380323);
nor I_22228 (I380204,I380315,I380408);
DFFARX1 I_22229 (I572857,I2507,I380221,I380448,);
nor I_22230 (I380456,I380448,I380315);
not I_22231 (I380473,I380456);
not I_22232 (I380490,I380448);
nor I_22233 (I380507,I380490,I380391);
DFFARX1 I_22234 (I380507,I2507,I380221,I380207,);
nand I_22235 (I380538,I572836,I572836);
and I_22236 (I380555,I380538,I572833);
DFFARX1 I_22237 (I380555,I2507,I380221,I380581,);
nor I_22238 (I380589,I380581,I380448);
DFFARX1 I_22239 (I380589,I2507,I380221,I380189,);
nand I_22240 (I380620,I380581,I380490);
nand I_22241 (I380198,I380473,I380620);
not I_22242 (I380651,I380581);
nor I_22243 (I380668,I380651,I380391);
DFFARX1 I_22244 (I380668,I2507,I380221,I380210,);
nor I_22245 (I380699,I572854,I572836);
or I_22246 (I380201,I380448,I380699);
nor I_22247 (I380192,I380581,I380699);
or I_22248 (I380195,I380315,I380699);
DFFARX1 I_22249 (I380699,I2507,I380221,I380213,);
not I_22250 (I380799,I2514);
DFFARX1 I_22251 (I254721,I2507,I380799,I380825,);
not I_22252 (I380833,I380825);
nand I_22253 (I380850,I254712,I254730);
and I_22254 (I380867,I380850,I254733);
DFFARX1 I_22255 (I380867,I2507,I380799,I380893,);
not I_22256 (I380901,I254727);
DFFARX1 I_22257 (I254715,I2507,I380799,I380927,);
not I_22258 (I380935,I380927);
nor I_22259 (I380952,I380935,I380833);
and I_22260 (I380969,I380952,I254727);
nor I_22261 (I380986,I380935,I380901);
nor I_22262 (I380782,I380893,I380986);
DFFARX1 I_22263 (I254724,I2507,I380799,I381026,);
nor I_22264 (I381034,I381026,I380893);
not I_22265 (I381051,I381034);
not I_22266 (I381068,I381026);
nor I_22267 (I381085,I381068,I380969);
DFFARX1 I_22268 (I381085,I2507,I380799,I380785,);
nand I_22269 (I381116,I254739,I254736);
and I_22270 (I381133,I381116,I254718);
DFFARX1 I_22271 (I381133,I2507,I380799,I381159,);
nor I_22272 (I381167,I381159,I381026);
DFFARX1 I_22273 (I381167,I2507,I380799,I380767,);
nand I_22274 (I381198,I381159,I381068);
nand I_22275 (I380776,I381051,I381198);
not I_22276 (I381229,I381159);
nor I_22277 (I381246,I381229,I380969);
DFFARX1 I_22278 (I381246,I2507,I380799,I380788,);
nor I_22279 (I381277,I254712,I254736);
or I_22280 (I380779,I381026,I381277);
nor I_22281 (I380770,I381159,I381277);
or I_22282 (I380773,I380893,I381277);
DFFARX1 I_22283 (I381277,I2507,I380799,I380791,);
not I_22284 (I381377,I2514);
DFFARX1 I_22285 (I149074,I2507,I381377,I381403,);
not I_22286 (I381411,I381403);
nand I_22287 (I381428,I149077,I149098);
and I_22288 (I381445,I381428,I149086);
DFFARX1 I_22289 (I381445,I2507,I381377,I381471,);
not I_22290 (I381479,I149083);
DFFARX1 I_22291 (I149074,I2507,I381377,I381505,);
not I_22292 (I381513,I381505);
nor I_22293 (I381530,I381513,I381411);
and I_22294 (I381547,I381530,I149083);
nor I_22295 (I381564,I381513,I381479);
nor I_22296 (I381360,I381471,I381564);
DFFARX1 I_22297 (I149092,I2507,I381377,I381604,);
nor I_22298 (I381612,I381604,I381471);
not I_22299 (I381629,I381612);
not I_22300 (I381646,I381604);
nor I_22301 (I381663,I381646,I381547);
DFFARX1 I_22302 (I381663,I2507,I381377,I381363,);
nand I_22303 (I381694,I149077,I149080);
and I_22304 (I381711,I381694,I149089);
DFFARX1 I_22305 (I381711,I2507,I381377,I381737,);
nor I_22306 (I381745,I381737,I381604);
DFFARX1 I_22307 (I381745,I2507,I381377,I381345,);
nand I_22308 (I381776,I381737,I381646);
nand I_22309 (I381354,I381629,I381776);
not I_22310 (I381807,I381737);
nor I_22311 (I381824,I381807,I381547);
DFFARX1 I_22312 (I381824,I2507,I381377,I381366,);
nor I_22313 (I381855,I149095,I149080);
or I_22314 (I381357,I381604,I381855);
nor I_22315 (I381348,I381737,I381855);
or I_22316 (I381351,I381471,I381855);
DFFARX1 I_22317 (I381855,I2507,I381377,I381369,);
not I_22318 (I381955,I2514);
DFFARX1 I_22319 (I261793,I2507,I381955,I381981,);
not I_22320 (I381989,I381981);
nand I_22321 (I382006,I261784,I261802);
and I_22322 (I382023,I382006,I261805);
DFFARX1 I_22323 (I382023,I2507,I381955,I382049,);
not I_22324 (I382057,I261799);
DFFARX1 I_22325 (I261787,I2507,I381955,I382083,);
not I_22326 (I382091,I382083);
nor I_22327 (I382108,I382091,I381989);
and I_22328 (I382125,I382108,I261799);
nor I_22329 (I382142,I382091,I382057);
nor I_22330 (I381938,I382049,I382142);
DFFARX1 I_22331 (I261796,I2507,I381955,I382182,);
nor I_22332 (I382190,I382182,I382049);
not I_22333 (I382207,I382190);
not I_22334 (I382224,I382182);
nor I_22335 (I382241,I382224,I382125);
DFFARX1 I_22336 (I382241,I2507,I381955,I381941,);
nand I_22337 (I382272,I261811,I261808);
and I_22338 (I382289,I382272,I261790);
DFFARX1 I_22339 (I382289,I2507,I381955,I382315,);
nor I_22340 (I382323,I382315,I382182);
DFFARX1 I_22341 (I382323,I2507,I381955,I381923,);
nand I_22342 (I382354,I382315,I382224);
nand I_22343 (I381932,I382207,I382354);
not I_22344 (I382385,I382315);
nor I_22345 (I382402,I382385,I382125);
DFFARX1 I_22346 (I382402,I2507,I381955,I381944,);
nor I_22347 (I382433,I261784,I261808);
or I_22348 (I381935,I382182,I382433);
nor I_22349 (I381926,I382315,I382433);
or I_22350 (I381929,I382049,I382433);
DFFARX1 I_22351 (I382433,I2507,I381955,I381947,);
not I_22352 (I382533,I2514);
DFFARX1 I_22353 (I337995,I2507,I382533,I382559,);
not I_22354 (I382567,I382559);
nand I_22355 (I382584,I338004,I338013);
and I_22356 (I382601,I382584,I338019);
DFFARX1 I_22357 (I382601,I2507,I382533,I382627,);
not I_22358 (I382635,I338016);
DFFARX1 I_22359 (I338001,I2507,I382533,I382661,);
not I_22360 (I382669,I382661);
nor I_22361 (I382686,I382669,I382567);
and I_22362 (I382703,I382686,I338016);
nor I_22363 (I382720,I382669,I382635);
nor I_22364 (I382516,I382627,I382720);
DFFARX1 I_22365 (I338010,I2507,I382533,I382760,);
nor I_22366 (I382768,I382760,I382627);
not I_22367 (I382785,I382768);
not I_22368 (I382802,I382760);
nor I_22369 (I382819,I382802,I382703);
DFFARX1 I_22370 (I382819,I2507,I382533,I382519,);
nand I_22371 (I382850,I338007,I337998);
and I_22372 (I382867,I382850,I337995);
DFFARX1 I_22373 (I382867,I2507,I382533,I382893,);
nor I_22374 (I382901,I382893,I382760);
DFFARX1 I_22375 (I382901,I2507,I382533,I382501,);
nand I_22376 (I382932,I382893,I382802);
nand I_22377 (I382510,I382785,I382932);
not I_22378 (I382963,I382893);
nor I_22379 (I382980,I382963,I382703);
DFFARX1 I_22380 (I382980,I2507,I382533,I382522,);
nor I_22381 (I383011,I337998,I337998);
or I_22382 (I382513,I382760,I383011);
nor I_22383 (I382504,I382893,I383011);
or I_22384 (I382507,I382627,I383011);
DFFARX1 I_22385 (I383011,I2507,I382533,I382525,);
not I_22386 (I383111,I2514);
DFFARX1 I_22387 (I559307,I2507,I383111,I383137,);
not I_22388 (I383145,I383137);
nand I_22389 (I383162,I559304,I559322);
and I_22390 (I383179,I383162,I559319);
DFFARX1 I_22391 (I383179,I2507,I383111,I383205,);
not I_22392 (I383213,I559301);
DFFARX1 I_22393 (I559304,I2507,I383111,I383239,);
not I_22394 (I383247,I383239);
nor I_22395 (I383264,I383247,I383145);
and I_22396 (I383281,I383264,I559301);
nor I_22397 (I383298,I383247,I383213);
nor I_22398 (I383094,I383205,I383298);
DFFARX1 I_22399 (I559313,I2507,I383111,I383338,);
nor I_22400 (I383346,I383338,I383205);
not I_22401 (I383363,I383346);
not I_22402 (I383380,I383338);
nor I_22403 (I383397,I383380,I383281);
DFFARX1 I_22404 (I383397,I2507,I383111,I383097,);
nand I_22405 (I383428,I559316,I559301);
and I_22406 (I383445,I383428,I559307);
DFFARX1 I_22407 (I383445,I2507,I383111,I383471,);
nor I_22408 (I383479,I383471,I383338);
DFFARX1 I_22409 (I383479,I2507,I383111,I383079,);
nand I_22410 (I383510,I383471,I383380);
nand I_22411 (I383088,I383363,I383510);
not I_22412 (I383541,I383471);
nor I_22413 (I383558,I383541,I383281);
DFFARX1 I_22414 (I383558,I2507,I383111,I383100,);
nor I_22415 (I383589,I559310,I559301);
or I_22416 (I383091,I383338,I383589);
nor I_22417 (I383082,I383471,I383589);
or I_22418 (I383085,I383205,I383589);
DFFARX1 I_22419 (I383589,I2507,I383111,I383103,);
not I_22420 (I383689,I2514);
DFFARX1 I_22421 (I255265,I2507,I383689,I383715,);
not I_22422 (I383723,I383715);
nand I_22423 (I383740,I255256,I255274);
and I_22424 (I383757,I383740,I255277);
DFFARX1 I_22425 (I383757,I2507,I383689,I383783,);
not I_22426 (I383791,I255271);
DFFARX1 I_22427 (I255259,I2507,I383689,I383817,);
not I_22428 (I383825,I383817);
nor I_22429 (I383842,I383825,I383723);
and I_22430 (I383859,I383842,I255271);
nor I_22431 (I383876,I383825,I383791);
nor I_22432 (I383672,I383783,I383876);
DFFARX1 I_22433 (I255268,I2507,I383689,I383916,);
nor I_22434 (I383924,I383916,I383783);
not I_22435 (I383941,I383924);
not I_22436 (I383958,I383916);
nor I_22437 (I383975,I383958,I383859);
DFFARX1 I_22438 (I383975,I2507,I383689,I383675,);
nand I_22439 (I384006,I255283,I255280);
and I_22440 (I384023,I384006,I255262);
DFFARX1 I_22441 (I384023,I2507,I383689,I384049,);
nor I_22442 (I384057,I384049,I383916);
DFFARX1 I_22443 (I384057,I2507,I383689,I383657,);
nand I_22444 (I384088,I384049,I383958);
nand I_22445 (I383666,I383941,I384088);
not I_22446 (I384119,I384049);
nor I_22447 (I384136,I384119,I383859);
DFFARX1 I_22448 (I384136,I2507,I383689,I383678,);
nor I_22449 (I384167,I255256,I255280);
or I_22450 (I383669,I383916,I384167);
nor I_22451 (I383660,I384049,I384167);
or I_22452 (I383663,I383783,I384167);
DFFARX1 I_22453 (I384167,I2507,I383689,I383681,);
not I_22454 (I384267,I2514);
DFFARX1 I_22455 (I181687,I2507,I384267,I384293,);
not I_22456 (I384301,I384293);
nand I_22457 (I384318,I181690,I181666);
and I_22458 (I384335,I384318,I181663);
DFFARX1 I_22459 (I384335,I2507,I384267,I384361,);
not I_22460 (I384369,I181669);
DFFARX1 I_22461 (I181663,I2507,I384267,I384395,);
not I_22462 (I384403,I384395);
nor I_22463 (I384420,I384403,I384301);
and I_22464 (I384437,I384420,I181669);
nor I_22465 (I384454,I384403,I384369);
nor I_22466 (I384250,I384361,I384454);
DFFARX1 I_22467 (I181672,I2507,I384267,I384494,);
nor I_22468 (I384502,I384494,I384361);
not I_22469 (I384519,I384502);
not I_22470 (I384536,I384494);
nor I_22471 (I384553,I384536,I384437);
DFFARX1 I_22472 (I384553,I2507,I384267,I384253,);
nand I_22473 (I384584,I181675,I181684);
and I_22474 (I384601,I384584,I181681);
DFFARX1 I_22475 (I384601,I2507,I384267,I384627,);
nor I_22476 (I384635,I384627,I384494);
DFFARX1 I_22477 (I384635,I2507,I384267,I384235,);
nand I_22478 (I384666,I384627,I384536);
nand I_22479 (I384244,I384519,I384666);
not I_22480 (I384697,I384627);
nor I_22481 (I384714,I384697,I384437);
DFFARX1 I_22482 (I384714,I2507,I384267,I384256,);
nor I_22483 (I384745,I181678,I181684);
or I_22484 (I384247,I384494,I384745);
nor I_22485 (I384238,I384627,I384745);
or I_22486 (I384241,I384361,I384745);
DFFARX1 I_22487 (I384745,I2507,I384267,I384259,);
not I_22488 (I384845,I2514);
DFFARX1 I_22489 (I706140,I2507,I384845,I384871,);
not I_22490 (I384879,I384871);
nand I_22491 (I384896,I706125,I706113);
and I_22492 (I384913,I384896,I706128);
DFFARX1 I_22493 (I384913,I2507,I384845,I384939,);
not I_22494 (I384947,I706113);
DFFARX1 I_22495 (I706131,I2507,I384845,I384973,);
not I_22496 (I384981,I384973);
nor I_22497 (I384998,I384981,I384879);
and I_22498 (I385015,I384998,I706113);
nor I_22499 (I385032,I384981,I384947);
nor I_22500 (I384828,I384939,I385032);
DFFARX1 I_22501 (I706119,I2507,I384845,I385072,);
nor I_22502 (I385080,I385072,I384939);
not I_22503 (I385097,I385080);
not I_22504 (I385114,I385072);
nor I_22505 (I385131,I385114,I385015);
DFFARX1 I_22506 (I385131,I2507,I384845,I384831,);
nand I_22507 (I385162,I706116,I706122);
and I_22508 (I385179,I385162,I706137);
DFFARX1 I_22509 (I385179,I2507,I384845,I385205,);
nor I_22510 (I385213,I385205,I385072);
DFFARX1 I_22511 (I385213,I2507,I384845,I384813,);
nand I_22512 (I385244,I385205,I385114);
nand I_22513 (I384822,I385097,I385244);
not I_22514 (I385275,I385205);
nor I_22515 (I385292,I385275,I385015);
DFFARX1 I_22516 (I385292,I2507,I384845,I384834,);
nor I_22517 (I385323,I706134,I706122);
or I_22518 (I384825,I385072,I385323);
nor I_22519 (I384816,I385205,I385323);
or I_22520 (I384819,I384939,I385323);
DFFARX1 I_22521 (I385323,I2507,I384845,I384837,);
not I_22522 (I385423,I2514);
DFFARX1 I_22523 (I454477,I2507,I385423,I385449,);
not I_22524 (I385457,I385449);
nand I_22525 (I385474,I454465,I454483);
and I_22526 (I385491,I385474,I454480);
DFFARX1 I_22527 (I385491,I2507,I385423,I385517,);
not I_22528 (I385525,I454471);
DFFARX1 I_22529 (I454468,I2507,I385423,I385551,);
not I_22530 (I385559,I385551);
nor I_22531 (I385576,I385559,I385457);
and I_22532 (I385593,I385576,I454471);
nor I_22533 (I385610,I385559,I385525);
nor I_22534 (I385406,I385517,I385610);
DFFARX1 I_22535 (I454462,I2507,I385423,I385650,);
nor I_22536 (I385658,I385650,I385517);
not I_22537 (I385675,I385658);
not I_22538 (I385692,I385650);
nor I_22539 (I385709,I385692,I385593);
DFFARX1 I_22540 (I385709,I2507,I385423,I385409,);
nand I_22541 (I385740,I454462,I454465);
and I_22542 (I385757,I385740,I454468);
DFFARX1 I_22543 (I385757,I2507,I385423,I385783,);
nor I_22544 (I385791,I385783,I385650);
DFFARX1 I_22545 (I385791,I2507,I385423,I385391,);
nand I_22546 (I385822,I385783,I385692);
nand I_22547 (I385400,I385675,I385822);
not I_22548 (I385853,I385783);
nor I_22549 (I385870,I385853,I385593);
DFFARX1 I_22550 (I385870,I2507,I385423,I385412,);
nor I_22551 (I385901,I454474,I454465);
or I_22552 (I385403,I385650,I385901);
nor I_22553 (I385394,I385783,I385901);
or I_22554 (I385397,I385517,I385901);
DFFARX1 I_22555 (I385901,I2507,I385423,I385415,);
not I_22556 (I386001,I2514);
DFFARX1 I_22557 (I274305,I2507,I386001,I386027,);
not I_22558 (I386035,I386027);
nand I_22559 (I386052,I274296,I274314);
and I_22560 (I386069,I386052,I274317);
DFFARX1 I_22561 (I386069,I2507,I386001,I386095,);
not I_22562 (I386103,I274311);
DFFARX1 I_22563 (I274299,I2507,I386001,I386129,);
not I_22564 (I386137,I386129);
nor I_22565 (I386154,I386137,I386035);
and I_22566 (I386171,I386154,I274311);
nor I_22567 (I386188,I386137,I386103);
nor I_22568 (I385984,I386095,I386188);
DFFARX1 I_22569 (I274308,I2507,I386001,I386228,);
nor I_22570 (I386236,I386228,I386095);
not I_22571 (I386253,I386236);
not I_22572 (I386270,I386228);
nor I_22573 (I386287,I386270,I386171);
DFFARX1 I_22574 (I386287,I2507,I386001,I385987,);
nand I_22575 (I386318,I274323,I274320);
and I_22576 (I386335,I386318,I274302);
DFFARX1 I_22577 (I386335,I2507,I386001,I386361,);
nor I_22578 (I386369,I386361,I386228);
DFFARX1 I_22579 (I386369,I2507,I386001,I385969,);
nand I_22580 (I386400,I386361,I386270);
nand I_22581 (I385978,I386253,I386400);
not I_22582 (I386431,I386361);
nor I_22583 (I386448,I386431,I386171);
DFFARX1 I_22584 (I386448,I2507,I386001,I385990,);
nor I_22585 (I386479,I274296,I274320);
or I_22586 (I385981,I386228,I386479);
nor I_22587 (I385972,I386361,I386479);
or I_22588 (I385975,I386095,I386479);
DFFARX1 I_22589 (I386479,I2507,I386001,I385993,);
not I_22590 (I386579,I2514);
DFFARX1 I_22591 (I530000,I2507,I386579,I386605,);
not I_22592 (I386613,I386605);
nand I_22593 (I386630,I529976,I529991);
and I_22594 (I386647,I386630,I530003);
DFFARX1 I_22595 (I386647,I2507,I386579,I386673,);
not I_22596 (I386681,I529988);
DFFARX1 I_22597 (I529979,I2507,I386579,I386707,);
not I_22598 (I386715,I386707);
nor I_22599 (I386732,I386715,I386613);
and I_22600 (I386749,I386732,I529988);
nor I_22601 (I386766,I386715,I386681);
nor I_22602 (I386562,I386673,I386766);
DFFARX1 I_22603 (I529976,I2507,I386579,I386806,);
nor I_22604 (I386814,I386806,I386673);
not I_22605 (I386831,I386814);
not I_22606 (I386848,I386806);
nor I_22607 (I386865,I386848,I386749);
DFFARX1 I_22608 (I386865,I2507,I386579,I386565,);
nand I_22609 (I386896,I529994,I529985);
and I_22610 (I386913,I386896,I529997);
DFFARX1 I_22611 (I386913,I2507,I386579,I386939,);
nor I_22612 (I386947,I386939,I386806);
DFFARX1 I_22613 (I386947,I2507,I386579,I386547,);
nand I_22614 (I386978,I386939,I386848);
nand I_22615 (I386556,I386831,I386978);
not I_22616 (I387009,I386939);
nor I_22617 (I387026,I387009,I386749);
DFFARX1 I_22618 (I387026,I2507,I386579,I386568,);
nor I_22619 (I387057,I529982,I529985);
or I_22620 (I386559,I386806,I387057);
nor I_22621 (I386550,I386939,I387057);
or I_22622 (I386553,I386673,I387057);
DFFARX1 I_22623 (I387057,I2507,I386579,I386571,);
not I_22624 (I387157,I2514);
DFFARX1 I_22625 (I251457,I2507,I387157,I387183,);
not I_22626 (I387191,I387183);
nand I_22627 (I387208,I251448,I251466);
and I_22628 (I387225,I387208,I251469);
DFFARX1 I_22629 (I387225,I2507,I387157,I387251,);
not I_22630 (I387259,I251463);
DFFARX1 I_22631 (I251451,I2507,I387157,I387285,);
not I_22632 (I387293,I387285);
nor I_22633 (I387310,I387293,I387191);
and I_22634 (I387327,I387310,I251463);
nor I_22635 (I387344,I387293,I387259);
nor I_22636 (I387140,I387251,I387344);
DFFARX1 I_22637 (I251460,I2507,I387157,I387384,);
nor I_22638 (I387392,I387384,I387251);
not I_22639 (I387409,I387392);
not I_22640 (I387426,I387384);
nor I_22641 (I387443,I387426,I387327);
DFFARX1 I_22642 (I387443,I2507,I387157,I387143,);
nand I_22643 (I387474,I251475,I251472);
and I_22644 (I387491,I387474,I251454);
DFFARX1 I_22645 (I387491,I2507,I387157,I387517,);
nor I_22646 (I387525,I387517,I387384);
DFFARX1 I_22647 (I387525,I2507,I387157,I387125,);
nand I_22648 (I387556,I387517,I387426);
nand I_22649 (I387134,I387409,I387556);
not I_22650 (I387587,I387517);
nor I_22651 (I387604,I387587,I387327);
DFFARX1 I_22652 (I387604,I2507,I387157,I387146,);
nor I_22653 (I387635,I251448,I251472);
or I_22654 (I387137,I387384,I387635);
nor I_22655 (I387128,I387517,I387635);
or I_22656 (I387131,I387251,I387635);
DFFARX1 I_22657 (I387635,I2507,I387157,I387149,);
not I_22658 (I387735,I2514);
DFFARX1 I_22659 (I250369,I2507,I387735,I387761,);
not I_22660 (I387769,I387761);
nand I_22661 (I387786,I250360,I250378);
and I_22662 (I387803,I387786,I250381);
DFFARX1 I_22663 (I387803,I2507,I387735,I387829,);
not I_22664 (I387837,I250375);
DFFARX1 I_22665 (I250363,I2507,I387735,I387863,);
not I_22666 (I387871,I387863);
nor I_22667 (I387888,I387871,I387769);
and I_22668 (I387905,I387888,I250375);
nor I_22669 (I387922,I387871,I387837);
nor I_22670 (I387718,I387829,I387922);
DFFARX1 I_22671 (I250372,I2507,I387735,I387962,);
nor I_22672 (I387970,I387962,I387829);
not I_22673 (I387987,I387970);
not I_22674 (I388004,I387962);
nor I_22675 (I388021,I388004,I387905);
DFFARX1 I_22676 (I388021,I2507,I387735,I387721,);
nand I_22677 (I388052,I250387,I250384);
and I_22678 (I388069,I388052,I250366);
DFFARX1 I_22679 (I388069,I2507,I387735,I388095,);
nor I_22680 (I388103,I388095,I387962);
DFFARX1 I_22681 (I388103,I2507,I387735,I387703,);
nand I_22682 (I388134,I388095,I388004);
nand I_22683 (I387712,I387987,I388134);
not I_22684 (I388165,I388095);
nor I_22685 (I388182,I388165,I387905);
DFFARX1 I_22686 (I388182,I2507,I387735,I387724,);
nor I_22687 (I388213,I250360,I250384);
or I_22688 (I387715,I387962,I388213);
nor I_22689 (I387706,I388095,I388213);
or I_22690 (I387709,I387829,I388213);
DFFARX1 I_22691 (I388213,I2507,I387735,I387727,);
not I_22692 (I388313,I2514);
DFFARX1 I_22693 (I638725,I2507,I388313,I388339,);
not I_22694 (I388347,I388339);
nand I_22695 (I388364,I638728,I638737);
and I_22696 (I388381,I388364,I638740);
DFFARX1 I_22697 (I388381,I2507,I388313,I388407,);
not I_22698 (I388415,I638749);
DFFARX1 I_22699 (I638731,I2507,I388313,I388441,);
not I_22700 (I388449,I388441);
nor I_22701 (I388466,I388449,I388347);
and I_22702 (I388483,I388466,I638749);
nor I_22703 (I388500,I388449,I388415);
nor I_22704 (I388296,I388407,I388500);
DFFARX1 I_22705 (I638728,I2507,I388313,I388540,);
nor I_22706 (I388548,I388540,I388407);
not I_22707 (I388565,I388548);
not I_22708 (I388582,I388540);
nor I_22709 (I388599,I388582,I388483);
DFFARX1 I_22710 (I388599,I2507,I388313,I388299,);
nand I_22711 (I388630,I638746,I638725);
and I_22712 (I388647,I388630,I638743);
DFFARX1 I_22713 (I388647,I2507,I388313,I388673,);
nor I_22714 (I388681,I388673,I388540);
DFFARX1 I_22715 (I388681,I2507,I388313,I388281,);
nand I_22716 (I388712,I388673,I388582);
nand I_22717 (I388290,I388565,I388712);
not I_22718 (I388743,I388673);
nor I_22719 (I388760,I388743,I388483);
DFFARX1 I_22720 (I388760,I2507,I388313,I388302,);
nor I_22721 (I388791,I638734,I638725);
or I_22722 (I388293,I388540,I388791);
nor I_22723 (I388284,I388673,I388791);
or I_22724 (I388287,I388407,I388791);
DFFARX1 I_22725 (I388791,I2507,I388313,I388305,);
not I_22726 (I388891,I2514);
DFFARX1 I_22727 (I289103,I2507,I388891,I388917,);
not I_22728 (I388925,I388917);
nand I_22729 (I388942,I289118,I289103);
and I_22730 (I388959,I388942,I289106);
DFFARX1 I_22731 (I388959,I2507,I388891,I388985,);
not I_22732 (I388993,I289106);
DFFARX1 I_22733 (I289115,I2507,I388891,I389019,);
not I_22734 (I389027,I389019);
nor I_22735 (I389044,I389027,I388925);
and I_22736 (I389061,I389044,I289106);
nor I_22737 (I389078,I389027,I388993);
nor I_22738 (I388874,I388985,I389078);
DFFARX1 I_22739 (I289109,I2507,I388891,I389118,);
nor I_22740 (I389126,I389118,I388985);
not I_22741 (I389143,I389126);
not I_22742 (I389160,I389118);
nor I_22743 (I389177,I389160,I389061);
DFFARX1 I_22744 (I389177,I2507,I388891,I388877,);
nand I_22745 (I389208,I289112,I289121);
and I_22746 (I389225,I389208,I289127);
DFFARX1 I_22747 (I389225,I2507,I388891,I389251,);
nor I_22748 (I389259,I389251,I389118);
DFFARX1 I_22749 (I389259,I2507,I388891,I388859,);
nand I_22750 (I389290,I389251,I389160);
nand I_22751 (I388868,I389143,I389290);
not I_22752 (I389321,I389251);
nor I_22753 (I389338,I389321,I389061);
DFFARX1 I_22754 (I389338,I2507,I388891,I388880,);
nor I_22755 (I389369,I289124,I289121);
or I_22756 (I388871,I389118,I389369);
nor I_22757 (I388862,I389251,I389369);
or I_22758 (I388865,I388985,I389369);
DFFARX1 I_22759 (I389369,I2507,I388891,I388883,);
not I_22760 (I389469,I2514);
DFFARX1 I_22761 (I489948,I2507,I389469,I389495,);
not I_22762 (I389503,I389495);
nand I_22763 (I389520,I489924,I489939);
and I_22764 (I389537,I389520,I489951);
DFFARX1 I_22765 (I389537,I2507,I389469,I389563,);
not I_22766 (I389571,I489936);
DFFARX1 I_22767 (I489927,I2507,I389469,I389597,);
not I_22768 (I389605,I389597);
nor I_22769 (I389622,I389605,I389503);
and I_22770 (I389639,I389622,I489936);
nor I_22771 (I389656,I389605,I389571);
nor I_22772 (I389452,I389563,I389656);
DFFARX1 I_22773 (I489924,I2507,I389469,I389696,);
nor I_22774 (I389704,I389696,I389563);
not I_22775 (I389721,I389704);
not I_22776 (I389738,I389696);
nor I_22777 (I389755,I389738,I389639);
DFFARX1 I_22778 (I389755,I2507,I389469,I389455,);
nand I_22779 (I389786,I489942,I489933);
and I_22780 (I389803,I389786,I489945);
DFFARX1 I_22781 (I389803,I2507,I389469,I389829,);
nor I_22782 (I389837,I389829,I389696);
DFFARX1 I_22783 (I389837,I2507,I389469,I389437,);
nand I_22784 (I389868,I389829,I389738);
nand I_22785 (I389446,I389721,I389868);
not I_22786 (I389899,I389829);
nor I_22787 (I389916,I389899,I389639);
DFFARX1 I_22788 (I389916,I2507,I389469,I389458,);
nor I_22789 (I389947,I489930,I489933);
or I_22790 (I389449,I389696,I389947);
nor I_22791 (I389440,I389829,I389947);
or I_22792 (I389443,I389563,I389947);
DFFARX1 I_22793 (I389947,I2507,I389469,I389461,);
not I_22794 (I390047,I2514);
DFFARX1 I_22795 (I270497,I2507,I390047,I390073,);
not I_22796 (I390081,I390073);
nand I_22797 (I390098,I270488,I270506);
and I_22798 (I390115,I390098,I270509);
DFFARX1 I_22799 (I390115,I2507,I390047,I390141,);
not I_22800 (I390149,I270503);
DFFARX1 I_22801 (I270491,I2507,I390047,I390175,);
not I_22802 (I390183,I390175);
nor I_22803 (I390200,I390183,I390081);
and I_22804 (I390217,I390200,I270503);
nor I_22805 (I390234,I390183,I390149);
nor I_22806 (I390030,I390141,I390234);
DFFARX1 I_22807 (I270500,I2507,I390047,I390274,);
nor I_22808 (I390282,I390274,I390141);
not I_22809 (I390299,I390282);
not I_22810 (I390316,I390274);
nor I_22811 (I390333,I390316,I390217);
DFFARX1 I_22812 (I390333,I2507,I390047,I390033,);
nand I_22813 (I390364,I270515,I270512);
and I_22814 (I390381,I390364,I270494);
DFFARX1 I_22815 (I390381,I2507,I390047,I390407,);
nor I_22816 (I390415,I390407,I390274);
DFFARX1 I_22817 (I390415,I2507,I390047,I390015,);
nand I_22818 (I390446,I390407,I390316);
nand I_22819 (I390024,I390299,I390446);
not I_22820 (I390477,I390407);
nor I_22821 (I390494,I390477,I390217);
DFFARX1 I_22822 (I390494,I2507,I390047,I390036,);
nor I_22823 (I390525,I270488,I270512);
or I_22824 (I390027,I390274,I390525);
nor I_22825 (I390018,I390407,I390525);
or I_22826 (I390021,I390141,I390525);
DFFARX1 I_22827 (I390525,I2507,I390047,I390039,);
not I_22828 (I390625,I2514);
DFFARX1 I_22829 (I552014,I2507,I390625,I390651,);
not I_22830 (I390659,I390651);
nand I_22831 (I390676,I552011,I552029);
and I_22832 (I390693,I390676,I552026);
DFFARX1 I_22833 (I390693,I2507,I390625,I390719,);
not I_22834 (I390727,I552008);
DFFARX1 I_22835 (I552011,I2507,I390625,I390753,);
not I_22836 (I390761,I390753);
nor I_22837 (I390778,I390761,I390659);
and I_22838 (I390795,I390778,I552008);
nor I_22839 (I390812,I390761,I390727);
nor I_22840 (I390608,I390719,I390812);
DFFARX1 I_22841 (I552020,I2507,I390625,I390852,);
nor I_22842 (I390860,I390852,I390719);
not I_22843 (I390877,I390860);
not I_22844 (I390894,I390852);
nor I_22845 (I390911,I390894,I390795);
DFFARX1 I_22846 (I390911,I2507,I390625,I390611,);
nand I_22847 (I390942,I552023,I552008);
and I_22848 (I390959,I390942,I552014);
DFFARX1 I_22849 (I390959,I2507,I390625,I390985,);
nor I_22850 (I390993,I390985,I390852);
DFFARX1 I_22851 (I390993,I2507,I390625,I390593,);
nand I_22852 (I391024,I390985,I390894);
nand I_22853 (I390602,I390877,I391024);
not I_22854 (I391055,I390985);
nor I_22855 (I391072,I391055,I390795);
DFFARX1 I_22856 (I391072,I2507,I390625,I390614,);
nor I_22857 (I391103,I552017,I552008);
or I_22858 (I390605,I390852,I391103);
nor I_22859 (I390596,I390985,I391103);
or I_22860 (I390599,I390719,I391103);
DFFARX1 I_22861 (I391103,I2507,I390625,I390617,);
not I_22862 (I391203,I2514);
DFFARX1 I_22863 (I448680,I2507,I391203,I391229,);
not I_22864 (I391237,I391229);
nand I_22865 (I391254,I448668,I448686);
and I_22866 (I391271,I391254,I448683);
DFFARX1 I_22867 (I391271,I2507,I391203,I391297,);
not I_22868 (I391305,I448674);
DFFARX1 I_22869 (I448671,I2507,I391203,I391331,);
not I_22870 (I391339,I391331);
nor I_22871 (I391356,I391339,I391237);
and I_22872 (I391373,I391356,I448674);
nor I_22873 (I391390,I391339,I391305);
nor I_22874 (I391186,I391297,I391390);
DFFARX1 I_22875 (I448665,I2507,I391203,I391430,);
nor I_22876 (I391438,I391430,I391297);
not I_22877 (I391455,I391438);
not I_22878 (I391472,I391430);
nor I_22879 (I391489,I391472,I391373);
DFFARX1 I_22880 (I391489,I2507,I391203,I391189,);
nand I_22881 (I391520,I448665,I448668);
and I_22882 (I391537,I391520,I448671);
DFFARX1 I_22883 (I391537,I2507,I391203,I391563,);
nor I_22884 (I391571,I391563,I391430);
DFFARX1 I_22885 (I391571,I2507,I391203,I391171,);
nand I_22886 (I391602,I391563,I391472);
nand I_22887 (I391180,I391455,I391602);
not I_22888 (I391633,I391563);
nor I_22889 (I391650,I391633,I391373);
DFFARX1 I_22890 (I391650,I2507,I391203,I391192,);
nor I_22891 (I391681,I448677,I448668);
or I_22892 (I391183,I391430,I391681);
nor I_22893 (I391174,I391563,I391681);
or I_22894 (I391177,I391297,I391681);
DFFARX1 I_22895 (I391681,I2507,I391203,I391195,);
not I_22896 (I391781,I2514);
DFFARX1 I_22897 (I441829,I2507,I391781,I391807,);
not I_22898 (I391815,I391807);
nand I_22899 (I391832,I441817,I441835);
and I_22900 (I391849,I391832,I441832);
DFFARX1 I_22901 (I391849,I2507,I391781,I391875,);
not I_22902 (I391883,I441823);
DFFARX1 I_22903 (I441820,I2507,I391781,I391909,);
not I_22904 (I391917,I391909);
nor I_22905 (I391934,I391917,I391815);
and I_22906 (I391951,I391934,I441823);
nor I_22907 (I391968,I391917,I391883);
nor I_22908 (I391764,I391875,I391968);
DFFARX1 I_22909 (I441814,I2507,I391781,I392008,);
nor I_22910 (I392016,I392008,I391875);
not I_22911 (I392033,I392016);
not I_22912 (I392050,I392008);
nor I_22913 (I392067,I392050,I391951);
DFFARX1 I_22914 (I392067,I2507,I391781,I391767,);
nand I_22915 (I392098,I441814,I441817);
and I_22916 (I392115,I392098,I441820);
DFFARX1 I_22917 (I392115,I2507,I391781,I392141,);
nor I_22918 (I392149,I392141,I392008);
DFFARX1 I_22919 (I392149,I2507,I391781,I391749,);
nand I_22920 (I392180,I392141,I392050);
nand I_22921 (I391758,I392033,I392180);
not I_22922 (I392211,I392141);
nor I_22923 (I392228,I392211,I391951);
DFFARX1 I_22924 (I392228,I2507,I391781,I391770,);
nor I_22925 (I392259,I441826,I441817);
or I_22926 (I391761,I392008,I392259);
nor I_22927 (I391752,I392141,I392259);
or I_22928 (I391755,I391875,I392259);
DFFARX1 I_22929 (I392259,I2507,I391781,I391773,);
not I_22930 (I392359,I2514);
DFFARX1 I_22931 (I162188,I2507,I392359,I392385,);
not I_22932 (I392393,I392385);
nand I_22933 (I392410,I162191,I162167);
and I_22934 (I392427,I392410,I162164);
DFFARX1 I_22935 (I392427,I2507,I392359,I392453,);
not I_22936 (I392461,I162170);
DFFARX1 I_22937 (I162164,I2507,I392359,I392487,);
not I_22938 (I392495,I392487);
nor I_22939 (I392512,I392495,I392393);
and I_22940 (I392529,I392512,I162170);
nor I_22941 (I392546,I392495,I392461);
nor I_22942 (I392342,I392453,I392546);
DFFARX1 I_22943 (I162173,I2507,I392359,I392586,);
nor I_22944 (I392594,I392586,I392453);
not I_22945 (I392611,I392594);
not I_22946 (I392628,I392586);
nor I_22947 (I392645,I392628,I392529);
DFFARX1 I_22948 (I392645,I2507,I392359,I392345,);
nand I_22949 (I392676,I162176,I162185);
and I_22950 (I392693,I392676,I162182);
DFFARX1 I_22951 (I392693,I2507,I392359,I392719,);
nor I_22952 (I392727,I392719,I392586);
DFFARX1 I_22953 (I392727,I2507,I392359,I392327,);
nand I_22954 (I392758,I392719,I392628);
nand I_22955 (I392336,I392611,I392758);
not I_22956 (I392789,I392719);
nor I_22957 (I392806,I392789,I392529);
DFFARX1 I_22958 (I392806,I2507,I392359,I392348,);
nor I_22959 (I392837,I162179,I162185);
or I_22960 (I392339,I392586,I392837);
nor I_22961 (I392330,I392719,I392837);
or I_22962 (I392333,I392453,I392837);
DFFARX1 I_22963 (I392837,I2507,I392359,I392351,);
not I_22964 (I392937,I2514);
DFFARX1 I_22965 (I650149,I2507,I392937,I392963,);
not I_22966 (I392971,I392963);
nand I_22967 (I392988,I650152,I650161);
and I_22968 (I393005,I392988,I650164);
DFFARX1 I_22969 (I393005,I2507,I392937,I393031,);
not I_22970 (I393039,I650173);
DFFARX1 I_22971 (I650155,I2507,I392937,I393065,);
not I_22972 (I393073,I393065);
nor I_22973 (I393090,I393073,I392971);
and I_22974 (I393107,I393090,I650173);
nor I_22975 (I393124,I393073,I393039);
nor I_22976 (I392920,I393031,I393124);
DFFARX1 I_22977 (I650152,I2507,I392937,I393164,);
nor I_22978 (I393172,I393164,I393031);
not I_22979 (I393189,I393172);
not I_22980 (I393206,I393164);
nor I_22981 (I393223,I393206,I393107);
DFFARX1 I_22982 (I393223,I2507,I392937,I392923,);
nand I_22983 (I393254,I650170,I650149);
and I_22984 (I393271,I393254,I650167);
DFFARX1 I_22985 (I393271,I2507,I392937,I393297,);
nor I_22986 (I393305,I393297,I393164);
DFFARX1 I_22987 (I393305,I2507,I392937,I392905,);
nand I_22988 (I393336,I393297,I393206);
nand I_22989 (I392914,I393189,I393336);
not I_22990 (I393367,I393297);
nor I_22991 (I393384,I393367,I393107);
DFFARX1 I_22992 (I393384,I2507,I392937,I392926,);
nor I_22993 (I393415,I650158,I650149);
or I_22994 (I392917,I393164,I393415);
nor I_22995 (I392908,I393297,I393415);
or I_22996 (I392911,I393031,I393415);
DFFARX1 I_22997 (I393415,I2507,I392937,I392929,);
not I_22998 (I393515,I2514);
DFFARX1 I_22999 (I210145,I2507,I393515,I393541,);
not I_23000 (I393549,I393541);
nand I_23001 (I393566,I210148,I210124);
and I_23002 (I393583,I393566,I210121);
DFFARX1 I_23003 (I393583,I2507,I393515,I393609,);
not I_23004 (I393617,I210127);
DFFARX1 I_23005 (I210121,I2507,I393515,I393643,);
not I_23006 (I393651,I393643);
nor I_23007 (I393668,I393651,I393549);
and I_23008 (I393685,I393668,I210127);
nor I_23009 (I393702,I393651,I393617);
nor I_23010 (I393498,I393609,I393702);
DFFARX1 I_23011 (I210130,I2507,I393515,I393742,);
nor I_23012 (I393750,I393742,I393609);
not I_23013 (I393767,I393750);
not I_23014 (I393784,I393742);
nor I_23015 (I393801,I393784,I393685);
DFFARX1 I_23016 (I393801,I2507,I393515,I393501,);
nand I_23017 (I393832,I210133,I210142);
and I_23018 (I393849,I393832,I210139);
DFFARX1 I_23019 (I393849,I2507,I393515,I393875,);
nor I_23020 (I393883,I393875,I393742);
DFFARX1 I_23021 (I393883,I2507,I393515,I393483,);
nand I_23022 (I393914,I393875,I393784);
nand I_23023 (I393492,I393767,I393914);
not I_23024 (I393945,I393875);
nor I_23025 (I393962,I393945,I393685);
DFFARX1 I_23026 (I393962,I2507,I393515,I393504,);
nor I_23027 (I393993,I210136,I210142);
or I_23028 (I393495,I393742,I393993);
nor I_23029 (I393486,I393875,I393993);
or I_23030 (I393489,I393609,I393993);
DFFARX1 I_23031 (I393993,I2507,I393515,I393507,);
not I_23032 (I394093,I2514);
DFFARX1 I_23033 (I118729,I2507,I394093,I394119,);
not I_23034 (I394127,I394119);
nand I_23035 (I394144,I118732,I118753);
and I_23036 (I394161,I394144,I118741);
DFFARX1 I_23037 (I394161,I2507,I394093,I394187,);
not I_23038 (I394195,I118738);
DFFARX1 I_23039 (I118729,I2507,I394093,I394221,);
not I_23040 (I394229,I394221);
nor I_23041 (I394246,I394229,I394127);
and I_23042 (I394263,I394246,I118738);
nor I_23043 (I394280,I394229,I394195);
nor I_23044 (I394076,I394187,I394280);
DFFARX1 I_23045 (I118747,I2507,I394093,I394320,);
nor I_23046 (I394328,I394320,I394187);
not I_23047 (I394345,I394328);
not I_23048 (I394362,I394320);
nor I_23049 (I394379,I394362,I394263);
DFFARX1 I_23050 (I394379,I2507,I394093,I394079,);
nand I_23051 (I394410,I118732,I118735);
and I_23052 (I394427,I394410,I118744);
DFFARX1 I_23053 (I394427,I2507,I394093,I394453,);
nor I_23054 (I394461,I394453,I394320);
DFFARX1 I_23055 (I394461,I2507,I394093,I394061,);
nand I_23056 (I394492,I394453,I394362);
nand I_23057 (I394070,I394345,I394492);
not I_23058 (I394523,I394453);
nor I_23059 (I394540,I394523,I394263);
DFFARX1 I_23060 (I394540,I2507,I394093,I394082,);
nor I_23061 (I394571,I118750,I118735);
or I_23062 (I394073,I394320,I394571);
nor I_23063 (I394064,I394453,I394571);
or I_23064 (I394067,I394187,I394571);
DFFARX1 I_23065 (I394571,I2507,I394093,I394085,);
not I_23066 (I394671,I2514);
DFFARX1 I_23067 (I432870,I2507,I394671,I394697,);
not I_23068 (I394705,I394697);
nand I_23069 (I394722,I432858,I432876);
and I_23070 (I394739,I394722,I432873);
DFFARX1 I_23071 (I394739,I2507,I394671,I394765,);
not I_23072 (I394773,I432864);
DFFARX1 I_23073 (I432861,I2507,I394671,I394799,);
not I_23074 (I394807,I394799);
nor I_23075 (I394824,I394807,I394705);
and I_23076 (I394841,I394824,I432864);
nor I_23077 (I394858,I394807,I394773);
nor I_23078 (I394654,I394765,I394858);
DFFARX1 I_23079 (I432855,I2507,I394671,I394898,);
nor I_23080 (I394906,I394898,I394765);
not I_23081 (I394923,I394906);
not I_23082 (I394940,I394898);
nor I_23083 (I394957,I394940,I394841);
DFFARX1 I_23084 (I394957,I2507,I394671,I394657,);
nand I_23085 (I394988,I432855,I432858);
and I_23086 (I395005,I394988,I432861);
DFFARX1 I_23087 (I395005,I2507,I394671,I395031,);
nor I_23088 (I395039,I395031,I394898);
DFFARX1 I_23089 (I395039,I2507,I394671,I394639,);
nand I_23090 (I395070,I395031,I394940);
nand I_23091 (I394648,I394923,I395070);
not I_23092 (I395101,I395031);
nor I_23093 (I395118,I395101,I394841);
DFFARX1 I_23094 (I395118,I2507,I394671,I394660,);
nor I_23095 (I395149,I432867,I432858);
or I_23096 (I394651,I394898,I395149);
nor I_23097 (I394642,I395031,I395149);
or I_23098 (I394645,I394765,I395149);
DFFARX1 I_23099 (I395149,I2507,I394671,I394663,);
not I_23100 (I395249,I2514);
DFFARX1 I_23101 (I653413,I2507,I395249,I395275,);
not I_23102 (I395283,I395275);
nand I_23103 (I395300,I653416,I653425);
and I_23104 (I395317,I395300,I653428);
DFFARX1 I_23105 (I395317,I2507,I395249,I395343,);
not I_23106 (I395351,I653437);
DFFARX1 I_23107 (I653419,I2507,I395249,I395377,);
not I_23108 (I395385,I395377);
nor I_23109 (I395402,I395385,I395283);
and I_23110 (I395419,I395402,I653437);
nor I_23111 (I395436,I395385,I395351);
nor I_23112 (I395232,I395343,I395436);
DFFARX1 I_23113 (I653416,I2507,I395249,I395476,);
nor I_23114 (I395484,I395476,I395343);
not I_23115 (I395501,I395484);
not I_23116 (I395518,I395476);
nor I_23117 (I395535,I395518,I395419);
DFFARX1 I_23118 (I395535,I2507,I395249,I395235,);
nand I_23119 (I395566,I653434,I653413);
and I_23120 (I395583,I395566,I653431);
DFFARX1 I_23121 (I395583,I2507,I395249,I395609,);
nor I_23122 (I395617,I395609,I395476);
DFFARX1 I_23123 (I395617,I2507,I395249,I395217,);
nand I_23124 (I395648,I395609,I395518);
nand I_23125 (I395226,I395501,I395648);
not I_23126 (I395679,I395609);
nor I_23127 (I395696,I395679,I395419);
DFFARX1 I_23128 (I395696,I2507,I395249,I395238,);
nor I_23129 (I395727,I653422,I653413);
or I_23130 (I395229,I395476,I395727);
nor I_23131 (I395220,I395609,I395727);
or I_23132 (I395223,I395343,I395727);
DFFARX1 I_23133 (I395727,I2507,I395249,I395241,);
not I_23134 (I395827,I2514);
DFFARX1 I_23135 (I80992,I2507,I395827,I395853,);
not I_23136 (I395861,I395853);
nand I_23137 (I395878,I81001,I81010);
and I_23138 (I395895,I395878,I80989);
DFFARX1 I_23139 (I395895,I2507,I395827,I395921,);
not I_23140 (I395929,I80992);
DFFARX1 I_23141 (I81007,I2507,I395827,I395955,);
not I_23142 (I395963,I395955);
nor I_23143 (I395980,I395963,I395861);
and I_23144 (I395997,I395980,I80992);
nor I_23145 (I396014,I395963,I395929);
nor I_23146 (I395810,I395921,I396014);
DFFARX1 I_23147 (I80998,I2507,I395827,I396054,);
nor I_23148 (I396062,I396054,I395921);
not I_23149 (I396079,I396062);
not I_23150 (I396096,I396054);
nor I_23151 (I396113,I396096,I395997);
DFFARX1 I_23152 (I396113,I2507,I395827,I395813,);
nand I_23153 (I396144,I81013,I80989);
and I_23154 (I396161,I396144,I80995);
DFFARX1 I_23155 (I396161,I2507,I395827,I396187,);
nor I_23156 (I396195,I396187,I396054);
DFFARX1 I_23157 (I396195,I2507,I395827,I395795,);
nand I_23158 (I396226,I396187,I396096);
nand I_23159 (I395804,I396079,I396226);
not I_23160 (I396257,I396187);
nor I_23161 (I396274,I396257,I395997);
DFFARX1 I_23162 (I396274,I2507,I395827,I395816,);
nor I_23163 (I396305,I81004,I80989);
or I_23164 (I395807,I396054,I396305);
nor I_23165 (I395798,I396187,I396305);
or I_23166 (I395801,I395921,I396305);
DFFARX1 I_23167 (I396305,I2507,I395827,I395819,);
not I_23168 (I396405,I2514);
DFFARX1 I_23169 (I119324,I2507,I396405,I396431,);
not I_23170 (I396439,I396431);
nand I_23171 (I396456,I119327,I119348);
and I_23172 (I396473,I396456,I119336);
DFFARX1 I_23173 (I396473,I2507,I396405,I396499,);
not I_23174 (I396507,I119333);
DFFARX1 I_23175 (I119324,I2507,I396405,I396533,);
not I_23176 (I396541,I396533);
nor I_23177 (I396558,I396541,I396439);
and I_23178 (I396575,I396558,I119333);
nor I_23179 (I396592,I396541,I396507);
nor I_23180 (I396388,I396499,I396592);
DFFARX1 I_23181 (I119342,I2507,I396405,I396632,);
nor I_23182 (I396640,I396632,I396499);
not I_23183 (I396657,I396640);
not I_23184 (I396674,I396632);
nor I_23185 (I396691,I396674,I396575);
DFFARX1 I_23186 (I396691,I2507,I396405,I396391,);
nand I_23187 (I396722,I119327,I119330);
and I_23188 (I396739,I396722,I119339);
DFFARX1 I_23189 (I396739,I2507,I396405,I396765,);
nor I_23190 (I396773,I396765,I396632);
DFFARX1 I_23191 (I396773,I2507,I396405,I396373,);
nand I_23192 (I396804,I396765,I396674);
nand I_23193 (I396382,I396657,I396804);
not I_23194 (I396835,I396765);
nor I_23195 (I396852,I396835,I396575);
DFFARX1 I_23196 (I396852,I2507,I396405,I396394,);
nor I_23197 (I396883,I119345,I119330);
or I_23198 (I396385,I396632,I396883);
nor I_23199 (I396376,I396765,I396883);
or I_23200 (I396379,I396499,I396883);
DFFARX1 I_23201 (I396883,I2507,I396405,I396397,);
not I_23202 (I396983,I2514);
DFFARX1 I_23203 (I268321,I2507,I396983,I397009,);
not I_23204 (I397017,I397009);
nand I_23205 (I397034,I268312,I268330);
and I_23206 (I397051,I397034,I268333);
DFFARX1 I_23207 (I397051,I2507,I396983,I397077,);
not I_23208 (I397085,I268327);
DFFARX1 I_23209 (I268315,I2507,I396983,I397111,);
not I_23210 (I397119,I397111);
nor I_23211 (I397136,I397119,I397017);
and I_23212 (I397153,I397136,I268327);
nor I_23213 (I397170,I397119,I397085);
nor I_23214 (I396966,I397077,I397170);
DFFARX1 I_23215 (I268324,I2507,I396983,I397210,);
nor I_23216 (I397218,I397210,I397077);
not I_23217 (I397235,I397218);
not I_23218 (I397252,I397210);
nor I_23219 (I397269,I397252,I397153);
DFFARX1 I_23220 (I397269,I2507,I396983,I396969,);
nand I_23221 (I397300,I268339,I268336);
and I_23222 (I397317,I397300,I268318);
DFFARX1 I_23223 (I397317,I2507,I396983,I397343,);
nor I_23224 (I397351,I397343,I397210);
DFFARX1 I_23225 (I397351,I2507,I396983,I396951,);
nand I_23226 (I397382,I397343,I397252);
nand I_23227 (I396960,I397235,I397382);
not I_23228 (I397413,I397343);
nor I_23229 (I397430,I397413,I397153);
DFFARX1 I_23230 (I397430,I2507,I396983,I396972,);
nor I_23231 (I397461,I268312,I268336);
or I_23232 (I396963,I397210,I397461);
nor I_23233 (I396954,I397343,I397461);
or I_23234 (I396957,I397077,I397461);
DFFARX1 I_23235 (I397461,I2507,I396983,I396975,);
not I_23236 (I397561,I2514);
DFFARX1 I_23237 (I683265,I2507,I397561,I397587,);
not I_23238 (I397595,I397587);
nand I_23239 (I397612,I683289,I683271);
and I_23240 (I397629,I397612,I683277);
DFFARX1 I_23241 (I397629,I2507,I397561,I397655,);
not I_23242 (I397663,I683283);
DFFARX1 I_23243 (I683268,I2507,I397561,I397689,);
not I_23244 (I397697,I397689);
nor I_23245 (I397714,I397697,I397595);
and I_23246 (I397731,I397714,I683283);
nor I_23247 (I397748,I397697,I397663);
nor I_23248 (I397544,I397655,I397748);
DFFARX1 I_23249 (I683280,I2507,I397561,I397788,);
nor I_23250 (I397796,I397788,I397655);
not I_23251 (I397813,I397796);
not I_23252 (I397830,I397788);
nor I_23253 (I397847,I397830,I397731);
DFFARX1 I_23254 (I397847,I2507,I397561,I397547,);
nand I_23255 (I397878,I683286,I683274);
and I_23256 (I397895,I397878,I683268);
DFFARX1 I_23257 (I397895,I2507,I397561,I397921,);
nor I_23258 (I397929,I397921,I397788);
DFFARX1 I_23259 (I397929,I2507,I397561,I397529,);
nand I_23260 (I397960,I397921,I397830);
nand I_23261 (I397538,I397813,I397960);
not I_23262 (I397991,I397921);
nor I_23263 (I398008,I397991,I397731);
DFFARX1 I_23264 (I398008,I2507,I397561,I397550,);
nor I_23265 (I398039,I683265,I683274);
or I_23266 (I397541,I397788,I398039);
nor I_23267 (I397532,I397921,I398039);
or I_23268 (I397535,I397655,I398039);
DFFARX1 I_23269 (I398039,I2507,I397561,I397553,);
not I_23270 (I398139,I2514);
DFFARX1 I_23271 (I646341,I2507,I398139,I398165,);
not I_23272 (I398173,I398165);
nand I_23273 (I398190,I646344,I646353);
and I_23274 (I398207,I398190,I646356);
DFFARX1 I_23275 (I398207,I2507,I398139,I398233,);
not I_23276 (I398241,I646365);
DFFARX1 I_23277 (I646347,I2507,I398139,I398267,);
not I_23278 (I398275,I398267);
nor I_23279 (I398292,I398275,I398173);
and I_23280 (I398309,I398292,I646365);
nor I_23281 (I398326,I398275,I398241);
nor I_23282 (I398122,I398233,I398326);
DFFARX1 I_23283 (I646344,I2507,I398139,I398366,);
nor I_23284 (I398374,I398366,I398233);
not I_23285 (I398391,I398374);
not I_23286 (I398408,I398366);
nor I_23287 (I398425,I398408,I398309);
DFFARX1 I_23288 (I398425,I2507,I398139,I398125,);
nand I_23289 (I398456,I646362,I646341);
and I_23290 (I398473,I398456,I646359);
DFFARX1 I_23291 (I398473,I2507,I398139,I398499,);
nor I_23292 (I398507,I398499,I398366);
DFFARX1 I_23293 (I398507,I2507,I398139,I398107,);
nand I_23294 (I398538,I398499,I398408);
nand I_23295 (I398116,I398391,I398538);
not I_23296 (I398569,I398499);
nor I_23297 (I398586,I398569,I398309);
DFFARX1 I_23298 (I398586,I2507,I398139,I398128,);
nor I_23299 (I398617,I646350,I646341);
or I_23300 (I398119,I398366,I398617);
nor I_23301 (I398110,I398499,I398617);
or I_23302 (I398113,I398233,I398617);
DFFARX1 I_23303 (I398617,I2507,I398139,I398131,);
not I_23304 (I398717,I2514);
DFFARX1 I_23305 (I589613,I2507,I398717,I398743,);
not I_23306 (I398751,I398743);
nand I_23307 (I398768,I589595,I589607);
and I_23308 (I398785,I398768,I589610);
DFFARX1 I_23309 (I398785,I2507,I398717,I398811,);
not I_23310 (I398819,I589604);
DFFARX1 I_23311 (I589601,I2507,I398717,I398845,);
not I_23312 (I398853,I398845);
nor I_23313 (I398870,I398853,I398751);
and I_23314 (I398887,I398870,I589604);
nor I_23315 (I398904,I398853,I398819);
nor I_23316 (I398700,I398811,I398904);
DFFARX1 I_23317 (I589619,I2507,I398717,I398944,);
nor I_23318 (I398952,I398944,I398811);
not I_23319 (I398969,I398952);
not I_23320 (I398986,I398944);
nor I_23321 (I399003,I398986,I398887);
DFFARX1 I_23322 (I399003,I2507,I398717,I398703,);
nand I_23323 (I399034,I589598,I589598);
and I_23324 (I399051,I399034,I589595);
DFFARX1 I_23325 (I399051,I2507,I398717,I399077,);
nor I_23326 (I399085,I399077,I398944);
DFFARX1 I_23327 (I399085,I2507,I398717,I398685,);
nand I_23328 (I399116,I399077,I398986);
nand I_23329 (I398694,I398969,I399116);
not I_23330 (I399147,I399077);
nor I_23331 (I399164,I399147,I398887);
DFFARX1 I_23332 (I399164,I2507,I398717,I398706,);
nor I_23333 (I399195,I589616,I589598);
or I_23334 (I398697,I398944,I399195);
nor I_23335 (I398688,I399077,I399195);
or I_23336 (I398691,I398811,I399195);
DFFARX1 I_23337 (I399195,I2507,I398717,I398709,);
not I_23338 (I399295,I2514);
DFFARX1 I_23339 (I31463,I2507,I399295,I399321,);
not I_23340 (I399329,I399321);
nand I_23341 (I399346,I31460,I31451);
and I_23342 (I399363,I399346,I31451);
DFFARX1 I_23343 (I399363,I2507,I399295,I399389,);
not I_23344 (I399397,I31454);
DFFARX1 I_23345 (I31469,I2507,I399295,I399423,);
not I_23346 (I399431,I399423);
nor I_23347 (I399448,I399431,I399329);
and I_23348 (I399465,I399448,I31454);
nor I_23349 (I399482,I399431,I399397);
nor I_23350 (I399278,I399389,I399482);
DFFARX1 I_23351 (I31454,I2507,I399295,I399522,);
nor I_23352 (I399530,I399522,I399389);
not I_23353 (I399547,I399530);
not I_23354 (I399564,I399522);
nor I_23355 (I399581,I399564,I399465);
DFFARX1 I_23356 (I399581,I2507,I399295,I399281,);
nand I_23357 (I399612,I31472,I31457);
and I_23358 (I399629,I399612,I31475);
DFFARX1 I_23359 (I399629,I2507,I399295,I399655,);
nor I_23360 (I399663,I399655,I399522);
DFFARX1 I_23361 (I399663,I2507,I399295,I399263,);
nand I_23362 (I399694,I399655,I399564);
nand I_23363 (I399272,I399547,I399694);
not I_23364 (I399725,I399655);
nor I_23365 (I399742,I399725,I399465);
DFFARX1 I_23366 (I399742,I2507,I399295,I399284,);
nor I_23367 (I399773,I31466,I31457);
or I_23368 (I399275,I399522,I399773);
nor I_23369 (I399266,I399655,I399773);
or I_23370 (I399269,I399389,I399773);
DFFARX1 I_23371 (I399773,I2507,I399295,I399287,);
not I_23372 (I399873,I2514);
DFFARX1 I_23373 (I90764,I2507,I399873,I399899,);
not I_23374 (I399907,I399899);
nand I_23375 (I399924,I90767,I90788);
and I_23376 (I399941,I399924,I90776);
DFFARX1 I_23377 (I399941,I2507,I399873,I399967,);
not I_23378 (I399975,I90773);
DFFARX1 I_23379 (I90764,I2507,I399873,I400001,);
not I_23380 (I400009,I400001);
nor I_23381 (I400026,I400009,I399907);
and I_23382 (I400043,I400026,I90773);
nor I_23383 (I400060,I400009,I399975);
nor I_23384 (I399856,I399967,I400060);
DFFARX1 I_23385 (I90782,I2507,I399873,I400100,);
nor I_23386 (I400108,I400100,I399967);
not I_23387 (I400125,I400108);
not I_23388 (I400142,I400100);
nor I_23389 (I400159,I400142,I400043);
DFFARX1 I_23390 (I400159,I2507,I399873,I399859,);
nand I_23391 (I400190,I90767,I90770);
and I_23392 (I400207,I400190,I90779);
DFFARX1 I_23393 (I400207,I2507,I399873,I400233,);
nor I_23394 (I400241,I400233,I400100);
DFFARX1 I_23395 (I400241,I2507,I399873,I399841,);
nand I_23396 (I400272,I400233,I400142);
nand I_23397 (I399850,I400125,I400272);
not I_23398 (I400303,I400233);
nor I_23399 (I400320,I400303,I400043);
DFFARX1 I_23400 (I400320,I2507,I399873,I399862,);
nor I_23401 (I400351,I90785,I90770);
or I_23402 (I399853,I400100,I400351);
nor I_23403 (I399844,I400233,I400351);
or I_23404 (I399847,I399967,I400351);
DFFARX1 I_23405 (I400351,I2507,I399873,I399865,);
not I_23406 (I400451,I2514);
DFFARX1 I_23407 (I237313,I2507,I400451,I400477,);
not I_23408 (I400485,I400477);
nand I_23409 (I400502,I237304,I237322);
and I_23410 (I400519,I400502,I237325);
DFFARX1 I_23411 (I400519,I2507,I400451,I400545,);
not I_23412 (I400553,I237319);
DFFARX1 I_23413 (I237307,I2507,I400451,I400579,);
not I_23414 (I400587,I400579);
nor I_23415 (I400604,I400587,I400485);
and I_23416 (I400621,I400604,I237319);
nor I_23417 (I400638,I400587,I400553);
nor I_23418 (I400434,I400545,I400638);
DFFARX1 I_23419 (I237316,I2507,I400451,I400678,);
nor I_23420 (I400686,I400678,I400545);
not I_23421 (I400703,I400686);
not I_23422 (I400720,I400678);
nor I_23423 (I400737,I400720,I400621);
DFFARX1 I_23424 (I400737,I2507,I400451,I400437,);
nand I_23425 (I400768,I237331,I237328);
and I_23426 (I400785,I400768,I237310);
DFFARX1 I_23427 (I400785,I2507,I400451,I400811,);
nor I_23428 (I400819,I400811,I400678);
DFFARX1 I_23429 (I400819,I2507,I400451,I400419,);
nand I_23430 (I400850,I400811,I400720);
nand I_23431 (I400428,I400703,I400850);
not I_23432 (I400881,I400811);
nor I_23433 (I400898,I400881,I400621);
DFFARX1 I_23434 (I400898,I2507,I400451,I400440,);
nor I_23435 (I400929,I237304,I237328);
or I_23436 (I400431,I400678,I400929);
nor I_23437 (I400422,I400811,I400929);
or I_23438 (I400425,I400545,I400929);
DFFARX1 I_23439 (I400929,I2507,I400451,I400443,);
not I_23440 (I401029,I2514);
DFFARX1 I_23441 (I474503,I2507,I401029,I401055,);
not I_23442 (I401063,I401055);
nand I_23443 (I401080,I474491,I474509);
and I_23444 (I401097,I401080,I474506);
DFFARX1 I_23445 (I401097,I2507,I401029,I401123,);
not I_23446 (I401131,I474497);
DFFARX1 I_23447 (I474494,I2507,I401029,I401157,);
not I_23448 (I401165,I401157);
nor I_23449 (I401182,I401165,I401063);
and I_23450 (I401199,I401182,I474497);
nor I_23451 (I401216,I401165,I401131);
nor I_23452 (I401012,I401123,I401216);
DFFARX1 I_23453 (I474488,I2507,I401029,I401256,);
nor I_23454 (I401264,I401256,I401123);
not I_23455 (I401281,I401264);
not I_23456 (I401298,I401256);
nor I_23457 (I401315,I401298,I401199);
DFFARX1 I_23458 (I401315,I2507,I401029,I401015,);
nand I_23459 (I401346,I474488,I474491);
and I_23460 (I401363,I401346,I474494);
DFFARX1 I_23461 (I401363,I2507,I401029,I401389,);
nor I_23462 (I401397,I401389,I401256);
DFFARX1 I_23463 (I401397,I2507,I401029,I400997,);
nand I_23464 (I401428,I401389,I401298);
nand I_23465 (I401006,I401281,I401428);
not I_23466 (I401459,I401389);
nor I_23467 (I401476,I401459,I401199);
DFFARX1 I_23468 (I401476,I2507,I401029,I401018,);
nor I_23469 (I401507,I474500,I474491);
or I_23470 (I401009,I401256,I401507);
nor I_23471 (I401000,I401389,I401507);
or I_23472 (I401003,I401123,I401507);
DFFARX1 I_23473 (I401507,I2507,I401029,I401021,);
not I_23474 (I401607,I2514);
DFFARX1 I_23475 (I202240,I2507,I401607,I401633,);
not I_23476 (I401641,I401633);
nand I_23477 (I401658,I202243,I202219);
and I_23478 (I401675,I401658,I202216);
DFFARX1 I_23479 (I401675,I2507,I401607,I401701,);
not I_23480 (I401709,I202222);
DFFARX1 I_23481 (I202216,I2507,I401607,I401735,);
not I_23482 (I401743,I401735);
nor I_23483 (I401760,I401743,I401641);
and I_23484 (I401777,I401760,I202222);
nor I_23485 (I401794,I401743,I401709);
nor I_23486 (I401590,I401701,I401794);
DFFARX1 I_23487 (I202225,I2507,I401607,I401834,);
nor I_23488 (I401842,I401834,I401701);
not I_23489 (I401859,I401842);
not I_23490 (I401876,I401834);
nor I_23491 (I401893,I401876,I401777);
DFFARX1 I_23492 (I401893,I2507,I401607,I401593,);
nand I_23493 (I401924,I202228,I202237);
and I_23494 (I401941,I401924,I202234);
DFFARX1 I_23495 (I401941,I2507,I401607,I401967,);
nor I_23496 (I401975,I401967,I401834);
DFFARX1 I_23497 (I401975,I2507,I401607,I401575,);
nand I_23498 (I402006,I401967,I401876);
nand I_23499 (I401584,I401859,I402006);
not I_23500 (I402037,I401967);
nor I_23501 (I402054,I402037,I401777);
DFFARX1 I_23502 (I402054,I2507,I401607,I401596,);
nor I_23503 (I402085,I202231,I202237);
or I_23504 (I401587,I401834,I402085);
nor I_23505 (I401578,I401967,I402085);
or I_23506 (I401581,I401701,I402085);
DFFARX1 I_23507 (I402085,I2507,I401607,I401599,);
not I_23508 (I402185,I2514);
DFFARX1 I_23509 (I22504,I2507,I402185,I402211,);
not I_23510 (I402219,I402211);
nand I_23511 (I402236,I22501,I22492);
and I_23512 (I402253,I402236,I22492);
DFFARX1 I_23513 (I402253,I2507,I402185,I402279,);
not I_23514 (I402287,I22495);
DFFARX1 I_23515 (I22510,I2507,I402185,I402313,);
not I_23516 (I402321,I402313);
nor I_23517 (I402338,I402321,I402219);
and I_23518 (I402355,I402338,I22495);
nor I_23519 (I402372,I402321,I402287);
nor I_23520 (I402168,I402279,I402372);
DFFARX1 I_23521 (I22495,I2507,I402185,I402412,);
nor I_23522 (I402420,I402412,I402279);
not I_23523 (I402437,I402420);
not I_23524 (I402454,I402412);
nor I_23525 (I402471,I402454,I402355);
DFFARX1 I_23526 (I402471,I2507,I402185,I402171,);
nand I_23527 (I402502,I22513,I22498);
and I_23528 (I402519,I402502,I22516);
DFFARX1 I_23529 (I402519,I2507,I402185,I402545,);
nor I_23530 (I402553,I402545,I402412);
DFFARX1 I_23531 (I402553,I2507,I402185,I402153,);
nand I_23532 (I402584,I402545,I402454);
nand I_23533 (I402162,I402437,I402584);
not I_23534 (I402615,I402545);
nor I_23535 (I402632,I402615,I402355);
DFFARX1 I_23536 (I402632,I2507,I402185,I402174,);
nor I_23537 (I402663,I22507,I22498);
or I_23538 (I402165,I402412,I402663);
nor I_23539 (I402156,I402545,I402663);
or I_23540 (I402159,I402279,I402663);
DFFARX1 I_23541 (I402663,I2507,I402185,I402177,);
not I_23542 (I402763,I2514);
DFFARX1 I_23543 (I477138,I2507,I402763,I402789,);
not I_23544 (I402797,I402789);
nand I_23545 (I402814,I477126,I477144);
and I_23546 (I402831,I402814,I477141);
DFFARX1 I_23547 (I402831,I2507,I402763,I402857,);
not I_23548 (I402865,I477132);
DFFARX1 I_23549 (I477129,I2507,I402763,I402891,);
not I_23550 (I402899,I402891);
nor I_23551 (I402916,I402899,I402797);
and I_23552 (I402933,I402916,I477132);
nor I_23553 (I402950,I402899,I402865);
nor I_23554 (I402746,I402857,I402950);
DFFARX1 I_23555 (I477123,I2507,I402763,I402990,);
nor I_23556 (I402998,I402990,I402857);
not I_23557 (I403015,I402998);
not I_23558 (I403032,I402990);
nor I_23559 (I403049,I403032,I402933);
DFFARX1 I_23560 (I403049,I2507,I402763,I402749,);
nand I_23561 (I403080,I477123,I477126);
and I_23562 (I403097,I403080,I477129);
DFFARX1 I_23563 (I403097,I2507,I402763,I403123,);
nor I_23564 (I403131,I403123,I402990);
DFFARX1 I_23565 (I403131,I2507,I402763,I402731,);
nand I_23566 (I403162,I403123,I403032);
nand I_23567 (I402740,I403015,I403162);
not I_23568 (I403193,I403123);
nor I_23569 (I403210,I403193,I402933);
DFFARX1 I_23570 (I403210,I2507,I402763,I402752,);
nor I_23571 (I403241,I477135,I477126);
or I_23572 (I402743,I402990,I403241);
nor I_23573 (I402734,I403123,I403241);
or I_23574 (I402737,I402857,I403241);
DFFARX1 I_23575 (I403241,I2507,I402763,I402755,);
not I_23576 (I403341,I2514);
DFFARX1 I_23577 (I116944,I2507,I403341,I403367,);
not I_23578 (I403375,I403367);
nand I_23579 (I403392,I116947,I116968);
and I_23580 (I403409,I403392,I116956);
DFFARX1 I_23581 (I403409,I2507,I403341,I403435,);
not I_23582 (I403443,I116953);
DFFARX1 I_23583 (I116944,I2507,I403341,I403469,);
not I_23584 (I403477,I403469);
nor I_23585 (I403494,I403477,I403375);
and I_23586 (I403511,I403494,I116953);
nor I_23587 (I403528,I403477,I403443);
nor I_23588 (I403324,I403435,I403528);
DFFARX1 I_23589 (I116962,I2507,I403341,I403568,);
nor I_23590 (I403576,I403568,I403435);
not I_23591 (I403593,I403576);
not I_23592 (I403610,I403568);
nor I_23593 (I403627,I403610,I403511);
DFFARX1 I_23594 (I403627,I2507,I403341,I403327,);
nand I_23595 (I403658,I116947,I116950);
and I_23596 (I403675,I403658,I116959);
DFFARX1 I_23597 (I403675,I2507,I403341,I403701,);
nor I_23598 (I403709,I403701,I403568);
DFFARX1 I_23599 (I403709,I2507,I403341,I403309,);
nand I_23600 (I403740,I403701,I403610);
nand I_23601 (I403318,I403593,I403740);
not I_23602 (I403771,I403701);
nor I_23603 (I403788,I403771,I403511);
DFFARX1 I_23604 (I403788,I2507,I403341,I403330,);
nor I_23605 (I403819,I116965,I116950);
or I_23606 (I403321,I403568,I403819);
nor I_23607 (I403312,I403701,I403819);
or I_23608 (I403315,I403435,I403819);
DFFARX1 I_23609 (I403819,I2507,I403341,I403333,);
not I_23610 (I403919,I2514);
DFFARX1 I_23611 (I697810,I2507,I403919,I403945,);
not I_23612 (I403953,I403945);
nand I_23613 (I403970,I697795,I697783);
and I_23614 (I403987,I403970,I697798);
DFFARX1 I_23615 (I403987,I2507,I403919,I404013,);
not I_23616 (I404021,I697783);
DFFARX1 I_23617 (I697801,I2507,I403919,I404047,);
not I_23618 (I404055,I404047);
nor I_23619 (I404072,I404055,I403953);
and I_23620 (I404089,I404072,I697783);
nor I_23621 (I404106,I404055,I404021);
nor I_23622 (I403902,I404013,I404106);
DFFARX1 I_23623 (I697789,I2507,I403919,I404146,);
nor I_23624 (I404154,I404146,I404013);
not I_23625 (I404171,I404154);
not I_23626 (I404188,I404146);
nor I_23627 (I404205,I404188,I404089);
DFFARX1 I_23628 (I404205,I2507,I403919,I403905,);
nand I_23629 (I404236,I697786,I697792);
and I_23630 (I404253,I404236,I697807);
DFFARX1 I_23631 (I404253,I2507,I403919,I404279,);
nor I_23632 (I404287,I404279,I404146);
DFFARX1 I_23633 (I404287,I2507,I403919,I403887,);
nand I_23634 (I404318,I404279,I404188);
nand I_23635 (I403896,I404171,I404318);
not I_23636 (I404349,I404279);
nor I_23637 (I404366,I404349,I404089);
DFFARX1 I_23638 (I404366,I2507,I403919,I403908,);
nor I_23639 (I404397,I697804,I697792);
or I_23640 (I403899,I404146,I404397);
nor I_23641 (I403890,I404279,I404397);
or I_23642 (I403893,I404013,I404397);
DFFARX1 I_23643 (I404397,I2507,I403919,I403911,);
not I_23644 (I404497,I2514);
DFFARX1 I_23645 (I715065,I2507,I404497,I404523,);
not I_23646 (I404531,I404523);
nand I_23647 (I404548,I715050,I715038);
and I_23648 (I404565,I404548,I715053);
DFFARX1 I_23649 (I404565,I2507,I404497,I404591,);
not I_23650 (I404599,I715038);
DFFARX1 I_23651 (I715056,I2507,I404497,I404625,);
not I_23652 (I404633,I404625);
nor I_23653 (I404650,I404633,I404531);
and I_23654 (I404667,I404650,I715038);
nor I_23655 (I404684,I404633,I404599);
nor I_23656 (I404480,I404591,I404684);
DFFARX1 I_23657 (I715044,I2507,I404497,I404724,);
nor I_23658 (I404732,I404724,I404591);
not I_23659 (I404749,I404732);
not I_23660 (I404766,I404724);
nor I_23661 (I404783,I404766,I404667);
DFFARX1 I_23662 (I404783,I2507,I404497,I404483,);
nand I_23663 (I404814,I715041,I715047);
and I_23664 (I404831,I404814,I715062);
DFFARX1 I_23665 (I404831,I2507,I404497,I404857,);
nor I_23666 (I404865,I404857,I404724);
DFFARX1 I_23667 (I404865,I2507,I404497,I404465,);
nand I_23668 (I404896,I404857,I404766);
nand I_23669 (I404474,I404749,I404896);
not I_23670 (I404927,I404857);
nor I_23671 (I404944,I404927,I404667);
DFFARX1 I_23672 (I404944,I2507,I404497,I404486,);
nor I_23673 (I404975,I715059,I715047);
or I_23674 (I404477,I404724,I404975);
nor I_23675 (I404468,I404857,I404975);
or I_23676 (I404471,I404591,I404975);
DFFARX1 I_23677 (I404975,I2507,I404497,I404489,);
not I_23678 (I405075,I2514);
DFFARX1 I_23679 (I246017,I2507,I405075,I405101,);
not I_23680 (I405109,I405101);
nand I_23681 (I405126,I246008,I246026);
and I_23682 (I405143,I405126,I246029);
DFFARX1 I_23683 (I405143,I2507,I405075,I405169,);
not I_23684 (I405177,I246023);
DFFARX1 I_23685 (I246011,I2507,I405075,I405203,);
not I_23686 (I405211,I405203);
nor I_23687 (I405228,I405211,I405109);
and I_23688 (I405245,I405228,I246023);
nor I_23689 (I405262,I405211,I405177);
nor I_23690 (I405058,I405169,I405262);
DFFARX1 I_23691 (I246020,I2507,I405075,I405302,);
nor I_23692 (I405310,I405302,I405169);
not I_23693 (I405327,I405310);
not I_23694 (I405344,I405302);
nor I_23695 (I405361,I405344,I405245);
DFFARX1 I_23696 (I405361,I2507,I405075,I405061,);
nand I_23697 (I405392,I246035,I246032);
and I_23698 (I405409,I405392,I246014);
DFFARX1 I_23699 (I405409,I2507,I405075,I405435,);
nor I_23700 (I405443,I405435,I405302);
DFFARX1 I_23701 (I405443,I2507,I405075,I405043,);
nand I_23702 (I405474,I405435,I405344);
nand I_23703 (I405052,I405327,I405474);
not I_23704 (I405505,I405435);
nor I_23705 (I405522,I405505,I405245);
DFFARX1 I_23706 (I405522,I2507,I405075,I405064,);
nor I_23707 (I405553,I246008,I246032);
or I_23708 (I405055,I405302,I405553);
nor I_23709 (I405046,I405435,I405553);
or I_23710 (I405049,I405169,I405553);
DFFARX1 I_23711 (I405553,I2507,I405075,I405067,);
not I_23712 (I405653,I2514);
DFFARX1 I_23713 (I459747,I2507,I405653,I405679,);
not I_23714 (I405687,I405679);
nand I_23715 (I405704,I459735,I459753);
and I_23716 (I405721,I405704,I459750);
DFFARX1 I_23717 (I405721,I2507,I405653,I405747,);
not I_23718 (I405755,I459741);
DFFARX1 I_23719 (I459738,I2507,I405653,I405781,);
not I_23720 (I405789,I405781);
nor I_23721 (I405806,I405789,I405687);
and I_23722 (I405823,I405806,I459741);
nor I_23723 (I405840,I405789,I405755);
nor I_23724 (I405636,I405747,I405840);
DFFARX1 I_23725 (I459732,I2507,I405653,I405880,);
nor I_23726 (I405888,I405880,I405747);
not I_23727 (I405905,I405888);
not I_23728 (I405922,I405880);
nor I_23729 (I405939,I405922,I405823);
DFFARX1 I_23730 (I405939,I2507,I405653,I405639,);
nand I_23731 (I405970,I459732,I459735);
and I_23732 (I405987,I405970,I459738);
DFFARX1 I_23733 (I405987,I2507,I405653,I406013,);
nor I_23734 (I406021,I406013,I405880);
DFFARX1 I_23735 (I406021,I2507,I405653,I405621,);
nand I_23736 (I406052,I406013,I405922);
nand I_23737 (I405630,I405905,I406052);
not I_23738 (I406083,I406013);
nor I_23739 (I406100,I406083,I405823);
DFFARX1 I_23740 (I406100,I2507,I405653,I405642,);
nor I_23741 (I406131,I459744,I459735);
or I_23742 (I405633,I405880,I406131);
nor I_23743 (I405624,I406013,I406131);
or I_23744 (I405627,I405747,I406131);
DFFARX1 I_23745 (I406131,I2507,I405653,I405645,);
not I_23746 (I406231,I2514);
DFFARX1 I_23747 (I546965,I2507,I406231,I406257,);
not I_23748 (I406265,I406257);
nand I_23749 (I406282,I546962,I546980);
and I_23750 (I406299,I406282,I546977);
DFFARX1 I_23751 (I406299,I2507,I406231,I406325,);
not I_23752 (I406333,I546959);
DFFARX1 I_23753 (I546962,I2507,I406231,I406359,);
not I_23754 (I406367,I406359);
nor I_23755 (I406384,I406367,I406265);
and I_23756 (I406401,I406384,I546959);
nor I_23757 (I406418,I406367,I406333);
nor I_23758 (I406214,I406325,I406418);
DFFARX1 I_23759 (I546971,I2507,I406231,I406458,);
nor I_23760 (I406466,I406458,I406325);
not I_23761 (I406483,I406466);
not I_23762 (I406500,I406458);
nor I_23763 (I406517,I406500,I406401);
DFFARX1 I_23764 (I406517,I2507,I406231,I406217,);
nand I_23765 (I406548,I546974,I546959);
and I_23766 (I406565,I406548,I546965);
DFFARX1 I_23767 (I406565,I2507,I406231,I406591,);
nor I_23768 (I406599,I406591,I406458);
DFFARX1 I_23769 (I406599,I2507,I406231,I406199,);
nand I_23770 (I406630,I406591,I406500);
nand I_23771 (I406208,I406483,I406630);
not I_23772 (I406661,I406591);
nor I_23773 (I406678,I406661,I406401);
DFFARX1 I_23774 (I406678,I2507,I406231,I406220,);
nor I_23775 (I406709,I546968,I546959);
or I_23776 (I406211,I406458,I406709);
nor I_23777 (I406202,I406591,I406709);
or I_23778 (I406205,I406325,I406709);
DFFARX1 I_23779 (I406709,I2507,I406231,I406223,);
not I_23780 (I406809,I2514);
DFFARX1 I_23781 (I119919,I2507,I406809,I406835,);
not I_23782 (I406843,I406835);
nand I_23783 (I406860,I119922,I119943);
and I_23784 (I406877,I406860,I119931);
DFFARX1 I_23785 (I406877,I2507,I406809,I406903,);
not I_23786 (I406911,I119928);
DFFARX1 I_23787 (I119919,I2507,I406809,I406937,);
not I_23788 (I406945,I406937);
nor I_23789 (I406962,I406945,I406843);
and I_23790 (I406979,I406962,I119928);
nor I_23791 (I406996,I406945,I406911);
nor I_23792 (I406792,I406903,I406996);
DFFARX1 I_23793 (I119937,I2507,I406809,I407036,);
nor I_23794 (I407044,I407036,I406903);
not I_23795 (I407061,I407044);
not I_23796 (I407078,I407036);
nor I_23797 (I407095,I407078,I406979);
DFFARX1 I_23798 (I407095,I2507,I406809,I406795,);
nand I_23799 (I407126,I119922,I119925);
and I_23800 (I407143,I407126,I119934);
DFFARX1 I_23801 (I407143,I2507,I406809,I407169,);
nor I_23802 (I407177,I407169,I407036);
DFFARX1 I_23803 (I407177,I2507,I406809,I406777,);
nand I_23804 (I407208,I407169,I407078);
nand I_23805 (I406786,I407061,I407208);
not I_23806 (I407239,I407169);
nor I_23807 (I407256,I407239,I406979);
DFFARX1 I_23808 (I407256,I2507,I406809,I406798,);
nor I_23809 (I407287,I119940,I119925);
or I_23810 (I406789,I407036,I407287);
nor I_23811 (I406780,I407169,I407287);
or I_23812 (I406783,I406903,I407287);
DFFARX1 I_23813 (I407287,I2507,I406809,I406801,);
not I_23814 (I407387,I2514);
DFFARX1 I_23815 (I503514,I2507,I407387,I407413,);
not I_23816 (I407421,I407413);
nand I_23817 (I407438,I503490,I503505);
and I_23818 (I407455,I407438,I503517);
DFFARX1 I_23819 (I407455,I2507,I407387,I407481,);
not I_23820 (I407489,I503502);
DFFARX1 I_23821 (I503493,I2507,I407387,I407515,);
not I_23822 (I407523,I407515);
nor I_23823 (I407540,I407523,I407421);
and I_23824 (I407557,I407540,I503502);
nor I_23825 (I407574,I407523,I407489);
nor I_23826 (I407370,I407481,I407574);
DFFARX1 I_23827 (I503490,I2507,I407387,I407614,);
nor I_23828 (I407622,I407614,I407481);
not I_23829 (I407639,I407622);
not I_23830 (I407656,I407614);
nor I_23831 (I407673,I407656,I407557);
DFFARX1 I_23832 (I407673,I2507,I407387,I407373,);
nand I_23833 (I407704,I503508,I503499);
and I_23834 (I407721,I407704,I503511);
DFFARX1 I_23835 (I407721,I2507,I407387,I407747,);
nor I_23836 (I407755,I407747,I407614);
DFFARX1 I_23837 (I407755,I2507,I407387,I407355,);
nand I_23838 (I407786,I407747,I407656);
nand I_23839 (I407364,I407639,I407786);
not I_23840 (I407817,I407747);
nor I_23841 (I407834,I407817,I407557);
DFFARX1 I_23842 (I407834,I2507,I407387,I407376,);
nor I_23843 (I407865,I503496,I503499);
or I_23844 (I407367,I407614,I407865);
nor I_23845 (I407358,I407747,I407865);
or I_23846 (I407361,I407481,I407865);
DFFARX1 I_23847 (I407865,I2507,I407387,I407379,);
not I_23848 (I407965,I2514);
DFFARX1 I_23849 (I509328,I2507,I407965,I407991,);
not I_23850 (I407999,I407991);
nand I_23851 (I408016,I509304,I509319);
and I_23852 (I408033,I408016,I509331);
DFFARX1 I_23853 (I408033,I2507,I407965,I408059,);
not I_23854 (I408067,I509316);
DFFARX1 I_23855 (I509307,I2507,I407965,I408093,);
not I_23856 (I408101,I408093);
nor I_23857 (I408118,I408101,I407999);
and I_23858 (I408135,I408118,I509316);
nor I_23859 (I408152,I408101,I408067);
nor I_23860 (I407948,I408059,I408152);
DFFARX1 I_23861 (I509304,I2507,I407965,I408192,);
nor I_23862 (I408200,I408192,I408059);
not I_23863 (I408217,I408200);
not I_23864 (I408234,I408192);
nor I_23865 (I408251,I408234,I408135);
DFFARX1 I_23866 (I408251,I2507,I407965,I407951,);
nand I_23867 (I408282,I509322,I509313);
and I_23868 (I408299,I408282,I509325);
DFFARX1 I_23869 (I408299,I2507,I407965,I408325,);
nor I_23870 (I408333,I408325,I408192);
DFFARX1 I_23871 (I408333,I2507,I407965,I407933,);
nand I_23872 (I408364,I408325,I408234);
nand I_23873 (I407942,I408217,I408364);
not I_23874 (I408395,I408325);
nor I_23875 (I408412,I408395,I408135);
DFFARX1 I_23876 (I408412,I2507,I407965,I407954,);
nor I_23877 (I408443,I509310,I509313);
or I_23878 (I407945,I408192,I408443);
nor I_23879 (I407936,I408325,I408443);
or I_23880 (I407939,I408059,I408443);
DFFARX1 I_23881 (I408443,I2507,I407965,I407957,);
not I_23882 (I408543,I2514);
DFFARX1 I_23883 (I555380,I2507,I408543,I408569,);
not I_23884 (I408577,I408569);
nand I_23885 (I408594,I555377,I555395);
and I_23886 (I408611,I408594,I555392);
DFFARX1 I_23887 (I408611,I2507,I408543,I408637,);
not I_23888 (I408645,I555374);
DFFARX1 I_23889 (I555377,I2507,I408543,I408671,);
not I_23890 (I408679,I408671);
nor I_23891 (I408696,I408679,I408577);
and I_23892 (I408713,I408696,I555374);
nor I_23893 (I408730,I408679,I408645);
nor I_23894 (I408526,I408637,I408730);
DFFARX1 I_23895 (I555386,I2507,I408543,I408770,);
nor I_23896 (I408778,I408770,I408637);
not I_23897 (I408795,I408778);
not I_23898 (I408812,I408770);
nor I_23899 (I408829,I408812,I408713);
DFFARX1 I_23900 (I408829,I2507,I408543,I408529,);
nand I_23901 (I408860,I555389,I555374);
and I_23902 (I408877,I408860,I555380);
DFFARX1 I_23903 (I408877,I2507,I408543,I408903,);
nor I_23904 (I408911,I408903,I408770);
DFFARX1 I_23905 (I408911,I2507,I408543,I408511,);
nand I_23906 (I408942,I408903,I408812);
nand I_23907 (I408520,I408795,I408942);
not I_23908 (I408973,I408903);
nor I_23909 (I408990,I408973,I408713);
DFFARX1 I_23910 (I408990,I2507,I408543,I408532,);
nor I_23911 (I409021,I555383,I555374);
or I_23912 (I408523,I408770,I409021);
nor I_23913 (I408514,I408903,I409021);
or I_23914 (I408517,I408637,I409021);
DFFARX1 I_23915 (I409021,I2507,I408543,I408535,);
not I_23916 (I409121,I2514);
DFFARX1 I_23917 (I656133,I2507,I409121,I409147,);
not I_23918 (I409155,I409147);
nand I_23919 (I409172,I656136,I656145);
and I_23920 (I409189,I409172,I656148);
DFFARX1 I_23921 (I409189,I2507,I409121,I409215,);
not I_23922 (I409223,I656157);
DFFARX1 I_23923 (I656139,I2507,I409121,I409249,);
not I_23924 (I409257,I409249);
nor I_23925 (I409274,I409257,I409155);
and I_23926 (I409291,I409274,I656157);
nor I_23927 (I409308,I409257,I409223);
nor I_23928 (I409104,I409215,I409308);
DFFARX1 I_23929 (I656136,I2507,I409121,I409348,);
nor I_23930 (I409356,I409348,I409215);
not I_23931 (I409373,I409356);
not I_23932 (I409390,I409348);
nor I_23933 (I409407,I409390,I409291);
DFFARX1 I_23934 (I409407,I2507,I409121,I409107,);
nand I_23935 (I409438,I656154,I656133);
and I_23936 (I409455,I409438,I656151);
DFFARX1 I_23937 (I409455,I2507,I409121,I409481,);
nor I_23938 (I409489,I409481,I409348);
DFFARX1 I_23939 (I409489,I2507,I409121,I409089,);
nand I_23940 (I409520,I409481,I409390);
nand I_23941 (I409098,I409373,I409520);
not I_23942 (I409551,I409481);
nor I_23943 (I409568,I409551,I409291);
DFFARX1 I_23944 (I409568,I2507,I409121,I409110,);
nor I_23945 (I409599,I656142,I656133);
or I_23946 (I409101,I409348,I409599);
nor I_23947 (I409092,I409481,I409599);
or I_23948 (I409095,I409215,I409599);
DFFARX1 I_23949 (I409599,I2507,I409121,I409113,);
not I_23950 (I409699,I2514);
DFFARX1 I_23951 (I164296,I2507,I409699,I409725,);
not I_23952 (I409733,I409725);
nand I_23953 (I409750,I164299,I164275);
and I_23954 (I409767,I409750,I164272);
DFFARX1 I_23955 (I409767,I2507,I409699,I409793,);
not I_23956 (I409801,I164278);
DFFARX1 I_23957 (I164272,I2507,I409699,I409827,);
not I_23958 (I409835,I409827);
nor I_23959 (I409852,I409835,I409733);
and I_23960 (I409869,I409852,I164278);
nor I_23961 (I409886,I409835,I409801);
nor I_23962 (I409682,I409793,I409886);
DFFARX1 I_23963 (I164281,I2507,I409699,I409926,);
nor I_23964 (I409934,I409926,I409793);
not I_23965 (I409951,I409934);
not I_23966 (I409968,I409926);
nor I_23967 (I409985,I409968,I409869);
DFFARX1 I_23968 (I409985,I2507,I409699,I409685,);
nand I_23969 (I410016,I164284,I164293);
and I_23970 (I410033,I410016,I164290);
DFFARX1 I_23971 (I410033,I2507,I409699,I410059,);
nor I_23972 (I410067,I410059,I409926);
DFFARX1 I_23973 (I410067,I2507,I409699,I409667,);
nand I_23974 (I410098,I410059,I409968);
nand I_23975 (I409676,I409951,I410098);
not I_23976 (I410129,I410059);
nor I_23977 (I410146,I410129,I409869);
DFFARX1 I_23978 (I410146,I2507,I409699,I409688,);
nor I_23979 (I410177,I164287,I164293);
or I_23980 (I409679,I409926,I410177);
nor I_23981 (I409670,I410059,I410177);
or I_23982 (I409673,I409793,I410177);
DFFARX1 I_23983 (I410177,I2507,I409699,I409691,);
not I_23984 (I410277,I2514);
DFFARX1 I_23985 (I693645,I2507,I410277,I410303,);
not I_23986 (I410311,I410303);
nand I_23987 (I410328,I693630,I693618);
and I_23988 (I410345,I410328,I693633);
DFFARX1 I_23989 (I410345,I2507,I410277,I410371,);
not I_23990 (I410379,I693618);
DFFARX1 I_23991 (I693636,I2507,I410277,I410405,);
not I_23992 (I410413,I410405);
nor I_23993 (I410430,I410413,I410311);
and I_23994 (I410447,I410430,I693618);
nor I_23995 (I410464,I410413,I410379);
nor I_23996 (I410260,I410371,I410464);
DFFARX1 I_23997 (I693624,I2507,I410277,I410504,);
nor I_23998 (I410512,I410504,I410371);
not I_23999 (I410529,I410512);
not I_24000 (I410546,I410504);
nor I_24001 (I410563,I410546,I410447);
DFFARX1 I_24002 (I410563,I2507,I410277,I410263,);
nand I_24003 (I410594,I693621,I693627);
and I_24004 (I410611,I410594,I693642);
DFFARX1 I_24005 (I410611,I2507,I410277,I410637,);
nor I_24006 (I410645,I410637,I410504);
DFFARX1 I_24007 (I410645,I2507,I410277,I410245,);
nand I_24008 (I410676,I410637,I410546);
nand I_24009 (I410254,I410529,I410676);
not I_24010 (I410707,I410637);
nor I_24011 (I410724,I410707,I410447);
DFFARX1 I_24012 (I410724,I2507,I410277,I410266,);
nor I_24013 (I410755,I693639,I693627);
or I_24014 (I410257,I410504,I410755);
nor I_24015 (I410248,I410637,I410755);
or I_24016 (I410251,I410371,I410755);
DFFARX1 I_24017 (I410755,I2507,I410277,I410269,);
not I_24018 (I410855,I2514);
DFFARX1 I_24019 (I204875,I2507,I410855,I410881,);
not I_24020 (I410889,I410881);
nand I_24021 (I410906,I204878,I204854);
and I_24022 (I410923,I410906,I204851);
DFFARX1 I_24023 (I410923,I2507,I410855,I410949,);
not I_24024 (I410957,I204857);
DFFARX1 I_24025 (I204851,I2507,I410855,I410983,);
not I_24026 (I410991,I410983);
nor I_24027 (I411008,I410991,I410889);
and I_24028 (I411025,I411008,I204857);
nor I_24029 (I411042,I410991,I410957);
nor I_24030 (I410838,I410949,I411042);
DFFARX1 I_24031 (I204860,I2507,I410855,I411082,);
nor I_24032 (I411090,I411082,I410949);
not I_24033 (I411107,I411090);
not I_24034 (I411124,I411082);
nor I_24035 (I411141,I411124,I411025);
DFFARX1 I_24036 (I411141,I2507,I410855,I410841,);
nand I_24037 (I411172,I204863,I204872);
and I_24038 (I411189,I411172,I204869);
DFFARX1 I_24039 (I411189,I2507,I410855,I411215,);
nor I_24040 (I411223,I411215,I411082);
DFFARX1 I_24041 (I411223,I2507,I410855,I410823,);
nand I_24042 (I411254,I411215,I411124);
nand I_24043 (I410832,I411107,I411254);
not I_24044 (I411285,I411215);
nor I_24045 (I411302,I411285,I411025);
DFFARX1 I_24046 (I411302,I2507,I410855,I410844,);
nor I_24047 (I411333,I204866,I204872);
or I_24048 (I410835,I411082,I411333);
nor I_24049 (I410826,I411215,I411333);
or I_24050 (I410829,I410949,I411333);
DFFARX1 I_24051 (I411333,I2507,I410855,I410847,);
not I_24052 (I411433,I2514);
DFFARX1 I_24053 (I176417,I2507,I411433,I411459,);
not I_24054 (I411467,I411459);
nand I_24055 (I411484,I176420,I176396);
and I_24056 (I411501,I411484,I176393);
DFFARX1 I_24057 (I411501,I2507,I411433,I411527,);
not I_24058 (I411535,I176399);
DFFARX1 I_24059 (I176393,I2507,I411433,I411561,);
not I_24060 (I411569,I411561);
nor I_24061 (I411586,I411569,I411467);
and I_24062 (I411603,I411586,I176399);
nor I_24063 (I411620,I411569,I411535);
nor I_24064 (I411416,I411527,I411620);
DFFARX1 I_24065 (I176402,I2507,I411433,I411660,);
nor I_24066 (I411668,I411660,I411527);
not I_24067 (I411685,I411668);
not I_24068 (I411702,I411660);
nor I_24069 (I411719,I411702,I411603);
DFFARX1 I_24070 (I411719,I2507,I411433,I411419,);
nand I_24071 (I411750,I176405,I176414);
and I_24072 (I411767,I411750,I176411);
DFFARX1 I_24073 (I411767,I2507,I411433,I411793,);
nor I_24074 (I411801,I411793,I411660);
DFFARX1 I_24075 (I411801,I2507,I411433,I411401,);
nand I_24076 (I411832,I411793,I411702);
nand I_24077 (I411410,I411685,I411832);
not I_24078 (I411863,I411793);
nor I_24079 (I411880,I411863,I411603);
DFFARX1 I_24080 (I411880,I2507,I411433,I411422,);
nor I_24081 (I411911,I176408,I176414);
or I_24082 (I411413,I411660,I411911);
nor I_24083 (I411404,I411793,I411911);
or I_24084 (I411407,I411527,I411911);
DFFARX1 I_24085 (I411911,I2507,I411433,I411425,);
not I_24086 (I412011,I2514);
DFFARX1 I_24087 (I314297,I2507,I412011,I412037,);
not I_24088 (I412045,I412037);
nand I_24089 (I412062,I314306,I314315);
and I_24090 (I412079,I412062,I314321);
DFFARX1 I_24091 (I412079,I2507,I412011,I412105,);
not I_24092 (I412113,I314318);
DFFARX1 I_24093 (I314303,I2507,I412011,I412139,);
not I_24094 (I412147,I412139);
nor I_24095 (I412164,I412147,I412045);
and I_24096 (I412181,I412164,I314318);
nor I_24097 (I412198,I412147,I412113);
nor I_24098 (I411994,I412105,I412198);
DFFARX1 I_24099 (I314312,I2507,I412011,I412238,);
nor I_24100 (I412246,I412238,I412105);
not I_24101 (I412263,I412246);
not I_24102 (I412280,I412238);
nor I_24103 (I412297,I412280,I412181);
DFFARX1 I_24104 (I412297,I2507,I412011,I411997,);
nand I_24105 (I412328,I314309,I314300);
and I_24106 (I412345,I412328,I314297);
DFFARX1 I_24107 (I412345,I2507,I412011,I412371,);
nor I_24108 (I412379,I412371,I412238);
DFFARX1 I_24109 (I412379,I2507,I412011,I411979,);
nand I_24110 (I412410,I412371,I412280);
nand I_24111 (I411988,I412263,I412410);
not I_24112 (I412441,I412371);
nor I_24113 (I412458,I412441,I412181);
DFFARX1 I_24114 (I412458,I2507,I412011,I412000,);
nor I_24115 (I412489,I314300,I314300);
or I_24116 (I411991,I412238,I412489);
nor I_24117 (I411982,I412371,I412489);
or I_24118 (I411985,I412105,I412489);
DFFARX1 I_24119 (I412489,I2507,I412011,I412003,);
not I_24120 (I412589,I2514);
DFFARX1 I_24121 (I688346,I2507,I412589,I412615,);
not I_24122 (I412623,I412615);
nand I_24123 (I412640,I688334,I688352);
and I_24124 (I412657,I412640,I688343);
DFFARX1 I_24125 (I412657,I2507,I412589,I412683,);
not I_24126 (I412691,I688358);
DFFARX1 I_24127 (I688355,I2507,I412589,I412717,);
not I_24128 (I412725,I412717);
nor I_24129 (I412742,I412725,I412623);
and I_24130 (I412759,I412742,I688358);
nor I_24131 (I412776,I412725,I412691);
nor I_24132 (I412572,I412683,I412776);
DFFARX1 I_24133 (I688337,I2507,I412589,I412816,);
nor I_24134 (I412824,I412816,I412683);
not I_24135 (I412841,I412824);
not I_24136 (I412858,I412816);
nor I_24137 (I412875,I412858,I412759);
DFFARX1 I_24138 (I412875,I2507,I412589,I412575,);
nand I_24139 (I412906,I688331,I688331);
and I_24140 (I412923,I412906,I688340);
DFFARX1 I_24141 (I412923,I2507,I412589,I412949,);
nor I_24142 (I412957,I412949,I412816);
DFFARX1 I_24143 (I412957,I2507,I412589,I412557,);
nand I_24144 (I412988,I412949,I412858);
nand I_24145 (I412566,I412841,I412988);
not I_24146 (I413019,I412949);
nor I_24147 (I413036,I413019,I412759);
DFFARX1 I_24148 (I413036,I2507,I412589,I412578,);
nor I_24149 (I413067,I688349,I688331);
or I_24150 (I412569,I412816,I413067);
nor I_24151 (I412560,I412949,I413067);
or I_24152 (I412563,I412683,I413067);
DFFARX1 I_24153 (I413067,I2507,I412589,I412581,);
not I_24154 (I413167,I2514);
DFFARX1 I_24155 (I227009,I2507,I413167,I413193,);
not I_24156 (I413201,I413193);
nand I_24157 (I413218,I227012,I226988);
and I_24158 (I413235,I413218,I226985);
DFFARX1 I_24159 (I413235,I2507,I413167,I413261,);
not I_24160 (I413269,I226991);
DFFARX1 I_24161 (I226985,I2507,I413167,I413295,);
not I_24162 (I413303,I413295);
nor I_24163 (I413320,I413303,I413201);
and I_24164 (I413337,I413320,I226991);
nor I_24165 (I413354,I413303,I413269);
nor I_24166 (I413150,I413261,I413354);
DFFARX1 I_24167 (I226994,I2507,I413167,I413394,);
nor I_24168 (I413402,I413394,I413261);
not I_24169 (I413419,I413402);
not I_24170 (I413436,I413394);
nor I_24171 (I413453,I413436,I413337);
DFFARX1 I_24172 (I413453,I2507,I413167,I413153,);
nand I_24173 (I413484,I226997,I227006);
and I_24174 (I413501,I413484,I227003);
DFFARX1 I_24175 (I413501,I2507,I413167,I413527,);
nor I_24176 (I413535,I413527,I413394);
DFFARX1 I_24177 (I413535,I2507,I413167,I413135,);
nand I_24178 (I413566,I413527,I413436);
nand I_24179 (I413144,I413419,I413566);
not I_24180 (I413597,I413527);
nor I_24181 (I413614,I413597,I413337);
DFFARX1 I_24182 (I413614,I2507,I413167,I413156,);
nor I_24183 (I413645,I227000,I227006);
or I_24184 (I413147,I413394,I413645);
nor I_24185 (I413138,I413527,I413645);
or I_24186 (I413141,I413261,I413645);
DFFARX1 I_24187 (I413645,I2507,I413167,I413159,);
not I_24188 (I413745,I2514);
DFFARX1 I_24189 (I482196,I2507,I413745,I413771,);
not I_24190 (I413779,I413771);
nand I_24191 (I413796,I482172,I482187);
and I_24192 (I413813,I413796,I482199);
DFFARX1 I_24193 (I413813,I2507,I413745,I413839,);
not I_24194 (I413847,I482184);
DFFARX1 I_24195 (I482175,I2507,I413745,I413873,);
not I_24196 (I413881,I413873);
nor I_24197 (I413898,I413881,I413779);
and I_24198 (I413915,I413898,I482184);
nor I_24199 (I413932,I413881,I413847);
nor I_24200 (I413728,I413839,I413932);
DFFARX1 I_24201 (I482172,I2507,I413745,I413972,);
nor I_24202 (I413980,I413972,I413839);
not I_24203 (I413997,I413980);
not I_24204 (I414014,I413972);
nor I_24205 (I414031,I414014,I413915);
DFFARX1 I_24206 (I414031,I2507,I413745,I413731,);
nand I_24207 (I414062,I482190,I482181);
and I_24208 (I414079,I414062,I482193);
DFFARX1 I_24209 (I414079,I2507,I413745,I414105,);
nor I_24210 (I414113,I414105,I413972);
DFFARX1 I_24211 (I414113,I2507,I413745,I413713,);
nand I_24212 (I414144,I414105,I414014);
nand I_24213 (I413722,I413997,I414144);
not I_24214 (I414175,I414105);
nor I_24215 (I414192,I414175,I413915);
DFFARX1 I_24216 (I414192,I2507,I413745,I413734,);
nor I_24217 (I414223,I482178,I482181);
or I_24218 (I413725,I413972,I414223);
nor I_24219 (I413716,I414105,I414223);
or I_24220 (I413719,I413839,I414223);
DFFARX1 I_24221 (I414223,I2507,I413745,I413737,);
not I_24222 (I414323,I2514);
DFFARX1 I_24223 (I623715,I2507,I414323,I414349,);
not I_24224 (I414357,I414349);
nand I_24225 (I414374,I623697,I623709);
and I_24226 (I414391,I414374,I623712);
DFFARX1 I_24227 (I414391,I2507,I414323,I414417,);
not I_24228 (I414425,I623706);
DFFARX1 I_24229 (I623703,I2507,I414323,I414451,);
not I_24230 (I414459,I414451);
nor I_24231 (I414476,I414459,I414357);
and I_24232 (I414493,I414476,I623706);
nor I_24233 (I414510,I414459,I414425);
nor I_24234 (I414306,I414417,I414510);
DFFARX1 I_24235 (I623721,I2507,I414323,I414550,);
nor I_24236 (I414558,I414550,I414417);
not I_24237 (I414575,I414558);
not I_24238 (I414592,I414550);
nor I_24239 (I414609,I414592,I414493);
DFFARX1 I_24240 (I414609,I2507,I414323,I414309,);
nand I_24241 (I414640,I623700,I623700);
and I_24242 (I414657,I414640,I623697);
DFFARX1 I_24243 (I414657,I2507,I414323,I414683,);
nor I_24244 (I414691,I414683,I414550);
DFFARX1 I_24245 (I414691,I2507,I414323,I414291,);
nand I_24246 (I414722,I414683,I414592);
nand I_24247 (I414300,I414575,I414722);
not I_24248 (I414753,I414683);
nor I_24249 (I414770,I414753,I414493);
DFFARX1 I_24250 (I414770,I2507,I414323,I414312,);
nor I_24251 (I414801,I623718,I623700);
or I_24252 (I414303,I414550,I414801);
nor I_24253 (I414294,I414683,I414801);
or I_24254 (I414297,I414417,I414801);
DFFARX1 I_24255 (I414801,I2507,I414323,I414315,);
not I_24256 (I414901,I2514);
DFFARX1 I_24257 (I70979,I2507,I414901,I414927,);
not I_24258 (I414935,I414927);
nand I_24259 (I414952,I70988,I70997);
and I_24260 (I414969,I414952,I70976);
DFFARX1 I_24261 (I414969,I2507,I414901,I414995,);
not I_24262 (I415003,I70979);
DFFARX1 I_24263 (I70994,I2507,I414901,I415029,);
not I_24264 (I415037,I415029);
nor I_24265 (I415054,I415037,I414935);
and I_24266 (I415071,I415054,I70979);
nor I_24267 (I415088,I415037,I415003);
nor I_24268 (I414884,I414995,I415088);
DFFARX1 I_24269 (I70985,I2507,I414901,I415128,);
nor I_24270 (I415136,I415128,I414995);
not I_24271 (I415153,I415136);
not I_24272 (I415170,I415128);
nor I_24273 (I415187,I415170,I415071);
DFFARX1 I_24274 (I415187,I2507,I414901,I414887,);
nand I_24275 (I415218,I71000,I70976);
and I_24276 (I415235,I415218,I70982);
DFFARX1 I_24277 (I415235,I2507,I414901,I415261,);
nor I_24278 (I415269,I415261,I415128);
DFFARX1 I_24279 (I415269,I2507,I414901,I414869,);
nand I_24280 (I415300,I415261,I415170);
nand I_24281 (I414878,I415153,I415300);
not I_24282 (I415331,I415261);
nor I_24283 (I415348,I415331,I415071);
DFFARX1 I_24284 (I415348,I2507,I414901,I414890,);
nor I_24285 (I415379,I70991,I70976);
or I_24286 (I414881,I415128,I415379);
nor I_24287 (I414872,I415261,I415379);
or I_24288 (I414875,I414995,I415379);
DFFARX1 I_24289 (I415379,I2507,I414901,I414893,);
not I_24290 (I415479,I2514);
DFFARX1 I_24291 (I449207,I2507,I415479,I415505,);
not I_24292 (I415513,I415505);
nand I_24293 (I415530,I449195,I449213);
and I_24294 (I415547,I415530,I449210);
DFFARX1 I_24295 (I415547,I2507,I415479,I415573,);
not I_24296 (I415581,I449201);
DFFARX1 I_24297 (I449198,I2507,I415479,I415607,);
not I_24298 (I415615,I415607);
nor I_24299 (I415632,I415615,I415513);
and I_24300 (I415649,I415632,I449201);
nor I_24301 (I415666,I415615,I415581);
nor I_24302 (I415462,I415573,I415666);
DFFARX1 I_24303 (I449192,I2507,I415479,I415706,);
nor I_24304 (I415714,I415706,I415573);
not I_24305 (I415731,I415714);
not I_24306 (I415748,I415706);
nor I_24307 (I415765,I415748,I415649);
DFFARX1 I_24308 (I415765,I2507,I415479,I415465,);
nand I_24309 (I415796,I449192,I449195);
and I_24310 (I415813,I415796,I449198);
DFFARX1 I_24311 (I415813,I2507,I415479,I415839,);
nor I_24312 (I415847,I415839,I415706);
DFFARX1 I_24313 (I415847,I2507,I415479,I415447,);
nand I_24314 (I415878,I415839,I415748);
nand I_24315 (I415456,I415731,I415878);
not I_24316 (I415909,I415839);
nor I_24317 (I415926,I415909,I415649);
DFFARX1 I_24318 (I415926,I2507,I415479,I415468,);
nor I_24319 (I415957,I449204,I449195);
or I_24320 (I415459,I415706,I415957);
nor I_24321 (I415450,I415839,I415957);
or I_24322 (I415453,I415573,I415957);
DFFARX1 I_24323 (I415957,I2507,I415479,I415471,);
not I_24324 (I416057,I2514);
DFFARX1 I_24325 (I556502,I2507,I416057,I416083,);
not I_24326 (I416091,I416083);
nand I_24327 (I416108,I556499,I556517);
and I_24328 (I416125,I416108,I556514);
DFFARX1 I_24329 (I416125,I2507,I416057,I416151,);
not I_24330 (I416159,I556496);
DFFARX1 I_24331 (I556499,I2507,I416057,I416185,);
not I_24332 (I416193,I416185);
nor I_24333 (I416210,I416193,I416091);
and I_24334 (I416227,I416210,I556496);
nor I_24335 (I416244,I416193,I416159);
nor I_24336 (I416040,I416151,I416244);
DFFARX1 I_24337 (I556508,I2507,I416057,I416284,);
nor I_24338 (I416292,I416284,I416151);
not I_24339 (I416309,I416292);
not I_24340 (I416326,I416284);
nor I_24341 (I416343,I416326,I416227);
DFFARX1 I_24342 (I416343,I2507,I416057,I416043,);
nand I_24343 (I416374,I556511,I556496);
and I_24344 (I416391,I416374,I556502);
DFFARX1 I_24345 (I416391,I2507,I416057,I416417,);
nor I_24346 (I416425,I416417,I416284);
DFFARX1 I_24347 (I416425,I2507,I416057,I416025,);
nand I_24348 (I416456,I416417,I416326);
nand I_24349 (I416034,I416309,I416456);
not I_24350 (I416487,I416417);
nor I_24351 (I416504,I416487,I416227);
DFFARX1 I_24352 (I416504,I2507,I416057,I416046,);
nor I_24353 (I416535,I556505,I556496);
or I_24354 (I416037,I416284,I416535);
nor I_24355 (I416028,I416417,I416535);
or I_24356 (I416031,I416151,I416535);
DFFARX1 I_24357 (I416535,I2507,I416057,I416049,);
not I_24358 (I416635,I2514);
DFFARX1 I_24359 (I290888,I2507,I416635,I416661,);
not I_24360 (I416669,I416661);
nand I_24361 (I416686,I290903,I290888);
and I_24362 (I416703,I416686,I290891);
DFFARX1 I_24363 (I416703,I2507,I416635,I416729,);
not I_24364 (I416737,I290891);
DFFARX1 I_24365 (I290900,I2507,I416635,I416763,);
not I_24366 (I416771,I416763);
nor I_24367 (I416788,I416771,I416669);
and I_24368 (I416805,I416788,I290891);
nor I_24369 (I416822,I416771,I416737);
nor I_24370 (I416618,I416729,I416822);
DFFARX1 I_24371 (I290894,I2507,I416635,I416862,);
nor I_24372 (I416870,I416862,I416729);
not I_24373 (I416887,I416870);
not I_24374 (I416904,I416862);
nor I_24375 (I416921,I416904,I416805);
DFFARX1 I_24376 (I416921,I2507,I416635,I416621,);
nand I_24377 (I416952,I290897,I290906);
and I_24378 (I416969,I416952,I290912);
DFFARX1 I_24379 (I416969,I2507,I416635,I416995,);
nor I_24380 (I417003,I416995,I416862);
DFFARX1 I_24381 (I417003,I2507,I416635,I416603,);
nand I_24382 (I417034,I416995,I416904);
nand I_24383 (I416612,I416887,I417034);
not I_24384 (I417065,I416995);
nor I_24385 (I417082,I417065,I416805);
DFFARX1 I_24386 (I417082,I2507,I416635,I416624,);
nor I_24387 (I417113,I290909,I290906);
or I_24388 (I416615,I416862,I417113);
nor I_24389 (I416606,I416995,I417113);
or I_24390 (I416609,I416729,I417113);
DFFARX1 I_24391 (I417113,I2507,I416635,I416627,);
not I_24392 (I417213,I2514);
DFFARX1 I_24393 (I184849,I2507,I417213,I417239,);
not I_24394 (I417247,I417239);
nand I_24395 (I417264,I184852,I184828);
and I_24396 (I417281,I417264,I184825);
DFFARX1 I_24397 (I417281,I2507,I417213,I417307,);
not I_24398 (I417315,I184831);
DFFARX1 I_24399 (I184825,I2507,I417213,I417341,);
not I_24400 (I417349,I417341);
nor I_24401 (I417366,I417349,I417247);
and I_24402 (I417383,I417366,I184831);
nor I_24403 (I417400,I417349,I417315);
nor I_24404 (I417196,I417307,I417400);
DFFARX1 I_24405 (I184834,I2507,I417213,I417440,);
nor I_24406 (I417448,I417440,I417307);
not I_24407 (I417465,I417448);
not I_24408 (I417482,I417440);
nor I_24409 (I417499,I417482,I417383);
DFFARX1 I_24410 (I417499,I2507,I417213,I417199,);
nand I_24411 (I417530,I184837,I184846);
and I_24412 (I417547,I417530,I184843);
DFFARX1 I_24413 (I417547,I2507,I417213,I417573,);
nor I_24414 (I417581,I417573,I417440);
DFFARX1 I_24415 (I417581,I2507,I417213,I417181,);
nand I_24416 (I417612,I417573,I417482);
nand I_24417 (I417190,I417465,I417612);
not I_24418 (I417643,I417573);
nor I_24419 (I417660,I417643,I417383);
DFFARX1 I_24420 (I417660,I2507,I417213,I417202,);
nor I_24421 (I417691,I184840,I184846);
or I_24422 (I417193,I417440,I417691);
nor I_24423 (I417184,I417573,I417691);
or I_24424 (I417187,I417307,I417691);
DFFARX1 I_24425 (I417691,I2507,I417213,I417205,);
not I_24426 (I417791,I2514);
DFFARX1 I_24427 (I550892,I2507,I417791,I417817,);
not I_24428 (I417825,I417817);
nand I_24429 (I417842,I550889,I550907);
and I_24430 (I417859,I417842,I550904);
DFFARX1 I_24431 (I417859,I2507,I417791,I417885,);
not I_24432 (I417893,I550886);
DFFARX1 I_24433 (I550889,I2507,I417791,I417919,);
not I_24434 (I417927,I417919);
nor I_24435 (I417944,I417927,I417825);
and I_24436 (I417961,I417944,I550886);
nor I_24437 (I417978,I417927,I417893);
nor I_24438 (I417774,I417885,I417978);
DFFARX1 I_24439 (I550898,I2507,I417791,I418018,);
nor I_24440 (I418026,I418018,I417885);
not I_24441 (I418043,I418026);
not I_24442 (I418060,I418018);
nor I_24443 (I418077,I418060,I417961);
DFFARX1 I_24444 (I418077,I2507,I417791,I417777,);
nand I_24445 (I418108,I550901,I550886);
and I_24446 (I418125,I418108,I550892);
DFFARX1 I_24447 (I418125,I2507,I417791,I418151,);
nor I_24448 (I418159,I418151,I418018);
DFFARX1 I_24449 (I418159,I2507,I417791,I417759,);
nand I_24450 (I418190,I418151,I418060);
nand I_24451 (I417768,I418043,I418190);
not I_24452 (I418221,I418151);
nor I_24453 (I418238,I418221,I417961);
DFFARX1 I_24454 (I418238,I2507,I417791,I417780,);
nor I_24455 (I418269,I550895,I550886);
or I_24456 (I417771,I418018,I418269);
nor I_24457 (I417762,I418151,I418269);
or I_24458 (I417765,I417885,I418269);
DFFARX1 I_24459 (I418269,I2507,I417791,I417783,);
not I_24460 (I418369,I2514);
DFFARX1 I_24461 (I523540,I2507,I418369,I418395,);
not I_24462 (I418403,I418395);
nand I_24463 (I418420,I523516,I523531);
and I_24464 (I418437,I418420,I523543);
DFFARX1 I_24465 (I418437,I2507,I418369,I418463,);
not I_24466 (I418471,I523528);
DFFARX1 I_24467 (I523519,I2507,I418369,I418497,);
not I_24468 (I418505,I418497);
nor I_24469 (I418522,I418505,I418403);
and I_24470 (I418539,I418522,I523528);
nor I_24471 (I418556,I418505,I418471);
nor I_24472 (I418352,I418463,I418556);
DFFARX1 I_24473 (I523516,I2507,I418369,I418596,);
nor I_24474 (I418604,I418596,I418463);
not I_24475 (I418621,I418604);
not I_24476 (I418638,I418596);
nor I_24477 (I418655,I418638,I418539);
DFFARX1 I_24478 (I418655,I2507,I418369,I418355,);
nand I_24479 (I418686,I523534,I523525);
and I_24480 (I418703,I418686,I523537);
DFFARX1 I_24481 (I418703,I2507,I418369,I418729,);
nor I_24482 (I418737,I418729,I418596);
DFFARX1 I_24483 (I418737,I2507,I418369,I418337,);
nand I_24484 (I418768,I418729,I418638);
nand I_24485 (I418346,I418621,I418768);
not I_24486 (I418799,I418729);
nor I_24487 (I418816,I418799,I418539);
DFFARX1 I_24488 (I418816,I2507,I418369,I418358,);
nor I_24489 (I418847,I523522,I523525);
or I_24490 (I418349,I418596,I418847);
nor I_24491 (I418340,I418729,I418847);
or I_24492 (I418343,I418463,I418847);
DFFARX1 I_24493 (I418847,I2507,I418369,I418361,);
not I_24494 (I418947,I2514);
DFFARX1 I_24495 (I455004,I2507,I418947,I418973,);
not I_24496 (I418981,I418973);
nand I_24497 (I418998,I454992,I455010);
and I_24498 (I419015,I418998,I455007);
DFFARX1 I_24499 (I419015,I2507,I418947,I419041,);
not I_24500 (I419049,I454998);
DFFARX1 I_24501 (I454995,I2507,I418947,I419075,);
not I_24502 (I419083,I419075);
nor I_24503 (I419100,I419083,I418981);
and I_24504 (I419117,I419100,I454998);
nor I_24505 (I419134,I419083,I419049);
nor I_24506 (I418930,I419041,I419134);
DFFARX1 I_24507 (I454989,I2507,I418947,I419174,);
nor I_24508 (I419182,I419174,I419041);
not I_24509 (I419199,I419182);
not I_24510 (I419216,I419174);
nor I_24511 (I419233,I419216,I419117);
DFFARX1 I_24512 (I419233,I2507,I418947,I418933,);
nand I_24513 (I419264,I454989,I454992);
and I_24514 (I419281,I419264,I454995);
DFFARX1 I_24515 (I419281,I2507,I418947,I419307,);
nor I_24516 (I419315,I419307,I419174);
DFFARX1 I_24517 (I419315,I2507,I418947,I418915,);
nand I_24518 (I419346,I419307,I419216);
nand I_24519 (I418924,I419199,I419346);
not I_24520 (I419377,I419307);
nor I_24521 (I419394,I419377,I419117);
DFFARX1 I_24522 (I419394,I2507,I418947,I418936,);
nor I_24523 (I419425,I455001,I454992);
or I_24524 (I418927,I419174,I419425);
nor I_24525 (I418918,I419307,I419425);
or I_24526 (I418921,I419041,I419425);
DFFARX1 I_24527 (I419425,I2507,I418947,I418939,);
not I_24528 (I419525,I2514);
DFFARX1 I_24529 (I37251,I2507,I419525,I419551,);
not I_24530 (I419559,I419551);
nand I_24531 (I419576,I37260,I37269);
and I_24532 (I419593,I419576,I37248);
DFFARX1 I_24533 (I419593,I2507,I419525,I419619,);
not I_24534 (I419627,I37251);
DFFARX1 I_24535 (I37266,I2507,I419525,I419653,);
not I_24536 (I419661,I419653);
nor I_24537 (I419678,I419661,I419559);
and I_24538 (I419695,I419678,I37251);
nor I_24539 (I419712,I419661,I419627);
nor I_24540 (I419508,I419619,I419712);
DFFARX1 I_24541 (I37257,I2507,I419525,I419752,);
nor I_24542 (I419760,I419752,I419619);
not I_24543 (I419777,I419760);
not I_24544 (I419794,I419752);
nor I_24545 (I419811,I419794,I419695);
DFFARX1 I_24546 (I419811,I2507,I419525,I419511,);
nand I_24547 (I419842,I37272,I37248);
and I_24548 (I419859,I419842,I37254);
DFFARX1 I_24549 (I419859,I2507,I419525,I419885,);
nor I_24550 (I419893,I419885,I419752);
DFFARX1 I_24551 (I419893,I2507,I419525,I419493,);
nand I_24552 (I419924,I419885,I419794);
nand I_24553 (I419502,I419777,I419924);
not I_24554 (I419955,I419885);
nor I_24555 (I419972,I419955,I419695);
DFFARX1 I_24556 (I419972,I2507,I419525,I419514,);
nor I_24557 (I420003,I37263,I37248);
or I_24558 (I419505,I419752,I420003);
nor I_24559 (I419496,I419885,I420003);
or I_24560 (I419499,I419619,I420003);
DFFARX1 I_24561 (I420003,I2507,I419525,I419517,);
not I_24562 (I420103,I2514);
DFFARX1 I_24563 (I513204,I2507,I420103,I420129,);
not I_24564 (I420137,I420129);
nand I_24565 (I420154,I513180,I513195);
and I_24566 (I420171,I420154,I513207);
DFFARX1 I_24567 (I420171,I2507,I420103,I420197,);
not I_24568 (I420205,I513192);
DFFARX1 I_24569 (I513183,I2507,I420103,I420231,);
not I_24570 (I420239,I420231);
nor I_24571 (I420256,I420239,I420137);
and I_24572 (I420273,I420256,I513192);
nor I_24573 (I420290,I420239,I420205);
nor I_24574 (I420086,I420197,I420290);
DFFARX1 I_24575 (I513180,I2507,I420103,I420330,);
nor I_24576 (I420338,I420330,I420197);
not I_24577 (I420355,I420338);
not I_24578 (I420372,I420330);
nor I_24579 (I420389,I420372,I420273);
DFFARX1 I_24580 (I420389,I2507,I420103,I420089,);
nand I_24581 (I420420,I513198,I513189);
and I_24582 (I420437,I420420,I513201);
DFFARX1 I_24583 (I420437,I2507,I420103,I420463,);
nor I_24584 (I420471,I420463,I420330);
DFFARX1 I_24585 (I420471,I2507,I420103,I420071,);
nand I_24586 (I420502,I420463,I420372);
nand I_24587 (I420080,I420355,I420502);
not I_24588 (I420533,I420463);
nor I_24589 (I420550,I420533,I420273);
DFFARX1 I_24590 (I420550,I2507,I420103,I420092,);
nor I_24591 (I420581,I513186,I513189);
or I_24592 (I420083,I420330,I420581);
nor I_24593 (I420074,I420463,I420581);
or I_24594 (I420077,I420197,I420581);
DFFARX1 I_24595 (I420581,I2507,I420103,I420095,);
not I_24596 (I420681,I2514);
DFFARX1 I_24597 (I248193,I2507,I420681,I420707,);
not I_24598 (I420715,I420707);
nand I_24599 (I420732,I248184,I248202);
and I_24600 (I420749,I420732,I248205);
DFFARX1 I_24601 (I420749,I2507,I420681,I420775,);
not I_24602 (I420783,I248199);
DFFARX1 I_24603 (I248187,I2507,I420681,I420809,);
not I_24604 (I420817,I420809);
nor I_24605 (I420834,I420817,I420715);
and I_24606 (I420851,I420834,I248199);
nor I_24607 (I420868,I420817,I420783);
nor I_24608 (I420664,I420775,I420868);
DFFARX1 I_24609 (I248196,I2507,I420681,I420908,);
nor I_24610 (I420916,I420908,I420775);
not I_24611 (I420933,I420916);
not I_24612 (I420950,I420908);
nor I_24613 (I420967,I420950,I420851);
DFFARX1 I_24614 (I420967,I2507,I420681,I420667,);
nand I_24615 (I420998,I248211,I248208);
and I_24616 (I421015,I420998,I248190);
DFFARX1 I_24617 (I421015,I2507,I420681,I421041,);
nor I_24618 (I421049,I421041,I420908);
DFFARX1 I_24619 (I421049,I2507,I420681,I420649,);
nand I_24620 (I421080,I421041,I420950);
nand I_24621 (I420658,I420933,I421080);
not I_24622 (I421111,I421041);
nor I_24623 (I421128,I421111,I420851);
DFFARX1 I_24624 (I421128,I2507,I420681,I420670,);
nor I_24625 (I421159,I248184,I248208);
or I_24626 (I420661,I420908,I421159);
nor I_24627 (I420652,I421041,I421159);
or I_24628 (I420655,I420775,I421159);
DFFARX1 I_24629 (I421159,I2507,I420681,I420673,);
not I_24630 (I421259,I2514);
DFFARX1 I_24631 (I632385,I2507,I421259,I421285,);
not I_24632 (I421293,I421285);
nand I_24633 (I421310,I632367,I632379);
and I_24634 (I421327,I421310,I632382);
DFFARX1 I_24635 (I421327,I2507,I421259,I421353,);
not I_24636 (I421361,I632376);
DFFARX1 I_24637 (I632373,I2507,I421259,I421387,);
not I_24638 (I421395,I421387);
nor I_24639 (I421412,I421395,I421293);
and I_24640 (I421429,I421412,I632376);
nor I_24641 (I421446,I421395,I421361);
nor I_24642 (I421242,I421353,I421446);
DFFARX1 I_24643 (I632391,I2507,I421259,I421486,);
nor I_24644 (I421494,I421486,I421353);
not I_24645 (I421511,I421494);
not I_24646 (I421528,I421486);
nor I_24647 (I421545,I421528,I421429);
DFFARX1 I_24648 (I421545,I2507,I421259,I421245,);
nand I_24649 (I421576,I632370,I632370);
and I_24650 (I421593,I421576,I632367);
DFFARX1 I_24651 (I421593,I2507,I421259,I421619,);
nor I_24652 (I421627,I421619,I421486);
DFFARX1 I_24653 (I421627,I2507,I421259,I421227,);
nand I_24654 (I421658,I421619,I421528);
nand I_24655 (I421236,I421511,I421658);
not I_24656 (I421689,I421619);
nor I_24657 (I421706,I421689,I421429);
DFFARX1 I_24658 (I421706,I2507,I421259,I421248,);
nor I_24659 (I421737,I632388,I632370);
or I_24660 (I421239,I421486,I421737);
nor I_24661 (I421230,I421619,I421737);
or I_24662 (I421233,I421353,I421737);
DFFARX1 I_24663 (I421737,I2507,I421259,I421251,);
not I_24664 (I421837,I2514);
DFFARX1 I_24665 (I664293,I2507,I421837,I421863,);
not I_24666 (I421871,I421863);
nand I_24667 (I421888,I664296,I664305);
and I_24668 (I421905,I421888,I664308);
DFFARX1 I_24669 (I421905,I2507,I421837,I421931,);
not I_24670 (I421939,I664317);
DFFARX1 I_24671 (I664299,I2507,I421837,I421965,);
not I_24672 (I421973,I421965);
nor I_24673 (I421990,I421973,I421871);
and I_24674 (I422007,I421990,I664317);
nor I_24675 (I422024,I421973,I421939);
nor I_24676 (I421820,I421931,I422024);
DFFARX1 I_24677 (I664296,I2507,I421837,I422064,);
nor I_24678 (I422072,I422064,I421931);
not I_24679 (I422089,I422072);
not I_24680 (I422106,I422064);
nor I_24681 (I422123,I422106,I422007);
DFFARX1 I_24682 (I422123,I2507,I421837,I421823,);
nand I_24683 (I422154,I664314,I664293);
and I_24684 (I422171,I422154,I664311);
DFFARX1 I_24685 (I422171,I2507,I421837,I422197,);
nor I_24686 (I422205,I422197,I422064);
DFFARX1 I_24687 (I422205,I2507,I421837,I421805,);
nand I_24688 (I422236,I422197,I422106);
nand I_24689 (I421814,I422089,I422236);
not I_24690 (I422267,I422197);
nor I_24691 (I422284,I422267,I422007);
DFFARX1 I_24692 (I422284,I2507,I421837,I421826,);
nor I_24693 (I422315,I664302,I664293);
or I_24694 (I421817,I422064,I422315);
nor I_24695 (I421808,I422197,I422315);
or I_24696 (I421811,I421931,I422315);
DFFARX1 I_24697 (I422315,I2507,I421837,I421829,);
not I_24698 (I422415,I2514);
DFFARX1 I_24699 (I604063,I2507,I422415,I422441,);
not I_24700 (I422449,I422441);
nand I_24701 (I422466,I604045,I604057);
and I_24702 (I422483,I422466,I604060);
DFFARX1 I_24703 (I422483,I2507,I422415,I422509,);
not I_24704 (I422517,I604054);
DFFARX1 I_24705 (I604051,I2507,I422415,I422543,);
not I_24706 (I422551,I422543);
nor I_24707 (I422568,I422551,I422449);
and I_24708 (I422585,I422568,I604054);
nor I_24709 (I422602,I422551,I422517);
nor I_24710 (I422398,I422509,I422602);
DFFARX1 I_24711 (I604069,I2507,I422415,I422642,);
nor I_24712 (I422650,I422642,I422509);
not I_24713 (I422667,I422650);
not I_24714 (I422684,I422642);
nor I_24715 (I422701,I422684,I422585);
DFFARX1 I_24716 (I422701,I2507,I422415,I422401,);
nand I_24717 (I422732,I604048,I604048);
and I_24718 (I422749,I422732,I604045);
DFFARX1 I_24719 (I422749,I2507,I422415,I422775,);
nor I_24720 (I422783,I422775,I422642);
DFFARX1 I_24721 (I422783,I2507,I422415,I422383,);
nand I_24722 (I422814,I422775,I422684);
nand I_24723 (I422392,I422667,I422814);
not I_24724 (I422845,I422775);
nor I_24725 (I422862,I422845,I422585);
DFFARX1 I_24726 (I422862,I2507,I422415,I422404,);
nor I_24727 (I422893,I604066,I604048);
or I_24728 (I422395,I422642,I422893);
nor I_24729 (I422386,I422775,I422893);
or I_24730 (I422389,I422509,I422893);
DFFARX1 I_24731 (I422893,I2507,I422415,I422407,);
not I_24732 (I422993,I2514);
DFFARX1 I_24733 (I195916,I2507,I422993,I423019,);
not I_24734 (I423027,I423019);
nand I_24735 (I423044,I195919,I195895);
and I_24736 (I423061,I423044,I195892);
DFFARX1 I_24737 (I423061,I2507,I422993,I423087,);
not I_24738 (I423095,I195898);
DFFARX1 I_24739 (I195892,I2507,I422993,I423121,);
not I_24740 (I423129,I423121);
nor I_24741 (I423146,I423129,I423027);
and I_24742 (I423163,I423146,I195898);
nor I_24743 (I423180,I423129,I423095);
nor I_24744 (I422976,I423087,I423180);
DFFARX1 I_24745 (I195901,I2507,I422993,I423220,);
nor I_24746 (I423228,I423220,I423087);
not I_24747 (I423245,I423228);
not I_24748 (I423262,I423220);
nor I_24749 (I423279,I423262,I423163);
DFFARX1 I_24750 (I423279,I2507,I422993,I422979,);
nand I_24751 (I423310,I195904,I195913);
and I_24752 (I423327,I423310,I195910);
DFFARX1 I_24753 (I423327,I2507,I422993,I423353,);
nor I_24754 (I423361,I423353,I423220);
DFFARX1 I_24755 (I423361,I2507,I422993,I422961,);
nand I_24756 (I423392,I423353,I423262);
nand I_24757 (I422970,I423245,I423392);
not I_24758 (I423423,I423353);
nor I_24759 (I423440,I423423,I423163);
DFFARX1 I_24760 (I423440,I2507,I422993,I422982,);
nor I_24761 (I423471,I195907,I195913);
or I_24762 (I422973,I423220,I423471);
nor I_24763 (I422964,I423353,I423471);
or I_24764 (I422967,I423087,I423471);
DFFARX1 I_24765 (I423471,I2507,I422993,I422985,);
not I_24766 (I423571,I2514);
DFFARX1 I_24767 (I542477,I2507,I423571,I423597,);
not I_24768 (I423605,I423597);
nand I_24769 (I423622,I542474,I542492);
and I_24770 (I423639,I423622,I542489);
DFFARX1 I_24771 (I423639,I2507,I423571,I423665,);
not I_24772 (I423673,I542471);
DFFARX1 I_24773 (I542474,I2507,I423571,I423699,);
not I_24774 (I423707,I423699);
nor I_24775 (I423724,I423707,I423605);
and I_24776 (I423741,I423724,I542471);
nor I_24777 (I423758,I423707,I423673);
nor I_24778 (I423554,I423665,I423758);
DFFARX1 I_24779 (I542483,I2507,I423571,I423798,);
nor I_24780 (I423806,I423798,I423665);
not I_24781 (I423823,I423806);
not I_24782 (I423840,I423798);
nor I_24783 (I423857,I423840,I423741);
DFFARX1 I_24784 (I423857,I2507,I423571,I423557,);
nand I_24785 (I423888,I542486,I542471);
and I_24786 (I423905,I423888,I542477);
DFFARX1 I_24787 (I423905,I2507,I423571,I423931,);
nor I_24788 (I423939,I423931,I423798);
DFFARX1 I_24789 (I423939,I2507,I423571,I423539,);
nand I_24790 (I423970,I423931,I423840);
nand I_24791 (I423548,I423823,I423970);
not I_24792 (I424001,I423931);
nor I_24793 (I424018,I424001,I423741);
DFFARX1 I_24794 (I424018,I2507,I423571,I423560,);
nor I_24795 (I424049,I542480,I542471);
or I_24796 (I423551,I423798,I424049);
nor I_24797 (I423542,I423931,I424049);
or I_24798 (I423545,I423665,I424049);
DFFARX1 I_24799 (I424049,I2507,I423571,I423563,);
not I_24800 (I424149,I2514);
DFFARX1 I_24801 (I452896,I2507,I424149,I424175,);
not I_24802 (I424183,I424175);
nand I_24803 (I424200,I452884,I452902);
and I_24804 (I424217,I424200,I452899);
DFFARX1 I_24805 (I424217,I2507,I424149,I424243,);
not I_24806 (I424251,I452890);
DFFARX1 I_24807 (I452887,I2507,I424149,I424277,);
not I_24808 (I424285,I424277);
nor I_24809 (I424302,I424285,I424183);
and I_24810 (I424319,I424302,I452890);
nor I_24811 (I424336,I424285,I424251);
nor I_24812 (I424132,I424243,I424336);
DFFARX1 I_24813 (I452881,I2507,I424149,I424376,);
nor I_24814 (I424384,I424376,I424243);
not I_24815 (I424401,I424384);
not I_24816 (I424418,I424376);
nor I_24817 (I424435,I424418,I424319);
DFFARX1 I_24818 (I424435,I2507,I424149,I424135,);
nand I_24819 (I424466,I452881,I452884);
and I_24820 (I424483,I424466,I452887);
DFFARX1 I_24821 (I424483,I2507,I424149,I424509,);
nor I_24822 (I424517,I424509,I424376);
DFFARX1 I_24823 (I424517,I2507,I424149,I424117,);
nand I_24824 (I424548,I424509,I424418);
nand I_24825 (I424126,I424401,I424548);
not I_24826 (I424579,I424509);
nor I_24827 (I424596,I424579,I424319);
DFFARX1 I_24828 (I424596,I2507,I424149,I424138,);
nor I_24829 (I424627,I452893,I452884);
or I_24830 (I424129,I424376,I424627);
nor I_24831 (I424120,I424509,I424627);
or I_24832 (I424123,I424243,I424627);
DFFARX1 I_24833 (I424627,I2507,I424149,I424141,);
not I_24834 (I424727,I2514);
DFFARX1 I_24835 (I298623,I2507,I424727,I424753,);
not I_24836 (I424761,I424753);
nand I_24837 (I424778,I298638,I298623);
and I_24838 (I424795,I424778,I298626);
DFFARX1 I_24839 (I424795,I2507,I424727,I424821,);
not I_24840 (I424829,I298626);
DFFARX1 I_24841 (I298635,I2507,I424727,I424855,);
not I_24842 (I424863,I424855);
nor I_24843 (I424880,I424863,I424761);
and I_24844 (I424897,I424880,I298626);
nor I_24845 (I424914,I424863,I424829);
nor I_24846 (I424710,I424821,I424914);
DFFARX1 I_24847 (I298629,I2507,I424727,I424954,);
nor I_24848 (I424962,I424954,I424821);
not I_24849 (I424979,I424962);
not I_24850 (I424996,I424954);
nor I_24851 (I425013,I424996,I424897);
DFFARX1 I_24852 (I425013,I2507,I424727,I424713,);
nand I_24853 (I425044,I298632,I298641);
and I_24854 (I425061,I425044,I298647);
DFFARX1 I_24855 (I425061,I2507,I424727,I425087,);
nor I_24856 (I425095,I425087,I424954);
DFFARX1 I_24857 (I425095,I2507,I424727,I424695,);
nand I_24858 (I425126,I425087,I424996);
nand I_24859 (I424704,I424979,I425126);
not I_24860 (I425157,I425087);
nor I_24861 (I425174,I425157,I424897);
DFFARX1 I_24862 (I425174,I2507,I424727,I424716,);
nor I_24863 (I425205,I298644,I298641);
or I_24864 (I424707,I424954,I425205);
nor I_24865 (I424698,I425087,I425205);
or I_24866 (I424701,I424821,I425205);
DFFARX1 I_24867 (I425205,I2507,I424727,I424719,);
not I_24868 (I425305,I2514);
DFFARX1 I_24869 (I627761,I2507,I425305,I425331,);
not I_24870 (I425339,I425331);
nand I_24871 (I425356,I627743,I627755);
and I_24872 (I425373,I425356,I627758);
DFFARX1 I_24873 (I425373,I2507,I425305,I425399,);
not I_24874 (I425407,I627752);
DFFARX1 I_24875 (I627749,I2507,I425305,I425433,);
not I_24876 (I425441,I425433);
nor I_24877 (I425458,I425441,I425339);
and I_24878 (I425475,I425458,I627752);
nor I_24879 (I425492,I425441,I425407);
nor I_24880 (I425288,I425399,I425492);
DFFARX1 I_24881 (I627767,I2507,I425305,I425532,);
nor I_24882 (I425540,I425532,I425399);
not I_24883 (I425557,I425540);
not I_24884 (I425574,I425532);
nor I_24885 (I425591,I425574,I425475);
DFFARX1 I_24886 (I425591,I2507,I425305,I425291,);
nand I_24887 (I425622,I627746,I627746);
and I_24888 (I425639,I425622,I627743);
DFFARX1 I_24889 (I425639,I2507,I425305,I425665,);
nor I_24890 (I425673,I425665,I425532);
DFFARX1 I_24891 (I425673,I2507,I425305,I425273,);
nand I_24892 (I425704,I425665,I425574);
nand I_24893 (I425282,I425557,I425704);
not I_24894 (I425735,I425665);
nor I_24895 (I425752,I425735,I425475);
DFFARX1 I_24896 (I425752,I2507,I425305,I425294,);
nor I_24897 (I425783,I627764,I627746);
or I_24898 (I425285,I425532,I425783);
nor I_24899 (I425276,I425665,I425783);
or I_24900 (I425279,I425399,I425783);
DFFARX1 I_24901 (I425783,I2507,I425305,I425297,);
not I_24902 (I425883,I2514);
DFFARX1 I_24903 (I529354,I2507,I425883,I425909,);
not I_24904 (I425917,I425909);
nand I_24905 (I425934,I529330,I529345);
and I_24906 (I425951,I425934,I529357);
DFFARX1 I_24907 (I425951,I2507,I425883,I425977,);
not I_24908 (I425985,I529342);
DFFARX1 I_24909 (I529333,I2507,I425883,I426011,);
not I_24910 (I426019,I426011);
nor I_24911 (I426036,I426019,I425917);
and I_24912 (I426053,I426036,I529342);
nor I_24913 (I426070,I426019,I425985);
nor I_24914 (I425866,I425977,I426070);
DFFARX1 I_24915 (I529330,I2507,I425883,I426110,);
nor I_24916 (I426118,I426110,I425977);
not I_24917 (I426135,I426118);
not I_24918 (I426152,I426110);
nor I_24919 (I426169,I426152,I426053);
DFFARX1 I_24920 (I426169,I2507,I425883,I425869,);
nand I_24921 (I426200,I529348,I529339);
and I_24922 (I426217,I426200,I529351);
DFFARX1 I_24923 (I426217,I2507,I425883,I426243,);
nor I_24924 (I426251,I426243,I426110);
DFFARX1 I_24925 (I426251,I2507,I425883,I425851,);
nand I_24926 (I426282,I426243,I426152);
nand I_24927 (I425860,I426135,I426282);
not I_24928 (I426313,I426243);
nor I_24929 (I426330,I426313,I426053);
DFFARX1 I_24930 (I426330,I2507,I425883,I425872,);
nor I_24931 (I426361,I529336,I529339);
or I_24932 (I425863,I426110,I426361);
nor I_24933 (I425854,I426243,I426361);
or I_24934 (I425857,I425977,I426361);
DFFARX1 I_24935 (I426361,I2507,I425883,I425875,);
not I_24936 (I426461,I2514);
DFFARX1 I_24937 (I220158,I2507,I426461,I426487,);
not I_24938 (I426495,I426487);
nand I_24939 (I426512,I220161,I220137);
and I_24940 (I426529,I426512,I220134);
DFFARX1 I_24941 (I426529,I2507,I426461,I426555,);
not I_24942 (I426563,I220140);
DFFARX1 I_24943 (I220134,I2507,I426461,I426589,);
not I_24944 (I426597,I426589);
nor I_24945 (I426614,I426597,I426495);
and I_24946 (I426631,I426614,I220140);
nor I_24947 (I426648,I426597,I426563);
nor I_24948 (I426444,I426555,I426648);
DFFARX1 I_24949 (I220143,I2507,I426461,I426688,);
nor I_24950 (I426696,I426688,I426555);
not I_24951 (I426713,I426696);
not I_24952 (I426730,I426688);
nor I_24953 (I426747,I426730,I426631);
DFFARX1 I_24954 (I426747,I2507,I426461,I426447,);
nand I_24955 (I426778,I220146,I220155);
and I_24956 (I426795,I426778,I220152);
DFFARX1 I_24957 (I426795,I2507,I426461,I426821,);
nor I_24958 (I426829,I426821,I426688);
DFFARX1 I_24959 (I426829,I2507,I426461,I426429,);
nand I_24960 (I426860,I426821,I426730);
nand I_24961 (I426438,I426713,I426860);
not I_24962 (I426891,I426821);
nor I_24963 (I426908,I426891,I426631);
DFFARX1 I_24964 (I426908,I2507,I426461,I426450,);
nor I_24965 (I426939,I220149,I220155);
or I_24966 (I426441,I426688,I426939);
nor I_24967 (I426432,I426821,I426939);
or I_24968 (I426435,I426555,I426939);
DFFARX1 I_24969 (I426939,I2507,I426461,I426453,);
not I_24970 (I427039,I2514);
DFFARX1 I_24971 (I120514,I2507,I427039,I427065,);
not I_24972 (I427073,I427065);
nand I_24973 (I427090,I120517,I120538);
and I_24974 (I427107,I427090,I120526);
DFFARX1 I_24975 (I427107,I2507,I427039,I427133,);
not I_24976 (I427141,I120523);
DFFARX1 I_24977 (I120514,I2507,I427039,I427167,);
not I_24978 (I427175,I427167);
nor I_24979 (I427192,I427175,I427073);
and I_24980 (I427209,I427192,I120523);
nor I_24981 (I427226,I427175,I427141);
nor I_24982 (I427022,I427133,I427226);
DFFARX1 I_24983 (I120532,I2507,I427039,I427266,);
nor I_24984 (I427274,I427266,I427133);
not I_24985 (I427291,I427274);
not I_24986 (I427308,I427266);
nor I_24987 (I427325,I427308,I427209);
DFFARX1 I_24988 (I427325,I2507,I427039,I427025,);
nand I_24989 (I427356,I120517,I120520);
and I_24990 (I427373,I427356,I120529);
DFFARX1 I_24991 (I427373,I2507,I427039,I427399,);
nor I_24992 (I427407,I427399,I427266);
DFFARX1 I_24993 (I427407,I2507,I427039,I427007,);
nand I_24994 (I427438,I427399,I427308);
nand I_24995 (I427016,I427291,I427438);
not I_24996 (I427469,I427399);
nor I_24997 (I427486,I427469,I427209);
DFFARX1 I_24998 (I427486,I2507,I427039,I427028,);
nor I_24999 (I427517,I120535,I120520);
or I_25000 (I427019,I427266,I427517);
nor I_25001 (I427010,I427399,I427517);
or I_25002 (I427013,I427133,I427517);
DFFARX1 I_25003 (I427517,I2507,I427039,I427031,);
not I_25004 (I427614,I2514);
DFFARX1 I_25005 (I388281,I2507,I427614,I427640,);
not I_25006 (I427648,I427640);
nand I_25007 (I427665,I388284,I388281);
and I_25008 (I427682,I427665,I388293);
DFFARX1 I_25009 (I427682,I2507,I427614,I427708,);
DFFARX1 I_25010 (I427708,I2507,I427614,I427603,);
DFFARX1 I_25011 (I388290,I2507,I427614,I427739,);
nand I_25012 (I427747,I427739,I388296);
not I_25013 (I427764,I427747);
DFFARX1 I_25014 (I427764,I2507,I427614,I427790,);
not I_25015 (I427798,I427790);
nor I_25016 (I427606,I427648,I427798);
DFFARX1 I_25017 (I388305,I2507,I427614,I427838,);
nor I_25018 (I427597,I427838,I427708);
nor I_25019 (I427588,I427838,I427764);
nand I_25020 (I427874,I388299,I388287);
and I_25021 (I427891,I427874,I388284);
DFFARX1 I_25022 (I427891,I2507,I427614,I427917,);
not I_25023 (I427925,I427917);
nand I_25024 (I427942,I427925,I427838);
nand I_25025 (I427591,I427925,I427747);
nor I_25026 (I427973,I388302,I388287);
and I_25027 (I427990,I427838,I427973);
nor I_25028 (I428007,I427925,I427990);
DFFARX1 I_25029 (I428007,I2507,I427614,I427600,);
nor I_25030 (I428038,I427640,I427973);
DFFARX1 I_25031 (I428038,I2507,I427614,I427585,);
nor I_25032 (I428069,I427917,I427973);
not I_25033 (I428086,I428069);
nand I_25034 (I427594,I428086,I427942);
not I_25035 (I428141,I2514);
DFFARX1 I_25036 (I8799,I2507,I428141,I428167,);
not I_25037 (I428175,I428167);
nand I_25038 (I428192,I8811,I8814);
and I_25039 (I428209,I428192,I8790);
DFFARX1 I_25040 (I428209,I2507,I428141,I428235,);
DFFARX1 I_25041 (I428235,I2507,I428141,I428130,);
DFFARX1 I_25042 (I8808,I2507,I428141,I428266,);
nand I_25043 (I428274,I428266,I8796);
not I_25044 (I428291,I428274);
DFFARX1 I_25045 (I428291,I2507,I428141,I428317,);
not I_25046 (I428325,I428317);
nor I_25047 (I428133,I428175,I428325);
DFFARX1 I_25048 (I8793,I2507,I428141,I428365,);
nor I_25049 (I428124,I428365,I428235);
nor I_25050 (I428115,I428365,I428291);
nand I_25051 (I428401,I8802,I8793);
and I_25052 (I428418,I428401,I8790);
DFFARX1 I_25053 (I428418,I2507,I428141,I428444,);
not I_25054 (I428452,I428444);
nand I_25055 (I428469,I428452,I428365);
nand I_25056 (I428118,I428452,I428274);
nor I_25057 (I428500,I8805,I8793);
and I_25058 (I428517,I428365,I428500);
nor I_25059 (I428534,I428452,I428517);
DFFARX1 I_25060 (I428534,I2507,I428141,I428127,);
nor I_25061 (I428565,I428167,I428500);
DFFARX1 I_25062 (I428565,I2507,I428141,I428112,);
nor I_25063 (I428596,I428444,I428500);
not I_25064 (I428613,I428596);
nand I_25065 (I428121,I428613,I428469);
not I_25066 (I428668,I2514);
DFFARX1 I_25067 (I80486,I2507,I428668,I428694,);
not I_25068 (I428702,I428694);
nand I_25069 (I428719,I80462,I80471);
and I_25070 (I428736,I428719,I80465);
DFFARX1 I_25071 (I428736,I2507,I428668,I428762,);
DFFARX1 I_25072 (I428762,I2507,I428668,I428657,);
DFFARX1 I_25073 (I80483,I2507,I428668,I428793,);
nand I_25074 (I428801,I428793,I80474);
not I_25075 (I428818,I428801);
DFFARX1 I_25076 (I428818,I2507,I428668,I428844,);
not I_25077 (I428852,I428844);
nor I_25078 (I428660,I428702,I428852);
DFFARX1 I_25079 (I80468,I2507,I428668,I428892,);
nor I_25080 (I428651,I428892,I428762);
nor I_25081 (I428642,I428892,I428818);
nand I_25082 (I428928,I80480,I80477);
and I_25083 (I428945,I428928,I80465);
DFFARX1 I_25084 (I428945,I2507,I428668,I428971,);
not I_25085 (I428979,I428971);
nand I_25086 (I428996,I428979,I428892);
nand I_25087 (I428645,I428979,I428801);
nor I_25088 (I429027,I80462,I80477);
and I_25089 (I429044,I428892,I429027);
nor I_25090 (I429061,I428979,I429044);
DFFARX1 I_25091 (I429061,I2507,I428668,I428654,);
nor I_25092 (I429092,I428694,I429027);
DFFARX1 I_25093 (I429092,I2507,I428668,I428639,);
nor I_25094 (I429123,I428971,I429027);
not I_25095 (I429140,I429123);
nand I_25096 (I428648,I429140,I428996);
not I_25097 (I429195,I2514);
DFFARX1 I_25098 (I422961,I2507,I429195,I429221,);
not I_25099 (I429229,I429221);
nand I_25100 (I429246,I422964,I422961);
and I_25101 (I429263,I429246,I422973);
DFFARX1 I_25102 (I429263,I2507,I429195,I429289,);
DFFARX1 I_25103 (I429289,I2507,I429195,I429184,);
DFFARX1 I_25104 (I422970,I2507,I429195,I429320,);
nand I_25105 (I429328,I429320,I422976);
not I_25106 (I429345,I429328);
DFFARX1 I_25107 (I429345,I2507,I429195,I429371,);
not I_25108 (I429379,I429371);
nor I_25109 (I429187,I429229,I429379);
DFFARX1 I_25110 (I422985,I2507,I429195,I429419,);
nor I_25111 (I429178,I429419,I429289);
nor I_25112 (I429169,I429419,I429345);
nand I_25113 (I429455,I422979,I422967);
and I_25114 (I429472,I429455,I422964);
DFFARX1 I_25115 (I429472,I2507,I429195,I429498,);
not I_25116 (I429506,I429498);
nand I_25117 (I429523,I429506,I429419);
nand I_25118 (I429172,I429506,I429328);
nor I_25119 (I429554,I422982,I422967);
and I_25120 (I429571,I429419,I429554);
nor I_25121 (I429588,I429506,I429571);
DFFARX1 I_25122 (I429588,I2507,I429195,I429181,);
nor I_25123 (I429619,I429221,I429554);
DFFARX1 I_25124 (I429619,I2507,I429195,I429166,);
nor I_25125 (I429650,I429498,I429554);
not I_25126 (I429667,I429650);
nand I_25127 (I429175,I429667,I429523);
not I_25128 (I429722,I2514);
DFFARX1 I_25129 (I359381,I2507,I429722,I429748,);
not I_25130 (I429756,I429748);
nand I_25131 (I429773,I359384,I359381);
and I_25132 (I429790,I429773,I359393);
DFFARX1 I_25133 (I429790,I2507,I429722,I429816,);
DFFARX1 I_25134 (I429816,I2507,I429722,I429711,);
DFFARX1 I_25135 (I359390,I2507,I429722,I429847,);
nand I_25136 (I429855,I429847,I359396);
not I_25137 (I429872,I429855);
DFFARX1 I_25138 (I429872,I2507,I429722,I429898,);
not I_25139 (I429906,I429898);
nor I_25140 (I429714,I429756,I429906);
DFFARX1 I_25141 (I359405,I2507,I429722,I429946,);
nor I_25142 (I429705,I429946,I429816);
nor I_25143 (I429696,I429946,I429872);
nand I_25144 (I429982,I359399,I359387);
and I_25145 (I429999,I429982,I359384);
DFFARX1 I_25146 (I429999,I2507,I429722,I430025,);
not I_25147 (I430033,I430025);
nand I_25148 (I430050,I430033,I429946);
nand I_25149 (I429699,I430033,I429855);
nor I_25150 (I430081,I359402,I359387);
and I_25151 (I430098,I429946,I430081);
nor I_25152 (I430115,I430033,I430098);
DFFARX1 I_25153 (I430115,I2507,I429722,I429708,);
nor I_25154 (I430146,I429748,I430081);
DFFARX1 I_25155 (I430146,I2507,I429722,I429693,);
nor I_25156 (I430177,I430025,I430081);
not I_25157 (I430194,I430177);
nand I_25158 (I429702,I430194,I430050);
not I_25159 (I430249,I2514);
DFFARX1 I_25160 (I568286,I2507,I430249,I430275,);
not I_25161 (I430283,I430275);
nand I_25162 (I430300,I568295,I568283);
and I_25163 (I430317,I430300,I568280);
DFFARX1 I_25164 (I430317,I2507,I430249,I430343,);
DFFARX1 I_25165 (I430343,I2507,I430249,I430238,);
DFFARX1 I_25166 (I568280,I2507,I430249,I430374,);
nand I_25167 (I430382,I430374,I568277);
not I_25168 (I430399,I430382);
DFFARX1 I_25169 (I430399,I2507,I430249,I430425,);
not I_25170 (I430433,I430425);
nor I_25171 (I430241,I430283,I430433);
DFFARX1 I_25172 (I568283,I2507,I430249,I430473,);
nor I_25173 (I430232,I430473,I430343);
nor I_25174 (I430223,I430473,I430399);
nand I_25175 (I430509,I568298,I568289);
and I_25176 (I430526,I430509,I568292);
DFFARX1 I_25177 (I430526,I2507,I430249,I430552,);
not I_25178 (I430560,I430552);
nand I_25179 (I430577,I430560,I430473);
nand I_25180 (I430226,I430560,I430382);
nor I_25181 (I430608,I568277,I568289);
and I_25182 (I430625,I430473,I430608);
nor I_25183 (I430642,I430560,I430625);
DFFARX1 I_25184 (I430642,I2507,I430249,I430235,);
nor I_25185 (I430673,I430275,I430608);
DFFARX1 I_25186 (I430673,I2507,I430249,I430220,);
nor I_25187 (I430704,I430552,I430608);
not I_25188 (I430721,I430704);
nand I_25189 (I430229,I430721,I430577);
not I_25190 (I430776,I2514);
DFFARX1 I_25191 (I392905,I2507,I430776,I430802,);
not I_25192 (I430810,I430802);
nand I_25193 (I430827,I392908,I392905);
and I_25194 (I430844,I430827,I392917);
DFFARX1 I_25195 (I430844,I2507,I430776,I430870,);
DFFARX1 I_25196 (I430870,I2507,I430776,I430765,);
DFFARX1 I_25197 (I392914,I2507,I430776,I430901,);
nand I_25198 (I430909,I430901,I392920);
not I_25199 (I430926,I430909);
DFFARX1 I_25200 (I430926,I2507,I430776,I430952,);
not I_25201 (I430960,I430952);
nor I_25202 (I430768,I430810,I430960);
DFFARX1 I_25203 (I392929,I2507,I430776,I431000,);
nor I_25204 (I430759,I431000,I430870);
nor I_25205 (I430750,I431000,I430926);
nand I_25206 (I431036,I392923,I392911);
and I_25207 (I431053,I431036,I392908);
DFFARX1 I_25208 (I431053,I2507,I430776,I431079,);
not I_25209 (I431087,I431079);
nand I_25210 (I431104,I431087,I431000);
nand I_25211 (I430753,I431087,I430909);
nor I_25212 (I431135,I392926,I392911);
and I_25213 (I431152,I431000,I431135);
nor I_25214 (I431169,I431087,I431152);
DFFARX1 I_25215 (I431169,I2507,I430776,I430762,);
nor I_25216 (I431200,I430802,I431135);
DFFARX1 I_25217 (I431200,I2507,I430776,I430747,);
nor I_25218 (I431231,I431079,I431135);
not I_25219 (I431248,I431231);
nand I_25220 (I430756,I431248,I431104);
not I_25221 (I431303,I2514);
DFFARX1 I_25222 (I620247,I2507,I431303,I431329,);
not I_25223 (I431337,I431329);
nand I_25224 (I431354,I620229,I620229);
and I_25225 (I431371,I431354,I620235);
DFFARX1 I_25226 (I431371,I2507,I431303,I431397,);
DFFARX1 I_25227 (I431397,I2507,I431303,I431292,);
DFFARX1 I_25228 (I620232,I2507,I431303,I431428,);
nand I_25229 (I431436,I431428,I620241);
not I_25230 (I431453,I431436);
DFFARX1 I_25231 (I431453,I2507,I431303,I431479,);
not I_25232 (I431487,I431479);
nor I_25233 (I431295,I431337,I431487);
DFFARX1 I_25234 (I620253,I2507,I431303,I431527,);
nor I_25235 (I431286,I431527,I431397);
nor I_25236 (I431277,I431527,I431453);
nand I_25237 (I431563,I620244,I620238);
and I_25238 (I431580,I431563,I620232);
DFFARX1 I_25239 (I431580,I2507,I431303,I431606,);
not I_25240 (I431614,I431606);
nand I_25241 (I431631,I431614,I431527);
nand I_25242 (I431280,I431614,I431436);
nor I_25243 (I431662,I620250,I620238);
and I_25244 (I431679,I431527,I431662);
nor I_25245 (I431696,I431614,I431679);
DFFARX1 I_25246 (I431696,I2507,I431303,I431289,);
nor I_25247 (I431727,I431329,I431662);
DFFARX1 I_25248 (I431727,I2507,I431303,I431274,);
nor I_25249 (I431758,I431606,I431662);
not I_25250 (I431775,I431758);
nand I_25251 (I431283,I431775,I431631);
not I_25252 (I431830,I2514);
DFFARX1 I_25253 (I332808,I2507,I431830,I431856,);
not I_25254 (I431864,I431856);
nand I_25255 (I431881,I332793,I332814);
and I_25256 (I431898,I431881,I332802);
DFFARX1 I_25257 (I431898,I2507,I431830,I431924,);
DFFARX1 I_25258 (I431924,I2507,I431830,I431819,);
DFFARX1 I_25259 (I332796,I2507,I431830,I431955,);
nand I_25260 (I431963,I431955,I332805);
not I_25261 (I431980,I431963);
DFFARX1 I_25262 (I431980,I2507,I431830,I432006,);
not I_25263 (I432014,I432006);
nor I_25264 (I431822,I431864,I432014);
DFFARX1 I_25265 (I332811,I2507,I431830,I432054,);
nor I_25266 (I431813,I432054,I431924);
nor I_25267 (I431804,I432054,I431980);
nand I_25268 (I432090,I332793,I332796);
and I_25269 (I432107,I432090,I332817);
DFFARX1 I_25270 (I432107,I2507,I431830,I432133,);
not I_25271 (I432141,I432133);
nand I_25272 (I432158,I432141,I432054);
nand I_25273 (I431807,I432141,I431963);
nor I_25274 (I432189,I332799,I332796);
and I_25275 (I432206,I432054,I432189);
nor I_25276 (I432223,I432141,I432206);
DFFARX1 I_25277 (I432223,I2507,I431830,I431816,);
nor I_25278 (I432254,I431856,I432189);
DFFARX1 I_25279 (I432254,I2507,I431830,I431801,);
nor I_25280 (I432285,I432133,I432189);
not I_25281 (I432302,I432285);
nand I_25282 (I431810,I432302,I432158);
not I_25283 (I432357,I2514);
DFFARX1 I_25284 (I231870,I2507,I432357,I432383,);
not I_25285 (I432391,I432383);
nand I_25286 (I432408,I231867,I231876);
and I_25287 (I432425,I432408,I231885);
DFFARX1 I_25288 (I432425,I2507,I432357,I432451,);
DFFARX1 I_25289 (I432451,I2507,I432357,I432346,);
DFFARX1 I_25290 (I231888,I2507,I432357,I432482,);
nand I_25291 (I432490,I432482,I231891);
not I_25292 (I432507,I432490);
DFFARX1 I_25293 (I432507,I2507,I432357,I432533,);
not I_25294 (I432541,I432533);
nor I_25295 (I432349,I432391,I432541);
DFFARX1 I_25296 (I231864,I2507,I432357,I432581,);
nor I_25297 (I432340,I432581,I432451);
nor I_25298 (I432331,I432581,I432507);
nand I_25299 (I432617,I231879,I231882);
and I_25300 (I432634,I432617,I231873);
DFFARX1 I_25301 (I432634,I2507,I432357,I432660,);
not I_25302 (I432668,I432660);
nand I_25303 (I432685,I432668,I432581);
nand I_25304 (I432334,I432668,I432490);
nor I_25305 (I432716,I231864,I231882);
and I_25306 (I432733,I432581,I432716);
nor I_25307 (I432750,I432668,I432733);
DFFARX1 I_25308 (I432750,I2507,I432357,I432343,);
nor I_25309 (I432781,I432383,I432716);
DFFARX1 I_25310 (I432781,I2507,I432357,I432328,);
nor I_25311 (I432812,I432660,I432716);
not I_25312 (I432829,I432812);
nand I_25313 (I432337,I432829,I432685);
not I_25314 (I432884,I2514);
DFFARX1 I_25315 (I267774,I2507,I432884,I432910,);
not I_25316 (I432918,I432910);
nand I_25317 (I432935,I267771,I267780);
and I_25318 (I432952,I432935,I267789);
DFFARX1 I_25319 (I432952,I2507,I432884,I432978,);
DFFARX1 I_25320 (I432978,I2507,I432884,I432873,);
DFFARX1 I_25321 (I267792,I2507,I432884,I433009,);
nand I_25322 (I433017,I433009,I267795);
not I_25323 (I433034,I433017);
DFFARX1 I_25324 (I433034,I2507,I432884,I433060,);
not I_25325 (I433068,I433060);
nor I_25326 (I432876,I432918,I433068);
DFFARX1 I_25327 (I267768,I2507,I432884,I433108,);
nor I_25328 (I432867,I433108,I432978);
nor I_25329 (I432858,I433108,I433034);
nand I_25330 (I433144,I267783,I267786);
and I_25331 (I433161,I433144,I267777);
DFFARX1 I_25332 (I433161,I2507,I432884,I433187,);
not I_25333 (I433195,I433187);
nand I_25334 (I433212,I433195,I433108);
nand I_25335 (I432861,I433195,I433017);
nor I_25336 (I433243,I267768,I267786);
and I_25337 (I433260,I433108,I433243);
nor I_25338 (I433277,I433195,I433260);
DFFARX1 I_25339 (I433277,I2507,I432884,I432870,);
nor I_25340 (I433308,I432910,I433243);
DFFARX1 I_25341 (I433308,I2507,I432884,I432855,);
nor I_25342 (I433339,I433187,I433243);
not I_25343 (I433356,I433339);
nand I_25344 (I432864,I433356,I433212);
not I_25345 (I433411,I2514);
DFFARX1 I_25346 (I410245,I2507,I433411,I433437,);
not I_25347 (I433445,I433437);
nand I_25348 (I433462,I410248,I410245);
and I_25349 (I433479,I433462,I410257);
DFFARX1 I_25350 (I433479,I2507,I433411,I433505,);
DFFARX1 I_25351 (I433505,I2507,I433411,I433400,);
DFFARX1 I_25352 (I410254,I2507,I433411,I433536,);
nand I_25353 (I433544,I433536,I410260);
not I_25354 (I433561,I433544);
DFFARX1 I_25355 (I433561,I2507,I433411,I433587,);
not I_25356 (I433595,I433587);
nor I_25357 (I433403,I433445,I433595);
DFFARX1 I_25358 (I410269,I2507,I433411,I433635,);
nor I_25359 (I433394,I433635,I433505);
nor I_25360 (I433385,I433635,I433561);
nand I_25361 (I433671,I410263,I410251);
and I_25362 (I433688,I433671,I410248);
DFFARX1 I_25363 (I433688,I2507,I433411,I433714,);
not I_25364 (I433722,I433714);
nand I_25365 (I433739,I433722,I433635);
nand I_25366 (I433388,I433722,I433544);
nor I_25367 (I433770,I410266,I410251);
and I_25368 (I433787,I433635,I433770);
nor I_25369 (I433804,I433722,I433787);
DFFARX1 I_25370 (I433804,I2507,I433411,I433397,);
nor I_25371 (I433835,I433437,I433770);
DFFARX1 I_25372 (I433835,I2507,I433411,I433382,);
nor I_25373 (I433866,I433714,I433770);
not I_25374 (I433883,I433866);
nand I_25375 (I433391,I433883,I433739);
not I_25376 (I433938,I2514);
DFFARX1 I_25377 (I287324,I2507,I433938,I433964,);
not I_25378 (I433972,I433964);
nand I_25379 (I433989,I287342,I287333);
and I_25380 (I434006,I433989,I287336);
DFFARX1 I_25381 (I434006,I2507,I433938,I434032,);
DFFARX1 I_25382 (I434032,I2507,I433938,I433927,);
DFFARX1 I_25383 (I287330,I2507,I433938,I434063,);
nand I_25384 (I434071,I434063,I287321);
not I_25385 (I434088,I434071);
DFFARX1 I_25386 (I434088,I2507,I433938,I434114,);
not I_25387 (I434122,I434114);
nor I_25388 (I433930,I433972,I434122);
DFFARX1 I_25389 (I287327,I2507,I433938,I434162,);
nor I_25390 (I433921,I434162,I434032);
nor I_25391 (I433912,I434162,I434088);
nand I_25392 (I434198,I287321,I287318);
and I_25393 (I434215,I434198,I287339);
DFFARX1 I_25394 (I434215,I2507,I433938,I434241,);
not I_25395 (I434249,I434241);
nand I_25396 (I434266,I434249,I434162);
nand I_25397 (I433915,I434249,I434071);
nor I_25398 (I434297,I287318,I287318);
and I_25399 (I434314,I434162,I434297);
nor I_25400 (I434331,I434249,I434314);
DFFARX1 I_25401 (I434331,I2507,I433938,I433924,);
nor I_25402 (I434362,I433964,I434297);
DFFARX1 I_25403 (I434362,I2507,I433938,I433909,);
nor I_25404 (I434393,I434241,I434297);
not I_25405 (I434410,I434393);
nand I_25406 (I433918,I434410,I434266);
not I_25407 (I434465,I2514);
DFFARX1 I_25408 (I8272,I2507,I434465,I434491,);
not I_25409 (I434499,I434491);
nand I_25410 (I434516,I8284,I8287);
and I_25411 (I434533,I434516,I8263);
DFFARX1 I_25412 (I434533,I2507,I434465,I434559,);
DFFARX1 I_25413 (I434559,I2507,I434465,I434454,);
DFFARX1 I_25414 (I8281,I2507,I434465,I434590,);
nand I_25415 (I434598,I434590,I8269);
not I_25416 (I434615,I434598);
DFFARX1 I_25417 (I434615,I2507,I434465,I434641,);
not I_25418 (I434649,I434641);
nor I_25419 (I434457,I434499,I434649);
DFFARX1 I_25420 (I8266,I2507,I434465,I434689,);
nor I_25421 (I434448,I434689,I434559);
nor I_25422 (I434439,I434689,I434615);
nand I_25423 (I434725,I8275,I8266);
and I_25424 (I434742,I434725,I8263);
DFFARX1 I_25425 (I434742,I2507,I434465,I434768,);
not I_25426 (I434776,I434768);
nand I_25427 (I434793,I434776,I434689);
nand I_25428 (I434442,I434776,I434598);
nor I_25429 (I434824,I8278,I8266);
and I_25430 (I434841,I434689,I434824);
nor I_25431 (I434858,I434776,I434841);
DFFARX1 I_25432 (I434858,I2507,I434465,I434451,);
nor I_25433 (I434889,I434491,I434824);
DFFARX1 I_25434 (I434889,I2507,I434465,I434436,);
nor I_25435 (I434920,I434768,I434824);
not I_25436 (I434937,I434920);
nand I_25437 (I434445,I434937,I434793);
not I_25438 (I434992,I2514);
DFFARX1 I_25439 (I116355,I2507,I434992,I435018,);
not I_25440 (I435026,I435018);
nand I_25441 (I435043,I116352,I116370);
and I_25442 (I435060,I435043,I116361);
DFFARX1 I_25443 (I435060,I2507,I434992,I435086,);
DFFARX1 I_25444 (I435086,I2507,I434992,I434981,);
DFFARX1 I_25445 (I116367,I2507,I434992,I435117,);
nand I_25446 (I435125,I435117,I116364);
not I_25447 (I435142,I435125);
DFFARX1 I_25448 (I435142,I2507,I434992,I435168,);
not I_25449 (I435176,I435168);
nor I_25450 (I434984,I435026,I435176);
DFFARX1 I_25451 (I116358,I2507,I434992,I435216,);
nor I_25452 (I434975,I435216,I435086);
nor I_25453 (I434966,I435216,I435142);
nand I_25454 (I435252,I116349,I116373);
and I_25455 (I435269,I435252,I116352);
DFFARX1 I_25456 (I435269,I2507,I434992,I435295,);
not I_25457 (I435303,I435295);
nand I_25458 (I435320,I435303,I435216);
nand I_25459 (I434969,I435303,I435125);
nor I_25460 (I435351,I116349,I116373);
and I_25461 (I435368,I435216,I435351);
nor I_25462 (I435385,I435303,I435368);
DFFARX1 I_25463 (I435385,I2507,I434992,I434978,);
nor I_25464 (I435416,I435018,I435351);
DFFARX1 I_25465 (I435416,I2507,I434992,I434963,);
nor I_25466 (I435447,I435295,I435351);
not I_25467 (I435464,I435447);
nand I_25468 (I434972,I435464,I435320);
not I_25469 (I435519,I2514);
DFFARX1 I_25470 (I691848,I2507,I435519,I435545,);
not I_25471 (I435553,I435545);
nand I_25472 (I435570,I691845,I691854);
and I_25473 (I435587,I435570,I691833);
DFFARX1 I_25474 (I435587,I2507,I435519,I435613,);
DFFARX1 I_25475 (I435613,I2507,I435519,I435508,);
DFFARX1 I_25476 (I691836,I2507,I435519,I435644,);
nand I_25477 (I435652,I435644,I691851);
not I_25478 (I435669,I435652);
DFFARX1 I_25479 (I435669,I2507,I435519,I435695,);
not I_25480 (I435703,I435695);
nor I_25481 (I435511,I435553,I435703);
DFFARX1 I_25482 (I691857,I2507,I435519,I435743,);
nor I_25483 (I435502,I435743,I435613);
nor I_25484 (I435493,I435743,I435669);
nand I_25485 (I435779,I691839,I691860);
and I_25486 (I435796,I435779,I691842);
DFFARX1 I_25487 (I435796,I2507,I435519,I435822,);
not I_25488 (I435830,I435822);
nand I_25489 (I435847,I435830,I435743);
nand I_25490 (I435496,I435830,I435652);
nor I_25491 (I435878,I691833,I691860);
and I_25492 (I435895,I435743,I435878);
nor I_25493 (I435912,I435830,I435895);
DFFARX1 I_25494 (I435912,I2507,I435519,I435505,);
nor I_25495 (I435943,I435545,I435878);
DFFARX1 I_25496 (I435943,I2507,I435519,I435490,);
nor I_25497 (I435974,I435822,I435878);
not I_25498 (I435991,I435974);
nand I_25499 (I435499,I435991,I435847);
not I_25500 (I436046,I2514);
DFFARX1 I_25501 (I82594,I2507,I436046,I436072,);
not I_25502 (I436080,I436072);
nand I_25503 (I436097,I82570,I82579);
and I_25504 (I436114,I436097,I82573);
DFFARX1 I_25505 (I436114,I2507,I436046,I436140,);
DFFARX1 I_25506 (I436140,I2507,I436046,I436035,);
DFFARX1 I_25507 (I82591,I2507,I436046,I436171,);
nand I_25508 (I436179,I436171,I82582);
not I_25509 (I436196,I436179);
DFFARX1 I_25510 (I436196,I2507,I436046,I436222,);
not I_25511 (I436230,I436222);
nor I_25512 (I436038,I436080,I436230);
DFFARX1 I_25513 (I82576,I2507,I436046,I436270,);
nor I_25514 (I436029,I436270,I436140);
nor I_25515 (I436020,I436270,I436196);
nand I_25516 (I436306,I82588,I82585);
and I_25517 (I436323,I436306,I82573);
DFFARX1 I_25518 (I436323,I2507,I436046,I436349,);
not I_25519 (I436357,I436349);
nand I_25520 (I436374,I436357,I436270);
nand I_25521 (I436023,I436357,I436179);
nor I_25522 (I436405,I82570,I82585);
and I_25523 (I436422,I436270,I436405);
nor I_25524 (I436439,I436357,I436422);
DFFARX1 I_25525 (I436439,I2507,I436046,I436032,);
nor I_25526 (I436470,I436072,I436405);
DFFARX1 I_25527 (I436470,I2507,I436046,I436017,);
nor I_25528 (I436501,I436349,I436405);
not I_25529 (I436518,I436501);
nand I_25530 (I436026,I436518,I436374);
not I_25531 (I436573,I2514);
DFFARX1 I_25532 (I267230,I2507,I436573,I436599,);
not I_25533 (I436607,I436599);
nand I_25534 (I436624,I267227,I267236);
and I_25535 (I436641,I436624,I267245);
DFFARX1 I_25536 (I436641,I2507,I436573,I436667,);
DFFARX1 I_25537 (I436667,I2507,I436573,I436562,);
DFFARX1 I_25538 (I267248,I2507,I436573,I436698,);
nand I_25539 (I436706,I436698,I267251);
not I_25540 (I436723,I436706);
DFFARX1 I_25541 (I436723,I2507,I436573,I436749,);
not I_25542 (I436757,I436749);
nor I_25543 (I436565,I436607,I436757);
DFFARX1 I_25544 (I267224,I2507,I436573,I436797,);
nor I_25545 (I436556,I436797,I436667);
nor I_25546 (I436547,I436797,I436723);
nand I_25547 (I436833,I267239,I267242);
and I_25548 (I436850,I436833,I267233);
DFFARX1 I_25549 (I436850,I2507,I436573,I436876,);
not I_25550 (I436884,I436876);
nand I_25551 (I436901,I436884,I436797);
nand I_25552 (I436550,I436884,I436706);
nor I_25553 (I436932,I267224,I267242);
and I_25554 (I436949,I436797,I436932);
nor I_25555 (I436966,I436884,I436949);
DFFARX1 I_25556 (I436966,I2507,I436573,I436559,);
nor I_25557 (I436997,I436599,I436932);
DFFARX1 I_25558 (I436997,I2507,I436573,I436544,);
nor I_25559 (I437028,I436876,I436932);
not I_25560 (I437045,I437028);
nand I_25561 (I436553,I437045,I436901);
not I_25562 (I437100,I2514);
DFFARX1 I_25563 (I727548,I2507,I437100,I437126,);
not I_25564 (I437134,I437126);
nand I_25565 (I437151,I727545,I727554);
and I_25566 (I437168,I437151,I727533);
DFFARX1 I_25567 (I437168,I2507,I437100,I437194,);
DFFARX1 I_25568 (I437194,I2507,I437100,I437089,);
DFFARX1 I_25569 (I727536,I2507,I437100,I437225,);
nand I_25570 (I437233,I437225,I727551);
not I_25571 (I437250,I437233);
DFFARX1 I_25572 (I437250,I2507,I437100,I437276,);
not I_25573 (I437284,I437276);
nor I_25574 (I437092,I437134,I437284);
DFFARX1 I_25575 (I727557,I2507,I437100,I437324,);
nor I_25576 (I437083,I437324,I437194);
nor I_25577 (I437074,I437324,I437250);
nand I_25578 (I437360,I727539,I727560);
and I_25579 (I437377,I437360,I727542);
DFFARX1 I_25580 (I437377,I2507,I437100,I437403,);
not I_25581 (I437411,I437403);
nand I_25582 (I437428,I437411,I437324);
nand I_25583 (I437077,I437411,I437233);
nor I_25584 (I437459,I727533,I727560);
and I_25585 (I437476,I437324,I437459);
nor I_25586 (I437493,I437411,I437476);
DFFARX1 I_25587 (I437493,I2507,I437100,I437086,);
nor I_25588 (I437524,I437126,I437459);
DFFARX1 I_25589 (I437524,I2507,I437100,I437071,);
nor I_25590 (I437555,I437403,I437459);
not I_25591 (I437572,I437555);
nand I_25592 (I437080,I437572,I437428);
not I_25593 (I437627,I2514);
DFFARX1 I_25594 (I520289,I2507,I437627,I437653,);
not I_25595 (I437661,I437653);
nand I_25596 (I437678,I520304,I520286);
and I_25597 (I437695,I437678,I520286);
DFFARX1 I_25598 (I437695,I2507,I437627,I437721,);
DFFARX1 I_25599 (I437721,I2507,I437627,I437616,);
DFFARX1 I_25600 (I520295,I2507,I437627,I437752,);
nand I_25601 (I437760,I437752,I520313);
not I_25602 (I437777,I437760);
DFFARX1 I_25603 (I437777,I2507,I437627,I437803,);
not I_25604 (I437811,I437803);
nor I_25605 (I437619,I437661,I437811);
DFFARX1 I_25606 (I520310,I2507,I437627,I437851,);
nor I_25607 (I437610,I437851,I437721);
nor I_25608 (I437601,I437851,I437777);
nand I_25609 (I437887,I520307,I520298);
and I_25610 (I437904,I437887,I520292);
DFFARX1 I_25611 (I437904,I2507,I437627,I437930,);
not I_25612 (I437938,I437930);
nand I_25613 (I437955,I437938,I437851);
nand I_25614 (I437604,I437938,I437760);
nor I_25615 (I437986,I520301,I520298);
and I_25616 (I438003,I437851,I437986);
nor I_25617 (I438020,I437938,I438003);
DFFARX1 I_25618 (I438020,I2507,I437627,I437613,);
nor I_25619 (I438051,I437653,I437986);
DFFARX1 I_25620 (I438051,I2507,I437627,I437598,);
nor I_25621 (I438082,I437930,I437986);
not I_25622 (I438099,I438082);
nand I_25623 (I437607,I438099,I437955);
not I_25624 (I438154,I2514);
DFFARX1 I_25625 (I519643,I2507,I438154,I438180,);
not I_25626 (I438188,I438180);
nand I_25627 (I438205,I519658,I519640);
and I_25628 (I438222,I438205,I519640);
DFFARX1 I_25629 (I438222,I2507,I438154,I438248,);
DFFARX1 I_25630 (I438248,I2507,I438154,I438143,);
DFFARX1 I_25631 (I519649,I2507,I438154,I438279,);
nand I_25632 (I438287,I438279,I519667);
not I_25633 (I438304,I438287);
DFFARX1 I_25634 (I438304,I2507,I438154,I438330,);
not I_25635 (I438338,I438330);
nor I_25636 (I438146,I438188,I438338);
DFFARX1 I_25637 (I519664,I2507,I438154,I438378,);
nor I_25638 (I438137,I438378,I438248);
nor I_25639 (I438128,I438378,I438304);
nand I_25640 (I438414,I519661,I519652);
and I_25641 (I438431,I438414,I519646);
DFFARX1 I_25642 (I438431,I2507,I438154,I438457,);
not I_25643 (I438465,I438457);
nand I_25644 (I438482,I438465,I438378);
nand I_25645 (I438131,I438465,I438287);
nor I_25646 (I438513,I519655,I519652);
and I_25647 (I438530,I438378,I438513);
nor I_25648 (I438547,I438465,I438530);
DFFARX1 I_25649 (I438547,I2507,I438154,I438140,);
nor I_25650 (I438578,I438180,I438513);
DFFARX1 I_25651 (I438578,I2507,I438154,I438125,);
nor I_25652 (I438609,I438457,I438513);
not I_25653 (I438626,I438609);
nand I_25654 (I438134,I438626,I438482);
not I_25655 (I438681,I2514);
DFFARX1 I_25656 (I62041,I2507,I438681,I438707,);
not I_25657 (I438715,I438707);
nand I_25658 (I438732,I62017,I62026);
and I_25659 (I438749,I438732,I62020);
DFFARX1 I_25660 (I438749,I2507,I438681,I438775,);
DFFARX1 I_25661 (I438775,I2507,I438681,I438670,);
DFFARX1 I_25662 (I62038,I2507,I438681,I438806,);
nand I_25663 (I438814,I438806,I62029);
not I_25664 (I438831,I438814);
DFFARX1 I_25665 (I438831,I2507,I438681,I438857,);
not I_25666 (I438865,I438857);
nor I_25667 (I438673,I438715,I438865);
DFFARX1 I_25668 (I62023,I2507,I438681,I438905,);
nor I_25669 (I438664,I438905,I438775);
nor I_25670 (I438655,I438905,I438831);
nand I_25671 (I438941,I62035,I62032);
and I_25672 (I438958,I438941,I62020);
DFFARX1 I_25673 (I438958,I2507,I438681,I438984,);
not I_25674 (I438992,I438984);
nand I_25675 (I439009,I438992,I438905);
nand I_25676 (I438658,I438992,I438814);
nor I_25677 (I439040,I62017,I62032);
and I_25678 (I439057,I438905,I439040);
nor I_25679 (I439074,I438992,I439057);
DFFARX1 I_25680 (I439074,I2507,I438681,I438667,);
nor I_25681 (I439105,I438707,I439040);
DFFARX1 I_25682 (I439105,I2507,I438681,I438652,);
nor I_25683 (I439136,I438984,I439040);
not I_25684 (I439153,I439136);
nand I_25685 (I438661,I439153,I439009);
not I_25686 (I439208,I2514);
DFFARX1 I_25687 (I340900,I2507,I439208,I439234,);
not I_25688 (I439242,I439234);
nand I_25689 (I439259,I340885,I340906);
and I_25690 (I439276,I439259,I340894);
DFFARX1 I_25691 (I439276,I2507,I439208,I439302,);
DFFARX1 I_25692 (I439302,I2507,I439208,I439197,);
DFFARX1 I_25693 (I340888,I2507,I439208,I439333,);
nand I_25694 (I439341,I439333,I340897);
not I_25695 (I439358,I439341);
DFFARX1 I_25696 (I439358,I2507,I439208,I439384,);
not I_25697 (I439392,I439384);
nor I_25698 (I439200,I439242,I439392);
DFFARX1 I_25699 (I340903,I2507,I439208,I439432,);
nor I_25700 (I439191,I439432,I439302);
nor I_25701 (I439182,I439432,I439358);
nand I_25702 (I439468,I340885,I340888);
and I_25703 (I439485,I439468,I340909);
DFFARX1 I_25704 (I439485,I2507,I439208,I439511,);
not I_25705 (I439519,I439511);
nand I_25706 (I439536,I439519,I439432);
nand I_25707 (I439185,I439519,I439341);
nor I_25708 (I439567,I340891,I340888);
and I_25709 (I439584,I439432,I439567);
nor I_25710 (I439601,I439519,I439584);
DFFARX1 I_25711 (I439601,I2507,I439208,I439194,);
nor I_25712 (I439632,I439234,I439567);
DFFARX1 I_25713 (I439632,I2507,I439208,I439179,);
nor I_25714 (I439663,I439511,I439567);
not I_25715 (I439680,I439663);
nand I_25716 (I439188,I439680,I439536);
not I_25717 (I439735,I2514);
DFFARX1 I_25718 (I695418,I2507,I439735,I439761,);
not I_25719 (I439769,I439761);
nand I_25720 (I439786,I695415,I695424);
and I_25721 (I439803,I439786,I695403);
DFFARX1 I_25722 (I439803,I2507,I439735,I439829,);
DFFARX1 I_25723 (I439829,I2507,I439735,I439724,);
DFFARX1 I_25724 (I695406,I2507,I439735,I439860,);
nand I_25725 (I439868,I439860,I695421);
not I_25726 (I439885,I439868);
DFFARX1 I_25727 (I439885,I2507,I439735,I439911,);
not I_25728 (I439919,I439911);
nor I_25729 (I439727,I439769,I439919);
DFFARX1 I_25730 (I695427,I2507,I439735,I439959,);
nor I_25731 (I439718,I439959,I439829);
nor I_25732 (I439709,I439959,I439885);
nand I_25733 (I439995,I695409,I695430);
and I_25734 (I440012,I439995,I695412);
DFFARX1 I_25735 (I440012,I2507,I439735,I440038,);
not I_25736 (I440046,I440038);
nand I_25737 (I440063,I440046,I439959);
nand I_25738 (I439712,I440046,I439868);
nor I_25739 (I440094,I695403,I695430);
and I_25740 (I440111,I439959,I440094);
nor I_25741 (I440128,I440046,I440111);
DFFARX1 I_25742 (I440128,I2507,I439735,I439721,);
nor I_25743 (I440159,I439761,I440094);
DFFARX1 I_25744 (I440159,I2507,I439735,I439706,);
nor I_25745 (I440190,I440038,I440094);
not I_25746 (I440207,I440190);
nand I_25747 (I439715,I440207,I440063);
not I_25748 (I440262,I2514);
DFFARX1 I_25749 (I687776,I2507,I440262,I440288,);
not I_25750 (I440296,I440288);
nand I_25751 (I440313,I687770,I687788);
and I_25752 (I440330,I440313,I687773);
DFFARX1 I_25753 (I440330,I2507,I440262,I440356,);
DFFARX1 I_25754 (I440356,I2507,I440262,I440251,);
DFFARX1 I_25755 (I687794,I2507,I440262,I440387,);
nand I_25756 (I440395,I440387,I687779);
not I_25757 (I440412,I440395);
DFFARX1 I_25758 (I440412,I2507,I440262,I440438,);
not I_25759 (I440446,I440438);
nor I_25760 (I440254,I440296,I440446);
DFFARX1 I_25761 (I687791,I2507,I440262,I440486,);
nor I_25762 (I440245,I440486,I440356);
nor I_25763 (I440236,I440486,I440412);
nand I_25764 (I440522,I687782,I687797);
and I_25765 (I440539,I440522,I687785);
DFFARX1 I_25766 (I440539,I2507,I440262,I440565,);
not I_25767 (I440573,I440565);
nand I_25768 (I440590,I440573,I440486);
nand I_25769 (I440239,I440573,I440395);
nor I_25770 (I440621,I687770,I687797);
and I_25771 (I440638,I440486,I440621);
nor I_25772 (I440655,I440573,I440638);
DFFARX1 I_25773 (I440655,I2507,I440262,I440248,);
nor I_25774 (I440686,I440288,I440621);
DFFARX1 I_25775 (I440686,I2507,I440262,I440233,);
nor I_25776 (I440717,I440565,I440621);
not I_25777 (I440734,I440717);
nand I_25778 (I440242,I440734,I440590);
not I_25779 (I440789,I2514);
DFFARX1 I_25780 (I336854,I2507,I440789,I440815,);
not I_25781 (I440823,I440815);
nand I_25782 (I440840,I336839,I336860);
and I_25783 (I440857,I440840,I336848);
DFFARX1 I_25784 (I440857,I2507,I440789,I440883,);
DFFARX1 I_25785 (I440883,I2507,I440789,I440778,);
DFFARX1 I_25786 (I336842,I2507,I440789,I440914,);
nand I_25787 (I440922,I440914,I336851);
not I_25788 (I440939,I440922);
DFFARX1 I_25789 (I440939,I2507,I440789,I440965,);
not I_25790 (I440973,I440965);
nor I_25791 (I440781,I440823,I440973);
DFFARX1 I_25792 (I336857,I2507,I440789,I441013,);
nor I_25793 (I440772,I441013,I440883);
nor I_25794 (I440763,I441013,I440939);
nand I_25795 (I441049,I336839,I336842);
and I_25796 (I441066,I441049,I336863);
DFFARX1 I_25797 (I441066,I2507,I440789,I441092,);
not I_25798 (I441100,I441092);
nand I_25799 (I441117,I441100,I441013);
nand I_25800 (I440766,I441100,I440922);
nor I_25801 (I441148,I336845,I336842);
and I_25802 (I441165,I441013,I441148);
nor I_25803 (I441182,I441100,I441165);
DFFARX1 I_25804 (I441182,I2507,I440789,I440775,);
nor I_25805 (I441213,I440815,I441148);
DFFARX1 I_25806 (I441213,I2507,I440789,I440760,);
nor I_25807 (I441244,I441092,I441148);
not I_25808 (I441261,I441244);
nand I_25809 (I440769,I441261,I441117);
not I_25810 (I441316,I2514);
DFFARX1 I_25811 (I39907,I2507,I441316,I441342,);
not I_25812 (I441350,I441342);
nand I_25813 (I441367,I39883,I39892);
and I_25814 (I441384,I441367,I39886);
DFFARX1 I_25815 (I441384,I2507,I441316,I441410,);
DFFARX1 I_25816 (I441410,I2507,I441316,I441305,);
DFFARX1 I_25817 (I39904,I2507,I441316,I441441,);
nand I_25818 (I441449,I441441,I39895);
not I_25819 (I441466,I441449);
DFFARX1 I_25820 (I441466,I2507,I441316,I441492,);
not I_25821 (I441500,I441492);
nor I_25822 (I441308,I441350,I441500);
DFFARX1 I_25823 (I39889,I2507,I441316,I441540,);
nor I_25824 (I441299,I441540,I441410);
nor I_25825 (I441290,I441540,I441466);
nand I_25826 (I441576,I39901,I39898);
and I_25827 (I441593,I441576,I39886);
DFFARX1 I_25828 (I441593,I2507,I441316,I441619,);
not I_25829 (I441627,I441619);
nand I_25830 (I441644,I441627,I441540);
nand I_25831 (I441293,I441627,I441449);
nor I_25832 (I441675,I39883,I39898);
and I_25833 (I441692,I441540,I441675);
nor I_25834 (I441709,I441627,I441692);
DFFARX1 I_25835 (I441709,I2507,I441316,I441302,);
nor I_25836 (I441740,I441342,I441675);
DFFARX1 I_25837 (I441740,I2507,I441316,I441287,);
nor I_25838 (I441771,I441619,I441675);
not I_25839 (I441788,I441771);
nand I_25840 (I441296,I441788,I441644);
not I_25841 (I441843,I2514);
DFFARX1 I_25842 (I320092,I2507,I441843,I441869,);
not I_25843 (I441877,I441869);
nand I_25844 (I441894,I320077,I320098);
and I_25845 (I441911,I441894,I320086);
DFFARX1 I_25846 (I441911,I2507,I441843,I441937,);
DFFARX1 I_25847 (I441937,I2507,I441843,I441832,);
DFFARX1 I_25848 (I320080,I2507,I441843,I441968,);
nand I_25849 (I441976,I441968,I320089);
not I_25850 (I441993,I441976);
DFFARX1 I_25851 (I441993,I2507,I441843,I442019,);
not I_25852 (I442027,I442019);
nor I_25853 (I441835,I441877,I442027);
DFFARX1 I_25854 (I320095,I2507,I441843,I442067,);
nor I_25855 (I441826,I442067,I441937);
nor I_25856 (I441817,I442067,I441993);
nand I_25857 (I442103,I320077,I320080);
and I_25858 (I442120,I442103,I320101);
DFFARX1 I_25859 (I442120,I2507,I441843,I442146,);
not I_25860 (I442154,I442146);
nand I_25861 (I442171,I442154,I442067);
nand I_25862 (I441820,I442154,I441976);
nor I_25863 (I442202,I320083,I320080);
and I_25864 (I442219,I442067,I442202);
nor I_25865 (I442236,I442154,I442219);
DFFARX1 I_25866 (I442236,I2507,I441843,I441829,);
nor I_25867 (I442267,I441869,I442202);
DFFARX1 I_25868 (I442267,I2507,I441843,I441814,);
nor I_25869 (I442298,I442146,I442202);
not I_25870 (I442315,I442298);
nand I_25871 (I441823,I442315,I442171);
not I_25872 (I442370,I2514);
DFFARX1 I_25873 (I3127,I2507,I442370,I442396,);
not I_25874 (I442404,I442396);
nand I_25875 (I442421,I3133,I3115);
and I_25876 (I442438,I442421,I3124);
DFFARX1 I_25877 (I442438,I2507,I442370,I442464,);
DFFARX1 I_25878 (I442464,I2507,I442370,I442359,);
DFFARX1 I_25879 (I3115,I2507,I442370,I442495,);
nand I_25880 (I442503,I442495,I3118);
not I_25881 (I442520,I442503);
DFFARX1 I_25882 (I442520,I2507,I442370,I442546,);
not I_25883 (I442554,I442546);
nor I_25884 (I442362,I442404,I442554);
DFFARX1 I_25885 (I3118,I2507,I442370,I442594,);
nor I_25886 (I442353,I442594,I442464);
nor I_25887 (I442344,I442594,I442520);
nand I_25888 (I442630,I3121,I3130);
and I_25889 (I442647,I442630,I3112);
DFFARX1 I_25890 (I442647,I2507,I442370,I442673,);
not I_25891 (I442681,I442673);
nand I_25892 (I442698,I442681,I442594);
nand I_25893 (I442347,I442681,I442503);
nor I_25894 (I442729,I3112,I3130);
and I_25895 (I442746,I442594,I442729);
nor I_25896 (I442763,I442681,I442746);
DFFARX1 I_25897 (I442763,I2507,I442370,I442356,);
nor I_25898 (I442794,I442396,I442729);
DFFARX1 I_25899 (I442794,I2507,I442370,I442341,);
nor I_25900 (I442825,I442673,I442729);
not I_25901 (I442842,I442825);
nand I_25902 (I442350,I442842,I442698);
not I_25903 (I442897,I2514);
DFFARX1 I_25904 (I155625,I2507,I442897,I442923,);
not I_25905 (I442931,I442923);
nand I_25906 (I442948,I155622,I155640);
and I_25907 (I442965,I442948,I155631);
DFFARX1 I_25908 (I442965,I2507,I442897,I442991,);
DFFARX1 I_25909 (I442991,I2507,I442897,I442886,);
DFFARX1 I_25910 (I155637,I2507,I442897,I443022,);
nand I_25911 (I443030,I443022,I155634);
not I_25912 (I443047,I443030);
DFFARX1 I_25913 (I443047,I2507,I442897,I443073,);
not I_25914 (I443081,I443073);
nor I_25915 (I442889,I442931,I443081);
DFFARX1 I_25916 (I155628,I2507,I442897,I443121,);
nor I_25917 (I442880,I443121,I442991);
nor I_25918 (I442871,I443121,I443047);
nand I_25919 (I443157,I155619,I155643);
and I_25920 (I443174,I443157,I155622);
DFFARX1 I_25921 (I443174,I2507,I442897,I443200,);
not I_25922 (I443208,I443200);
nand I_25923 (I443225,I443208,I443121);
nand I_25924 (I442874,I443208,I443030);
nor I_25925 (I443256,I155619,I155643);
and I_25926 (I443273,I443121,I443256);
nor I_25927 (I443290,I443208,I443273);
DFFARX1 I_25928 (I443290,I2507,I442897,I442883,);
nor I_25929 (I443321,I442923,I443256);
DFFARX1 I_25930 (I443321,I2507,I442897,I442868,);
nor I_25931 (I443352,I443200,I443256);
not I_25932 (I443369,I443352);
nand I_25933 (I442877,I443369,I443225);
not I_25934 (I443424,I2514);
DFFARX1 I_25935 (I185888,I2507,I443424,I443450,);
not I_25936 (I443458,I443450);
nand I_25937 (I443475,I185879,I185879);
and I_25938 (I443492,I443475,I185897);
DFFARX1 I_25939 (I443492,I2507,I443424,I443518,);
DFFARX1 I_25940 (I443518,I2507,I443424,I443413,);
DFFARX1 I_25941 (I185900,I2507,I443424,I443549,);
nand I_25942 (I443557,I443549,I185882);
not I_25943 (I443574,I443557);
DFFARX1 I_25944 (I443574,I2507,I443424,I443600,);
not I_25945 (I443608,I443600);
nor I_25946 (I443416,I443458,I443608);
DFFARX1 I_25947 (I185894,I2507,I443424,I443648,);
nor I_25948 (I443407,I443648,I443518);
nor I_25949 (I443398,I443648,I443574);
nand I_25950 (I443684,I185906,I185885);
and I_25951 (I443701,I443684,I185891);
DFFARX1 I_25952 (I443701,I2507,I443424,I443727,);
not I_25953 (I443735,I443727);
nand I_25954 (I443752,I443735,I443648);
nand I_25955 (I443401,I443735,I443557);
nor I_25956 (I443783,I185903,I185885);
and I_25957 (I443800,I443648,I443783);
nor I_25958 (I443817,I443735,I443800);
DFFARX1 I_25959 (I443817,I2507,I443424,I443410,);
nor I_25960 (I443848,I443450,I443783);
DFFARX1 I_25961 (I443848,I2507,I443424,I443395,);
nor I_25962 (I443879,I443727,I443783);
not I_25963 (I443896,I443879);
nand I_25964 (I443404,I443896,I443752);
not I_25965 (I443951,I2514);
DFFARX1 I_25966 (I705533,I2507,I443951,I443977,);
not I_25967 (I443985,I443977);
nand I_25968 (I444002,I705530,I705539);
and I_25969 (I444019,I444002,I705518);
DFFARX1 I_25970 (I444019,I2507,I443951,I444045,);
DFFARX1 I_25971 (I444045,I2507,I443951,I443940,);
DFFARX1 I_25972 (I705521,I2507,I443951,I444076,);
nand I_25973 (I444084,I444076,I705536);
not I_25974 (I444101,I444084);
DFFARX1 I_25975 (I444101,I2507,I443951,I444127,);
not I_25976 (I444135,I444127);
nor I_25977 (I443943,I443985,I444135);
DFFARX1 I_25978 (I705542,I2507,I443951,I444175,);
nor I_25979 (I443934,I444175,I444045);
nor I_25980 (I443925,I444175,I444101);
nand I_25981 (I444211,I705524,I705545);
and I_25982 (I444228,I444211,I705527);
DFFARX1 I_25983 (I444228,I2507,I443951,I444254,);
not I_25984 (I444262,I444254);
nand I_25985 (I444279,I444262,I444175);
nand I_25986 (I443928,I444262,I444084);
nor I_25987 (I444310,I705518,I705545);
and I_25988 (I444327,I444175,I444310);
nor I_25989 (I444344,I444262,I444327);
DFFARX1 I_25990 (I444344,I2507,I443951,I443937,);
nor I_25991 (I444375,I443977,I444310);
DFFARX1 I_25992 (I444375,I2507,I443951,I443922,);
nor I_25993 (I444406,I444254,I444310);
not I_25994 (I444423,I444406);
nand I_25995 (I443931,I444423,I444279);
not I_25996 (I444478,I2514);
DFFARX1 I_25997 (I385969,I2507,I444478,I444504,);
not I_25998 (I444512,I444504);
nand I_25999 (I444529,I385972,I385969);
and I_26000 (I444546,I444529,I385981);
DFFARX1 I_26001 (I444546,I2507,I444478,I444572,);
DFFARX1 I_26002 (I444572,I2507,I444478,I444467,);
DFFARX1 I_26003 (I385978,I2507,I444478,I444603,);
nand I_26004 (I444611,I444603,I385984);
not I_26005 (I444628,I444611);
DFFARX1 I_26006 (I444628,I2507,I444478,I444654,);
not I_26007 (I444662,I444654);
nor I_26008 (I444470,I444512,I444662);
DFFARX1 I_26009 (I385993,I2507,I444478,I444702,);
nor I_26010 (I444461,I444702,I444572);
nor I_26011 (I444452,I444702,I444628);
nand I_26012 (I444738,I385987,I385975);
and I_26013 (I444755,I444738,I385972);
DFFARX1 I_26014 (I444755,I2507,I444478,I444781,);
not I_26015 (I444789,I444781);
nand I_26016 (I444806,I444789,I444702);
nand I_26017 (I444455,I444789,I444611);
nor I_26018 (I444837,I385990,I385975);
and I_26019 (I444854,I444702,I444837);
nor I_26020 (I444871,I444789,I444854);
DFFARX1 I_26021 (I444871,I2507,I444478,I444464,);
nor I_26022 (I444902,I444504,I444837);
DFFARX1 I_26023 (I444902,I2507,I444478,I444449,);
nor I_26024 (I444933,I444781,I444837);
not I_26025 (I444950,I444933);
nand I_26026 (I444458,I444950,I444806);
not I_26027 (I445005,I2514);
DFFARX1 I_26028 (I422383,I2507,I445005,I445031,);
not I_26029 (I445039,I445031);
nand I_26030 (I445056,I422386,I422383);
and I_26031 (I445073,I445056,I422395);
DFFARX1 I_26032 (I445073,I2507,I445005,I445099,);
DFFARX1 I_26033 (I445099,I2507,I445005,I444994,);
DFFARX1 I_26034 (I422392,I2507,I445005,I445130,);
nand I_26035 (I445138,I445130,I422398);
not I_26036 (I445155,I445138);
DFFARX1 I_26037 (I445155,I2507,I445005,I445181,);
not I_26038 (I445189,I445181);
nor I_26039 (I444997,I445039,I445189);
DFFARX1 I_26040 (I422407,I2507,I445005,I445229,);
nor I_26041 (I444988,I445229,I445099);
nor I_26042 (I444979,I445229,I445155);
nand I_26043 (I445265,I422401,I422389);
and I_26044 (I445282,I445265,I422386);
DFFARX1 I_26045 (I445282,I2507,I445005,I445308,);
not I_26046 (I445316,I445308);
nand I_26047 (I445333,I445316,I445229);
nand I_26048 (I444982,I445316,I445138);
nor I_26049 (I445364,I422404,I422389);
and I_26050 (I445381,I445229,I445364);
nor I_26051 (I445398,I445316,I445381);
DFFARX1 I_26052 (I445398,I2507,I445005,I444991,);
nor I_26053 (I445429,I445031,I445364);
DFFARX1 I_26054 (I445429,I2507,I445005,I444976,);
nor I_26055 (I445460,I445308,I445364);
not I_26056 (I445477,I445460);
nand I_26057 (I444985,I445477,I445333);
not I_26058 (I445532,I2514);
DFFARX1 I_26059 (I692443,I2507,I445532,I445558,);
not I_26060 (I445566,I445558);
nand I_26061 (I445583,I692440,I692449);
and I_26062 (I445600,I445583,I692428);
DFFARX1 I_26063 (I445600,I2507,I445532,I445626,);
DFFARX1 I_26064 (I445626,I2507,I445532,I445521,);
DFFARX1 I_26065 (I692431,I2507,I445532,I445657,);
nand I_26066 (I445665,I445657,I692446);
not I_26067 (I445682,I445665);
DFFARX1 I_26068 (I445682,I2507,I445532,I445708,);
not I_26069 (I445716,I445708);
nor I_26070 (I445524,I445566,I445716);
DFFARX1 I_26071 (I692452,I2507,I445532,I445756,);
nor I_26072 (I445515,I445756,I445626);
nor I_26073 (I445506,I445756,I445682);
nand I_26074 (I445792,I692434,I692455);
and I_26075 (I445809,I445792,I692437);
DFFARX1 I_26076 (I445809,I2507,I445532,I445835,);
not I_26077 (I445843,I445835);
nand I_26078 (I445860,I445843,I445756);
nand I_26079 (I445509,I445843,I445665);
nor I_26080 (I445891,I692428,I692455);
and I_26081 (I445908,I445756,I445891);
nor I_26082 (I445925,I445843,I445908);
DFFARX1 I_26083 (I445925,I2507,I445532,I445518,);
nor I_26084 (I445956,I445558,I445891);
DFFARX1 I_26085 (I445956,I2507,I445532,I445503,);
nor I_26086 (I445987,I445835,I445891);
not I_26087 (I446004,I445987);
nand I_26088 (I445512,I446004,I445860);
not I_26089 (I446059,I2514);
DFFARX1 I_26090 (I403309,I2507,I446059,I446085,);
not I_26091 (I446093,I446085);
nand I_26092 (I446110,I403312,I403309);
and I_26093 (I446127,I446110,I403321);
DFFARX1 I_26094 (I446127,I2507,I446059,I446153,);
DFFARX1 I_26095 (I446153,I2507,I446059,I446048,);
DFFARX1 I_26096 (I403318,I2507,I446059,I446184,);
nand I_26097 (I446192,I446184,I403324);
not I_26098 (I446209,I446192);
DFFARX1 I_26099 (I446209,I2507,I446059,I446235,);
not I_26100 (I446243,I446235);
nor I_26101 (I446051,I446093,I446243);
DFFARX1 I_26102 (I403333,I2507,I446059,I446283,);
nor I_26103 (I446042,I446283,I446153);
nor I_26104 (I446033,I446283,I446209);
nand I_26105 (I446319,I403327,I403315);
and I_26106 (I446336,I446319,I403312);
DFFARX1 I_26107 (I446336,I2507,I446059,I446362,);
not I_26108 (I446370,I446362);
nand I_26109 (I446387,I446370,I446283);
nand I_26110 (I446036,I446370,I446192);
nor I_26111 (I446418,I403330,I403315);
and I_26112 (I446435,I446283,I446418);
nor I_26113 (I446452,I446370,I446435);
DFFARX1 I_26114 (I446452,I2507,I446059,I446045,);
nor I_26115 (I446483,I446085,I446418);
DFFARX1 I_26116 (I446483,I2507,I446059,I446030,);
nor I_26117 (I446514,I446362,I446418);
not I_26118 (I446531,I446514);
nand I_26119 (I446039,I446531,I446387);
not I_26120 (I446586,I2514);
DFFARX1 I_26121 (I390015,I2507,I446586,I446612,);
not I_26122 (I446620,I446612);
nand I_26123 (I446637,I390018,I390015);
and I_26124 (I446654,I446637,I390027);
DFFARX1 I_26125 (I446654,I2507,I446586,I446680,);
DFFARX1 I_26126 (I446680,I2507,I446586,I446575,);
DFFARX1 I_26127 (I390024,I2507,I446586,I446711,);
nand I_26128 (I446719,I446711,I390030);
not I_26129 (I446736,I446719);
DFFARX1 I_26130 (I446736,I2507,I446586,I446762,);
not I_26131 (I446770,I446762);
nor I_26132 (I446578,I446620,I446770);
DFFARX1 I_26133 (I390039,I2507,I446586,I446810,);
nor I_26134 (I446569,I446810,I446680);
nor I_26135 (I446560,I446810,I446736);
nand I_26136 (I446846,I390033,I390021);
and I_26137 (I446863,I446846,I390018);
DFFARX1 I_26138 (I446863,I2507,I446586,I446889,);
not I_26139 (I446897,I446889);
nand I_26140 (I446914,I446897,I446810);
nand I_26141 (I446563,I446897,I446719);
nor I_26142 (I446945,I390036,I390021);
and I_26143 (I446962,I446810,I446945);
nor I_26144 (I446979,I446897,I446962);
DFFARX1 I_26145 (I446979,I2507,I446586,I446572,);
nor I_26146 (I447010,I446612,I446945);
DFFARX1 I_26147 (I447010,I2507,I446586,I446557,);
nor I_26148 (I447041,I446889,I446945);
not I_26149 (I447058,I447041);
nand I_26150 (I446566,I447058,I446914);
not I_26151 (I447113,I2514);
DFFARX1 I_26152 (I387125,I2507,I447113,I447139,);
not I_26153 (I447147,I447139);
nand I_26154 (I447164,I387128,I387125);
and I_26155 (I447181,I447164,I387137);
DFFARX1 I_26156 (I447181,I2507,I447113,I447207,);
DFFARX1 I_26157 (I447207,I2507,I447113,I447102,);
DFFARX1 I_26158 (I387134,I2507,I447113,I447238,);
nand I_26159 (I447246,I447238,I387140);
not I_26160 (I447263,I447246);
DFFARX1 I_26161 (I447263,I2507,I447113,I447289,);
not I_26162 (I447297,I447289);
nor I_26163 (I447105,I447147,I447297);
DFFARX1 I_26164 (I387149,I2507,I447113,I447337,);
nor I_26165 (I447096,I447337,I447207);
nor I_26166 (I447087,I447337,I447263);
nand I_26167 (I447373,I387143,I387131);
and I_26168 (I447390,I447373,I387128);
DFFARX1 I_26169 (I447390,I2507,I447113,I447416,);
not I_26170 (I447424,I447416);
nand I_26171 (I447441,I447424,I447337);
nand I_26172 (I447090,I447424,I447246);
nor I_26173 (I447472,I387146,I387131);
and I_26174 (I447489,I447337,I447472);
nor I_26175 (I447506,I447424,I447489);
DFFARX1 I_26176 (I447506,I2507,I447113,I447099,);
nor I_26177 (I447537,I447139,I447472);
DFFARX1 I_26178 (I447537,I2507,I447113,I447084,);
nor I_26179 (I447568,I447416,I447472);
not I_26180 (I447585,I447568);
nand I_26181 (I447093,I447585,I447441);
not I_26182 (I447640,I2514);
DFFARX1 I_26183 (I36218,I2507,I447640,I447666,);
not I_26184 (I447674,I447666);
nand I_26185 (I447691,I36194,I36203);
and I_26186 (I447708,I447691,I36197);
DFFARX1 I_26187 (I447708,I2507,I447640,I447734,);
DFFARX1 I_26188 (I447734,I2507,I447640,I447629,);
DFFARX1 I_26189 (I36215,I2507,I447640,I447765,);
nand I_26190 (I447773,I447765,I36206);
not I_26191 (I447790,I447773);
DFFARX1 I_26192 (I447790,I2507,I447640,I447816,);
not I_26193 (I447824,I447816);
nor I_26194 (I447632,I447674,I447824);
DFFARX1 I_26195 (I36200,I2507,I447640,I447864,);
nor I_26196 (I447623,I447864,I447734);
nor I_26197 (I447614,I447864,I447790);
nand I_26198 (I447900,I36212,I36209);
and I_26199 (I447917,I447900,I36197);
DFFARX1 I_26200 (I447917,I2507,I447640,I447943,);
not I_26201 (I447951,I447943);
nand I_26202 (I447968,I447951,I447864);
nand I_26203 (I447617,I447951,I447773);
nor I_26204 (I447999,I36194,I36209);
and I_26205 (I448016,I447864,I447999);
nor I_26206 (I448033,I447951,I448016);
DFFARX1 I_26207 (I448033,I2507,I447640,I447626,);
nor I_26208 (I448064,I447666,I447999);
DFFARX1 I_26209 (I448064,I2507,I447640,I447611,);
nor I_26210 (I448095,I447943,I447999);
not I_26211 (I448112,I448095);
nand I_26212 (I447620,I448112,I447968);
not I_26213 (I448167,I2514);
DFFARX1 I_26214 (I178510,I2507,I448167,I448193,);
not I_26215 (I448201,I448193);
nand I_26216 (I448218,I178501,I178501);
and I_26217 (I448235,I448218,I178519);
DFFARX1 I_26218 (I448235,I2507,I448167,I448261,);
DFFARX1 I_26219 (I448261,I2507,I448167,I448156,);
DFFARX1 I_26220 (I178522,I2507,I448167,I448292,);
nand I_26221 (I448300,I448292,I178504);
not I_26222 (I448317,I448300);
DFFARX1 I_26223 (I448317,I2507,I448167,I448343,);
not I_26224 (I448351,I448343);
nor I_26225 (I448159,I448201,I448351);
DFFARX1 I_26226 (I178516,I2507,I448167,I448391,);
nor I_26227 (I448150,I448391,I448261);
nor I_26228 (I448141,I448391,I448317);
nand I_26229 (I448427,I178528,I178507);
and I_26230 (I448444,I448427,I178513);
DFFARX1 I_26231 (I448444,I2507,I448167,I448470,);
not I_26232 (I448478,I448470);
nand I_26233 (I448495,I448478,I448391);
nand I_26234 (I448144,I448478,I448300);
nor I_26235 (I448526,I178525,I178507);
and I_26236 (I448543,I448391,I448526);
nor I_26237 (I448560,I448478,I448543);
DFFARX1 I_26238 (I448560,I2507,I448167,I448153,);
nor I_26239 (I448591,I448193,I448526);
DFFARX1 I_26240 (I448591,I2507,I448167,I448138,);
nor I_26241 (I448622,I448470,I448526);
not I_26242 (I448639,I448622);
nand I_26243 (I448147,I448639,I448495);
not I_26244 (I448694,I2514);
DFFARX1 I_26245 (I392327,I2507,I448694,I448720,);
not I_26246 (I448728,I448720);
nand I_26247 (I448745,I392330,I392327);
and I_26248 (I448762,I448745,I392339);
DFFARX1 I_26249 (I448762,I2507,I448694,I448788,);
DFFARX1 I_26250 (I448788,I2507,I448694,I448683,);
DFFARX1 I_26251 (I392336,I2507,I448694,I448819,);
nand I_26252 (I448827,I448819,I392342);
not I_26253 (I448844,I448827);
DFFARX1 I_26254 (I448844,I2507,I448694,I448870,);
not I_26255 (I448878,I448870);
nor I_26256 (I448686,I448728,I448878);
DFFARX1 I_26257 (I392351,I2507,I448694,I448918,);
nor I_26258 (I448677,I448918,I448788);
nor I_26259 (I448668,I448918,I448844);
nand I_26260 (I448954,I392345,I392333);
and I_26261 (I448971,I448954,I392330);
DFFARX1 I_26262 (I448971,I2507,I448694,I448997,);
not I_26263 (I449005,I448997);
nand I_26264 (I449022,I449005,I448918);
nand I_26265 (I448671,I449005,I448827);
nor I_26266 (I449053,I392348,I392333);
and I_26267 (I449070,I448918,I449053);
nor I_26268 (I449087,I449005,I449070);
DFFARX1 I_26269 (I449087,I2507,I448694,I448680,);
nor I_26270 (I449118,I448720,I449053);
DFFARX1 I_26271 (I449118,I2507,I448694,I448665,);
nor I_26272 (I449149,I448997,I449053);
not I_26273 (I449166,I449149);
nand I_26274 (I448674,I449166,I449022);
not I_26275 (I449221,I2514);
DFFARX1 I_26276 (I366317,I2507,I449221,I449247,);
not I_26277 (I449255,I449247);
nand I_26278 (I449272,I366320,I366317);
and I_26279 (I449289,I449272,I366329);
DFFARX1 I_26280 (I449289,I2507,I449221,I449315,);
DFFARX1 I_26281 (I449315,I2507,I449221,I449210,);
DFFARX1 I_26282 (I366326,I2507,I449221,I449346,);
nand I_26283 (I449354,I449346,I366332);
not I_26284 (I449371,I449354);
DFFARX1 I_26285 (I449371,I2507,I449221,I449397,);
not I_26286 (I449405,I449397);
nor I_26287 (I449213,I449255,I449405);
DFFARX1 I_26288 (I366341,I2507,I449221,I449445,);
nor I_26289 (I449204,I449445,I449315);
nor I_26290 (I449195,I449445,I449371);
nand I_26291 (I449481,I366335,I366323);
and I_26292 (I449498,I449481,I366320);
DFFARX1 I_26293 (I449498,I2507,I449221,I449524,);
not I_26294 (I449532,I449524);
nand I_26295 (I449549,I449532,I449445);
nand I_26296 (I449198,I449532,I449354);
nor I_26297 (I449580,I366338,I366323);
and I_26298 (I449597,I449445,I449580);
nor I_26299 (I449614,I449532,I449597);
DFFARX1 I_26300 (I449614,I2507,I449221,I449207,);
nor I_26301 (I449645,I449247,I449580);
DFFARX1 I_26302 (I449645,I2507,I449221,I449192,);
nor I_26303 (I449676,I449524,I449580);
not I_26304 (I449693,I449676);
nand I_26305 (I449201,I449693,I449549);
not I_26306 (I449748,I2514);
DFFARX1 I_26307 (I143130,I2507,I449748,I449774,);
not I_26308 (I449782,I449774);
nand I_26309 (I449799,I143127,I143145);
and I_26310 (I449816,I449799,I143136);
DFFARX1 I_26311 (I449816,I2507,I449748,I449842,);
DFFARX1 I_26312 (I449842,I2507,I449748,I449737,);
DFFARX1 I_26313 (I143142,I2507,I449748,I449873,);
nand I_26314 (I449881,I449873,I143139);
not I_26315 (I449898,I449881);
DFFARX1 I_26316 (I449898,I2507,I449748,I449924,);
not I_26317 (I449932,I449924);
nor I_26318 (I449740,I449782,I449932);
DFFARX1 I_26319 (I143133,I2507,I449748,I449972,);
nor I_26320 (I449731,I449972,I449842);
nor I_26321 (I449722,I449972,I449898);
nand I_26322 (I450008,I143124,I143148);
and I_26323 (I450025,I450008,I143127);
DFFARX1 I_26324 (I450025,I2507,I449748,I450051,);
not I_26325 (I450059,I450051);
nand I_26326 (I450076,I450059,I449972);
nand I_26327 (I449725,I450059,I449881);
nor I_26328 (I450107,I143124,I143148);
and I_26329 (I450124,I449972,I450107);
nor I_26330 (I450141,I450059,I450124);
DFFARX1 I_26331 (I450141,I2507,I449748,I449734,);
nor I_26332 (I450172,I449774,I450107);
DFFARX1 I_26333 (I450172,I2507,I449748,I449719,);
nor I_26334 (I450203,I450051,I450107);
not I_26335 (I450220,I450203);
nand I_26336 (I449728,I450220,I450076);
not I_26337 (I450275,I2514);
DFFARX1 I_26338 (I194847,I2507,I450275,I450301,);
not I_26339 (I450309,I450301);
nand I_26340 (I450326,I194838,I194838);
and I_26341 (I450343,I450326,I194856);
DFFARX1 I_26342 (I450343,I2507,I450275,I450369,);
DFFARX1 I_26343 (I450369,I2507,I450275,I450264,);
DFFARX1 I_26344 (I194859,I2507,I450275,I450400,);
nand I_26345 (I450408,I450400,I194841);
not I_26346 (I450425,I450408);
DFFARX1 I_26347 (I450425,I2507,I450275,I450451,);
not I_26348 (I450459,I450451);
nor I_26349 (I450267,I450309,I450459);
DFFARX1 I_26350 (I194853,I2507,I450275,I450499,);
nor I_26351 (I450258,I450499,I450369);
nor I_26352 (I450249,I450499,I450425);
nand I_26353 (I450535,I194865,I194844);
and I_26354 (I450552,I450535,I194850);
DFFARX1 I_26355 (I450552,I2507,I450275,I450578,);
not I_26356 (I450586,I450578);
nand I_26357 (I450603,I450586,I450499);
nand I_26358 (I450252,I450586,I450408);
nor I_26359 (I450634,I194862,I194844);
and I_26360 (I450651,I450499,I450634);
nor I_26361 (I450668,I450586,I450651);
DFFARX1 I_26362 (I450668,I2507,I450275,I450261,);
nor I_26363 (I450699,I450301,I450634);
DFFARX1 I_26364 (I450699,I2507,I450275,I450246,);
nor I_26365 (I450730,I450578,I450634);
not I_26366 (I450747,I450730);
nand I_26367 (I450255,I450747,I450603);
not I_26368 (I450802,I2514);
DFFARX1 I_26369 (I216454,I2507,I450802,I450828,);
not I_26370 (I450836,I450828);
nand I_26371 (I450853,I216445,I216445);
and I_26372 (I450870,I450853,I216463);
DFFARX1 I_26373 (I450870,I2507,I450802,I450896,);
DFFARX1 I_26374 (I450896,I2507,I450802,I450791,);
DFFARX1 I_26375 (I216466,I2507,I450802,I450927,);
nand I_26376 (I450935,I450927,I216448);
not I_26377 (I450952,I450935);
DFFARX1 I_26378 (I450952,I2507,I450802,I450978,);
not I_26379 (I450986,I450978);
nor I_26380 (I450794,I450836,I450986);
DFFARX1 I_26381 (I216460,I2507,I450802,I451026,);
nor I_26382 (I450785,I451026,I450896);
nor I_26383 (I450776,I451026,I450952);
nand I_26384 (I451062,I216472,I216451);
and I_26385 (I451079,I451062,I216457);
DFFARX1 I_26386 (I451079,I2507,I450802,I451105,);
not I_26387 (I451113,I451105);
nand I_26388 (I451130,I451113,I451026);
nand I_26389 (I450779,I451113,I450935);
nor I_26390 (I451161,I216469,I216451);
and I_26391 (I451178,I451026,I451161);
nor I_26392 (I451195,I451113,I451178);
DFFARX1 I_26393 (I451195,I2507,I450802,I450788,);
nor I_26394 (I451226,I450828,I451161);
DFFARX1 I_26395 (I451226,I2507,I450802,I450773,);
nor I_26396 (I451257,I451105,I451161);
not I_26397 (I451274,I451257);
nand I_26398 (I450782,I451274,I451130);
not I_26399 (I451329,I2514);
DFFARX1 I_26400 (I717433,I2507,I451329,I451355,);
not I_26401 (I451363,I451355);
nand I_26402 (I451380,I717430,I717439);
and I_26403 (I451397,I451380,I717418);
DFFARX1 I_26404 (I451397,I2507,I451329,I451423,);
DFFARX1 I_26405 (I451423,I2507,I451329,I451318,);
DFFARX1 I_26406 (I717421,I2507,I451329,I451454,);
nand I_26407 (I451462,I451454,I717436);
not I_26408 (I451479,I451462);
DFFARX1 I_26409 (I451479,I2507,I451329,I451505,);
not I_26410 (I451513,I451505);
nor I_26411 (I451321,I451363,I451513);
DFFARX1 I_26412 (I717442,I2507,I451329,I451553,);
nor I_26413 (I451312,I451553,I451423);
nor I_26414 (I451303,I451553,I451479);
nand I_26415 (I451589,I717424,I717445);
and I_26416 (I451606,I451589,I717427);
DFFARX1 I_26417 (I451606,I2507,I451329,I451632,);
not I_26418 (I451640,I451632);
nand I_26419 (I451657,I451640,I451553);
nand I_26420 (I451306,I451640,I451462);
nor I_26421 (I451688,I717418,I717445);
and I_26422 (I451705,I451553,I451688);
nor I_26423 (I451722,I451640,I451705);
DFFARX1 I_26424 (I451722,I2507,I451329,I451315,);
nor I_26425 (I451753,I451355,I451688);
DFFARX1 I_26426 (I451753,I2507,I451329,I451300,);
nor I_26427 (I451784,I451632,I451688);
not I_26428 (I451801,I451784);
nand I_26429 (I451309,I451801,I451657);
not I_26430 (I451856,I2514);
DFFARX1 I_26431 (I21974,I2507,I451856,I451882,);
not I_26432 (I451890,I451882);
nand I_26433 (I451907,I21986,I21989);
and I_26434 (I451924,I451907,I21965);
DFFARX1 I_26435 (I451924,I2507,I451856,I451950,);
DFFARX1 I_26436 (I451950,I2507,I451856,I451845,);
DFFARX1 I_26437 (I21983,I2507,I451856,I451981,);
nand I_26438 (I451989,I451981,I21971);
not I_26439 (I452006,I451989);
DFFARX1 I_26440 (I452006,I2507,I451856,I452032,);
not I_26441 (I452040,I452032);
nor I_26442 (I451848,I451890,I452040);
DFFARX1 I_26443 (I21968,I2507,I451856,I452080,);
nor I_26444 (I451839,I452080,I451950);
nor I_26445 (I451830,I452080,I452006);
nand I_26446 (I452116,I21977,I21968);
and I_26447 (I452133,I452116,I21965);
DFFARX1 I_26448 (I452133,I2507,I451856,I452159,);
not I_26449 (I452167,I452159);
nand I_26450 (I452184,I452167,I452080);
nand I_26451 (I451833,I452167,I451989);
nor I_26452 (I452215,I21980,I21968);
and I_26453 (I452232,I452080,I452215);
nor I_26454 (I452249,I452167,I452232);
DFFARX1 I_26455 (I452249,I2507,I451856,I451842,);
nor I_26456 (I452280,I451882,I452215);
DFFARX1 I_26457 (I452280,I2507,I451856,I451827,);
nor I_26458 (I452311,I452159,I452215);
not I_26459 (I452328,I452311);
nand I_26460 (I451836,I452328,I452184);
not I_26461 (I452383,I2514);
DFFARX1 I_26462 (I586723,I2507,I452383,I452409,);
not I_26463 (I452417,I452409);
nand I_26464 (I452434,I586705,I586705);
and I_26465 (I452451,I452434,I586711);
DFFARX1 I_26466 (I452451,I2507,I452383,I452477,);
DFFARX1 I_26467 (I452477,I2507,I452383,I452372,);
DFFARX1 I_26468 (I586708,I2507,I452383,I452508,);
nand I_26469 (I452516,I452508,I586717);
not I_26470 (I452533,I452516);
DFFARX1 I_26471 (I452533,I2507,I452383,I452559,);
not I_26472 (I452567,I452559);
nor I_26473 (I452375,I452417,I452567);
DFFARX1 I_26474 (I586729,I2507,I452383,I452607,);
nor I_26475 (I452366,I452607,I452477);
nor I_26476 (I452357,I452607,I452533);
nand I_26477 (I452643,I586720,I586714);
and I_26478 (I452660,I452643,I586708);
DFFARX1 I_26479 (I452660,I2507,I452383,I452686,);
not I_26480 (I452694,I452686);
nand I_26481 (I452711,I452694,I452607);
nand I_26482 (I452360,I452694,I452516);
nor I_26483 (I452742,I586726,I586714);
and I_26484 (I452759,I452607,I452742);
nor I_26485 (I452776,I452694,I452759);
DFFARX1 I_26486 (I452776,I2507,I452383,I452369,);
nor I_26487 (I452807,I452409,I452742);
DFFARX1 I_26488 (I452807,I2507,I452383,I452354,);
nor I_26489 (I452838,I452686,I452742);
not I_26490 (I452855,I452838);
nand I_26491 (I452363,I452855,I452711);
not I_26492 (I452910,I2514);
DFFARX1 I_26493 (I377877,I2507,I452910,I452936,);
not I_26494 (I452944,I452936);
nand I_26495 (I452961,I377880,I377877);
and I_26496 (I452978,I452961,I377889);
DFFARX1 I_26497 (I452978,I2507,I452910,I453004,);
DFFARX1 I_26498 (I453004,I2507,I452910,I452899,);
DFFARX1 I_26499 (I377886,I2507,I452910,I453035,);
nand I_26500 (I453043,I453035,I377892);
not I_26501 (I453060,I453043);
DFFARX1 I_26502 (I453060,I2507,I452910,I453086,);
not I_26503 (I453094,I453086);
nor I_26504 (I452902,I452944,I453094);
DFFARX1 I_26505 (I377901,I2507,I452910,I453134,);
nor I_26506 (I452893,I453134,I453004);
nor I_26507 (I452884,I453134,I453060);
nand I_26508 (I453170,I377895,I377883);
and I_26509 (I453187,I453170,I377880);
DFFARX1 I_26510 (I453187,I2507,I452910,I453213,);
not I_26511 (I453221,I453213);
nand I_26512 (I453238,I453221,I453134);
nand I_26513 (I452887,I453221,I453043);
nor I_26514 (I453269,I377898,I377883);
and I_26515 (I453286,I453134,I453269);
nor I_26516 (I453303,I453221,I453286);
DFFARX1 I_26517 (I453303,I2507,I452910,I452896,);
nor I_26518 (I453334,I452936,I453269);
DFFARX1 I_26519 (I453334,I2507,I452910,I452881,);
nor I_26520 (I453365,I453213,I453269);
not I_26521 (I453382,I453365);
nand I_26522 (I452890,I453382,I453238);
not I_26523 (I453437,I2514);
DFFARX1 I_26524 (I676925,I2507,I453437,I453463,);
not I_26525 (I453471,I453463);
nand I_26526 (I453488,I676907,I676910);
and I_26527 (I453505,I453488,I676922);
DFFARX1 I_26528 (I453505,I2507,I453437,I453531,);
DFFARX1 I_26529 (I453531,I2507,I453437,I453426,);
DFFARX1 I_26530 (I676931,I2507,I453437,I453562,);
nand I_26531 (I453570,I453562,I676916);
not I_26532 (I453587,I453570);
DFFARX1 I_26533 (I453587,I2507,I453437,I453613,);
not I_26534 (I453621,I453613);
nor I_26535 (I453429,I453471,I453621);
DFFARX1 I_26536 (I676928,I2507,I453437,I453661,);
nor I_26537 (I453420,I453661,I453531);
nor I_26538 (I453411,I453661,I453587);
nand I_26539 (I453697,I676919,I676913);
and I_26540 (I453714,I453697,I676907);
DFFARX1 I_26541 (I453714,I2507,I453437,I453740,);
not I_26542 (I453748,I453740);
nand I_26543 (I453765,I453748,I453661);
nand I_26544 (I453414,I453748,I453570);
nor I_26545 (I453796,I676910,I676913);
and I_26546 (I453813,I453661,I453796);
nor I_26547 (I453830,I453748,I453813);
DFFARX1 I_26548 (I453830,I2507,I453437,I453423,);
nor I_26549 (I453861,I453463,I453796);
DFFARX1 I_26550 (I453861,I2507,I453437,I453408,);
nor I_26551 (I453892,I453740,I453796);
not I_26552 (I453909,I453892);
nand I_26553 (I453417,I453909,I453765);
not I_26554 (I453964,I2514);
DFFARX1 I_26555 (I385391,I2507,I453964,I453990,);
not I_26556 (I453998,I453990);
nand I_26557 (I454015,I385394,I385391);
and I_26558 (I454032,I454015,I385403);
DFFARX1 I_26559 (I454032,I2507,I453964,I454058,);
DFFARX1 I_26560 (I454058,I2507,I453964,I453953,);
DFFARX1 I_26561 (I385400,I2507,I453964,I454089,);
nand I_26562 (I454097,I454089,I385406);
not I_26563 (I454114,I454097);
DFFARX1 I_26564 (I454114,I2507,I453964,I454140,);
not I_26565 (I454148,I454140);
nor I_26566 (I453956,I453998,I454148);
DFFARX1 I_26567 (I385415,I2507,I453964,I454188,);
nor I_26568 (I453947,I454188,I454058);
nor I_26569 (I453938,I454188,I454114);
nand I_26570 (I454224,I385409,I385397);
and I_26571 (I454241,I454224,I385394);
DFFARX1 I_26572 (I454241,I2507,I453964,I454267,);
not I_26573 (I454275,I454267);
nand I_26574 (I454292,I454275,I454188);
nand I_26575 (I453941,I454275,I454097);
nor I_26576 (I454323,I385412,I385397);
and I_26577 (I454340,I454188,I454323);
nor I_26578 (I454357,I454275,I454340);
DFFARX1 I_26579 (I454357,I2507,I453964,I453950,);
nor I_26580 (I454388,I453990,I454323);
DFFARX1 I_26581 (I454388,I2507,I453964,I453935,);
nor I_26582 (I454419,I454267,I454323);
not I_26583 (I454436,I454419);
nand I_26584 (I453944,I454436,I454292);
not I_26585 (I454491,I2514);
DFFARX1 I_26586 (I69946,I2507,I454491,I454517,);
not I_26587 (I454525,I454517);
nand I_26588 (I454542,I69922,I69931);
and I_26589 (I454559,I454542,I69925);
DFFARX1 I_26590 (I454559,I2507,I454491,I454585,);
DFFARX1 I_26591 (I454585,I2507,I454491,I454480,);
DFFARX1 I_26592 (I69943,I2507,I454491,I454616,);
nand I_26593 (I454624,I454616,I69934);
not I_26594 (I454641,I454624);
DFFARX1 I_26595 (I454641,I2507,I454491,I454667,);
not I_26596 (I454675,I454667);
nor I_26597 (I454483,I454525,I454675);
DFFARX1 I_26598 (I69928,I2507,I454491,I454715,);
nor I_26599 (I454474,I454715,I454585);
nor I_26600 (I454465,I454715,I454641);
nand I_26601 (I454751,I69940,I69937);
and I_26602 (I454768,I454751,I69925);
DFFARX1 I_26603 (I454768,I2507,I454491,I454794,);
not I_26604 (I454802,I454794);
nand I_26605 (I454819,I454802,I454715);
nand I_26606 (I454468,I454802,I454624);
nor I_26607 (I454850,I69922,I69937);
and I_26608 (I454867,I454715,I454850);
nor I_26609 (I454884,I454802,I454867);
DFFARX1 I_26610 (I454884,I2507,I454491,I454477,);
nor I_26611 (I454915,I454517,I454850);
DFFARX1 I_26612 (I454915,I2507,I454491,I454462,);
nor I_26613 (I454946,I454794,I454850);
not I_26614 (I454963,I454946);
nand I_26615 (I454471,I454963,I454819);
not I_26616 (I455018,I2514);
DFFARX1 I_26617 (I27771,I2507,I455018,I455044,);
not I_26618 (I455052,I455044);
nand I_26619 (I455069,I27783,I27786);
and I_26620 (I455086,I455069,I27762);
DFFARX1 I_26621 (I455086,I2507,I455018,I455112,);
DFFARX1 I_26622 (I455112,I2507,I455018,I455007,);
DFFARX1 I_26623 (I27780,I2507,I455018,I455143,);
nand I_26624 (I455151,I455143,I27768);
not I_26625 (I455168,I455151);
DFFARX1 I_26626 (I455168,I2507,I455018,I455194,);
not I_26627 (I455202,I455194);
nor I_26628 (I455010,I455052,I455202);
DFFARX1 I_26629 (I27765,I2507,I455018,I455242,);
nor I_26630 (I455001,I455242,I455112);
nor I_26631 (I454992,I455242,I455168);
nand I_26632 (I455278,I27774,I27765);
and I_26633 (I455295,I455278,I27762);
DFFARX1 I_26634 (I455295,I2507,I455018,I455321,);
not I_26635 (I455329,I455321);
nand I_26636 (I455346,I455329,I455242);
nand I_26637 (I454995,I455329,I455151);
nor I_26638 (I455377,I27777,I27765);
and I_26639 (I455394,I455242,I455377);
nor I_26640 (I455411,I455329,I455394);
DFFARX1 I_26641 (I455411,I2507,I455018,I455004,);
nor I_26642 (I455442,I455044,I455377);
DFFARX1 I_26643 (I455442,I2507,I455018,I454989,);
nor I_26644 (I455473,I455321,I455377);
not I_26645 (I455490,I455473);
nand I_26646 (I454998,I455490,I455346);
not I_26647 (I455545,I2514);
DFFARX1 I_26648 (I205914,I2507,I455545,I455571,);
not I_26649 (I455579,I455571);
nand I_26650 (I455596,I205905,I205905);
and I_26651 (I455613,I455596,I205923);
DFFARX1 I_26652 (I455613,I2507,I455545,I455639,);
DFFARX1 I_26653 (I455639,I2507,I455545,I455534,);
DFFARX1 I_26654 (I205926,I2507,I455545,I455670,);
nand I_26655 (I455678,I455670,I205908);
not I_26656 (I455695,I455678);
DFFARX1 I_26657 (I455695,I2507,I455545,I455721,);
not I_26658 (I455729,I455721);
nor I_26659 (I455537,I455579,I455729);
DFFARX1 I_26660 (I205920,I2507,I455545,I455769,);
nor I_26661 (I455528,I455769,I455639);
nor I_26662 (I455519,I455769,I455695);
nand I_26663 (I455805,I205932,I205911);
and I_26664 (I455822,I455805,I205917);
DFFARX1 I_26665 (I455822,I2507,I455545,I455848,);
not I_26666 (I455856,I455848);
nand I_26667 (I455873,I455856,I455769);
nand I_26668 (I455522,I455856,I455678);
nor I_26669 (I455904,I205929,I205911);
and I_26670 (I455921,I455769,I455904);
nor I_26671 (I455938,I455856,I455921);
DFFARX1 I_26672 (I455938,I2507,I455545,I455531,);
nor I_26673 (I455969,I455571,I455904);
DFFARX1 I_26674 (I455969,I2507,I455545,I455516,);
nor I_26675 (I456000,I455848,I455904);
not I_26676 (I456017,I456000);
nand I_26677 (I455525,I456017,I455873);
not I_26678 (I456072,I2514);
DFFARX1 I_26679 (I416603,I2507,I456072,I456098,);
not I_26680 (I456106,I456098);
nand I_26681 (I456123,I416606,I416603);
and I_26682 (I456140,I456123,I416615);
DFFARX1 I_26683 (I456140,I2507,I456072,I456166,);
DFFARX1 I_26684 (I456166,I2507,I456072,I456061,);
DFFARX1 I_26685 (I416612,I2507,I456072,I456197,);
nand I_26686 (I456205,I456197,I416618);
not I_26687 (I456222,I456205);
DFFARX1 I_26688 (I456222,I2507,I456072,I456248,);
not I_26689 (I456256,I456248);
nor I_26690 (I456064,I456106,I456256);
DFFARX1 I_26691 (I416627,I2507,I456072,I456296,);
nor I_26692 (I456055,I456296,I456166);
nor I_26693 (I456046,I456296,I456222);
nand I_26694 (I456332,I416621,I416609);
and I_26695 (I456349,I456332,I416606);
DFFARX1 I_26696 (I456349,I2507,I456072,I456375,);
not I_26697 (I456383,I456375);
nand I_26698 (I456400,I456383,I456296);
nand I_26699 (I456049,I456383,I456205);
nor I_26700 (I456431,I416624,I416609);
and I_26701 (I456448,I456296,I456431);
nor I_26702 (I456465,I456383,I456448);
DFFARX1 I_26703 (I456465,I2507,I456072,I456058,);
nor I_26704 (I456496,I456098,I456431);
DFFARX1 I_26705 (I456496,I2507,I456072,I456043,);
nor I_26706 (I456527,I456375,I456431);
not I_26707 (I456544,I456527);
nand I_26708 (I456052,I456544,I456400);
not I_26709 (I456599,I2514);
DFFARX1 I_26710 (I68892,I2507,I456599,I456625,);
not I_26711 (I456633,I456625);
nand I_26712 (I456650,I68868,I68877);
and I_26713 (I456667,I456650,I68871);
DFFARX1 I_26714 (I456667,I2507,I456599,I456693,);
DFFARX1 I_26715 (I456693,I2507,I456599,I456588,);
DFFARX1 I_26716 (I68889,I2507,I456599,I456724,);
nand I_26717 (I456732,I456724,I68880);
not I_26718 (I456749,I456732);
DFFARX1 I_26719 (I456749,I2507,I456599,I456775,);
not I_26720 (I456783,I456775);
nor I_26721 (I456591,I456633,I456783);
DFFARX1 I_26722 (I68874,I2507,I456599,I456823,);
nor I_26723 (I456582,I456823,I456693);
nor I_26724 (I456573,I456823,I456749);
nand I_26725 (I456859,I68886,I68883);
and I_26726 (I456876,I456859,I68871);
DFFARX1 I_26727 (I456876,I2507,I456599,I456902,);
not I_26728 (I456910,I456902);
nand I_26729 (I456927,I456910,I456823);
nand I_26730 (I456576,I456910,I456732);
nor I_26731 (I456958,I68868,I68883);
and I_26732 (I456975,I456823,I456958);
nor I_26733 (I456992,I456910,I456975);
DFFARX1 I_26734 (I456992,I2507,I456599,I456585,);
nor I_26735 (I457023,I456625,I456958);
DFFARX1 I_26736 (I457023,I2507,I456599,I456570,);
nor I_26737 (I457054,I456902,I456958);
not I_26738 (I457071,I457054);
nand I_26739 (I456579,I457071,I456927);
not I_26740 (I457126,I2514);
DFFARX1 I_26741 (I193793,I2507,I457126,I457152,);
not I_26742 (I457160,I457152);
nand I_26743 (I457177,I193784,I193784);
and I_26744 (I457194,I457177,I193802);
DFFARX1 I_26745 (I457194,I2507,I457126,I457220,);
DFFARX1 I_26746 (I457220,I2507,I457126,I457115,);
DFFARX1 I_26747 (I193805,I2507,I457126,I457251,);
nand I_26748 (I457259,I457251,I193787);
not I_26749 (I457276,I457259);
DFFARX1 I_26750 (I457276,I2507,I457126,I457302,);
not I_26751 (I457310,I457302);
nor I_26752 (I457118,I457160,I457310);
DFFARX1 I_26753 (I193799,I2507,I457126,I457350,);
nor I_26754 (I457109,I457350,I457220);
nor I_26755 (I457100,I457350,I457276);
nand I_26756 (I457386,I193811,I193790);
and I_26757 (I457403,I457386,I193796);
DFFARX1 I_26758 (I457403,I2507,I457126,I457429,);
not I_26759 (I457437,I457429);
nand I_26760 (I457454,I457437,I457350);
nand I_26761 (I457103,I457437,I457259);
nor I_26762 (I457485,I193808,I193790);
and I_26763 (I457502,I457350,I457485);
nor I_26764 (I457519,I457437,I457502);
DFFARX1 I_26765 (I457519,I2507,I457126,I457112,);
nor I_26766 (I457550,I457152,I457485);
DFFARX1 I_26767 (I457550,I2507,I457126,I457097,);
nor I_26768 (I457581,I457429,I457485);
not I_26769 (I457598,I457581);
nand I_26770 (I457106,I457598,I457454);
not I_26771 (I457653,I2514);
DFFARX1 I_26772 (I621981,I2507,I457653,I457679,);
not I_26773 (I457687,I457679);
nand I_26774 (I457704,I621963,I621963);
and I_26775 (I457721,I457704,I621969);
DFFARX1 I_26776 (I457721,I2507,I457653,I457747,);
DFFARX1 I_26777 (I457747,I2507,I457653,I457642,);
DFFARX1 I_26778 (I621966,I2507,I457653,I457778,);
nand I_26779 (I457786,I457778,I621975);
not I_26780 (I457803,I457786);
DFFARX1 I_26781 (I457803,I2507,I457653,I457829,);
not I_26782 (I457837,I457829);
nor I_26783 (I457645,I457687,I457837);
DFFARX1 I_26784 (I621987,I2507,I457653,I457877,);
nor I_26785 (I457636,I457877,I457747);
nor I_26786 (I457627,I457877,I457803);
nand I_26787 (I457913,I621978,I621972);
and I_26788 (I457930,I457913,I621966);
DFFARX1 I_26789 (I457930,I2507,I457653,I457956,);
not I_26790 (I457964,I457956);
nand I_26791 (I457981,I457964,I457877);
nand I_26792 (I457630,I457964,I457786);
nor I_26793 (I458012,I621984,I621972);
and I_26794 (I458029,I457877,I458012);
nor I_26795 (I458046,I457964,I458029);
DFFARX1 I_26796 (I458046,I2507,I457653,I457639,);
nor I_26797 (I458077,I457679,I458012);
DFFARX1 I_26798 (I458077,I2507,I457653,I457624,);
nor I_26799 (I458108,I457956,I458012);
not I_26800 (I458125,I458108);
nand I_26801 (I457633,I458125,I457981);
not I_26802 (I458180,I2514);
DFFARX1 I_26803 (I593081,I2507,I458180,I458206,);
not I_26804 (I458214,I458206);
nand I_26805 (I458231,I593063,I593063);
and I_26806 (I458248,I458231,I593069);
DFFARX1 I_26807 (I458248,I2507,I458180,I458274,);
DFFARX1 I_26808 (I458274,I2507,I458180,I458169,);
DFFARX1 I_26809 (I593066,I2507,I458180,I458305,);
nand I_26810 (I458313,I458305,I593075);
not I_26811 (I458330,I458313);
DFFARX1 I_26812 (I458330,I2507,I458180,I458356,);
not I_26813 (I458364,I458356);
nor I_26814 (I458172,I458214,I458364);
DFFARX1 I_26815 (I593087,I2507,I458180,I458404,);
nor I_26816 (I458163,I458404,I458274);
nor I_26817 (I458154,I458404,I458330);
nand I_26818 (I458440,I593078,I593072);
and I_26819 (I458457,I458440,I593066);
DFFARX1 I_26820 (I458457,I2507,I458180,I458483,);
not I_26821 (I458491,I458483);
nand I_26822 (I458508,I458491,I458404);
nand I_26823 (I458157,I458491,I458313);
nor I_26824 (I458539,I593084,I593072);
and I_26825 (I458556,I458404,I458539);
nor I_26826 (I458573,I458491,I458556);
DFFARX1 I_26827 (I458573,I2507,I458180,I458166,);
nor I_26828 (I458604,I458206,I458539);
DFFARX1 I_26829 (I458604,I2507,I458180,I458151,);
nor I_26830 (I458635,I458483,I458539);
not I_26831 (I458652,I458635);
nand I_26832 (I458160,I458652,I458508);
not I_26833 (I458707,I2514);
DFFARX1 I_26834 (I175348,I2507,I458707,I458733,);
not I_26835 (I458741,I458733);
nand I_26836 (I458758,I175339,I175339);
and I_26837 (I458775,I458758,I175357);
DFFARX1 I_26838 (I458775,I2507,I458707,I458801,);
DFFARX1 I_26839 (I458801,I2507,I458707,I458696,);
DFFARX1 I_26840 (I175360,I2507,I458707,I458832,);
nand I_26841 (I458840,I458832,I175342);
not I_26842 (I458857,I458840);
DFFARX1 I_26843 (I458857,I2507,I458707,I458883,);
not I_26844 (I458891,I458883);
nor I_26845 (I458699,I458741,I458891);
DFFARX1 I_26846 (I175354,I2507,I458707,I458931,);
nor I_26847 (I458690,I458931,I458801);
nor I_26848 (I458681,I458931,I458857);
nand I_26849 (I458967,I175366,I175345);
and I_26850 (I458984,I458967,I175351);
DFFARX1 I_26851 (I458984,I2507,I458707,I459010,);
not I_26852 (I459018,I459010);
nand I_26853 (I459035,I459018,I458931);
nand I_26854 (I458684,I459018,I458840);
nor I_26855 (I459066,I175363,I175345);
and I_26856 (I459083,I458931,I459066);
nor I_26857 (I459100,I459018,I459083);
DFFARX1 I_26858 (I459100,I2507,I458707,I458693,);
nor I_26859 (I459131,I458733,I459066);
DFFARX1 I_26860 (I459131,I2507,I458707,I458678,);
nor I_26861 (I459162,I459010,I459066);
not I_26862 (I459179,I459162);
nand I_26863 (I458687,I459179,I459035);
not I_26864 (I459234,I2514);
DFFARX1 I_26865 (I343790,I2507,I459234,I459260,);
not I_26866 (I459268,I459260);
nand I_26867 (I459285,I343775,I343796);
and I_26868 (I459302,I459285,I343784);
DFFARX1 I_26869 (I459302,I2507,I459234,I459328,);
DFFARX1 I_26870 (I459328,I2507,I459234,I459223,);
DFFARX1 I_26871 (I343778,I2507,I459234,I459359,);
nand I_26872 (I459367,I459359,I343787);
not I_26873 (I459384,I459367);
DFFARX1 I_26874 (I459384,I2507,I459234,I459410,);
not I_26875 (I459418,I459410);
nor I_26876 (I459226,I459268,I459418);
DFFARX1 I_26877 (I343793,I2507,I459234,I459458,);
nor I_26878 (I459217,I459458,I459328);
nor I_26879 (I459208,I459458,I459384);
nand I_26880 (I459494,I343775,I343778);
and I_26881 (I459511,I459494,I343799);
DFFARX1 I_26882 (I459511,I2507,I459234,I459537,);
not I_26883 (I459545,I459537);
nand I_26884 (I459562,I459545,I459458);
nand I_26885 (I459211,I459545,I459367);
nor I_26886 (I459593,I343781,I343778);
and I_26887 (I459610,I459458,I459593);
nor I_26888 (I459627,I459545,I459610);
DFFARX1 I_26889 (I459627,I2507,I459234,I459220,);
nor I_26890 (I459658,I459260,I459593);
DFFARX1 I_26891 (I459658,I2507,I459234,I459205,);
nor I_26892 (I459689,I459537,I459593);
not I_26893 (I459706,I459689);
nand I_26894 (I459214,I459706,I459562);
not I_26895 (I459761,I2514);
DFFARX1 I_26896 (I114570,I2507,I459761,I459787,);
not I_26897 (I459795,I459787);
nand I_26898 (I459812,I114567,I114585);
and I_26899 (I459829,I459812,I114576);
DFFARX1 I_26900 (I459829,I2507,I459761,I459855,);
DFFARX1 I_26901 (I459855,I2507,I459761,I459750,);
DFFARX1 I_26902 (I114582,I2507,I459761,I459886,);
nand I_26903 (I459894,I459886,I114579);
not I_26904 (I459911,I459894);
DFFARX1 I_26905 (I459911,I2507,I459761,I459937,);
not I_26906 (I459945,I459937);
nor I_26907 (I459753,I459795,I459945);
DFFARX1 I_26908 (I114573,I2507,I459761,I459985,);
nor I_26909 (I459744,I459985,I459855);
nor I_26910 (I459735,I459985,I459911);
nand I_26911 (I460021,I114564,I114588);
and I_26912 (I460038,I460021,I114567);
DFFARX1 I_26913 (I460038,I2507,I459761,I460064,);
not I_26914 (I460072,I460064);
nand I_26915 (I460089,I460072,I459985);
nand I_26916 (I459738,I460072,I459894);
nor I_26917 (I460120,I114564,I114588);
and I_26918 (I460137,I459985,I460120);
nor I_26919 (I460154,I460072,I460137);
DFFARX1 I_26920 (I460154,I2507,I459761,I459747,);
nor I_26921 (I460185,I459787,I460120);
DFFARX1 I_26922 (I460185,I2507,I459761,I459732,);
nor I_26923 (I460216,I460064,I460120);
not I_26924 (I460233,I460216);
nand I_26925 (I459741,I460233,I460089);
not I_26926 (I460288,I2514);
DFFARX1 I_26927 (I99100,I2507,I460288,I460314,);
not I_26928 (I460322,I460314);
nand I_26929 (I460339,I99097,I99115);
and I_26930 (I460356,I460339,I99106);
DFFARX1 I_26931 (I460356,I2507,I460288,I460382,);
DFFARX1 I_26932 (I460382,I2507,I460288,I460277,);
DFFARX1 I_26933 (I99112,I2507,I460288,I460413,);
nand I_26934 (I460421,I460413,I99109);
not I_26935 (I460438,I460421);
DFFARX1 I_26936 (I460438,I2507,I460288,I460464,);
not I_26937 (I460472,I460464);
nor I_26938 (I460280,I460322,I460472);
DFFARX1 I_26939 (I99103,I2507,I460288,I460512,);
nor I_26940 (I460271,I460512,I460382);
nor I_26941 (I460262,I460512,I460438);
nand I_26942 (I460548,I99094,I99118);
and I_26943 (I460565,I460548,I99097);
DFFARX1 I_26944 (I460565,I2507,I460288,I460591,);
not I_26945 (I460599,I460591);
nand I_26946 (I460616,I460599,I460512);
nand I_26947 (I460265,I460599,I460421);
nor I_26948 (I460647,I99094,I99118);
and I_26949 (I460664,I460512,I460647);
nor I_26950 (I460681,I460599,I460664);
DFFARX1 I_26951 (I460681,I2507,I460288,I460274,);
nor I_26952 (I460712,I460314,I460647);
DFFARX1 I_26953 (I460712,I2507,I460288,I460259,);
nor I_26954 (I460743,I460591,I460647);
not I_26955 (I460760,I460743);
nand I_26956 (I460268,I460760,I460616);
not I_26957 (I460815,I2514);
DFFARX1 I_26958 (I518997,I2507,I460815,I460841,);
not I_26959 (I460849,I460841);
nand I_26960 (I460866,I519012,I518994);
and I_26961 (I460883,I460866,I518994);
DFFARX1 I_26962 (I460883,I2507,I460815,I460909,);
DFFARX1 I_26963 (I460909,I2507,I460815,I460804,);
DFFARX1 I_26964 (I519003,I2507,I460815,I460940,);
nand I_26965 (I460948,I460940,I519021);
not I_26966 (I460965,I460948);
DFFARX1 I_26967 (I460965,I2507,I460815,I460991,);
not I_26968 (I460999,I460991);
nor I_26969 (I460807,I460849,I460999);
DFFARX1 I_26970 (I519018,I2507,I460815,I461039,);
nor I_26971 (I460798,I461039,I460909);
nor I_26972 (I460789,I461039,I460965);
nand I_26973 (I461075,I519015,I519006);
and I_26974 (I461092,I461075,I519000);
DFFARX1 I_26975 (I461092,I2507,I460815,I461118,);
not I_26976 (I461126,I461118);
nand I_26977 (I461143,I461126,I461039);
nand I_26978 (I460792,I461126,I460948);
nor I_26979 (I461174,I519009,I519006);
and I_26980 (I461191,I461039,I461174);
nor I_26981 (I461208,I461126,I461191);
DFFARX1 I_26982 (I461208,I2507,I460815,I460801,);
nor I_26983 (I461239,I460841,I461174);
DFFARX1 I_26984 (I461239,I2507,I460815,I460786,);
nor I_26985 (I461270,I461118,I461174);
not I_26986 (I461287,I461270);
nand I_26987 (I460795,I461287,I461143);
not I_26988 (I461342,I2514);
DFFARX1 I_26989 (I284944,I2507,I461342,I461368,);
not I_26990 (I461376,I461368);
nand I_26991 (I461393,I284962,I284953);
and I_26992 (I461410,I461393,I284956);
DFFARX1 I_26993 (I461410,I2507,I461342,I461436,);
DFFARX1 I_26994 (I461436,I2507,I461342,I461331,);
DFFARX1 I_26995 (I284950,I2507,I461342,I461467,);
nand I_26996 (I461475,I461467,I284941);
not I_26997 (I461492,I461475);
DFFARX1 I_26998 (I461492,I2507,I461342,I461518,);
not I_26999 (I461526,I461518);
nor I_27000 (I461334,I461376,I461526);
DFFARX1 I_27001 (I284947,I2507,I461342,I461566,);
nor I_27002 (I461325,I461566,I461436);
nor I_27003 (I461316,I461566,I461492);
nand I_27004 (I461602,I284941,I284938);
and I_27005 (I461619,I461602,I284959);
DFFARX1 I_27006 (I461619,I2507,I461342,I461645,);
not I_27007 (I461653,I461645);
nand I_27008 (I461670,I461653,I461566);
nand I_27009 (I461319,I461653,I461475);
nor I_27010 (I461701,I284938,I284938);
and I_27011 (I461718,I461566,I461701);
nor I_27012 (I461735,I461653,I461718);
DFFARX1 I_27013 (I461735,I2507,I461342,I461328,);
nor I_27014 (I461766,I461368,I461701);
DFFARX1 I_27015 (I461766,I2507,I461342,I461313,);
nor I_27016 (I461797,I461645,I461701);
not I_27017 (I461814,I461797);
nand I_27018 (I461322,I461814,I461670);
not I_27019 (I461869,I2514);
DFFARX1 I_27020 (I349555,I2507,I461869,I461895,);
not I_27021 (I461903,I461895);
nand I_27022 (I461920,I349558,I349555);
and I_27023 (I461937,I461920,I349567);
DFFARX1 I_27024 (I461937,I2507,I461869,I461963,);
DFFARX1 I_27025 (I461963,I2507,I461869,I461858,);
DFFARX1 I_27026 (I349564,I2507,I461869,I461994,);
nand I_27027 (I462002,I461994,I349570);
not I_27028 (I462019,I462002);
DFFARX1 I_27029 (I462019,I2507,I461869,I462045,);
not I_27030 (I462053,I462045);
nor I_27031 (I461861,I461903,I462053);
DFFARX1 I_27032 (I349579,I2507,I461869,I462093,);
nor I_27033 (I461852,I462093,I461963);
nor I_27034 (I461843,I462093,I462019);
nand I_27035 (I462129,I349573,I349561);
and I_27036 (I462146,I462129,I349558);
DFFARX1 I_27037 (I462146,I2507,I461869,I462172,);
not I_27038 (I462180,I462172);
nand I_27039 (I462197,I462180,I462093);
nand I_27040 (I461846,I462180,I462002);
nor I_27041 (I462228,I349576,I349561);
and I_27042 (I462245,I462093,I462228);
nor I_27043 (I462262,I462180,I462245);
DFFARX1 I_27044 (I462262,I2507,I461869,I461855,);
nor I_27045 (I462293,I461895,I462228);
DFFARX1 I_27046 (I462293,I2507,I461869,I461840,);
nor I_27047 (I462324,I462172,I462228);
not I_27048 (I462341,I462324);
nand I_27049 (I461849,I462341,I462197);
not I_27050 (I462396,I2514);
DFFARX1 I_27051 (I508661,I2507,I462396,I462422,);
not I_27052 (I462430,I462422);
nand I_27053 (I462447,I508676,I508658);
and I_27054 (I462464,I462447,I508658);
DFFARX1 I_27055 (I462464,I2507,I462396,I462490,);
DFFARX1 I_27056 (I462490,I2507,I462396,I462385,);
DFFARX1 I_27057 (I508667,I2507,I462396,I462521,);
nand I_27058 (I462529,I462521,I508685);
not I_27059 (I462546,I462529);
DFFARX1 I_27060 (I462546,I2507,I462396,I462572,);
not I_27061 (I462580,I462572);
nor I_27062 (I462388,I462430,I462580);
DFFARX1 I_27063 (I508682,I2507,I462396,I462620,);
nor I_27064 (I462379,I462620,I462490);
nor I_27065 (I462370,I462620,I462546);
nand I_27066 (I462656,I508679,I508670);
and I_27067 (I462673,I462656,I508664);
DFFARX1 I_27068 (I462673,I2507,I462396,I462699,);
not I_27069 (I462707,I462699);
nand I_27070 (I462724,I462707,I462620);
nand I_27071 (I462373,I462707,I462529);
nor I_27072 (I462755,I508673,I508670);
and I_27073 (I462772,I462620,I462755);
nor I_27074 (I462789,I462707,I462772);
DFFARX1 I_27075 (I462789,I2507,I462396,I462382,);
nor I_27076 (I462820,I462422,I462755);
DFFARX1 I_27077 (I462820,I2507,I462396,I462367,);
nor I_27078 (I462851,I462699,I462755);
not I_27079 (I462868,I462851);
nand I_27080 (I462376,I462868,I462724);
not I_27081 (I462923,I2514);
DFFARX1 I_27082 (I284349,I2507,I462923,I462949,);
not I_27083 (I462957,I462949);
nand I_27084 (I462974,I284367,I284358);
and I_27085 (I462991,I462974,I284361);
DFFARX1 I_27086 (I462991,I2507,I462923,I463017,);
DFFARX1 I_27087 (I463017,I2507,I462923,I462912,);
DFFARX1 I_27088 (I284355,I2507,I462923,I463048,);
nand I_27089 (I463056,I463048,I284346);
not I_27090 (I463073,I463056);
DFFARX1 I_27091 (I463073,I2507,I462923,I463099,);
not I_27092 (I463107,I463099);
nor I_27093 (I462915,I462957,I463107);
DFFARX1 I_27094 (I284352,I2507,I462923,I463147,);
nor I_27095 (I462906,I463147,I463017);
nor I_27096 (I462897,I463147,I463073);
nand I_27097 (I463183,I284346,I284343);
and I_27098 (I463200,I463183,I284364);
DFFARX1 I_27099 (I463200,I2507,I462923,I463226,);
not I_27100 (I463234,I463226);
nand I_27101 (I463251,I463234,I463147);
nand I_27102 (I462900,I463234,I463056);
nor I_27103 (I463282,I284343,I284343);
and I_27104 (I463299,I463147,I463282);
nor I_27105 (I463316,I463234,I463299);
DFFARX1 I_27106 (I463316,I2507,I462923,I462909,);
nor I_27107 (I463347,I462949,I463282);
DFFARX1 I_27108 (I463347,I2507,I462923,I462894,);
nor I_27109 (I463378,I463226,I463282);
not I_27110 (I463395,I463378);
nand I_27111 (I462903,I463395,I463251);
not I_27112 (I463450,I2514);
DFFARX1 I_27113 (I318358,I2507,I463450,I463476,);
not I_27114 (I463484,I463476);
nand I_27115 (I463501,I318343,I318364);
and I_27116 (I463518,I463501,I318352);
DFFARX1 I_27117 (I463518,I2507,I463450,I463544,);
DFFARX1 I_27118 (I463544,I2507,I463450,I463439,);
DFFARX1 I_27119 (I318346,I2507,I463450,I463575,);
nand I_27120 (I463583,I463575,I318355);
not I_27121 (I463600,I463583);
DFFARX1 I_27122 (I463600,I2507,I463450,I463626,);
not I_27123 (I463634,I463626);
nor I_27124 (I463442,I463484,I463634);
DFFARX1 I_27125 (I318361,I2507,I463450,I463674,);
nor I_27126 (I463433,I463674,I463544);
nor I_27127 (I463424,I463674,I463600);
nand I_27128 (I463710,I318343,I318346);
and I_27129 (I463727,I463710,I318367);
DFFARX1 I_27130 (I463727,I2507,I463450,I463753,);
not I_27131 (I463761,I463753);
nand I_27132 (I463778,I463761,I463674);
nand I_27133 (I463427,I463761,I463583);
nor I_27134 (I463809,I318349,I318346);
and I_27135 (I463826,I463674,I463809);
nor I_27136 (I463843,I463761,I463826);
DFFARX1 I_27137 (I463843,I2507,I463450,I463436,);
nor I_27138 (I463874,I463476,I463809);
DFFARX1 I_27139 (I463874,I2507,I463450,I463421,);
nor I_27140 (I463905,I463753,I463809);
not I_27141 (I463922,I463905);
nand I_27142 (I463430,I463922,I463778);
not I_27143 (I463977,I2514);
DFFARX1 I_27144 (I107430,I2507,I463977,I464003,);
not I_27145 (I464011,I464003);
nand I_27146 (I464028,I107427,I107445);
and I_27147 (I464045,I464028,I107436);
DFFARX1 I_27148 (I464045,I2507,I463977,I464071,);
DFFARX1 I_27149 (I464071,I2507,I463977,I463966,);
DFFARX1 I_27150 (I107442,I2507,I463977,I464102,);
nand I_27151 (I464110,I464102,I107439);
not I_27152 (I464127,I464110);
DFFARX1 I_27153 (I464127,I2507,I463977,I464153,);
not I_27154 (I464161,I464153);
nor I_27155 (I463969,I464011,I464161);
DFFARX1 I_27156 (I107433,I2507,I463977,I464201,);
nor I_27157 (I463960,I464201,I464071);
nor I_27158 (I463951,I464201,I464127);
nand I_27159 (I464237,I107424,I107448);
and I_27160 (I464254,I464237,I107427);
DFFARX1 I_27161 (I464254,I2507,I463977,I464280,);
not I_27162 (I464288,I464280);
nand I_27163 (I464305,I464288,I464201);
nand I_27164 (I463954,I464288,I464110);
nor I_27165 (I464336,I107424,I107448);
and I_27166 (I464353,I464201,I464336);
nor I_27167 (I464370,I464288,I464353);
DFFARX1 I_27168 (I464370,I2507,I463977,I463963,);
nor I_27169 (I464401,I464003,I464336);
DFFARX1 I_27170 (I464401,I2507,I463977,I463948,);
nor I_27171 (I464432,I464280,I464336);
not I_27172 (I464449,I464432);
nand I_27173 (I463957,I464449,I464305);
not I_27174 (I464504,I2514);
DFFARX1 I_27175 (I644721,I2507,I464504,I464530,);
not I_27176 (I464538,I464530);
nand I_27177 (I464555,I644727,I644709);
and I_27178 (I464572,I464555,I644718);
DFFARX1 I_27179 (I464572,I2507,I464504,I464598,);
DFFARX1 I_27180 (I464598,I2507,I464504,I464493,);
DFFARX1 I_27181 (I644724,I2507,I464504,I464629,);
nand I_27182 (I464637,I464629,I644712);
not I_27183 (I464654,I464637);
DFFARX1 I_27184 (I464654,I2507,I464504,I464680,);
not I_27185 (I464688,I464680);
nor I_27186 (I464496,I464538,I464688);
DFFARX1 I_27187 (I644730,I2507,I464504,I464728,);
nor I_27188 (I464487,I464728,I464598);
nor I_27189 (I464478,I464728,I464654);
nand I_27190 (I464764,I644709,I644715);
and I_27191 (I464781,I464764,I644733);
DFFARX1 I_27192 (I464781,I2507,I464504,I464807,);
not I_27193 (I464815,I464807);
nand I_27194 (I464832,I464815,I464728);
nand I_27195 (I464481,I464815,I464637);
nor I_27196 (I464863,I644712,I644715);
and I_27197 (I464880,I464728,I464863);
nor I_27198 (I464897,I464815,I464880);
DFFARX1 I_27199 (I464897,I2507,I464504,I464490,);
nor I_27200 (I464928,I464530,I464863);
DFFARX1 I_27201 (I464928,I2507,I464504,I464475,);
nor I_27202 (I464959,I464807,I464863);
not I_27203 (I464976,I464959);
nand I_27204 (I464484,I464976,I464832);
not I_27205 (I465031,I2514);
DFFARX1 I_27206 (I303908,I2507,I465031,I465057,);
not I_27207 (I465065,I465057);
nand I_27208 (I465082,I303893,I303914);
and I_27209 (I465099,I465082,I303902);
DFFARX1 I_27210 (I465099,I2507,I465031,I465125,);
DFFARX1 I_27211 (I465125,I2507,I465031,I465020,);
DFFARX1 I_27212 (I303896,I2507,I465031,I465156,);
nand I_27213 (I465164,I465156,I303905);
not I_27214 (I465181,I465164);
DFFARX1 I_27215 (I465181,I2507,I465031,I465207,);
not I_27216 (I465215,I465207);
nor I_27217 (I465023,I465065,I465215);
DFFARX1 I_27218 (I303911,I2507,I465031,I465255,);
nor I_27219 (I465014,I465255,I465125);
nor I_27220 (I465005,I465255,I465181);
nand I_27221 (I465291,I303893,I303896);
and I_27222 (I465308,I465291,I303917);
DFFARX1 I_27223 (I465308,I2507,I465031,I465334,);
not I_27224 (I465342,I465334);
nand I_27225 (I465359,I465342,I465255);
nand I_27226 (I465008,I465342,I465164);
nor I_27227 (I465390,I303899,I303896);
and I_27228 (I465407,I465255,I465390);
nor I_27229 (I465424,I465342,I465407);
DFFARX1 I_27230 (I465424,I2507,I465031,I465017,);
nor I_27231 (I465455,I465057,I465390);
DFFARX1 I_27232 (I465455,I2507,I465031,I465002,);
nor I_27233 (I465486,I465334,I465390);
not I_27234 (I465503,I465486);
nand I_27235 (I465011,I465503,I465359);
not I_27236 (I465558,I2514);
DFFARX1 I_27237 (I164808,I2507,I465558,I465584,);
not I_27238 (I465592,I465584);
nand I_27239 (I465609,I164799,I164799);
and I_27240 (I465626,I465609,I164817);
DFFARX1 I_27241 (I465626,I2507,I465558,I465652,);
DFFARX1 I_27242 (I465652,I2507,I465558,I465547,);
DFFARX1 I_27243 (I164820,I2507,I465558,I465683,);
nand I_27244 (I465691,I465683,I164802);
not I_27245 (I465708,I465691);
DFFARX1 I_27246 (I465708,I2507,I465558,I465734,);
not I_27247 (I465742,I465734);
nor I_27248 (I465550,I465592,I465742);
DFFARX1 I_27249 (I164814,I2507,I465558,I465782,);
nor I_27250 (I465541,I465782,I465652);
nor I_27251 (I465532,I465782,I465708);
nand I_27252 (I465818,I164826,I164805);
and I_27253 (I465835,I465818,I164811);
DFFARX1 I_27254 (I465835,I2507,I465558,I465861,);
not I_27255 (I465869,I465861);
nand I_27256 (I465886,I465869,I465782);
nand I_27257 (I465535,I465869,I465691);
nor I_27258 (I465917,I164823,I164805);
and I_27259 (I465934,I465782,I465917);
nor I_27260 (I465951,I465869,I465934);
DFFARX1 I_27261 (I465951,I2507,I465558,I465544,);
nor I_27262 (I465982,I465584,I465917);
DFFARX1 I_27263 (I465982,I2507,I465558,I465529,);
nor I_27264 (I466013,I465861,I465917);
not I_27265 (I466030,I466013);
nand I_27266 (I465538,I466030,I465886);
not I_27267 (I466085,I2514);
DFFARX1 I_27268 (I335120,I2507,I466085,I466111,);
not I_27269 (I466119,I466111);
nand I_27270 (I466136,I335105,I335126);
and I_27271 (I466153,I466136,I335114);
DFFARX1 I_27272 (I466153,I2507,I466085,I466179,);
DFFARX1 I_27273 (I466179,I2507,I466085,I466074,);
DFFARX1 I_27274 (I335108,I2507,I466085,I466210,);
nand I_27275 (I466218,I466210,I335117);
not I_27276 (I466235,I466218);
DFFARX1 I_27277 (I466235,I2507,I466085,I466261,);
not I_27278 (I466269,I466261);
nor I_27279 (I466077,I466119,I466269);
DFFARX1 I_27280 (I335123,I2507,I466085,I466309,);
nor I_27281 (I466068,I466309,I466179);
nor I_27282 (I466059,I466309,I466235);
nand I_27283 (I466345,I335105,I335108);
and I_27284 (I466362,I466345,I335129);
DFFARX1 I_27285 (I466362,I2507,I466085,I466388,);
not I_27286 (I466396,I466388);
nand I_27287 (I466413,I466396,I466309);
nand I_27288 (I466062,I466396,I466218);
nor I_27289 (I466444,I335111,I335108);
and I_27290 (I466461,I466309,I466444);
nor I_27291 (I466478,I466396,I466461);
DFFARX1 I_27292 (I466478,I2507,I466085,I466071,);
nor I_27293 (I466509,I466111,I466444);
DFFARX1 I_27294 (I466509,I2507,I466085,I466056,);
nor I_27295 (I466540,I466388,I466444);
not I_27296 (I466557,I466540);
nand I_27297 (I466065,I466557,I466413);
not I_27298 (I466612,I2514);
DFFARX1 I_27299 (I707913,I2507,I466612,I466638,);
not I_27300 (I466646,I466638);
nand I_27301 (I466663,I707910,I707919);
and I_27302 (I466680,I466663,I707898);
DFFARX1 I_27303 (I466680,I2507,I466612,I466706,);
DFFARX1 I_27304 (I466706,I2507,I466612,I466601,);
DFFARX1 I_27305 (I707901,I2507,I466612,I466737,);
nand I_27306 (I466745,I466737,I707916);
not I_27307 (I466762,I466745);
DFFARX1 I_27308 (I466762,I2507,I466612,I466788,);
not I_27309 (I466796,I466788);
nor I_27310 (I466604,I466646,I466796);
DFFARX1 I_27311 (I707922,I2507,I466612,I466836,);
nor I_27312 (I466595,I466836,I466706);
nor I_27313 (I466586,I466836,I466762);
nand I_27314 (I466872,I707904,I707925);
and I_27315 (I466889,I466872,I707907);
DFFARX1 I_27316 (I466889,I2507,I466612,I466915,);
not I_27317 (I466923,I466915);
nand I_27318 (I466940,I466923,I466836);
nand I_27319 (I466589,I466923,I466745);
nor I_27320 (I466971,I707898,I707925);
and I_27321 (I466988,I466836,I466971);
nor I_27322 (I467005,I466923,I466988);
DFFARX1 I_27323 (I467005,I2507,I466612,I466598,);
nor I_27324 (I467036,I466638,I466971);
DFFARX1 I_27325 (I467036,I2507,I466612,I466583,);
nor I_27326 (I467067,I466915,I466971);
not I_27327 (I467084,I467067);
nand I_27328 (I466592,I467084,I466940);
not I_27329 (I467139,I2514);
DFFARX1 I_27330 (I382501,I2507,I467139,I467165,);
not I_27331 (I467173,I467165);
nand I_27332 (I467190,I382504,I382501);
and I_27333 (I467207,I467190,I382513);
DFFARX1 I_27334 (I467207,I2507,I467139,I467233,);
DFFARX1 I_27335 (I467233,I2507,I467139,I467128,);
DFFARX1 I_27336 (I382510,I2507,I467139,I467264,);
nand I_27337 (I467272,I467264,I382516);
not I_27338 (I467289,I467272);
DFFARX1 I_27339 (I467289,I2507,I467139,I467315,);
not I_27340 (I467323,I467315);
nor I_27341 (I467131,I467173,I467323);
DFFARX1 I_27342 (I382525,I2507,I467139,I467363,);
nor I_27343 (I467122,I467363,I467233);
nor I_27344 (I467113,I467363,I467289);
nand I_27345 (I467399,I382519,I382507);
and I_27346 (I467416,I467399,I382504);
DFFARX1 I_27347 (I467416,I2507,I467139,I467442,);
not I_27348 (I467450,I467442);
nand I_27349 (I467467,I467450,I467363);
nand I_27350 (I467116,I467450,I467272);
nor I_27351 (I467498,I382522,I382507);
and I_27352 (I467515,I467363,I467498);
nor I_27353 (I467532,I467450,I467515);
DFFARX1 I_27354 (I467532,I2507,I467139,I467125,);
nor I_27355 (I467563,I467165,I467498);
DFFARX1 I_27356 (I467563,I2507,I467139,I467110,);
nor I_27357 (I467594,I467442,I467498);
not I_27358 (I467611,I467594);
nand I_27359 (I467119,I467611,I467467);
not I_27360 (I467666,I2514);
DFFARX1 I_27361 (I484759,I2507,I467666,I467692,);
not I_27362 (I467700,I467692);
nand I_27363 (I467717,I484774,I484756);
and I_27364 (I467734,I467717,I484756);
DFFARX1 I_27365 (I467734,I2507,I467666,I467760,);
DFFARX1 I_27366 (I467760,I2507,I467666,I467655,);
DFFARX1 I_27367 (I484765,I2507,I467666,I467791,);
nand I_27368 (I467799,I467791,I484783);
not I_27369 (I467816,I467799);
DFFARX1 I_27370 (I467816,I2507,I467666,I467842,);
not I_27371 (I467850,I467842);
nor I_27372 (I467658,I467700,I467850);
DFFARX1 I_27373 (I484780,I2507,I467666,I467890,);
nor I_27374 (I467649,I467890,I467760);
nor I_27375 (I467640,I467890,I467816);
nand I_27376 (I467926,I484777,I484768);
and I_27377 (I467943,I467926,I484762);
DFFARX1 I_27378 (I467943,I2507,I467666,I467969,);
not I_27379 (I467977,I467969);
nand I_27380 (I467994,I467977,I467890);
nand I_27381 (I467643,I467977,I467799);
nor I_27382 (I468025,I484771,I484768);
and I_27383 (I468042,I467890,I468025);
nor I_27384 (I468059,I467977,I468042);
DFFARX1 I_27385 (I468059,I2507,I467666,I467652,);
nor I_27386 (I468090,I467692,I468025);
DFFARX1 I_27387 (I468090,I2507,I467666,I467637,);
nor I_27388 (I468121,I467969,I468025);
not I_27389 (I468138,I468121);
nand I_27390 (I467646,I468138,I467994);
not I_27391 (I468193,I2514);
DFFARX1 I_27392 (I50447,I2507,I468193,I468219,);
not I_27393 (I468227,I468219);
nand I_27394 (I468244,I50423,I50432);
and I_27395 (I468261,I468244,I50426);
DFFARX1 I_27396 (I468261,I2507,I468193,I468287,);
DFFARX1 I_27397 (I468287,I2507,I468193,I468182,);
DFFARX1 I_27398 (I50444,I2507,I468193,I468318,);
nand I_27399 (I468326,I468318,I50435);
not I_27400 (I468343,I468326);
DFFARX1 I_27401 (I468343,I2507,I468193,I468369,);
not I_27402 (I468377,I468369);
nor I_27403 (I468185,I468227,I468377);
DFFARX1 I_27404 (I50429,I2507,I468193,I468417,);
nor I_27405 (I468176,I468417,I468287);
nor I_27406 (I468167,I468417,I468343);
nand I_27407 (I468453,I50441,I50438);
and I_27408 (I468470,I468453,I50426);
DFFARX1 I_27409 (I468470,I2507,I468193,I468496,);
not I_27410 (I468504,I468496);
nand I_27411 (I468521,I468504,I468417);
nand I_27412 (I468170,I468504,I468326);
nor I_27413 (I468552,I50423,I50438);
and I_27414 (I468569,I468417,I468552);
nor I_27415 (I468586,I468504,I468569);
DFFARX1 I_27416 (I468586,I2507,I468193,I468179,);
nor I_27417 (I468617,I468219,I468552);
DFFARX1 I_27418 (I468617,I2507,I468193,I468164,);
nor I_27419 (I468648,I468496,I468552);
not I_27420 (I468665,I468648);
nand I_27421 (I468173,I468665,I468521);
not I_27422 (I468720,I2514);
DFFARX1 I_27423 (I265598,I2507,I468720,I468746,);
not I_27424 (I468754,I468746);
nand I_27425 (I468771,I265595,I265604);
and I_27426 (I468788,I468771,I265613);
DFFARX1 I_27427 (I468788,I2507,I468720,I468814,);
DFFARX1 I_27428 (I468814,I2507,I468720,I468709,);
DFFARX1 I_27429 (I265616,I2507,I468720,I468845,);
nand I_27430 (I468853,I468845,I265619);
not I_27431 (I468870,I468853);
DFFARX1 I_27432 (I468870,I2507,I468720,I468896,);
not I_27433 (I468904,I468896);
nor I_27434 (I468712,I468754,I468904);
DFFARX1 I_27435 (I265592,I2507,I468720,I468944,);
nor I_27436 (I468703,I468944,I468814);
nor I_27437 (I468694,I468944,I468870);
nand I_27438 (I468980,I265607,I265610);
and I_27439 (I468997,I468980,I265601);
DFFARX1 I_27440 (I468997,I2507,I468720,I469023,);
not I_27441 (I469031,I469023);
nand I_27442 (I469048,I469031,I468944);
nand I_27443 (I468697,I469031,I468853);
nor I_27444 (I469079,I265592,I265610);
and I_27445 (I469096,I468944,I469079);
nor I_27446 (I469113,I469031,I469096);
DFFARX1 I_27447 (I469113,I2507,I468720,I468706,);
nor I_27448 (I469144,I468746,I469079);
DFFARX1 I_27449 (I469144,I2507,I468720,I468691,);
nor I_27450 (I469175,I469023,I469079);
not I_27451 (I469192,I469175);
nand I_27452 (I468700,I469192,I469048);
not I_27453 (I469247,I2514);
DFFARX1 I_27454 (I690063,I2507,I469247,I469273,);
not I_27455 (I469281,I469273);
nand I_27456 (I469298,I690060,I690069);
and I_27457 (I469315,I469298,I690048);
DFFARX1 I_27458 (I469315,I2507,I469247,I469341,);
DFFARX1 I_27459 (I469341,I2507,I469247,I469236,);
DFFARX1 I_27460 (I690051,I2507,I469247,I469372,);
nand I_27461 (I469380,I469372,I690066);
not I_27462 (I469397,I469380);
DFFARX1 I_27463 (I469397,I2507,I469247,I469423,);
not I_27464 (I469431,I469423);
nor I_27465 (I469239,I469281,I469431);
DFFARX1 I_27466 (I690072,I2507,I469247,I469471,);
nor I_27467 (I469230,I469471,I469341);
nor I_27468 (I469221,I469471,I469397);
nand I_27469 (I469507,I690054,I690075);
and I_27470 (I469524,I469507,I690057);
DFFARX1 I_27471 (I469524,I2507,I469247,I469550,);
not I_27472 (I469558,I469550);
nand I_27473 (I469575,I469558,I469471);
nand I_27474 (I469224,I469558,I469380);
nor I_27475 (I469606,I690048,I690075);
and I_27476 (I469623,I469471,I469606);
nor I_27477 (I469640,I469558,I469623);
DFFARX1 I_27478 (I469640,I2507,I469247,I469233,);
nor I_27479 (I469671,I469273,I469606);
DFFARX1 I_27480 (I469671,I2507,I469247,I469218,);
nor I_27481 (I469702,I469550,I469606);
not I_27482 (I469719,I469702);
nand I_27483 (I469227,I469719,I469575);
not I_27484 (I469774,I2514);
DFFARX1 I_27485 (I86623,I2507,I469774,I469800,);
not I_27486 (I469808,I469800);
nand I_27487 (I469825,I86599,I86617);
and I_27488 (I469842,I469825,I86605);
DFFARX1 I_27489 (I469842,I2507,I469774,I469868,);
DFFARX1 I_27490 (I469868,I2507,I469774,I469763,);
DFFARX1 I_27491 (I86614,I2507,I469774,I469899,);
nand I_27492 (I469907,I469899,I86620);
not I_27493 (I469924,I469907);
DFFARX1 I_27494 (I469924,I2507,I469774,I469950,);
not I_27495 (I469958,I469950);
nor I_27496 (I469766,I469808,I469958);
DFFARX1 I_27497 (I86599,I2507,I469774,I469998,);
nor I_27498 (I469757,I469998,I469868);
nor I_27499 (I469748,I469998,I469924);
nand I_27500 (I470034,I86611,I86602);
and I_27501 (I470051,I470034,I86626);
DFFARX1 I_27502 (I470051,I2507,I469774,I470077,);
not I_27503 (I470085,I470077);
nand I_27504 (I470102,I470085,I469998);
nand I_27505 (I469751,I470085,I469907);
nor I_27506 (I470133,I86608,I86602);
and I_27507 (I470150,I469998,I470133);
nor I_27508 (I470167,I470085,I470150);
DFFARX1 I_27509 (I470167,I2507,I469774,I469760,);
nor I_27510 (I470198,I469800,I470133);
DFFARX1 I_27511 (I470198,I2507,I469774,I469745,);
nor I_27512 (I470229,I470077,I470133);
not I_27513 (I470246,I470229);
nand I_27514 (I469754,I470246,I470102);
not I_27515 (I470301,I2514);
DFFARX1 I_27516 (I9853,I2507,I470301,I470327,);
not I_27517 (I470335,I470327);
nand I_27518 (I470352,I9865,I9868);
and I_27519 (I470369,I470352,I9844);
DFFARX1 I_27520 (I470369,I2507,I470301,I470395,);
DFFARX1 I_27521 (I470395,I2507,I470301,I470290,);
DFFARX1 I_27522 (I9862,I2507,I470301,I470426,);
nand I_27523 (I470434,I470426,I9850);
not I_27524 (I470451,I470434);
DFFARX1 I_27525 (I470451,I2507,I470301,I470477,);
not I_27526 (I470485,I470477);
nor I_27527 (I470293,I470335,I470485);
DFFARX1 I_27528 (I9847,I2507,I470301,I470525,);
nor I_27529 (I470284,I470525,I470395);
nor I_27530 (I470275,I470525,I470451);
nand I_27531 (I470561,I9856,I9847);
and I_27532 (I470578,I470561,I9844);
DFFARX1 I_27533 (I470578,I2507,I470301,I470604,);
not I_27534 (I470612,I470604);
nand I_27535 (I470629,I470612,I470525);
nand I_27536 (I470278,I470612,I470434);
nor I_27537 (I470660,I9859,I9847);
and I_27538 (I470677,I470525,I470660);
nor I_27539 (I470694,I470612,I470677);
DFFARX1 I_27540 (I470694,I2507,I470301,I470287,);
nor I_27541 (I470725,I470327,I470660);
DFFARX1 I_27542 (I470725,I2507,I470301,I470272,);
nor I_27543 (I470756,I470604,I470660);
not I_27544 (I470773,I470756);
nand I_27545 (I470281,I470773,I470629);
not I_27546 (I470828,I2514);
DFFARX1 I_27547 (I669989,I2507,I470828,I470854,);
not I_27548 (I470862,I470854);
nand I_27549 (I470879,I669971,I669974);
and I_27550 (I470896,I470879,I669986);
DFFARX1 I_27551 (I470896,I2507,I470828,I470922,);
DFFARX1 I_27552 (I470922,I2507,I470828,I470817,);
DFFARX1 I_27553 (I669995,I2507,I470828,I470953,);
nand I_27554 (I470961,I470953,I669980);
not I_27555 (I470978,I470961);
DFFARX1 I_27556 (I470978,I2507,I470828,I471004,);
not I_27557 (I471012,I471004);
nor I_27558 (I470820,I470862,I471012);
DFFARX1 I_27559 (I669992,I2507,I470828,I471052,);
nor I_27560 (I470811,I471052,I470922);
nor I_27561 (I470802,I471052,I470978);
nand I_27562 (I471088,I669983,I669977);
and I_27563 (I471105,I471088,I669971);
DFFARX1 I_27564 (I471105,I2507,I470828,I471131,);
not I_27565 (I471139,I471131);
nand I_27566 (I471156,I471139,I471052);
nand I_27567 (I470805,I471139,I470961);
nor I_27568 (I471187,I669974,I669977);
and I_27569 (I471204,I471052,I471187);
nor I_27570 (I471221,I471139,I471204);
DFFARX1 I_27571 (I471221,I2507,I470828,I470814,);
nor I_27572 (I471252,I470854,I471187);
DFFARX1 I_27573 (I471252,I2507,I470828,I470799,);
nor I_27574 (I471283,I471131,I471187);
not I_27575 (I471300,I471283);
nand I_27576 (I470808,I471300,I471156);
not I_27577 (I471355,I2514);
DFFARX1 I_27578 (I635275,I2507,I471355,I471381,);
not I_27579 (I471389,I471381);
nand I_27580 (I471406,I635257,I635257);
and I_27581 (I471423,I471406,I635263);
DFFARX1 I_27582 (I471423,I2507,I471355,I471449,);
DFFARX1 I_27583 (I471449,I2507,I471355,I471344,);
DFFARX1 I_27584 (I635260,I2507,I471355,I471480,);
nand I_27585 (I471488,I471480,I635269);
not I_27586 (I471505,I471488);
DFFARX1 I_27587 (I471505,I2507,I471355,I471531,);
not I_27588 (I471539,I471531);
nor I_27589 (I471347,I471389,I471539);
DFFARX1 I_27590 (I635281,I2507,I471355,I471579,);
nor I_27591 (I471338,I471579,I471449);
nor I_27592 (I471329,I471579,I471505);
nand I_27593 (I471615,I635272,I635266);
and I_27594 (I471632,I471615,I635260);
DFFARX1 I_27595 (I471632,I2507,I471355,I471658,);
not I_27596 (I471666,I471658);
nand I_27597 (I471683,I471666,I471579);
nand I_27598 (I471332,I471666,I471488);
nor I_27599 (I471714,I635278,I635266);
and I_27600 (I471731,I471579,I471714);
nor I_27601 (I471748,I471666,I471731);
DFFARX1 I_27602 (I471748,I2507,I471355,I471341,);
nor I_27603 (I471779,I471381,I471714);
DFFARX1 I_27604 (I471779,I2507,I471355,I471326,);
nor I_27605 (I471810,I471658,I471714);
not I_27606 (I471827,I471810);
nand I_27607 (I471335,I471827,I471683);
not I_27608 (I471882,I2514);
DFFARX1 I_27609 (I426429,I2507,I471882,I471908,);
not I_27610 (I471916,I471908);
nand I_27611 (I471933,I426432,I426429);
and I_27612 (I471950,I471933,I426441);
DFFARX1 I_27613 (I471950,I2507,I471882,I471976,);
DFFARX1 I_27614 (I471976,I2507,I471882,I471871,);
DFFARX1 I_27615 (I426438,I2507,I471882,I472007,);
nand I_27616 (I472015,I472007,I426444);
not I_27617 (I472032,I472015);
DFFARX1 I_27618 (I472032,I2507,I471882,I472058,);
not I_27619 (I472066,I472058);
nor I_27620 (I471874,I471916,I472066);
DFFARX1 I_27621 (I426453,I2507,I471882,I472106,);
nor I_27622 (I471865,I472106,I471976);
nor I_27623 (I471856,I472106,I472032);
nand I_27624 (I472142,I426447,I426435);
and I_27625 (I472159,I472142,I426432);
DFFARX1 I_27626 (I472159,I2507,I471882,I472185,);
not I_27627 (I472193,I472185);
nand I_27628 (I472210,I472193,I472106);
nand I_27629 (I471859,I472193,I472015);
nor I_27630 (I472241,I426450,I426435);
and I_27631 (I472258,I472106,I472241);
nor I_27632 (I472275,I472193,I472258);
DFFARX1 I_27633 (I472275,I2507,I471882,I471868,);
nor I_27634 (I472306,I471908,I472241);
DFFARX1 I_27635 (I472306,I2507,I471882,I471853,);
nor I_27636 (I472337,I472185,I472241);
not I_27637 (I472354,I472337);
nand I_27638 (I471862,I472354,I472210);
not I_27639 (I472409,I2514);
DFFARX1 I_27640 (I189050,I2507,I472409,I472435,);
not I_27641 (I472443,I472435);
nand I_27642 (I472460,I189041,I189041);
and I_27643 (I472477,I472460,I189059);
DFFARX1 I_27644 (I472477,I2507,I472409,I472503,);
DFFARX1 I_27645 (I472503,I2507,I472409,I472398,);
DFFARX1 I_27646 (I189062,I2507,I472409,I472534,);
nand I_27647 (I472542,I472534,I189044);
not I_27648 (I472559,I472542);
DFFARX1 I_27649 (I472559,I2507,I472409,I472585,);
not I_27650 (I472593,I472585);
nor I_27651 (I472401,I472443,I472593);
DFFARX1 I_27652 (I189056,I2507,I472409,I472633,);
nor I_27653 (I472392,I472633,I472503);
nor I_27654 (I472383,I472633,I472559);
nand I_27655 (I472669,I189068,I189047);
and I_27656 (I472686,I472669,I189053);
DFFARX1 I_27657 (I472686,I2507,I472409,I472712,);
not I_27658 (I472720,I472712);
nand I_27659 (I472737,I472720,I472633);
nand I_27660 (I472386,I472720,I472542);
nor I_27661 (I472768,I189065,I189047);
and I_27662 (I472785,I472633,I472768);
nor I_27663 (I472802,I472720,I472785);
DFFARX1 I_27664 (I472802,I2507,I472409,I472395,);
nor I_27665 (I472833,I472435,I472768);
DFFARX1 I_27666 (I472833,I2507,I472409,I472380,);
nor I_27667 (I472864,I472712,I472768);
not I_27668 (I472881,I472864);
nand I_27669 (I472389,I472881,I472737);
not I_27670 (I472936,I2514);
DFFARX1 I_27671 (I394639,I2507,I472936,I472962,);
not I_27672 (I472970,I472962);
nand I_27673 (I472987,I394642,I394639);
and I_27674 (I473004,I472987,I394651);
DFFARX1 I_27675 (I473004,I2507,I472936,I473030,);
DFFARX1 I_27676 (I473030,I2507,I472936,I472925,);
DFFARX1 I_27677 (I394648,I2507,I472936,I473061,);
nand I_27678 (I473069,I473061,I394654);
not I_27679 (I473086,I473069);
DFFARX1 I_27680 (I473086,I2507,I472936,I473112,);
not I_27681 (I473120,I473112);
nor I_27682 (I472928,I472970,I473120);
DFFARX1 I_27683 (I394663,I2507,I472936,I473160,);
nor I_27684 (I472919,I473160,I473030);
nor I_27685 (I472910,I473160,I473086);
nand I_27686 (I473196,I394657,I394645);
and I_27687 (I473213,I473196,I394642);
DFFARX1 I_27688 (I473213,I2507,I472936,I473239,);
not I_27689 (I473247,I473239);
nand I_27690 (I473264,I473247,I473160);
nand I_27691 (I472913,I473247,I473069);
nor I_27692 (I473295,I394660,I394645);
and I_27693 (I473312,I473160,I473295);
nor I_27694 (I473329,I473247,I473312);
DFFARX1 I_27695 (I473329,I2507,I472936,I472922,);
nor I_27696 (I473360,I472962,I473295);
DFFARX1 I_27697 (I473360,I2507,I472936,I472907,);
nor I_27698 (I473391,I473239,I473295);
not I_27699 (I473408,I473391);
nand I_27700 (I472916,I473408,I473264);
not I_27701 (I473463,I2514);
DFFARX1 I_27702 (I477653,I2507,I473463,I473489,);
not I_27703 (I473497,I473489);
nand I_27704 (I473514,I477668,I477650);
and I_27705 (I473531,I473514,I477650);
DFFARX1 I_27706 (I473531,I2507,I473463,I473557,);
DFFARX1 I_27707 (I473557,I2507,I473463,I473452,);
DFFARX1 I_27708 (I477659,I2507,I473463,I473588,);
nand I_27709 (I473596,I473588,I477677);
not I_27710 (I473613,I473596);
DFFARX1 I_27711 (I473613,I2507,I473463,I473639,);
not I_27712 (I473647,I473639);
nor I_27713 (I473455,I473497,I473647);
DFFARX1 I_27714 (I477674,I2507,I473463,I473687,);
nor I_27715 (I473446,I473687,I473557);
nor I_27716 (I473437,I473687,I473613);
nand I_27717 (I473723,I477671,I477662);
and I_27718 (I473740,I473723,I477656);
DFFARX1 I_27719 (I473740,I2507,I473463,I473766,);
not I_27720 (I473774,I473766);
nand I_27721 (I473791,I473774,I473687);
nand I_27722 (I473440,I473774,I473596);
nor I_27723 (I473822,I477665,I477662);
and I_27724 (I473839,I473687,I473822);
nor I_27725 (I473856,I473774,I473839);
DFFARX1 I_27726 (I473856,I2507,I473463,I473449,);
nor I_27727 (I473887,I473489,I473822);
DFFARX1 I_27728 (I473887,I2507,I473463,I473434,);
nor I_27729 (I473918,I473766,I473822);
not I_27730 (I473935,I473918);
nand I_27731 (I473443,I473935,I473791);
not I_27732 (I473990,I2514);
DFFARX1 I_27733 (I229694,I2507,I473990,I474016,);
not I_27734 (I474024,I474016);
nand I_27735 (I474041,I229691,I229700);
and I_27736 (I474058,I474041,I229709);
DFFARX1 I_27737 (I474058,I2507,I473990,I474084,);
DFFARX1 I_27738 (I474084,I2507,I473990,I473979,);
DFFARX1 I_27739 (I229712,I2507,I473990,I474115,);
nand I_27740 (I474123,I474115,I229715);
not I_27741 (I474140,I474123);
DFFARX1 I_27742 (I474140,I2507,I473990,I474166,);
not I_27743 (I474174,I474166);
nor I_27744 (I473982,I474024,I474174);
DFFARX1 I_27745 (I229688,I2507,I473990,I474214,);
nor I_27746 (I473973,I474214,I474084);
nor I_27747 (I473964,I474214,I474140);
nand I_27748 (I474250,I229703,I229706);
and I_27749 (I474267,I474250,I229697);
DFFARX1 I_27750 (I474267,I2507,I473990,I474293,);
not I_27751 (I474301,I474293);
nand I_27752 (I474318,I474301,I474214);
nand I_27753 (I473967,I474301,I474123);
nor I_27754 (I474349,I229688,I229706);
and I_27755 (I474366,I474214,I474349);
nor I_27756 (I474383,I474301,I474366);
DFFARX1 I_27757 (I474383,I2507,I473990,I473976,);
nor I_27758 (I474414,I474016,I474349);
DFFARX1 I_27759 (I474414,I2507,I473990,I473961,);
nor I_27760 (I474445,I474293,I474349);
not I_27761 (I474462,I474445);
nand I_27762 (I473970,I474462,I474318);
not I_27763 (I474517,I2514);
DFFARX1 I_27764 (I356491,I2507,I474517,I474543,);
not I_27765 (I474551,I474543);
nand I_27766 (I474568,I356494,I356491);
and I_27767 (I474585,I474568,I356503);
DFFARX1 I_27768 (I474585,I2507,I474517,I474611,);
DFFARX1 I_27769 (I474611,I2507,I474517,I474506,);
DFFARX1 I_27770 (I356500,I2507,I474517,I474642,);
nand I_27771 (I474650,I474642,I356506);
not I_27772 (I474667,I474650);
DFFARX1 I_27773 (I474667,I2507,I474517,I474693,);
not I_27774 (I474701,I474693);
nor I_27775 (I474509,I474551,I474701);
DFFARX1 I_27776 (I356515,I2507,I474517,I474741,);
nor I_27777 (I474500,I474741,I474611);
nor I_27778 (I474491,I474741,I474667);
nand I_27779 (I474777,I356509,I356497);
and I_27780 (I474794,I474777,I356494);
DFFARX1 I_27781 (I474794,I2507,I474517,I474820,);
not I_27782 (I474828,I474820);
nand I_27783 (I474845,I474828,I474741);
nand I_27784 (I474494,I474828,I474650);
nor I_27785 (I474876,I356512,I356497);
and I_27786 (I474893,I474741,I474876);
nor I_27787 (I474910,I474828,I474893);
DFFARX1 I_27788 (I474910,I2507,I474517,I474503,);
nor I_27789 (I474941,I474543,I474876);
DFFARX1 I_27790 (I474941,I2507,I474517,I474488,);
nor I_27791 (I474972,I474820,I474876);
not I_27792 (I474989,I474972);
nand I_27793 (I474497,I474989,I474845);
not I_27794 (I475044,I2514);
DFFARX1 I_27795 (I624871,I2507,I475044,I475070,);
not I_27796 (I475078,I475070);
nand I_27797 (I475095,I624853,I624853);
and I_27798 (I475112,I475095,I624859);
DFFARX1 I_27799 (I475112,I2507,I475044,I475138,);
DFFARX1 I_27800 (I475138,I2507,I475044,I475033,);
DFFARX1 I_27801 (I624856,I2507,I475044,I475169,);
nand I_27802 (I475177,I475169,I624865);
not I_27803 (I475194,I475177);
DFFARX1 I_27804 (I475194,I2507,I475044,I475220,);
not I_27805 (I475228,I475220);
nor I_27806 (I475036,I475078,I475228);
DFFARX1 I_27807 (I624877,I2507,I475044,I475268,);
nor I_27808 (I475027,I475268,I475138);
nor I_27809 (I475018,I475268,I475194);
nand I_27810 (I475304,I624868,I624862);
and I_27811 (I475321,I475304,I624856);
DFFARX1 I_27812 (I475321,I2507,I475044,I475347,);
not I_27813 (I475355,I475347);
nand I_27814 (I475372,I475355,I475268);
nand I_27815 (I475021,I475355,I475177);
nor I_27816 (I475403,I624874,I624862);
and I_27817 (I475420,I475268,I475403);
nor I_27818 (I475437,I475355,I475420);
DFFARX1 I_27819 (I475437,I2507,I475044,I475030,);
nor I_27820 (I475468,I475070,I475403);
DFFARX1 I_27821 (I475468,I2507,I475044,I475015,);
nor I_27822 (I475499,I475347,I475403);
not I_27823 (I475516,I475499);
nand I_27824 (I475024,I475516,I475372);
not I_27825 (I475571,I2514);
DFFARX1 I_27826 (I144320,I2507,I475571,I475597,);
not I_27827 (I475605,I475597);
nand I_27828 (I475622,I144317,I144335);
and I_27829 (I475639,I475622,I144326);
DFFARX1 I_27830 (I475639,I2507,I475571,I475665,);
DFFARX1 I_27831 (I475665,I2507,I475571,I475560,);
DFFARX1 I_27832 (I144332,I2507,I475571,I475696,);
nand I_27833 (I475704,I475696,I144329);
not I_27834 (I475721,I475704);
DFFARX1 I_27835 (I475721,I2507,I475571,I475747,);
not I_27836 (I475755,I475747);
nor I_27837 (I475563,I475605,I475755);
DFFARX1 I_27838 (I144323,I2507,I475571,I475795,);
nor I_27839 (I475554,I475795,I475665);
nor I_27840 (I475545,I475795,I475721);
nand I_27841 (I475831,I144314,I144338);
and I_27842 (I475848,I475831,I144317);
DFFARX1 I_27843 (I475848,I2507,I475571,I475874,);
not I_27844 (I475882,I475874);
nand I_27845 (I475899,I475882,I475795);
nand I_27846 (I475548,I475882,I475704);
nor I_27847 (I475930,I144314,I144338);
and I_27848 (I475947,I475795,I475930);
nor I_27849 (I475964,I475882,I475947);
DFFARX1 I_27850 (I475964,I2507,I475571,I475557,);
nor I_27851 (I475995,I475597,I475930);
DFFARX1 I_27852 (I475995,I2507,I475571,I475542,);
nor I_27853 (I476026,I475874,I475930);
not I_27854 (I476043,I476026);
nand I_27855 (I475551,I476043,I475899);
not I_27856 (I476098,I2514);
DFFARX1 I_27857 (I176929,I2507,I476098,I476124,);
not I_27858 (I476132,I476124);
nand I_27859 (I476149,I176920,I176920);
and I_27860 (I476166,I476149,I176938);
DFFARX1 I_27861 (I476166,I2507,I476098,I476192,);
DFFARX1 I_27862 (I476192,I2507,I476098,I476087,);
DFFARX1 I_27863 (I176941,I2507,I476098,I476223,);
nand I_27864 (I476231,I476223,I176923);
not I_27865 (I476248,I476231);
DFFARX1 I_27866 (I476248,I2507,I476098,I476274,);
not I_27867 (I476282,I476274);
nor I_27868 (I476090,I476132,I476282);
DFFARX1 I_27869 (I176935,I2507,I476098,I476322,);
nor I_27870 (I476081,I476322,I476192);
nor I_27871 (I476072,I476322,I476248);
nand I_27872 (I476358,I176947,I176926);
and I_27873 (I476375,I476358,I176932);
DFFARX1 I_27874 (I476375,I2507,I476098,I476401,);
not I_27875 (I476409,I476401);
nand I_27876 (I476426,I476409,I476322);
nand I_27877 (I476075,I476409,I476231);
nor I_27878 (I476457,I176944,I176926);
and I_27879 (I476474,I476322,I476457);
nor I_27880 (I476491,I476409,I476474);
DFFARX1 I_27881 (I476491,I2507,I476098,I476084,);
nor I_27882 (I476522,I476124,I476457);
DFFARX1 I_27883 (I476522,I2507,I476098,I476069,);
nor I_27884 (I476553,I476401,I476457);
not I_27885 (I476570,I476553);
nand I_27886 (I476078,I476570,I476426);
not I_27887 (I476625,I2514);
DFFARX1 I_27888 (I215400,I2507,I476625,I476651,);
not I_27889 (I476659,I476651);
nand I_27890 (I476676,I215391,I215391);
and I_27891 (I476693,I476676,I215409);
DFFARX1 I_27892 (I476693,I2507,I476625,I476719,);
DFFARX1 I_27893 (I476719,I2507,I476625,I476614,);
DFFARX1 I_27894 (I215412,I2507,I476625,I476750,);
nand I_27895 (I476758,I476750,I215394);
not I_27896 (I476775,I476758);
DFFARX1 I_27897 (I476775,I2507,I476625,I476801,);
not I_27898 (I476809,I476801);
nor I_27899 (I476617,I476659,I476809);
DFFARX1 I_27900 (I215406,I2507,I476625,I476849,);
nor I_27901 (I476608,I476849,I476719);
nor I_27902 (I476599,I476849,I476775);
nand I_27903 (I476885,I215418,I215397);
and I_27904 (I476902,I476885,I215403);
DFFARX1 I_27905 (I476902,I2507,I476625,I476928,);
not I_27906 (I476936,I476928);
nand I_27907 (I476953,I476936,I476849);
nand I_27908 (I476602,I476936,I476758);
nor I_27909 (I476984,I215415,I215397);
and I_27910 (I477001,I476849,I476984);
nor I_27911 (I477018,I476936,I477001);
DFFARX1 I_27912 (I477018,I2507,I476625,I476611,);
nor I_27913 (I477049,I476651,I476984);
DFFARX1 I_27914 (I477049,I2507,I476625,I476596,);
nor I_27915 (I477080,I476928,I476984);
not I_27916 (I477097,I477080);
nand I_27917 (I476605,I477097,I476953);
not I_27918 (I477152,I2514);
DFFARX1 I_27919 (I165862,I2507,I477152,I477178,);
not I_27920 (I477186,I477178);
nand I_27921 (I477203,I165853,I165853);
and I_27922 (I477220,I477203,I165871);
DFFARX1 I_27923 (I477220,I2507,I477152,I477246,);
DFFARX1 I_27924 (I477246,I2507,I477152,I477141,);
DFFARX1 I_27925 (I165874,I2507,I477152,I477277,);
nand I_27926 (I477285,I477277,I165856);
not I_27927 (I477302,I477285);
DFFARX1 I_27928 (I477302,I2507,I477152,I477328,);
not I_27929 (I477336,I477328);
nor I_27930 (I477144,I477186,I477336);
DFFARX1 I_27931 (I165868,I2507,I477152,I477376,);
nor I_27932 (I477135,I477376,I477246);
nor I_27933 (I477126,I477376,I477302);
nand I_27934 (I477412,I165880,I165859);
and I_27935 (I477429,I477412,I165865);
DFFARX1 I_27936 (I477429,I2507,I477152,I477455,);
not I_27937 (I477463,I477455);
nand I_27938 (I477480,I477463,I477376);
nand I_27939 (I477129,I477463,I477285);
nor I_27940 (I477511,I165877,I165859);
and I_27941 (I477528,I477376,I477511);
nor I_27942 (I477545,I477463,I477528);
DFFARX1 I_27943 (I477545,I2507,I477152,I477138,);
nor I_27944 (I477576,I477178,I477511);
DFFARX1 I_27945 (I477576,I2507,I477152,I477123,);
nor I_27946 (I477607,I477455,I477511);
not I_27947 (I477624,I477607);
nand I_27948 (I477132,I477624,I477480);
not I_27949 (I477685,I2514);
DFFARX1 I_27950 (I584411,I2507,I477685,I477711,);
DFFARX1 I_27951 (I584393,I2507,I477685,I477728,);
not I_27952 (I477736,I477728);
not I_27953 (I477753,I584402);
nor I_27954 (I477770,I477753,I584414);
not I_27955 (I477787,I584396);
nor I_27956 (I477804,I477770,I584405);
nor I_27957 (I477821,I477728,I477804);
DFFARX1 I_27958 (I477821,I2507,I477685,I477671,);
nor I_27959 (I477852,I584405,I584414);
nand I_27960 (I477869,I477852,I584402);
DFFARX1 I_27961 (I477869,I2507,I477685,I477674,);
nor I_27962 (I477900,I477787,I584405);
nand I_27963 (I477917,I477900,I584417);
nor I_27964 (I477934,I477711,I477917);
DFFARX1 I_27965 (I477934,I2507,I477685,I477650,);
not I_27966 (I477965,I477917);
nand I_27967 (I477662,I477728,I477965);
DFFARX1 I_27968 (I477917,I2507,I477685,I478005,);
not I_27969 (I478013,I478005);
not I_27970 (I478030,I584405);
not I_27971 (I478047,I584393);
nor I_27972 (I478064,I478047,I584396);
nor I_27973 (I477677,I478013,I478064);
nor I_27974 (I478095,I478047,I584399);
and I_27975 (I478112,I478095,I584408);
or I_27976 (I478129,I478112,I584396);
DFFARX1 I_27977 (I478129,I2507,I477685,I478155,);
nor I_27978 (I477665,I478155,I477711);
not I_27979 (I478177,I478155);
and I_27980 (I478194,I478177,I477711);
nor I_27981 (I477659,I477736,I478194);
nand I_27982 (I478225,I478177,I477787);
nor I_27983 (I477653,I478047,I478225);
nand I_27984 (I477656,I478177,I477965);
nand I_27985 (I478270,I477787,I584393);
nor I_27986 (I477668,I478030,I478270);
not I_27987 (I478331,I2514);
DFFARX1 I_27988 (I272126,I2507,I478331,I478357,);
DFFARX1 I_27989 (I272123,I2507,I478331,I478374,);
not I_27990 (I478382,I478374);
not I_27991 (I478399,I272138);
nor I_27992 (I478416,I478399,I272141);
not I_27993 (I478433,I272129);
nor I_27994 (I478450,I478416,I272135);
nor I_27995 (I478467,I478374,I478450);
DFFARX1 I_27996 (I478467,I2507,I478331,I478317,);
nor I_27997 (I478498,I272135,I272141);
nand I_27998 (I478515,I478498,I272138);
DFFARX1 I_27999 (I478515,I2507,I478331,I478320,);
nor I_28000 (I478546,I478433,I272135);
nand I_28001 (I478563,I478546,I272147);
nor I_28002 (I478580,I478357,I478563);
DFFARX1 I_28003 (I478580,I2507,I478331,I478296,);
not I_28004 (I478611,I478563);
nand I_28005 (I478308,I478374,I478611);
DFFARX1 I_28006 (I478563,I2507,I478331,I478651,);
not I_28007 (I478659,I478651);
not I_28008 (I478676,I272135);
not I_28009 (I478693,I272120);
nor I_28010 (I478710,I478693,I272129);
nor I_28011 (I478323,I478659,I478710);
nor I_28012 (I478741,I478693,I272132);
and I_28013 (I478758,I478741,I272120);
or I_28014 (I478775,I478758,I272144);
DFFARX1 I_28015 (I478775,I2507,I478331,I478801,);
nor I_28016 (I478311,I478801,I478357);
not I_28017 (I478823,I478801);
and I_28018 (I478840,I478823,I478357);
nor I_28019 (I478305,I478382,I478840);
nand I_28020 (I478871,I478823,I478433);
nor I_28021 (I478299,I478693,I478871);
nand I_28022 (I478302,I478823,I478611);
nand I_28023 (I478916,I478433,I272120);
nor I_28024 (I478314,I478676,I478916);
not I_28025 (I478977,I2514);
DFFARX1 I_28026 (I406205,I2507,I478977,I479003,);
DFFARX1 I_28027 (I406199,I2507,I478977,I479020,);
not I_28028 (I479028,I479020);
not I_28029 (I479045,I406214);
nor I_28030 (I479062,I479045,I406199);
not I_28031 (I479079,I406208);
nor I_28032 (I479096,I479062,I406217);
nor I_28033 (I479113,I479020,I479096);
DFFARX1 I_28034 (I479113,I2507,I478977,I478963,);
nor I_28035 (I479144,I406217,I406199);
nand I_28036 (I479161,I479144,I406214);
DFFARX1 I_28037 (I479161,I2507,I478977,I478966,);
nor I_28038 (I479192,I479079,I406217);
nand I_28039 (I479209,I479192,I406202);
nor I_28040 (I479226,I479003,I479209);
DFFARX1 I_28041 (I479226,I2507,I478977,I478942,);
not I_28042 (I479257,I479209);
nand I_28043 (I478954,I479020,I479257);
DFFARX1 I_28044 (I479209,I2507,I478977,I479297,);
not I_28045 (I479305,I479297);
not I_28046 (I479322,I406217);
not I_28047 (I479339,I406211);
nor I_28048 (I479356,I479339,I406208);
nor I_28049 (I478969,I479305,I479356);
nor I_28050 (I479387,I479339,I406220);
and I_28051 (I479404,I479387,I406223);
or I_28052 (I479421,I479404,I406202);
DFFARX1 I_28053 (I479421,I2507,I478977,I479447,);
nor I_28054 (I478957,I479447,I479003);
not I_28055 (I479469,I479447);
and I_28056 (I479486,I479469,I479003);
nor I_28057 (I478951,I479028,I479486);
nand I_28058 (I479517,I479469,I479079);
nor I_28059 (I478945,I479339,I479517);
nand I_28060 (I478948,I479469,I479257);
nand I_28061 (I479562,I479079,I406211);
nor I_28062 (I478960,I479322,I479562);
not I_28063 (I479623,I2514);
DFFARX1 I_28064 (I192203,I2507,I479623,I479649,);
DFFARX1 I_28065 (I192209,I2507,I479623,I479666,);
not I_28066 (I479674,I479666);
not I_28067 (I479691,I192230);
nor I_28068 (I479708,I479691,I192218);
not I_28069 (I479725,I192227);
nor I_28070 (I479742,I479708,I192212);
nor I_28071 (I479759,I479666,I479742);
DFFARX1 I_28072 (I479759,I2507,I479623,I479609,);
nor I_28073 (I479790,I192212,I192218);
nand I_28074 (I479807,I479790,I192230);
DFFARX1 I_28075 (I479807,I2507,I479623,I479612,);
nor I_28076 (I479838,I479725,I192212);
nand I_28077 (I479855,I479838,I192203);
nor I_28078 (I479872,I479649,I479855);
DFFARX1 I_28079 (I479872,I2507,I479623,I479588,);
not I_28080 (I479903,I479855);
nand I_28081 (I479600,I479666,I479903);
DFFARX1 I_28082 (I479855,I2507,I479623,I479943,);
not I_28083 (I479951,I479943);
not I_28084 (I479968,I192212);
not I_28085 (I479985,I192215);
nor I_28086 (I480002,I479985,I192227);
nor I_28087 (I479615,I479951,I480002);
nor I_28088 (I480033,I479985,I192224);
and I_28089 (I480050,I480033,I192206);
or I_28090 (I480067,I480050,I192221);
DFFARX1 I_28091 (I480067,I2507,I479623,I480093,);
nor I_28092 (I479603,I480093,I479649);
not I_28093 (I480115,I480093);
and I_28094 (I480132,I480115,I479649);
nor I_28095 (I479597,I479674,I480132);
nand I_28096 (I480163,I480115,I479725);
nor I_28097 (I479591,I479985,I480163);
nand I_28098 (I479594,I480115,I479903);
nand I_28099 (I480208,I479725,I192215);
nor I_28100 (I479606,I479968,I480208);
not I_28101 (I480269,I2514);
DFFARX1 I_28102 (I167961,I2507,I480269,I480295,);
DFFARX1 I_28103 (I167967,I2507,I480269,I480312,);
not I_28104 (I480320,I480312);
not I_28105 (I480337,I167988);
nor I_28106 (I480354,I480337,I167976);
not I_28107 (I480371,I167985);
nor I_28108 (I480388,I480354,I167970);
nor I_28109 (I480405,I480312,I480388);
DFFARX1 I_28110 (I480405,I2507,I480269,I480255,);
nor I_28111 (I480436,I167970,I167976);
nand I_28112 (I480453,I480436,I167988);
DFFARX1 I_28113 (I480453,I2507,I480269,I480258,);
nor I_28114 (I480484,I480371,I167970);
nand I_28115 (I480501,I480484,I167961);
nor I_28116 (I480518,I480295,I480501);
DFFARX1 I_28117 (I480518,I2507,I480269,I480234,);
not I_28118 (I480549,I480501);
nand I_28119 (I480246,I480312,I480549);
DFFARX1 I_28120 (I480501,I2507,I480269,I480589,);
not I_28121 (I480597,I480589);
not I_28122 (I480614,I167970);
not I_28123 (I480631,I167973);
nor I_28124 (I480648,I480631,I167985);
nor I_28125 (I480261,I480597,I480648);
nor I_28126 (I480679,I480631,I167982);
and I_28127 (I480696,I480679,I167964);
or I_28128 (I480713,I480696,I167979);
DFFARX1 I_28129 (I480713,I2507,I480269,I480739,);
nor I_28130 (I480249,I480739,I480295);
not I_28131 (I480761,I480739);
and I_28132 (I480778,I480761,I480295);
nor I_28133 (I480243,I480320,I480778);
nand I_28134 (I480809,I480761,I480371);
nor I_28135 (I480237,I480631,I480809);
nand I_28136 (I480240,I480761,I480549);
nand I_28137 (I480854,I480371,I167973);
nor I_28138 (I480252,I480614,I480854);
not I_28139 (I480915,I2514);
DFFARX1 I_28140 (I140750,I2507,I480915,I480941,);
DFFARX1 I_28141 (I140762,I2507,I480915,I480958,);
not I_28142 (I480966,I480958);
not I_28143 (I480983,I140768);
nor I_28144 (I481000,I480983,I140753);
not I_28145 (I481017,I140744);
nor I_28146 (I481034,I481000,I140765);
nor I_28147 (I481051,I480958,I481034);
DFFARX1 I_28148 (I481051,I2507,I480915,I480901,);
nor I_28149 (I481082,I140765,I140753);
nand I_28150 (I481099,I481082,I140768);
DFFARX1 I_28151 (I481099,I2507,I480915,I480904,);
nor I_28152 (I481130,I481017,I140765);
nand I_28153 (I481147,I481130,I140747);
nor I_28154 (I481164,I480941,I481147);
DFFARX1 I_28155 (I481164,I2507,I480915,I480880,);
not I_28156 (I481195,I481147);
nand I_28157 (I480892,I480958,I481195);
DFFARX1 I_28158 (I481147,I2507,I480915,I481235,);
not I_28159 (I481243,I481235);
not I_28160 (I481260,I140765);
not I_28161 (I481277,I140756);
nor I_28162 (I481294,I481277,I140744);
nor I_28163 (I480907,I481243,I481294);
nor I_28164 (I481325,I481277,I140759);
and I_28165 (I481342,I481325,I140747);
or I_28166 (I481359,I481342,I140744);
DFFARX1 I_28167 (I481359,I2507,I480915,I481385,);
nor I_28168 (I480895,I481385,I480941);
not I_28169 (I481407,I481385);
and I_28170 (I481424,I481407,I480941);
nor I_28171 (I480889,I480966,I481424);
nand I_28172 (I481455,I481407,I481017);
nor I_28173 (I480883,I481277,I481455);
nand I_28174 (I480886,I481407,I481195);
nand I_28175 (I481500,I481017,I140756);
nor I_28176 (I480898,I481260,I481500);
not I_28177 (I481561,I2514);
DFFARX1 I_28178 (I629495,I2507,I481561,I481587,);
DFFARX1 I_28179 (I629477,I2507,I481561,I481604,);
not I_28180 (I481612,I481604);
not I_28181 (I481629,I629486);
nor I_28182 (I481646,I481629,I629498);
not I_28183 (I481663,I629480);
nor I_28184 (I481680,I481646,I629489);
nor I_28185 (I481697,I481604,I481680);
DFFARX1 I_28186 (I481697,I2507,I481561,I481547,);
nor I_28187 (I481728,I629489,I629498);
nand I_28188 (I481745,I481728,I629486);
DFFARX1 I_28189 (I481745,I2507,I481561,I481550,);
nor I_28190 (I481776,I481663,I629489);
nand I_28191 (I481793,I481776,I629501);
nor I_28192 (I481810,I481587,I481793);
DFFARX1 I_28193 (I481810,I2507,I481561,I481526,);
not I_28194 (I481841,I481793);
nand I_28195 (I481538,I481604,I481841);
DFFARX1 I_28196 (I481793,I2507,I481561,I481881,);
not I_28197 (I481889,I481881);
not I_28198 (I481906,I629489);
not I_28199 (I481923,I629477);
nor I_28200 (I481940,I481923,I629480);
nor I_28201 (I481553,I481889,I481940);
nor I_28202 (I481971,I481923,I629483);
and I_28203 (I481988,I481971,I629492);
or I_28204 (I482005,I481988,I629480);
DFFARX1 I_28205 (I482005,I2507,I481561,I482031,);
nor I_28206 (I481541,I482031,I481587);
not I_28207 (I482053,I482031);
and I_28208 (I482070,I482053,I481587);
nor I_28209 (I481535,I481612,I482070);
nand I_28210 (I482101,I482053,I481663);
nor I_28211 (I481529,I481923,I482101);
nand I_28212 (I481532,I482053,I481841);
nand I_28213 (I482146,I481663,I629477);
nor I_28214 (I481544,I481906,I482146);
not I_28215 (I482207,I2514);
DFFARX1 I_28216 (I153245,I2507,I482207,I482233,);
DFFARX1 I_28217 (I153257,I2507,I482207,I482250,);
not I_28218 (I482258,I482250);
not I_28219 (I482275,I153263);
nor I_28220 (I482292,I482275,I153248);
not I_28221 (I482309,I153239);
nor I_28222 (I482326,I482292,I153260);
nor I_28223 (I482343,I482250,I482326);
DFFARX1 I_28224 (I482343,I2507,I482207,I482193,);
nor I_28225 (I482374,I153260,I153248);
nand I_28226 (I482391,I482374,I153263);
DFFARX1 I_28227 (I482391,I2507,I482207,I482196,);
nor I_28228 (I482422,I482309,I153260);
nand I_28229 (I482439,I482422,I153242);
nor I_28230 (I482456,I482233,I482439);
DFFARX1 I_28231 (I482456,I2507,I482207,I482172,);
not I_28232 (I482487,I482439);
nand I_28233 (I482184,I482250,I482487);
DFFARX1 I_28234 (I482439,I2507,I482207,I482527,);
not I_28235 (I482535,I482527);
not I_28236 (I482552,I153260);
not I_28237 (I482569,I153251);
nor I_28238 (I482586,I482569,I153239);
nor I_28239 (I482199,I482535,I482586);
nor I_28240 (I482617,I482569,I153254);
and I_28241 (I482634,I482617,I153242);
or I_28242 (I482651,I482634,I153239);
DFFARX1 I_28243 (I482651,I2507,I482207,I482677,);
nor I_28244 (I482187,I482677,I482233);
not I_28245 (I482699,I482677);
and I_28246 (I482716,I482699,I482233);
nor I_28247 (I482181,I482258,I482716);
nand I_28248 (I482747,I482699,I482309);
nor I_28249 (I482175,I482569,I482747);
nand I_28250 (I482178,I482699,I482487);
nand I_28251 (I482792,I482309,I153251);
nor I_28252 (I482190,I482552,I482792);
not I_28253 (I482853,I2514);
DFFARX1 I_28254 (I452360,I2507,I482853,I482879,);
DFFARX1 I_28255 (I452357,I2507,I482853,I482896,);
not I_28256 (I482904,I482896);
not I_28257 (I482921,I452357);
nor I_28258 (I482938,I482921,I452360);
not I_28259 (I482955,I452372);
nor I_28260 (I482972,I482938,I452366);
nor I_28261 (I482989,I482896,I482972);
DFFARX1 I_28262 (I482989,I2507,I482853,I482839,);
nor I_28263 (I483020,I452366,I452360);
nand I_28264 (I483037,I483020,I452357);
DFFARX1 I_28265 (I483037,I2507,I482853,I482842,);
nor I_28266 (I483068,I482955,I452366);
nand I_28267 (I483085,I483068,I452354);
nor I_28268 (I483102,I482879,I483085);
DFFARX1 I_28269 (I483102,I2507,I482853,I482818,);
not I_28270 (I483133,I483085);
nand I_28271 (I482830,I482896,I483133);
DFFARX1 I_28272 (I483085,I2507,I482853,I483173,);
not I_28273 (I483181,I483173);
not I_28274 (I483198,I452366);
not I_28275 (I483215,I452363);
nor I_28276 (I483232,I483215,I452372);
nor I_28277 (I482845,I483181,I483232);
nor I_28278 (I483263,I483215,I452369);
and I_28279 (I483280,I483263,I452375);
or I_28280 (I483297,I483280,I452354);
DFFARX1 I_28281 (I483297,I2507,I482853,I483323,);
nor I_28282 (I482833,I483323,I482879);
not I_28283 (I483345,I483323);
and I_28284 (I483362,I483345,I482879);
nor I_28285 (I482827,I482904,I483362);
nand I_28286 (I483393,I483345,I482955);
nor I_28287 (I482821,I483215,I483393);
nand I_28288 (I482824,I483345,I483133);
nand I_28289 (I483438,I482955,I452363);
nor I_28290 (I482836,I483198,I483438);
not I_28291 (I483499,I2514);
DFFARX1 I_28292 (I654519,I2507,I483499,I483525,);
DFFARX1 I_28293 (I654525,I2507,I483499,I483542,);
not I_28294 (I483550,I483542);
not I_28295 (I483567,I654522);
nor I_28296 (I483584,I483567,I654501);
not I_28297 (I483601,I654504);
nor I_28298 (I483618,I483584,I654510);
nor I_28299 (I483635,I483542,I483618);
DFFARX1 I_28300 (I483635,I2507,I483499,I483485,);
nor I_28301 (I483666,I654510,I654501);
nand I_28302 (I483683,I483666,I654522);
DFFARX1 I_28303 (I483683,I2507,I483499,I483488,);
nor I_28304 (I483714,I483601,I654510);
nand I_28305 (I483731,I483714,I654504);
nor I_28306 (I483748,I483525,I483731);
DFFARX1 I_28307 (I483748,I2507,I483499,I483464,);
not I_28308 (I483779,I483731);
nand I_28309 (I483476,I483542,I483779);
DFFARX1 I_28310 (I483731,I2507,I483499,I483819,);
not I_28311 (I483827,I483819);
not I_28312 (I483844,I654510);
not I_28313 (I483861,I654513);
nor I_28314 (I483878,I483861,I654504);
nor I_28315 (I483491,I483827,I483878);
nor I_28316 (I483909,I483861,I654501);
and I_28317 (I483926,I483909,I654507);
or I_28318 (I483943,I483926,I654516);
DFFARX1 I_28319 (I483943,I2507,I483499,I483969,);
nor I_28320 (I483479,I483969,I483525);
not I_28321 (I483991,I483969);
and I_28322 (I484008,I483991,I483525);
nor I_28323 (I483473,I483550,I484008);
nand I_28324 (I484039,I483991,I483601);
nor I_28325 (I483467,I483861,I484039);
nand I_28326 (I483470,I483991,I483779);
nand I_28327 (I484084,I483601,I654513);
nor I_28328 (I483482,I483844,I484084);
not I_28329 (I484145,I2514);
DFFARX1 I_28330 (I177447,I2507,I484145,I484171,);
DFFARX1 I_28331 (I177453,I2507,I484145,I484188,);
not I_28332 (I484196,I484188);
not I_28333 (I484213,I177474);
nor I_28334 (I484230,I484213,I177462);
not I_28335 (I484247,I177471);
nor I_28336 (I484264,I484230,I177456);
nor I_28337 (I484281,I484188,I484264);
DFFARX1 I_28338 (I484281,I2507,I484145,I484131,);
nor I_28339 (I484312,I177456,I177462);
nand I_28340 (I484329,I484312,I177474);
DFFARX1 I_28341 (I484329,I2507,I484145,I484134,);
nor I_28342 (I484360,I484247,I177456);
nand I_28343 (I484377,I484360,I177447);
nor I_28344 (I484394,I484171,I484377);
DFFARX1 I_28345 (I484394,I2507,I484145,I484110,);
not I_28346 (I484425,I484377);
nand I_28347 (I484122,I484188,I484425);
DFFARX1 I_28348 (I484377,I2507,I484145,I484465,);
not I_28349 (I484473,I484465);
not I_28350 (I484490,I177456);
not I_28351 (I484507,I177459);
nor I_28352 (I484524,I484507,I177471);
nor I_28353 (I484137,I484473,I484524);
nor I_28354 (I484555,I484507,I177468);
and I_28355 (I484572,I484555,I177450);
or I_28356 (I484589,I484572,I177465);
DFFARX1 I_28357 (I484589,I2507,I484145,I484615,);
nor I_28358 (I484125,I484615,I484171);
not I_28359 (I484637,I484615);
and I_28360 (I484654,I484637,I484171);
nor I_28361 (I484119,I484196,I484654);
nand I_28362 (I484685,I484637,I484247);
nor I_28363 (I484113,I484507,I484685);
nand I_28364 (I484116,I484637,I484425);
nand I_28365 (I484730,I484247,I177459);
nor I_28366 (I484128,I484490,I484730);
not I_28367 (I484791,I2514);
DFFARX1 I_28368 (I567155,I2507,I484791,I484817,);
DFFARX1 I_28369 (I567158,I2507,I484791,I484834,);
not I_28370 (I484842,I484834);
not I_28371 (I484859,I567155);
nor I_28372 (I484876,I484859,I567167);
not I_28373 (I484893,I567176);
nor I_28374 (I484910,I484876,I567164);
nor I_28375 (I484927,I484834,I484910);
DFFARX1 I_28376 (I484927,I2507,I484791,I484777,);
nor I_28377 (I484958,I567164,I567167);
nand I_28378 (I484975,I484958,I567155);
DFFARX1 I_28379 (I484975,I2507,I484791,I484780,);
nor I_28380 (I485006,I484893,I567164);
nand I_28381 (I485023,I485006,I567170);
nor I_28382 (I485040,I484817,I485023);
DFFARX1 I_28383 (I485040,I2507,I484791,I484756,);
not I_28384 (I485071,I485023);
nand I_28385 (I484768,I484834,I485071);
DFFARX1 I_28386 (I485023,I2507,I484791,I485111,);
not I_28387 (I485119,I485111);
not I_28388 (I485136,I567164);
not I_28389 (I485153,I567161);
nor I_28390 (I485170,I485153,I567176);
nor I_28391 (I484783,I485119,I485170);
nor I_28392 (I485201,I485153,I567173);
and I_28393 (I485218,I485201,I567161);
or I_28394 (I485235,I485218,I567158);
DFFARX1 I_28395 (I485235,I2507,I484791,I485261,);
nor I_28396 (I484771,I485261,I484817);
not I_28397 (I485283,I485261);
and I_28398 (I485300,I485283,I484817);
nor I_28399 (I484765,I484842,I485300);
nand I_28400 (I485331,I485283,I484893);
nor I_28401 (I484759,I485153,I485331);
nand I_28402 (I484762,I485283,I485071);
nand I_28403 (I485376,I484893,I567161);
nor I_28404 (I484774,I485136,I485376);
not I_28405 (I485437,I2514);
DFFARX1 I_28406 (I359965,I2507,I485437,I485463,);
DFFARX1 I_28407 (I359959,I2507,I485437,I485480,);
not I_28408 (I485488,I485480);
not I_28409 (I485505,I359974);
nor I_28410 (I485522,I485505,I359959);
not I_28411 (I485539,I359968);
nor I_28412 (I485556,I485522,I359977);
nor I_28413 (I485573,I485480,I485556);
DFFARX1 I_28414 (I485573,I2507,I485437,I485423,);
nor I_28415 (I485604,I359977,I359959);
nand I_28416 (I485621,I485604,I359974);
DFFARX1 I_28417 (I485621,I2507,I485437,I485426,);
nor I_28418 (I485652,I485539,I359977);
nand I_28419 (I485669,I485652,I359962);
nor I_28420 (I485686,I485463,I485669);
DFFARX1 I_28421 (I485686,I2507,I485437,I485402,);
not I_28422 (I485717,I485669);
nand I_28423 (I485414,I485480,I485717);
DFFARX1 I_28424 (I485669,I2507,I485437,I485757,);
not I_28425 (I485765,I485757);
not I_28426 (I485782,I359977);
not I_28427 (I485799,I359971);
nor I_28428 (I485816,I485799,I359968);
nor I_28429 (I485429,I485765,I485816);
nor I_28430 (I485847,I485799,I359980);
and I_28431 (I485864,I485847,I359983);
or I_28432 (I485881,I485864,I359962);
DFFARX1 I_28433 (I485881,I2507,I485437,I485907,);
nor I_28434 (I485417,I485907,I485463);
not I_28435 (I485929,I485907);
and I_28436 (I485946,I485929,I485463);
nor I_28437 (I485411,I485488,I485946);
nand I_28438 (I485977,I485929,I485539);
nor I_28439 (I485405,I485799,I485977);
nand I_28440 (I485408,I485929,I485717);
nand I_28441 (I486022,I485539,I359971);
nor I_28442 (I485420,I485782,I486022);
not I_28443 (I486083,I2514);
DFFARX1 I_28444 (I79408,I2507,I486083,I486109,);
DFFARX1 I_28445 (I79414,I2507,I486083,I486126,);
not I_28446 (I486134,I486126);
not I_28447 (I486151,I79432);
nor I_28448 (I486168,I486151,I79411);
not I_28449 (I486185,I79417);
nor I_28450 (I486202,I486168,I79423);
nor I_28451 (I486219,I486126,I486202);
DFFARX1 I_28452 (I486219,I2507,I486083,I486069,);
nor I_28453 (I486250,I79423,I79411);
nand I_28454 (I486267,I486250,I79432);
DFFARX1 I_28455 (I486267,I2507,I486083,I486072,);
nor I_28456 (I486298,I486185,I79423);
nand I_28457 (I486315,I486298,I79429);
nor I_28458 (I486332,I486109,I486315);
DFFARX1 I_28459 (I486332,I2507,I486083,I486048,);
not I_28460 (I486363,I486315);
nand I_28461 (I486060,I486126,I486363);
DFFARX1 I_28462 (I486315,I2507,I486083,I486403,);
not I_28463 (I486411,I486403);
not I_28464 (I486428,I79423);
not I_28465 (I486445,I79411);
nor I_28466 (I486462,I486445,I79417);
nor I_28467 (I486075,I486411,I486462);
nor I_28468 (I486493,I486445,I79420);
and I_28469 (I486510,I486493,I79408);
or I_28470 (I486527,I486510,I79426);
DFFARX1 I_28471 (I486527,I2507,I486083,I486553,);
nor I_28472 (I486063,I486553,I486109);
not I_28473 (I486575,I486553);
and I_28474 (I486592,I486575,I486109);
nor I_28475 (I486057,I486134,I486592);
nand I_28476 (I486623,I486575,I486185);
nor I_28477 (I486051,I486445,I486623);
nand I_28478 (I486054,I486575,I486363);
nand I_28479 (I486668,I486185,I79411);
nor I_28480 (I486066,I486428,I486668);
not I_28481 (I486729,I2514);
DFFARX1 I_28482 (I438131,I2507,I486729,I486755,);
DFFARX1 I_28483 (I438128,I2507,I486729,I486772,);
not I_28484 (I486780,I486772);
not I_28485 (I486797,I438128);
nor I_28486 (I486814,I486797,I438131);
not I_28487 (I486831,I438143);
nor I_28488 (I486848,I486814,I438137);
nor I_28489 (I486865,I486772,I486848);
DFFARX1 I_28490 (I486865,I2507,I486729,I486715,);
nor I_28491 (I486896,I438137,I438131);
nand I_28492 (I486913,I486896,I438128);
DFFARX1 I_28493 (I486913,I2507,I486729,I486718,);
nor I_28494 (I486944,I486831,I438137);
nand I_28495 (I486961,I486944,I438125);
nor I_28496 (I486978,I486755,I486961);
DFFARX1 I_28497 (I486978,I2507,I486729,I486694,);
not I_28498 (I487009,I486961);
nand I_28499 (I486706,I486772,I487009);
DFFARX1 I_28500 (I486961,I2507,I486729,I487049,);
not I_28501 (I487057,I487049);
not I_28502 (I487074,I438137);
not I_28503 (I487091,I438134);
nor I_28504 (I487108,I487091,I438143);
nor I_28505 (I486721,I487057,I487108);
nor I_28506 (I487139,I487091,I438140);
and I_28507 (I487156,I487139,I438146);
or I_28508 (I487173,I487156,I438125);
DFFARX1 I_28509 (I487173,I2507,I486729,I487199,);
nor I_28510 (I486709,I487199,I486755);
not I_28511 (I487221,I487199);
and I_28512 (I487238,I487221,I486755);
nor I_28513 (I486703,I486780,I487238);
nand I_28514 (I487269,I487221,I486831);
nor I_28515 (I486697,I487091,I487269);
nand I_28516 (I486700,I487221,I487009);
nand I_28517 (I487314,I486831,I438134);
nor I_28518 (I486712,I487074,I487314);
not I_28519 (I487375,I2514);
DFFARX1 I_28520 (I364589,I2507,I487375,I487401,);
DFFARX1 I_28521 (I364583,I2507,I487375,I487418,);
not I_28522 (I487426,I487418);
not I_28523 (I487443,I364598);
nor I_28524 (I487460,I487443,I364583);
not I_28525 (I487477,I364592);
nor I_28526 (I487494,I487460,I364601);
nor I_28527 (I487511,I487418,I487494);
DFFARX1 I_28528 (I487511,I2507,I487375,I487361,);
nor I_28529 (I487542,I364601,I364583);
nand I_28530 (I487559,I487542,I364598);
DFFARX1 I_28531 (I487559,I2507,I487375,I487364,);
nor I_28532 (I487590,I487477,I364601);
nand I_28533 (I487607,I487590,I364586);
nor I_28534 (I487624,I487401,I487607);
DFFARX1 I_28535 (I487624,I2507,I487375,I487340,);
not I_28536 (I487655,I487607);
nand I_28537 (I487352,I487418,I487655);
DFFARX1 I_28538 (I487607,I2507,I487375,I487695,);
not I_28539 (I487703,I487695);
not I_28540 (I487720,I364601);
not I_28541 (I487737,I364595);
nor I_28542 (I487754,I487737,I364592);
nor I_28543 (I487367,I487703,I487754);
nor I_28544 (I487785,I487737,I364604);
and I_28545 (I487802,I487785,I364607);
or I_28546 (I487819,I487802,I364586);
DFFARX1 I_28547 (I487819,I2507,I487375,I487845,);
nor I_28548 (I487355,I487845,I487401);
not I_28549 (I487867,I487845);
and I_28550 (I487884,I487867,I487401);
nor I_28551 (I487349,I487426,I487884);
nand I_28552 (I487915,I487867,I487477);
nor I_28553 (I487343,I487737,I487915);
nand I_28554 (I487346,I487867,I487655);
nand I_28555 (I487960,I487477,I364595);
nor I_28556 (I487358,I487720,I487960);
not I_28557 (I488021,I2514);
DFFARX1 I_28558 (I135990,I2507,I488021,I488047,);
DFFARX1 I_28559 (I136002,I2507,I488021,I488064,);
not I_28560 (I488072,I488064);
not I_28561 (I488089,I136008);
nor I_28562 (I488106,I488089,I135993);
not I_28563 (I488123,I135984);
nor I_28564 (I488140,I488106,I136005);
nor I_28565 (I488157,I488064,I488140);
DFFARX1 I_28566 (I488157,I2507,I488021,I488007,);
nor I_28567 (I488188,I136005,I135993);
nand I_28568 (I488205,I488188,I136008);
DFFARX1 I_28569 (I488205,I2507,I488021,I488010,);
nor I_28570 (I488236,I488123,I136005);
nand I_28571 (I488253,I488236,I135987);
nor I_28572 (I488270,I488047,I488253);
DFFARX1 I_28573 (I488270,I2507,I488021,I487986,);
not I_28574 (I488301,I488253);
nand I_28575 (I487998,I488064,I488301);
DFFARX1 I_28576 (I488253,I2507,I488021,I488341,);
not I_28577 (I488349,I488341);
not I_28578 (I488366,I136005);
not I_28579 (I488383,I135996);
nor I_28580 (I488400,I488383,I135984);
nor I_28581 (I488013,I488349,I488400);
nor I_28582 (I488431,I488383,I135999);
and I_28583 (I488448,I488431,I135987);
or I_28584 (I488465,I488448,I135984);
DFFARX1 I_28585 (I488465,I2507,I488021,I488491,);
nor I_28586 (I488001,I488491,I488047);
not I_28587 (I488513,I488491);
and I_28588 (I488530,I488513,I488047);
nor I_28589 (I487995,I488072,I488530);
nand I_28590 (I488561,I488513,I488123);
nor I_28591 (I487989,I488383,I488561);
nand I_28592 (I487992,I488513,I488301);
nand I_28593 (I488606,I488123,I135996);
nor I_28594 (I488004,I488366,I488606);
not I_28595 (I488667,I2514);
DFFARX1 I_28596 (I601173,I2507,I488667,I488693,);
DFFARX1 I_28597 (I601155,I2507,I488667,I488710,);
not I_28598 (I488718,I488710);
not I_28599 (I488735,I601164);
nor I_28600 (I488752,I488735,I601176);
not I_28601 (I488769,I601158);
nor I_28602 (I488786,I488752,I601167);
nor I_28603 (I488803,I488710,I488786);
DFFARX1 I_28604 (I488803,I2507,I488667,I488653,);
nor I_28605 (I488834,I601167,I601176);
nand I_28606 (I488851,I488834,I601164);
DFFARX1 I_28607 (I488851,I2507,I488667,I488656,);
nor I_28608 (I488882,I488769,I601167);
nand I_28609 (I488899,I488882,I601179);
nor I_28610 (I488916,I488693,I488899);
DFFARX1 I_28611 (I488916,I2507,I488667,I488632,);
not I_28612 (I488947,I488899);
nand I_28613 (I488644,I488710,I488947);
DFFARX1 I_28614 (I488899,I2507,I488667,I488987,);
not I_28615 (I488995,I488987);
not I_28616 (I489012,I601167);
not I_28617 (I489029,I601155);
nor I_28618 (I489046,I489029,I601158);
nor I_28619 (I488659,I488995,I489046);
nor I_28620 (I489077,I489029,I601161);
and I_28621 (I489094,I489077,I601170);
or I_28622 (I489111,I489094,I601158);
DFFARX1 I_28623 (I489111,I2507,I488667,I489137,);
nor I_28624 (I488647,I489137,I488693);
not I_28625 (I489159,I489137);
and I_28626 (I489176,I489159,I488693);
nor I_28627 (I488641,I488718,I489176);
nand I_28628 (I489207,I489159,I488769);
nor I_28629 (I488635,I489029,I489207);
nand I_28630 (I488638,I489159,I488947);
nand I_28631 (I489252,I488769,I601155);
nor I_28632 (I488650,I489012,I489252);
not I_28633 (I489313,I2514);
DFFARX1 I_28634 (I462900,I2507,I489313,I489339,);
DFFARX1 I_28635 (I462897,I2507,I489313,I489356,);
not I_28636 (I489364,I489356);
not I_28637 (I489381,I462897);
nor I_28638 (I489398,I489381,I462900);
not I_28639 (I489415,I462912);
nor I_28640 (I489432,I489398,I462906);
nor I_28641 (I489449,I489356,I489432);
DFFARX1 I_28642 (I489449,I2507,I489313,I489299,);
nor I_28643 (I489480,I462906,I462900);
nand I_28644 (I489497,I489480,I462897);
DFFARX1 I_28645 (I489497,I2507,I489313,I489302,);
nor I_28646 (I489528,I489415,I462906);
nand I_28647 (I489545,I489528,I462894);
nor I_28648 (I489562,I489339,I489545);
DFFARX1 I_28649 (I489562,I2507,I489313,I489278,);
not I_28650 (I489593,I489545);
nand I_28651 (I489290,I489356,I489593);
DFFARX1 I_28652 (I489545,I2507,I489313,I489633,);
not I_28653 (I489641,I489633);
not I_28654 (I489658,I462906);
not I_28655 (I489675,I462903);
nor I_28656 (I489692,I489675,I462912);
nor I_28657 (I489305,I489641,I489692);
nor I_28658 (I489723,I489675,I462909);
and I_28659 (I489740,I489723,I462915);
or I_28660 (I489757,I489740,I462894);
DFFARX1 I_28661 (I489757,I2507,I489313,I489783,);
nor I_28662 (I489293,I489783,I489339);
not I_28663 (I489805,I489783);
and I_28664 (I489822,I489805,I489339);
nor I_28665 (I489287,I489364,I489822);
nand I_28666 (I489853,I489805,I489415);
nor I_28667 (I489281,I489675,I489853);
nand I_28668 (I489284,I489805,I489593);
nand I_28669 (I489898,I489415,I462903);
nor I_28670 (I489296,I489658,I489898);
not I_28671 (I489959,I2514);
DFFARX1 I_28672 (I649079,I2507,I489959,I489985,);
DFFARX1 I_28673 (I649085,I2507,I489959,I490002,);
not I_28674 (I490010,I490002);
not I_28675 (I490027,I649082);
nor I_28676 (I490044,I490027,I649061);
not I_28677 (I490061,I649064);
nor I_28678 (I490078,I490044,I649070);
nor I_28679 (I490095,I490002,I490078);
DFFARX1 I_28680 (I490095,I2507,I489959,I489945,);
nor I_28681 (I490126,I649070,I649061);
nand I_28682 (I490143,I490126,I649082);
DFFARX1 I_28683 (I490143,I2507,I489959,I489948,);
nor I_28684 (I490174,I490061,I649070);
nand I_28685 (I490191,I490174,I649064);
nor I_28686 (I490208,I489985,I490191);
DFFARX1 I_28687 (I490208,I2507,I489959,I489924,);
not I_28688 (I490239,I490191);
nand I_28689 (I489936,I490002,I490239);
DFFARX1 I_28690 (I490191,I2507,I489959,I490279,);
not I_28691 (I490287,I490279);
not I_28692 (I490304,I649070);
not I_28693 (I490321,I649073);
nor I_28694 (I490338,I490321,I649064);
nor I_28695 (I489951,I490287,I490338);
nor I_28696 (I490369,I490321,I649061);
and I_28697 (I490386,I490369,I649067);
or I_28698 (I490403,I490386,I649076);
DFFARX1 I_28699 (I490403,I2507,I489959,I490429,);
nor I_28700 (I489939,I490429,I489985);
not I_28701 (I490451,I490429);
and I_28702 (I490468,I490451,I489985);
nor I_28703 (I489933,I490010,I490468);
nand I_28704 (I490499,I490451,I490061);
nor I_28705 (I489927,I490321,I490499);
nand I_28706 (I489930,I490451,I490239);
nand I_28707 (I490544,I490061,I649073);
nor I_28708 (I489942,I490304,I490544);
not I_28709 (I490605,I2514);
DFFARX1 I_28710 (I18276,I2507,I490605,I490631,);
DFFARX1 I_28711 (I18282,I2507,I490605,I490648,);
not I_28712 (I490656,I490648);
not I_28713 (I490673,I18276);
nor I_28714 (I490690,I490673,I18288);
not I_28715 (I490707,I18300);
nor I_28716 (I490724,I490690,I18294);
nor I_28717 (I490741,I490648,I490724);
DFFARX1 I_28718 (I490741,I2507,I490605,I490591,);
nor I_28719 (I490772,I18294,I18288);
nand I_28720 (I490789,I490772,I18276);
DFFARX1 I_28721 (I490789,I2507,I490605,I490594,);
nor I_28722 (I490820,I490707,I18294);
nand I_28723 (I490837,I490820,I18279);
nor I_28724 (I490854,I490631,I490837);
DFFARX1 I_28725 (I490854,I2507,I490605,I490570,);
not I_28726 (I490885,I490837);
nand I_28727 (I490582,I490648,I490885);
DFFARX1 I_28728 (I490837,I2507,I490605,I490925,);
not I_28729 (I490933,I490925);
not I_28730 (I490950,I18294);
not I_28731 (I490967,I18279);
nor I_28732 (I490984,I490967,I18300);
nor I_28733 (I490597,I490933,I490984);
nor I_28734 (I491015,I490967,I18297);
and I_28735 (I491032,I491015,I18291);
or I_28736 (I491049,I491032,I18285);
DFFARX1 I_28737 (I491049,I2507,I490605,I491075,);
nor I_28738 (I490585,I491075,I490631);
not I_28739 (I491097,I491075);
and I_28740 (I491114,I491097,I490631);
nor I_28741 (I490579,I490656,I491114);
nand I_28742 (I491145,I491097,I490707);
nor I_28743 (I490573,I490967,I491145);
nand I_28744 (I490576,I491097,I490885);
nand I_28745 (I491190,I490707,I18279);
nor I_28746 (I490588,I490950,I491190);
not I_28747 (I491251,I2514);
DFFARX1 I_28748 (I281371,I2507,I491251,I491277,);
DFFARX1 I_28749 (I281383,I2507,I491251,I491294,);
not I_28750 (I491302,I491294);
not I_28751 (I491319,I281368);
nor I_28752 (I491336,I491319,I281386);
not I_28753 (I491353,I281392);
nor I_28754 (I491370,I491336,I281374);
nor I_28755 (I491387,I491294,I491370);
DFFARX1 I_28756 (I491387,I2507,I491251,I491237,);
nor I_28757 (I491418,I281374,I281386);
nand I_28758 (I491435,I491418,I281368);
DFFARX1 I_28759 (I491435,I2507,I491251,I491240,);
nor I_28760 (I491466,I491353,I281374);
nand I_28761 (I491483,I491466,I281377);
nor I_28762 (I491500,I491277,I491483);
DFFARX1 I_28763 (I491500,I2507,I491251,I491216,);
not I_28764 (I491531,I491483);
nand I_28765 (I491228,I491294,I491531);
DFFARX1 I_28766 (I491483,I2507,I491251,I491571,);
not I_28767 (I491579,I491571);
not I_28768 (I491596,I281374);
not I_28769 (I491613,I281380);
nor I_28770 (I491630,I491613,I281392);
nor I_28771 (I491243,I491579,I491630);
nor I_28772 (I491661,I491613,I281389);
and I_28773 (I491678,I491661,I281368);
or I_28774 (I491695,I491678,I281371);
DFFARX1 I_28775 (I491695,I2507,I491251,I491721,);
nor I_28776 (I491231,I491721,I491277);
not I_28777 (I491743,I491721);
and I_28778 (I491760,I491743,I491277);
nor I_28779 (I491225,I491302,I491760);
nand I_28780 (I491791,I491743,I491353);
nor I_28781 (I491219,I491613,I491791);
nand I_28782 (I491222,I491743,I491531);
nand I_28783 (I491836,I491353,I281380);
nor I_28784 (I491234,I491596,I491836);
not I_28785 (I491897,I2514);
DFFARX1 I_28786 (I697188,I2507,I491897,I491923,);
DFFARX1 I_28787 (I697212,I2507,I491897,I491940,);
not I_28788 (I491948,I491940);
not I_28789 (I491965,I697194);
nor I_28790 (I491982,I491965,I697203);
not I_28791 (I491999,I697188);
nor I_28792 (I492016,I491982,I697209);
nor I_28793 (I492033,I491940,I492016);
DFFARX1 I_28794 (I492033,I2507,I491897,I491883,);
nor I_28795 (I492064,I697209,I697203);
nand I_28796 (I492081,I492064,I697194);
DFFARX1 I_28797 (I492081,I2507,I491897,I491886,);
nor I_28798 (I492112,I491999,I697209);
nand I_28799 (I492129,I492112,I697206);
nor I_28800 (I492146,I491923,I492129);
DFFARX1 I_28801 (I492146,I2507,I491897,I491862,);
not I_28802 (I492177,I492129);
nand I_28803 (I491874,I491940,I492177);
DFFARX1 I_28804 (I492129,I2507,I491897,I492217,);
not I_28805 (I492225,I492217);
not I_28806 (I492242,I697209);
not I_28807 (I492259,I697200);
nor I_28808 (I492276,I492259,I697188);
nor I_28809 (I491889,I492225,I492276);
nor I_28810 (I492307,I492259,I697191);
and I_28811 (I492324,I492307,I697215);
or I_28812 (I492341,I492324,I697197);
DFFARX1 I_28813 (I492341,I2507,I491897,I492367,);
nor I_28814 (I491877,I492367,I491923);
not I_28815 (I492389,I492367);
and I_28816 (I492406,I492389,I491923);
nor I_28817 (I491871,I491948,I492406);
nand I_28818 (I492437,I492389,I491999);
nor I_28819 (I491865,I492259,I492437);
nand I_28820 (I491868,I492389,I492177);
nand I_28821 (I492482,I491999,I697200);
nor I_28822 (I491880,I492242,I492482);
not I_28823 (I492543,I2514);
DFFARX1 I_28824 (I322970,I2507,I492543,I492569,);
DFFARX1 I_28825 (I322982,I2507,I492543,I492586,);
not I_28826 (I492594,I492586);
not I_28827 (I492611,I322991);
nor I_28828 (I492628,I492611,I322967);
not I_28829 (I492645,I322985);
nor I_28830 (I492662,I492628,I322979);
nor I_28831 (I492679,I492586,I492662);
DFFARX1 I_28832 (I492679,I2507,I492543,I492529,);
nor I_28833 (I492710,I322979,I322967);
nand I_28834 (I492727,I492710,I322991);
DFFARX1 I_28835 (I492727,I2507,I492543,I492532,);
nor I_28836 (I492758,I492645,I322979);
nand I_28837 (I492775,I492758,I322973);
nor I_28838 (I492792,I492569,I492775);
DFFARX1 I_28839 (I492792,I2507,I492543,I492508,);
not I_28840 (I492823,I492775);
nand I_28841 (I492520,I492586,I492823);
DFFARX1 I_28842 (I492775,I2507,I492543,I492863,);
not I_28843 (I492871,I492863);
not I_28844 (I492888,I322979);
not I_28845 (I492905,I322988);
nor I_28846 (I492922,I492905,I322985);
nor I_28847 (I492535,I492871,I492922);
nor I_28848 (I492953,I492905,I322970);
and I_28849 (I492970,I492953,I322967);
or I_28850 (I492987,I492970,I322976);
DFFARX1 I_28851 (I492987,I2507,I492543,I493013,);
nor I_28852 (I492523,I493013,I492569);
not I_28853 (I493035,I493013);
and I_28854 (I493052,I493035,I492569);
nor I_28855 (I492517,I492594,I493052);
nand I_28856 (I493083,I493035,I492645);
nor I_28857 (I492511,I492905,I493083);
nand I_28858 (I492514,I493035,I492823);
nand I_28859 (I493128,I492645,I322988);
nor I_28860 (I492526,I492888,I493128);
not I_28861 (I493189,I2514);
DFFARX1 I_28862 (I635853,I2507,I493189,I493215,);
DFFARX1 I_28863 (I635835,I2507,I493189,I493232,);
not I_28864 (I493240,I493232);
not I_28865 (I493257,I635844);
nor I_28866 (I493274,I493257,I635856);
not I_28867 (I493291,I635838);
nor I_28868 (I493308,I493274,I635847);
nor I_28869 (I493325,I493232,I493308);
DFFARX1 I_28870 (I493325,I2507,I493189,I493175,);
nor I_28871 (I493356,I635847,I635856);
nand I_28872 (I493373,I493356,I635844);
DFFARX1 I_28873 (I493373,I2507,I493189,I493178,);
nor I_28874 (I493404,I493291,I635847);
nand I_28875 (I493421,I493404,I635859);
nor I_28876 (I493438,I493215,I493421);
DFFARX1 I_28877 (I493438,I2507,I493189,I493154,);
not I_28878 (I493469,I493421);
nand I_28879 (I493166,I493232,I493469);
DFFARX1 I_28880 (I493421,I2507,I493189,I493509,);
not I_28881 (I493517,I493509);
not I_28882 (I493534,I635847);
not I_28883 (I493551,I635835);
nor I_28884 (I493568,I493551,I635838);
nor I_28885 (I493181,I493517,I493568);
nor I_28886 (I493599,I493551,I635841);
and I_28887 (I493616,I493599,I635850);
or I_28888 (I493633,I493616,I635838);
DFFARX1 I_28889 (I493633,I2507,I493189,I493659,);
nor I_28890 (I493169,I493659,I493215);
not I_28891 (I493681,I493659);
and I_28892 (I493698,I493681,I493215);
nor I_28893 (I493163,I493240,I493698);
nand I_28894 (I493729,I493681,I493291);
nor I_28895 (I493157,I493551,I493729);
nand I_28896 (I493160,I493681,I493469);
nand I_28897 (I493774,I493291,I635835);
nor I_28898 (I493172,I493534,I493774);
not I_28899 (I493835,I2514);
DFFARX1 I_28900 (I613311,I2507,I493835,I493861,);
DFFARX1 I_28901 (I613293,I2507,I493835,I493878,);
not I_28902 (I493886,I493878);
not I_28903 (I493903,I613302);
nor I_28904 (I493920,I493903,I613314);
not I_28905 (I493937,I613296);
nor I_28906 (I493954,I493920,I613305);
nor I_28907 (I493971,I493878,I493954);
DFFARX1 I_28908 (I493971,I2507,I493835,I493821,);
nor I_28909 (I494002,I613305,I613314);
nand I_28910 (I494019,I494002,I613302);
DFFARX1 I_28911 (I494019,I2507,I493835,I493824,);
nor I_28912 (I494050,I493937,I613305);
nand I_28913 (I494067,I494050,I613317);
nor I_28914 (I494084,I493861,I494067);
DFFARX1 I_28915 (I494084,I2507,I493835,I493800,);
not I_28916 (I494115,I494067);
nand I_28917 (I493812,I493878,I494115);
DFFARX1 I_28918 (I494067,I2507,I493835,I494155,);
not I_28919 (I494163,I494155);
not I_28920 (I494180,I613305);
not I_28921 (I494197,I613293);
nor I_28922 (I494214,I494197,I613296);
nor I_28923 (I493827,I494163,I494214);
nor I_28924 (I494245,I494197,I613299);
and I_28925 (I494262,I494245,I613308);
or I_28926 (I494279,I494262,I613296);
DFFARX1 I_28927 (I494279,I2507,I493835,I494305,);
nor I_28928 (I493815,I494305,I493861);
not I_28929 (I494327,I494305);
and I_28930 (I494344,I494327,I493861);
nor I_28931 (I493809,I493886,I494344);
nand I_28932 (I494375,I494327,I493937);
nor I_28933 (I493803,I494197,I494375);
nand I_28934 (I493806,I494327,I494115);
nand I_28935 (I494420,I493937,I613293);
nor I_28936 (I493818,I494180,I494420);
not I_28937 (I494481,I2514);
DFFARX1 I_28938 (I208013,I2507,I494481,I494507,);
DFFARX1 I_28939 (I208019,I2507,I494481,I494524,);
not I_28940 (I494532,I494524);
not I_28941 (I494549,I208040);
nor I_28942 (I494566,I494549,I208028);
not I_28943 (I494583,I208037);
nor I_28944 (I494600,I494566,I208022);
nor I_28945 (I494617,I494524,I494600);
DFFARX1 I_28946 (I494617,I2507,I494481,I494467,);
nor I_28947 (I494648,I208022,I208028);
nand I_28948 (I494665,I494648,I208040);
DFFARX1 I_28949 (I494665,I2507,I494481,I494470,);
nor I_28950 (I494696,I494583,I208022);
nand I_28951 (I494713,I494696,I208013);
nor I_28952 (I494730,I494507,I494713);
DFFARX1 I_28953 (I494730,I2507,I494481,I494446,);
not I_28954 (I494761,I494713);
nand I_28955 (I494458,I494524,I494761);
DFFARX1 I_28956 (I494713,I2507,I494481,I494801,);
not I_28957 (I494809,I494801);
not I_28958 (I494826,I208022);
not I_28959 (I494843,I208025);
nor I_28960 (I494860,I494843,I208037);
nor I_28961 (I494473,I494809,I494860);
nor I_28962 (I494891,I494843,I208034);
and I_28963 (I494908,I494891,I208016);
or I_28964 (I494925,I494908,I208031);
DFFARX1 I_28965 (I494925,I2507,I494481,I494951,);
nor I_28966 (I494461,I494951,I494507);
not I_28967 (I494973,I494951);
and I_28968 (I494990,I494973,I494507);
nor I_28969 (I494455,I494532,I494990);
nand I_28970 (I495021,I494973,I494583);
nor I_28971 (I494449,I494843,I495021);
nand I_28972 (I494452,I494973,I494761);
nand I_28973 (I495066,I494583,I208025);
nor I_28974 (I494464,I494826,I495066);
not I_28975 (I495127,I2514);
DFFARX1 I_28976 (I175866,I2507,I495127,I495153,);
DFFARX1 I_28977 (I175872,I2507,I495127,I495170,);
not I_28978 (I495178,I495170);
not I_28979 (I495195,I175893);
nor I_28980 (I495212,I495195,I175881);
not I_28981 (I495229,I175890);
nor I_28982 (I495246,I495212,I175875);
nor I_28983 (I495263,I495170,I495246);
DFFARX1 I_28984 (I495263,I2507,I495127,I495113,);
nor I_28985 (I495294,I175875,I175881);
nand I_28986 (I495311,I495294,I175893);
DFFARX1 I_28987 (I495311,I2507,I495127,I495116,);
nor I_28988 (I495342,I495229,I175875);
nand I_28989 (I495359,I495342,I175866);
nor I_28990 (I495376,I495153,I495359);
DFFARX1 I_28991 (I495376,I2507,I495127,I495092,);
not I_28992 (I495407,I495359);
nand I_28993 (I495104,I495170,I495407);
DFFARX1 I_28994 (I495359,I2507,I495127,I495447,);
not I_28995 (I495455,I495447);
not I_28996 (I495472,I175875);
not I_28997 (I495489,I175878);
nor I_28998 (I495506,I495489,I175890);
nor I_28999 (I495119,I495455,I495506);
nor I_29000 (I495537,I495489,I175887);
and I_29001 (I495554,I495537,I175869);
or I_29002 (I495571,I495554,I175884);
DFFARX1 I_29003 (I495571,I2507,I495127,I495597,);
nor I_29004 (I495107,I495597,I495153);
not I_29005 (I495619,I495597);
and I_29006 (I495636,I495619,I495153);
nor I_29007 (I495101,I495178,I495636);
nand I_29008 (I495667,I495619,I495229);
nor I_29009 (I495095,I495489,I495667);
nand I_29010 (I495098,I495619,I495407);
nand I_29011 (I495712,I495229,I175878);
nor I_29012 (I495110,I495472,I495712);
not I_29013 (I495773,I2514);
DFFARX1 I_29014 (I59382,I2507,I495773,I495799,);
DFFARX1 I_29015 (I59388,I2507,I495773,I495816,);
not I_29016 (I495824,I495816);
not I_29017 (I495841,I59406);
nor I_29018 (I495858,I495841,I59385);
not I_29019 (I495875,I59391);
nor I_29020 (I495892,I495858,I59397);
nor I_29021 (I495909,I495816,I495892);
DFFARX1 I_29022 (I495909,I2507,I495773,I495759,);
nor I_29023 (I495940,I59397,I59385);
nand I_29024 (I495957,I495940,I59406);
DFFARX1 I_29025 (I495957,I2507,I495773,I495762,);
nor I_29026 (I495988,I495875,I59397);
nand I_29027 (I496005,I495988,I59403);
nor I_29028 (I496022,I495799,I496005);
DFFARX1 I_29029 (I496022,I2507,I495773,I495738,);
not I_29030 (I496053,I496005);
nand I_29031 (I495750,I495816,I496053);
DFFARX1 I_29032 (I496005,I2507,I495773,I496093,);
not I_29033 (I496101,I496093);
not I_29034 (I496118,I59397);
not I_29035 (I496135,I59385);
nor I_29036 (I496152,I496135,I59391);
nor I_29037 (I495765,I496101,I496152);
nor I_29038 (I496183,I496135,I59394);
and I_29039 (I496200,I496183,I59382);
or I_29040 (I496217,I496200,I59400);
DFFARX1 I_29041 (I496217,I2507,I495773,I496243,);
nor I_29042 (I495753,I496243,I495799);
not I_29043 (I496265,I496243);
and I_29044 (I496282,I496265,I495799);
nor I_29045 (I495747,I495824,I496282);
nand I_29046 (I496313,I496265,I495875);
nor I_29047 (I495741,I496135,I496313);
nand I_29048 (I495744,I496265,I496053);
nand I_29049 (I496358,I495875,I59385);
nor I_29050 (I495756,I496118,I496358);
not I_29051 (I496419,I2514);
DFFARX1 I_29052 (I78354,I2507,I496419,I496445,);
DFFARX1 I_29053 (I78360,I2507,I496419,I496462,);
not I_29054 (I496470,I496462);
not I_29055 (I496487,I78378);
nor I_29056 (I496504,I496487,I78357);
not I_29057 (I496521,I78363);
nor I_29058 (I496538,I496504,I78369);
nor I_29059 (I496555,I496462,I496538);
DFFARX1 I_29060 (I496555,I2507,I496419,I496405,);
nor I_29061 (I496586,I78369,I78357);
nand I_29062 (I496603,I496586,I78378);
DFFARX1 I_29063 (I496603,I2507,I496419,I496408,);
nor I_29064 (I496634,I496521,I78369);
nand I_29065 (I496651,I496634,I78375);
nor I_29066 (I496668,I496445,I496651);
DFFARX1 I_29067 (I496668,I2507,I496419,I496384,);
not I_29068 (I496699,I496651);
nand I_29069 (I496396,I496462,I496699);
DFFARX1 I_29070 (I496651,I2507,I496419,I496739,);
not I_29071 (I496747,I496739);
not I_29072 (I496764,I78369);
not I_29073 (I496781,I78357);
nor I_29074 (I496798,I496781,I78363);
nor I_29075 (I496411,I496747,I496798);
nor I_29076 (I496829,I496781,I78366);
and I_29077 (I496846,I496829,I78354);
or I_29078 (I496863,I496846,I78372);
DFFARX1 I_29079 (I496863,I2507,I496419,I496889,);
nor I_29080 (I496399,I496889,I496445);
not I_29081 (I496911,I496889);
and I_29082 (I496928,I496911,I496445);
nor I_29083 (I496393,I496470,I496928);
nand I_29084 (I496959,I496911,I496521);
nor I_29085 (I496387,I496781,I496959);
nand I_29086 (I496390,I496911,I496699);
nand I_29087 (I497004,I496521,I78357);
nor I_29088 (I496402,I496764,I497004);
not I_29089 (I497065,I2514);
DFFARX1 I_29090 (I196946,I2507,I497065,I497091,);
DFFARX1 I_29091 (I196952,I2507,I497065,I497108,);
not I_29092 (I497116,I497108);
not I_29093 (I497133,I196973);
nor I_29094 (I497150,I497133,I196961);
not I_29095 (I497167,I196970);
nor I_29096 (I497184,I497150,I196955);
nor I_29097 (I497201,I497108,I497184);
DFFARX1 I_29098 (I497201,I2507,I497065,I497051,);
nor I_29099 (I497232,I196955,I196961);
nand I_29100 (I497249,I497232,I196973);
DFFARX1 I_29101 (I497249,I2507,I497065,I497054,);
nor I_29102 (I497280,I497167,I196955);
nand I_29103 (I497297,I497280,I196946);
nor I_29104 (I497314,I497091,I497297);
DFFARX1 I_29105 (I497314,I2507,I497065,I497030,);
not I_29106 (I497345,I497297);
nand I_29107 (I497042,I497108,I497345);
DFFARX1 I_29108 (I497297,I2507,I497065,I497385,);
not I_29109 (I497393,I497385);
not I_29110 (I497410,I196955);
not I_29111 (I497427,I196958);
nor I_29112 (I497444,I497427,I196970);
nor I_29113 (I497057,I497393,I497444);
nor I_29114 (I497475,I497427,I196967);
and I_29115 (I497492,I497475,I196949);
or I_29116 (I497509,I497492,I196964);
DFFARX1 I_29117 (I497509,I2507,I497065,I497535,);
nor I_29118 (I497045,I497535,I497091);
not I_29119 (I497557,I497535);
and I_29120 (I497574,I497557,I497091);
nor I_29121 (I497039,I497116,I497574);
nand I_29122 (I497605,I497557,I497167);
nor I_29123 (I497033,I497427,I497605);
nand I_29124 (I497036,I497557,I497345);
nand I_29125 (I497650,I497167,I196958);
nor I_29126 (I497048,I497410,I497650);
not I_29127 (I497711,I2514);
DFFARX1 I_29128 (I304474,I2507,I497711,I497737,);
DFFARX1 I_29129 (I304486,I2507,I497711,I497754,);
not I_29130 (I497762,I497754);
not I_29131 (I497779,I304495);
nor I_29132 (I497796,I497779,I304471);
not I_29133 (I497813,I304489);
nor I_29134 (I497830,I497796,I304483);
nor I_29135 (I497847,I497754,I497830);
DFFARX1 I_29136 (I497847,I2507,I497711,I497697,);
nor I_29137 (I497878,I304483,I304471);
nand I_29138 (I497895,I497878,I304495);
DFFARX1 I_29139 (I497895,I2507,I497711,I497700,);
nor I_29140 (I497926,I497813,I304483);
nand I_29141 (I497943,I497926,I304477);
nor I_29142 (I497960,I497737,I497943);
DFFARX1 I_29143 (I497960,I2507,I497711,I497676,);
not I_29144 (I497991,I497943);
nand I_29145 (I497688,I497754,I497991);
DFFARX1 I_29146 (I497943,I2507,I497711,I498031,);
not I_29147 (I498039,I498031);
not I_29148 (I498056,I304483);
not I_29149 (I498073,I304492);
nor I_29150 (I498090,I498073,I304489);
nor I_29151 (I497703,I498039,I498090);
nor I_29152 (I498121,I498073,I304474);
and I_29153 (I498138,I498121,I304471);
or I_29154 (I498155,I498138,I304480);
DFFARX1 I_29155 (I498155,I2507,I497711,I498181,);
nor I_29156 (I497691,I498181,I497737);
not I_29157 (I498203,I498181);
and I_29158 (I498220,I498203,I497737);
nor I_29159 (I497685,I497762,I498220);
nand I_29160 (I498251,I498203,I497813);
nor I_29161 (I497679,I498073,I498251);
nand I_29162 (I497682,I498203,I497991);
nand I_29163 (I498296,I497813,I304492);
nor I_29164 (I497694,I498056,I498296);
not I_29165 (I498357,I2514);
DFFARX1 I_29166 (I640919,I2507,I498357,I498383,);
DFFARX1 I_29167 (I640925,I2507,I498357,I498400,);
not I_29168 (I498408,I498400);
not I_29169 (I498425,I640922);
nor I_29170 (I498442,I498425,I640901);
not I_29171 (I498459,I640904);
nor I_29172 (I498476,I498442,I640910);
nor I_29173 (I498493,I498400,I498476);
DFFARX1 I_29174 (I498493,I2507,I498357,I498343,);
nor I_29175 (I498524,I640910,I640901);
nand I_29176 (I498541,I498524,I640922);
DFFARX1 I_29177 (I498541,I2507,I498357,I498346,);
nor I_29178 (I498572,I498459,I640910);
nand I_29179 (I498589,I498572,I640904);
nor I_29180 (I498606,I498383,I498589);
DFFARX1 I_29181 (I498606,I2507,I498357,I498322,);
not I_29182 (I498637,I498589);
nand I_29183 (I498334,I498400,I498637);
DFFARX1 I_29184 (I498589,I2507,I498357,I498677,);
not I_29185 (I498685,I498677);
not I_29186 (I498702,I640910);
not I_29187 (I498719,I640913);
nor I_29188 (I498736,I498719,I640904);
nor I_29189 (I498349,I498685,I498736);
nor I_29190 (I498767,I498719,I640901);
and I_29191 (I498784,I498767,I640907);
or I_29192 (I498801,I498784,I640916);
DFFARX1 I_29193 (I498801,I2507,I498357,I498827,);
nor I_29194 (I498337,I498827,I498383);
not I_29195 (I498849,I498827);
and I_29196 (I498866,I498849,I498383);
nor I_29197 (I498331,I498408,I498866);
nand I_29198 (I498897,I498849,I498459);
nor I_29199 (I498325,I498719,I498897);
nand I_29200 (I498328,I498849,I498637);
nand I_29201 (I498942,I498459,I640913);
nor I_29202 (I498340,I498702,I498942);
not I_29203 (I499003,I2514);
DFFARX1 I_29204 (I285536,I2507,I499003,I499029,);
DFFARX1 I_29205 (I285548,I2507,I499003,I499046,);
not I_29206 (I499054,I499046);
not I_29207 (I499071,I285533);
nor I_29208 (I499088,I499071,I285551);
not I_29209 (I499105,I285557);
nor I_29210 (I499122,I499088,I285539);
nor I_29211 (I499139,I499046,I499122);
DFFARX1 I_29212 (I499139,I2507,I499003,I498989,);
nor I_29213 (I499170,I285539,I285551);
nand I_29214 (I499187,I499170,I285533);
DFFARX1 I_29215 (I499187,I2507,I499003,I498992,);
nor I_29216 (I499218,I499105,I285539);
nand I_29217 (I499235,I499218,I285542);
nor I_29218 (I499252,I499029,I499235);
DFFARX1 I_29219 (I499252,I2507,I499003,I498968,);
not I_29220 (I499283,I499235);
nand I_29221 (I498980,I499046,I499283);
DFFARX1 I_29222 (I499235,I2507,I499003,I499323,);
not I_29223 (I499331,I499323);
not I_29224 (I499348,I285539);
not I_29225 (I499365,I285545);
nor I_29226 (I499382,I499365,I285557);
nor I_29227 (I498995,I499331,I499382);
nor I_29228 (I499413,I499365,I285554);
and I_29229 (I499430,I499413,I285533);
or I_29230 (I499447,I499430,I285536);
DFFARX1 I_29231 (I499447,I2507,I499003,I499473,);
nor I_29232 (I498983,I499473,I499029);
not I_29233 (I499495,I499473);
and I_29234 (I499512,I499495,I499029);
nor I_29235 (I498977,I499054,I499512);
nand I_29236 (I499543,I499495,I499105);
nor I_29237 (I498971,I499365,I499543);
nand I_29238 (I498974,I499495,I499283);
nand I_29239 (I499588,I499105,I285545);
nor I_29240 (I498986,I499348,I499588);
not I_29241 (I499649,I2514);
DFFARX1 I_29242 (I222242,I2507,I499649,I499675,);
DFFARX1 I_29243 (I222248,I2507,I499649,I499692,);
not I_29244 (I499700,I499692);
not I_29245 (I499717,I222269);
nor I_29246 (I499734,I499717,I222257);
not I_29247 (I499751,I222266);
nor I_29248 (I499768,I499734,I222251);
nor I_29249 (I499785,I499692,I499768);
DFFARX1 I_29250 (I499785,I2507,I499649,I499635,);
nor I_29251 (I499816,I222251,I222257);
nand I_29252 (I499833,I499816,I222269);
DFFARX1 I_29253 (I499833,I2507,I499649,I499638,);
nor I_29254 (I499864,I499751,I222251);
nand I_29255 (I499881,I499864,I222242);
nor I_29256 (I499898,I499675,I499881);
DFFARX1 I_29257 (I499898,I2507,I499649,I499614,);
not I_29258 (I499929,I499881);
nand I_29259 (I499626,I499692,I499929);
DFFARX1 I_29260 (I499881,I2507,I499649,I499969,);
not I_29261 (I499977,I499969);
not I_29262 (I499994,I222251);
not I_29263 (I500011,I222254);
nor I_29264 (I500028,I500011,I222266);
nor I_29265 (I499641,I499977,I500028);
nor I_29266 (I500059,I500011,I222263);
and I_29267 (I500076,I500059,I222245);
or I_29268 (I500093,I500076,I222260);
DFFARX1 I_29269 (I500093,I2507,I499649,I500119,);
nor I_29270 (I499629,I500119,I499675);
not I_29271 (I500141,I500119);
and I_29272 (I500158,I500141,I499675);
nor I_29273 (I499623,I499700,I500158);
nand I_29274 (I500189,I500141,I499751);
nor I_29275 (I499617,I500011,I500189);
nand I_29276 (I499620,I500141,I499929);
nand I_29277 (I500234,I499751,I222254);
nor I_29278 (I499632,I499994,I500234);
not I_29279 (I500295,I2514);
DFFARX1 I_29280 (I710278,I2507,I500295,I500321,);
DFFARX1 I_29281 (I710302,I2507,I500295,I500338,);
not I_29282 (I500346,I500338);
not I_29283 (I500363,I710284);
nor I_29284 (I500380,I500363,I710293);
not I_29285 (I500397,I710278);
nor I_29286 (I500414,I500380,I710299);
nor I_29287 (I500431,I500338,I500414);
DFFARX1 I_29288 (I500431,I2507,I500295,I500281,);
nor I_29289 (I500462,I710299,I710293);
nand I_29290 (I500479,I500462,I710284);
DFFARX1 I_29291 (I500479,I2507,I500295,I500284,);
nor I_29292 (I500510,I500397,I710299);
nand I_29293 (I500527,I500510,I710296);
nor I_29294 (I500544,I500321,I500527);
DFFARX1 I_29295 (I500544,I2507,I500295,I500260,);
not I_29296 (I500575,I500527);
nand I_29297 (I500272,I500338,I500575);
DFFARX1 I_29298 (I500527,I2507,I500295,I500615,);
not I_29299 (I500623,I500615);
not I_29300 (I500640,I710299);
not I_29301 (I500657,I710290);
nor I_29302 (I500674,I500657,I710278);
nor I_29303 (I500287,I500623,I500674);
nor I_29304 (I500705,I500657,I710281);
and I_29305 (I500722,I500705,I710305);
or I_29306 (I500739,I500722,I710287);
DFFARX1 I_29307 (I500739,I2507,I500295,I500765,);
nor I_29308 (I500275,I500765,I500321);
not I_29309 (I500787,I500765);
and I_29310 (I500804,I500787,I500321);
nor I_29311 (I500269,I500346,I500804);
nand I_29312 (I500835,I500787,I500397);
nor I_29313 (I500263,I500657,I500835);
nand I_29314 (I500266,I500787,I500575);
nand I_29315 (I500880,I500397,I710290);
nor I_29316 (I500278,I500640,I500880);
not I_29317 (I500941,I2514);
DFFARX1 I_29318 (I600595,I2507,I500941,I500967,);
DFFARX1 I_29319 (I600577,I2507,I500941,I500984,);
not I_29320 (I500992,I500984);
not I_29321 (I501009,I600586);
nor I_29322 (I501026,I501009,I600598);
not I_29323 (I501043,I600580);
nor I_29324 (I501060,I501026,I600589);
nor I_29325 (I501077,I500984,I501060);
DFFARX1 I_29326 (I501077,I2507,I500941,I500927,);
nor I_29327 (I501108,I600589,I600598);
nand I_29328 (I501125,I501108,I600586);
DFFARX1 I_29329 (I501125,I2507,I500941,I500930,);
nor I_29330 (I501156,I501043,I600589);
nand I_29331 (I501173,I501156,I600601);
nor I_29332 (I501190,I500967,I501173);
DFFARX1 I_29333 (I501190,I2507,I500941,I500906,);
not I_29334 (I501221,I501173);
nand I_29335 (I500918,I500984,I501221);
DFFARX1 I_29336 (I501173,I2507,I500941,I501261,);
not I_29337 (I501269,I501261);
not I_29338 (I501286,I600589);
not I_29339 (I501303,I600577);
nor I_29340 (I501320,I501303,I600580);
nor I_29341 (I500933,I501269,I501320);
nor I_29342 (I501351,I501303,I600583);
and I_29343 (I501368,I501351,I600592);
or I_29344 (I501385,I501368,I600580);
DFFARX1 I_29345 (I501385,I2507,I500941,I501411,);
nor I_29346 (I500921,I501411,I500967);
not I_29347 (I501433,I501411);
and I_29348 (I501450,I501433,I500967);
nor I_29349 (I500915,I500992,I501450);
nand I_29350 (I501481,I501433,I501043);
nor I_29351 (I500909,I501303,I501481);
nand I_29352 (I500912,I501433,I501221);
nand I_29353 (I501526,I501043,I600577);
nor I_29354 (I500924,I501286,I501526);
not I_29355 (I501587,I2514);
DFFARX1 I_29356 (I224877,I2507,I501587,I501613,);
DFFARX1 I_29357 (I224883,I2507,I501587,I501630,);
not I_29358 (I501638,I501630);
not I_29359 (I501655,I224904);
nor I_29360 (I501672,I501655,I224892);
not I_29361 (I501689,I224901);
nor I_29362 (I501706,I501672,I224886);
nor I_29363 (I501723,I501630,I501706);
DFFARX1 I_29364 (I501723,I2507,I501587,I501573,);
nor I_29365 (I501754,I224886,I224892);
nand I_29366 (I501771,I501754,I224904);
DFFARX1 I_29367 (I501771,I2507,I501587,I501576,);
nor I_29368 (I501802,I501689,I224886);
nand I_29369 (I501819,I501802,I224877);
nor I_29370 (I501836,I501613,I501819);
DFFARX1 I_29371 (I501836,I2507,I501587,I501552,);
not I_29372 (I501867,I501819);
nand I_29373 (I501564,I501630,I501867);
DFFARX1 I_29374 (I501819,I2507,I501587,I501907,);
not I_29375 (I501915,I501907);
not I_29376 (I501932,I224886);
not I_29377 (I501949,I224889);
nor I_29378 (I501966,I501949,I224901);
nor I_29379 (I501579,I501915,I501966);
nor I_29380 (I501997,I501949,I224898);
and I_29381 (I502014,I501997,I224880);
or I_29382 (I502031,I502014,I224895);
DFFARX1 I_29383 (I502031,I2507,I501587,I502057,);
nor I_29384 (I501567,I502057,I501613);
not I_29385 (I502079,I502057);
and I_29386 (I502096,I502079,I501613);
nor I_29387 (I501561,I501638,I502096);
nand I_29388 (I502127,I502079,I501689);
nor I_29389 (I501555,I501949,I502127);
nand I_29390 (I501558,I502079,I501867);
nand I_29391 (I502172,I501689,I224889);
nor I_29392 (I501570,I501932,I502172);
not I_29393 (I502233,I2514);
DFFARX1 I_29394 (I255806,I2507,I502233,I502259,);
DFFARX1 I_29395 (I255803,I2507,I502233,I502276,);
not I_29396 (I502284,I502276);
not I_29397 (I502301,I255818);
nor I_29398 (I502318,I502301,I255821);
not I_29399 (I502335,I255809);
nor I_29400 (I502352,I502318,I255815);
nor I_29401 (I502369,I502276,I502352);
DFFARX1 I_29402 (I502369,I2507,I502233,I502219,);
nor I_29403 (I502400,I255815,I255821);
nand I_29404 (I502417,I502400,I255818);
DFFARX1 I_29405 (I502417,I2507,I502233,I502222,);
nor I_29406 (I502448,I502335,I255815);
nand I_29407 (I502465,I502448,I255827);
nor I_29408 (I502482,I502259,I502465);
DFFARX1 I_29409 (I502482,I2507,I502233,I502198,);
not I_29410 (I502513,I502465);
nand I_29411 (I502210,I502276,I502513);
DFFARX1 I_29412 (I502465,I2507,I502233,I502553,);
not I_29413 (I502561,I502553);
not I_29414 (I502578,I255815);
not I_29415 (I502595,I255800);
nor I_29416 (I502612,I502595,I255809);
nor I_29417 (I502225,I502561,I502612);
nor I_29418 (I502643,I502595,I255812);
and I_29419 (I502660,I502643,I255800);
or I_29420 (I502677,I502660,I255824);
DFFARX1 I_29421 (I502677,I2507,I502233,I502703,);
nor I_29422 (I502213,I502703,I502259);
not I_29423 (I502725,I502703);
and I_29424 (I502742,I502725,I502259);
nor I_29425 (I502207,I502284,I502742);
nand I_29426 (I502773,I502725,I502335);
nor I_29427 (I502201,I502595,I502773);
nand I_29428 (I502204,I502725,I502513);
nand I_29429 (I502818,I502335,I255800);
nor I_29430 (I502216,I502578,I502818);
not I_29431 (I502879,I2514);
DFFARX1 I_29432 (I2204,I2507,I502879,I502905,);
DFFARX1 I_29433 (I2236,I2507,I502879,I502922,);
not I_29434 (I502930,I502922);
not I_29435 (I502947,I2212);
nor I_29436 (I502964,I502947,I2124);
not I_29437 (I502981,I2100);
nor I_29438 (I502998,I502964,I2412);
nor I_29439 (I503015,I502922,I502998);
DFFARX1 I_29440 (I503015,I2507,I502879,I502865,);
nor I_29441 (I503046,I2412,I2124);
nand I_29442 (I503063,I503046,I2212);
DFFARX1 I_29443 (I503063,I2507,I502879,I502868,);
nor I_29444 (I503094,I502981,I2412);
nand I_29445 (I503111,I503094,I1828);
nor I_29446 (I503128,I502905,I503111);
DFFARX1 I_29447 (I503128,I2507,I502879,I502844,);
not I_29448 (I503159,I503111);
nand I_29449 (I502856,I502922,I503159);
DFFARX1 I_29450 (I503111,I2507,I502879,I503199,);
not I_29451 (I503207,I503199);
not I_29452 (I503224,I2412);
not I_29453 (I503241,I2388);
nor I_29454 (I503258,I503241,I2100);
nor I_29455 (I502871,I503207,I503258);
nor I_29456 (I503289,I503241,I2108);
and I_29457 (I503306,I503289,I2500);
or I_29458 (I503323,I503306,I2164);
DFFARX1 I_29459 (I503323,I2507,I502879,I503349,);
nor I_29460 (I502859,I503349,I502905);
not I_29461 (I503371,I503349);
and I_29462 (I503388,I503371,I502905);
nor I_29463 (I502853,I502930,I503388);
nand I_29464 (I503419,I503371,I502981);
nor I_29465 (I502847,I503241,I503419);
nand I_29466 (I502850,I503371,I503159);
nand I_29467 (I503464,I502981,I2388);
nor I_29468 (I502862,I503224,I503464);
not I_29469 (I503525,I2514);
DFFARX1 I_29470 (I545837,I2507,I503525,I503551,);
DFFARX1 I_29471 (I545840,I2507,I503525,I503568,);
not I_29472 (I503576,I503568);
not I_29473 (I503593,I545837);
nor I_29474 (I503610,I503593,I545849);
not I_29475 (I503627,I545858);
nor I_29476 (I503644,I503610,I545846);
nor I_29477 (I503661,I503568,I503644);
DFFARX1 I_29478 (I503661,I2507,I503525,I503511,);
nor I_29479 (I503692,I545846,I545849);
nand I_29480 (I503709,I503692,I545837);
DFFARX1 I_29481 (I503709,I2507,I503525,I503514,);
nor I_29482 (I503740,I503627,I545846);
nand I_29483 (I503757,I503740,I545852);
nor I_29484 (I503774,I503551,I503757);
DFFARX1 I_29485 (I503774,I2507,I503525,I503490,);
not I_29486 (I503805,I503757);
nand I_29487 (I503502,I503568,I503805);
DFFARX1 I_29488 (I503757,I2507,I503525,I503845,);
not I_29489 (I503853,I503845);
not I_29490 (I503870,I545846);
not I_29491 (I503887,I545843);
nor I_29492 (I503904,I503887,I545858);
nor I_29493 (I503517,I503853,I503904);
nor I_29494 (I503935,I503887,I545855);
and I_29495 (I503952,I503935,I545843);
or I_29496 (I503969,I503952,I545840);
DFFARX1 I_29497 (I503969,I2507,I503525,I503995,);
nor I_29498 (I503505,I503995,I503551);
not I_29499 (I504017,I503995);
and I_29500 (I504034,I504017,I503551);
nor I_29501 (I503499,I503576,I504034);
nand I_29502 (I504065,I504017,I503627);
nor I_29503 (I503493,I503887,I504065);
nand I_29504 (I503496,I504017,I503805);
nand I_29505 (I504110,I503627,I545843);
nor I_29506 (I503508,I503870,I504110);
not I_29507 (I504171,I2514);
DFFARX1 I_29508 (I198000,I2507,I504171,I504197,);
DFFARX1 I_29509 (I198006,I2507,I504171,I504214,);
not I_29510 (I504222,I504214);
not I_29511 (I504239,I198027);
nor I_29512 (I504256,I504239,I198015);
not I_29513 (I504273,I198024);
nor I_29514 (I504290,I504256,I198009);
nor I_29515 (I504307,I504214,I504290);
DFFARX1 I_29516 (I504307,I2507,I504171,I504157,);
nor I_29517 (I504338,I198009,I198015);
nand I_29518 (I504355,I504338,I198027);
DFFARX1 I_29519 (I504355,I2507,I504171,I504160,);
nor I_29520 (I504386,I504273,I198009);
nand I_29521 (I504403,I504386,I198000);
nor I_29522 (I504420,I504197,I504403);
DFFARX1 I_29523 (I504420,I2507,I504171,I504136,);
not I_29524 (I504451,I504403);
nand I_29525 (I504148,I504214,I504451);
DFFARX1 I_29526 (I504403,I2507,I504171,I504491,);
not I_29527 (I504499,I504491);
not I_29528 (I504516,I198009);
not I_29529 (I504533,I198012);
nor I_29530 (I504550,I504533,I198024);
nor I_29531 (I504163,I504499,I504550);
nor I_29532 (I504581,I504533,I198021);
and I_29533 (I504598,I504581,I198003);
or I_29534 (I504615,I504598,I198018);
DFFARX1 I_29535 (I504615,I2507,I504171,I504641,);
nor I_29536 (I504151,I504641,I504197);
not I_29537 (I504663,I504641);
and I_29538 (I504680,I504663,I504197);
nor I_29539 (I504145,I504222,I504680);
nand I_29540 (I504711,I504663,I504273);
nor I_29541 (I504139,I504533,I504711);
nand I_29542 (I504142,I504663,I504451);
nand I_29543 (I504756,I504273,I198012);
nor I_29544 (I504154,I504516,I504756);
not I_29545 (I504817,I2514);
DFFARX1 I_29546 (I264510,I2507,I504817,I504843,);
DFFARX1 I_29547 (I264507,I2507,I504817,I504860,);
not I_29548 (I504868,I504860);
not I_29549 (I504885,I264522);
nor I_29550 (I504902,I504885,I264525);
not I_29551 (I504919,I264513);
nor I_29552 (I504936,I504902,I264519);
nor I_29553 (I504953,I504860,I504936);
DFFARX1 I_29554 (I504953,I2507,I504817,I504803,);
nor I_29555 (I504984,I264519,I264525);
nand I_29556 (I505001,I504984,I264522);
DFFARX1 I_29557 (I505001,I2507,I504817,I504806,);
nor I_29558 (I505032,I504919,I264519);
nand I_29559 (I505049,I505032,I264531);
nor I_29560 (I505066,I504843,I505049);
DFFARX1 I_29561 (I505066,I2507,I504817,I504782,);
not I_29562 (I505097,I505049);
nand I_29563 (I504794,I504860,I505097);
DFFARX1 I_29564 (I505049,I2507,I504817,I505137,);
not I_29565 (I505145,I505137);
not I_29566 (I505162,I264519);
not I_29567 (I505179,I264504);
nor I_29568 (I505196,I505179,I264513);
nor I_29569 (I504809,I505145,I505196);
nor I_29570 (I505227,I505179,I264516);
and I_29571 (I505244,I505227,I264504);
or I_29572 (I505261,I505244,I264528);
DFFARX1 I_29573 (I505261,I2507,I504817,I505287,);
nor I_29574 (I504797,I505287,I504843);
not I_29575 (I505309,I505287);
and I_29576 (I505326,I505309,I504843);
nor I_29577 (I504791,I504868,I505326);
nand I_29578 (I505357,I505309,I504919);
nor I_29579 (I504785,I505179,I505357);
nand I_29580 (I504788,I505309,I505097);
nand I_29581 (I505402,I504919,I264504);
nor I_29582 (I504800,I505162,I505402);
not I_29583 (I505463,I2514);
DFFARX1 I_29584 (I405627,I2507,I505463,I505489,);
DFFARX1 I_29585 (I405621,I2507,I505463,I505506,);
not I_29586 (I505514,I505506);
not I_29587 (I505531,I405636);
nor I_29588 (I505548,I505531,I405621);
not I_29589 (I505565,I405630);
nor I_29590 (I505582,I505548,I405639);
nor I_29591 (I505599,I505506,I505582);
DFFARX1 I_29592 (I505599,I2507,I505463,I505449,);
nor I_29593 (I505630,I405639,I405621);
nand I_29594 (I505647,I505630,I405636);
DFFARX1 I_29595 (I505647,I2507,I505463,I505452,);
nor I_29596 (I505678,I505565,I405639);
nand I_29597 (I505695,I505678,I405624);
nor I_29598 (I505712,I505489,I505695);
DFFARX1 I_29599 (I505712,I2507,I505463,I505428,);
not I_29600 (I505743,I505695);
nand I_29601 (I505440,I505506,I505743);
DFFARX1 I_29602 (I505695,I2507,I505463,I505783,);
not I_29603 (I505791,I505783);
not I_29604 (I505808,I405639);
not I_29605 (I505825,I405633);
nor I_29606 (I505842,I505825,I405630);
nor I_29607 (I505455,I505791,I505842);
nor I_29608 (I505873,I505825,I405642);
and I_29609 (I505890,I505873,I405645);
or I_29610 (I505907,I505890,I405624);
DFFARX1 I_29611 (I505907,I2507,I505463,I505933,);
nor I_29612 (I505443,I505933,I505489);
not I_29613 (I505955,I505933);
and I_29614 (I505972,I505955,I505489);
nor I_29615 (I505437,I505514,I505972);
nand I_29616 (I506003,I505955,I505565);
nor I_29617 (I505431,I505825,I506003);
nand I_29618 (I505434,I505955,I505743);
nand I_29619 (I506048,I505565,I405633);
nor I_29620 (I505446,I505808,I506048);
not I_29621 (I506109,I2514);
DFFARX1 I_29622 (I449725,I2507,I506109,I506135,);
DFFARX1 I_29623 (I449722,I2507,I506109,I506152,);
not I_29624 (I506160,I506152);
not I_29625 (I506177,I449722);
nor I_29626 (I506194,I506177,I449725);
not I_29627 (I506211,I449737);
nor I_29628 (I506228,I506194,I449731);
nor I_29629 (I506245,I506152,I506228);
DFFARX1 I_29630 (I506245,I2507,I506109,I506095,);
nor I_29631 (I506276,I449731,I449725);
nand I_29632 (I506293,I506276,I449722);
DFFARX1 I_29633 (I506293,I2507,I506109,I506098,);
nor I_29634 (I506324,I506211,I449731);
nand I_29635 (I506341,I506324,I449719);
nor I_29636 (I506358,I506135,I506341);
DFFARX1 I_29637 (I506358,I2507,I506109,I506074,);
not I_29638 (I506389,I506341);
nand I_29639 (I506086,I506152,I506389);
DFFARX1 I_29640 (I506341,I2507,I506109,I506429,);
not I_29641 (I506437,I506429);
not I_29642 (I506454,I449731);
not I_29643 (I506471,I449728);
nor I_29644 (I506488,I506471,I449737);
nor I_29645 (I506101,I506437,I506488);
nor I_29646 (I506519,I506471,I449734);
and I_29647 (I506536,I506519,I449740);
or I_29648 (I506553,I506536,I449719);
DFFARX1 I_29649 (I506553,I2507,I506109,I506579,);
nor I_29650 (I506089,I506579,I506135);
not I_29651 (I506601,I506579);
and I_29652 (I506618,I506601,I506135);
nor I_29653 (I506083,I506160,I506618);
nand I_29654 (I506649,I506601,I506211);
nor I_29655 (I506077,I506471,I506649);
nand I_29656 (I506080,I506601,I506389);
nand I_29657 (I506694,I506211,I449728);
nor I_29658 (I506092,I506454,I506694);
not I_29659 (I506755,I2514);
DFFARX1 I_29660 (I694808,I2507,I506755,I506781,);
DFFARX1 I_29661 (I694832,I2507,I506755,I506798,);
not I_29662 (I506806,I506798);
not I_29663 (I506823,I694814);
nor I_29664 (I506840,I506823,I694823);
not I_29665 (I506857,I694808);
nor I_29666 (I506874,I506840,I694829);
nor I_29667 (I506891,I506798,I506874);
DFFARX1 I_29668 (I506891,I2507,I506755,I506741,);
nor I_29669 (I506922,I694829,I694823);
nand I_29670 (I506939,I506922,I694814);
DFFARX1 I_29671 (I506939,I2507,I506755,I506744,);
nor I_29672 (I506970,I506857,I694829);
nand I_29673 (I506987,I506970,I694826);
nor I_29674 (I507004,I506781,I506987);
DFFARX1 I_29675 (I507004,I2507,I506755,I506720,);
not I_29676 (I507035,I506987);
nand I_29677 (I506732,I506798,I507035);
DFFARX1 I_29678 (I506987,I2507,I506755,I507075,);
not I_29679 (I507083,I507075);
not I_29680 (I507100,I694829);
not I_29681 (I507117,I694820);
nor I_29682 (I507134,I507117,I694808);
nor I_29683 (I506747,I507083,I507134);
nor I_29684 (I507165,I507117,I694811);
and I_29685 (I507182,I507165,I694835);
or I_29686 (I507199,I507182,I694817);
DFFARX1 I_29687 (I507199,I2507,I506755,I507225,);
nor I_29688 (I506735,I507225,I506781);
not I_29689 (I507247,I507225);
and I_29690 (I507264,I507247,I506781);
nor I_29691 (I506729,I506806,I507264);
nand I_29692 (I507295,I507247,I506857);
nor I_29693 (I506723,I507117,I507295);
nand I_29694 (I506726,I507247,I507035);
nand I_29695 (I507340,I506857,I694820);
nor I_29696 (I506738,I507100,I507340);
not I_29697 (I507401,I2514);
DFFARX1 I_29698 (I212229,I2507,I507401,I507427,);
DFFARX1 I_29699 (I212235,I2507,I507401,I507444,);
not I_29700 (I507452,I507444);
not I_29701 (I507469,I212256);
nor I_29702 (I507486,I507469,I212244);
not I_29703 (I507503,I212253);
nor I_29704 (I507520,I507486,I212238);
nor I_29705 (I507537,I507444,I507520);
DFFARX1 I_29706 (I507537,I2507,I507401,I507387,);
nor I_29707 (I507568,I212238,I212244);
nand I_29708 (I507585,I507568,I212256);
DFFARX1 I_29709 (I507585,I2507,I507401,I507390,);
nor I_29710 (I507616,I507503,I212238);
nand I_29711 (I507633,I507616,I212229);
nor I_29712 (I507650,I507427,I507633);
DFFARX1 I_29713 (I507650,I2507,I507401,I507366,);
not I_29714 (I507681,I507633);
nand I_29715 (I507378,I507444,I507681);
DFFARX1 I_29716 (I507633,I2507,I507401,I507721,);
not I_29717 (I507729,I507721);
not I_29718 (I507746,I212238);
not I_29719 (I507763,I212241);
nor I_29720 (I507780,I507763,I212253);
nor I_29721 (I507393,I507729,I507780);
nor I_29722 (I507811,I507763,I212250);
and I_29723 (I507828,I507811,I212232);
or I_29724 (I507845,I507828,I212247);
DFFARX1 I_29725 (I507845,I2507,I507401,I507871,);
nor I_29726 (I507381,I507871,I507427);
not I_29727 (I507893,I507871);
and I_29728 (I507910,I507893,I507427);
nor I_29729 (I507375,I507452,I507910);
nand I_29730 (I507941,I507893,I507503);
nor I_29731 (I507369,I507763,I507941);
nand I_29732 (I507372,I507893,I507681);
nand I_29733 (I507986,I507503,I212241);
nor I_29734 (I507384,I507746,I507986);
not I_29735 (I508047,I2514);
DFFARX1 I_29736 (I571695,I2507,I508047,I508073,);
DFFARX1 I_29737 (I571677,I2507,I508047,I508090,);
not I_29738 (I508098,I508090);
not I_29739 (I508115,I571686);
nor I_29740 (I508132,I508115,I571698);
not I_29741 (I508149,I571680);
nor I_29742 (I508166,I508132,I571689);
nor I_29743 (I508183,I508090,I508166);
DFFARX1 I_29744 (I508183,I2507,I508047,I508033,);
nor I_29745 (I508214,I571689,I571698);
nand I_29746 (I508231,I508214,I571686);
DFFARX1 I_29747 (I508231,I2507,I508047,I508036,);
nor I_29748 (I508262,I508149,I571689);
nand I_29749 (I508279,I508262,I571701);
nor I_29750 (I508296,I508073,I508279);
DFFARX1 I_29751 (I508296,I2507,I508047,I508012,);
not I_29752 (I508327,I508279);
nand I_29753 (I508024,I508090,I508327);
DFFARX1 I_29754 (I508279,I2507,I508047,I508367,);
not I_29755 (I508375,I508367);
not I_29756 (I508392,I571689);
not I_29757 (I508409,I571677);
nor I_29758 (I508426,I508409,I571680);
nor I_29759 (I508039,I508375,I508426);
nor I_29760 (I508457,I508409,I571683);
and I_29761 (I508474,I508457,I571692);
or I_29762 (I508491,I508474,I571680);
DFFARX1 I_29763 (I508491,I2507,I508047,I508517,);
nor I_29764 (I508027,I508517,I508073);
not I_29765 (I508539,I508517);
and I_29766 (I508556,I508539,I508073);
nor I_29767 (I508021,I508098,I508556);
nand I_29768 (I508587,I508539,I508149);
nor I_29769 (I508015,I508409,I508587);
nand I_29770 (I508018,I508539,I508327);
nand I_29771 (I508632,I508149,I571677);
nor I_29772 (I508030,I508392,I508632);
not I_29773 (I508693,I2514);
DFFARX1 I_29774 (I151460,I2507,I508693,I508719,);
DFFARX1 I_29775 (I151472,I2507,I508693,I508736,);
not I_29776 (I508744,I508736);
not I_29777 (I508761,I151478);
nor I_29778 (I508778,I508761,I151463);
not I_29779 (I508795,I151454);
nor I_29780 (I508812,I508778,I151475);
nor I_29781 (I508829,I508736,I508812);
DFFARX1 I_29782 (I508829,I2507,I508693,I508679,);
nor I_29783 (I508860,I151475,I151463);
nand I_29784 (I508877,I508860,I151478);
DFFARX1 I_29785 (I508877,I2507,I508693,I508682,);
nor I_29786 (I508908,I508795,I151475);
nand I_29787 (I508925,I508908,I151457);
nor I_29788 (I508942,I508719,I508925);
DFFARX1 I_29789 (I508942,I2507,I508693,I508658,);
not I_29790 (I508973,I508925);
nand I_29791 (I508670,I508736,I508973);
DFFARX1 I_29792 (I508925,I2507,I508693,I509013,);
not I_29793 (I509021,I509013);
not I_29794 (I509038,I151475);
not I_29795 (I509055,I151466);
nor I_29796 (I509072,I509055,I151454);
nor I_29797 (I508685,I509021,I509072);
nor I_29798 (I509103,I509055,I151469);
and I_29799 (I509120,I509103,I151457);
or I_29800 (I509137,I509120,I151454);
DFFARX1 I_29801 (I509137,I2507,I508693,I509163,);
nor I_29802 (I508673,I509163,I508719);
not I_29803 (I509185,I509163);
and I_29804 (I509202,I509185,I508719);
nor I_29805 (I508667,I508744,I509202);
nand I_29806 (I509233,I509185,I508795);
nor I_29807 (I508661,I509055,I509233);
nand I_29808 (I508664,I509185,I508973);
nand I_29809 (I509278,I508795,I151466);
nor I_29810 (I508676,I509038,I509278);
not I_29811 (I509339,I2514);
DFFARX1 I_29812 (I571117,I2507,I509339,I509365,);
DFFARX1 I_29813 (I571099,I2507,I509339,I509382,);
not I_29814 (I509390,I509382);
not I_29815 (I509407,I571108);
nor I_29816 (I509424,I509407,I571120);
not I_29817 (I509441,I571102);
nor I_29818 (I509458,I509424,I571111);
nor I_29819 (I509475,I509382,I509458);
DFFARX1 I_29820 (I509475,I2507,I509339,I509325,);
nor I_29821 (I509506,I571111,I571120);
nand I_29822 (I509523,I509506,I571108);
DFFARX1 I_29823 (I509523,I2507,I509339,I509328,);
nor I_29824 (I509554,I509441,I571111);
nand I_29825 (I509571,I509554,I571123);
nor I_29826 (I509588,I509365,I509571);
DFFARX1 I_29827 (I509588,I2507,I509339,I509304,);
not I_29828 (I509619,I509571);
nand I_29829 (I509316,I509382,I509619);
DFFARX1 I_29830 (I509571,I2507,I509339,I509659,);
not I_29831 (I509667,I509659);
not I_29832 (I509684,I571111);
not I_29833 (I509701,I571099);
nor I_29834 (I509718,I509701,I571102);
nor I_29835 (I509331,I509667,I509718);
nor I_29836 (I509749,I509701,I571105);
and I_29837 (I509766,I509749,I571114);
or I_29838 (I509783,I509766,I571102);
DFFARX1 I_29839 (I509783,I2507,I509339,I509809,);
nor I_29840 (I509319,I509809,I509365);
not I_29841 (I509831,I509809);
and I_29842 (I509848,I509831,I509365);
nor I_29843 (I509313,I509390,I509848);
nand I_29844 (I509879,I509831,I509441);
nor I_29845 (I509307,I509701,I509879);
nand I_29846 (I509310,I509831,I509619);
nand I_29847 (I509924,I509441,I571099);
nor I_29848 (I509322,I509684,I509924);
not I_29849 (I509985,I2514);
DFFARX1 I_29850 (I715633,I2507,I509985,I510011,);
DFFARX1 I_29851 (I715657,I2507,I509985,I510028,);
not I_29852 (I510036,I510028);
not I_29853 (I510053,I715639);
nor I_29854 (I510070,I510053,I715648);
not I_29855 (I510087,I715633);
nor I_29856 (I510104,I510070,I715654);
nor I_29857 (I510121,I510028,I510104);
DFFARX1 I_29858 (I510121,I2507,I509985,I509971,);
nor I_29859 (I510152,I715654,I715648);
nand I_29860 (I510169,I510152,I715639);
DFFARX1 I_29861 (I510169,I2507,I509985,I509974,);
nor I_29862 (I510200,I510087,I715654);
nand I_29863 (I510217,I510200,I715651);
nor I_29864 (I510234,I510011,I510217);
DFFARX1 I_29865 (I510234,I2507,I509985,I509950,);
not I_29866 (I510265,I510217);
nand I_29867 (I509962,I510028,I510265);
DFFARX1 I_29868 (I510217,I2507,I509985,I510305,);
not I_29869 (I510313,I510305);
not I_29870 (I510330,I715654);
not I_29871 (I510347,I715645);
nor I_29872 (I510364,I510347,I715633);
nor I_29873 (I509977,I510313,I510364);
nor I_29874 (I510395,I510347,I715636);
and I_29875 (I510412,I510395,I715660);
or I_29876 (I510429,I510412,I715642);
DFFARX1 I_29877 (I510429,I2507,I509985,I510455,);
nor I_29878 (I509965,I510455,I510011);
not I_29879 (I510477,I510455);
and I_29880 (I510494,I510477,I510011);
nor I_29881 (I509959,I510036,I510494);
nand I_29882 (I510525,I510477,I510087);
nor I_29883 (I509953,I510347,I510525);
nand I_29884 (I509956,I510477,I510265);
nand I_29885 (I510570,I510087,I715645);
nor I_29886 (I509968,I510330,I510570);
not I_29887 (I510631,I2514);
DFFARX1 I_29888 (I310254,I2507,I510631,I510657,);
DFFARX1 I_29889 (I310266,I2507,I510631,I510674,);
not I_29890 (I510682,I510674);
not I_29891 (I510699,I310275);
nor I_29892 (I510716,I510699,I310251);
not I_29893 (I510733,I310269);
nor I_29894 (I510750,I510716,I310263);
nor I_29895 (I510767,I510674,I510750);
DFFARX1 I_29896 (I510767,I2507,I510631,I510617,);
nor I_29897 (I510798,I310263,I310251);
nand I_29898 (I510815,I510798,I310275);
DFFARX1 I_29899 (I510815,I2507,I510631,I510620,);
nor I_29900 (I510846,I510733,I310263);
nand I_29901 (I510863,I510846,I310257);
nor I_29902 (I510880,I510657,I510863);
DFFARX1 I_29903 (I510880,I2507,I510631,I510596,);
not I_29904 (I510911,I510863);
nand I_29905 (I510608,I510674,I510911);
DFFARX1 I_29906 (I510863,I2507,I510631,I510951,);
not I_29907 (I510959,I510951);
not I_29908 (I510976,I310263);
not I_29909 (I510993,I310272);
nor I_29910 (I511010,I510993,I310269);
nor I_29911 (I510623,I510959,I511010);
nor I_29912 (I511041,I510993,I310254);
and I_29913 (I511058,I511041,I310251);
or I_29914 (I511075,I511058,I310260);
DFFARX1 I_29915 (I511075,I2507,I510631,I511101,);
nor I_29916 (I510611,I511101,I510657);
not I_29917 (I511123,I511101);
and I_29918 (I511140,I511123,I510657);
nor I_29919 (I510605,I510682,I511140);
nand I_29920 (I511171,I511123,I510733);
nor I_29921 (I510599,I510993,I511171);
nand I_29922 (I510602,I511123,I510911);
nand I_29923 (I511216,I510733,I310272);
nor I_29924 (I510614,I510976,I511216);
not I_29925 (I511277,I2514);
DFFARX1 I_29926 (I416031,I2507,I511277,I511303,);
DFFARX1 I_29927 (I416025,I2507,I511277,I511320,);
not I_29928 (I511328,I511320);
not I_29929 (I511345,I416040);
nor I_29930 (I511362,I511345,I416025);
not I_29931 (I511379,I416034);
nor I_29932 (I511396,I511362,I416043);
nor I_29933 (I511413,I511320,I511396);
DFFARX1 I_29934 (I511413,I2507,I511277,I511263,);
nor I_29935 (I511444,I416043,I416025);
nand I_29936 (I511461,I511444,I416040);
DFFARX1 I_29937 (I511461,I2507,I511277,I511266,);
nor I_29938 (I511492,I511379,I416043);
nand I_29939 (I511509,I511492,I416028);
nor I_29940 (I511526,I511303,I511509);
DFFARX1 I_29941 (I511526,I2507,I511277,I511242,);
not I_29942 (I511557,I511509);
nand I_29943 (I511254,I511320,I511557);
DFFARX1 I_29944 (I511509,I2507,I511277,I511597,);
not I_29945 (I511605,I511597);
not I_29946 (I511622,I416043);
not I_29947 (I511639,I416037);
nor I_29948 (I511656,I511639,I416034);
nor I_29949 (I511269,I511605,I511656);
nor I_29950 (I511687,I511639,I416046);
and I_29951 (I511704,I511687,I416049);
or I_29952 (I511721,I511704,I416028);
DFFARX1 I_29953 (I511721,I2507,I511277,I511747,);
nor I_29954 (I511257,I511747,I511303);
not I_29955 (I511769,I511747);
and I_29956 (I511786,I511769,I511303);
nor I_29957 (I511251,I511328,I511786);
nand I_29958 (I511817,I511769,I511379);
nor I_29959 (I511245,I511639,I511817);
nand I_29960 (I511248,I511769,I511557);
nand I_29961 (I511862,I511379,I416037);
nor I_29962 (I511260,I511622,I511862);
not I_29963 (I511923,I2514);
DFFARX1 I_29964 (I72557,I2507,I511923,I511949,);
DFFARX1 I_29965 (I72563,I2507,I511923,I511966,);
not I_29966 (I511974,I511966);
not I_29967 (I511991,I72581);
nor I_29968 (I512008,I511991,I72560);
not I_29969 (I512025,I72566);
nor I_29970 (I512042,I512008,I72572);
nor I_29971 (I512059,I511966,I512042);
DFFARX1 I_29972 (I512059,I2507,I511923,I511909,);
nor I_29973 (I512090,I72572,I72560);
nand I_29974 (I512107,I512090,I72581);
DFFARX1 I_29975 (I512107,I2507,I511923,I511912,);
nor I_29976 (I512138,I512025,I72572);
nand I_29977 (I512155,I512138,I72578);
nor I_29978 (I512172,I511949,I512155);
DFFARX1 I_29979 (I512172,I2507,I511923,I511888,);
not I_29980 (I512203,I512155);
nand I_29981 (I511900,I511966,I512203);
DFFARX1 I_29982 (I512155,I2507,I511923,I512243,);
not I_29983 (I512251,I512243);
not I_29984 (I512268,I72572);
not I_29985 (I512285,I72560);
nor I_29986 (I512302,I512285,I72566);
nor I_29987 (I511915,I512251,I512302);
nor I_29988 (I512333,I512285,I72569);
and I_29989 (I512350,I512333,I72557);
or I_29990 (I512367,I512350,I72575);
DFFARX1 I_29991 (I512367,I2507,I511923,I512393,);
nor I_29992 (I511903,I512393,I511949);
not I_29993 (I512415,I512393);
and I_29994 (I512432,I512415,I511949);
nor I_29995 (I511897,I511974,I512432);
nand I_29996 (I512463,I512415,I512025);
nor I_29997 (I511891,I512285,I512463);
nand I_29998 (I511894,I512415,I512203);
nand I_29999 (I512508,I512025,I72560);
nor I_30000 (I511906,I512268,I512508);
not I_30001 (I512569,I2514);
DFFARX1 I_30002 (I292081,I2507,I512569,I512595,);
DFFARX1 I_30003 (I292093,I2507,I512569,I512612,);
not I_30004 (I512620,I512612);
not I_30005 (I512637,I292078);
nor I_30006 (I512654,I512637,I292096);
not I_30007 (I512671,I292102);
nor I_30008 (I512688,I512654,I292084);
nor I_30009 (I512705,I512612,I512688);
DFFARX1 I_30010 (I512705,I2507,I512569,I512555,);
nor I_30011 (I512736,I292084,I292096);
nand I_30012 (I512753,I512736,I292078);
DFFARX1 I_30013 (I512753,I2507,I512569,I512558,);
nor I_30014 (I512784,I512671,I292084);
nand I_30015 (I512801,I512784,I292087);
nor I_30016 (I512818,I512595,I512801);
DFFARX1 I_30017 (I512818,I2507,I512569,I512534,);
not I_30018 (I512849,I512801);
nand I_30019 (I512546,I512612,I512849);
DFFARX1 I_30020 (I512801,I2507,I512569,I512889,);
not I_30021 (I512897,I512889);
not I_30022 (I512914,I292084);
not I_30023 (I512931,I292090);
nor I_30024 (I512948,I512931,I292102);
nor I_30025 (I512561,I512897,I512948);
nor I_30026 (I512979,I512931,I292099);
and I_30027 (I512996,I512979,I292078);
or I_30028 (I513013,I512996,I292081);
DFFARX1 I_30029 (I513013,I2507,I512569,I513039,);
nor I_30030 (I512549,I513039,I512595);
not I_30031 (I513061,I513039);
and I_30032 (I513078,I513061,I512595);
nor I_30033 (I512543,I512620,I513078);
nand I_30034 (I513109,I513061,I512671);
nor I_30035 (I512537,I512931,I513109);
nand I_30036 (I512540,I513061,I512849);
nand I_30037 (I513154,I512671,I292090);
nor I_30038 (I512552,I512914,I513154);
not I_30039 (I513215,I2514);
DFFARX1 I_30040 (I443928,I2507,I513215,I513241,);
DFFARX1 I_30041 (I443925,I2507,I513215,I513258,);
not I_30042 (I513266,I513258);
not I_30043 (I513283,I443925);
nor I_30044 (I513300,I513283,I443928);
not I_30045 (I513317,I443940);
nor I_30046 (I513334,I513300,I443934);
nor I_30047 (I513351,I513258,I513334);
DFFARX1 I_30048 (I513351,I2507,I513215,I513201,);
nor I_30049 (I513382,I443934,I443928);
nand I_30050 (I513399,I513382,I443925);
DFFARX1 I_30051 (I513399,I2507,I513215,I513204,);
nor I_30052 (I513430,I513317,I443934);
nand I_30053 (I513447,I513430,I443922);
nor I_30054 (I513464,I513241,I513447);
DFFARX1 I_30055 (I513464,I2507,I513215,I513180,);
not I_30056 (I513495,I513447);
nand I_30057 (I513192,I513258,I513495);
DFFARX1 I_30058 (I513447,I2507,I513215,I513535,);
not I_30059 (I513543,I513535);
not I_30060 (I513560,I443934);
not I_30061 (I513577,I443931);
nor I_30062 (I513594,I513577,I443940);
nor I_30063 (I513207,I513543,I513594);
nor I_30064 (I513625,I513577,I443937);
and I_30065 (I513642,I513625,I443943);
or I_30066 (I513659,I513642,I443922);
DFFARX1 I_30067 (I513659,I2507,I513215,I513685,);
nor I_30068 (I513195,I513685,I513241);
not I_30069 (I513707,I513685);
and I_30070 (I513724,I513707,I513241);
nor I_30071 (I513189,I513266,I513724);
nand I_30072 (I513755,I513707,I513317);
nor I_30073 (I513183,I513577,I513755);
nand I_30074 (I513186,I513707,I513495);
nand I_30075 (I513800,I513317,I443931);
nor I_30076 (I513198,I513560,I513800);
not I_30077 (I513861,I2514);
DFFARX1 I_30078 (I414297,I2507,I513861,I513887,);
DFFARX1 I_30079 (I414291,I2507,I513861,I513904,);
not I_30080 (I513912,I513904);
not I_30081 (I513929,I414306);
nor I_30082 (I513946,I513929,I414291);
not I_30083 (I513963,I414300);
nor I_30084 (I513980,I513946,I414309);
nor I_30085 (I513997,I513904,I513980);
DFFARX1 I_30086 (I513997,I2507,I513861,I513847,);
nor I_30087 (I514028,I414309,I414291);
nand I_30088 (I514045,I514028,I414306);
DFFARX1 I_30089 (I514045,I2507,I513861,I513850,);
nor I_30090 (I514076,I513963,I414309);
nand I_30091 (I514093,I514076,I414294);
nor I_30092 (I514110,I513887,I514093);
DFFARX1 I_30093 (I514110,I2507,I513861,I513826,);
not I_30094 (I514141,I514093);
nand I_30095 (I513838,I513904,I514141);
DFFARX1 I_30096 (I514093,I2507,I513861,I514181,);
not I_30097 (I514189,I514181);
not I_30098 (I514206,I414309);
not I_30099 (I514223,I414303);
nor I_30100 (I514240,I514223,I414300);
nor I_30101 (I513853,I514189,I514240);
nor I_30102 (I514271,I514223,I414312);
and I_30103 (I514288,I514271,I414315);
or I_30104 (I514305,I514288,I414294);
DFFARX1 I_30105 (I514305,I2507,I513861,I514331,);
nor I_30106 (I513841,I514331,I513887);
not I_30107 (I514353,I514331);
and I_30108 (I514370,I514353,I513887);
nor I_30109 (I513835,I513912,I514370);
nand I_30110 (I514401,I514353,I513963);
nor I_30111 (I513829,I514223,I514401);
nand I_30112 (I513832,I514353,I514141);
nand I_30113 (I514446,I513963,I414303);
nor I_30114 (I513844,I514206,I514446);
not I_30115 (I514507,I2514);
DFFARX1 I_30116 (I83642,I2507,I514507,I514533,);
DFFARX1 I_30117 (I83645,I2507,I514507,I514550,);
not I_30118 (I514558,I514550);
not I_30119 (I514575,I83630);
nor I_30120 (I514592,I514575,I83624);
not I_30121 (I514609,I83633);
nor I_30122 (I514626,I514592,I83648);
nor I_30123 (I514643,I514550,I514626);
DFFARX1 I_30124 (I514643,I2507,I514507,I514493,);
nor I_30125 (I514674,I83648,I83624);
nand I_30126 (I514691,I514674,I83630);
DFFARX1 I_30127 (I514691,I2507,I514507,I514496,);
nor I_30128 (I514722,I514609,I83648);
nand I_30129 (I514739,I514722,I83651);
nor I_30130 (I514756,I514533,I514739);
DFFARX1 I_30131 (I514756,I2507,I514507,I514472,);
not I_30132 (I514787,I514739);
nand I_30133 (I514484,I514550,I514787);
DFFARX1 I_30134 (I514739,I2507,I514507,I514827,);
not I_30135 (I514835,I514827);
not I_30136 (I514852,I83648);
not I_30137 (I514869,I83627);
nor I_30138 (I514886,I514869,I83633);
nor I_30139 (I514499,I514835,I514886);
nor I_30140 (I514917,I514869,I83636);
and I_30141 (I514934,I514917,I83624);
or I_30142 (I514951,I514934,I83639);
DFFARX1 I_30143 (I514951,I2507,I514507,I514977,);
nor I_30144 (I514487,I514977,I514533);
not I_30145 (I514999,I514977);
and I_30146 (I515016,I514999,I514533);
nor I_30147 (I514481,I514558,I515016);
nand I_30148 (I515047,I514999,I514609);
nor I_30149 (I514475,I514869,I515047);
nand I_30150 (I514478,I514999,I514787);
nand I_30151 (I515092,I514609,I83627);
nor I_30152 (I514490,I514852,I515092);
not I_30153 (I515153,I2514);
DFFARX1 I_30154 (I691238,I2507,I515153,I515179,);
DFFARX1 I_30155 (I691262,I2507,I515153,I515196,);
not I_30156 (I515204,I515196);
not I_30157 (I515221,I691244);
nor I_30158 (I515238,I515221,I691253);
not I_30159 (I515255,I691238);
nor I_30160 (I515272,I515238,I691259);
nor I_30161 (I515289,I515196,I515272);
DFFARX1 I_30162 (I515289,I2507,I515153,I515139,);
nor I_30163 (I515320,I691259,I691253);
nand I_30164 (I515337,I515320,I691244);
DFFARX1 I_30165 (I515337,I2507,I515153,I515142,);
nor I_30166 (I515368,I515255,I691259);
nand I_30167 (I515385,I515368,I691256);
nor I_30168 (I515402,I515179,I515385);
DFFARX1 I_30169 (I515402,I2507,I515153,I515118,);
not I_30170 (I515433,I515385);
nand I_30171 (I515130,I515196,I515433);
DFFARX1 I_30172 (I515385,I2507,I515153,I515473,);
not I_30173 (I515481,I515473);
not I_30174 (I515498,I691259);
not I_30175 (I515515,I691250);
nor I_30176 (I515532,I515515,I691238);
nor I_30177 (I515145,I515481,I515532);
nor I_30178 (I515563,I515515,I691241);
and I_30179 (I515580,I515563,I691265);
or I_30180 (I515597,I515580,I691247);
DFFARX1 I_30181 (I515597,I2507,I515153,I515623,);
nor I_30182 (I515133,I515623,I515179);
not I_30183 (I515645,I515623);
and I_30184 (I515662,I515645,I515179);
nor I_30185 (I515127,I515204,I515662);
nand I_30186 (I515693,I515645,I515255);
nor I_30187 (I515121,I515515,I515693);
nand I_30188 (I515124,I515645,I515433);
nand I_30189 (I515738,I515255,I691250);
nor I_30190 (I515136,I515498,I515738);
not I_30191 (I515799,I2514);
DFFARX1 I_30192 (I268862,I2507,I515799,I515825,);
DFFARX1 I_30193 (I268859,I2507,I515799,I515842,);
not I_30194 (I515850,I515842);
not I_30195 (I515867,I268874);
nor I_30196 (I515884,I515867,I268877);
not I_30197 (I515901,I268865);
nor I_30198 (I515918,I515884,I268871);
nor I_30199 (I515935,I515842,I515918);
DFFARX1 I_30200 (I515935,I2507,I515799,I515785,);
nor I_30201 (I515966,I268871,I268877);
nand I_30202 (I515983,I515966,I268874);
DFFARX1 I_30203 (I515983,I2507,I515799,I515788,);
nor I_30204 (I516014,I515901,I268871);
nand I_30205 (I516031,I516014,I268883);
nor I_30206 (I516048,I515825,I516031);
DFFARX1 I_30207 (I516048,I2507,I515799,I515764,);
not I_30208 (I516079,I516031);
nand I_30209 (I515776,I515842,I516079);
DFFARX1 I_30210 (I516031,I2507,I515799,I516119,);
not I_30211 (I516127,I516119);
not I_30212 (I516144,I268871);
not I_30213 (I516161,I268856);
nor I_30214 (I516178,I516161,I268865);
nor I_30215 (I515791,I516127,I516178);
nor I_30216 (I516209,I516161,I268868);
and I_30217 (I516226,I516209,I268856);
or I_30218 (I516243,I516226,I268880);
DFFARX1 I_30219 (I516243,I2507,I515799,I516269,);
nor I_30220 (I515779,I516269,I515825);
not I_30221 (I516291,I516269);
and I_30222 (I516308,I516291,I515825);
nor I_30223 (I515773,I515850,I516308);
nand I_30224 (I516339,I516291,I515901);
nor I_30225 (I515767,I516161,I516339);
nand I_30226 (I515770,I516291,I516079);
nand I_30227 (I516384,I515901,I268856);
nor I_30228 (I515782,I516144,I516384);
not I_30229 (I516445,I2514);
DFFARX1 I_30230 (I16695,I2507,I516445,I516471,);
DFFARX1 I_30231 (I16701,I2507,I516445,I516488,);
not I_30232 (I516496,I516488);
not I_30233 (I516513,I16695);
nor I_30234 (I516530,I516513,I16707);
not I_30235 (I516547,I16719);
nor I_30236 (I516564,I516530,I16713);
nor I_30237 (I516581,I516488,I516564);
DFFARX1 I_30238 (I516581,I2507,I516445,I516431,);
nor I_30239 (I516612,I16713,I16707);
nand I_30240 (I516629,I516612,I16695);
DFFARX1 I_30241 (I516629,I2507,I516445,I516434,);
nor I_30242 (I516660,I516547,I16713);
nand I_30243 (I516677,I516660,I16698);
nor I_30244 (I516694,I516471,I516677);
DFFARX1 I_30245 (I516694,I2507,I516445,I516410,);
not I_30246 (I516725,I516677);
nand I_30247 (I516422,I516488,I516725);
DFFARX1 I_30248 (I516677,I2507,I516445,I516765,);
not I_30249 (I516773,I516765);
not I_30250 (I516790,I16713);
not I_30251 (I516807,I16698);
nor I_30252 (I516824,I516807,I16719);
nor I_30253 (I516437,I516773,I516824);
nor I_30254 (I516855,I516807,I16716);
and I_30255 (I516872,I516855,I16710);
or I_30256 (I516889,I516872,I16704);
DFFARX1 I_30257 (I516889,I2507,I516445,I516915,);
nor I_30258 (I516425,I516915,I516471);
not I_30259 (I516937,I516915);
and I_30260 (I516954,I516937,I516471);
nor I_30261 (I516419,I516496,I516954);
nand I_30262 (I516985,I516937,I516547);
nor I_30263 (I516413,I516807,I516985);
nand I_30264 (I516416,I516937,I516725);
nand I_30265 (I517030,I516547,I16698);
nor I_30266 (I516428,I516790,I517030);
not I_30267 (I517091,I2514);
DFFARX1 I_30268 (I395801,I2507,I517091,I517117,);
DFFARX1 I_30269 (I395795,I2507,I517091,I517134,);
not I_30270 (I517142,I517134);
not I_30271 (I517159,I395810);
nor I_30272 (I517176,I517159,I395795);
not I_30273 (I517193,I395804);
nor I_30274 (I517210,I517176,I395813);
nor I_30275 (I517227,I517134,I517210);
DFFARX1 I_30276 (I517227,I2507,I517091,I517077,);
nor I_30277 (I517258,I395813,I395795);
nand I_30278 (I517275,I517258,I395810);
DFFARX1 I_30279 (I517275,I2507,I517091,I517080,);
nor I_30280 (I517306,I517193,I395813);
nand I_30281 (I517323,I517306,I395798);
nor I_30282 (I517340,I517117,I517323);
DFFARX1 I_30283 (I517340,I2507,I517091,I517056,);
not I_30284 (I517371,I517323);
nand I_30285 (I517068,I517134,I517371);
DFFARX1 I_30286 (I517323,I2507,I517091,I517411,);
not I_30287 (I517419,I517411);
not I_30288 (I517436,I395813);
not I_30289 (I517453,I395807);
nor I_30290 (I517470,I517453,I395804);
nor I_30291 (I517083,I517419,I517470);
nor I_30292 (I517501,I517453,I395816);
and I_30293 (I517518,I517501,I395819);
or I_30294 (I517535,I517518,I395798);
DFFARX1 I_30295 (I517535,I2507,I517091,I517561,);
nor I_30296 (I517071,I517561,I517117);
not I_30297 (I517583,I517561);
and I_30298 (I517600,I517583,I517117);
nor I_30299 (I517065,I517142,I517600);
nand I_30300 (I517631,I517583,I517193);
nor I_30301 (I517059,I517453,I517631);
nand I_30302 (I517062,I517583,I517371);
nand I_30303 (I517676,I517193,I395807);
nor I_30304 (I517074,I517436,I517676);
not I_30305 (I517737,I2514);
DFFARX1 I_30306 (I256350,I2507,I517737,I517763,);
DFFARX1 I_30307 (I256347,I2507,I517737,I517780,);
not I_30308 (I517788,I517780);
not I_30309 (I517805,I256362);
nor I_30310 (I517822,I517805,I256365);
not I_30311 (I517839,I256353);
nor I_30312 (I517856,I517822,I256359);
nor I_30313 (I517873,I517780,I517856);
DFFARX1 I_30314 (I517873,I2507,I517737,I517723,);
nor I_30315 (I517904,I256359,I256365);
nand I_30316 (I517921,I517904,I256362);
DFFARX1 I_30317 (I517921,I2507,I517737,I517726,);
nor I_30318 (I517952,I517839,I256359);
nand I_30319 (I517969,I517952,I256371);
nor I_30320 (I517986,I517763,I517969);
DFFARX1 I_30321 (I517986,I2507,I517737,I517702,);
not I_30322 (I518017,I517969);
nand I_30323 (I517714,I517780,I518017);
DFFARX1 I_30324 (I517969,I2507,I517737,I518057,);
not I_30325 (I518065,I518057);
not I_30326 (I518082,I256359);
not I_30327 (I518099,I256344);
nor I_30328 (I518116,I518099,I256353);
nor I_30329 (I517729,I518065,I518116);
nor I_30330 (I518147,I518099,I256356);
and I_30331 (I518164,I518147,I256344);
or I_30332 (I518181,I518164,I256368);
DFFARX1 I_30333 (I518181,I2507,I517737,I518207,);
nor I_30334 (I517717,I518207,I517763);
not I_30335 (I518229,I518207);
and I_30336 (I518246,I518229,I517763);
nor I_30337 (I517711,I517788,I518246);
nand I_30338 (I518277,I518229,I517839);
nor I_30339 (I517705,I518099,I518277);
nand I_30340 (I517708,I518229,I518017);
nand I_30341 (I518322,I517839,I256344);
nor I_30342 (I517720,I518082,I518322);
not I_30343 (I518383,I2514);
DFFARX1 I_30344 (I475021,I2507,I518383,I518409,);
DFFARX1 I_30345 (I475018,I2507,I518383,I518426,);
not I_30346 (I518434,I518426);
not I_30347 (I518451,I475018);
nor I_30348 (I518468,I518451,I475021);
not I_30349 (I518485,I475033);
nor I_30350 (I518502,I518468,I475027);
nor I_30351 (I518519,I518426,I518502);
DFFARX1 I_30352 (I518519,I2507,I518383,I518369,);
nor I_30353 (I518550,I475027,I475021);
nand I_30354 (I518567,I518550,I475018);
DFFARX1 I_30355 (I518567,I2507,I518383,I518372,);
nor I_30356 (I518598,I518485,I475027);
nand I_30357 (I518615,I518598,I475015);
nor I_30358 (I518632,I518409,I518615);
DFFARX1 I_30359 (I518632,I2507,I518383,I518348,);
not I_30360 (I518663,I518615);
nand I_30361 (I518360,I518426,I518663);
DFFARX1 I_30362 (I518615,I2507,I518383,I518703,);
not I_30363 (I518711,I518703);
not I_30364 (I518728,I475027);
not I_30365 (I518745,I475024);
nor I_30366 (I518762,I518745,I475033);
nor I_30367 (I518375,I518711,I518762);
nor I_30368 (I518793,I518745,I475030);
and I_30369 (I518810,I518793,I475036);
or I_30370 (I518827,I518810,I475015);
DFFARX1 I_30371 (I518827,I2507,I518383,I518853,);
nor I_30372 (I518363,I518853,I518409);
not I_30373 (I518875,I518853);
and I_30374 (I518892,I518875,I518409);
nor I_30375 (I518357,I518434,I518892);
nand I_30376 (I518923,I518875,I518485);
nor I_30377 (I518351,I518745,I518923);
nand I_30378 (I518354,I518875,I518663);
nand I_30379 (I518968,I518485,I475024);
nor I_30380 (I518366,I518728,I518968);
not I_30381 (I519029,I2514);
DFFARX1 I_30382 (I383663,I2507,I519029,I519055,);
DFFARX1 I_30383 (I383657,I2507,I519029,I519072,);
not I_30384 (I519080,I519072);
not I_30385 (I519097,I383672);
nor I_30386 (I519114,I519097,I383657);
not I_30387 (I519131,I383666);
nor I_30388 (I519148,I519114,I383675);
nor I_30389 (I519165,I519072,I519148);
DFFARX1 I_30390 (I519165,I2507,I519029,I519015,);
nor I_30391 (I519196,I383675,I383657);
nand I_30392 (I519213,I519196,I383672);
DFFARX1 I_30393 (I519213,I2507,I519029,I519018,);
nor I_30394 (I519244,I519131,I383675);
nand I_30395 (I519261,I519244,I383660);
nor I_30396 (I519278,I519055,I519261);
DFFARX1 I_30397 (I519278,I2507,I519029,I518994,);
not I_30398 (I519309,I519261);
nand I_30399 (I519006,I519072,I519309);
DFFARX1 I_30400 (I519261,I2507,I519029,I519349,);
not I_30401 (I519357,I519349);
not I_30402 (I519374,I383675);
not I_30403 (I519391,I383669);
nor I_30404 (I519408,I519391,I383666);
nor I_30405 (I519021,I519357,I519408);
nor I_30406 (I519439,I519391,I383678);
and I_30407 (I519456,I519439,I383681);
or I_30408 (I519473,I519456,I383660);
DFFARX1 I_30409 (I519473,I2507,I519029,I519499,);
nor I_30410 (I519009,I519499,I519055);
not I_30411 (I519521,I519499);
and I_30412 (I519538,I519521,I519055);
nor I_30413 (I519003,I519080,I519538);
nand I_30414 (I519569,I519521,I519131);
nor I_30415 (I518997,I519391,I519569);
nand I_30416 (I519000,I519521,I519309);
nand I_30417 (I519614,I519131,I383669);
nor I_30418 (I519012,I519374,I519614);
not I_30419 (I519675,I2514);
DFFARX1 I_30420 (I431807,I2507,I519675,I519701,);
DFFARX1 I_30421 (I431804,I2507,I519675,I519718,);
not I_30422 (I519726,I519718);
not I_30423 (I519743,I431804);
nor I_30424 (I519760,I519743,I431807);
not I_30425 (I519777,I431819);
nor I_30426 (I519794,I519760,I431813);
nor I_30427 (I519811,I519718,I519794);
DFFARX1 I_30428 (I519811,I2507,I519675,I519661,);
nor I_30429 (I519842,I431813,I431807);
nand I_30430 (I519859,I519842,I431804);
DFFARX1 I_30431 (I519859,I2507,I519675,I519664,);
nor I_30432 (I519890,I519777,I431813);
nand I_30433 (I519907,I519890,I431801);
nor I_30434 (I519924,I519701,I519907);
DFFARX1 I_30435 (I519924,I2507,I519675,I519640,);
not I_30436 (I519955,I519907);
nand I_30437 (I519652,I519718,I519955);
DFFARX1 I_30438 (I519907,I2507,I519675,I519995,);
not I_30439 (I520003,I519995);
not I_30440 (I520020,I431813);
not I_30441 (I520037,I431810);
nor I_30442 (I520054,I520037,I431819);
nor I_30443 (I519667,I520003,I520054);
nor I_30444 (I520085,I520037,I431816);
and I_30445 (I520102,I520085,I431822);
or I_30446 (I520119,I520102,I431801);
DFFARX1 I_30447 (I520119,I2507,I519675,I520145,);
nor I_30448 (I519655,I520145,I519701);
not I_30449 (I520167,I520145);
and I_30450 (I520184,I520167,I519701);
nor I_30451 (I519649,I519726,I520184);
nand I_30452 (I520215,I520167,I519777);
nor I_30453 (I519643,I520037,I520215);
nand I_30454 (I519646,I520167,I519955);
nand I_30455 (I520260,I519777,I431810);
nor I_30456 (I519658,I520020,I520260);
not I_30457 (I520321,I2514);
DFFARX1 I_30458 (I50950,I2507,I520321,I520347,);
DFFARX1 I_30459 (I50956,I2507,I520321,I520364,);
not I_30460 (I520372,I520364);
not I_30461 (I520389,I50974);
nor I_30462 (I520406,I520389,I50953);
not I_30463 (I520423,I50959);
nor I_30464 (I520440,I520406,I50965);
nor I_30465 (I520457,I520364,I520440);
DFFARX1 I_30466 (I520457,I2507,I520321,I520307,);
nor I_30467 (I520488,I50965,I50953);
nand I_30468 (I520505,I520488,I50974);
DFFARX1 I_30469 (I520505,I2507,I520321,I520310,);
nor I_30470 (I520536,I520423,I50965);
nand I_30471 (I520553,I520536,I50971);
nor I_30472 (I520570,I520347,I520553);
DFFARX1 I_30473 (I520570,I2507,I520321,I520286,);
not I_30474 (I520601,I520553);
nand I_30475 (I520298,I520364,I520601);
DFFARX1 I_30476 (I520553,I2507,I520321,I520641,);
not I_30477 (I520649,I520641);
not I_30478 (I520666,I50965);
not I_30479 (I520683,I50953);
nor I_30480 (I520700,I520683,I50959);
nor I_30481 (I520313,I520649,I520700);
nor I_30482 (I520731,I520683,I50962);
and I_30483 (I520748,I520731,I50950);
or I_30484 (I520765,I520748,I50968);
DFFARX1 I_30485 (I520765,I2507,I520321,I520791,);
nor I_30486 (I520301,I520791,I520347);
not I_30487 (I520813,I520791);
and I_30488 (I520830,I520813,I520347);
nor I_30489 (I520295,I520372,I520830);
nand I_30490 (I520861,I520813,I520423);
nor I_30491 (I520289,I520683,I520861);
nand I_30492 (I520292,I520813,I520601);
nand I_30493 (I520906,I520423,I50953);
nor I_30494 (I520304,I520666,I520906);
not I_30495 (I520967,I2514);
DFFARX1 I_30496 (I228606,I2507,I520967,I520993,);
DFFARX1 I_30497 (I228603,I2507,I520967,I521010,);
not I_30498 (I521018,I521010);
not I_30499 (I521035,I228618);
nor I_30500 (I521052,I521035,I228621);
not I_30501 (I521069,I228609);
nor I_30502 (I521086,I521052,I228615);
nor I_30503 (I521103,I521010,I521086);
DFFARX1 I_30504 (I521103,I2507,I520967,I520953,);
nor I_30505 (I521134,I228615,I228621);
nand I_30506 (I521151,I521134,I228618);
DFFARX1 I_30507 (I521151,I2507,I520967,I520956,);
nor I_30508 (I521182,I521069,I228615);
nand I_30509 (I521199,I521182,I228627);
nor I_30510 (I521216,I520993,I521199);
DFFARX1 I_30511 (I521216,I2507,I520967,I520932,);
not I_30512 (I521247,I521199);
nand I_30513 (I520944,I521010,I521247);
DFFARX1 I_30514 (I521199,I2507,I520967,I521287,);
not I_30515 (I521295,I521287);
not I_30516 (I521312,I228615);
not I_30517 (I521329,I228600);
nor I_30518 (I521346,I521329,I228609);
nor I_30519 (I520959,I521295,I521346);
nor I_30520 (I521377,I521329,I228612);
and I_30521 (I521394,I521377,I228600);
or I_30522 (I521411,I521394,I228624);
DFFARX1 I_30523 (I521411,I2507,I520967,I521437,);
nor I_30524 (I520947,I521437,I520993);
not I_30525 (I521459,I521437);
and I_30526 (I521476,I521459,I520993);
nor I_30527 (I520941,I521018,I521476);
nand I_30528 (I521507,I521459,I521069);
nor I_30529 (I520935,I521329,I521507);
nand I_30530 (I520938,I521459,I521247);
nand I_30531 (I521552,I521069,I228600);
nor I_30532 (I520950,I521312,I521552);
not I_30533 (I521613,I2514);
DFFARX1 I_30534 (I293271,I2507,I521613,I521639,);
DFFARX1 I_30535 (I293283,I2507,I521613,I521656,);
not I_30536 (I521664,I521656);
not I_30537 (I521681,I293268);
nor I_30538 (I521698,I521681,I293286);
not I_30539 (I521715,I293292);
nor I_30540 (I521732,I521698,I293274);
nor I_30541 (I521749,I521656,I521732);
DFFARX1 I_30542 (I521749,I2507,I521613,I521599,);
nor I_30543 (I521780,I293274,I293286);
nand I_30544 (I521797,I521780,I293268);
DFFARX1 I_30545 (I521797,I2507,I521613,I521602,);
nor I_30546 (I521828,I521715,I293274);
nand I_30547 (I521845,I521828,I293277);
nor I_30548 (I521862,I521639,I521845);
DFFARX1 I_30549 (I521862,I2507,I521613,I521578,);
not I_30550 (I521893,I521845);
nand I_30551 (I521590,I521656,I521893);
DFFARX1 I_30552 (I521845,I2507,I521613,I521933,);
not I_30553 (I521941,I521933);
not I_30554 (I521958,I293274);
not I_30555 (I521975,I293280);
nor I_30556 (I521992,I521975,I293292);
nor I_30557 (I521605,I521941,I521992);
nor I_30558 (I522023,I521975,I293289);
and I_30559 (I522040,I522023,I293268);
or I_30560 (I522057,I522040,I293271);
DFFARX1 I_30561 (I522057,I2507,I521613,I522083,);
nor I_30562 (I521593,I522083,I521639);
not I_30563 (I522105,I522083);
and I_30564 (I522122,I522105,I521639);
nor I_30565 (I521587,I521664,I522122);
nand I_30566 (I522153,I522105,I521715);
nor I_30567 (I521581,I521975,I522153);
nand I_30568 (I521584,I522105,I521893);
nand I_30569 (I522198,I521715,I293280);
nor I_30570 (I521596,I521958,I522198);
not I_30571 (I522259,I2514);
DFFARX1 I_30572 (I651799,I2507,I522259,I522285,);
DFFARX1 I_30573 (I651805,I2507,I522259,I522302,);
not I_30574 (I522310,I522302);
not I_30575 (I522327,I651802);
nor I_30576 (I522344,I522327,I651781);
not I_30577 (I522361,I651784);
nor I_30578 (I522378,I522344,I651790);
nor I_30579 (I522395,I522302,I522378);
DFFARX1 I_30580 (I522395,I2507,I522259,I522245,);
nor I_30581 (I522426,I651790,I651781);
nand I_30582 (I522443,I522426,I651802);
DFFARX1 I_30583 (I522443,I2507,I522259,I522248,);
nor I_30584 (I522474,I522361,I651790);
nand I_30585 (I522491,I522474,I651784);
nor I_30586 (I522508,I522285,I522491);
DFFARX1 I_30587 (I522508,I2507,I522259,I522224,);
not I_30588 (I522539,I522491);
nand I_30589 (I522236,I522302,I522539);
DFFARX1 I_30590 (I522491,I2507,I522259,I522579,);
not I_30591 (I522587,I522579);
not I_30592 (I522604,I651790);
not I_30593 (I522621,I651793);
nor I_30594 (I522638,I522621,I651784);
nor I_30595 (I522251,I522587,I522638);
nor I_30596 (I522669,I522621,I651781);
and I_30597 (I522686,I522669,I651787);
or I_30598 (I522703,I522686,I651796);
DFFARX1 I_30599 (I522703,I2507,I522259,I522729,);
nor I_30600 (I522239,I522729,I522285);
not I_30601 (I522751,I522729);
and I_30602 (I522768,I522751,I522285);
nor I_30603 (I522233,I522310,I522768);
nand I_30604 (I522799,I522751,I522361);
nor I_30605 (I522227,I522621,I522799);
nand I_30606 (I522230,I522751,I522539);
nand I_30607 (I522844,I522361,I651793);
nor I_30608 (I522242,I522604,I522844);
not I_30609 (I522905,I2514);
DFFARX1 I_30610 (I313144,I2507,I522905,I522931,);
DFFARX1 I_30611 (I313156,I2507,I522905,I522948,);
not I_30612 (I522956,I522948);
not I_30613 (I522973,I313165);
nor I_30614 (I522990,I522973,I313141);
not I_30615 (I523007,I313159);
nor I_30616 (I523024,I522990,I313153);
nor I_30617 (I523041,I522948,I523024);
DFFARX1 I_30618 (I523041,I2507,I522905,I522891,);
nor I_30619 (I523072,I313153,I313141);
nand I_30620 (I523089,I523072,I313165);
DFFARX1 I_30621 (I523089,I2507,I522905,I522894,);
nor I_30622 (I523120,I523007,I313153);
nand I_30623 (I523137,I523120,I313147);
nor I_30624 (I523154,I522931,I523137);
DFFARX1 I_30625 (I523154,I2507,I522905,I522870,);
not I_30626 (I523185,I523137);
nand I_30627 (I522882,I522948,I523185);
DFFARX1 I_30628 (I523137,I2507,I522905,I523225,);
not I_30629 (I523233,I523225);
not I_30630 (I523250,I313153);
not I_30631 (I523267,I313162);
nor I_30632 (I523284,I523267,I313159);
nor I_30633 (I522897,I523233,I523284);
nor I_30634 (I523315,I523267,I313144);
and I_30635 (I523332,I523315,I313141);
or I_30636 (I523349,I523332,I313150);
DFFARX1 I_30637 (I523349,I2507,I522905,I523375,);
nor I_30638 (I522885,I523375,I522931);
not I_30639 (I523397,I523375);
and I_30640 (I523414,I523397,I522931);
nor I_30641 (I522879,I522956,I523414);
nand I_30642 (I523445,I523397,I523007);
nor I_30643 (I522873,I523267,I523445);
nand I_30644 (I522876,I523397,I523185);
nand I_30645 (I523490,I523007,I313162);
nor I_30646 (I522888,I523250,I523490);
not I_30647 (I523551,I2514);
DFFARX1 I_30648 (I232958,I2507,I523551,I523577,);
DFFARX1 I_30649 (I232955,I2507,I523551,I523594,);
not I_30650 (I523602,I523594);
not I_30651 (I523619,I232970);
nor I_30652 (I523636,I523619,I232973);
not I_30653 (I523653,I232961);
nor I_30654 (I523670,I523636,I232967);
nor I_30655 (I523687,I523594,I523670);
DFFARX1 I_30656 (I523687,I2507,I523551,I523537,);
nor I_30657 (I523718,I232967,I232973);
nand I_30658 (I523735,I523718,I232970);
DFFARX1 I_30659 (I523735,I2507,I523551,I523540,);
nor I_30660 (I523766,I523653,I232967);
nand I_30661 (I523783,I523766,I232979);
nor I_30662 (I523800,I523577,I523783);
DFFARX1 I_30663 (I523800,I2507,I523551,I523516,);
not I_30664 (I523831,I523783);
nand I_30665 (I523528,I523594,I523831);
DFFARX1 I_30666 (I523783,I2507,I523551,I523871,);
not I_30667 (I523879,I523871);
not I_30668 (I523896,I232967);
not I_30669 (I523913,I232952);
nor I_30670 (I523930,I523913,I232961);
nor I_30671 (I523543,I523879,I523930);
nor I_30672 (I523961,I523913,I232964);
and I_30673 (I523978,I523961,I232952);
or I_30674 (I523995,I523978,I232976);
DFFARX1 I_30675 (I523995,I2507,I523551,I524021,);
nor I_30676 (I523531,I524021,I523577);
not I_30677 (I524043,I524021);
and I_30678 (I524060,I524043,I523577);
nor I_30679 (I523525,I523602,I524060);
nand I_30680 (I524091,I524043,I523653);
nor I_30681 (I523519,I523913,I524091);
nand I_30682 (I523522,I524043,I523831);
nand I_30683 (I524136,I523653,I232952);
nor I_30684 (I523534,I523896,I524136);
not I_30685 (I524197,I2514);
DFFARX1 I_30686 (I262334,I2507,I524197,I524223,);
DFFARX1 I_30687 (I262331,I2507,I524197,I524240,);
not I_30688 (I524248,I524240);
not I_30689 (I524265,I262346);
nor I_30690 (I524282,I524265,I262349);
not I_30691 (I524299,I262337);
nor I_30692 (I524316,I524282,I262343);
nor I_30693 (I524333,I524240,I524316);
DFFARX1 I_30694 (I524333,I2507,I524197,I524183,);
nor I_30695 (I524364,I262343,I262349);
nand I_30696 (I524381,I524364,I262346);
DFFARX1 I_30697 (I524381,I2507,I524197,I524186,);
nor I_30698 (I524412,I524299,I262343);
nand I_30699 (I524429,I524412,I262355);
nor I_30700 (I524446,I524223,I524429);
DFFARX1 I_30701 (I524446,I2507,I524197,I524162,);
not I_30702 (I524477,I524429);
nand I_30703 (I524174,I524240,I524477);
DFFARX1 I_30704 (I524429,I2507,I524197,I524517,);
not I_30705 (I524525,I524517);
not I_30706 (I524542,I262343);
not I_30707 (I524559,I262328);
nor I_30708 (I524576,I524559,I262337);
nor I_30709 (I524189,I524525,I524576);
nor I_30710 (I524607,I524559,I262340);
and I_30711 (I524624,I524607,I262328);
or I_30712 (I524641,I524624,I262352);
DFFARX1 I_30713 (I524641,I2507,I524197,I524667,);
nor I_30714 (I524177,I524667,I524223);
not I_30715 (I524689,I524667);
and I_30716 (I524706,I524689,I524223);
nor I_30717 (I524171,I524248,I524706);
nand I_30718 (I524737,I524689,I524299);
nor I_30719 (I524165,I524559,I524737);
nand I_30720 (I524168,I524689,I524477);
nand I_30721 (I524782,I524299,I262328);
nor I_30722 (I524180,I524542,I524782);
not I_30723 (I524843,I2514);
DFFARX1 I_30724 (I379039,I2507,I524843,I524869,);
DFFARX1 I_30725 (I379033,I2507,I524843,I524886,);
not I_30726 (I524894,I524886);
not I_30727 (I524911,I379048);
nor I_30728 (I524928,I524911,I379033);
not I_30729 (I524945,I379042);
nor I_30730 (I524962,I524928,I379051);
nor I_30731 (I524979,I524886,I524962);
DFFARX1 I_30732 (I524979,I2507,I524843,I524829,);
nor I_30733 (I525010,I379051,I379033);
nand I_30734 (I525027,I525010,I379048);
DFFARX1 I_30735 (I525027,I2507,I524843,I524832,);
nor I_30736 (I525058,I524945,I379051);
nand I_30737 (I525075,I525058,I379036);
nor I_30738 (I525092,I524869,I525075);
DFFARX1 I_30739 (I525092,I2507,I524843,I524808,);
not I_30740 (I525123,I525075);
nand I_30741 (I524820,I524886,I525123);
DFFARX1 I_30742 (I525075,I2507,I524843,I525163,);
not I_30743 (I525171,I525163);
not I_30744 (I525188,I379051);
not I_30745 (I525205,I379045);
nor I_30746 (I525222,I525205,I379042);
nor I_30747 (I524835,I525171,I525222);
nor I_30748 (I525253,I525205,I379054);
and I_30749 (I525270,I525253,I379057);
or I_30750 (I525287,I525270,I379036);
DFFARX1 I_30751 (I525287,I2507,I524843,I525313,);
nor I_30752 (I524823,I525313,I524869);
not I_30753 (I525335,I525313);
and I_30754 (I525352,I525335,I524869);
nor I_30755 (I524817,I524894,I525352);
nand I_30756 (I525383,I525335,I524945);
nor I_30757 (I524811,I525205,I525383);
nand I_30758 (I524814,I525335,I525123);
nand I_30759 (I525428,I524945,I379045);
nor I_30760 (I524826,I525188,I525428);
not I_30761 (I525489,I2514);
DFFARX1 I_30762 (I292676,I2507,I525489,I525515,);
DFFARX1 I_30763 (I292688,I2507,I525489,I525532,);
not I_30764 (I525540,I525532);
not I_30765 (I525557,I292673);
nor I_30766 (I525574,I525557,I292691);
not I_30767 (I525591,I292697);
nor I_30768 (I525608,I525574,I292679);
nor I_30769 (I525625,I525532,I525608);
DFFARX1 I_30770 (I525625,I2507,I525489,I525475,);
nor I_30771 (I525656,I292679,I292691);
nand I_30772 (I525673,I525656,I292673);
DFFARX1 I_30773 (I525673,I2507,I525489,I525478,);
nor I_30774 (I525704,I525591,I292679);
nand I_30775 (I525721,I525704,I292682);
nor I_30776 (I525738,I525515,I525721);
DFFARX1 I_30777 (I525738,I2507,I525489,I525454,);
not I_30778 (I525769,I525721);
nand I_30779 (I525466,I525532,I525769);
DFFARX1 I_30780 (I525721,I2507,I525489,I525809,);
not I_30781 (I525817,I525809);
not I_30782 (I525834,I292679);
not I_30783 (I525851,I292685);
nor I_30784 (I525868,I525851,I292697);
nor I_30785 (I525481,I525817,I525868);
nor I_30786 (I525899,I525851,I292694);
and I_30787 (I525916,I525899,I292673);
or I_30788 (I525933,I525916,I292676);
DFFARX1 I_30789 (I525933,I2507,I525489,I525959,);
nor I_30790 (I525469,I525959,I525515);
not I_30791 (I525981,I525959);
and I_30792 (I525998,I525981,I525515);
nor I_30793 (I525463,I525540,I525998);
nand I_30794 (I526029,I525981,I525591);
nor I_30795 (I525457,I525851,I526029);
nand I_30796 (I525460,I525981,I525769);
nand I_30797 (I526074,I525591,I292685);
nor I_30798 (I525472,I525834,I526074);
not I_30799 (I526135,I2514);
DFFARX1 I_30800 (I83097,I2507,I526135,I526161,);
DFFARX1 I_30801 (I83103,I2507,I526135,I526178,);
not I_30802 (I526186,I526178);
not I_30803 (I526203,I83121);
nor I_30804 (I526220,I526203,I83100);
not I_30805 (I526237,I83106);
nor I_30806 (I526254,I526220,I83112);
nor I_30807 (I526271,I526178,I526254);
DFFARX1 I_30808 (I526271,I2507,I526135,I526121,);
nor I_30809 (I526302,I83112,I83100);
nand I_30810 (I526319,I526302,I83121);
DFFARX1 I_30811 (I526319,I2507,I526135,I526124,);
nor I_30812 (I526350,I526237,I83112);
nand I_30813 (I526367,I526350,I83118);
nor I_30814 (I526384,I526161,I526367);
DFFARX1 I_30815 (I526384,I2507,I526135,I526100,);
not I_30816 (I526415,I526367);
nand I_30817 (I526112,I526178,I526415);
DFFARX1 I_30818 (I526367,I2507,I526135,I526455,);
not I_30819 (I526463,I526455);
not I_30820 (I526480,I83112);
not I_30821 (I526497,I83100);
nor I_30822 (I526514,I526497,I83106);
nor I_30823 (I526127,I526463,I526514);
nor I_30824 (I526545,I526497,I83109);
and I_30825 (I526562,I526545,I83097);
or I_30826 (I526579,I526562,I83115);
DFFARX1 I_30827 (I526579,I2507,I526135,I526605,);
nor I_30828 (I526115,I526605,I526161);
not I_30829 (I526627,I526605);
and I_30830 (I526644,I526627,I526161);
nor I_30831 (I526109,I526186,I526644);
nand I_30832 (I526675,I526627,I526237);
nor I_30833 (I526103,I526497,I526675);
nand I_30834 (I526106,I526627,I526415);
nand I_30835 (I526720,I526237,I83100);
nor I_30836 (I526118,I526480,I526720);
not I_30837 (I526781,I2514);
DFFARX1 I_30838 (I370947,I2507,I526781,I526807,);
DFFARX1 I_30839 (I370941,I2507,I526781,I526824,);
not I_30840 (I526832,I526824);
not I_30841 (I526849,I370956);
nor I_30842 (I526866,I526849,I370941);
not I_30843 (I526883,I370950);
nor I_30844 (I526900,I526866,I370959);
nor I_30845 (I526917,I526824,I526900);
DFFARX1 I_30846 (I526917,I2507,I526781,I526767,);
nor I_30847 (I526948,I370959,I370941);
nand I_30848 (I526965,I526948,I370956);
DFFARX1 I_30849 (I526965,I2507,I526781,I526770,);
nor I_30850 (I526996,I526883,I370959);
nand I_30851 (I527013,I526996,I370944);
nor I_30852 (I527030,I526807,I527013);
DFFARX1 I_30853 (I527030,I2507,I526781,I526746,);
not I_30854 (I527061,I527013);
nand I_30855 (I526758,I526824,I527061);
DFFARX1 I_30856 (I527013,I2507,I526781,I527101,);
not I_30857 (I527109,I527101);
not I_30858 (I527126,I370959);
not I_30859 (I527143,I370953);
nor I_30860 (I527160,I527143,I370950);
nor I_30861 (I526773,I527109,I527160);
nor I_30862 (I527191,I527143,I370962);
and I_30863 (I527208,I527191,I370965);
or I_30864 (I527225,I527208,I370944);
DFFARX1 I_30865 (I527225,I2507,I526781,I527251,);
nor I_30866 (I526761,I527251,I526807);
not I_30867 (I527273,I527251);
and I_30868 (I527290,I527273,I526807);
nor I_30869 (I526755,I526832,I527290);
nand I_30870 (I527321,I527273,I526883);
nor I_30871 (I526749,I527143,I527321);
nand I_30872 (I526752,I527273,I527061);
nand I_30873 (I527366,I526883,I370953);
nor I_30874 (I526764,I527126,I527366);
not I_30875 (I527427,I2514);
DFFARX1 I_30876 (I121710,I2507,I527427,I527453,);
DFFARX1 I_30877 (I121722,I2507,I527427,I527470,);
not I_30878 (I527478,I527470);
not I_30879 (I527495,I121728);
nor I_30880 (I527512,I527495,I121713);
not I_30881 (I527529,I121704);
nor I_30882 (I527546,I527512,I121725);
nor I_30883 (I527563,I527470,I527546);
DFFARX1 I_30884 (I527563,I2507,I527427,I527413,);
nor I_30885 (I527594,I121725,I121713);
nand I_30886 (I527611,I527594,I121728);
DFFARX1 I_30887 (I527611,I2507,I527427,I527416,);
nor I_30888 (I527642,I527529,I121725);
nand I_30889 (I527659,I527642,I121707);
nor I_30890 (I527676,I527453,I527659);
DFFARX1 I_30891 (I527676,I2507,I527427,I527392,);
not I_30892 (I527707,I527659);
nand I_30893 (I527404,I527470,I527707);
DFFARX1 I_30894 (I527659,I2507,I527427,I527747,);
not I_30895 (I527755,I527747);
not I_30896 (I527772,I121725);
not I_30897 (I527789,I121716);
nor I_30898 (I527806,I527789,I121704);
nor I_30899 (I527419,I527755,I527806);
nor I_30900 (I527837,I527789,I121719);
and I_30901 (I527854,I527837,I121707);
or I_30902 (I527871,I527854,I121704);
DFFARX1 I_30903 (I527871,I2507,I527427,I527897,);
nor I_30904 (I527407,I527897,I527453);
not I_30905 (I527919,I527897);
and I_30906 (I527936,I527919,I527453);
nor I_30907 (I527401,I527478,I527936);
nand I_30908 (I527967,I527919,I527529);
nor I_30909 (I527395,I527789,I527967);
nand I_30910 (I527398,I527919,I527707);
nand I_30911 (I528012,I527529,I121716);
nor I_30912 (I527410,I527772,I528012);
not I_30913 (I528073,I2514);
DFFARX1 I_30914 (I85427,I2507,I528073,I528099,);
DFFARX1 I_30915 (I85430,I2507,I528073,I528116,);
not I_30916 (I528124,I528116);
not I_30917 (I528141,I85415);
nor I_30918 (I528158,I528141,I85409);
not I_30919 (I528175,I85418);
nor I_30920 (I528192,I528158,I85433);
nor I_30921 (I528209,I528116,I528192);
DFFARX1 I_30922 (I528209,I2507,I528073,I528059,);
nor I_30923 (I528240,I85433,I85409);
nand I_30924 (I528257,I528240,I85415);
DFFARX1 I_30925 (I528257,I2507,I528073,I528062,);
nor I_30926 (I528288,I528175,I85433);
nand I_30927 (I528305,I528288,I85436);
nor I_30928 (I528322,I528099,I528305);
DFFARX1 I_30929 (I528322,I2507,I528073,I528038,);
not I_30930 (I528353,I528305);
nand I_30931 (I528050,I528116,I528353);
DFFARX1 I_30932 (I528305,I2507,I528073,I528393,);
not I_30933 (I528401,I528393);
not I_30934 (I528418,I85433);
not I_30935 (I528435,I85412);
nor I_30936 (I528452,I528435,I85418);
nor I_30937 (I528065,I528401,I528452);
nor I_30938 (I528483,I528435,I85421);
and I_30939 (I528500,I528483,I85409);
or I_30940 (I528517,I528500,I85424);
DFFARX1 I_30941 (I528517,I2507,I528073,I528543,);
nor I_30942 (I528053,I528543,I528099);
not I_30943 (I528565,I528543);
and I_30944 (I528582,I528565,I528099);
nor I_30945 (I528047,I528124,I528582);
nand I_30946 (I528613,I528565,I528175);
nor I_30947 (I528041,I528435,I528613);
nand I_30948 (I528044,I528565,I528353);
nand I_30949 (I528658,I528175,I85412);
nor I_30950 (I528056,I528418,I528658);
not I_30951 (I528719,I2514);
DFFARX1 I_30952 (I413719,I2507,I528719,I528745,);
DFFARX1 I_30953 (I413713,I2507,I528719,I528762,);
not I_30954 (I528770,I528762);
not I_30955 (I528787,I413728);
nor I_30956 (I528804,I528787,I413713);
not I_30957 (I528821,I413722);
nor I_30958 (I528838,I528804,I413731);
nor I_30959 (I528855,I528762,I528838);
DFFARX1 I_30960 (I528855,I2507,I528719,I528705,);
nor I_30961 (I528886,I413731,I413713);
nand I_30962 (I528903,I528886,I413728);
DFFARX1 I_30963 (I528903,I2507,I528719,I528708,);
nor I_30964 (I528934,I528821,I413731);
nand I_30965 (I528951,I528934,I413716);
nor I_30966 (I528968,I528745,I528951);
DFFARX1 I_30967 (I528968,I2507,I528719,I528684,);
not I_30968 (I528999,I528951);
nand I_30969 (I528696,I528762,I528999);
DFFARX1 I_30970 (I528951,I2507,I528719,I529039,);
not I_30971 (I529047,I529039);
not I_30972 (I529064,I413731);
not I_30973 (I529081,I413725);
nor I_30974 (I529098,I529081,I413722);
nor I_30975 (I528711,I529047,I529098);
nor I_30976 (I529129,I529081,I413734);
and I_30977 (I529146,I529129,I413737);
or I_30978 (I529163,I529146,I413716);
DFFARX1 I_30979 (I529163,I2507,I528719,I529189,);
nor I_30980 (I528699,I529189,I528745);
not I_30981 (I529211,I529189);
and I_30982 (I529228,I529211,I528745);
nor I_30983 (I528693,I528770,I529228);
nand I_30984 (I529259,I529211,I528821);
nor I_30985 (I528687,I529081,I529259);
nand I_30986 (I528690,I529211,I528999);
nand I_30987 (I529304,I528821,I413725);
nor I_30988 (I528702,I529064,I529304);
not I_30989 (I529365,I2514);
DFFARX1 I_30990 (I248734,I2507,I529365,I529391,);
DFFARX1 I_30991 (I248731,I2507,I529365,I529408,);
not I_30992 (I529416,I529408);
not I_30993 (I529433,I248746);
nor I_30994 (I529450,I529433,I248749);
not I_30995 (I529467,I248737);
nor I_30996 (I529484,I529450,I248743);
nor I_30997 (I529501,I529408,I529484);
DFFARX1 I_30998 (I529501,I2507,I529365,I529351,);
nor I_30999 (I529532,I248743,I248749);
nand I_31000 (I529549,I529532,I248746);
DFFARX1 I_31001 (I529549,I2507,I529365,I529354,);
nor I_31002 (I529580,I529467,I248743);
nand I_31003 (I529597,I529580,I248755);
nor I_31004 (I529614,I529391,I529597);
DFFARX1 I_31005 (I529614,I2507,I529365,I529330,);
not I_31006 (I529645,I529597);
nand I_31007 (I529342,I529408,I529645);
DFFARX1 I_31008 (I529597,I2507,I529365,I529685,);
not I_31009 (I529693,I529685);
not I_31010 (I529710,I248743);
not I_31011 (I529727,I248728);
nor I_31012 (I529744,I529727,I248737);
nor I_31013 (I529357,I529693,I529744);
nor I_31014 (I529775,I529727,I248740);
and I_31015 (I529792,I529775,I248728);
or I_31016 (I529809,I529792,I248752);
DFFARX1 I_31017 (I529809,I2507,I529365,I529835,);
nor I_31018 (I529345,I529835,I529391);
not I_31019 (I529857,I529835);
and I_31020 (I529874,I529857,I529391);
nor I_31021 (I529339,I529416,I529874);
nand I_31022 (I529905,I529857,I529467);
nor I_31023 (I529333,I529727,I529905);
nand I_31024 (I529336,I529857,I529645);
nand I_31025 (I529950,I529467,I248728);
nor I_31026 (I529348,I529710,I529950);
not I_31027 (I530011,I2514);
DFFARX1 I_31028 (I240574,I2507,I530011,I530037,);
DFFARX1 I_31029 (I240571,I2507,I530011,I530054,);
not I_31030 (I530062,I530054);
not I_31031 (I530079,I240586);
nor I_31032 (I530096,I530079,I240589);
not I_31033 (I530113,I240577);
nor I_31034 (I530130,I530096,I240583);
nor I_31035 (I530147,I530054,I530130);
DFFARX1 I_31036 (I530147,I2507,I530011,I529997,);
nor I_31037 (I530178,I240583,I240589);
nand I_31038 (I530195,I530178,I240586);
DFFARX1 I_31039 (I530195,I2507,I530011,I530000,);
nor I_31040 (I530226,I530113,I240583);
nand I_31041 (I530243,I530226,I240595);
nor I_31042 (I530260,I530037,I530243);
DFFARX1 I_31043 (I530260,I2507,I530011,I529976,);
not I_31044 (I530291,I530243);
nand I_31045 (I529988,I530054,I530291);
DFFARX1 I_31046 (I530243,I2507,I530011,I530331,);
not I_31047 (I530339,I530331);
not I_31048 (I530356,I240583);
not I_31049 (I530373,I240568);
nor I_31050 (I530390,I530373,I240577);
nor I_31051 (I530003,I530339,I530390);
nor I_31052 (I530421,I530373,I240580);
and I_31053 (I530438,I530421,I240568);
or I_31054 (I530455,I530438,I240592);
DFFARX1 I_31055 (I530455,I2507,I530011,I530481,);
nor I_31056 (I529991,I530481,I530037);
not I_31057 (I530503,I530481);
and I_31058 (I530520,I530503,I530037);
nor I_31059 (I529985,I530062,I530520);
nand I_31060 (I530551,I530503,I530113);
nor I_31061 (I529979,I530373,I530551);
nand I_31062 (I529982,I530503,I530291);
nand I_31063 (I530596,I530113,I240568);
nor I_31064 (I529994,I530356,I530596);
not I_31065 (I530657,I2514);
DFFARX1 I_31066 (I6090,I2507,I530657,I530683,);
DFFARX1 I_31067 (I6087,I2507,I530657,I530700,);
not I_31068 (I530708,I530700);
not I_31069 (I530725,I6099);
nor I_31070 (I530742,I530725,I6096);
not I_31071 (I530759,I6105);
nor I_31072 (I530776,I530742,I6102);
nor I_31073 (I530793,I530700,I530776);
DFFARX1 I_31074 (I530793,I2507,I530657,I530643,);
nor I_31075 (I530824,I6102,I6096);
nand I_31076 (I530841,I530824,I6099);
DFFARX1 I_31077 (I530841,I2507,I530657,I530646,);
nor I_31078 (I530872,I530759,I6102);
nand I_31079 (I530889,I530872,I6093);
nor I_31080 (I530906,I530683,I530889);
DFFARX1 I_31081 (I530906,I2507,I530657,I530622,);
not I_31082 (I530937,I530889);
nand I_31083 (I530634,I530700,I530937);
DFFARX1 I_31084 (I530889,I2507,I530657,I530977,);
not I_31085 (I530985,I530977);
not I_31086 (I531002,I6102);
not I_31087 (I531019,I6093);
nor I_31088 (I531036,I531019,I6105);
nor I_31089 (I530649,I530985,I531036);
nor I_31090 (I531067,I531019,I6087);
and I_31091 (I531084,I531067,I6108);
or I_31092 (I531101,I531084,I6090);
DFFARX1 I_31093 (I531101,I2507,I530657,I531127,);
nor I_31094 (I530637,I531127,I530683);
not I_31095 (I531149,I531127);
and I_31096 (I531166,I531149,I530683);
nor I_31097 (I530631,I530708,I531166);
nand I_31098 (I531197,I531149,I530759);
nor I_31099 (I530625,I531019,I531197);
nand I_31100 (I530628,I531149,I530937);
nand I_31101 (I531242,I530759,I6093);
nor I_31102 (I530640,I531002,I531242);
not I_31103 (I531303,I2514);
DFFARX1 I_31104 (I544154,I2507,I531303,I531329,);
DFFARX1 I_31105 (I544157,I2507,I531303,I531346,);
not I_31106 (I531354,I531346);
not I_31107 (I531371,I544154);
nor I_31108 (I531388,I531371,I544166);
not I_31109 (I531405,I544175);
nor I_31110 (I531422,I531388,I544163);
nor I_31111 (I531439,I531346,I531422);
DFFARX1 I_31112 (I531439,I2507,I531303,I531289,);
nor I_31113 (I531470,I544163,I544166);
nand I_31114 (I531487,I531470,I544154);
DFFARX1 I_31115 (I531487,I2507,I531303,I531292,);
nor I_31116 (I531518,I531405,I544163);
nand I_31117 (I531535,I531518,I544169);
nor I_31118 (I531552,I531329,I531535);
DFFARX1 I_31119 (I531552,I2507,I531303,I531268,);
not I_31120 (I531583,I531535);
nand I_31121 (I531280,I531346,I531583);
DFFARX1 I_31122 (I531535,I2507,I531303,I531623,);
not I_31123 (I531631,I531623);
not I_31124 (I531648,I544163);
not I_31125 (I531665,I544160);
nor I_31126 (I531682,I531665,I544175);
nor I_31127 (I531295,I531631,I531682);
nor I_31128 (I531713,I531665,I544172);
and I_31129 (I531730,I531713,I544160);
or I_31130 (I531747,I531730,I544157);
DFFARX1 I_31131 (I531747,I2507,I531303,I531773,);
nor I_31132 (I531283,I531773,I531329);
not I_31133 (I531795,I531773);
and I_31134 (I531812,I531795,I531329);
nor I_31135 (I531277,I531354,I531812);
nand I_31136 (I531843,I531795,I531405);
nor I_31137 (I531271,I531665,I531843);
nand I_31138 (I531274,I531795,I531583);
nand I_31139 (I531888,I531405,I544160);
nor I_31140 (I531286,I531648,I531888);
not I_31141 (I531949,I2514);
DFFARX1 I_31142 (I647991,I2507,I531949,I531975,);
DFFARX1 I_31143 (I647997,I2507,I531949,I531992,);
not I_31144 (I532000,I531992);
not I_31145 (I532017,I647994);
nor I_31146 (I532034,I532017,I647973);
not I_31147 (I532051,I647976);
nor I_31148 (I532068,I532034,I647982);
nor I_31149 (I532085,I531992,I532068);
DFFARX1 I_31150 (I532085,I2507,I531949,I531935,);
nor I_31151 (I532116,I647982,I647973);
nand I_31152 (I532133,I532116,I647994);
DFFARX1 I_31153 (I532133,I2507,I531949,I531938,);
nor I_31154 (I532164,I532051,I647982);
nand I_31155 (I532181,I532164,I647976);
nor I_31156 (I532198,I531975,I532181);
DFFARX1 I_31157 (I532198,I2507,I531949,I531914,);
not I_31158 (I532229,I532181);
nand I_31159 (I531926,I531992,I532229);
DFFARX1 I_31160 (I532181,I2507,I531949,I532269,);
not I_31161 (I532277,I532269);
not I_31162 (I532294,I647982);
not I_31163 (I532311,I647985);
nor I_31164 (I532328,I532311,I647976);
nor I_31165 (I531941,I532277,I532328);
nor I_31166 (I532359,I532311,I647973);
and I_31167 (I532376,I532359,I647979);
or I_31168 (I532393,I532376,I647988);
DFFARX1 I_31169 (I532393,I2507,I531949,I532419,);
nor I_31170 (I531929,I532419,I531975);
not I_31171 (I532441,I532419);
and I_31172 (I532458,I532441,I531975);
nor I_31173 (I531923,I532000,I532458);
nand I_31174 (I532489,I532441,I532051);
nor I_31175 (I531917,I532311,I532489);
nand I_31176 (I531920,I532441,I532229);
nand I_31177 (I532534,I532051,I647985);
nor I_31178 (I531932,I532294,I532534);
not I_31179 (I532595,I2514);
DFFARX1 I_31180 (I716228,I2507,I532595,I532621,);
DFFARX1 I_31181 (I716252,I2507,I532595,I532638,);
not I_31182 (I532646,I532638);
not I_31183 (I532663,I716234);
nor I_31184 (I532680,I532663,I716243);
not I_31185 (I532697,I716228);
nor I_31186 (I532714,I532680,I716249);
nor I_31187 (I532731,I532638,I532714);
DFFARX1 I_31188 (I532731,I2507,I532595,I532581,);
nor I_31189 (I532762,I716249,I716243);
nand I_31190 (I532779,I532762,I716234);
DFFARX1 I_31191 (I532779,I2507,I532595,I532584,);
nor I_31192 (I532810,I532697,I716249);
nand I_31193 (I532827,I532810,I716246);
nor I_31194 (I532844,I532621,I532827);
DFFARX1 I_31195 (I532844,I2507,I532595,I532560,);
not I_31196 (I532875,I532827);
nand I_31197 (I532572,I532638,I532875);
DFFARX1 I_31198 (I532827,I2507,I532595,I532915,);
not I_31199 (I532923,I532915);
not I_31200 (I532940,I716249);
not I_31201 (I532957,I716240);
nor I_31202 (I532974,I532957,I716228);
nor I_31203 (I532587,I532923,I532974);
nor I_31204 (I533005,I532957,I716231);
and I_31205 (I533022,I533005,I716255);
or I_31206 (I533039,I533022,I716237);
DFFARX1 I_31207 (I533039,I2507,I532595,I533065,);
nor I_31208 (I532575,I533065,I532621);
not I_31209 (I533087,I533065);
and I_31210 (I533104,I533087,I532621);
nor I_31211 (I532569,I532646,I533104);
nand I_31212 (I533135,I533087,I532697);
nor I_31213 (I532563,I532957,I533135);
nand I_31214 (I532566,I533087,I532875);
nand I_31215 (I533180,I532697,I716240);
nor I_31216 (I532578,I532940,I533180);
not I_31217 (I533241,I2514);
DFFARX1 I_31218 (I350717,I2507,I533241,I533267,);
DFFARX1 I_31219 (I350711,I2507,I533241,I533284,);
not I_31220 (I533292,I533284);
not I_31221 (I533309,I350726);
nor I_31222 (I533326,I533309,I350711);
not I_31223 (I533343,I350720);
nor I_31224 (I533360,I533326,I350729);
nor I_31225 (I533377,I533284,I533360);
DFFARX1 I_31226 (I533377,I2507,I533241,I533227,);
nor I_31227 (I533408,I350729,I350711);
nand I_31228 (I533425,I533408,I350726);
DFFARX1 I_31229 (I533425,I2507,I533241,I533230,);
nor I_31230 (I533456,I533343,I350729);
nand I_31231 (I533473,I533456,I350714);
nor I_31232 (I533490,I533267,I533473);
DFFARX1 I_31233 (I533490,I2507,I533241,I533206,);
not I_31234 (I533521,I533473);
nand I_31235 (I533218,I533284,I533521);
DFFARX1 I_31236 (I533473,I2507,I533241,I533561,);
not I_31237 (I533569,I533561);
not I_31238 (I533586,I350729);
not I_31239 (I533603,I350723);
nor I_31240 (I533620,I533603,I350720);
nor I_31241 (I533233,I533569,I533620);
nor I_31242 (I533651,I533603,I350732);
and I_31243 (I533668,I533651,I350735);
or I_31244 (I533685,I533668,I350714);
DFFARX1 I_31245 (I533685,I2507,I533241,I533711,);
nor I_31246 (I533221,I533711,I533267);
not I_31247 (I533733,I533711);
and I_31248 (I533750,I533733,I533267);
nor I_31249 (I533215,I533292,I533750);
nand I_31250 (I533781,I533733,I533343);
nor I_31251 (I533209,I533603,I533781);
nand I_31252 (I533212,I533733,I533521);
nand I_31253 (I533826,I533343,I350723);
nor I_31254 (I533224,I533586,I533826);
not I_31255 (I533887,I2514);
DFFARX1 I_31256 (I64125,I2507,I533887,I533913,);
DFFARX1 I_31257 (I64131,I2507,I533887,I533930,);
not I_31258 (I533938,I533930);
not I_31259 (I533955,I64149);
nor I_31260 (I533972,I533955,I64128);
not I_31261 (I533989,I64134);
nor I_31262 (I534006,I533972,I64140);
nor I_31263 (I534023,I533930,I534006);
DFFARX1 I_31264 (I534023,I2507,I533887,I533873,);
nor I_31265 (I534054,I64140,I64128);
nand I_31266 (I534071,I534054,I64149);
DFFARX1 I_31267 (I534071,I2507,I533887,I533876,);
nor I_31268 (I534102,I533989,I64140);
nand I_31269 (I534119,I534102,I64146);
nor I_31270 (I534136,I533913,I534119);
DFFARX1 I_31271 (I534136,I2507,I533887,I533852,);
not I_31272 (I534167,I534119);
nand I_31273 (I533864,I533930,I534167);
DFFARX1 I_31274 (I534119,I2507,I533887,I534207,);
not I_31275 (I534215,I534207);
not I_31276 (I534232,I64140);
not I_31277 (I534249,I64128);
nor I_31278 (I534266,I534249,I64134);
nor I_31279 (I533879,I534215,I534266);
nor I_31280 (I534297,I534249,I64137);
and I_31281 (I534314,I534297,I64125);
or I_31282 (I534331,I534314,I64143);
DFFARX1 I_31283 (I534331,I2507,I533887,I534357,);
nor I_31284 (I533867,I534357,I533913);
not I_31285 (I534379,I534357);
and I_31286 (I534396,I534379,I533913);
nor I_31287 (I533861,I533938,I534396);
nand I_31288 (I534427,I534379,I533989);
nor I_31289 (I533855,I534249,I534427);
nand I_31290 (I533858,I534379,I534167);
nand I_31291 (I534472,I533989,I64128);
nor I_31292 (I533870,I534232,I534472);
not I_31293 (I534533,I2514);
DFFARX1 I_31294 (I409673,I2507,I534533,I534559,);
DFFARX1 I_31295 (I409667,I2507,I534533,I534576,);
not I_31296 (I534584,I534576);
not I_31297 (I534601,I409682);
nor I_31298 (I534618,I534601,I409667);
not I_31299 (I534635,I409676);
nor I_31300 (I534652,I534618,I409685);
nor I_31301 (I534669,I534576,I534652);
DFFARX1 I_31302 (I534669,I2507,I534533,I534519,);
nor I_31303 (I534700,I409685,I409667);
nand I_31304 (I534717,I534700,I409682);
DFFARX1 I_31305 (I534717,I2507,I534533,I534522,);
nor I_31306 (I534748,I534635,I409685);
nand I_31307 (I534765,I534748,I409670);
nor I_31308 (I534782,I534559,I534765);
DFFARX1 I_31309 (I534782,I2507,I534533,I534498,);
not I_31310 (I534813,I534765);
nand I_31311 (I534510,I534576,I534813);
DFFARX1 I_31312 (I534765,I2507,I534533,I534853,);
not I_31313 (I534861,I534853);
not I_31314 (I534878,I409685);
not I_31315 (I534895,I409679);
nor I_31316 (I534912,I534895,I409676);
nor I_31317 (I534525,I534861,I534912);
nor I_31318 (I534943,I534895,I409688);
and I_31319 (I534960,I534943,I409691);
or I_31320 (I534977,I534960,I409670);
DFFARX1 I_31321 (I534977,I2507,I534533,I535003,);
nor I_31322 (I534513,I535003,I534559);
not I_31323 (I535025,I535003);
and I_31324 (I535042,I535025,I534559);
nor I_31325 (I534507,I534584,I535042);
nand I_31326 (I535073,I535025,I534635);
nor I_31327 (I534501,I534895,I535073);
nand I_31328 (I534504,I535025,I534813);
nand I_31329 (I535118,I534635,I409679);
nor I_31330 (I534516,I534878,I535118);
not I_31331 (I535179,I2514);
DFFARX1 I_31332 (I67287,I2507,I535179,I535205,);
DFFARX1 I_31333 (I67293,I2507,I535179,I535222,);
not I_31334 (I535230,I535222);
not I_31335 (I535247,I67311);
nor I_31336 (I535264,I535247,I67290);
not I_31337 (I535281,I67296);
nor I_31338 (I535298,I535264,I67302);
nor I_31339 (I535315,I535222,I535298);
DFFARX1 I_31340 (I535315,I2507,I535179,I535165,);
nor I_31341 (I535346,I67302,I67290);
nand I_31342 (I535363,I535346,I67311);
DFFARX1 I_31343 (I535363,I2507,I535179,I535168,);
nor I_31344 (I535394,I535281,I67302);
nand I_31345 (I535411,I535394,I67308);
nor I_31346 (I535428,I535205,I535411);
DFFARX1 I_31347 (I535428,I2507,I535179,I535144,);
not I_31348 (I535459,I535411);
nand I_31349 (I535156,I535222,I535459);
DFFARX1 I_31350 (I535411,I2507,I535179,I535499,);
not I_31351 (I535507,I535499);
not I_31352 (I535524,I67302);
not I_31353 (I535541,I67290);
nor I_31354 (I535558,I535541,I67296);
nor I_31355 (I535171,I535507,I535558);
nor I_31356 (I535589,I535541,I67299);
and I_31357 (I535606,I535589,I67287);
or I_31358 (I535623,I535606,I67305);
DFFARX1 I_31359 (I535623,I2507,I535179,I535649,);
nor I_31360 (I535159,I535649,I535205);
not I_31361 (I535671,I535649);
and I_31362 (I535688,I535671,I535205);
nor I_31363 (I535153,I535230,I535688);
nand I_31364 (I535719,I535671,I535281);
nor I_31365 (I535147,I535541,I535719);
nand I_31366 (I535150,I535671,I535459);
nand I_31367 (I535764,I535281,I67290);
nor I_31368 (I535162,I535524,I535764);
not I_31369 (I535825,I2514);
DFFARX1 I_31370 (I247646,I2507,I535825,I535851,);
DFFARX1 I_31371 (I247643,I2507,I535825,I535868,);
not I_31372 (I535876,I535868);
not I_31373 (I535893,I247658);
nor I_31374 (I535910,I535893,I247661);
not I_31375 (I535927,I247649);
nor I_31376 (I535944,I535910,I247655);
nor I_31377 (I535961,I535868,I535944);
DFFARX1 I_31378 (I535961,I2507,I535825,I535811,);
nor I_31379 (I535992,I247655,I247661);
nand I_31380 (I536009,I535992,I247658);
DFFARX1 I_31381 (I536009,I2507,I535825,I535814,);
nor I_31382 (I536040,I535927,I247655);
nand I_31383 (I536057,I536040,I247667);
nor I_31384 (I536074,I535851,I536057);
DFFARX1 I_31385 (I536074,I2507,I535825,I535790,);
not I_31386 (I536105,I536057);
nand I_31387 (I535802,I535868,I536105);
DFFARX1 I_31388 (I536057,I2507,I535825,I536145,);
not I_31389 (I536153,I536145);
not I_31390 (I536170,I247655);
not I_31391 (I536187,I247640);
nor I_31392 (I536204,I536187,I247649);
nor I_31393 (I535817,I536153,I536204);
nor I_31394 (I536235,I536187,I247652);
and I_31395 (I536252,I536235,I247640);
or I_31396 (I536269,I536252,I247664);
DFFARX1 I_31397 (I536269,I2507,I535825,I536295,);
nor I_31398 (I535805,I536295,I535851);
not I_31399 (I536317,I536295);
and I_31400 (I536334,I536317,I535851);
nor I_31401 (I535799,I535876,I536334);
nand I_31402 (I536365,I536317,I535927);
nor I_31403 (I535793,I536187,I536365);
nand I_31404 (I535796,I536317,I536105);
nand I_31405 (I536410,I535927,I247640);
nor I_31406 (I535808,I536170,I536410);
not I_31407 (I536471,I2514);
DFFARX1 I_31408 (I354185,I2507,I536471,I536497,);
DFFARX1 I_31409 (I354179,I2507,I536471,I536514,);
not I_31410 (I536522,I536514);
not I_31411 (I536539,I354194);
nor I_31412 (I536556,I536539,I354179);
not I_31413 (I536573,I354188);
nor I_31414 (I536590,I536556,I354197);
nor I_31415 (I536607,I536514,I536590);
DFFARX1 I_31416 (I536607,I2507,I536471,I536457,);
nor I_31417 (I536638,I354197,I354179);
nand I_31418 (I536655,I536638,I354194);
DFFARX1 I_31419 (I536655,I2507,I536471,I536460,);
nor I_31420 (I536686,I536573,I354197);
nand I_31421 (I536703,I536686,I354182);
nor I_31422 (I536720,I536497,I536703);
DFFARX1 I_31423 (I536720,I2507,I536471,I536436,);
not I_31424 (I536751,I536703);
nand I_31425 (I536448,I536514,I536751);
DFFARX1 I_31426 (I536703,I2507,I536471,I536791,);
not I_31427 (I536799,I536791);
not I_31428 (I536816,I354197);
not I_31429 (I536833,I354191);
nor I_31430 (I536850,I536833,I354188);
nor I_31431 (I536463,I536799,I536850);
nor I_31432 (I536881,I536833,I354200);
and I_31433 (I536898,I536881,I354203);
or I_31434 (I536915,I536898,I354182);
DFFARX1 I_31435 (I536915,I2507,I536471,I536941,);
nor I_31436 (I536451,I536941,I536497);
not I_31437 (I536963,I536941);
and I_31438 (I536980,I536963,I536497);
nor I_31439 (I536445,I536522,I536980);
nand I_31440 (I537011,I536963,I536573);
nor I_31441 (I536439,I536833,I537011);
nand I_31442 (I536442,I536963,I536751);
nand I_31443 (I537056,I536573,I354191);
nor I_31444 (I536454,I536816,I537056);
not I_31445 (I537117,I2514);
DFFARX1 I_31446 (I662135,I2507,I537117,I537143,);
DFFARX1 I_31447 (I662141,I2507,I537117,I537160,);
not I_31448 (I537168,I537160);
not I_31449 (I537185,I662138);
nor I_31450 (I537202,I537185,I662117);
not I_31451 (I537219,I662120);
nor I_31452 (I537236,I537202,I662126);
nor I_31453 (I537253,I537160,I537236);
DFFARX1 I_31454 (I537253,I2507,I537117,I537103,);
nor I_31455 (I537284,I662126,I662117);
nand I_31456 (I537301,I537284,I662138);
DFFARX1 I_31457 (I537301,I2507,I537117,I537106,);
nor I_31458 (I537332,I537219,I662126);
nand I_31459 (I537349,I537332,I662120);
nor I_31460 (I537366,I537143,I537349);
DFFARX1 I_31461 (I537366,I2507,I537117,I537082,);
not I_31462 (I537397,I537349);
nand I_31463 (I537094,I537160,I537397);
DFFARX1 I_31464 (I537349,I2507,I537117,I537437,);
not I_31465 (I537445,I537437);
not I_31466 (I537462,I662126);
not I_31467 (I537479,I662129);
nor I_31468 (I537496,I537479,I662120);
nor I_31469 (I537109,I537445,I537496);
nor I_31470 (I537527,I537479,I662117);
and I_31471 (I537544,I537527,I662123);
or I_31472 (I537561,I537544,I662132);
DFFARX1 I_31473 (I537561,I2507,I537117,I537587,);
nor I_31474 (I537097,I537587,I537143);
not I_31475 (I537609,I537587);
and I_31476 (I537626,I537609,I537143);
nor I_31477 (I537091,I537168,I537626);
nand I_31478 (I537657,I537609,I537219);
nor I_31479 (I537085,I537479,I537657);
nand I_31480 (I537088,I537609,I537397);
nand I_31481 (I537702,I537219,I662129);
nor I_31482 (I537100,I537462,I537702);
not I_31483 (I537763,I2514);
DFFARX1 I_31484 (I687224,I2507,I537763,I537789,);
DFFARX1 I_31485 (I687221,I2507,I537763,I537806,);
not I_31486 (I537814,I537806);
not I_31487 (I537831,I687218);
nor I_31488 (I537848,I537831,I687209);
not I_31489 (I537865,I687230);
nor I_31490 (I537882,I537848,I687209);
nor I_31491 (I537899,I537806,I537882);
DFFARX1 I_31492 (I537899,I2507,I537763,I537749,);
nor I_31493 (I537930,I687209,I687209);
nand I_31494 (I537947,I537930,I687218);
DFFARX1 I_31495 (I537947,I2507,I537763,I537752,);
nor I_31496 (I537978,I537865,I687209);
nand I_31497 (I537995,I537978,I687233);
nor I_31498 (I538012,I537789,I537995);
DFFARX1 I_31499 (I538012,I2507,I537763,I537728,);
not I_31500 (I538043,I537995);
nand I_31501 (I537740,I537806,I538043);
DFFARX1 I_31502 (I537995,I2507,I537763,I538083,);
not I_31503 (I538091,I538083);
not I_31504 (I538108,I687209);
not I_31505 (I538125,I687212);
nor I_31506 (I538142,I538125,I687230);
nor I_31507 (I537755,I538091,I538142);
nor I_31508 (I538173,I538125,I687215);
and I_31509 (I538190,I538173,I687236);
or I_31510 (I538207,I538190,I687227);
DFFARX1 I_31511 (I538207,I2507,I537763,I538233,);
nor I_31512 (I537743,I538233,I537789);
not I_31513 (I538255,I538233);
and I_31514 (I538272,I538255,I537789);
nor I_31515 (I537737,I537814,I538272);
nand I_31516 (I538303,I538255,I537865);
nor I_31517 (I537731,I538125,I538303);
nand I_31518 (I537734,I538255,I538043);
nand I_31519 (I538348,I537865,I687212);
nor I_31520 (I537746,I538108,I538348);
not I_31521 (I538409,I2514);
DFFARX1 I_31522 (I263966,I2507,I538409,I538435,);
DFFARX1 I_31523 (I263963,I2507,I538409,I538452,);
not I_31524 (I538460,I538452);
not I_31525 (I538477,I263978);
nor I_31526 (I538494,I538477,I263981);
not I_31527 (I538511,I263969);
nor I_31528 (I538528,I538494,I263975);
nor I_31529 (I538545,I538452,I538528);
DFFARX1 I_31530 (I538545,I2507,I538409,I538395,);
nor I_31531 (I538576,I263975,I263981);
nand I_31532 (I538593,I538576,I263978);
DFFARX1 I_31533 (I538593,I2507,I538409,I538398,);
nor I_31534 (I538624,I538511,I263975);
nand I_31535 (I538641,I538624,I263987);
nor I_31536 (I538658,I538435,I538641);
DFFARX1 I_31537 (I538658,I2507,I538409,I538374,);
not I_31538 (I538689,I538641);
nand I_31539 (I538386,I538452,I538689);
DFFARX1 I_31540 (I538641,I2507,I538409,I538729,);
not I_31541 (I538737,I538729);
not I_31542 (I538754,I263975);
not I_31543 (I538771,I263960);
nor I_31544 (I538788,I538771,I263969);
nor I_31545 (I538401,I538737,I538788);
nor I_31546 (I538819,I538771,I263972);
and I_31547 (I538836,I538819,I263960);
or I_31548 (I538853,I538836,I263984);
DFFARX1 I_31549 (I538853,I2507,I538409,I538879,);
nor I_31550 (I538389,I538879,I538435);
not I_31551 (I538901,I538879);
and I_31552 (I538918,I538901,I538435);
nor I_31553 (I538383,I538460,I538918);
nand I_31554 (I538949,I538901,I538511);
nor I_31555 (I538377,I538771,I538949);
nand I_31556 (I538380,I538901,I538689);
nand I_31557 (I538994,I538511,I263960);
nor I_31558 (I538392,I538754,I538994);
not I_31559 (I539055,I2514);
DFFARX1 I_31560 (I331062,I2507,I539055,I539081,);
DFFARX1 I_31561 (I331074,I2507,I539055,I539098,);
not I_31562 (I539106,I539098);
not I_31563 (I539123,I331083);
nor I_31564 (I539140,I539123,I331059);
not I_31565 (I539157,I331077);
nor I_31566 (I539174,I539140,I331071);
nor I_31567 (I539191,I539098,I539174);
DFFARX1 I_31568 (I539191,I2507,I539055,I539041,);
nor I_31569 (I539222,I331071,I331059);
nand I_31570 (I539239,I539222,I331083);
DFFARX1 I_31571 (I539239,I2507,I539055,I539044,);
nor I_31572 (I539270,I539157,I331071);
nand I_31573 (I539287,I539270,I331065);
nor I_31574 (I539304,I539081,I539287);
DFFARX1 I_31575 (I539304,I2507,I539055,I539020,);
not I_31576 (I539335,I539287);
nand I_31577 (I539032,I539098,I539335);
DFFARX1 I_31578 (I539287,I2507,I539055,I539375,);
not I_31579 (I539383,I539375);
not I_31580 (I539400,I331071);
not I_31581 (I539417,I331080);
nor I_31582 (I539434,I539417,I331077);
nor I_31583 (I539047,I539383,I539434);
nor I_31584 (I539465,I539417,I331062);
and I_31585 (I539482,I539465,I331059);
or I_31586 (I539499,I539482,I331068);
DFFARX1 I_31587 (I539499,I2507,I539055,I539525,);
nor I_31588 (I539035,I539525,I539081);
not I_31589 (I539547,I539525);
and I_31590 (I539564,I539547,I539081);
nor I_31591 (I539029,I539106,I539564);
nand I_31592 (I539595,I539547,I539157);
nor I_31593 (I539023,I539417,I539595);
nand I_31594 (I539026,I539547,I539335);
nand I_31595 (I539640,I539157,I331080);
nor I_31596 (I539038,I539400,I539640);
not I_31597 (I539695,I2514);
DFFARX1 I_31598 (I249840,I2507,I539695,I539721,);
DFFARX1 I_31599 (I539721,I2507,I539695,I539738,);
not I_31600 (I539687,I539738);
not I_31601 (I539760,I539721);
DFFARX1 I_31602 (I249828,I2507,I539695,I539786,);
nand I_31603 (I539794,I539786,I249834);
not I_31604 (I539811,I249834);
not I_31605 (I539828,I249831);
nand I_31606 (I539845,I249819,I249816);
and I_31607 (I539862,I249819,I249816);
not I_31608 (I539879,I249843);
nand I_31609 (I539896,I539879,I539828);
nor I_31610 (I539669,I539896,I539794);
nor I_31611 (I539927,I539811,I539896);
nand I_31612 (I539672,I539862,I539927);
not I_31613 (I539958,I249816);
nor I_31614 (I539975,I539958,I249819);
nor I_31615 (I539992,I539975,I249843);
nor I_31616 (I540009,I539760,I539992);
DFFARX1 I_31617 (I540009,I2507,I539695,I539681,);
not I_31618 (I540040,I539975);
DFFARX1 I_31619 (I540040,I2507,I539695,I539684,);
and I_31620 (I539678,I539786,I539975);
nor I_31621 (I540085,I539958,I249825);
and I_31622 (I540102,I540085,I249822);
or I_31623 (I540119,I540102,I249837);
DFFARX1 I_31624 (I540119,I2507,I539695,I540145,);
nor I_31625 (I540153,I540145,I539879);
DFFARX1 I_31626 (I540153,I2507,I539695,I539666,);
nand I_31627 (I540184,I540145,I539786);
nand I_31628 (I540201,I539879,I540184);
nor I_31629 (I539675,I540201,I539845);
not I_31630 (I540256,I2514);
DFFARX1 I_31631 (I20402,I2507,I540256,I540282,);
DFFARX1 I_31632 (I540282,I2507,I540256,I540299,);
not I_31633 (I540248,I540299);
not I_31634 (I540321,I540282);
DFFARX1 I_31635 (I20387,I2507,I540256,I540347,);
nand I_31636 (I540355,I540347,I20399);
not I_31637 (I540372,I20399);
not I_31638 (I540389,I20405);
nand I_31639 (I540406,I20393,I20384);
and I_31640 (I540423,I20393,I20384);
not I_31641 (I540440,I20390);
nand I_31642 (I540457,I540440,I540389);
nor I_31643 (I540230,I540457,I540355);
nor I_31644 (I540488,I540372,I540457);
nand I_31645 (I540233,I540423,I540488);
not I_31646 (I540519,I20396);
nor I_31647 (I540536,I540519,I20393);
nor I_31648 (I540553,I540536,I20390);
nor I_31649 (I540570,I540321,I540553);
DFFARX1 I_31650 (I540570,I2507,I540256,I540242,);
not I_31651 (I540601,I540536);
DFFARX1 I_31652 (I540601,I2507,I540256,I540245,);
and I_31653 (I540239,I540347,I540536);
nor I_31654 (I540646,I540519,I20384);
and I_31655 (I540663,I540646,I20408);
or I_31656 (I540680,I540663,I20387);
DFFARX1 I_31657 (I540680,I2507,I540256,I540706,);
nor I_31658 (I540714,I540706,I540440);
DFFARX1 I_31659 (I540714,I2507,I540256,I540227,);
nand I_31660 (I540745,I540706,I540347);
nand I_31661 (I540762,I540440,I540745);
nor I_31662 (I540236,I540762,I540406);
not I_31663 (I540817,I2514);
DFFARX1 I_31664 (I324701,I2507,I540817,I540843,);
DFFARX1 I_31665 (I540843,I2507,I540817,I540860,);
not I_31666 (I540809,I540860);
not I_31667 (I540882,I540843);
DFFARX1 I_31668 (I324716,I2507,I540817,I540908,);
nand I_31669 (I540916,I540908,I324707);
not I_31670 (I540933,I324707);
not I_31671 (I540950,I324713);
nand I_31672 (I540967,I324710,I324719);
and I_31673 (I540984,I324710,I324719);
not I_31674 (I541001,I324704);
nand I_31675 (I541018,I541001,I540950);
nor I_31676 (I540791,I541018,I540916);
nor I_31677 (I541049,I540933,I541018);
nand I_31678 (I540794,I540984,I541049);
not I_31679 (I541080,I324701);
nor I_31680 (I541097,I541080,I324710);
nor I_31681 (I541114,I541097,I324704);
nor I_31682 (I541131,I540882,I541114);
DFFARX1 I_31683 (I541131,I2507,I540817,I540803,);
not I_31684 (I541162,I541097);
DFFARX1 I_31685 (I541162,I2507,I540817,I540806,);
and I_31686 (I540800,I540908,I541097);
nor I_31687 (I541207,I541080,I324725);
and I_31688 (I541224,I541207,I324704);
or I_31689 (I541241,I541224,I324722);
DFFARX1 I_31690 (I541241,I2507,I540817,I541267,);
nor I_31691 (I541275,I541267,I541001);
DFFARX1 I_31692 (I541275,I2507,I540817,I540788,);
nand I_31693 (I541306,I541267,I540908);
nand I_31694 (I541323,I541001,I541306);
nor I_31695 (I540797,I541323,I540967);
not I_31696 (I541378,I2514);
DFFARX1 I_31697 (I396376,I2507,I541378,I541404,);
DFFARX1 I_31698 (I541404,I2507,I541378,I541421,);
not I_31699 (I541370,I541421);
not I_31700 (I541443,I541404);
DFFARX1 I_31701 (I396388,I2507,I541378,I541469,);
nand I_31702 (I541477,I541469,I396397);
not I_31703 (I541494,I396397);
not I_31704 (I541511,I396379);
nand I_31705 (I541528,I396382,I396373);
and I_31706 (I541545,I396382,I396373);
not I_31707 (I541562,I396391);
nand I_31708 (I541579,I541562,I541511);
nor I_31709 (I541352,I541579,I541477);
nor I_31710 (I541610,I541494,I541579);
nand I_31711 (I541355,I541545,I541610);
not I_31712 (I541641,I396394);
nor I_31713 (I541658,I541641,I396382);
nor I_31714 (I541675,I541658,I396391);
nor I_31715 (I541692,I541443,I541675);
DFFARX1 I_31716 (I541692,I2507,I541378,I541364,);
not I_31717 (I541723,I541658);
DFFARX1 I_31718 (I541723,I2507,I541378,I541367,);
and I_31719 (I541361,I541469,I541658);
nor I_31720 (I541768,I541641,I396373);
and I_31721 (I541785,I541768,I396385);
or I_31722 (I541802,I541785,I396376);
DFFARX1 I_31723 (I541802,I2507,I541378,I541828,);
nor I_31724 (I541836,I541828,I541562);
DFFARX1 I_31725 (I541836,I2507,I541378,I541349,);
nand I_31726 (I541867,I541828,I541469);
nand I_31727 (I541884,I541562,I541867);
nor I_31728 (I541358,I541884,I541528);
not I_31729 (I541939,I2514);
DFFARX1 I_31730 (I301003,I2507,I541939,I541965,);
DFFARX1 I_31731 (I541965,I2507,I541939,I541982,);
not I_31732 (I541931,I541982);
not I_31733 (I542004,I541965);
DFFARX1 I_31734 (I301018,I2507,I541939,I542030,);
nand I_31735 (I542038,I542030,I301009);
not I_31736 (I542055,I301009);
not I_31737 (I542072,I301015);
nand I_31738 (I542089,I301012,I301021);
and I_31739 (I542106,I301012,I301021);
not I_31740 (I542123,I301006);
nand I_31741 (I542140,I542123,I542072);
nor I_31742 (I541913,I542140,I542038);
nor I_31743 (I542171,I542055,I542140);
nand I_31744 (I541916,I542106,I542171);
not I_31745 (I542202,I301003);
nor I_31746 (I542219,I542202,I301012);
nor I_31747 (I542236,I542219,I301006);
nor I_31748 (I542253,I542004,I542236);
DFFARX1 I_31749 (I542253,I2507,I541939,I541925,);
not I_31750 (I542284,I542219);
DFFARX1 I_31751 (I542284,I2507,I541939,I541928,);
and I_31752 (I541922,I542030,I542219);
nor I_31753 (I542329,I542202,I301027);
and I_31754 (I542346,I542329,I301006);
or I_31755 (I542363,I542346,I301024);
DFFARX1 I_31756 (I542363,I2507,I541939,I542389,);
nor I_31757 (I542397,I542389,I542123);
DFFARX1 I_31758 (I542397,I2507,I541939,I541910,);
nand I_31759 (I542428,I542389,I542030);
nand I_31760 (I542445,I542123,I542428);
nor I_31761 (I541919,I542445,I542089);
not I_31762 (I542500,I2514);
DFFARX1 I_31763 (I615042,I2507,I542500,I542526,);
DFFARX1 I_31764 (I542526,I2507,I542500,I542543,);
not I_31765 (I542492,I542543);
not I_31766 (I542565,I542526);
DFFARX1 I_31767 (I615033,I2507,I542500,I542591,);
nand I_31768 (I542599,I542591,I615030);
not I_31769 (I542616,I615030);
not I_31770 (I542633,I615039);
nand I_31771 (I542650,I615048,I615030);
and I_31772 (I542667,I615048,I615030);
not I_31773 (I542684,I615027);
nand I_31774 (I542701,I542684,I542633);
nor I_31775 (I542474,I542701,I542599);
nor I_31776 (I542732,I542616,I542701);
nand I_31777 (I542477,I542667,I542732);
not I_31778 (I542763,I615036);
nor I_31779 (I542780,I542763,I615048);
nor I_31780 (I542797,I542780,I615027);
nor I_31781 (I542814,I542565,I542797);
DFFARX1 I_31782 (I542814,I2507,I542500,I542486,);
not I_31783 (I542845,I542780);
DFFARX1 I_31784 (I542845,I2507,I542500,I542489,);
and I_31785 (I542483,I542591,I542780);
nor I_31786 (I542890,I542763,I615051);
and I_31787 (I542907,I542890,I615027);
or I_31788 (I542924,I542907,I615045);
DFFARX1 I_31789 (I542924,I2507,I542500,I542950,);
nor I_31790 (I542958,I542950,I542684);
DFFARX1 I_31791 (I542958,I2507,I542500,I542471,);
nand I_31792 (I542989,I542950,I542591);
nand I_31793 (I543006,I542684,I542989);
nor I_31794 (I542480,I543006,I542650);
not I_31795 (I543061,I2514);
DFFARX1 I_31796 (I311407,I2507,I543061,I543087,);
DFFARX1 I_31797 (I543087,I2507,I543061,I543104,);
not I_31798 (I543053,I543104);
not I_31799 (I543126,I543087);
DFFARX1 I_31800 (I311422,I2507,I543061,I543152,);
nand I_31801 (I543160,I543152,I311413);
not I_31802 (I543177,I311413);
not I_31803 (I543194,I311419);
nand I_31804 (I543211,I311416,I311425);
and I_31805 (I543228,I311416,I311425);
not I_31806 (I543245,I311410);
nand I_31807 (I543262,I543245,I543194);
nor I_31808 (I543035,I543262,I543160);
nor I_31809 (I543293,I543177,I543262);
nand I_31810 (I543038,I543228,I543293);
not I_31811 (I543324,I311407);
nor I_31812 (I543341,I543324,I311416);
nor I_31813 (I543358,I543341,I311410);
nor I_31814 (I543375,I543126,I543358);
DFFARX1 I_31815 (I543375,I2507,I543061,I543047,);
not I_31816 (I543406,I543341);
DFFARX1 I_31817 (I543406,I2507,I543061,I543050,);
and I_31818 (I543044,I543152,I543341);
nor I_31819 (I543451,I543324,I311431);
and I_31820 (I543468,I543451,I311410);
or I_31821 (I543485,I543468,I311428);
DFFARX1 I_31822 (I543485,I2507,I543061,I543511,);
nor I_31823 (I543519,I543511,I543245);
DFFARX1 I_31824 (I543519,I2507,I543061,I543032,);
nand I_31825 (I543550,I543511,I543152);
nand I_31826 (I543567,I543245,I543550);
nor I_31827 (I543041,I543567,I543211);
not I_31828 (I543622,I2514);
DFFARX1 I_31829 (I162712,I2507,I543622,I543648,);
DFFARX1 I_31830 (I543648,I2507,I543622,I543665,);
not I_31831 (I543614,I543665);
not I_31832 (I543687,I543648);
DFFARX1 I_31833 (I162709,I2507,I543622,I543713,);
nand I_31834 (I543721,I543713,I162703);
not I_31835 (I543738,I162703);
not I_31836 (I543755,I162700);
nand I_31837 (I543772,I162694,I162691);
and I_31838 (I543789,I162694,I162691);
not I_31839 (I543806,I162706);
nand I_31840 (I543823,I543806,I543755);
nor I_31841 (I543596,I543823,I543721);
nor I_31842 (I543854,I543738,I543823);
nand I_31843 (I543599,I543789,I543854);
not I_31844 (I543885,I162718);
nor I_31845 (I543902,I543885,I162694);
nor I_31846 (I543919,I543902,I162706);
nor I_31847 (I543936,I543687,I543919);
DFFARX1 I_31848 (I543936,I2507,I543622,I543608,);
not I_31849 (I543967,I543902);
DFFARX1 I_31850 (I543967,I2507,I543622,I543611,);
and I_31851 (I543605,I543713,I543902);
nor I_31852 (I544012,I543885,I162715);
and I_31853 (I544029,I544012,I162691);
or I_31854 (I544046,I544029,I162697);
DFFARX1 I_31855 (I544046,I2507,I543622,I544072,);
nor I_31856 (I544080,I544072,I543806);
DFFARX1 I_31857 (I544080,I2507,I543622,I543593,);
nand I_31858 (I544111,I544072,I543713);
nand I_31859 (I544128,I543806,I544111);
nor I_31860 (I543602,I544128,I543772);
not I_31861 (I544183,I2514);
DFFARX1 I_31862 (I262896,I2507,I544183,I544209,);
DFFARX1 I_31863 (I544209,I2507,I544183,I544226,);
not I_31864 (I544175,I544226);
not I_31865 (I544248,I544209);
DFFARX1 I_31866 (I262884,I2507,I544183,I544274,);
nand I_31867 (I544282,I544274,I262890);
not I_31868 (I544299,I262890);
not I_31869 (I544316,I262887);
nand I_31870 (I544333,I262875,I262872);
and I_31871 (I544350,I262875,I262872);
not I_31872 (I544367,I262899);
nand I_31873 (I544384,I544367,I544316);
nor I_31874 (I544157,I544384,I544282);
nor I_31875 (I544415,I544299,I544384);
nand I_31876 (I544160,I544350,I544415);
not I_31877 (I544446,I262872);
nor I_31878 (I544463,I544446,I262875);
nor I_31879 (I544480,I544463,I262899);
nor I_31880 (I544497,I544248,I544480);
DFFARX1 I_31881 (I544497,I2507,I544183,I544169,);
not I_31882 (I544528,I544463);
DFFARX1 I_31883 (I544528,I2507,I544183,I544172,);
and I_31884 (I544166,I544274,I544463);
nor I_31885 (I544573,I544446,I262881);
and I_31886 (I544590,I544573,I262878);
or I_31887 (I544607,I544590,I262893);
DFFARX1 I_31888 (I544607,I2507,I544183,I544633,);
nor I_31889 (I544641,I544633,I544367);
DFFARX1 I_31890 (I544641,I2507,I544183,I544154,);
nand I_31891 (I544672,I544633,I544274);
nand I_31892 (I544689,I544367,I544672);
nor I_31893 (I544163,I544689,I544333);
not I_31894 (I544744,I2514);
DFFARX1 I_31895 (I495738,I2507,I544744,I544770,);
DFFARX1 I_31896 (I544770,I2507,I544744,I544787,);
not I_31897 (I544736,I544787);
not I_31898 (I544809,I544770);
DFFARX1 I_31899 (I495765,I2507,I544744,I544835,);
nand I_31900 (I544843,I544835,I495756);
not I_31901 (I544860,I495756);
not I_31902 (I544877,I495738);
nand I_31903 (I544894,I495750,I495753);
and I_31904 (I544911,I495750,I495753);
not I_31905 (I544928,I495762);
nand I_31906 (I544945,I544928,I544877);
nor I_31907 (I544718,I544945,I544843);
nor I_31908 (I544976,I544860,I544945);
nand I_31909 (I544721,I544911,I544976);
not I_31910 (I545007,I495747);
nor I_31911 (I545024,I545007,I495750);
nor I_31912 (I545041,I545024,I495762);
nor I_31913 (I545058,I544809,I545041);
DFFARX1 I_31914 (I545058,I2507,I544744,I544730,);
not I_31915 (I545089,I545024);
DFFARX1 I_31916 (I545089,I2507,I544744,I544733,);
and I_31917 (I544727,I544835,I545024);
nor I_31918 (I545134,I545007,I495741);
and I_31919 (I545151,I545134,I495744);
or I_31920 (I545168,I545151,I495759);
DFFARX1 I_31921 (I545168,I2507,I544744,I545194,);
nor I_31922 (I545202,I545194,I544928);
DFFARX1 I_31923 (I545202,I2507,I544744,I544715,);
nand I_31924 (I545233,I545194,I544835);
nand I_31925 (I545250,I544928,I545233);
nor I_31926 (I544724,I545250,I544894);
not I_31927 (I545305,I2514);
DFFARX1 I_31928 (I584986,I2507,I545305,I545331,);
DFFARX1 I_31929 (I545331,I2507,I545305,I545348,);
not I_31930 (I545297,I545348);
not I_31931 (I545370,I545331);
DFFARX1 I_31932 (I584977,I2507,I545305,I545396,);
nand I_31933 (I545404,I545396,I584974);
not I_31934 (I545421,I584974);
not I_31935 (I545438,I584983);
nand I_31936 (I545455,I584992,I584974);
and I_31937 (I545472,I584992,I584974);
not I_31938 (I545489,I584971);
nand I_31939 (I545506,I545489,I545438);
nor I_31940 (I545279,I545506,I545404);
nor I_31941 (I545537,I545421,I545506);
nand I_31942 (I545282,I545472,I545537);
not I_31943 (I545568,I584980);
nor I_31944 (I545585,I545568,I584992);
nor I_31945 (I545602,I545585,I584971);
nor I_31946 (I545619,I545370,I545602);
DFFARX1 I_31947 (I545619,I2507,I545305,I545291,);
not I_31948 (I545650,I545585);
DFFARX1 I_31949 (I545650,I2507,I545305,I545294,);
and I_31950 (I545288,I545396,I545585);
nor I_31951 (I545695,I545568,I584995);
and I_31952 (I545712,I545695,I584971);
or I_31953 (I545729,I545712,I584989);
DFFARX1 I_31954 (I545729,I2507,I545305,I545755,);
nor I_31955 (I545763,I545755,I545489);
DFFARX1 I_31956 (I545763,I2507,I545305,I545276,);
nand I_31957 (I545794,I545755,I545396);
nand I_31958 (I545811,I545489,I545794);
nor I_31959 (I545285,I545811,I545455);
not I_31960 (I545866,I2514);
DFFARX1 I_31961 (I372678,I2507,I545866,I545892,);
DFFARX1 I_31962 (I545892,I2507,I545866,I545909,);
not I_31963 (I545858,I545909);
not I_31964 (I545931,I545892);
DFFARX1 I_31965 (I372690,I2507,I545866,I545957,);
nand I_31966 (I545965,I545957,I372699);
not I_31967 (I545982,I372699);
not I_31968 (I545999,I372681);
nand I_31969 (I546016,I372684,I372675);
and I_31970 (I546033,I372684,I372675);
not I_31971 (I546050,I372693);
nand I_31972 (I546067,I546050,I545999);
nor I_31973 (I545840,I546067,I545965);
nor I_31974 (I546098,I545982,I546067);
nand I_31975 (I545843,I546033,I546098);
not I_31976 (I546129,I372696);
nor I_31977 (I546146,I546129,I372684);
nor I_31978 (I546163,I546146,I372693);
nor I_31979 (I546180,I545931,I546163);
DFFARX1 I_31980 (I546180,I2507,I545866,I545852,);
not I_31981 (I546211,I546146);
DFFARX1 I_31982 (I546211,I2507,I545866,I545855,);
and I_31983 (I545849,I545957,I546146);
nor I_31984 (I546256,I546129,I372675);
and I_31985 (I546273,I546256,I372687);
or I_31986 (I546290,I546273,I372678);
DFFARX1 I_31987 (I546290,I2507,I545866,I546316,);
nor I_31988 (I546324,I546316,I546050);
DFFARX1 I_31989 (I546324,I2507,I545866,I545837,);
nand I_31990 (I546355,I546316,I545957);
nand I_31991 (I546372,I546050,I546355);
nor I_31992 (I545846,I546372,I546016);
not I_31993 (I546427,I2514);
DFFARX1 I_31994 (I53597,I2507,I546427,I546453,);
DFFARX1 I_31995 (I546453,I2507,I546427,I546470,);
not I_31996 (I546419,I546470);
not I_31997 (I546492,I546453);
DFFARX1 I_31998 (I53585,I2507,I546427,I546518,);
nand I_31999 (I546526,I546518,I53600);
not I_32000 (I546543,I53600);
not I_32001 (I546560,I53588);
nand I_32002 (I546577,I53609,I53603);
and I_32003 (I546594,I53609,I53603);
not I_32004 (I546611,I53591);
nand I_32005 (I546628,I546611,I546560);
nor I_32006 (I546401,I546628,I546526);
nor I_32007 (I546659,I546543,I546628);
nand I_32008 (I546404,I546594,I546659);
not I_32009 (I546690,I53594);
nor I_32010 (I546707,I546690,I53609);
nor I_32011 (I546724,I546707,I53591);
nor I_32012 (I546741,I546492,I546724);
DFFARX1 I_32013 (I546741,I2507,I546427,I546413,);
not I_32014 (I546772,I546707);
DFFARX1 I_32015 (I546772,I2507,I546427,I546416,);
and I_32016 (I546410,I546518,I546707);
nor I_32017 (I546817,I546690,I53588);
and I_32018 (I546834,I546817,I53585);
or I_32019 (I546851,I546834,I53606);
DFFARX1 I_32020 (I546851,I2507,I546427,I546877,);
nor I_32021 (I546885,I546877,I546611);
DFFARX1 I_32022 (I546885,I2507,I546427,I546398,);
nand I_32023 (I546916,I546877,I546518);
nand I_32024 (I546933,I546611,I546916);
nor I_32025 (I546407,I546933,I546577);
not I_32026 (I546988,I2514);
DFFARX1 I_32027 (I395220,I2507,I546988,I547014,);
DFFARX1 I_32028 (I547014,I2507,I546988,I547031,);
not I_32029 (I546980,I547031);
not I_32030 (I547053,I547014);
DFFARX1 I_32031 (I395232,I2507,I546988,I547079,);
nand I_32032 (I547087,I547079,I395241);
not I_32033 (I547104,I395241);
not I_32034 (I547121,I395223);
nand I_32035 (I547138,I395226,I395217);
and I_32036 (I547155,I395226,I395217);
not I_32037 (I547172,I395235);
nand I_32038 (I547189,I547172,I547121);
nor I_32039 (I546962,I547189,I547087);
nor I_32040 (I547220,I547104,I547189);
nand I_32041 (I546965,I547155,I547220);
not I_32042 (I547251,I395238);
nor I_32043 (I547268,I547251,I395226);
nor I_32044 (I547285,I547268,I395235);
nor I_32045 (I547302,I547053,I547285);
DFFARX1 I_32046 (I547302,I2507,I546988,I546974,);
not I_32047 (I547333,I547268);
DFFARX1 I_32048 (I547333,I2507,I546988,I546977,);
and I_32049 (I546971,I547079,I547268);
nor I_32050 (I547378,I547251,I395217);
and I_32051 (I547395,I547378,I395229);
or I_32052 (I547412,I547395,I395220);
DFFARX1 I_32053 (I547412,I2507,I546988,I547438,);
nor I_32054 (I547446,I547438,I547172);
DFFARX1 I_32055 (I547446,I2507,I546988,I546959,);
nand I_32056 (I547477,I547438,I547079);
nand I_32057 (I547494,I547172,I547477);
nor I_32058 (I546968,I547494,I547138);
not I_32059 (I547549,I2514);
DFFARX1 I_32060 (I491216,I2507,I547549,I547575,);
DFFARX1 I_32061 (I547575,I2507,I547549,I547592,);
not I_32062 (I547541,I547592);
not I_32063 (I547614,I547575);
DFFARX1 I_32064 (I491243,I2507,I547549,I547640,);
nand I_32065 (I547648,I547640,I491234);
not I_32066 (I547665,I491234);
not I_32067 (I547682,I491216);
nand I_32068 (I547699,I491228,I491231);
and I_32069 (I547716,I491228,I491231);
not I_32070 (I547733,I491240);
nand I_32071 (I547750,I547733,I547682);
nor I_32072 (I547523,I547750,I547648);
nor I_32073 (I547781,I547665,I547750);
nand I_32074 (I547526,I547716,I547781);
not I_32075 (I547812,I491225);
nor I_32076 (I547829,I547812,I491228);
nor I_32077 (I547846,I547829,I491240);
nor I_32078 (I547863,I547614,I547846);
DFFARX1 I_32079 (I547863,I2507,I547549,I547535,);
not I_32080 (I547894,I547829);
DFFARX1 I_32081 (I547894,I2507,I547549,I547538,);
and I_32082 (I547532,I547640,I547829);
nor I_32083 (I547939,I547812,I491219);
and I_32084 (I547956,I547939,I491222);
or I_32085 (I547973,I547956,I491237);
DFFARX1 I_32086 (I547973,I2507,I547549,I547999,);
nor I_32087 (I548007,I547999,I547733);
DFFARX1 I_32088 (I548007,I2507,I547549,I547520,);
nand I_32089 (I548038,I547999,I547640);
nand I_32090 (I548055,I547733,I548038);
nor I_32091 (I547529,I548055,I547699);
not I_32092 (I548110,I2514);
DFFARX1 I_32093 (I29361,I2507,I548110,I548136,);
DFFARX1 I_32094 (I548136,I2507,I548110,I548153,);
not I_32095 (I548102,I548153);
not I_32096 (I548175,I548136);
DFFARX1 I_32097 (I29346,I2507,I548110,I548201,);
nand I_32098 (I548209,I548201,I29358);
not I_32099 (I548226,I29358);
not I_32100 (I548243,I29364);
nand I_32101 (I548260,I29352,I29343);
and I_32102 (I548277,I29352,I29343);
not I_32103 (I548294,I29349);
nand I_32104 (I548311,I548294,I548243);
nor I_32105 (I548084,I548311,I548209);
nor I_32106 (I548342,I548226,I548311);
nand I_32107 (I548087,I548277,I548342);
not I_32108 (I548373,I29355);
nor I_32109 (I548390,I548373,I29352);
nor I_32110 (I548407,I548390,I29349);
nor I_32111 (I548424,I548175,I548407);
DFFARX1 I_32112 (I548424,I2507,I548110,I548096,);
not I_32113 (I548455,I548390);
DFFARX1 I_32114 (I548455,I2507,I548110,I548099,);
and I_32115 (I548093,I548201,I548390);
nor I_32116 (I548500,I548373,I29343);
and I_32117 (I548517,I548500,I29367);
or I_32118 (I548534,I548517,I29346);
DFFARX1 I_32119 (I548534,I2507,I548110,I548560,);
nor I_32120 (I548568,I548560,I548294);
DFFARX1 I_32121 (I548568,I2507,I548110,I548081,);
nand I_32122 (I548599,I548560,I548201);
nand I_32123 (I548616,I548294,I548599);
nor I_32124 (I548090,I548616,I548260);
not I_32125 (I548671,I2514);
DFFARX1 I_32126 (I256912,I2507,I548671,I548697,);
DFFARX1 I_32127 (I548697,I2507,I548671,I548714,);
not I_32128 (I548663,I548714);
not I_32129 (I548736,I548697);
DFFARX1 I_32130 (I256900,I2507,I548671,I548762,);
nand I_32131 (I548770,I548762,I256906);
not I_32132 (I548787,I256906);
not I_32133 (I548804,I256903);
nand I_32134 (I548821,I256891,I256888);
and I_32135 (I548838,I256891,I256888);
not I_32136 (I548855,I256915);
nand I_32137 (I548872,I548855,I548804);
nor I_32138 (I548645,I548872,I548770);
nor I_32139 (I548903,I548787,I548872);
nand I_32140 (I548648,I548838,I548903);
not I_32141 (I548934,I256888);
nor I_32142 (I548951,I548934,I256891);
nor I_32143 (I548968,I548951,I256915);
nor I_32144 (I548985,I548736,I548968);
DFFARX1 I_32145 (I548985,I2507,I548671,I548657,);
not I_32146 (I549016,I548951);
DFFARX1 I_32147 (I549016,I2507,I548671,I548660,);
and I_32148 (I548654,I548762,I548951);
nor I_32149 (I549061,I548934,I256897);
and I_32150 (I549078,I549061,I256894);
or I_32151 (I549095,I549078,I256909);
DFFARX1 I_32152 (I549095,I2507,I548671,I549121,);
nor I_32153 (I549129,I549121,I548855);
DFFARX1 I_32154 (I549129,I2507,I548671,I548642,);
nand I_32155 (I549160,I549121,I548762);
nand I_32156 (I549177,I548855,I549160);
nor I_32157 (I548651,I549177,I548821);
not I_32158 (I549232,I2514);
DFFARX1 I_32159 (I672286,I2507,I549232,I549258,);
DFFARX1 I_32160 (I549258,I2507,I549232,I549275,);
not I_32161 (I549224,I549275);
not I_32162 (I549297,I549258);
DFFARX1 I_32163 (I672283,I2507,I549232,I549323,);
nand I_32164 (I549331,I549323,I672289);
not I_32165 (I549348,I672289);
not I_32166 (I549365,I672298);
nand I_32167 (I549382,I672292,I672286);
and I_32168 (I549399,I672292,I672286);
not I_32169 (I549416,I672304);
nand I_32170 (I549433,I549416,I549365);
nor I_32171 (I549206,I549433,I549331);
nor I_32172 (I549464,I549348,I549433);
nand I_32173 (I549209,I549399,I549464);
not I_32174 (I549495,I672301);
nor I_32175 (I549512,I549495,I672292);
nor I_32176 (I549529,I549512,I672304);
nor I_32177 (I549546,I549297,I549529);
DFFARX1 I_32178 (I549546,I2507,I549232,I549218,);
not I_32179 (I549577,I549512);
DFFARX1 I_32180 (I549577,I2507,I549232,I549221,);
and I_32181 (I549215,I549323,I549512);
nor I_32182 (I549622,I549495,I672295);
and I_32183 (I549639,I549622,I672307);
or I_32184 (I549656,I549639,I672283);
DFFARX1 I_32185 (I549656,I2507,I549232,I549682,);
nor I_32186 (I549690,I549682,I549416);
DFFARX1 I_32187 (I549690,I2507,I549232,I549203,);
nand I_32188 (I549721,I549682,I549323);
nand I_32189 (I549738,I549416,I549721);
nor I_32190 (I549212,I549738,I549382);
not I_32191 (I549793,I2514);
DFFARX1 I_32192 (I37787,I2507,I549793,I549819,);
DFFARX1 I_32193 (I549819,I2507,I549793,I549836,);
not I_32194 (I549785,I549836);
not I_32195 (I549858,I549819);
DFFARX1 I_32196 (I37775,I2507,I549793,I549884,);
nand I_32197 (I549892,I549884,I37790);
not I_32198 (I549909,I37790);
not I_32199 (I549926,I37778);
nand I_32200 (I549943,I37799,I37793);
and I_32201 (I549960,I37799,I37793);
not I_32202 (I549977,I37781);
nand I_32203 (I549994,I549977,I549926);
nor I_32204 (I549767,I549994,I549892);
nor I_32205 (I550025,I549909,I549994);
nand I_32206 (I549770,I549960,I550025);
not I_32207 (I550056,I37784);
nor I_32208 (I550073,I550056,I37799);
nor I_32209 (I550090,I550073,I37781);
nor I_32210 (I550107,I549858,I550090);
DFFARX1 I_32211 (I550107,I2507,I549793,I549779,);
not I_32212 (I550138,I550073);
DFFARX1 I_32213 (I550138,I2507,I549793,I549782,);
and I_32214 (I549776,I549884,I550073);
nor I_32215 (I550183,I550056,I37778);
and I_32216 (I550200,I550183,I37775);
or I_32217 (I550217,I550200,I37796);
DFFARX1 I_32218 (I550217,I2507,I549793,I550243,);
nor I_32219 (I550251,I550243,I549977);
DFFARX1 I_32220 (I550251,I2507,I549793,I549764,);
nand I_32221 (I550282,I550243,I549884);
nand I_32222 (I550299,I549977,I550282);
nor I_32223 (I549773,I550299,I549943);
not I_32224 (I550354,I2514);
DFFARX1 I_32225 (I518348,I2507,I550354,I550380,);
DFFARX1 I_32226 (I550380,I2507,I550354,I550397,);
not I_32227 (I550346,I550397);
not I_32228 (I550419,I550380);
DFFARX1 I_32229 (I518375,I2507,I550354,I550445,);
nand I_32230 (I550453,I550445,I518366);
not I_32231 (I550470,I518366);
not I_32232 (I550487,I518348);
nand I_32233 (I550504,I518360,I518363);
and I_32234 (I550521,I518360,I518363);
not I_32235 (I550538,I518372);
nand I_32236 (I550555,I550538,I550487);
nor I_32237 (I550328,I550555,I550453);
nor I_32238 (I550586,I550470,I550555);
nand I_32239 (I550331,I550521,I550586);
not I_32240 (I550617,I518357);
nor I_32241 (I550634,I550617,I518360);
nor I_32242 (I550651,I550634,I518372);
nor I_32243 (I550668,I550419,I550651);
DFFARX1 I_32244 (I550668,I2507,I550354,I550340,);
not I_32245 (I550699,I550634);
DFFARX1 I_32246 (I550699,I2507,I550354,I550343,);
and I_32247 (I550337,I550445,I550634);
nor I_32248 (I550744,I550617,I518351);
and I_32249 (I550761,I550744,I518354);
or I_32250 (I550778,I550761,I518369);
DFFARX1 I_32251 (I550778,I2507,I550354,I550804,);
nor I_32252 (I550812,I550804,I550538);
DFFARX1 I_32253 (I550812,I2507,I550354,I550325,);
nand I_32254 (I550843,I550804,I550445);
nand I_32255 (I550860,I550538,I550843);
nor I_32256 (I550334,I550860,I550504);
not I_32257 (I550915,I2514);
DFFARX1 I_32258 (I15132,I2507,I550915,I550941,);
DFFARX1 I_32259 (I550941,I2507,I550915,I550958,);
not I_32260 (I550907,I550958);
not I_32261 (I550980,I550941);
DFFARX1 I_32262 (I15117,I2507,I550915,I551006,);
nand I_32263 (I551014,I551006,I15129);
not I_32264 (I551031,I15129);
not I_32265 (I551048,I15135);
nand I_32266 (I551065,I15123,I15114);
and I_32267 (I551082,I15123,I15114);
not I_32268 (I551099,I15120);
nand I_32269 (I551116,I551099,I551048);
nor I_32270 (I550889,I551116,I551014);
nor I_32271 (I551147,I551031,I551116);
nand I_32272 (I550892,I551082,I551147);
not I_32273 (I551178,I15126);
nor I_32274 (I551195,I551178,I15123);
nor I_32275 (I551212,I551195,I15120);
nor I_32276 (I551229,I550980,I551212);
DFFARX1 I_32277 (I551229,I2507,I550915,I550901,);
not I_32278 (I551260,I551195);
DFFARX1 I_32279 (I551260,I2507,I550915,I550904,);
and I_32280 (I550898,I551006,I551195);
nor I_32281 (I551305,I551178,I15114);
and I_32282 (I551322,I551305,I15138);
or I_32283 (I551339,I551322,I15117);
DFFARX1 I_32284 (I551339,I2507,I550915,I551365,);
nor I_32285 (I551373,I551365,I551099);
DFFARX1 I_32286 (I551373,I2507,I550915,I550886,);
nand I_32287 (I551404,I551365,I551006);
nand I_32288 (I551421,I551099,I551404);
nor I_32289 (I550895,I551421,I551065);
not I_32290 (I551476,I2514);
DFFARX1 I_32291 (I505428,I2507,I551476,I551502,);
DFFARX1 I_32292 (I551502,I2507,I551476,I551519,);
not I_32293 (I551468,I551519);
not I_32294 (I551541,I551502);
DFFARX1 I_32295 (I505455,I2507,I551476,I551567,);
nand I_32296 (I551575,I551567,I505446);
not I_32297 (I551592,I505446);
not I_32298 (I551609,I505428);
nand I_32299 (I551626,I505440,I505443);
and I_32300 (I551643,I505440,I505443);
not I_32301 (I551660,I505452);
nand I_32302 (I551677,I551660,I551609);
nor I_32303 (I551450,I551677,I551575);
nor I_32304 (I551708,I551592,I551677);
nand I_32305 (I551453,I551643,I551708);
not I_32306 (I551739,I505437);
nor I_32307 (I551756,I551739,I505440);
nor I_32308 (I551773,I551756,I505452);
nor I_32309 (I551790,I551541,I551773);
DFFARX1 I_32310 (I551790,I2507,I551476,I551462,);
not I_32311 (I551821,I551756);
DFFARX1 I_32312 (I551821,I2507,I551476,I551465,);
and I_32313 (I551459,I551567,I551756);
nor I_32314 (I551866,I551739,I505431);
and I_32315 (I551883,I551866,I505434);
or I_32316 (I551900,I551883,I505449);
DFFARX1 I_32317 (I551900,I2507,I551476,I551926,);
nor I_32318 (I551934,I551926,I551660);
DFFARX1 I_32319 (I551934,I2507,I551476,I551447,);
nand I_32320 (I551965,I551926,I551567);
nand I_32321 (I551982,I551660,I551965);
nor I_32322 (I551456,I551982,I551626);
not I_32323 (I552037,I2514);
DFFARX1 I_32324 (I627180,I2507,I552037,I552063,);
DFFARX1 I_32325 (I552063,I2507,I552037,I552080,);
not I_32326 (I552029,I552080);
not I_32327 (I552102,I552063);
DFFARX1 I_32328 (I627171,I2507,I552037,I552128,);
nand I_32329 (I552136,I552128,I627168);
not I_32330 (I552153,I627168);
not I_32331 (I552170,I627177);
nand I_32332 (I552187,I627186,I627168);
and I_32333 (I552204,I627186,I627168);
not I_32334 (I552221,I627165);
nand I_32335 (I552238,I552221,I552170);
nor I_32336 (I552011,I552238,I552136);
nor I_32337 (I552269,I552153,I552238);
nand I_32338 (I552014,I552204,I552269);
not I_32339 (I552300,I627174);
nor I_32340 (I552317,I552300,I627186);
nor I_32341 (I552334,I552317,I627165);
nor I_32342 (I552351,I552102,I552334);
DFFARX1 I_32343 (I552351,I2507,I552037,I552023,);
not I_32344 (I552382,I552317);
DFFARX1 I_32345 (I552382,I2507,I552037,I552026,);
and I_32346 (I552020,I552128,I552317);
nor I_32347 (I552427,I552300,I627189);
and I_32348 (I552444,I552427,I627165);
or I_32349 (I552461,I552444,I627183);
DFFARX1 I_32350 (I552461,I2507,I552037,I552487,);
nor I_32351 (I552495,I552487,I552221);
DFFARX1 I_32352 (I552495,I2507,I552037,I552008,);
nand I_32353 (I552526,I552487,I552128);
nand I_32354 (I552543,I552221,I552526);
nor I_32355 (I552017,I552543,I552187);
not I_32356 (I552598,I2514);
DFFARX1 I_32357 (I502844,I2507,I552598,I552624,);
DFFARX1 I_32358 (I552624,I2507,I552598,I552641,);
not I_32359 (I552590,I552641);
not I_32360 (I552663,I552624);
DFFARX1 I_32361 (I502871,I2507,I552598,I552689,);
nand I_32362 (I552697,I552689,I502862);
not I_32363 (I552714,I502862);
not I_32364 (I552731,I502844);
nand I_32365 (I552748,I502856,I502859);
and I_32366 (I552765,I502856,I502859);
not I_32367 (I552782,I502868);
nand I_32368 (I552799,I552782,I552731);
nor I_32369 (I552572,I552799,I552697);
nor I_32370 (I552830,I552714,I552799);
nand I_32371 (I552575,I552765,I552830);
not I_32372 (I552861,I502853);
nor I_32373 (I552878,I552861,I502856);
nor I_32374 (I552895,I552878,I502868);
nor I_32375 (I552912,I552663,I552895);
DFFARX1 I_32376 (I552912,I2507,I552598,I552584,);
not I_32377 (I552943,I552878);
DFFARX1 I_32378 (I552943,I2507,I552598,I552587,);
and I_32379 (I552581,I552689,I552878);
nor I_32380 (I552988,I552861,I502847);
and I_32381 (I553005,I552988,I502850);
or I_32382 (I553022,I553005,I502865);
DFFARX1 I_32383 (I553022,I2507,I552598,I553048,);
nor I_32384 (I553056,I553048,I552782);
DFFARX1 I_32385 (I553056,I2507,I552598,I552569,);
nand I_32386 (I553087,I553048,I552689);
nand I_32387 (I553104,I552782,I553087);
nor I_32388 (I552578,I553104,I552748);
not I_32389 (I553159,I2514);
DFFARX1 I_32390 (I526746,I2507,I553159,I553185,);
DFFARX1 I_32391 (I553185,I2507,I553159,I553202,);
not I_32392 (I553151,I553202);
not I_32393 (I553224,I553185);
DFFARX1 I_32394 (I526773,I2507,I553159,I553250,);
nand I_32395 (I553258,I553250,I526764);
not I_32396 (I553275,I526764);
not I_32397 (I553292,I526746);
nand I_32398 (I553309,I526758,I526761);
and I_32399 (I553326,I526758,I526761);
not I_32400 (I553343,I526770);
nand I_32401 (I553360,I553343,I553292);
nor I_32402 (I553133,I553360,I553258);
nor I_32403 (I553391,I553275,I553360);
nand I_32404 (I553136,I553326,I553391);
not I_32405 (I553422,I526755);
nor I_32406 (I553439,I553422,I526758);
nor I_32407 (I553456,I553439,I526770);
nor I_32408 (I553473,I553224,I553456);
DFFARX1 I_32409 (I553473,I2507,I553159,I553145,);
not I_32410 (I553504,I553439);
DFFARX1 I_32411 (I553504,I2507,I553159,I553148,);
and I_32412 (I553142,I553250,I553439);
nor I_32413 (I553549,I553422,I526749);
and I_32414 (I553566,I553549,I526752);
or I_32415 (I553583,I553566,I526767);
DFFARX1 I_32416 (I553583,I2507,I553159,I553609,);
nor I_32417 (I553617,I553609,I553343);
DFFARX1 I_32418 (I553617,I2507,I553159,I553130,);
nand I_32419 (I553648,I553609,I553250);
nand I_32420 (I553665,I553343,I553648);
nor I_32421 (I553139,I553665,I553309);
not I_32422 (I553720,I2514);
DFFARX1 I_32423 (I177995,I2507,I553720,I553746,);
DFFARX1 I_32424 (I553746,I2507,I553720,I553763,);
not I_32425 (I553712,I553763);
not I_32426 (I553785,I553746);
DFFARX1 I_32427 (I177992,I2507,I553720,I553811,);
nand I_32428 (I553819,I553811,I177986);
not I_32429 (I553836,I177986);
not I_32430 (I553853,I177983);
nand I_32431 (I553870,I177977,I177974);
and I_32432 (I553887,I177977,I177974);
not I_32433 (I553904,I177989);
nand I_32434 (I553921,I553904,I553853);
nor I_32435 (I553694,I553921,I553819);
nor I_32436 (I553952,I553836,I553921);
nand I_32437 (I553697,I553887,I553952);
not I_32438 (I553983,I178001);
nor I_32439 (I554000,I553983,I177977);
nor I_32440 (I554017,I554000,I177989);
nor I_32441 (I554034,I553785,I554017);
DFFARX1 I_32442 (I554034,I2507,I553720,I553706,);
not I_32443 (I554065,I554000);
DFFARX1 I_32444 (I554065,I2507,I553720,I553709,);
and I_32445 (I553703,I553811,I554000);
nor I_32446 (I554110,I553983,I177998);
and I_32447 (I554127,I554110,I177974);
or I_32448 (I554144,I554127,I177980);
DFFARX1 I_32449 (I554144,I2507,I553720,I554170,);
nor I_32450 (I554178,I554170,I553904);
DFFARX1 I_32451 (I554178,I2507,I553720,I553691,);
nand I_32452 (I554209,I554170,I553811);
nand I_32453 (I554226,I553904,I554209);
nor I_32454 (I553700,I554226,I553870);
not I_32455 (I554281,I2514);
DFFARX1 I_32456 (I77839,I2507,I554281,I554307,);
DFFARX1 I_32457 (I554307,I2507,I554281,I554324,);
not I_32458 (I554273,I554324);
not I_32459 (I554346,I554307);
DFFARX1 I_32460 (I77827,I2507,I554281,I554372,);
nand I_32461 (I554380,I554372,I77842);
not I_32462 (I554397,I77842);
not I_32463 (I554414,I77830);
nand I_32464 (I554431,I77851,I77845);
and I_32465 (I554448,I77851,I77845);
not I_32466 (I554465,I77833);
nand I_32467 (I554482,I554465,I554414);
nor I_32468 (I554255,I554482,I554380);
nor I_32469 (I554513,I554397,I554482);
nand I_32470 (I554258,I554448,I554513);
not I_32471 (I554544,I77836);
nor I_32472 (I554561,I554544,I77851);
nor I_32473 (I554578,I554561,I77833);
nor I_32474 (I554595,I554346,I554578);
DFFARX1 I_32475 (I554595,I2507,I554281,I554267,);
not I_32476 (I554626,I554561);
DFFARX1 I_32477 (I554626,I2507,I554281,I554270,);
and I_32478 (I554264,I554372,I554561);
nor I_32479 (I554671,I554544,I77830);
and I_32480 (I554688,I554671,I77827);
or I_32481 (I554705,I554688,I77848);
DFFARX1 I_32482 (I554705,I2507,I554281,I554731,);
nor I_32483 (I554739,I554731,I554465);
DFFARX1 I_32484 (I554739,I2507,I554281,I554252,);
nand I_32485 (I554770,I554731,I554372);
nand I_32486 (I554787,I554465,I554770);
nor I_32487 (I554261,I554787,I554431);
not I_32488 (I554842,I2514);
DFFARX1 I_32489 (I672864,I2507,I554842,I554868,);
DFFARX1 I_32490 (I554868,I2507,I554842,I554885,);
not I_32491 (I554834,I554885);
not I_32492 (I554907,I554868);
DFFARX1 I_32493 (I672861,I2507,I554842,I554933,);
nand I_32494 (I554941,I554933,I672867);
not I_32495 (I554958,I672867);
not I_32496 (I554975,I672876);
nand I_32497 (I554992,I672870,I672864);
and I_32498 (I555009,I672870,I672864);
not I_32499 (I555026,I672882);
nand I_32500 (I555043,I555026,I554975);
nor I_32501 (I554816,I555043,I554941);
nor I_32502 (I555074,I554958,I555043);
nand I_32503 (I554819,I555009,I555074);
not I_32504 (I555105,I672879);
nor I_32505 (I555122,I555105,I672870);
nor I_32506 (I555139,I555122,I672882);
nor I_32507 (I555156,I554907,I555139);
DFFARX1 I_32508 (I555156,I2507,I554842,I554828,);
not I_32509 (I555187,I555122);
DFFARX1 I_32510 (I555187,I2507,I554842,I554831,);
and I_32511 (I554825,I554933,I555122);
nor I_32512 (I555232,I555105,I672873);
and I_32513 (I555249,I555232,I672885);
or I_32514 (I555266,I555249,I672861);
DFFARX1 I_32515 (I555266,I2507,I554842,I555292,);
nor I_32516 (I555300,I555292,I555026);
DFFARX1 I_32517 (I555300,I2507,I554842,I554813,);
nand I_32518 (I555331,I555292,I554933);
nand I_32519 (I555348,I555026,I555331);
nor I_32520 (I554822,I555348,I554992);
not I_32521 (I555403,I2514);
DFFARX1 I_32522 (I606950,I2507,I555403,I555429,);
DFFARX1 I_32523 (I555429,I2507,I555403,I555446,);
not I_32524 (I555395,I555446);
not I_32525 (I555468,I555429);
DFFARX1 I_32526 (I606941,I2507,I555403,I555494,);
nand I_32527 (I555502,I555494,I606938);
not I_32528 (I555519,I606938);
not I_32529 (I555536,I606947);
nand I_32530 (I555553,I606956,I606938);
and I_32531 (I555570,I606956,I606938);
not I_32532 (I555587,I606935);
nand I_32533 (I555604,I555587,I555536);
nor I_32534 (I555377,I555604,I555502);
nor I_32535 (I555635,I555519,I555604);
nand I_32536 (I555380,I555570,I555635);
not I_32537 (I555666,I606944);
nor I_32538 (I555683,I555666,I606956);
nor I_32539 (I555700,I555683,I606935);
nor I_32540 (I555717,I555468,I555700);
DFFARX1 I_32541 (I555717,I2507,I555403,I555389,);
not I_32542 (I555748,I555683);
DFFARX1 I_32543 (I555748,I2507,I555403,I555392,);
and I_32544 (I555386,I555494,I555683);
nor I_32545 (I555793,I555666,I606959);
and I_32546 (I555810,I555793,I606935);
or I_32547 (I555827,I555810,I606953);
DFFARX1 I_32548 (I555827,I2507,I555403,I555853,);
nor I_32549 (I555861,I555853,I555587);
DFFARX1 I_32550 (I555861,I2507,I555403,I555374,);
nand I_32551 (I555892,I555853,I555494);
nand I_32552 (I555909,I555587,I555892);
nor I_32553 (I555383,I555909,I555553);
not I_32554 (I555964,I2514);
DFFARX1 I_32555 (I640363,I2507,I555964,I555990,);
DFFARX1 I_32556 (I555990,I2507,I555964,I556007,);
not I_32557 (I555956,I556007);
not I_32558 (I556029,I555990);
DFFARX1 I_32559 (I640369,I2507,I555964,I556055,);
nand I_32560 (I556063,I556055,I640378);
not I_32561 (I556080,I640378);
not I_32562 (I556097,I640357);
nand I_32563 (I556114,I640360,I640360);
and I_32564 (I556131,I640360,I640360);
not I_32565 (I556148,I640372);
nand I_32566 (I556165,I556148,I556097);
nor I_32567 (I555938,I556165,I556063);
nor I_32568 (I556196,I556080,I556165);
nand I_32569 (I555941,I556131,I556196);
not I_32570 (I556227,I640366);
nor I_32571 (I556244,I556227,I640360);
nor I_32572 (I556261,I556244,I640372);
nor I_32573 (I556278,I556029,I556261);
DFFARX1 I_32574 (I556278,I2507,I555964,I555950,);
not I_32575 (I556309,I556244);
DFFARX1 I_32576 (I556309,I2507,I555964,I555953,);
and I_32577 (I555947,I556055,I556244);
nor I_32578 (I556354,I556227,I640381);
and I_32579 (I556371,I556354,I640357);
or I_32580 (I556388,I556371,I640375);
DFFARX1 I_32581 (I556388,I2507,I555964,I556414,);
nor I_32582 (I556422,I556414,I556148);
DFFARX1 I_32583 (I556422,I2507,I555964,I555935,);
nand I_32584 (I556453,I556414,I556055);
nand I_32585 (I556470,I556148,I556453);
nor I_32586 (I555944,I556470,I556114);
not I_32587 (I556525,I2514);
DFFARX1 I_32588 (I109807,I2507,I556525,I556551,);
DFFARX1 I_32589 (I556551,I2507,I556525,I556568,);
not I_32590 (I556517,I556568);
not I_32591 (I556590,I556551);
DFFARX1 I_32592 (I109822,I2507,I556525,I556616,);
nand I_32593 (I556624,I556616,I109804);
not I_32594 (I556641,I109804);
not I_32595 (I556658,I109813);
nand I_32596 (I556675,I109819,I109810);
and I_32597 (I556692,I109819,I109810);
not I_32598 (I556709,I109807);
nand I_32599 (I556726,I556709,I556658);
nor I_32600 (I556499,I556726,I556624);
nor I_32601 (I556757,I556641,I556726);
nand I_32602 (I556502,I556692,I556757);
not I_32603 (I556788,I109804);
nor I_32604 (I556805,I556788,I109819);
nor I_32605 (I556822,I556805,I109807);
nor I_32606 (I556839,I556590,I556822);
DFFARX1 I_32607 (I556839,I2507,I556525,I556511,);
not I_32608 (I556870,I556805);
DFFARX1 I_32609 (I556870,I2507,I556525,I556514,);
and I_32610 (I556508,I556616,I556805);
nor I_32611 (I556915,I556788,I109828);
and I_32612 (I556932,I556915,I109825);
or I_32613 (I556949,I556932,I109816);
DFFARX1 I_32614 (I556949,I2507,I556525,I556975,);
nor I_32615 (I556983,I556975,I556709);
DFFARX1 I_32616 (I556983,I2507,I556525,I556496,);
nand I_32617 (I557014,I556975,I556616);
nand I_32618 (I557031,I556709,I557014);
nor I_32619 (I556505,I557031,I556675);
not I_32620 (I557086,I2514);
DFFARX1 I_32621 (I327013,I2507,I557086,I557112,);
DFFARX1 I_32622 (I557112,I2507,I557086,I557129,);
not I_32623 (I557078,I557129);
not I_32624 (I557151,I557112);
DFFARX1 I_32625 (I327028,I2507,I557086,I557177,);
nand I_32626 (I557185,I557177,I327019);
not I_32627 (I557202,I327019);
not I_32628 (I557219,I327025);
nand I_32629 (I557236,I327022,I327031);
and I_32630 (I557253,I327022,I327031);
not I_32631 (I557270,I327016);
nand I_32632 (I557287,I557270,I557219);
nor I_32633 (I557060,I557287,I557185);
nor I_32634 (I557318,I557202,I557287);
nand I_32635 (I557063,I557253,I557318);
not I_32636 (I557349,I327013);
nor I_32637 (I557366,I557349,I327022);
nor I_32638 (I557383,I557366,I327016);
nor I_32639 (I557400,I557151,I557383);
DFFARX1 I_32640 (I557400,I2507,I557086,I557072,);
not I_32641 (I557431,I557366);
DFFARX1 I_32642 (I557431,I2507,I557086,I557075,);
and I_32643 (I557069,I557177,I557366);
nor I_32644 (I557476,I557349,I327037);
and I_32645 (I557493,I557476,I327016);
or I_32646 (I557510,I557493,I327034);
DFFARX1 I_32647 (I557510,I2507,I557086,I557536,);
nor I_32648 (I557544,I557536,I557270);
DFFARX1 I_32649 (I557544,I2507,I557086,I557057,);
nand I_32650 (I557575,I557536,I557177);
nand I_32651 (I557592,I557270,I557575);
nor I_32652 (I557066,I557592,I557236);
not I_32653 (I557647,I2514);
DFFARX1 I_32654 (I158002,I2507,I557647,I557673,);
DFFARX1 I_32655 (I557673,I2507,I557647,I557690,);
not I_32656 (I557639,I557690);
not I_32657 (I557712,I557673);
DFFARX1 I_32658 (I158017,I2507,I557647,I557738,);
nand I_32659 (I557746,I557738,I157999);
not I_32660 (I557763,I157999);
not I_32661 (I557780,I158008);
nand I_32662 (I557797,I158014,I158005);
and I_32663 (I557814,I158014,I158005);
not I_32664 (I557831,I158002);
nand I_32665 (I557848,I557831,I557780);
nor I_32666 (I557621,I557848,I557746);
nor I_32667 (I557879,I557763,I557848);
nand I_32668 (I557624,I557814,I557879);
not I_32669 (I557910,I157999);
nor I_32670 (I557927,I557910,I158014);
nor I_32671 (I557944,I557927,I158002);
nor I_32672 (I557961,I557712,I557944);
DFFARX1 I_32673 (I557961,I2507,I557647,I557633,);
not I_32674 (I557992,I557927);
DFFARX1 I_32675 (I557992,I2507,I557647,I557636,);
and I_32676 (I557630,I557738,I557927);
nor I_32677 (I558037,I557910,I158023);
and I_32678 (I558054,I558037,I158020);
or I_32679 (I558071,I558054,I158011);
DFFARX1 I_32680 (I558071,I2507,I557647,I558097,);
nor I_32681 (I558105,I558097,I557831);
DFFARX1 I_32682 (I558105,I2507,I557647,I557618,);
nand I_32683 (I558136,I558097,I557738);
nand I_32684 (I558153,I557831,I558136);
nor I_32685 (I557627,I558153,I557797);
not I_32686 (I558208,I2514);
DFFARX1 I_32687 (I504136,I2507,I558208,I558234,);
DFFARX1 I_32688 (I558234,I2507,I558208,I558251,);
not I_32689 (I558200,I558251);
not I_32690 (I558273,I558234);
DFFARX1 I_32691 (I504163,I2507,I558208,I558299,);
nand I_32692 (I558307,I558299,I504154);
not I_32693 (I558324,I504154);
not I_32694 (I558341,I504136);
nand I_32695 (I558358,I504148,I504151);
and I_32696 (I558375,I504148,I504151);
not I_32697 (I558392,I504160);
nand I_32698 (I558409,I558392,I558341);
nor I_32699 (I558182,I558409,I558307);
nor I_32700 (I558440,I558324,I558409);
nand I_32701 (I558185,I558375,I558440);
not I_32702 (I558471,I504145);
nor I_32703 (I558488,I558471,I504148);
nor I_32704 (I558505,I558488,I504160);
nor I_32705 (I558522,I558273,I558505);
DFFARX1 I_32706 (I558522,I2507,I558208,I558194,);
not I_32707 (I558553,I558488);
DFFARX1 I_32708 (I558553,I2507,I558208,I558197,);
and I_32709 (I558191,I558299,I558488);
nor I_32710 (I558598,I558471,I504139);
and I_32711 (I558615,I558598,I504142);
or I_32712 (I558632,I558615,I504157);
DFFARX1 I_32713 (I558632,I2507,I558208,I558658,);
nor I_32714 (I558666,I558658,I558392);
DFFARX1 I_32715 (I558666,I2507,I558208,I558179,);
nand I_32716 (I558697,I558658,I558299);
nand I_32717 (I558714,I558392,I558697);
nor I_32718 (I558188,I558714,I558358);
not I_32719 (I558769,I2514);
DFFARX1 I_32720 (I174306,I2507,I558769,I558795,);
DFFARX1 I_32721 (I558795,I2507,I558769,I558812,);
not I_32722 (I558761,I558812);
not I_32723 (I558834,I558795);
DFFARX1 I_32724 (I174303,I2507,I558769,I558860,);
nand I_32725 (I558868,I558860,I174297);
not I_32726 (I558885,I174297);
not I_32727 (I558902,I174294);
nand I_32728 (I558919,I174288,I174285);
and I_32729 (I558936,I174288,I174285);
not I_32730 (I558953,I174300);
nand I_32731 (I558970,I558953,I558902);
nor I_32732 (I558743,I558970,I558868);
nor I_32733 (I559001,I558885,I558970);
nand I_32734 (I558746,I558936,I559001);
not I_32735 (I559032,I174312);
nor I_32736 (I559049,I559032,I174288);
nor I_32737 (I559066,I559049,I174300);
nor I_32738 (I559083,I558834,I559066);
DFFARX1 I_32739 (I559083,I2507,I558769,I558755,);
not I_32740 (I559114,I559049);
DFFARX1 I_32741 (I559114,I2507,I558769,I558758,);
and I_32742 (I558752,I558860,I559049);
nor I_32743 (I559159,I559032,I174309);
and I_32744 (I559176,I559159,I174285);
or I_32745 (I559193,I559176,I174291);
DFFARX1 I_32746 (I559193,I2507,I558769,I559219,);
nor I_32747 (I559227,I559219,I558953);
DFFARX1 I_32748 (I559227,I2507,I558769,I558740,);
nand I_32749 (I559258,I559219,I558860);
nand I_32750 (I559275,I558953,I559258);
nor I_32751 (I558749,I559275,I558919);
not I_32752 (I559330,I2514);
DFFARX1 I_32753 (I42003,I2507,I559330,I559356,);
DFFARX1 I_32754 (I559356,I2507,I559330,I559373,);
not I_32755 (I559322,I559373);
not I_32756 (I559395,I559356);
DFFARX1 I_32757 (I41991,I2507,I559330,I559421,);
nand I_32758 (I559429,I559421,I42006);
not I_32759 (I559446,I42006);
not I_32760 (I559463,I41994);
nand I_32761 (I559480,I42015,I42009);
and I_32762 (I559497,I42015,I42009);
not I_32763 (I559514,I41997);
nand I_32764 (I559531,I559514,I559463);
nor I_32765 (I559304,I559531,I559429);
nor I_32766 (I559562,I559446,I559531);
nand I_32767 (I559307,I559497,I559562);
not I_32768 (I559593,I42000);
nor I_32769 (I559610,I559593,I42015);
nor I_32770 (I559627,I559610,I41997);
nor I_32771 (I559644,I559395,I559627);
DFFARX1 I_32772 (I559644,I2507,I559330,I559316,);
not I_32773 (I559675,I559610);
DFFARX1 I_32774 (I559675,I2507,I559330,I559319,);
and I_32775 (I559313,I559421,I559610);
nor I_32776 (I559720,I559593,I41994);
and I_32777 (I559737,I559720,I41991);
or I_32778 (I559754,I559737,I42012);
DFFARX1 I_32779 (I559754,I2507,I559330,I559780,);
nor I_32780 (I559788,I559780,I559514);
DFFARX1 I_32781 (I559788,I2507,I559330,I559301,);
nand I_32782 (I559819,I559780,I559421);
nand I_32783 (I559836,I559514,I559819);
nor I_32784 (I559310,I559836,I559480);
not I_32785 (I559891,I2514);
DFFARX1 I_32786 (I1948,I2507,I559891,I559917,);
DFFARX1 I_32787 (I559917,I2507,I559891,I559934,);
not I_32788 (I559883,I559934);
not I_32789 (I559956,I559917);
DFFARX1 I_32790 (I2372,I2507,I559891,I559982,);
nand I_32791 (I559990,I559982,I1764);
not I_32792 (I560007,I1764);
not I_32793 (I560024,I2172);
nand I_32794 (I560041,I1884,I2252);
and I_32795 (I560058,I1884,I2252);
not I_32796 (I560075,I1756);
nand I_32797 (I560092,I560075,I560024);
nor I_32798 (I559865,I560092,I559990);
nor I_32799 (I560123,I560007,I560092);
nand I_32800 (I559868,I560058,I560123);
not I_32801 (I560154,I1796);
nor I_32802 (I560171,I560154,I1884);
nor I_32803 (I560188,I560171,I1756);
nor I_32804 (I560205,I559956,I560188);
DFFARX1 I_32805 (I560205,I2507,I559891,I559877,);
not I_32806 (I560236,I560171);
DFFARX1 I_32807 (I560236,I2507,I559891,I559880,);
and I_32808 (I559874,I559982,I560171);
nor I_32809 (I560281,I560154,I2308);
and I_32810 (I560298,I560281,I1916);
or I_32811 (I560315,I560298,I2188);
DFFARX1 I_32812 (I560315,I2507,I559891,I560341,);
nor I_32813 (I560349,I560341,I560075);
DFFARX1 I_32814 (I560349,I2507,I559891,I559862,);
nand I_32815 (I560380,I560341,I559982);
nand I_32816 (I560397,I560075,I560380);
nor I_32817 (I559871,I560397,I560041);
not I_32818 (I560452,I2514);
DFFARX1 I_32819 (I272688,I2507,I560452,I560478,);
DFFARX1 I_32820 (I560478,I2507,I560452,I560495,);
not I_32821 (I560444,I560495);
not I_32822 (I560517,I560478);
DFFARX1 I_32823 (I272676,I2507,I560452,I560543,);
nand I_32824 (I560551,I560543,I272682);
not I_32825 (I560568,I272682);
not I_32826 (I560585,I272679);
nand I_32827 (I560602,I272667,I272664);
and I_32828 (I560619,I272667,I272664);
not I_32829 (I560636,I272691);
nand I_32830 (I560653,I560636,I560585);
nor I_32831 (I560426,I560653,I560551);
nor I_32832 (I560684,I560568,I560653);
nand I_32833 (I560429,I560619,I560684);
not I_32834 (I560715,I272664);
nor I_32835 (I560732,I560715,I272667);
nor I_32836 (I560749,I560732,I272691);
nor I_32837 (I560766,I560517,I560749);
DFFARX1 I_32838 (I560766,I2507,I560452,I560438,);
not I_32839 (I560797,I560732);
DFFARX1 I_32840 (I560797,I2507,I560452,I560441,);
and I_32841 (I560435,I560543,I560732);
nor I_32842 (I560842,I560715,I272673);
and I_32843 (I560859,I560842,I272670);
or I_32844 (I560876,I560859,I272685);
DFFARX1 I_32845 (I560876,I2507,I560452,I560902,);
nor I_32846 (I560910,I560902,I560636);
DFFARX1 I_32847 (I560910,I2507,I560452,I560423,);
nand I_32848 (I560941,I560902,I560543);
nand I_32849 (I560958,I560636,I560941);
nor I_32850 (I560432,I560958,I560602);
not I_32851 (I561013,I2514);
DFFARX1 I_32852 (I384238,I2507,I561013,I561039,);
DFFARX1 I_32853 (I561039,I2507,I561013,I561056,);
not I_32854 (I561005,I561056);
not I_32855 (I561078,I561039);
DFFARX1 I_32856 (I384250,I2507,I561013,I561104,);
nand I_32857 (I561112,I561104,I384259);
not I_32858 (I561129,I384259);
not I_32859 (I561146,I384241);
nand I_32860 (I561163,I384244,I384235);
and I_32861 (I561180,I384244,I384235);
not I_32862 (I561197,I384253);
nand I_32863 (I561214,I561197,I561146);
nor I_32864 (I560987,I561214,I561112);
nor I_32865 (I561245,I561129,I561214);
nand I_32866 (I560990,I561180,I561245);
not I_32867 (I561276,I384256);
nor I_32868 (I561293,I561276,I384244);
nor I_32869 (I561310,I561293,I384253);
nor I_32870 (I561327,I561078,I561310);
DFFARX1 I_32871 (I561327,I2507,I561013,I560999,);
not I_32872 (I561358,I561293);
DFFARX1 I_32873 (I561358,I2507,I561013,I561002,);
and I_32874 (I560996,I561104,I561293);
nor I_32875 (I561403,I561276,I384235);
and I_32876 (I561420,I561403,I384247);
or I_32877 (I561437,I561420,I384238);
DFFARX1 I_32878 (I561437,I2507,I561013,I561463,);
nor I_32879 (I561471,I561463,I561197);
DFFARX1 I_32880 (I561471,I2507,I561013,I560984,);
nand I_32881 (I561502,I561463,I561104);
nand I_32882 (I561519,I561197,I561502);
nor I_32883 (I560993,I561519,I561163);
not I_32884 (I561574,I2514);
DFFARX1 I_32885 (I330481,I2507,I561574,I561600,);
DFFARX1 I_32886 (I561600,I2507,I561574,I561617,);
not I_32887 (I561566,I561617);
not I_32888 (I561639,I561600);
DFFARX1 I_32889 (I330496,I2507,I561574,I561665,);
nand I_32890 (I561673,I561665,I330487);
not I_32891 (I561690,I330487);
not I_32892 (I561707,I330493);
nand I_32893 (I561724,I330490,I330499);
and I_32894 (I561741,I330490,I330499);
not I_32895 (I561758,I330484);
nand I_32896 (I561775,I561758,I561707);
nor I_32897 (I561548,I561775,I561673);
nor I_32898 (I561806,I561690,I561775);
nand I_32899 (I561551,I561741,I561806);
not I_32900 (I561837,I330481);
nor I_32901 (I561854,I561837,I330490);
nor I_32902 (I561871,I561854,I330484);
nor I_32903 (I561888,I561639,I561871);
DFFARX1 I_32904 (I561888,I2507,I561574,I561560,);
not I_32905 (I561919,I561854);
DFFARX1 I_32906 (I561919,I2507,I561574,I561563,);
and I_32907 (I561557,I561665,I561854);
nor I_32908 (I561964,I561837,I330505);
and I_32909 (I561981,I561964,I330484);
or I_32910 (I561998,I561981,I330502);
DFFARX1 I_32911 (I561998,I2507,I561574,I562024,);
nor I_32912 (I562032,I562024,I561758);
DFFARX1 I_32913 (I562032,I2507,I561574,I561545,);
nand I_32914 (I562063,I562024,I561665);
nand I_32915 (I562080,I561758,I562063);
nor I_32916 (I561554,I562080,I561724);
not I_32917 (I562135,I2514);
DFFARX1 I_32918 (I461849,I2507,I562135,I562161,);
DFFARX1 I_32919 (I562161,I2507,I562135,I562178,);
not I_32920 (I562127,I562178);
not I_32921 (I562200,I562161);
DFFARX1 I_32922 (I461846,I2507,I562135,I562226,);
nand I_32923 (I562234,I562226,I461861);
not I_32924 (I562251,I461861);
not I_32925 (I562268,I461858);
nand I_32926 (I562285,I461855,I461843);
and I_32927 (I562302,I461855,I461843);
not I_32928 (I562319,I461840);
nand I_32929 (I562336,I562319,I562268);
nor I_32930 (I562109,I562336,I562234);
nor I_32931 (I562367,I562251,I562336);
nand I_32932 (I562112,I562302,I562367);
not I_32933 (I562398,I461846);
nor I_32934 (I562415,I562398,I461855);
nor I_32935 (I562432,I562415,I461840);
nor I_32936 (I562449,I562200,I562432);
DFFARX1 I_32937 (I562449,I2507,I562135,I562121,);
not I_32938 (I562480,I562415);
DFFARX1 I_32939 (I562480,I2507,I562135,I562124,);
and I_32940 (I562118,I562226,I562415);
nor I_32941 (I562525,I562398,I461852);
and I_32942 (I562542,I562525,I461840);
or I_32943 (I562559,I562542,I461843);
DFFARX1 I_32944 (I562559,I2507,I562135,I562585,);
nor I_32945 (I562593,I562585,I562319);
DFFARX1 I_32946 (I562593,I2507,I562135,I562106,);
nand I_32947 (I562624,I562585,I562226);
nand I_32948 (I562641,I562319,I562624);
nor I_32949 (I562115,I562641,I562285);
not I_32950 (I562696,I2514);
DFFARX1 I_32951 (I15659,I2507,I562696,I562722,);
DFFARX1 I_32952 (I562722,I2507,I562696,I562739,);
not I_32953 (I562688,I562739);
not I_32954 (I562761,I562722);
DFFARX1 I_32955 (I15644,I2507,I562696,I562787,);
nand I_32956 (I562795,I562787,I15656);
not I_32957 (I562812,I15656);
not I_32958 (I562829,I15662);
nand I_32959 (I562846,I15650,I15641);
and I_32960 (I562863,I15650,I15641);
not I_32961 (I562880,I15647);
nand I_32962 (I562897,I562880,I562829);
nor I_32963 (I562670,I562897,I562795);
nor I_32964 (I562928,I562812,I562897);
nand I_32965 (I562673,I562863,I562928);
not I_32966 (I562959,I15653);
nor I_32967 (I562976,I562959,I15650);
nor I_32968 (I562993,I562976,I15647);
nor I_32969 (I563010,I562761,I562993);
DFFARX1 I_32970 (I563010,I2507,I562696,I562682,);
not I_32971 (I563041,I562976);
DFFARX1 I_32972 (I563041,I2507,I562696,I562685,);
and I_32973 (I562679,I562787,I562976);
nor I_32974 (I563086,I562959,I15641);
and I_32975 (I563103,I563086,I15665);
or I_32976 (I563120,I563103,I15644);
DFFARX1 I_32977 (I563120,I2507,I562696,I563146,);
nor I_32978 (I563154,I563146,I562880);
DFFARX1 I_32979 (I563154,I2507,I562696,I562667,);
nand I_32980 (I563185,I563146,I562787);
nand I_32981 (I563202,I562880,I563185);
nor I_32982 (I562676,I563202,I562846);
not I_32983 (I563257,I2514);
DFFARX1 I_32984 (I20929,I2507,I563257,I563283,);
DFFARX1 I_32985 (I563283,I2507,I563257,I563300,);
not I_32986 (I563249,I563300);
not I_32987 (I563322,I563283);
DFFARX1 I_32988 (I20914,I2507,I563257,I563348,);
nand I_32989 (I563356,I563348,I20926);
not I_32990 (I563373,I20926);
not I_32991 (I563390,I20932);
nand I_32992 (I563407,I20920,I20911);
and I_32993 (I563424,I20920,I20911);
not I_32994 (I563441,I20917);
nand I_32995 (I563458,I563441,I563390);
nor I_32996 (I563231,I563458,I563356);
nor I_32997 (I563489,I563373,I563458);
nand I_32998 (I563234,I563424,I563489);
not I_32999 (I563520,I20923);
nor I_33000 (I563537,I563520,I20920);
nor I_33001 (I563554,I563537,I20917);
nor I_33002 (I563571,I563322,I563554);
DFFARX1 I_33003 (I563571,I2507,I563257,I563243,);
not I_33004 (I563602,I563537);
DFFARX1 I_33005 (I563602,I2507,I563257,I563246,);
and I_33006 (I563240,I563348,I563537);
nor I_33007 (I563647,I563520,I20911);
and I_33008 (I563664,I563647,I20935);
or I_33009 (I563681,I563664,I20914);
DFFARX1 I_33010 (I563681,I2507,I563257,I563707,);
nor I_33011 (I563715,I563707,I563441);
DFFARX1 I_33012 (I563715,I2507,I563257,I563228,);
nand I_33013 (I563746,I563707,I563348);
nand I_33014 (I563763,I563441,I563746);
nor I_33015 (I563237,I563763,I563407);
not I_33016 (I563818,I2514);
DFFARX1 I_33017 (I725763,I2507,I563818,I563844,);
DFFARX1 I_33018 (I563844,I2507,I563818,I563861,);
not I_33019 (I563810,I563861);
not I_33020 (I563883,I563844);
DFFARX1 I_33021 (I725757,I2507,I563818,I563909,);
nand I_33022 (I563917,I563909,I725748);
not I_33023 (I563934,I725748);
not I_33024 (I563951,I725775);
nand I_33025 (I563968,I725760,I725769);
and I_33026 (I563985,I725760,I725769);
not I_33027 (I564002,I725754);
nand I_33028 (I564019,I564002,I563951);
nor I_33029 (I563792,I564019,I563917);
nor I_33030 (I564050,I563934,I564019);
nand I_33031 (I563795,I563985,I564050);
not I_33032 (I564081,I725772);
nor I_33033 (I564098,I564081,I725760);
nor I_33034 (I564115,I564098,I725754);
nor I_33035 (I564132,I563883,I564115);
DFFARX1 I_33036 (I564132,I2507,I563818,I563804,);
not I_33037 (I564163,I564098);
DFFARX1 I_33038 (I564163,I2507,I563818,I563807,);
and I_33039 (I563801,I563909,I564098);
nor I_33040 (I564208,I564081,I725766);
and I_33041 (I564225,I564208,I725748);
or I_33042 (I564242,I564225,I725751);
DFFARX1 I_33043 (I564242,I2507,I563818,I564268,);
nor I_33044 (I564276,I564268,I564002);
DFFARX1 I_33045 (I564276,I2507,I563818,I563789,);
nand I_33046 (I564307,I564268,I563909);
nand I_33047 (I564324,I564002,I564307);
nor I_33048 (I563798,I564324,I563968);
not I_33049 (I564379,I2514);
DFFARX1 I_33050 (I699583,I2507,I564379,I564405,);
DFFARX1 I_33051 (I564405,I2507,I564379,I564422,);
not I_33052 (I564371,I564422);
not I_33053 (I564444,I564405);
DFFARX1 I_33054 (I699577,I2507,I564379,I564470,);
nand I_33055 (I564478,I564470,I699568);
not I_33056 (I564495,I699568);
not I_33057 (I564512,I699595);
nand I_33058 (I564529,I699580,I699589);
and I_33059 (I564546,I699580,I699589);
not I_33060 (I564563,I699574);
nand I_33061 (I564580,I564563,I564512);
nor I_33062 (I564353,I564580,I564478);
nor I_33063 (I564611,I564495,I564580);
nand I_33064 (I564356,I564546,I564611);
not I_33065 (I564642,I699592);
nor I_33066 (I564659,I564642,I699580);
nor I_33067 (I564676,I564659,I699574);
nor I_33068 (I564693,I564444,I564676);
DFFARX1 I_33069 (I564693,I2507,I564379,I564365,);
not I_33070 (I564724,I564659);
DFFARX1 I_33071 (I564724,I2507,I564379,I564368,);
and I_33072 (I564362,I564470,I564659);
nor I_33073 (I564769,I564642,I699586);
and I_33074 (I564786,I564769,I699568);
or I_33075 (I564803,I564786,I699571);
DFFARX1 I_33076 (I564803,I2507,I564379,I564829,);
nor I_33077 (I564837,I564829,I564563);
DFFARX1 I_33078 (I564837,I2507,I564379,I564350,);
nand I_33079 (I564868,I564829,I564470);
nand I_33080 (I564885,I564563,I564868);
nor I_33081 (I564359,I564885,I564529);
not I_33082 (I564940,I2514);
DFFARX1 I_33083 (I637584,I2507,I564940,I564966,);
DFFARX1 I_33084 (I564966,I2507,I564940,I564983,);
not I_33085 (I564932,I564983);
not I_33086 (I565005,I564966);
DFFARX1 I_33087 (I637575,I2507,I564940,I565031,);
nand I_33088 (I565039,I565031,I637572);
not I_33089 (I565056,I637572);
not I_33090 (I565073,I637581);
nand I_33091 (I565090,I637590,I637572);
and I_33092 (I565107,I637590,I637572);
not I_33093 (I565124,I637569);
nand I_33094 (I565141,I565124,I565073);
nor I_33095 (I564914,I565141,I565039);
nor I_33096 (I565172,I565056,I565141);
nand I_33097 (I564917,I565107,I565172);
not I_33098 (I565203,I637578);
nor I_33099 (I565220,I565203,I637590);
nor I_33100 (I565237,I565220,I637569);
nor I_33101 (I565254,I565005,I565237);
DFFARX1 I_33102 (I565254,I2507,I564940,I564926,);
not I_33103 (I565285,I565220);
DFFARX1 I_33104 (I565285,I2507,I564940,I564929,);
and I_33105 (I564923,I565031,I565220);
nor I_33106 (I565330,I565203,I637593);
and I_33107 (I565347,I565330,I637569);
or I_33108 (I565364,I565347,I637587);
DFFARX1 I_33109 (I565364,I2507,I564940,I565390,);
nor I_33110 (I565398,I565390,I565124);
DFFARX1 I_33111 (I565398,I2507,I564940,I564911,);
nand I_33112 (I565429,I565390,I565031);
nand I_33113 (I565446,I565124,I565429);
nor I_33114 (I564920,I565446,I565090);
not I_33115 (I565501,I2514);
DFFARX1 I_33116 (I134202,I2507,I565501,I565527,);
DFFARX1 I_33117 (I565527,I2507,I565501,I565544,);
not I_33118 (I565493,I565544);
not I_33119 (I565566,I565527);
DFFARX1 I_33120 (I134217,I2507,I565501,I565592,);
nand I_33121 (I565600,I565592,I134199);
not I_33122 (I565617,I134199);
not I_33123 (I565634,I134208);
nand I_33124 (I565651,I134214,I134205);
and I_33125 (I565668,I134214,I134205);
not I_33126 (I565685,I134202);
nand I_33127 (I565702,I565685,I565634);
nor I_33128 (I565475,I565702,I565600);
nor I_33129 (I565733,I565617,I565702);
nand I_33130 (I565478,I565668,I565733);
not I_33131 (I565764,I134199);
nor I_33132 (I565781,I565764,I134214);
nor I_33133 (I565798,I565781,I134202);
nor I_33134 (I565815,I565566,I565798);
DFFARX1 I_33135 (I565815,I2507,I565501,I565487,);
not I_33136 (I565846,I565781);
DFFARX1 I_33137 (I565846,I2507,I565501,I565490,);
and I_33138 (I565484,I565592,I565781);
nor I_33139 (I565891,I565764,I134223);
and I_33140 (I565908,I565891,I134220);
or I_33141 (I565925,I565908,I134211);
DFFARX1 I_33142 (I565925,I2507,I565501,I565951,);
nor I_33143 (I565959,I565951,I565685);
DFFARX1 I_33144 (I565959,I2507,I565501,I565472,);
nand I_33145 (I565990,I565951,I565592);
nand I_33146 (I566007,I565685,I565990);
nor I_33147 (I565481,I566007,I565651);
not I_33148 (I566062,I2514);
DFFARX1 I_33149 (I179049,I2507,I566062,I566088,);
DFFARX1 I_33150 (I566088,I2507,I566062,I566105,);
not I_33151 (I566054,I566105);
not I_33152 (I566127,I566088);
DFFARX1 I_33153 (I179046,I2507,I566062,I566153,);
nand I_33154 (I566161,I566153,I179040);
not I_33155 (I566178,I179040);
not I_33156 (I566195,I179037);
nand I_33157 (I566212,I179031,I179028);
and I_33158 (I566229,I179031,I179028);
not I_33159 (I566246,I179043);
nand I_33160 (I566263,I566246,I566195);
nor I_33161 (I566036,I566263,I566161);
nor I_33162 (I566294,I566178,I566263);
nand I_33163 (I566039,I566229,I566294);
not I_33164 (I566325,I179055);
nor I_33165 (I566342,I566325,I179031);
nor I_33166 (I566359,I566342,I179043);
nor I_33167 (I566376,I566127,I566359);
DFFARX1 I_33168 (I566376,I2507,I566062,I566048,);
not I_33169 (I566407,I566342);
DFFARX1 I_33170 (I566407,I2507,I566062,I566051,);
and I_33171 (I566045,I566153,I566342);
nor I_33172 (I566452,I566325,I179052);
and I_33173 (I566469,I566452,I179028);
or I_33174 (I566486,I566469,I179034);
DFFARX1 I_33175 (I566486,I2507,I566062,I566512,);
nor I_33176 (I566520,I566512,I566246);
DFFARX1 I_33177 (I566520,I2507,I566062,I566033,);
nand I_33178 (I566551,I566512,I566153);
nand I_33179 (I566568,I566246,I566551);
nor I_33180 (I566042,I566568,I566212);
not I_33181 (I566623,I2514);
DFFARX1 I_33182 (I238960,I2507,I566623,I566649,);
DFFARX1 I_33183 (I566649,I2507,I566623,I566666,);
not I_33184 (I566615,I566666);
not I_33185 (I566688,I566649);
DFFARX1 I_33186 (I238948,I2507,I566623,I566714,);
nand I_33187 (I566722,I566714,I238954);
not I_33188 (I566739,I238954);
not I_33189 (I566756,I238951);
nand I_33190 (I566773,I238939,I238936);
and I_33191 (I566790,I238939,I238936);
not I_33192 (I566807,I238963);
nand I_33193 (I566824,I566807,I566756);
nor I_33194 (I566597,I566824,I566722);
nor I_33195 (I566855,I566739,I566824);
nand I_33196 (I566600,I566790,I566855);
not I_33197 (I566886,I238936);
nor I_33198 (I566903,I566886,I238939);
nor I_33199 (I566920,I566903,I238963);
nor I_33200 (I566937,I566688,I566920);
DFFARX1 I_33201 (I566937,I2507,I566623,I566609,);
not I_33202 (I566968,I566903);
DFFARX1 I_33203 (I566968,I2507,I566623,I566612,);
and I_33204 (I566606,I566714,I566903);
nor I_33205 (I567013,I566886,I238945);
and I_33206 (I567030,I567013,I238942);
or I_33207 (I567047,I567030,I238957);
DFFARX1 I_33208 (I567047,I2507,I566623,I567073,);
nor I_33209 (I567081,I567073,I566807);
DFFARX1 I_33210 (I567081,I2507,I566623,I566594,);
nand I_33211 (I567112,I567073,I566714);
nand I_33212 (I567129,I566807,I567112);
nor I_33213 (I566603,I567129,I566773);
not I_33214 (I567184,I2514);
DFFARX1 I_33215 (I288526,I2507,I567184,I567210,);
DFFARX1 I_33216 (I567210,I2507,I567184,I567227,);
not I_33217 (I567176,I567227);
not I_33218 (I567249,I567210);
DFFARX1 I_33219 (I288523,I2507,I567184,I567275,);
nand I_33220 (I567283,I567275,I288517);
not I_33221 (I567300,I288517);
not I_33222 (I567317,I288529);
nand I_33223 (I567334,I288532,I288511);
and I_33224 (I567351,I288532,I288511);
not I_33225 (I567368,I288508);
nand I_33226 (I567385,I567368,I567317);
nor I_33227 (I567158,I567385,I567283);
nor I_33228 (I567416,I567300,I567385);
nand I_33229 (I567161,I567351,I567416);
not I_33230 (I567447,I288514);
nor I_33231 (I567464,I567447,I288532);
nor I_33232 (I567481,I567464,I288508);
nor I_33233 (I567498,I567249,I567481);
DFFARX1 I_33234 (I567498,I2507,I567184,I567170,);
not I_33235 (I567529,I567464);
DFFARX1 I_33236 (I567529,I2507,I567184,I567173,);
and I_33237 (I567167,I567275,I567464);
nor I_33238 (I567574,I567447,I288508);
and I_33239 (I567591,I567574,I288520);
or I_33240 (I567608,I567591,I288511);
DFFARX1 I_33241 (I567608,I2507,I567184,I567634,);
nor I_33242 (I567642,I567634,I567368);
DFFARX1 I_33243 (I567642,I2507,I567184,I567155,);
nand I_33244 (I567673,I567634,I567275);
nand I_33245 (I567690,I567368,I567673);
nor I_33246 (I567164,I567690,I567334);
not I_33247 (I567745,I2514);
DFFARX1 I_33248 (I341463,I2507,I567745,I567771,);
DFFARX1 I_33249 (I567771,I2507,I567745,I567788,);
not I_33250 (I567737,I567788);
not I_33251 (I567810,I567771);
DFFARX1 I_33252 (I341478,I2507,I567745,I567836,);
nand I_33253 (I567844,I567836,I341469);
not I_33254 (I567861,I341469);
not I_33255 (I567878,I341475);
nand I_33256 (I567895,I341472,I341481);
and I_33257 (I567912,I341472,I341481);
not I_33258 (I567929,I341466);
nand I_33259 (I567946,I567929,I567878);
nor I_33260 (I567719,I567946,I567844);
nor I_33261 (I567977,I567861,I567946);
nand I_33262 (I567722,I567912,I567977);
not I_33263 (I568008,I341463);
nor I_33264 (I568025,I568008,I341472);
nor I_33265 (I568042,I568025,I341466);
nor I_33266 (I568059,I567810,I568042);
DFFARX1 I_33267 (I568059,I2507,I567745,I567731,);
not I_33268 (I568090,I568025);
DFFARX1 I_33269 (I568090,I2507,I567745,I567734,);
and I_33270 (I567728,I567836,I568025);
nor I_33271 (I568135,I568008,I341487);
and I_33272 (I568152,I568135,I341466);
or I_33273 (I568169,I568152,I341484);
DFFARX1 I_33274 (I568169,I2507,I567745,I568195,);
nor I_33275 (I568203,I568195,I567929);
DFFARX1 I_33276 (I568203,I2507,I567745,I567716,);
nand I_33277 (I568234,I568195,I567836);
nand I_33278 (I568251,I567929,I568234);
nor I_33279 (I567725,I568251,I567895);
not I_33280 (I568306,I2514);
DFFARX1 I_33281 (I358806,I2507,I568306,I568332,);
DFFARX1 I_33282 (I568332,I2507,I568306,I568349,);
not I_33283 (I568298,I568349);
not I_33284 (I568371,I568332);
DFFARX1 I_33285 (I358818,I2507,I568306,I568397,);
nand I_33286 (I568405,I568397,I358827);
not I_33287 (I568422,I358827);
not I_33288 (I568439,I358809);
nand I_33289 (I568456,I358812,I358803);
and I_33290 (I568473,I358812,I358803);
not I_33291 (I568490,I358821);
nand I_33292 (I568507,I568490,I568439);
nor I_33293 (I568280,I568507,I568405);
nor I_33294 (I568538,I568422,I568507);
nand I_33295 (I568283,I568473,I568538);
not I_33296 (I568569,I358824);
nor I_33297 (I568586,I568569,I358812);
nor I_33298 (I568603,I568586,I358821);
nor I_33299 (I568620,I568371,I568603);
DFFARX1 I_33300 (I568620,I2507,I568306,I568292,);
not I_33301 (I568651,I568586);
DFFARX1 I_33302 (I568651,I2507,I568306,I568295,);
and I_33303 (I568289,I568397,I568586);
nor I_33304 (I568696,I568569,I358803);
and I_33305 (I568713,I568696,I358815);
or I_33306 (I568730,I568713,I358806);
DFFARX1 I_33307 (I568730,I2507,I568306,I568756,);
nor I_33308 (I568764,I568756,I568490);
DFFARX1 I_33309 (I568764,I2507,I568306,I568277,);
nand I_33310 (I568795,I568756,I568397);
nand I_33311 (I568812,I568490,I568795);
nor I_33312 (I568286,I568812,I568456);
not I_33313 (I568867,I2514);
DFFARX1 I_33314 (I42530,I2507,I568867,I568893,);
DFFARX1 I_33315 (I568893,I2507,I568867,I568910,);
not I_33316 (I568859,I568910);
not I_33317 (I568932,I568893);
DFFARX1 I_33318 (I42518,I2507,I568867,I568958,);
nand I_33319 (I568966,I568958,I42533);
not I_33320 (I568983,I42533);
not I_33321 (I569000,I42521);
nand I_33322 (I569017,I42542,I42536);
and I_33323 (I569034,I42542,I42536);
not I_33324 (I569051,I42524);
nand I_33325 (I569068,I569051,I569000);
nor I_33326 (I568841,I569068,I568966);
nor I_33327 (I569099,I568983,I569068);
nand I_33328 (I568844,I569034,I569099);
not I_33329 (I569130,I42527);
nor I_33330 (I569147,I569130,I42542);
nor I_33331 (I569164,I569147,I42524);
nor I_33332 (I569181,I568932,I569164);
DFFARX1 I_33333 (I569181,I2507,I568867,I568853,);
not I_33334 (I569212,I569147);
DFFARX1 I_33335 (I569212,I2507,I568867,I568856,);
and I_33336 (I568850,I568958,I569147);
nor I_33337 (I569257,I569130,I42521);
and I_33338 (I569274,I569257,I42518);
or I_33339 (I569291,I569274,I42539);
DFFARX1 I_33340 (I569291,I2507,I568867,I569317,);
nor I_33341 (I569325,I569317,I569051);
DFFARX1 I_33342 (I569325,I2507,I568867,I568838,);
nand I_33343 (I569356,I569317,I568958);
nand I_33344 (I569373,I569051,I569356);
nor I_33345 (I568847,I569373,I569017);
not I_33346 (I569428,I2514);
DFFARX1 I_33347 (I200129,I2507,I569428,I569454,);
DFFARX1 I_33348 (I569454,I2507,I569428,I569471,);
not I_33349 (I569420,I569471);
not I_33350 (I569493,I569454);
DFFARX1 I_33351 (I200126,I2507,I569428,I569519,);
nand I_33352 (I569527,I569519,I200120);
not I_33353 (I569544,I200120);
not I_33354 (I569561,I200117);
nand I_33355 (I569578,I200111,I200108);
and I_33356 (I569595,I200111,I200108);
not I_33357 (I569612,I200123);
nand I_33358 (I569629,I569612,I569561);
nor I_33359 (I569402,I569629,I569527);
nor I_33360 (I569660,I569544,I569629);
nand I_33361 (I569405,I569595,I569660);
not I_33362 (I569691,I200135);
nor I_33363 (I569708,I569691,I200111);
nor I_33364 (I569725,I569708,I200123);
nor I_33365 (I569742,I569493,I569725);
DFFARX1 I_33366 (I569742,I2507,I569428,I569414,);
not I_33367 (I569773,I569708);
DFFARX1 I_33368 (I569773,I2507,I569428,I569417,);
and I_33369 (I569411,I569519,I569708);
nor I_33370 (I569818,I569691,I200132);
and I_33371 (I569835,I569818,I200108);
or I_33372 (I569852,I569835,I200114);
DFFARX1 I_33373 (I569852,I2507,I569428,I569878,);
nor I_33374 (I569886,I569878,I569612);
DFFARX1 I_33375 (I569886,I2507,I569428,I569399,);
nand I_33376 (I569917,I569878,I569519);
nand I_33377 (I569934,I569612,I569917);
nor I_33378 (I569408,I569934,I569578);
not I_33379 (I569989,I2514);
DFFARX1 I_33380 (I128847,I2507,I569989,I570015,);
DFFARX1 I_33381 (I570015,I2507,I569989,I570032,);
not I_33382 (I569981,I570032);
not I_33383 (I570054,I570015);
DFFARX1 I_33384 (I128862,I2507,I569989,I570080,);
nand I_33385 (I570088,I570080,I128844);
not I_33386 (I570105,I128844);
not I_33387 (I570122,I128853);
nand I_33388 (I570139,I128859,I128850);
and I_33389 (I570156,I128859,I128850);
not I_33390 (I570173,I128847);
nand I_33391 (I570190,I570173,I570122);
nor I_33392 (I569963,I570190,I570088);
nor I_33393 (I570221,I570105,I570190);
nand I_33394 (I569966,I570156,I570221);
not I_33395 (I570252,I128844);
nor I_33396 (I570269,I570252,I128859);
nor I_33397 (I570286,I570269,I128847);
nor I_33398 (I570303,I570054,I570286);
DFFARX1 I_33399 (I570303,I2507,I569989,I569975,);
not I_33400 (I570334,I570269);
DFFARX1 I_33401 (I570334,I2507,I569989,I569978,);
and I_33402 (I569972,I570080,I570269);
nor I_33403 (I570379,I570252,I128868);
and I_33404 (I570396,I570379,I128865);
or I_33405 (I570413,I570396,I128856);
DFFARX1 I_33406 (I570413,I2507,I569989,I570439,);
nor I_33407 (I570447,I570439,I570173);
DFFARX1 I_33408 (I570447,I2507,I569989,I569960,);
nand I_33409 (I570478,I570439,I570080);
nand I_33410 (I570495,I570173,I570478);
nor I_33411 (I569969,I570495,I570139);
not I_33412 (I570553,I2514);
DFFARX1 I_33413 (I276472,I2507,I570553,I570579,);
and I_33414 (I570587,I570579,I276487);
DFFARX1 I_33415 (I570587,I2507,I570553,I570536,);
DFFARX1 I_33416 (I276490,I2507,I570553,I570627,);
not I_33417 (I570635,I276484);
not I_33418 (I570652,I276499);
nand I_33419 (I570669,I570652,I570635);
nor I_33420 (I570524,I570627,I570669);
DFFARX1 I_33421 (I570669,I2507,I570553,I570709,);
not I_33422 (I570545,I570709);
not I_33423 (I570731,I276475);
nand I_33424 (I570748,I570652,I570731);
DFFARX1 I_33425 (I570748,I2507,I570553,I570774,);
not I_33426 (I570782,I570774);
not I_33427 (I570799,I276478);
nand I_33428 (I570816,I570799,I276472);
and I_33429 (I570833,I570635,I570816);
nor I_33430 (I570850,I570748,I570833);
DFFARX1 I_33431 (I570850,I2507,I570553,I570521,);
DFFARX1 I_33432 (I570833,I2507,I570553,I570542,);
nor I_33433 (I570895,I276478,I276481);
nor I_33434 (I570533,I570748,I570895);
or I_33435 (I570926,I276478,I276481);
nor I_33436 (I570943,I276496,I276493);
DFFARX1 I_33437 (I570943,I2507,I570553,I570969,);
not I_33438 (I570977,I570969);
nor I_33439 (I570539,I570977,I570782);
nand I_33440 (I571008,I570977,I570627);
not I_33441 (I571025,I276496);
nand I_33442 (I571042,I571025,I570731);
nand I_33443 (I571059,I570977,I571042);
nand I_33444 (I570530,I571059,I571008);
nand I_33445 (I570527,I571042,I570926);
not I_33446 (I571131,I2514);
DFFARX1 I_33447 (I694240,I2507,I571131,I571157,);
and I_33448 (I571165,I571157,I694222);
DFFARX1 I_33449 (I571165,I2507,I571131,I571114,);
DFFARX1 I_33450 (I694213,I2507,I571131,I571205,);
not I_33451 (I571213,I694228);
not I_33452 (I571230,I694216);
nand I_33453 (I571247,I571230,I571213);
nor I_33454 (I571102,I571205,I571247);
DFFARX1 I_33455 (I571247,I2507,I571131,I571287,);
not I_33456 (I571123,I571287);
not I_33457 (I571309,I694225);
nand I_33458 (I571326,I571230,I571309);
DFFARX1 I_33459 (I571326,I2507,I571131,I571352,);
not I_33460 (I571360,I571352);
not I_33461 (I571377,I694234);
nand I_33462 (I571394,I571377,I694213);
and I_33463 (I571411,I571213,I571394);
nor I_33464 (I571428,I571326,I571411);
DFFARX1 I_33465 (I571428,I2507,I571131,I571099,);
DFFARX1 I_33466 (I571411,I2507,I571131,I571120,);
nor I_33467 (I571473,I694234,I694237);
nor I_33468 (I571111,I571326,I571473);
or I_33469 (I571504,I694234,I694237);
nor I_33470 (I571521,I694231,I694219);
DFFARX1 I_33471 (I571521,I2507,I571131,I571547,);
not I_33472 (I571555,I571547);
nor I_33473 (I571117,I571555,I571360);
nand I_33474 (I571586,I571555,I571205);
not I_33475 (I571603,I694231);
nand I_33476 (I571620,I571603,I571309);
nand I_33477 (I571637,I571555,I571620);
nand I_33478 (I571108,I571637,I571586);
nand I_33479 (I571105,I571620,I571504);
not I_33480 (I571709,I2514);
DFFARX1 I_33481 (I528044,I2507,I571709,I571735,);
and I_33482 (I571743,I571735,I528038);
DFFARX1 I_33483 (I571743,I2507,I571709,I571692,);
DFFARX1 I_33484 (I528056,I2507,I571709,I571783,);
not I_33485 (I571791,I528047);
not I_33486 (I571808,I528059);
nand I_33487 (I571825,I571808,I571791);
nor I_33488 (I571680,I571783,I571825);
DFFARX1 I_33489 (I571825,I2507,I571709,I571865,);
not I_33490 (I571701,I571865);
not I_33491 (I571887,I528065);
nand I_33492 (I571904,I571808,I571887);
DFFARX1 I_33493 (I571904,I2507,I571709,I571930,);
not I_33494 (I571938,I571930);
not I_33495 (I571955,I528041);
nand I_33496 (I571972,I571955,I528062);
and I_33497 (I571989,I571791,I571972);
nor I_33498 (I572006,I571904,I571989);
DFFARX1 I_33499 (I572006,I2507,I571709,I571677,);
DFFARX1 I_33500 (I571989,I2507,I571709,I571698,);
nor I_33501 (I572051,I528041,I528053);
nor I_33502 (I571689,I571904,I572051);
or I_33503 (I572082,I528041,I528053);
nor I_33504 (I572099,I528038,I528050);
DFFARX1 I_33505 (I572099,I2507,I571709,I572125,);
not I_33506 (I572133,I572125);
nor I_33507 (I571695,I572133,I571938);
nand I_33508 (I572164,I572133,I571783);
not I_33509 (I572181,I528038);
nand I_33510 (I572198,I572181,I571887);
nand I_33511 (I572215,I572133,I572198);
nand I_33512 (I571686,I572215,I572164);
nand I_33513 (I571683,I572198,I572082);
not I_33514 (I572287,I2514);
DFFARX1 I_33515 (I243288,I2507,I572287,I572313,);
and I_33516 (I572321,I572313,I243303);
DFFARX1 I_33517 (I572321,I2507,I572287,I572270,);
DFFARX1 I_33518 (I243306,I2507,I572287,I572361,);
not I_33519 (I572369,I243300);
not I_33520 (I572386,I243315);
nand I_33521 (I572403,I572386,I572369);
nor I_33522 (I572258,I572361,I572403);
DFFARX1 I_33523 (I572403,I2507,I572287,I572443,);
not I_33524 (I572279,I572443);
not I_33525 (I572465,I243291);
nand I_33526 (I572482,I572386,I572465);
DFFARX1 I_33527 (I572482,I2507,I572287,I572508,);
not I_33528 (I572516,I572508);
not I_33529 (I572533,I243294);
nand I_33530 (I572550,I572533,I243288);
and I_33531 (I572567,I572369,I572550);
nor I_33532 (I572584,I572482,I572567);
DFFARX1 I_33533 (I572584,I2507,I572287,I572255,);
DFFARX1 I_33534 (I572567,I2507,I572287,I572276,);
nor I_33535 (I572629,I243294,I243297);
nor I_33536 (I572267,I572482,I572629);
or I_33537 (I572660,I243294,I243297);
nor I_33538 (I572677,I243312,I243309);
DFFARX1 I_33539 (I572677,I2507,I572287,I572703,);
not I_33540 (I572711,I572703);
nor I_33541 (I572273,I572711,I572516);
nand I_33542 (I572742,I572711,I572361);
not I_33543 (I572759,I243312);
nand I_33544 (I572776,I572759,I572465);
nand I_33545 (I572793,I572711,I572776);
nand I_33546 (I572264,I572793,I572742);
nand I_33547 (I572261,I572776,I572660);
not I_33548 (I572865,I2514);
DFFARX1 I_33549 (I258520,I2507,I572865,I572891,);
and I_33550 (I572899,I572891,I258535);
DFFARX1 I_33551 (I572899,I2507,I572865,I572848,);
DFFARX1 I_33552 (I258538,I2507,I572865,I572939,);
not I_33553 (I572947,I258532);
not I_33554 (I572964,I258547);
nand I_33555 (I572981,I572964,I572947);
nor I_33556 (I572836,I572939,I572981);
DFFARX1 I_33557 (I572981,I2507,I572865,I573021,);
not I_33558 (I572857,I573021);
not I_33559 (I573043,I258523);
nand I_33560 (I573060,I572964,I573043);
DFFARX1 I_33561 (I573060,I2507,I572865,I573086,);
not I_33562 (I573094,I573086);
not I_33563 (I573111,I258526);
nand I_33564 (I573128,I573111,I258520);
and I_33565 (I573145,I572947,I573128);
nor I_33566 (I573162,I573060,I573145);
DFFARX1 I_33567 (I573162,I2507,I572865,I572833,);
DFFARX1 I_33568 (I573145,I2507,I572865,I572854,);
nor I_33569 (I573207,I258526,I258529);
nor I_33570 (I572845,I573060,I573207);
or I_33571 (I573238,I258526,I258529);
nor I_33572 (I573255,I258544,I258541);
DFFARX1 I_33573 (I573255,I2507,I572865,I573281,);
not I_33574 (I573289,I573281);
nor I_33575 (I572851,I573289,I573094);
nand I_33576 (I573320,I573289,I572939);
not I_33577 (I573337,I258544);
nand I_33578 (I573354,I573337,I573043);
nand I_33579 (I573371,I573289,I573354);
nand I_33580 (I572842,I573371,I573320);
nand I_33581 (I572839,I573354,I573238);
not I_33582 (I573443,I2514);
DFFARX1 I_33583 (I566036,I2507,I573443,I573469,);
and I_33584 (I573477,I573469,I566033);
DFFARX1 I_33585 (I573477,I2507,I573443,I573426,);
DFFARX1 I_33586 (I566039,I2507,I573443,I573517,);
not I_33587 (I573525,I566042);
not I_33588 (I573542,I566036);
nand I_33589 (I573559,I573542,I573525);
nor I_33590 (I573414,I573517,I573559);
DFFARX1 I_33591 (I573559,I2507,I573443,I573599,);
not I_33592 (I573435,I573599);
not I_33593 (I573621,I566051);
nand I_33594 (I573638,I573542,I573621);
DFFARX1 I_33595 (I573638,I2507,I573443,I573664,);
not I_33596 (I573672,I573664);
not I_33597 (I573689,I566048);
nand I_33598 (I573706,I573689,I566054);
and I_33599 (I573723,I573525,I573706);
nor I_33600 (I573740,I573638,I573723);
DFFARX1 I_33601 (I573740,I2507,I573443,I573411,);
DFFARX1 I_33602 (I573723,I2507,I573443,I573432,);
nor I_33603 (I573785,I566048,I566033);
nor I_33604 (I573423,I573638,I573785);
or I_33605 (I573816,I566048,I566033);
nor I_33606 (I573833,I566045,I566039);
DFFARX1 I_33607 (I573833,I2507,I573443,I573859,);
not I_33608 (I573867,I573859);
nor I_33609 (I573429,I573867,I573672);
nand I_33610 (I573898,I573867,I573517);
not I_33611 (I573915,I566045);
nand I_33612 (I573932,I573915,I573621);
nand I_33613 (I573949,I573867,I573932);
nand I_33614 (I573420,I573949,I573898);
nand I_33615 (I573417,I573932,I573816);
not I_33616 (I574021,I2514);
DFFARX1 I_33617 (I190649,I2507,I574021,I574047,);
and I_33618 (I574055,I574047,I190634);
DFFARX1 I_33619 (I574055,I2507,I574021,I574004,);
DFFARX1 I_33620 (I190640,I2507,I574021,I574095,);
not I_33621 (I574103,I190622);
not I_33622 (I574120,I190643);
nand I_33623 (I574137,I574120,I574103);
nor I_33624 (I573992,I574095,I574137);
DFFARX1 I_33625 (I574137,I2507,I574021,I574177,);
not I_33626 (I574013,I574177);
not I_33627 (I574199,I190646);
nand I_33628 (I574216,I574120,I574199);
DFFARX1 I_33629 (I574216,I2507,I574021,I574242,);
not I_33630 (I574250,I574242);
not I_33631 (I574267,I190637);
nand I_33632 (I574284,I574267,I190625);
and I_33633 (I574301,I574103,I574284);
nor I_33634 (I574318,I574216,I574301);
DFFARX1 I_33635 (I574318,I2507,I574021,I573989,);
DFFARX1 I_33636 (I574301,I2507,I574021,I574010,);
nor I_33637 (I574363,I190637,I190631);
nor I_33638 (I574001,I574216,I574363);
or I_33639 (I574394,I190637,I190631);
nor I_33640 (I574411,I190628,I190622);
DFFARX1 I_33641 (I574411,I2507,I574021,I574437,);
not I_33642 (I574445,I574437);
nor I_33643 (I574007,I574445,I574250);
nand I_33644 (I574476,I574445,I574095);
not I_33645 (I574493,I190628);
nand I_33646 (I574510,I574493,I574199);
nand I_33647 (I574527,I574445,I574510);
nand I_33648 (I573998,I574527,I574476);
nand I_33649 (I573995,I574510,I574394);
not I_33650 (I574599,I2514);
DFFARX1 I_33651 (I150264,I2507,I574599,I574625,);
and I_33652 (I574633,I574625,I150267);
DFFARX1 I_33653 (I574633,I2507,I574599,I574582,);
DFFARX1 I_33654 (I150267,I2507,I574599,I574673,);
not I_33655 (I574681,I150282);
not I_33656 (I574698,I150288);
nand I_33657 (I574715,I574698,I574681);
nor I_33658 (I574570,I574673,I574715);
DFFARX1 I_33659 (I574715,I2507,I574599,I574755,);
not I_33660 (I574591,I574755);
not I_33661 (I574777,I150276);
nand I_33662 (I574794,I574698,I574777);
DFFARX1 I_33663 (I574794,I2507,I574599,I574820,);
not I_33664 (I574828,I574820);
not I_33665 (I574845,I150273);
nand I_33666 (I574862,I574845,I150270);
and I_33667 (I574879,I574681,I574862);
nor I_33668 (I574896,I574794,I574879);
DFFARX1 I_33669 (I574896,I2507,I574599,I574567,);
DFFARX1 I_33670 (I574879,I2507,I574599,I574588,);
nor I_33671 (I574941,I150273,I150264);
nor I_33672 (I574579,I574794,I574941);
or I_33673 (I574972,I150273,I150264);
nor I_33674 (I574989,I150279,I150285);
DFFARX1 I_33675 (I574989,I2507,I574599,I575015,);
not I_33676 (I575023,I575015);
nor I_33677 (I574585,I575023,I574828);
nand I_33678 (I575054,I575023,I574673);
not I_33679 (I575071,I150279);
nand I_33680 (I575088,I575071,I574777);
nand I_33681 (I575105,I575023,I575088);
nand I_33682 (I574576,I575105,I575054);
nand I_33683 (I574573,I575088,I574972);
not I_33684 (I575177,I2514);
DFFARX1 I_33685 (I14060,I2507,I575177,I575203,);
and I_33686 (I575211,I575203,I14063);
DFFARX1 I_33687 (I575211,I2507,I575177,I575160,);
DFFARX1 I_33688 (I14063,I2507,I575177,I575251,);
not I_33689 (I575259,I14066);
not I_33690 (I575276,I14081);
nand I_33691 (I575293,I575276,I575259);
nor I_33692 (I575148,I575251,I575293);
DFFARX1 I_33693 (I575293,I2507,I575177,I575333,);
not I_33694 (I575169,I575333);
not I_33695 (I575355,I14075);
nand I_33696 (I575372,I575276,I575355);
DFFARX1 I_33697 (I575372,I2507,I575177,I575398,);
not I_33698 (I575406,I575398);
not I_33699 (I575423,I14078);
nand I_33700 (I575440,I575423,I14060);
and I_33701 (I575457,I575259,I575440);
nor I_33702 (I575474,I575372,I575457);
DFFARX1 I_33703 (I575474,I2507,I575177,I575145,);
DFFARX1 I_33704 (I575457,I2507,I575177,I575166,);
nor I_33705 (I575519,I14078,I14072);
nor I_33706 (I575157,I575372,I575519);
or I_33707 (I575550,I14078,I14072);
nor I_33708 (I575567,I14069,I14084);
DFFARX1 I_33709 (I575567,I2507,I575177,I575593,);
not I_33710 (I575601,I575593);
nor I_33711 (I575163,I575601,I575406);
nand I_33712 (I575632,I575601,I575251);
not I_33713 (I575649,I14069);
nand I_33714 (I575666,I575649,I575355);
nand I_33715 (I575683,I575601,I575666);
nand I_33716 (I575154,I575683,I575632);
nand I_33717 (I575151,I575666,I575550);
not I_33718 (I575755,I2514);
DFFARX1 I_33719 (I180109,I2507,I575755,I575781,);
and I_33720 (I575789,I575781,I180094);
DFFARX1 I_33721 (I575789,I2507,I575755,I575738,);
DFFARX1 I_33722 (I180100,I2507,I575755,I575829,);
not I_33723 (I575837,I180082);
not I_33724 (I575854,I180103);
nand I_33725 (I575871,I575854,I575837);
nor I_33726 (I575726,I575829,I575871);
DFFARX1 I_33727 (I575871,I2507,I575755,I575911,);
not I_33728 (I575747,I575911);
not I_33729 (I575933,I180106);
nand I_33730 (I575950,I575854,I575933);
DFFARX1 I_33731 (I575950,I2507,I575755,I575976,);
not I_33732 (I575984,I575976);
not I_33733 (I576001,I180097);
nand I_33734 (I576018,I576001,I180085);
and I_33735 (I576035,I575837,I576018);
nor I_33736 (I576052,I575950,I576035);
DFFARX1 I_33737 (I576052,I2507,I575755,I575723,);
DFFARX1 I_33738 (I576035,I2507,I575755,I575744,);
nor I_33739 (I576097,I180097,I180091);
nor I_33740 (I575735,I575950,I576097);
or I_33741 (I576128,I180097,I180091);
nor I_33742 (I576145,I180088,I180082);
DFFARX1 I_33743 (I576145,I2507,I575755,I576171,);
not I_33744 (I576179,I576171);
nor I_33745 (I575741,I576179,I575984);
nand I_33746 (I576210,I576179,I575829);
not I_33747 (I576227,I180088);
nand I_33748 (I576244,I576227,I575933);
nand I_33749 (I576261,I576179,I576244);
nand I_33750 (I575732,I576261,I576210);
nand I_33751 (I575729,I576244,I576128);
not I_33752 (I576333,I2514);
DFFARX1 I_33753 (I389452,I2507,I576333,I576359,);
and I_33754 (I576367,I576359,I389440);
DFFARX1 I_33755 (I576367,I2507,I576333,I576316,);
DFFARX1 I_33756 (I389443,I2507,I576333,I576407,);
not I_33757 (I576415,I389437);
not I_33758 (I576432,I389461);
nand I_33759 (I576449,I576432,I576415);
nor I_33760 (I576304,I576407,I576449);
DFFARX1 I_33761 (I576449,I2507,I576333,I576489,);
not I_33762 (I576325,I576489);
not I_33763 (I576511,I389449);
nand I_33764 (I576528,I576432,I576511);
DFFARX1 I_33765 (I576528,I2507,I576333,I576554,);
not I_33766 (I576562,I576554);
not I_33767 (I576579,I389458);
nand I_33768 (I576596,I576579,I389455);
and I_33769 (I576613,I576415,I576596);
nor I_33770 (I576630,I576528,I576613);
DFFARX1 I_33771 (I576630,I2507,I576333,I576301,);
DFFARX1 I_33772 (I576613,I2507,I576333,I576322,);
nor I_33773 (I576675,I389458,I389446);
nor I_33774 (I576313,I576528,I576675);
or I_33775 (I576706,I389458,I389446);
nor I_33776 (I576723,I389437,I389440);
DFFARX1 I_33777 (I576723,I2507,I576333,I576749,);
not I_33778 (I576757,I576749);
nor I_33779 (I576319,I576757,I576562);
nand I_33780 (I576788,I576757,I576407);
not I_33781 (I576805,I389437);
nand I_33782 (I576822,I576805,I576511);
nand I_33783 (I576839,I576757,I576822);
nand I_33784 (I576310,I576839,I576788);
nand I_33785 (I576307,I576822,I576706);
not I_33786 (I576911,I2514);
DFFARX1 I_33787 (I726370,I2507,I576911,I576937,);
and I_33788 (I576945,I576937,I726352);
DFFARX1 I_33789 (I576945,I2507,I576911,I576894,);
DFFARX1 I_33790 (I726343,I2507,I576911,I576985,);
not I_33791 (I576993,I726358);
not I_33792 (I577010,I726346);
nand I_33793 (I577027,I577010,I576993);
nor I_33794 (I576882,I576985,I577027);
DFFARX1 I_33795 (I577027,I2507,I576911,I577067,);
not I_33796 (I576903,I577067);
not I_33797 (I577089,I726355);
nand I_33798 (I577106,I577010,I577089);
DFFARX1 I_33799 (I577106,I2507,I576911,I577132,);
not I_33800 (I577140,I577132);
not I_33801 (I577157,I726364);
nand I_33802 (I577174,I577157,I726343);
and I_33803 (I577191,I576993,I577174);
nor I_33804 (I577208,I577106,I577191);
DFFARX1 I_33805 (I577208,I2507,I576911,I576879,);
DFFARX1 I_33806 (I577191,I2507,I576911,I576900,);
nor I_33807 (I577253,I726364,I726367);
nor I_33808 (I576891,I577106,I577253);
or I_33809 (I577284,I726364,I726367);
nor I_33810 (I577301,I726361,I726349);
DFFARX1 I_33811 (I577301,I2507,I576911,I577327,);
not I_33812 (I577335,I577327);
nor I_33813 (I576897,I577335,I577140);
nand I_33814 (I577366,I577335,I576985);
not I_33815 (I577383,I726361);
nand I_33816 (I577400,I577383,I577089);
nand I_33817 (I577417,I577335,I577400);
nand I_33818 (I576888,I577417,I577366);
nand I_33819 (I576885,I577400,I577284);
not I_33820 (I577489,I2514);
DFFARX1 I_33821 (I16168,I2507,I577489,I577515,);
and I_33822 (I577523,I577515,I16171);
DFFARX1 I_33823 (I577523,I2507,I577489,I577472,);
DFFARX1 I_33824 (I16171,I2507,I577489,I577563,);
not I_33825 (I577571,I16174);
not I_33826 (I577588,I16189);
nand I_33827 (I577605,I577588,I577571);
nor I_33828 (I577460,I577563,I577605);
DFFARX1 I_33829 (I577605,I2507,I577489,I577645,);
not I_33830 (I577481,I577645);
not I_33831 (I577667,I16183);
nand I_33832 (I577684,I577588,I577667);
DFFARX1 I_33833 (I577684,I2507,I577489,I577710,);
not I_33834 (I577718,I577710);
not I_33835 (I577735,I16186);
nand I_33836 (I577752,I577735,I16168);
and I_33837 (I577769,I577571,I577752);
nor I_33838 (I577786,I577684,I577769);
DFFARX1 I_33839 (I577786,I2507,I577489,I577457,);
DFFARX1 I_33840 (I577769,I2507,I577489,I577478,);
nor I_33841 (I577831,I16186,I16180);
nor I_33842 (I577469,I577684,I577831);
or I_33843 (I577862,I16186,I16180);
nor I_33844 (I577879,I16177,I16192);
DFFARX1 I_33845 (I577879,I2507,I577489,I577905,);
not I_33846 (I577913,I577905);
nor I_33847 (I577475,I577913,I577718);
nand I_33848 (I577944,I577913,I577563);
not I_33849 (I577961,I16177);
nand I_33850 (I577978,I577961,I577667);
nand I_33851 (I577995,I577913,I577978);
nand I_33852 (I577466,I577995,I577944);
nand I_33853 (I577463,I577978,I577862);
not I_33854 (I578067,I2514);
DFFARX1 I_33855 (I2148,I2507,I578067,I578093,);
and I_33856 (I578101,I578093,I2428);
DFFARX1 I_33857 (I578101,I2507,I578067,I578050,);
DFFARX1 I_33858 (I2180,I2507,I578067,I578141,);
not I_33859 (I578149,I1804);
not I_33860 (I578166,I2436);
nand I_33861 (I578183,I578166,I578149);
nor I_33862 (I578038,I578141,I578183);
DFFARX1 I_33863 (I578183,I2507,I578067,I578223,);
not I_33864 (I578059,I578223);
not I_33865 (I578245,I1380);
nand I_33866 (I578262,I578166,I578245);
DFFARX1 I_33867 (I578262,I2507,I578067,I578288,);
not I_33868 (I578296,I578288);
not I_33869 (I578313,I1860);
nand I_33870 (I578330,I578313,I1996);
and I_33871 (I578347,I578149,I578330);
nor I_33872 (I578364,I578262,I578347);
DFFARX1 I_33873 (I578364,I2507,I578067,I578035,);
DFFARX1 I_33874 (I578347,I2507,I578067,I578056,);
nor I_33875 (I578409,I1860,I1556);
nor I_33876 (I578047,I578262,I578409);
or I_33877 (I578440,I1860,I1556);
nor I_33878 (I578457,I1812,I2356);
DFFARX1 I_33879 (I578457,I2507,I578067,I578483,);
not I_33880 (I578491,I578483);
nor I_33881 (I578053,I578491,I578296);
nand I_33882 (I578522,I578491,I578141);
not I_33883 (I578539,I1812);
nand I_33884 (I578556,I578539,I578245);
nand I_33885 (I578573,I578491,I578556);
nand I_33886 (I578044,I578573,I578522);
nand I_33887 (I578041,I578556,I578440);
not I_33888 (I578645,I2514);
DFFARX1 I_33889 (I211202,I2507,I578645,I578671,);
and I_33890 (I578679,I578671,I211187);
DFFARX1 I_33891 (I578679,I2507,I578645,I578628,);
DFFARX1 I_33892 (I211193,I2507,I578645,I578719,);
not I_33893 (I578727,I211175);
not I_33894 (I578744,I211196);
nand I_33895 (I578761,I578744,I578727);
nor I_33896 (I578616,I578719,I578761);
DFFARX1 I_33897 (I578761,I2507,I578645,I578801,);
not I_33898 (I578637,I578801);
not I_33899 (I578823,I211199);
nand I_33900 (I578840,I578744,I578823);
DFFARX1 I_33901 (I578840,I2507,I578645,I578866,);
not I_33902 (I578874,I578866);
not I_33903 (I578891,I211190);
nand I_33904 (I578908,I578891,I211178);
and I_33905 (I578925,I578727,I578908);
nor I_33906 (I578942,I578840,I578925);
DFFARX1 I_33907 (I578942,I2507,I578645,I578613,);
DFFARX1 I_33908 (I578925,I2507,I578645,I578634,);
nor I_33909 (I578987,I211190,I211184);
nor I_33910 (I578625,I578840,I578987);
or I_33911 (I579018,I211190,I211184);
nor I_33912 (I579035,I211181,I211175);
DFFARX1 I_33913 (I579035,I2507,I578645,I579061,);
not I_33914 (I579069,I579061);
nor I_33915 (I578631,I579069,I578874);
nand I_33916 (I579100,I579069,I578719);
not I_33917 (I579117,I211181);
nand I_33918 (I579134,I579117,I578823);
nand I_33919 (I579151,I579069,I579134);
nand I_33920 (I578622,I579151,I579100);
nand I_33921 (I578619,I579134,I579018);
not I_33922 (I579223,I2514);
DFFARX1 I_33923 (I1668,I2507,I579223,I579249,);
and I_33924 (I579257,I579249,I2004);
DFFARX1 I_33925 (I579257,I2507,I579223,I579206,);
DFFARX1 I_33926 (I1644,I2507,I579223,I579297,);
not I_33927 (I579305,I2012);
not I_33928 (I579322,I1452);
nand I_33929 (I579339,I579322,I579305);
nor I_33930 (I579194,I579297,I579339);
DFFARX1 I_33931 (I579339,I2507,I579223,I579379,);
not I_33932 (I579215,I579379);
not I_33933 (I579401,I1892);
nand I_33934 (I579418,I579322,I579401);
DFFARX1 I_33935 (I579418,I2507,I579223,I579444,);
not I_33936 (I579452,I579444);
not I_33937 (I579469,I2364);
nand I_33938 (I579486,I579469,I1564);
and I_33939 (I579503,I579305,I579486);
nor I_33940 (I579520,I579418,I579503);
DFFARX1 I_33941 (I579520,I2507,I579223,I579191,);
DFFARX1 I_33942 (I579503,I2507,I579223,I579212,);
nor I_33943 (I579565,I2364,I2060);
nor I_33944 (I579203,I579418,I579565);
or I_33945 (I579596,I2364,I2060);
nor I_33946 (I579613,I1580,I1596);
DFFARX1 I_33947 (I579613,I2507,I579223,I579639,);
not I_33948 (I579647,I579639);
nor I_33949 (I579209,I579647,I579452);
nand I_33950 (I579678,I579647,I579297);
not I_33951 (I579695,I1580);
nand I_33952 (I579712,I579695,I579401);
nand I_33953 (I579729,I579647,I579712);
nand I_33954 (I579200,I579729,I579678);
nand I_33955 (I579197,I579712,I579596);
not I_33956 (I579801,I2514);
DFFARX1 I_33957 (I368644,I2507,I579801,I579827,);
and I_33958 (I579835,I579827,I368632);
DFFARX1 I_33959 (I579835,I2507,I579801,I579784,);
DFFARX1 I_33960 (I368635,I2507,I579801,I579875,);
not I_33961 (I579883,I368629);
not I_33962 (I579900,I368653);
nand I_33963 (I579917,I579900,I579883);
nor I_33964 (I579772,I579875,I579917);
DFFARX1 I_33965 (I579917,I2507,I579801,I579957,);
not I_33966 (I579793,I579957);
not I_33967 (I579979,I368641);
nand I_33968 (I579996,I579900,I579979);
DFFARX1 I_33969 (I579996,I2507,I579801,I580022,);
not I_33970 (I580030,I580022);
not I_33971 (I580047,I368650);
nand I_33972 (I580064,I580047,I368647);
and I_33973 (I580081,I579883,I580064);
nor I_33974 (I580098,I579996,I580081);
DFFARX1 I_33975 (I580098,I2507,I579801,I579769,);
DFFARX1 I_33976 (I580081,I2507,I579801,I579790,);
nor I_33977 (I580143,I368650,I368638);
nor I_33978 (I579781,I579996,I580143);
or I_33979 (I580174,I368650,I368638);
nor I_33980 (I580191,I368629,I368632);
DFFARX1 I_33981 (I580191,I2507,I579801,I580217,);
not I_33982 (I580225,I580217);
nor I_33983 (I579787,I580225,I580030);
nand I_33984 (I580256,I580225,I579875);
not I_33985 (I580273,I368629);
nand I_33986 (I580290,I580273,I579979);
nand I_33987 (I580307,I580225,I580290);
nand I_33988 (I579778,I580307,I580256);
nand I_33989 (I579775,I580290,I580174);
not I_33990 (I580379,I2514);
DFFARX1 I_33991 (I713280,I2507,I580379,I580405,);
and I_33992 (I580413,I580405,I713262);
DFFARX1 I_33993 (I580413,I2507,I580379,I580362,);
DFFARX1 I_33994 (I713253,I2507,I580379,I580453,);
not I_33995 (I580461,I713268);
not I_33996 (I580478,I713256);
nand I_33997 (I580495,I580478,I580461);
nor I_33998 (I580350,I580453,I580495);
DFFARX1 I_33999 (I580495,I2507,I580379,I580535,);
not I_34000 (I580371,I580535);
not I_34001 (I580557,I713265);
nand I_34002 (I580574,I580478,I580557);
DFFARX1 I_34003 (I580574,I2507,I580379,I580600,);
not I_34004 (I580608,I580600);
not I_34005 (I580625,I713274);
nand I_34006 (I580642,I580625,I713253);
and I_34007 (I580659,I580461,I580642);
nor I_34008 (I580676,I580574,I580659);
DFFARX1 I_34009 (I580676,I2507,I580379,I580347,);
DFFARX1 I_34010 (I580659,I2507,I580379,I580368,);
nor I_34011 (I580721,I713274,I713277);
nor I_34012 (I580359,I580574,I580721);
or I_34013 (I580752,I713274,I713277);
nor I_34014 (I580769,I713271,I713259);
DFFARX1 I_34015 (I580769,I2507,I580379,I580795,);
not I_34016 (I580803,I580795);
nor I_34017 (I580365,I580803,I580608);
nand I_34018 (I580834,I580803,I580453);
not I_34019 (I580851,I713271);
nand I_34020 (I580868,I580851,I580557);
nand I_34021 (I580885,I580803,I580868);
nand I_34022 (I580356,I580885,I580834);
nand I_34023 (I580353,I580868,I580752);
not I_34024 (I580957,I2514);
DFFARX1 I_34025 (I723395,I2507,I580957,I580983,);
and I_34026 (I580991,I580983,I723377);
DFFARX1 I_34027 (I580991,I2507,I580957,I580940,);
DFFARX1 I_34028 (I723368,I2507,I580957,I581031,);
not I_34029 (I581039,I723383);
not I_34030 (I581056,I723371);
nand I_34031 (I581073,I581056,I581039);
nor I_34032 (I580928,I581031,I581073);
DFFARX1 I_34033 (I581073,I2507,I580957,I581113,);
not I_34034 (I580949,I581113);
not I_34035 (I581135,I723380);
nand I_34036 (I581152,I581056,I581135);
DFFARX1 I_34037 (I581152,I2507,I580957,I581178,);
not I_34038 (I581186,I581178);
not I_34039 (I581203,I723389);
nand I_34040 (I581220,I581203,I723368);
and I_34041 (I581237,I581039,I581220);
nor I_34042 (I581254,I581152,I581237);
DFFARX1 I_34043 (I581254,I2507,I580957,I580925,);
DFFARX1 I_34044 (I581237,I2507,I580957,I580946,);
nor I_34045 (I581299,I723389,I723392);
nor I_34046 (I580937,I581152,I581299);
or I_34047 (I581330,I723389,I723392);
nor I_34048 (I581347,I723386,I723374);
DFFARX1 I_34049 (I581347,I2507,I580957,I581373,);
not I_34050 (I581381,I581373);
nor I_34051 (I580943,I581381,I581186);
nand I_34052 (I581412,I581381,I581031);
not I_34053 (I581429,I723386);
nand I_34054 (I581446,I581429,I581135);
nand I_34055 (I581463,I581381,I581446);
nand I_34056 (I580934,I581463,I581412);
nand I_34057 (I580931,I581446,I581330);
not I_34058 (I581535,I2514);
DFFARX1 I_34059 (I68365,I2507,I581535,I581561,);
and I_34060 (I581569,I581561,I68341);
DFFARX1 I_34061 (I581569,I2507,I581535,I581518,);
DFFARX1 I_34062 (I68359,I2507,I581535,I581609,);
not I_34063 (I581617,I68347);
not I_34064 (I581634,I68344);
nand I_34065 (I581651,I581634,I581617);
nor I_34066 (I581506,I581609,I581651);
DFFARX1 I_34067 (I581651,I2507,I581535,I581691,);
not I_34068 (I581527,I581691);
not I_34069 (I581713,I68353);
nand I_34070 (I581730,I581634,I581713);
DFFARX1 I_34071 (I581730,I2507,I581535,I581756,);
not I_34072 (I581764,I581756);
not I_34073 (I581781,I68344);
nand I_34074 (I581798,I581781,I68362);
and I_34075 (I581815,I581617,I581798);
nor I_34076 (I581832,I581730,I581815);
DFFARX1 I_34077 (I581832,I2507,I581535,I581503,);
DFFARX1 I_34078 (I581815,I2507,I581535,I581524,);
nor I_34079 (I581877,I68344,I68356);
nor I_34080 (I581515,I581730,I581877);
or I_34081 (I581908,I68344,I68356);
nor I_34082 (I581925,I68350,I68341);
DFFARX1 I_34083 (I581925,I2507,I581535,I581951,);
not I_34084 (I581959,I581951);
nor I_34085 (I581521,I581959,I581764);
nand I_34086 (I581990,I581959,I581609);
not I_34087 (I582007,I68350);
nand I_34088 (I582024,I582007,I581713);
nand I_34089 (I582041,I581959,I582024);
nand I_34090 (I581512,I582041,I581990);
nand I_34091 (I581509,I582024,I581908);
not I_34092 (I582113,I2514);
DFFARX1 I_34093 (I378470,I2507,I582113,I582139,);
and I_34094 (I582147,I582139,I378458);
DFFARX1 I_34095 (I582147,I2507,I582113,I582096,);
DFFARX1 I_34096 (I378461,I2507,I582113,I582187,);
not I_34097 (I582195,I378455);
not I_34098 (I582212,I378479);
nand I_34099 (I582229,I582212,I582195);
nor I_34100 (I582084,I582187,I582229);
DFFARX1 I_34101 (I582229,I2507,I582113,I582269,);
not I_34102 (I582105,I582269);
not I_34103 (I582291,I378467);
nand I_34104 (I582308,I582212,I582291);
DFFARX1 I_34105 (I582308,I2507,I582113,I582334,);
not I_34106 (I582342,I582334);
not I_34107 (I582359,I378476);
nand I_34108 (I582376,I582359,I378473);
and I_34109 (I582393,I582195,I582376);
nor I_34110 (I582410,I582308,I582393);
DFFARX1 I_34111 (I582410,I2507,I582113,I582081,);
DFFARX1 I_34112 (I582393,I2507,I582113,I582102,);
nor I_34113 (I582455,I378476,I378464);
nor I_34114 (I582093,I582308,I582455);
or I_34115 (I582486,I378476,I378464);
nor I_34116 (I582503,I378455,I378458);
DFFARX1 I_34117 (I582503,I2507,I582113,I582529,);
not I_34118 (I582537,I582529);
nor I_34119 (I582099,I582537,I582342);
nand I_34120 (I582568,I582537,I582187);
not I_34121 (I582585,I378455);
nand I_34122 (I582602,I582585,I582291);
nand I_34123 (I582619,I582537,I582602);
nand I_34124 (I582090,I582619,I582568);
nand I_34125 (I582087,I582602,I582486);
not I_34126 (I582691,I2514);
DFFARX1 I_34127 (I420664,I2507,I582691,I582717,);
and I_34128 (I582725,I582717,I420652);
DFFARX1 I_34129 (I582725,I2507,I582691,I582674,);
DFFARX1 I_34130 (I420655,I2507,I582691,I582765,);
not I_34131 (I582773,I420649);
not I_34132 (I582790,I420673);
nand I_34133 (I582807,I582790,I582773);
nor I_34134 (I582662,I582765,I582807);
DFFARX1 I_34135 (I582807,I2507,I582691,I582847,);
not I_34136 (I582683,I582847);
not I_34137 (I582869,I420661);
nand I_34138 (I582886,I582790,I582869);
DFFARX1 I_34139 (I582886,I2507,I582691,I582912,);
not I_34140 (I582920,I582912);
not I_34141 (I582937,I420670);
nand I_34142 (I582954,I582937,I420667);
and I_34143 (I582971,I582773,I582954);
nor I_34144 (I582988,I582886,I582971);
DFFARX1 I_34145 (I582988,I2507,I582691,I582659,);
DFFARX1 I_34146 (I582971,I2507,I582691,I582680,);
nor I_34147 (I583033,I420670,I420658);
nor I_34148 (I582671,I582886,I583033);
or I_34149 (I583064,I420670,I420658);
nor I_34150 (I583081,I420649,I420652);
DFFARX1 I_34151 (I583081,I2507,I582691,I583107,);
not I_34152 (I583115,I583107);
nor I_34153 (I582677,I583115,I582920);
nand I_34154 (I583146,I583115,I582765);
not I_34155 (I583163,I420649);
nand I_34156 (I583180,I583163,I582869);
nand I_34157 (I583197,I583115,I583180);
nand I_34158 (I582668,I583197,I583146);
nand I_34159 (I582665,I583180,I583064);
not I_34160 (I583269,I2514);
DFFARX1 I_34161 (I74689,I2507,I583269,I583295,);
and I_34162 (I583303,I583295,I74665);
DFFARX1 I_34163 (I583303,I2507,I583269,I583252,);
DFFARX1 I_34164 (I74683,I2507,I583269,I583343,);
not I_34165 (I583351,I74671);
not I_34166 (I583368,I74668);
nand I_34167 (I583385,I583368,I583351);
nor I_34168 (I583240,I583343,I583385);
DFFARX1 I_34169 (I583385,I2507,I583269,I583425,);
not I_34170 (I583261,I583425);
not I_34171 (I583447,I74677);
nand I_34172 (I583464,I583368,I583447);
DFFARX1 I_34173 (I583464,I2507,I583269,I583490,);
not I_34174 (I583498,I583490);
not I_34175 (I583515,I74668);
nand I_34176 (I583532,I583515,I74686);
and I_34177 (I583549,I583351,I583532);
nor I_34178 (I583566,I583464,I583549);
DFFARX1 I_34179 (I583566,I2507,I583269,I583237,);
DFFARX1 I_34180 (I583549,I2507,I583269,I583258,);
nor I_34181 (I583611,I74668,I74680);
nor I_34182 (I583249,I583464,I583611);
or I_34183 (I583642,I74668,I74680);
nor I_34184 (I583659,I74674,I74665);
DFFARX1 I_34185 (I583659,I2507,I583269,I583685,);
not I_34186 (I583693,I583685);
nor I_34187 (I583255,I583693,I583498);
nand I_34188 (I583724,I583693,I583343);
not I_34189 (I583741,I74674);
nand I_34190 (I583758,I583741,I583447);
nand I_34191 (I583775,I583693,I583758);
nand I_34192 (I583246,I583775,I583724);
nand I_34193 (I583243,I583758,I583642);
not I_34194 (I583847,I2514);
DFFARX1 I_34195 (I113374,I2507,I583847,I583873,);
and I_34196 (I583881,I583873,I113377);
DFFARX1 I_34197 (I583881,I2507,I583847,I583830,);
DFFARX1 I_34198 (I113377,I2507,I583847,I583921,);
not I_34199 (I583929,I113392);
not I_34200 (I583946,I113398);
nand I_34201 (I583963,I583946,I583929);
nor I_34202 (I583818,I583921,I583963);
DFFARX1 I_34203 (I583963,I2507,I583847,I584003,);
not I_34204 (I583839,I584003);
not I_34205 (I584025,I113386);
nand I_34206 (I584042,I583946,I584025);
DFFARX1 I_34207 (I584042,I2507,I583847,I584068,);
not I_34208 (I584076,I584068);
not I_34209 (I584093,I113383);
nand I_34210 (I584110,I584093,I113380);
and I_34211 (I584127,I583929,I584110);
nor I_34212 (I584144,I584042,I584127);
DFFARX1 I_34213 (I584144,I2507,I583847,I583815,);
DFFARX1 I_34214 (I584127,I2507,I583847,I583836,);
nor I_34215 (I584189,I113383,I113374);
nor I_34216 (I583827,I584042,I584189);
or I_34217 (I584220,I113383,I113374);
nor I_34218 (I584237,I113389,I113395);
DFFARX1 I_34219 (I584237,I2507,I583847,I584263,);
not I_34220 (I584271,I584263);
nor I_34221 (I583833,I584271,I584076);
nand I_34222 (I584302,I584271,I583921);
not I_34223 (I584319,I113389);
nand I_34224 (I584336,I584319,I584025);
nand I_34225 (I584353,I584271,I584336);
nand I_34226 (I583824,I584353,I584302);
nand I_34227 (I583821,I584336,I584220);
not I_34228 (I584425,I2514);
DFFARX1 I_34229 (I721015,I2507,I584425,I584451,);
and I_34230 (I584459,I584451,I720997);
DFFARX1 I_34231 (I584459,I2507,I584425,I584408,);
DFFARX1 I_34232 (I720988,I2507,I584425,I584499,);
not I_34233 (I584507,I721003);
not I_34234 (I584524,I720991);
nand I_34235 (I584541,I584524,I584507);
nor I_34236 (I584396,I584499,I584541);
DFFARX1 I_34237 (I584541,I2507,I584425,I584581,);
not I_34238 (I584417,I584581);
not I_34239 (I584603,I721000);
nand I_34240 (I584620,I584524,I584603);
DFFARX1 I_34241 (I584620,I2507,I584425,I584646,);
not I_34242 (I584654,I584646);
not I_34243 (I584671,I721009);
nand I_34244 (I584688,I584671,I720988);
and I_34245 (I584705,I584507,I584688);
nor I_34246 (I584722,I584620,I584705);
DFFARX1 I_34247 (I584722,I2507,I584425,I584393,);
DFFARX1 I_34248 (I584705,I2507,I584425,I584414,);
nor I_34249 (I584767,I721009,I721012);
nor I_34250 (I584405,I584620,I584767);
or I_34251 (I584798,I721009,I721012);
nor I_34252 (I584815,I721006,I720994);
DFFARX1 I_34253 (I584815,I2507,I584425,I584841,);
not I_34254 (I584849,I584841);
nor I_34255 (I584411,I584849,I584654);
nand I_34256 (I584880,I584849,I584499);
not I_34257 (I584897,I721006);
nand I_34258 (I584914,I584897,I584603);
nand I_34259 (I584931,I584849,I584914);
nand I_34260 (I584402,I584931,I584880);
nand I_34261 (I584399,I584914,I584798);
not I_34262 (I585003,I2514);
DFFARX1 I_34263 (I4317,I2507,I585003,I585029,);
and I_34264 (I585037,I585029,I4323);
DFFARX1 I_34265 (I585037,I2507,I585003,I584986,);
DFFARX1 I_34266 (I4302,I2507,I585003,I585077,);
not I_34267 (I585085,I4308);
not I_34268 (I585102,I4314);
nand I_34269 (I585119,I585102,I585085);
nor I_34270 (I584974,I585077,I585119);
DFFARX1 I_34271 (I585119,I2507,I585003,I585159,);
not I_34272 (I584995,I585159);
not I_34273 (I585181,I4305);
nand I_34274 (I585198,I585102,I585181);
DFFARX1 I_34275 (I585198,I2507,I585003,I585224,);
not I_34276 (I585232,I585224);
not I_34277 (I585249,I4320);
nand I_34278 (I585266,I585249,I4305);
and I_34279 (I585283,I585085,I585266);
nor I_34280 (I585300,I585198,I585283);
DFFARX1 I_34281 (I585300,I2507,I585003,I584971,);
DFFARX1 I_34282 (I585283,I2507,I585003,I584992,);
nor I_34283 (I585345,I4320,I4308);
nor I_34284 (I584983,I585198,I585345);
or I_34285 (I585376,I4320,I4308);
nor I_34286 (I585393,I4311,I4302);
DFFARX1 I_34287 (I585393,I2507,I585003,I585419,);
not I_34288 (I585427,I585419);
nor I_34289 (I584989,I585427,I585232);
nand I_34290 (I585458,I585427,I585077);
not I_34291 (I585475,I4311);
nand I_34292 (I585492,I585475,I585181);
nand I_34293 (I585509,I585427,I585492);
nand I_34294 (I584980,I585509,I585458);
nand I_34295 (I584977,I585492,I585376);
not I_34296 (I585581,I2514);
DFFARX1 I_34297 (I480240,I2507,I585581,I585607,);
and I_34298 (I585615,I585607,I480234);
DFFARX1 I_34299 (I585615,I2507,I585581,I585564,);
DFFARX1 I_34300 (I480252,I2507,I585581,I585655,);
not I_34301 (I585663,I480243);
not I_34302 (I585680,I480255);
nand I_34303 (I585697,I585680,I585663);
nor I_34304 (I585552,I585655,I585697);
DFFARX1 I_34305 (I585697,I2507,I585581,I585737,);
not I_34306 (I585573,I585737);
not I_34307 (I585759,I480261);
nand I_34308 (I585776,I585680,I585759);
DFFARX1 I_34309 (I585776,I2507,I585581,I585802,);
not I_34310 (I585810,I585802);
not I_34311 (I585827,I480237);
nand I_34312 (I585844,I585827,I480258);
and I_34313 (I585861,I585663,I585844);
nor I_34314 (I585878,I585776,I585861);
DFFARX1 I_34315 (I585878,I2507,I585581,I585549,);
DFFARX1 I_34316 (I585861,I2507,I585581,I585570,);
nor I_34317 (I585923,I480237,I480249);
nor I_34318 (I585561,I585776,I585923);
or I_34319 (I585954,I480237,I480249);
nor I_34320 (I585971,I480234,I480246);
DFFARX1 I_34321 (I585971,I2507,I585581,I585997,);
not I_34322 (I586005,I585997);
nor I_34323 (I585567,I586005,I585810);
nand I_34324 (I586036,I586005,I585655);
not I_34325 (I586053,I480234);
nand I_34326 (I586070,I586053,I585759);
nand I_34327 (I586087,I586005,I586070);
nand I_34328 (I585558,I586087,I586036);
nand I_34329 (I585555,I586070,I585954);
not I_34330 (I586159,I2514);
DFFARX1 I_34331 (I30397,I2507,I586159,I586185,);
and I_34332 (I586193,I586185,I30400);
DFFARX1 I_34333 (I586193,I2507,I586159,I586142,);
DFFARX1 I_34334 (I30400,I2507,I586159,I586233,);
not I_34335 (I586241,I30403);
not I_34336 (I586258,I30418);
nand I_34337 (I586275,I586258,I586241);
nor I_34338 (I586130,I586233,I586275);
DFFARX1 I_34339 (I586275,I2507,I586159,I586315,);
not I_34340 (I586151,I586315);
not I_34341 (I586337,I30412);
nand I_34342 (I586354,I586258,I586337);
DFFARX1 I_34343 (I586354,I2507,I586159,I586380,);
not I_34344 (I586388,I586380);
not I_34345 (I586405,I30415);
nand I_34346 (I586422,I586405,I30397);
and I_34347 (I586439,I586241,I586422);
nor I_34348 (I586456,I586354,I586439);
DFFARX1 I_34349 (I586456,I2507,I586159,I586127,);
DFFARX1 I_34350 (I586439,I2507,I586159,I586148,);
nor I_34351 (I586501,I30415,I30409);
nor I_34352 (I586139,I586354,I586501);
or I_34353 (I586532,I30415,I30409);
nor I_34354 (I586549,I30406,I30421);
DFFARX1 I_34355 (I586549,I2507,I586159,I586575,);
not I_34356 (I586583,I586575);
nor I_34357 (I586145,I586583,I586388);
nand I_34358 (I586614,I586583,I586233);
not I_34359 (I586631,I30406);
nand I_34360 (I586648,I586631,I586337);
nand I_34361 (I586665,I586583,I586648);
nand I_34362 (I586136,I586665,I586614);
nand I_34363 (I586133,I586648,I586532);
not I_34364 (I586737,I2514);
DFFARX1 I_34365 (I230776,I2507,I586737,I586763,);
and I_34366 (I586771,I586763,I230791);
DFFARX1 I_34367 (I586771,I2507,I586737,I586720,);
DFFARX1 I_34368 (I230794,I2507,I586737,I586811,);
not I_34369 (I586819,I230788);
not I_34370 (I586836,I230803);
nand I_34371 (I586853,I586836,I586819);
nor I_34372 (I586708,I586811,I586853);
DFFARX1 I_34373 (I586853,I2507,I586737,I586893,);
not I_34374 (I586729,I586893);
not I_34375 (I586915,I230779);
nand I_34376 (I586932,I586836,I586915);
DFFARX1 I_34377 (I586932,I2507,I586737,I586958,);
not I_34378 (I586966,I586958);
not I_34379 (I586983,I230782);
nand I_34380 (I587000,I586983,I230776);
and I_34381 (I587017,I586819,I587000);
nor I_34382 (I587034,I586932,I587017);
DFFARX1 I_34383 (I587034,I2507,I586737,I586705,);
DFFARX1 I_34384 (I587017,I2507,I586737,I586726,);
nor I_34385 (I587079,I230782,I230785);
nor I_34386 (I586717,I586932,I587079);
or I_34387 (I587110,I230782,I230785);
nor I_34388 (I587127,I230800,I230797);
DFFARX1 I_34389 (I587127,I2507,I586737,I587153,);
not I_34390 (I587161,I587153);
nor I_34391 (I586723,I587161,I586966);
nand I_34392 (I587192,I587161,I586811);
not I_34393 (I587209,I230800);
nand I_34394 (I587226,I587209,I586915);
nand I_34395 (I587243,I587161,I587226);
nand I_34396 (I586714,I587243,I587192);
nand I_34397 (I586711,I587226,I587110);
not I_34398 (I587315,I2514);
DFFARX1 I_34399 (I223323,I2507,I587315,I587341,);
and I_34400 (I587349,I587341,I223308);
DFFARX1 I_34401 (I587349,I2507,I587315,I587298,);
DFFARX1 I_34402 (I223314,I2507,I587315,I587389,);
not I_34403 (I587397,I223296);
not I_34404 (I587414,I223317);
nand I_34405 (I587431,I587414,I587397);
nor I_34406 (I587286,I587389,I587431);
DFFARX1 I_34407 (I587431,I2507,I587315,I587471,);
not I_34408 (I587307,I587471);
not I_34409 (I587493,I223320);
nand I_34410 (I587510,I587414,I587493);
DFFARX1 I_34411 (I587510,I2507,I587315,I587536,);
not I_34412 (I587544,I587536);
not I_34413 (I587561,I223311);
nand I_34414 (I587578,I587561,I223299);
and I_34415 (I587595,I587397,I587578);
nor I_34416 (I587612,I587510,I587595);
DFFARX1 I_34417 (I587612,I2507,I587315,I587283,);
DFFARX1 I_34418 (I587595,I2507,I587315,I587304,);
nor I_34419 (I587657,I223311,I223305);
nor I_34420 (I587295,I587510,I587657);
or I_34421 (I587688,I223311,I223305);
nor I_34422 (I587705,I223302,I223296);
DFFARX1 I_34423 (I587705,I2507,I587315,I587731,);
not I_34424 (I587739,I587731);
nor I_34425 (I587301,I587739,I587544);
nand I_34426 (I587770,I587739,I587389);
not I_34427 (I587787,I223302);
nand I_34428 (I587804,I587787,I587493);
nand I_34429 (I587821,I587739,I587804);
nand I_34430 (I587292,I587821,I587770);
nand I_34431 (I587289,I587804,I587688);
not I_34432 (I587893,I2514);
DFFARX1 I_34433 (I659962,I2507,I587893,I587919,);
and I_34434 (I587927,I587919,I659956);
DFFARX1 I_34435 (I587927,I2507,I587893,I587876,);
DFFARX1 I_34436 (I659941,I2507,I587893,I587967,);
not I_34437 (I587975,I659947);
not I_34438 (I587992,I659959);
nand I_34439 (I588009,I587992,I587975);
nor I_34440 (I587864,I587967,I588009);
DFFARX1 I_34441 (I588009,I2507,I587893,I588049,);
not I_34442 (I587885,I588049);
not I_34443 (I588071,I659941);
nand I_34444 (I588088,I587992,I588071);
DFFARX1 I_34445 (I588088,I2507,I587893,I588114,);
not I_34446 (I588122,I588114);
not I_34447 (I588139,I659965);
nand I_34448 (I588156,I588139,I659953);
and I_34449 (I588173,I587975,I588156);
nor I_34450 (I588190,I588088,I588173);
DFFARX1 I_34451 (I588190,I2507,I587893,I587861,);
DFFARX1 I_34452 (I588173,I2507,I587893,I587882,);
nor I_34453 (I588235,I659965,I659944);
nor I_34454 (I587873,I588088,I588235);
or I_34455 (I588266,I659965,I659944);
nor I_34456 (I588283,I659950,I659944);
DFFARX1 I_34457 (I588283,I2507,I587893,I588309,);
not I_34458 (I588317,I588309);
nor I_34459 (I587879,I588317,I588122);
nand I_34460 (I588348,I588317,I587967);
not I_34461 (I588365,I659950);
nand I_34462 (I588382,I588365,I588071);
nand I_34463 (I588399,I588317,I588382);
nand I_34464 (I587870,I588399,I588348);
nand I_34465 (I587867,I588382,I588266);
not I_34466 (I588471,I2514);
DFFARX1 I_34467 (I2492,I2507,I588471,I588497,);
and I_34468 (I588505,I588497,I2276);
DFFARX1 I_34469 (I588505,I2507,I588471,I588454,);
DFFARX1 I_34470 (I2140,I2507,I588471,I588545,);
not I_34471 (I588553,I1900);
not I_34472 (I588570,I1372);
nand I_34473 (I588587,I588570,I588553);
nor I_34474 (I588442,I588545,I588587);
DFFARX1 I_34475 (I588587,I2507,I588471,I588627,);
not I_34476 (I588463,I588627);
not I_34477 (I588649,I1484);
nand I_34478 (I588666,I588570,I588649);
DFFARX1 I_34479 (I588666,I2507,I588471,I588692,);
not I_34480 (I588700,I588692);
not I_34481 (I588717,I1708);
nand I_34482 (I588734,I588717,I2220);
and I_34483 (I588751,I588553,I588734);
nor I_34484 (I588768,I588666,I588751);
DFFARX1 I_34485 (I588768,I2507,I588471,I588439,);
DFFARX1 I_34486 (I588751,I2507,I588471,I588460,);
nor I_34487 (I588813,I1708,I2084);
nor I_34488 (I588451,I588666,I588813);
or I_34489 (I588844,I1708,I2084);
nor I_34490 (I588861,I1748,I1500);
DFFARX1 I_34491 (I588861,I2507,I588471,I588887,);
not I_34492 (I588895,I588887);
nor I_34493 (I588457,I588895,I588700);
nand I_34494 (I588926,I588895,I588545);
not I_34495 (I588943,I1748);
nand I_34496 (I588960,I588943,I588649);
nand I_34497 (I588977,I588895,I588960);
nand I_34498 (I588448,I588977,I588926);
nand I_34499 (I588445,I588960,I588844);
not I_34500 (I589049,I2514);
DFFARX1 I_34501 (I253080,I2507,I589049,I589075,);
and I_34502 (I589083,I589075,I253095);
DFFARX1 I_34503 (I589083,I2507,I589049,I589032,);
DFFARX1 I_34504 (I253098,I2507,I589049,I589123,);
not I_34505 (I589131,I253092);
not I_34506 (I589148,I253107);
nand I_34507 (I589165,I589148,I589131);
nor I_34508 (I589020,I589123,I589165);
DFFARX1 I_34509 (I589165,I2507,I589049,I589205,);
not I_34510 (I589041,I589205);
not I_34511 (I589227,I253083);
nand I_34512 (I589244,I589148,I589227);
DFFARX1 I_34513 (I589244,I2507,I589049,I589270,);
not I_34514 (I589278,I589270);
not I_34515 (I589295,I253086);
nand I_34516 (I589312,I589295,I253080);
and I_34517 (I589329,I589131,I589312);
nor I_34518 (I589346,I589244,I589329);
DFFARX1 I_34519 (I589346,I2507,I589049,I589017,);
DFFARX1 I_34520 (I589329,I2507,I589049,I589038,);
nor I_34521 (I589391,I253086,I253089);
nor I_34522 (I589029,I589244,I589391);
or I_34523 (I589422,I253086,I253089);
nor I_34524 (I589439,I253104,I253101);
DFFARX1 I_34525 (I589439,I2507,I589049,I589465,);
not I_34526 (I589473,I589465);
nor I_34527 (I589035,I589473,I589278);
nand I_34528 (I589504,I589473,I589123);
not I_34529 (I589521,I253104);
nand I_34530 (I589538,I589521,I589227);
nand I_34531 (I589555,I589473,I589538);
nand I_34532 (I589026,I589555,I589504);
nand I_34533 (I589023,I589538,I589422);
not I_34534 (I589627,I2514);
DFFARX1 I_34535 (I52028,I2507,I589627,I589653,);
and I_34536 (I589661,I589653,I52004);
DFFARX1 I_34537 (I589661,I2507,I589627,I589610,);
DFFARX1 I_34538 (I52022,I2507,I589627,I589701,);
not I_34539 (I589709,I52010);
not I_34540 (I589726,I52007);
nand I_34541 (I589743,I589726,I589709);
nor I_34542 (I589598,I589701,I589743);
DFFARX1 I_34543 (I589743,I2507,I589627,I589783,);
not I_34544 (I589619,I589783);
not I_34545 (I589805,I52016);
nand I_34546 (I589822,I589726,I589805);
DFFARX1 I_34547 (I589822,I2507,I589627,I589848,);
not I_34548 (I589856,I589848);
not I_34549 (I589873,I52007);
nand I_34550 (I589890,I589873,I52025);
and I_34551 (I589907,I589709,I589890);
nor I_34552 (I589924,I589822,I589907);
DFFARX1 I_34553 (I589924,I2507,I589627,I589595,);
DFFARX1 I_34554 (I589907,I2507,I589627,I589616,);
nor I_34555 (I589969,I52007,I52019);
nor I_34556 (I589607,I589822,I589969);
or I_34557 (I590000,I52007,I52019);
nor I_34558 (I590017,I52013,I52004);
DFFARX1 I_34559 (I590017,I2507,I589627,I590043,);
not I_34560 (I590051,I590043);
nor I_34561 (I589613,I590051,I589856);
nand I_34562 (I590082,I590051,I589701);
not I_34563 (I590099,I52013);
nand I_34564 (I590116,I590099,I589805);
nand I_34565 (I590133,I590051,I590116);
nand I_34566 (I589604,I590133,I590082);
nand I_34567 (I589601,I590116,I590000);
not I_34568 (I590205,I2514);
DFFARX1 I_34569 (I334542,I2507,I590205,I590231,);
and I_34570 (I590239,I590231,I334530);
DFFARX1 I_34571 (I590239,I2507,I590205,I590188,);
DFFARX1 I_34572 (I334545,I2507,I590205,I590279,);
not I_34573 (I590287,I334536);
not I_34574 (I590304,I334527);
nand I_34575 (I590321,I590304,I590287);
nor I_34576 (I590176,I590279,I590321);
DFFARX1 I_34577 (I590321,I2507,I590205,I590361,);
not I_34578 (I590197,I590361);
not I_34579 (I590383,I334533);
nand I_34580 (I590400,I590304,I590383);
DFFARX1 I_34581 (I590400,I2507,I590205,I590426,);
not I_34582 (I590434,I590426);
not I_34583 (I590451,I334548);
nand I_34584 (I590468,I590451,I334551);
and I_34585 (I590485,I590287,I590468);
nor I_34586 (I590502,I590400,I590485);
DFFARX1 I_34587 (I590502,I2507,I590205,I590173,);
DFFARX1 I_34588 (I590485,I2507,I590205,I590194,);
nor I_34589 (I590547,I334548,I334527);
nor I_34590 (I590185,I590400,I590547);
or I_34591 (I590578,I334548,I334527);
nor I_34592 (I590595,I334539,I334530);
DFFARX1 I_34593 (I590595,I2507,I590205,I590621,);
not I_34594 (I590629,I590621);
nor I_34595 (I590191,I590629,I590434);
nand I_34596 (I590660,I590629,I590279);
not I_34597 (I590677,I334539);
nand I_34598 (I590694,I590677,I590383);
nand I_34599 (I590711,I590629,I590694);
nand I_34600 (I590182,I590711,I590660);
nand I_34601 (I590179,I590694,I590578);
not I_34602 (I590783,I2514);
DFFARX1 I_34603 (I729345,I2507,I590783,I590809,);
and I_34604 (I590817,I590809,I729327);
DFFARX1 I_34605 (I590817,I2507,I590783,I590766,);
DFFARX1 I_34606 (I729318,I2507,I590783,I590857,);
not I_34607 (I590865,I729333);
not I_34608 (I590882,I729321);
nand I_34609 (I590899,I590882,I590865);
nor I_34610 (I590754,I590857,I590899);
DFFARX1 I_34611 (I590899,I2507,I590783,I590939,);
not I_34612 (I590775,I590939);
not I_34613 (I590961,I729330);
nand I_34614 (I590978,I590882,I590961);
DFFARX1 I_34615 (I590978,I2507,I590783,I591004,);
not I_34616 (I591012,I591004);
not I_34617 (I591029,I729339);
nand I_34618 (I591046,I591029,I729318);
and I_34619 (I591063,I590865,I591046);
nor I_34620 (I591080,I590978,I591063);
DFFARX1 I_34621 (I591080,I2507,I590783,I590751,);
DFFARX1 I_34622 (I591063,I2507,I590783,I590772,);
nor I_34623 (I591125,I729339,I729342);
nor I_34624 (I590763,I590978,I591125);
or I_34625 (I591156,I729339,I729342);
nor I_34626 (I591173,I729336,I729324);
DFFARX1 I_34627 (I591173,I2507,I590783,I591199,);
not I_34628 (I591207,I591199);
nor I_34629 (I590769,I591207,I591012);
nand I_34630 (I591238,I591207,I590857);
not I_34631 (I591255,I729336);
nand I_34632 (I591272,I591255,I590961);
nand I_34633 (I591289,I591207,I591272);
nand I_34634 (I590760,I591289,I591238);
nand I_34635 (I590757,I591272,I591156);
not I_34636 (I591361,I2514);
DFFARX1 I_34637 (I696620,I2507,I591361,I591387,);
and I_34638 (I591395,I591387,I696602);
DFFARX1 I_34639 (I591395,I2507,I591361,I591344,);
DFFARX1 I_34640 (I696593,I2507,I591361,I591435,);
not I_34641 (I591443,I696608);
not I_34642 (I591460,I696596);
nand I_34643 (I591477,I591460,I591443);
nor I_34644 (I591332,I591435,I591477);
DFFARX1 I_34645 (I591477,I2507,I591361,I591517,);
not I_34646 (I591353,I591517);
not I_34647 (I591539,I696605);
nand I_34648 (I591556,I591460,I591539);
DFFARX1 I_34649 (I591556,I2507,I591361,I591582,);
not I_34650 (I591590,I591582);
not I_34651 (I591607,I696614);
nand I_34652 (I591624,I591607,I696593);
and I_34653 (I591641,I591443,I591624);
nor I_34654 (I591658,I591556,I591641);
DFFARX1 I_34655 (I591658,I2507,I591361,I591329,);
DFFARX1 I_34656 (I591641,I2507,I591361,I591350,);
nor I_34657 (I591703,I696614,I696617);
nor I_34658 (I591341,I591556,I591703);
or I_34659 (I591734,I696614,I696617);
nor I_34660 (I591751,I696611,I696599);
DFFARX1 I_34661 (I591751,I2507,I591361,I591777,);
not I_34662 (I591785,I591777);
nor I_34663 (I591347,I591785,I591590);
nand I_34664 (I591816,I591785,I591435);
not I_34665 (I591833,I696611);
nand I_34666 (I591850,I591833,I591539);
nand I_34667 (I591867,I591785,I591850);
nand I_34668 (I591338,I591867,I591816);
nand I_34669 (I591335,I591850,I591734);
not I_34670 (I591939,I2514);
DFFARX1 I_34671 (I148479,I2507,I591939,I591965,);
and I_34672 (I591973,I591965,I148482);
DFFARX1 I_34673 (I591973,I2507,I591939,I591922,);
DFFARX1 I_34674 (I148482,I2507,I591939,I592013,);
not I_34675 (I592021,I148497);
not I_34676 (I592038,I148503);
nand I_34677 (I592055,I592038,I592021);
nor I_34678 (I591910,I592013,I592055);
DFFARX1 I_34679 (I592055,I2507,I591939,I592095,);
not I_34680 (I591931,I592095);
not I_34681 (I592117,I148491);
nand I_34682 (I592134,I592038,I592117);
DFFARX1 I_34683 (I592134,I2507,I591939,I592160,);
not I_34684 (I592168,I592160);
not I_34685 (I592185,I148488);
nand I_34686 (I592202,I592185,I148485);
and I_34687 (I592219,I592021,I592202);
nor I_34688 (I592236,I592134,I592219);
DFFARX1 I_34689 (I592236,I2507,I591939,I591907,);
DFFARX1 I_34690 (I592219,I2507,I591939,I591928,);
nor I_34691 (I592281,I148488,I148479);
nor I_34692 (I591919,I592134,I592281);
or I_34693 (I592312,I148488,I148479);
nor I_34694 (I592329,I148494,I148500);
DFFARX1 I_34695 (I592329,I2507,I591939,I592355,);
not I_34696 (I592363,I592355);
nor I_34697 (I591925,I592363,I592168);
nand I_34698 (I592394,I592363,I592013);
not I_34699 (I592411,I148494);
nand I_34700 (I592428,I592411,I592117);
nand I_34701 (I592445,I592363,I592428);
nand I_34702 (I591916,I592445,I592394);
nand I_34703 (I591913,I592428,I592312);
not I_34704 (I592517,I2514);
DFFARX1 I_34705 (I24073,I2507,I592517,I592543,);
and I_34706 (I592551,I592543,I24076);
DFFARX1 I_34707 (I592551,I2507,I592517,I592500,);
DFFARX1 I_34708 (I24076,I2507,I592517,I592591,);
not I_34709 (I592599,I24079);
not I_34710 (I592616,I24094);
nand I_34711 (I592633,I592616,I592599);
nor I_34712 (I592488,I592591,I592633);
DFFARX1 I_34713 (I592633,I2507,I592517,I592673,);
not I_34714 (I592509,I592673);
not I_34715 (I592695,I24088);
nand I_34716 (I592712,I592616,I592695);
DFFARX1 I_34717 (I592712,I2507,I592517,I592738,);
not I_34718 (I592746,I592738);
not I_34719 (I592763,I24091);
nand I_34720 (I592780,I592763,I24073);
and I_34721 (I592797,I592599,I592780);
nor I_34722 (I592814,I592712,I592797);
DFFARX1 I_34723 (I592814,I2507,I592517,I592485,);
DFFARX1 I_34724 (I592797,I2507,I592517,I592506,);
nor I_34725 (I592859,I24091,I24085);
nor I_34726 (I592497,I592712,I592859);
or I_34727 (I592890,I24091,I24085);
nor I_34728 (I592907,I24082,I24097);
DFFARX1 I_34729 (I592907,I2507,I592517,I592933,);
not I_34730 (I592941,I592933);
nor I_34731 (I592503,I592941,I592746);
nand I_34732 (I592972,I592941,I592591);
not I_34733 (I592989,I24082);
nand I_34734 (I593006,I592989,I592695);
nand I_34735 (I593023,I592941,I593006);
nand I_34736 (I592494,I593023,I592972);
nand I_34737 (I592491,I593006,I592890);
not I_34738 (I593095,I2514);
DFFARX1 I_34739 (I463424,I2507,I593095,I593121,);
and I_34740 (I593129,I593121,I463430);
DFFARX1 I_34741 (I593129,I2507,I593095,I593078,);
DFFARX1 I_34742 (I463436,I2507,I593095,I593169,);
not I_34743 (I593177,I463421);
not I_34744 (I593194,I463421);
nand I_34745 (I593211,I593194,I593177);
nor I_34746 (I593066,I593169,I593211);
DFFARX1 I_34747 (I593211,I2507,I593095,I593251,);
not I_34748 (I593087,I593251);
not I_34749 (I593273,I463439);
nand I_34750 (I593290,I593194,I593273);
DFFARX1 I_34751 (I593290,I2507,I593095,I593316,);
not I_34752 (I593324,I593316);
not I_34753 (I593341,I463433);
nand I_34754 (I593358,I593341,I463424);
and I_34755 (I593375,I593177,I593358);
nor I_34756 (I593392,I593290,I593375);
DFFARX1 I_34757 (I593392,I2507,I593095,I593063,);
DFFARX1 I_34758 (I593375,I2507,I593095,I593084,);
nor I_34759 (I593437,I463433,I463442);
nor I_34760 (I593075,I593290,I593437);
or I_34761 (I593468,I463433,I463442);
nor I_34762 (I593485,I463427,I463427);
DFFARX1 I_34763 (I593485,I2507,I593095,I593511,);
not I_34764 (I593519,I593511);
nor I_34765 (I593081,I593519,I593324);
nand I_34766 (I593550,I593519,I593169);
not I_34767 (I593567,I463427);
nand I_34768 (I593584,I593567,I593273);
nand I_34769 (I593601,I593519,I593584);
nand I_34770 (I593072,I593601,I593550);
nand I_34771 (I593069,I593584,I593468);
not I_34772 (I593673,I2514);
DFFARX1 I_34773 (I167461,I2507,I593673,I593699,);
and I_34774 (I593707,I593699,I167446);
DFFARX1 I_34775 (I593707,I2507,I593673,I593656,);
DFFARX1 I_34776 (I167452,I2507,I593673,I593747,);
not I_34777 (I593755,I167434);
not I_34778 (I593772,I167455);
nand I_34779 (I593789,I593772,I593755);
nor I_34780 (I593644,I593747,I593789);
DFFARX1 I_34781 (I593789,I2507,I593673,I593829,);
not I_34782 (I593665,I593829);
not I_34783 (I593851,I167458);
nand I_34784 (I593868,I593772,I593851);
DFFARX1 I_34785 (I593868,I2507,I593673,I593894,);
not I_34786 (I593902,I593894);
not I_34787 (I593919,I167449);
nand I_34788 (I593936,I593919,I167437);
and I_34789 (I593953,I593755,I593936);
nor I_34790 (I593970,I593868,I593953);
DFFARX1 I_34791 (I593970,I2507,I593673,I593641,);
DFFARX1 I_34792 (I593953,I2507,I593673,I593662,);
nor I_34793 (I594015,I167449,I167443);
nor I_34794 (I593653,I593868,I594015);
or I_34795 (I594046,I167449,I167443);
nor I_34796 (I594063,I167440,I167434);
DFFARX1 I_34797 (I594063,I2507,I593673,I594089,);
not I_34798 (I594097,I594089);
nor I_34799 (I593659,I594097,I593902);
nand I_34800 (I594128,I594097,I593747);
not I_34801 (I594145,I167440);
nand I_34802 (I594162,I594145,I593851);
nand I_34803 (I594179,I594097,I594162);
nand I_34804 (I593650,I594179,I594128);
nand I_34805 (I593647,I594162,I594046);
not I_34806 (I594251,I2514);
DFFARX1 I_34807 (I325294,I2507,I594251,I594277,);
and I_34808 (I594285,I594277,I325282);
DFFARX1 I_34809 (I594285,I2507,I594251,I594234,);
DFFARX1 I_34810 (I325297,I2507,I594251,I594325,);
not I_34811 (I594333,I325288);
not I_34812 (I594350,I325279);
nand I_34813 (I594367,I594350,I594333);
nor I_34814 (I594222,I594325,I594367);
DFFARX1 I_34815 (I594367,I2507,I594251,I594407,);
not I_34816 (I594243,I594407);
not I_34817 (I594429,I325285);
nand I_34818 (I594446,I594350,I594429);
DFFARX1 I_34819 (I594446,I2507,I594251,I594472,);
not I_34820 (I594480,I594472);
not I_34821 (I594497,I325300);
nand I_34822 (I594514,I594497,I325303);
and I_34823 (I594531,I594333,I594514);
nor I_34824 (I594548,I594446,I594531);
DFFARX1 I_34825 (I594548,I2507,I594251,I594219,);
DFFARX1 I_34826 (I594531,I2507,I594251,I594240,);
nor I_34827 (I594593,I325300,I325279);
nor I_34828 (I594231,I594446,I594593);
or I_34829 (I594624,I325300,I325279);
nor I_34830 (I594641,I325291,I325282);
DFFARX1 I_34831 (I594641,I2507,I594251,I594667,);
not I_34832 (I594675,I594667);
nor I_34833 (I594237,I594675,I594480);
nand I_34834 (I594706,I594675,I594325);
not I_34835 (I594723,I325291);
nand I_34836 (I594740,I594723,I594429);
nand I_34837 (I594757,I594675,I594740);
nand I_34838 (I594228,I594757,I594706);
nand I_34839 (I594225,I594740,I594624);
not I_34840 (I594829,I2514);
DFFARX1 I_34841 (I135389,I2507,I594829,I594855,);
and I_34842 (I594863,I594855,I135392);
DFFARX1 I_34843 (I594863,I2507,I594829,I594812,);
DFFARX1 I_34844 (I135392,I2507,I594829,I594903,);
not I_34845 (I594911,I135407);
not I_34846 (I594928,I135413);
nand I_34847 (I594945,I594928,I594911);
nor I_34848 (I594800,I594903,I594945);
DFFARX1 I_34849 (I594945,I2507,I594829,I594985,);
not I_34850 (I594821,I594985);
not I_34851 (I595007,I135401);
nand I_34852 (I595024,I594928,I595007);
DFFARX1 I_34853 (I595024,I2507,I594829,I595050,);
not I_34854 (I595058,I595050);
not I_34855 (I595075,I135398);
nand I_34856 (I595092,I595075,I135395);
and I_34857 (I595109,I594911,I595092);
nor I_34858 (I595126,I595024,I595109);
DFFARX1 I_34859 (I595126,I2507,I594829,I594797,);
DFFARX1 I_34860 (I595109,I2507,I594829,I594818,);
nor I_34861 (I595171,I135398,I135389);
nor I_34862 (I594809,I595024,I595171);
or I_34863 (I595202,I135398,I135389);
nor I_34864 (I595219,I135404,I135410);
DFFARX1 I_34865 (I595219,I2507,I594829,I595245,);
not I_34866 (I595253,I595245);
nor I_34867 (I594815,I595253,I595058);
nand I_34868 (I595284,I595253,I594903);
not I_34869 (I595301,I135404);
nand I_34870 (I595318,I595301,I595007);
nand I_34871 (I595335,I595253,I595318);
nand I_34872 (I594806,I595335,I595284);
nand I_34873 (I594803,I595318,I595202);
not I_34874 (I595407,I2514);
DFFARX1 I_34875 (I103259,I2507,I595407,I595433,);
and I_34876 (I595441,I595433,I103262);
DFFARX1 I_34877 (I595441,I2507,I595407,I595390,);
DFFARX1 I_34878 (I103262,I2507,I595407,I595481,);
not I_34879 (I595489,I103277);
not I_34880 (I595506,I103283);
nand I_34881 (I595523,I595506,I595489);
nor I_34882 (I595378,I595481,I595523);
DFFARX1 I_34883 (I595523,I2507,I595407,I595563,);
not I_34884 (I595399,I595563);
not I_34885 (I595585,I103271);
nand I_34886 (I595602,I595506,I595585);
DFFARX1 I_34887 (I595602,I2507,I595407,I595628,);
not I_34888 (I595636,I595628);
not I_34889 (I595653,I103268);
nand I_34890 (I595670,I595653,I103265);
and I_34891 (I595687,I595489,I595670);
nor I_34892 (I595704,I595602,I595687);
DFFARX1 I_34893 (I595704,I2507,I595407,I595375,);
DFFARX1 I_34894 (I595687,I2507,I595407,I595396,);
nor I_34895 (I595749,I103268,I103259);
nor I_34896 (I595387,I595602,I595749);
or I_34897 (I595780,I103268,I103259);
nor I_34898 (I595797,I103274,I103280);
DFFARX1 I_34899 (I595797,I2507,I595407,I595823,);
not I_34900 (I595831,I595823);
nor I_34901 (I595393,I595831,I595636);
nand I_34902 (I595862,I595831,I595481);
not I_34903 (I595879,I103274);
nand I_34904 (I595896,I595879,I595585);
nand I_34905 (I595913,I595831,I595896);
nand I_34906 (I595384,I595913,I595862);
nand I_34907 (I595381,I595896,I595780);
not I_34908 (I595985,I2514);
DFFARX1 I_34909 (I246552,I2507,I595985,I596011,);
and I_34910 (I596019,I596011,I246567);
DFFARX1 I_34911 (I596019,I2507,I595985,I595968,);
DFFARX1 I_34912 (I246570,I2507,I595985,I596059,);
not I_34913 (I596067,I246564);
not I_34914 (I596084,I246579);
nand I_34915 (I596101,I596084,I596067);
nor I_34916 (I595956,I596059,I596101);
DFFARX1 I_34917 (I596101,I2507,I595985,I596141,);
not I_34918 (I595977,I596141);
not I_34919 (I596163,I246555);
nand I_34920 (I596180,I596084,I596163);
DFFARX1 I_34921 (I596180,I2507,I595985,I596206,);
not I_34922 (I596214,I596206);
not I_34923 (I596231,I246558);
nand I_34924 (I596248,I596231,I246552);
and I_34925 (I596265,I596067,I596248);
nor I_34926 (I596282,I596180,I596265);
DFFARX1 I_34927 (I596282,I2507,I595985,I595953,);
DFFARX1 I_34928 (I596265,I2507,I595985,I595974,);
nor I_34929 (I596327,I246558,I246561);
nor I_34930 (I595965,I596180,I596327);
or I_34931 (I596358,I246558,I246561);
nor I_34932 (I596375,I246576,I246573);
DFFARX1 I_34933 (I596375,I2507,I595985,I596401,);
not I_34934 (I596409,I596401);
nor I_34935 (I595971,I596409,I596214);
nand I_34936 (I596440,I596409,I596059);
not I_34937 (I596457,I246576);
nand I_34938 (I596474,I596457,I596163);
nand I_34939 (I596491,I596409,I596474);
nand I_34940 (I595962,I596491,I596440);
nand I_34941 (I595959,I596474,I596358);
not I_34942 (I596563,I2514);
DFFARX1 I_34943 (I310844,I2507,I596563,I596589,);
and I_34944 (I596597,I596589,I310832);
DFFARX1 I_34945 (I596597,I2507,I596563,I596546,);
DFFARX1 I_34946 (I310847,I2507,I596563,I596637,);
not I_34947 (I596645,I310838);
not I_34948 (I596662,I310829);
nand I_34949 (I596679,I596662,I596645);
nor I_34950 (I596534,I596637,I596679);
DFFARX1 I_34951 (I596679,I2507,I596563,I596719,);
not I_34952 (I596555,I596719);
not I_34953 (I596741,I310835);
nand I_34954 (I596758,I596662,I596741);
DFFARX1 I_34955 (I596758,I2507,I596563,I596784,);
not I_34956 (I596792,I596784);
not I_34957 (I596809,I310850);
nand I_34958 (I596826,I596809,I310853);
and I_34959 (I596843,I596645,I596826);
nor I_34960 (I596860,I596758,I596843);
DFFARX1 I_34961 (I596860,I2507,I596563,I596531,);
DFFARX1 I_34962 (I596843,I2507,I596563,I596552,);
nor I_34963 (I596905,I310850,I310829);
nor I_34964 (I596543,I596758,I596905);
or I_34965 (I596936,I310850,I310829);
nor I_34966 (I596953,I310841,I310832);
DFFARX1 I_34967 (I596953,I2507,I596563,I596979,);
not I_34968 (I596987,I596979);
nor I_34969 (I596549,I596987,I596792);
nand I_34970 (I597018,I596987,I596637);
not I_34971 (I597035,I310841);
nand I_34972 (I597052,I597035,I596741);
nand I_34973 (I597069,I596987,I597052);
nand I_34974 (I596540,I597069,I597018);
nand I_34975 (I596537,I597052,I596936);
not I_34976 (I597141,I2514);
DFFARX1 I_34977 (I411994,I2507,I597141,I597167,);
and I_34978 (I597175,I597167,I411982);
DFFARX1 I_34979 (I597175,I2507,I597141,I597124,);
DFFARX1 I_34980 (I411985,I2507,I597141,I597215,);
not I_34981 (I597223,I411979);
not I_34982 (I597240,I412003);
nand I_34983 (I597257,I597240,I597223);
nor I_34984 (I597112,I597215,I597257);
DFFARX1 I_34985 (I597257,I2507,I597141,I597297,);
not I_34986 (I597133,I597297);
not I_34987 (I597319,I411991);
nand I_34988 (I597336,I597240,I597319);
DFFARX1 I_34989 (I597336,I2507,I597141,I597362,);
not I_34990 (I597370,I597362);
not I_34991 (I597387,I412000);
nand I_34992 (I597404,I597387,I411997);
and I_34993 (I597421,I597223,I597404);
nor I_34994 (I597438,I597336,I597421);
DFFARX1 I_34995 (I597438,I2507,I597141,I597109,);
DFFARX1 I_34996 (I597421,I2507,I597141,I597130,);
nor I_34997 (I597483,I412000,I411988);
nor I_34998 (I597121,I597336,I597483);
or I_34999 (I597514,I412000,I411988);
nor I_35000 (I597531,I411979,I411982);
DFFARX1 I_35001 (I597531,I2507,I597141,I597557,);
not I_35002 (I597565,I597557);
nor I_35003 (I597127,I597565,I597370);
nand I_35004 (I597596,I597565,I597215);
not I_35005 (I597613,I411979);
nand I_35006 (I597630,I597613,I597319);
nand I_35007 (I597647,I597565,I597630);
nand I_35008 (I597118,I597647,I597596);
nand I_35009 (I597115,I597630,I597514);
not I_35010 (I597719,I2514);
DFFARX1 I_35011 (I197500,I2507,I597719,I597745,);
and I_35012 (I597753,I597745,I197485);
DFFARX1 I_35013 (I597753,I2507,I597719,I597702,);
DFFARX1 I_35014 (I197491,I2507,I597719,I597793,);
not I_35015 (I597801,I197473);
not I_35016 (I597818,I197494);
nand I_35017 (I597835,I597818,I597801);
nor I_35018 (I597690,I597793,I597835);
DFFARX1 I_35019 (I597835,I2507,I597719,I597875,);
not I_35020 (I597711,I597875);
not I_35021 (I597897,I197497);
nand I_35022 (I597914,I597818,I597897);
DFFARX1 I_35023 (I597914,I2507,I597719,I597940,);
not I_35024 (I597948,I597940);
not I_35025 (I597965,I197488);
nand I_35026 (I597982,I597965,I197476);
and I_35027 (I597999,I597801,I597982);
nor I_35028 (I598016,I597914,I597999);
DFFARX1 I_35029 (I598016,I2507,I597719,I597687,);
DFFARX1 I_35030 (I597999,I2507,I597719,I597708,);
nor I_35031 (I598061,I197488,I197482);
nor I_35032 (I597699,I597914,I598061);
or I_35033 (I598092,I197488,I197482);
nor I_35034 (I598109,I197479,I197473);
DFFARX1 I_35035 (I598109,I2507,I597719,I598135,);
not I_35036 (I598143,I598135);
nor I_35037 (I597705,I598143,I597948);
nand I_35038 (I598174,I598143,I597793);
not I_35039 (I598191,I197479);
nand I_35040 (I598208,I598191,I597897);
nand I_35041 (I598225,I598143,I598208);
nand I_35042 (I597696,I598225,I598174);
nand I_35043 (I597693,I598208,I598092);
not I_35044 (I598297,I2514);
DFFARX1 I_35045 (I279192,I2507,I598297,I598323,);
and I_35046 (I598331,I598323,I279207);
DFFARX1 I_35047 (I598331,I2507,I598297,I598280,);
DFFARX1 I_35048 (I279210,I2507,I598297,I598371,);
not I_35049 (I598379,I279204);
not I_35050 (I598396,I279219);
nand I_35051 (I598413,I598396,I598379);
nor I_35052 (I598268,I598371,I598413);
DFFARX1 I_35053 (I598413,I2507,I598297,I598453,);
not I_35054 (I598289,I598453);
not I_35055 (I598475,I279195);
nand I_35056 (I598492,I598396,I598475);
DFFARX1 I_35057 (I598492,I2507,I598297,I598518,);
not I_35058 (I598526,I598518);
not I_35059 (I598543,I279198);
nand I_35060 (I598560,I598543,I279192);
and I_35061 (I598577,I598379,I598560);
nor I_35062 (I598594,I598492,I598577);
DFFARX1 I_35063 (I598594,I2507,I598297,I598265,);
DFFARX1 I_35064 (I598577,I2507,I598297,I598286,);
nor I_35065 (I598639,I279198,I279201);
nor I_35066 (I598277,I598492,I598639);
or I_35067 (I598670,I279198,I279201);
nor I_35068 (I598687,I279216,I279213);
DFFARX1 I_35069 (I598687,I2507,I598297,I598713,);
not I_35070 (I598721,I598713);
nor I_35071 (I598283,I598721,I598526);
nand I_35072 (I598752,I598721,I598371);
not I_35073 (I598769,I279216);
nand I_35074 (I598786,I598769,I598475);
nand I_35075 (I598803,I598721,I598786);
nand I_35076 (I598274,I598803,I598752);
nand I_35077 (I598271,I598786,I598670);
not I_35078 (I598875,I2514);
DFFARX1 I_35079 (I335698,I2507,I598875,I598901,);
and I_35080 (I598909,I598901,I335686);
DFFARX1 I_35081 (I598909,I2507,I598875,I598858,);
DFFARX1 I_35082 (I335701,I2507,I598875,I598949,);
not I_35083 (I598957,I335692);
not I_35084 (I598974,I335683);
nand I_35085 (I598991,I598974,I598957);
nor I_35086 (I598846,I598949,I598991);
DFFARX1 I_35087 (I598991,I2507,I598875,I599031,);
not I_35088 (I598867,I599031);
not I_35089 (I599053,I335689);
nand I_35090 (I599070,I598974,I599053);
DFFARX1 I_35091 (I599070,I2507,I598875,I599096,);
not I_35092 (I599104,I599096);
not I_35093 (I599121,I335704);
nand I_35094 (I599138,I599121,I335707);
and I_35095 (I599155,I598957,I599138);
nor I_35096 (I599172,I599070,I599155);
DFFARX1 I_35097 (I599172,I2507,I598875,I598843,);
DFFARX1 I_35098 (I599155,I2507,I598875,I598864,);
nor I_35099 (I599217,I335704,I335683);
nor I_35100 (I598855,I599070,I599217);
or I_35101 (I599248,I335704,I335683);
nor I_35102 (I599265,I335695,I335686);
DFFARX1 I_35103 (I599265,I2507,I598875,I599291,);
not I_35104 (I599299,I599291);
nor I_35105 (I598861,I599299,I599104);
nand I_35106 (I599330,I599299,I598949);
not I_35107 (I599347,I335695);
nand I_35108 (I599364,I599347,I599053);
nand I_35109 (I599381,I599299,I599364);
nand I_35110 (I598852,I599381,I599330);
nand I_35111 (I598849,I599364,I599248);
not I_35112 (I599453,I2514);
DFFARX1 I_35113 (I439709,I2507,I599453,I599479,);
and I_35114 (I599487,I599479,I439715);
DFFARX1 I_35115 (I599487,I2507,I599453,I599436,);
DFFARX1 I_35116 (I439721,I2507,I599453,I599527,);
not I_35117 (I599535,I439706);
not I_35118 (I599552,I439706);
nand I_35119 (I599569,I599552,I599535);
nor I_35120 (I599424,I599527,I599569);
DFFARX1 I_35121 (I599569,I2507,I599453,I599609,);
not I_35122 (I599445,I599609);
not I_35123 (I599631,I439724);
nand I_35124 (I599648,I599552,I599631);
DFFARX1 I_35125 (I599648,I2507,I599453,I599674,);
not I_35126 (I599682,I599674);
not I_35127 (I599699,I439718);
nand I_35128 (I599716,I599699,I439709);
and I_35129 (I599733,I599535,I599716);
nor I_35130 (I599750,I599648,I599733);
DFFARX1 I_35131 (I599750,I2507,I599453,I599421,);
DFFARX1 I_35132 (I599733,I2507,I599453,I599442,);
nor I_35133 (I599795,I439718,I439727);
nor I_35134 (I599433,I599648,I599795);
or I_35135 (I599826,I439718,I439727);
nor I_35136 (I599843,I439712,I439712);
DFFARX1 I_35137 (I599843,I2507,I599453,I599869,);
not I_35138 (I599877,I599869);
nor I_35139 (I599439,I599877,I599682);
nand I_35140 (I599908,I599877,I599527);
not I_35141 (I599925,I439712);
nand I_35142 (I599942,I599925,I599631);
nand I_35143 (I599959,I599877,I599942);
nand I_35144 (I599430,I599959,I599908);
nand I_35145 (I599427,I599942,I599826);
not I_35146 (I600031,I2514);
DFFARX1 I_35147 (I88384,I2507,I600031,I600057,);
and I_35148 (I600065,I600057,I88387);
DFFARX1 I_35149 (I600065,I2507,I600031,I600014,);
DFFARX1 I_35150 (I88387,I2507,I600031,I600105,);
not I_35151 (I600113,I88402);
not I_35152 (I600130,I88408);
nand I_35153 (I600147,I600130,I600113);
nor I_35154 (I600002,I600105,I600147);
DFFARX1 I_35155 (I600147,I2507,I600031,I600187,);
not I_35156 (I600023,I600187);
not I_35157 (I600209,I88396);
nand I_35158 (I600226,I600130,I600209);
DFFARX1 I_35159 (I600226,I2507,I600031,I600252,);
not I_35160 (I600260,I600252);
not I_35161 (I600277,I88393);
nand I_35162 (I600294,I600277,I88390);
and I_35163 (I600311,I600113,I600294);
nor I_35164 (I600328,I600226,I600311);
DFFARX1 I_35165 (I600328,I2507,I600031,I599999,);
DFFARX1 I_35166 (I600311,I2507,I600031,I600020,);
nor I_35167 (I600373,I88393,I88384);
nor I_35168 (I600011,I600226,I600373);
or I_35169 (I600404,I88393,I88384);
nor I_35170 (I600421,I88399,I88405);
DFFARX1 I_35171 (I600421,I2507,I600031,I600447,);
not I_35172 (I600455,I600447);
nor I_35173 (I600017,I600455,I600260);
nand I_35174 (I600486,I600455,I600105);
not I_35175 (I600503,I88399);
nand I_35176 (I600520,I600503,I600209);
nand I_35177 (I600537,I600455,I600520);
nand I_35178 (I600008,I600537,I600486);
nand I_35179 (I600005,I600520,I600404);
not I_35180 (I600609,I2514);
DFFARX1 I_35181 (I434966,I2507,I600609,I600635,);
and I_35182 (I600643,I600635,I434972);
DFFARX1 I_35183 (I600643,I2507,I600609,I600592,);
DFFARX1 I_35184 (I434978,I2507,I600609,I600683,);
not I_35185 (I600691,I434963);
not I_35186 (I600708,I434963);
nand I_35187 (I600725,I600708,I600691);
nor I_35188 (I600580,I600683,I600725);
DFFARX1 I_35189 (I600725,I2507,I600609,I600765,);
not I_35190 (I600601,I600765);
not I_35191 (I600787,I434981);
nand I_35192 (I600804,I600708,I600787);
DFFARX1 I_35193 (I600804,I2507,I600609,I600830,);
not I_35194 (I600838,I600830);
not I_35195 (I600855,I434975);
nand I_35196 (I600872,I600855,I434966);
and I_35197 (I600889,I600691,I600872);
nor I_35198 (I600906,I600804,I600889);
DFFARX1 I_35199 (I600906,I2507,I600609,I600577,);
DFFARX1 I_35200 (I600889,I2507,I600609,I600598,);
nor I_35201 (I600951,I434975,I434984);
nor I_35202 (I600589,I600804,I600951);
or I_35203 (I600982,I434975,I434984);
nor I_35204 (I600999,I434969,I434969);
DFFARX1 I_35205 (I600999,I2507,I600609,I601025,);
not I_35206 (I601033,I601025);
nor I_35207 (I600595,I601033,I600838);
nand I_35208 (I601064,I601033,I600683);
not I_35209 (I601081,I434969);
nand I_35210 (I601098,I601081,I600787);
nand I_35211 (I601115,I601033,I601098);
nand I_35212 (I600586,I601115,I601064);
nand I_35213 (I600583,I601098,I600982);
not I_35214 (I601187,I2514);
DFFARX1 I_35215 (I655066,I2507,I601187,I601213,);
and I_35216 (I601221,I601213,I655060);
DFFARX1 I_35217 (I601221,I2507,I601187,I601170,);
DFFARX1 I_35218 (I655045,I2507,I601187,I601261,);
not I_35219 (I601269,I655051);
not I_35220 (I601286,I655063);
nand I_35221 (I601303,I601286,I601269);
nor I_35222 (I601158,I601261,I601303);
DFFARX1 I_35223 (I601303,I2507,I601187,I601343,);
not I_35224 (I601179,I601343);
not I_35225 (I601365,I655045);
nand I_35226 (I601382,I601286,I601365);
DFFARX1 I_35227 (I601382,I2507,I601187,I601408,);
not I_35228 (I601416,I601408);
not I_35229 (I601433,I655069);
nand I_35230 (I601450,I601433,I655057);
and I_35231 (I601467,I601269,I601450);
nor I_35232 (I601484,I601382,I601467);
DFFARX1 I_35233 (I601484,I2507,I601187,I601155,);
DFFARX1 I_35234 (I601467,I2507,I601187,I601176,);
nor I_35235 (I601529,I655069,I655048);
nor I_35236 (I601167,I601382,I601529);
or I_35237 (I601560,I655069,I655048);
nor I_35238 (I601577,I655054,I655048);
DFFARX1 I_35239 (I601577,I2507,I601187,I601603,);
not I_35240 (I601611,I601603);
nor I_35241 (I601173,I601611,I601416);
nand I_35242 (I601642,I601611,I601261);
not I_35243 (I601659,I655054);
nand I_35244 (I601676,I601659,I601365);
nand I_35245 (I601693,I601611,I601676);
nand I_35246 (I601164,I601693,I601642);
nand I_35247 (I601161,I601676,I601560);
not I_35248 (I601765,I2514);
DFFARX1 I_35249 (I87789,I2507,I601765,I601791,);
and I_35250 (I601799,I601791,I87813);
DFFARX1 I_35251 (I601799,I2507,I601765,I601748,);
DFFARX1 I_35252 (I87789,I2507,I601765,I601839,);
not I_35253 (I601847,I87807);
not I_35254 (I601864,I87792);
nand I_35255 (I601881,I601864,I601847);
nor I_35256 (I601736,I601839,I601881);
DFFARX1 I_35257 (I601881,I2507,I601765,I601921,);
not I_35258 (I601757,I601921);
not I_35259 (I601943,I87801);
nand I_35260 (I601960,I601864,I601943);
DFFARX1 I_35261 (I601960,I2507,I601765,I601986,);
not I_35262 (I601994,I601986);
not I_35263 (I602011,I87798);
nand I_35264 (I602028,I602011,I87795);
and I_35265 (I602045,I601847,I602028);
nor I_35266 (I602062,I601960,I602045);
DFFARX1 I_35267 (I602062,I2507,I601765,I601733,);
DFFARX1 I_35268 (I602045,I2507,I601765,I601754,);
nor I_35269 (I602107,I87798,I87804);
nor I_35270 (I601745,I601960,I602107);
or I_35271 (I602138,I87798,I87804);
nor I_35272 (I602155,I87810,I87816);
DFFARX1 I_35273 (I602155,I2507,I601765,I602181,);
not I_35274 (I602189,I602181);
nor I_35275 (I601751,I602189,I601994);
nand I_35276 (I602220,I602189,I601839);
not I_35277 (I602237,I87810);
nand I_35278 (I602254,I602237,I601943);
nand I_35279 (I602271,I602189,I602254);
nand I_35280 (I601742,I602271,I602220);
nand I_35281 (I601739,I602254,I602138);
not I_35282 (I602343,I2514);
DFFARX1 I_35283 (I404480,I2507,I602343,I602369,);
and I_35284 (I602377,I602369,I404468);
DFFARX1 I_35285 (I602377,I2507,I602343,I602326,);
DFFARX1 I_35286 (I404471,I2507,I602343,I602417,);
not I_35287 (I602425,I404465);
not I_35288 (I602442,I404489);
nand I_35289 (I602459,I602442,I602425);
nor I_35290 (I602314,I602417,I602459);
DFFARX1 I_35291 (I602459,I2507,I602343,I602499,);
not I_35292 (I602335,I602499);
not I_35293 (I602521,I404477);
nand I_35294 (I602538,I602442,I602521);
DFFARX1 I_35295 (I602538,I2507,I602343,I602564,);
not I_35296 (I602572,I602564);
not I_35297 (I602589,I404486);
nand I_35298 (I602606,I602589,I404483);
and I_35299 (I602623,I602425,I602606);
nor I_35300 (I602640,I602538,I602623);
DFFARX1 I_35301 (I602640,I2507,I602343,I602311,);
DFFARX1 I_35302 (I602623,I2507,I602343,I602332,);
nor I_35303 (I602685,I404486,I404474);
nor I_35304 (I602323,I602538,I602685);
or I_35305 (I602716,I404486,I404474);
nor I_35306 (I602733,I404465,I404468);
DFFARX1 I_35307 (I602733,I2507,I602343,I602759,);
not I_35308 (I602767,I602759);
nor I_35309 (I602329,I602767,I602572);
nand I_35310 (I602798,I602767,I602417);
not I_35311 (I602815,I404465);
nand I_35312 (I602832,I602815,I602521);
nand I_35313 (I602849,I602767,I602832);
nand I_35314 (I602320,I602849,I602798);
nand I_35315 (I602317,I602832,I602716);
not I_35316 (I602921,I2514);
DFFARX1 I_35317 (I557621,I2507,I602921,I602947,);
and I_35318 (I602955,I602947,I557618);
DFFARX1 I_35319 (I602955,I2507,I602921,I602904,);
DFFARX1 I_35320 (I557624,I2507,I602921,I602995,);
not I_35321 (I603003,I557627);
not I_35322 (I603020,I557621);
nand I_35323 (I603037,I603020,I603003);
nor I_35324 (I602892,I602995,I603037);
DFFARX1 I_35325 (I603037,I2507,I602921,I603077,);
not I_35326 (I602913,I603077);
not I_35327 (I603099,I557636);
nand I_35328 (I603116,I603020,I603099);
DFFARX1 I_35329 (I603116,I2507,I602921,I603142,);
not I_35330 (I603150,I603142);
not I_35331 (I603167,I557633);
nand I_35332 (I603184,I603167,I557639);
and I_35333 (I603201,I603003,I603184);
nor I_35334 (I603218,I603116,I603201);
DFFARX1 I_35335 (I603218,I2507,I602921,I602889,);
DFFARX1 I_35336 (I603201,I2507,I602921,I602910,);
nor I_35337 (I603263,I557633,I557618);
nor I_35338 (I602901,I603116,I603263);
or I_35339 (I603294,I557633,I557618);
nor I_35340 (I603311,I557630,I557624);
DFFARX1 I_35341 (I603311,I2507,I602921,I603337,);
not I_35342 (I603345,I603337);
nor I_35343 (I602907,I603345,I603150);
nand I_35344 (I603376,I603345,I602995);
not I_35345 (I603393,I557630);
nand I_35346 (I603410,I603393,I603099);
nand I_35347 (I603427,I603345,I603410);
nand I_35348 (I602898,I603427,I603376);
nand I_35349 (I602895,I603410,I603294);
not I_35350 (I603499,I2514);
DFFARX1 I_35351 (I696025,I2507,I603499,I603525,);
and I_35352 (I603533,I603525,I696007);
DFFARX1 I_35353 (I603533,I2507,I603499,I603482,);
DFFARX1 I_35354 (I695998,I2507,I603499,I603573,);
not I_35355 (I603581,I696013);
not I_35356 (I603598,I696001);
nand I_35357 (I603615,I603598,I603581);
nor I_35358 (I603470,I603573,I603615);
DFFARX1 I_35359 (I603615,I2507,I603499,I603655,);
not I_35360 (I603491,I603655);
not I_35361 (I603677,I696010);
nand I_35362 (I603694,I603598,I603677);
DFFARX1 I_35363 (I603694,I2507,I603499,I603720,);
not I_35364 (I603728,I603720);
not I_35365 (I603745,I696019);
nand I_35366 (I603762,I603745,I695998);
and I_35367 (I603779,I603581,I603762);
nor I_35368 (I603796,I603694,I603779);
DFFARX1 I_35369 (I603796,I2507,I603499,I603467,);
DFFARX1 I_35370 (I603779,I2507,I603499,I603488,);
nor I_35371 (I603841,I696019,I696022);
nor I_35372 (I603479,I603694,I603841);
or I_35373 (I603872,I696019,I696022);
nor I_35374 (I603889,I696016,I696004);
DFFARX1 I_35375 (I603889,I2507,I603499,I603915,);
not I_35376 (I603923,I603915);
nor I_35377 (I603485,I603923,I603728);
nand I_35378 (I603954,I603923,I603573);
not I_35379 (I603971,I696016);
nand I_35380 (I603988,I603971,I603677);
nand I_35381 (I604005,I603923,I603988);
nand I_35382 (I603476,I604005,I603954);
nand I_35383 (I603473,I603988,I603872);
not I_35384 (I604077,I2514);
DFFARX1 I_35385 (I339744,I2507,I604077,I604103,);
and I_35386 (I604111,I604103,I339732);
DFFARX1 I_35387 (I604111,I2507,I604077,I604060,);
DFFARX1 I_35388 (I339747,I2507,I604077,I604151,);
not I_35389 (I604159,I339738);
not I_35390 (I604176,I339729);
nand I_35391 (I604193,I604176,I604159);
nor I_35392 (I604048,I604151,I604193);
DFFARX1 I_35393 (I604193,I2507,I604077,I604233,);
not I_35394 (I604069,I604233);
not I_35395 (I604255,I339735);
nand I_35396 (I604272,I604176,I604255);
DFFARX1 I_35397 (I604272,I2507,I604077,I604298,);
not I_35398 (I604306,I604298);
not I_35399 (I604323,I339750);
nand I_35400 (I604340,I604323,I339753);
and I_35401 (I604357,I604159,I604340);
nor I_35402 (I604374,I604272,I604357);
DFFARX1 I_35403 (I604374,I2507,I604077,I604045,);
DFFARX1 I_35404 (I604357,I2507,I604077,I604066,);
nor I_35405 (I604419,I339750,I339729);
nor I_35406 (I604057,I604272,I604419);
or I_35407 (I604450,I339750,I339729);
nor I_35408 (I604467,I339741,I339732);
DFFARX1 I_35409 (I604467,I2507,I604077,I604493,);
not I_35410 (I604501,I604493);
nor I_35411 (I604063,I604501,I604306);
nand I_35412 (I604532,I604501,I604151);
not I_35413 (I604549,I339741);
nand I_35414 (I604566,I604549,I604255);
nand I_35415 (I604583,I604501,I604566);
nand I_35416 (I604054,I604583,I604532);
nand I_35417 (I604051,I604566,I604450);
not I_35418 (I604655,I2514);
DFFARX1 I_35419 (I308532,I2507,I604655,I604681,);
and I_35420 (I604689,I604681,I308520);
DFFARX1 I_35421 (I604689,I2507,I604655,I604638,);
DFFARX1 I_35422 (I308535,I2507,I604655,I604729,);
not I_35423 (I604737,I308526);
not I_35424 (I604754,I308517);
nand I_35425 (I604771,I604754,I604737);
nor I_35426 (I604626,I604729,I604771);
DFFARX1 I_35427 (I604771,I2507,I604655,I604811,);
not I_35428 (I604647,I604811);
not I_35429 (I604833,I308523);
nand I_35430 (I604850,I604754,I604833);
DFFARX1 I_35431 (I604850,I2507,I604655,I604876,);
not I_35432 (I604884,I604876);
not I_35433 (I604901,I308538);
nand I_35434 (I604918,I604901,I308541);
and I_35435 (I604935,I604737,I604918);
nor I_35436 (I604952,I604850,I604935);
DFFARX1 I_35437 (I604952,I2507,I604655,I604623,);
DFFARX1 I_35438 (I604935,I2507,I604655,I604644,);
nor I_35439 (I604997,I308538,I308517);
nor I_35440 (I604635,I604850,I604997);
or I_35441 (I605028,I308538,I308517);
nor I_35442 (I605045,I308529,I308520);
DFFARX1 I_35443 (I605045,I2507,I604655,I605071,);
not I_35444 (I605079,I605071);
nor I_35445 (I604641,I605079,I604884);
nand I_35446 (I605110,I605079,I604729);
not I_35447 (I605127,I308529);
nand I_35448 (I605144,I605127,I604833);
nand I_35449 (I605161,I605079,I605144);
nand I_35450 (I604632,I605161,I605110);
nand I_35451 (I604629,I605144,I605028);
not I_35452 (I605233,I2514);
DFFARX1 I_35453 (I269400,I2507,I605233,I605259,);
and I_35454 (I605267,I605259,I269415);
DFFARX1 I_35455 (I605267,I2507,I605233,I605216,);
DFFARX1 I_35456 (I269418,I2507,I605233,I605307,);
not I_35457 (I605315,I269412);
not I_35458 (I605332,I269427);
nand I_35459 (I605349,I605332,I605315);
nor I_35460 (I605204,I605307,I605349);
DFFARX1 I_35461 (I605349,I2507,I605233,I605389,);
not I_35462 (I605225,I605389);
not I_35463 (I605411,I269403);
nand I_35464 (I605428,I605332,I605411);
DFFARX1 I_35465 (I605428,I2507,I605233,I605454,);
not I_35466 (I605462,I605454);
not I_35467 (I605479,I269406);
nand I_35468 (I605496,I605479,I269400);
and I_35469 (I605513,I605315,I605496);
nor I_35470 (I605530,I605428,I605513);
DFFARX1 I_35471 (I605530,I2507,I605233,I605201,);
DFFARX1 I_35472 (I605513,I2507,I605233,I605222,);
nor I_35473 (I605575,I269406,I269409);
nor I_35474 (I605213,I605428,I605575);
or I_35475 (I605606,I269406,I269409);
nor I_35476 (I605623,I269424,I269421);
DFFARX1 I_35477 (I605623,I2507,I605233,I605649,);
not I_35478 (I605657,I605649);
nor I_35479 (I605219,I605657,I605462);
nand I_35480 (I605688,I605657,I605307);
not I_35481 (I605705,I269424);
nand I_35482 (I605722,I605705,I605411);
nand I_35483 (I605739,I605657,I605722);
nand I_35484 (I605210,I605739,I605688);
nand I_35485 (I605207,I605722,I605606);
not I_35486 (I605811,I2514);
DFFARX1 I_35487 (I493806,I2507,I605811,I605837,);
and I_35488 (I605845,I605837,I493800);
DFFARX1 I_35489 (I605845,I2507,I605811,I605794,);
DFFARX1 I_35490 (I493818,I2507,I605811,I605885,);
not I_35491 (I605893,I493809);
not I_35492 (I605910,I493821);
nand I_35493 (I605927,I605910,I605893);
nor I_35494 (I605782,I605885,I605927);
DFFARX1 I_35495 (I605927,I2507,I605811,I605967,);
not I_35496 (I605803,I605967);
not I_35497 (I605989,I493827);
nand I_35498 (I606006,I605910,I605989);
DFFARX1 I_35499 (I606006,I2507,I605811,I606032,);
not I_35500 (I606040,I606032);
not I_35501 (I606057,I493803);
nand I_35502 (I606074,I606057,I493824);
and I_35503 (I606091,I605893,I606074);
nor I_35504 (I606108,I606006,I606091);
DFFARX1 I_35505 (I606108,I2507,I605811,I605779,);
DFFARX1 I_35506 (I606091,I2507,I605811,I605800,);
nor I_35507 (I606153,I493803,I493815);
nor I_35508 (I605791,I606006,I606153);
or I_35509 (I606184,I493803,I493815);
nor I_35510 (I606201,I493800,I493812);
DFFARX1 I_35511 (I606201,I2507,I605811,I606227,);
not I_35512 (I606235,I606227);
nor I_35513 (I605797,I606235,I606040);
nand I_35514 (I606266,I606235,I605885);
not I_35515 (I606283,I493800);
nand I_35516 (I606300,I606283,I605989);
nand I_35517 (I606317,I606235,I606300);
nand I_35518 (I605788,I606317,I606266);
nand I_35519 (I605785,I606300,I606184);
not I_35520 (I606389,I2514);
DFFARX1 I_35521 (I665402,I2507,I606389,I606415,);
and I_35522 (I606423,I606415,I665396);
DFFARX1 I_35523 (I606423,I2507,I606389,I606372,);
DFFARX1 I_35524 (I665381,I2507,I606389,I606463,);
not I_35525 (I606471,I665387);
not I_35526 (I606488,I665399);
nand I_35527 (I606505,I606488,I606471);
nor I_35528 (I606360,I606463,I606505);
DFFARX1 I_35529 (I606505,I2507,I606389,I606545,);
not I_35530 (I606381,I606545);
not I_35531 (I606567,I665381);
nand I_35532 (I606584,I606488,I606567);
DFFARX1 I_35533 (I606584,I2507,I606389,I606610,);
not I_35534 (I606618,I606610);
not I_35535 (I606635,I665405);
nand I_35536 (I606652,I606635,I665393);
and I_35537 (I606669,I606471,I606652);
nor I_35538 (I606686,I606584,I606669);
DFFARX1 I_35539 (I606686,I2507,I606389,I606357,);
DFFARX1 I_35540 (I606669,I2507,I606389,I606378,);
nor I_35541 (I606731,I665405,I665384);
nor I_35542 (I606369,I606584,I606731);
or I_35543 (I606762,I665405,I665384);
nor I_35544 (I606779,I665390,I665384);
DFFARX1 I_35545 (I606779,I2507,I606389,I606805,);
not I_35546 (I606813,I606805);
nor I_35547 (I606375,I606813,I606618);
nand I_35548 (I606844,I606813,I606463);
not I_35549 (I606861,I665390);
nand I_35550 (I606878,I606861,I606567);
nand I_35551 (I606895,I606813,I606878);
nand I_35552 (I606366,I606895,I606844);
nand I_35553 (I606363,I606878,I606762);
not I_35554 (I606967,I2514);
DFFARX1 I_35555 (I522230,I2507,I606967,I606993,);
and I_35556 (I607001,I606993,I522224);
DFFARX1 I_35557 (I607001,I2507,I606967,I606950,);
DFFARX1 I_35558 (I522242,I2507,I606967,I607041,);
not I_35559 (I607049,I522233);
not I_35560 (I607066,I522245);
nand I_35561 (I607083,I607066,I607049);
nor I_35562 (I606938,I607041,I607083);
DFFARX1 I_35563 (I607083,I2507,I606967,I607123,);
not I_35564 (I606959,I607123);
not I_35565 (I607145,I522251);
nand I_35566 (I607162,I607066,I607145);
DFFARX1 I_35567 (I607162,I2507,I606967,I607188,);
not I_35568 (I607196,I607188);
not I_35569 (I607213,I522227);
nand I_35570 (I607230,I607213,I522248);
and I_35571 (I607247,I607049,I607230);
nor I_35572 (I607264,I607162,I607247);
DFFARX1 I_35573 (I607264,I2507,I606967,I606935,);
DFFARX1 I_35574 (I607247,I2507,I606967,I606956,);
nor I_35575 (I607309,I522227,I522239);
nor I_35576 (I606947,I607162,I607309);
or I_35577 (I607340,I522227,I522239);
nor I_35578 (I607357,I522224,I522236);
DFFARX1 I_35579 (I607357,I2507,I606967,I607383,);
not I_35580 (I607391,I607383);
nor I_35581 (I606953,I607391,I607196);
nand I_35582 (I607422,I607391,I607041);
not I_35583 (I607439,I522224);
nand I_35584 (I607456,I607439,I607145);
nand I_35585 (I607473,I607391,I607456);
nand I_35586 (I606944,I607473,I607422);
nand I_35587 (I606941,I607456,I607340);
not I_35588 (I607545,I2514);
DFFARX1 I_35589 (I134794,I2507,I607545,I607571,);
and I_35590 (I607579,I607571,I134797);
DFFARX1 I_35591 (I607579,I2507,I607545,I607528,);
DFFARX1 I_35592 (I134797,I2507,I607545,I607619,);
not I_35593 (I607627,I134812);
not I_35594 (I607644,I134818);
nand I_35595 (I607661,I607644,I607627);
nor I_35596 (I607516,I607619,I607661);
DFFARX1 I_35597 (I607661,I2507,I607545,I607701,);
not I_35598 (I607537,I607701);
not I_35599 (I607723,I134806);
nand I_35600 (I607740,I607644,I607723);
DFFARX1 I_35601 (I607740,I2507,I607545,I607766,);
not I_35602 (I607774,I607766);
not I_35603 (I607791,I134803);
nand I_35604 (I607808,I607791,I134800);
and I_35605 (I607825,I607627,I607808);
nor I_35606 (I607842,I607740,I607825);
DFFARX1 I_35607 (I607842,I2507,I607545,I607513,);
DFFARX1 I_35608 (I607825,I2507,I607545,I607534,);
nor I_35609 (I607887,I134803,I134794);
nor I_35610 (I607525,I607740,I607887);
or I_35611 (I607918,I134803,I134794);
nor I_35612 (I607935,I134809,I134815);
DFFARX1 I_35613 (I607935,I2507,I607545,I607961,);
not I_35614 (I607969,I607961);
nor I_35615 (I607531,I607969,I607774);
nand I_35616 (I608000,I607969,I607619);
not I_35617 (I608017,I134809);
nand I_35618 (I608034,I608017,I607723);
nand I_35619 (I608051,I607969,I608034);
nand I_35620 (I607522,I608051,I608000);
nand I_35621 (I607519,I608034,I607918);
not I_35622 (I608123,I2514);
DFFARX1 I_35623 (I229144,I2507,I608123,I608149,);
and I_35624 (I608157,I608149,I229159);
DFFARX1 I_35625 (I608157,I2507,I608123,I608106,);
DFFARX1 I_35626 (I229162,I2507,I608123,I608197,);
not I_35627 (I608205,I229156);
not I_35628 (I608222,I229171);
nand I_35629 (I608239,I608222,I608205);
nor I_35630 (I608094,I608197,I608239);
DFFARX1 I_35631 (I608239,I2507,I608123,I608279,);
not I_35632 (I608115,I608279);
not I_35633 (I608301,I229147);
nand I_35634 (I608318,I608222,I608301);
DFFARX1 I_35635 (I608318,I2507,I608123,I608344,);
not I_35636 (I608352,I608344);
not I_35637 (I608369,I229150);
nand I_35638 (I608386,I608369,I229144);
and I_35639 (I608403,I608205,I608386);
nor I_35640 (I608420,I608318,I608403);
DFFARX1 I_35641 (I608420,I2507,I608123,I608091,);
DFFARX1 I_35642 (I608403,I2507,I608123,I608112,);
nor I_35643 (I608465,I229150,I229153);
nor I_35644 (I608103,I608318,I608465);
or I_35645 (I608496,I229150,I229153);
nor I_35646 (I608513,I229168,I229165);
DFFARX1 I_35647 (I608513,I2507,I608123,I608539,);
not I_35648 (I608547,I608539);
nor I_35649 (I608109,I608547,I608352);
nand I_35650 (I608578,I608547,I608197);
not I_35651 (I608595,I229168);
nand I_35652 (I608612,I608595,I608301);
nand I_35653 (I608629,I608547,I608612);
nand I_35654 (I608100,I608629,I608578);
nand I_35655 (I608097,I608612,I608496);
not I_35656 (I608701,I2514);
DFFARX1 I_35657 (I473964,I2507,I608701,I608727,);
and I_35658 (I608735,I608727,I473970);
DFFARX1 I_35659 (I608735,I2507,I608701,I608684,);
DFFARX1 I_35660 (I473976,I2507,I608701,I608775,);
not I_35661 (I608783,I473961);
not I_35662 (I608800,I473961);
nand I_35663 (I608817,I608800,I608783);
nor I_35664 (I608672,I608775,I608817);
DFFARX1 I_35665 (I608817,I2507,I608701,I608857,);
not I_35666 (I608693,I608857);
not I_35667 (I608879,I473979);
nand I_35668 (I608896,I608800,I608879);
DFFARX1 I_35669 (I608896,I2507,I608701,I608922,);
not I_35670 (I608930,I608922);
not I_35671 (I608947,I473973);
nand I_35672 (I608964,I608947,I473964);
and I_35673 (I608981,I608783,I608964);
nor I_35674 (I608998,I608896,I608981);
DFFARX1 I_35675 (I608998,I2507,I608701,I608669,);
DFFARX1 I_35676 (I608981,I2507,I608701,I608690,);
nor I_35677 (I609043,I473973,I473982);
nor I_35678 (I608681,I608896,I609043);
or I_35679 (I609074,I473973,I473982);
nor I_35680 (I609091,I473967,I473967);
DFFARX1 I_35681 (I609091,I2507,I608701,I609117,);
not I_35682 (I609125,I609117);
nor I_35683 (I608687,I609125,I608930);
nand I_35684 (I609156,I609125,I608775);
not I_35685 (I609173,I473967);
nand I_35686 (I609190,I609173,I608879);
nand I_35687 (I609207,I609125,I609190);
nand I_35688 (I608678,I609207,I609156);
nand I_35689 (I608675,I609190,I609074);
not I_35690 (I609279,I2514);
DFFARX1 I_35691 (I562109,I2507,I609279,I609305,);
and I_35692 (I609313,I609305,I562106);
DFFARX1 I_35693 (I609313,I2507,I609279,I609262,);
DFFARX1 I_35694 (I562112,I2507,I609279,I609353,);
not I_35695 (I609361,I562115);
not I_35696 (I609378,I562109);
nand I_35697 (I609395,I609378,I609361);
nor I_35698 (I609250,I609353,I609395);
DFFARX1 I_35699 (I609395,I2507,I609279,I609435,);
not I_35700 (I609271,I609435);
not I_35701 (I609457,I562124);
nand I_35702 (I609474,I609378,I609457);
DFFARX1 I_35703 (I609474,I2507,I609279,I609500,);
not I_35704 (I609508,I609500);
not I_35705 (I609525,I562121);
nand I_35706 (I609542,I609525,I562127);
and I_35707 (I609559,I609361,I609542);
nor I_35708 (I609576,I609474,I609559);
DFFARX1 I_35709 (I609576,I2507,I609279,I609247,);
DFFARX1 I_35710 (I609559,I2507,I609279,I609268,);
nor I_35711 (I609621,I562121,I562106);
nor I_35712 (I609259,I609474,I609621);
or I_35713 (I609652,I562121,I562106);
nor I_35714 (I609669,I562118,I562112);
DFFARX1 I_35715 (I609669,I2507,I609279,I609695,);
not I_35716 (I609703,I609695);
nor I_35717 (I609265,I609703,I609508);
nand I_35718 (I609734,I609703,I609353);
not I_35719 (I609751,I562118);
nand I_35720 (I609768,I609751,I609457);
nand I_35721 (I609785,I609703,I609768);
nand I_35722 (I609256,I609785,I609734);
nand I_35723 (I609253,I609768,I609652);
not I_35724 (I609857,I2514);
DFFARX1 I_35725 (I419508,I2507,I609857,I609883,);
and I_35726 (I609891,I609883,I419496);
DFFARX1 I_35727 (I609891,I2507,I609857,I609840,);
DFFARX1 I_35728 (I419499,I2507,I609857,I609931,);
not I_35729 (I609939,I419493);
not I_35730 (I609956,I419517);
nand I_35731 (I609973,I609956,I609939);
nor I_35732 (I609828,I609931,I609973);
DFFARX1 I_35733 (I609973,I2507,I609857,I610013,);
not I_35734 (I609849,I610013);
not I_35735 (I610035,I419505);
nand I_35736 (I610052,I609956,I610035);
DFFARX1 I_35737 (I610052,I2507,I609857,I610078,);
not I_35738 (I610086,I610078);
not I_35739 (I610103,I419514);
nand I_35740 (I610120,I610103,I419511);
and I_35741 (I610137,I609939,I610120);
nor I_35742 (I610154,I610052,I610137);
DFFARX1 I_35743 (I610154,I2507,I609857,I609825,);
DFFARX1 I_35744 (I610137,I2507,I609857,I609846,);
nor I_35745 (I610199,I419514,I419502);
nor I_35746 (I609837,I610052,I610199);
or I_35747 (I610230,I419514,I419502);
nor I_35748 (I610247,I419493,I419496);
DFFARX1 I_35749 (I610247,I2507,I609857,I610273,);
not I_35750 (I610281,I610273);
nor I_35751 (I609843,I610281,I610086);
nand I_35752 (I610312,I610281,I609931);
not I_35753 (I610329,I419493);
nand I_35754 (I610346,I610329,I610035);
nand I_35755 (I610363,I610281,I610346);
nand I_35756 (I609834,I610363,I610312);
nand I_35757 (I609831,I610346,I610230);
not I_35758 (I610435,I2514);
DFFARX1 I_35759 (I18803,I2507,I610435,I610461,);
and I_35760 (I610469,I610461,I18806);
DFFARX1 I_35761 (I610469,I2507,I610435,I610418,);
DFFARX1 I_35762 (I18806,I2507,I610435,I610509,);
not I_35763 (I610517,I18809);
not I_35764 (I610534,I18824);
nand I_35765 (I610551,I610534,I610517);
nor I_35766 (I610406,I610509,I610551);
DFFARX1 I_35767 (I610551,I2507,I610435,I610591,);
not I_35768 (I610427,I610591);
not I_35769 (I610613,I18818);
nand I_35770 (I610630,I610534,I610613);
DFFARX1 I_35771 (I610630,I2507,I610435,I610656,);
not I_35772 (I610664,I610656);
not I_35773 (I610681,I18821);
nand I_35774 (I610698,I610681,I18803);
and I_35775 (I610715,I610517,I610698);
nor I_35776 (I610732,I610630,I610715);
DFFARX1 I_35777 (I610732,I2507,I610435,I610403,);
DFFARX1 I_35778 (I610715,I2507,I610435,I610424,);
nor I_35779 (I610777,I18821,I18815);
nor I_35780 (I610415,I610630,I610777);
or I_35781 (I610808,I18821,I18815);
nor I_35782 (I610825,I18812,I18827);
DFFARX1 I_35783 (I610825,I2507,I610435,I610851,);
not I_35784 (I610859,I610851);
nor I_35785 (I610421,I610859,I610664);
nand I_35786 (I610890,I610859,I610509);
not I_35787 (I610907,I18812);
nand I_35788 (I610924,I610907,I610613);
nand I_35789 (I610941,I610859,I610924);
nand I_35790 (I610412,I610941,I610890);
nand I_35791 (I610409,I610924,I610808);
not I_35792 (I611013,I2514);
DFFARX1 I_35793 (I144909,I2507,I611013,I611039,);
and I_35794 (I611047,I611039,I144912);
DFFARX1 I_35795 (I611047,I2507,I611013,I610996,);
DFFARX1 I_35796 (I144912,I2507,I611013,I611087,);
not I_35797 (I611095,I144927);
not I_35798 (I611112,I144933);
nand I_35799 (I611129,I611112,I611095);
nor I_35800 (I610984,I611087,I611129);
DFFARX1 I_35801 (I611129,I2507,I611013,I611169,);
not I_35802 (I611005,I611169);
not I_35803 (I611191,I144921);
nand I_35804 (I611208,I611112,I611191);
DFFARX1 I_35805 (I611208,I2507,I611013,I611234,);
not I_35806 (I611242,I611234);
not I_35807 (I611259,I144918);
nand I_35808 (I611276,I611259,I144915);
and I_35809 (I611293,I611095,I611276);
nor I_35810 (I611310,I611208,I611293);
DFFARX1 I_35811 (I611310,I2507,I611013,I610981,);
DFFARX1 I_35812 (I611293,I2507,I611013,I611002,);
nor I_35813 (I611355,I144918,I144909);
nor I_35814 (I610993,I611208,I611355);
or I_35815 (I611386,I144918,I144909);
nor I_35816 (I611403,I144924,I144930);
DFFARX1 I_35817 (I611403,I2507,I611013,I611429,);
not I_35818 (I611437,I611429);
nor I_35819 (I610999,I611437,I611242);
nand I_35820 (I611468,I611437,I611087);
not I_35821 (I611485,I144924);
nand I_35822 (I611502,I611485,I611191);
nand I_35823 (I611519,I611437,I611502);
nand I_35824 (I610990,I611519,I611468);
nand I_35825 (I610987,I611502,I611386);
not I_35826 (I611591,I2514);
DFFARX1 I_35827 (I535796,I2507,I611591,I611617,);
and I_35828 (I611625,I611617,I535790);
DFFARX1 I_35829 (I611625,I2507,I611591,I611574,);
DFFARX1 I_35830 (I535808,I2507,I611591,I611665,);
not I_35831 (I611673,I535799);
not I_35832 (I611690,I535811);
nand I_35833 (I611707,I611690,I611673);
nor I_35834 (I611562,I611665,I611707);
DFFARX1 I_35835 (I611707,I2507,I611591,I611747,);
not I_35836 (I611583,I611747);
not I_35837 (I611769,I535817);
nand I_35838 (I611786,I611690,I611769);
DFFARX1 I_35839 (I611786,I2507,I611591,I611812,);
not I_35840 (I611820,I611812);
not I_35841 (I611837,I535793);
nand I_35842 (I611854,I611837,I535814);
and I_35843 (I611871,I611673,I611854);
nor I_35844 (I611888,I611786,I611871);
DFFARX1 I_35845 (I611888,I2507,I611591,I611559,);
DFFARX1 I_35846 (I611871,I2507,I611591,I611580,);
nor I_35847 (I611933,I535793,I535805);
nor I_35848 (I611571,I611786,I611933);
or I_35849 (I611964,I535793,I535805);
nor I_35850 (I611981,I535790,I535802);
DFFARX1 I_35851 (I611981,I2507,I611591,I612007,);
not I_35852 (I612015,I612007);
nor I_35853 (I611577,I612015,I611820);
nand I_35854 (I612046,I612015,I611665);
not I_35855 (I612063,I535790);
nand I_35856 (I612080,I612063,I611769);
nand I_35857 (I612097,I612015,I612080);
nand I_35858 (I611568,I612097,I612046);
nand I_35859 (I611565,I612080,I611964);
not I_35860 (I612169,I2514);
DFFARX1 I_35861 (I45704,I2507,I612169,I612195,);
and I_35862 (I612203,I612195,I45680);
DFFARX1 I_35863 (I612203,I2507,I612169,I612152,);
DFFARX1 I_35864 (I45698,I2507,I612169,I612243,);
not I_35865 (I612251,I45686);
not I_35866 (I612268,I45683);
nand I_35867 (I612285,I612268,I612251);
nor I_35868 (I612140,I612243,I612285);
DFFARX1 I_35869 (I612285,I2507,I612169,I612325,);
not I_35870 (I612161,I612325);
not I_35871 (I612347,I45692);
nand I_35872 (I612364,I612268,I612347);
DFFARX1 I_35873 (I612364,I2507,I612169,I612390,);
not I_35874 (I612398,I612390);
not I_35875 (I612415,I45683);
nand I_35876 (I612432,I612415,I45701);
and I_35877 (I612449,I612251,I612432);
nor I_35878 (I612466,I612364,I612449);
DFFARX1 I_35879 (I612466,I2507,I612169,I612137,);
DFFARX1 I_35880 (I612449,I2507,I612169,I612158,);
nor I_35881 (I612511,I45683,I45695);
nor I_35882 (I612149,I612364,I612511);
or I_35883 (I612542,I45683,I45695);
nor I_35884 (I612559,I45689,I45680);
DFFARX1 I_35885 (I612559,I2507,I612169,I612585,);
not I_35886 (I612593,I612585);
nor I_35887 (I612155,I612593,I612398);
nand I_35888 (I612624,I612593,I612243);
not I_35889 (I612641,I45689);
nand I_35890 (I612658,I612641,I612347);
nand I_35891 (I612675,I612593,I612658);
nand I_35892 (I612146,I612675,I612624);
nand I_35893 (I612143,I612658,I612542);
not I_35894 (I612747,I2514);
DFFARX1 I_35895 (I29870,I2507,I612747,I612773,);
and I_35896 (I612781,I612773,I29873);
DFFARX1 I_35897 (I612781,I2507,I612747,I612730,);
DFFARX1 I_35898 (I29873,I2507,I612747,I612821,);
not I_35899 (I612829,I29876);
not I_35900 (I612846,I29891);
nand I_35901 (I612863,I612846,I612829);
nor I_35902 (I612718,I612821,I612863);
DFFARX1 I_35903 (I612863,I2507,I612747,I612903,);
not I_35904 (I612739,I612903);
not I_35905 (I612925,I29885);
nand I_35906 (I612942,I612846,I612925);
DFFARX1 I_35907 (I612942,I2507,I612747,I612968,);
not I_35908 (I612976,I612968);
not I_35909 (I612993,I29888);
nand I_35910 (I613010,I612993,I29870);
and I_35911 (I613027,I612829,I613010);
nor I_35912 (I613044,I612942,I613027);
DFFARX1 I_35913 (I613044,I2507,I612747,I612715,);
DFFARX1 I_35914 (I613027,I2507,I612747,I612736,);
nor I_35915 (I613089,I29888,I29882);
nor I_35916 (I612727,I612942,I613089);
or I_35917 (I613120,I29888,I29882);
nor I_35918 (I613137,I29879,I29894);
DFFARX1 I_35919 (I613137,I2507,I612747,I613163,);
not I_35920 (I613171,I613163);
nor I_35921 (I612733,I613171,I612976);
nand I_35922 (I613202,I613171,I612821);
not I_35923 (I613219,I29879);
nand I_35924 (I613236,I613219,I612925);
nand I_35925 (I613253,I613171,I613236);
nand I_35926 (I612724,I613253,I613202);
nand I_35927 (I612721,I613236,I613120);
not I_35928 (I613325,I2514);
DFFARX1 I_35929 (I11425,I2507,I613325,I613351,);
and I_35930 (I613359,I613351,I11428);
DFFARX1 I_35931 (I613359,I2507,I613325,I613308,);
DFFARX1 I_35932 (I11428,I2507,I613325,I613399,);
not I_35933 (I613407,I11431);
not I_35934 (I613424,I11446);
nand I_35935 (I613441,I613424,I613407);
nor I_35936 (I613296,I613399,I613441);
DFFARX1 I_35937 (I613441,I2507,I613325,I613481,);
not I_35938 (I613317,I613481);
not I_35939 (I613503,I11440);
nand I_35940 (I613520,I613424,I613503);
DFFARX1 I_35941 (I613520,I2507,I613325,I613546,);
not I_35942 (I613554,I613546);
not I_35943 (I613571,I11443);
nand I_35944 (I613588,I613571,I11425);
and I_35945 (I613605,I613407,I613588);
nor I_35946 (I613622,I613520,I613605);
DFFARX1 I_35947 (I613622,I2507,I613325,I613293,);
DFFARX1 I_35948 (I613605,I2507,I613325,I613314,);
nor I_35949 (I613667,I11443,I11437);
nor I_35950 (I613305,I613520,I613667);
or I_35951 (I613698,I11443,I11437);
nor I_35952 (I613715,I11434,I11449);
DFFARX1 I_35953 (I613715,I2507,I613325,I613741,);
not I_35954 (I613749,I613741);
nor I_35955 (I613311,I613749,I613554);
nand I_35956 (I613780,I613749,I613399);
not I_35957 (I613797,I11434);
nand I_35958 (I613814,I613797,I613503);
nand I_35959 (I613831,I613749,I613814);
nand I_35960 (I613302,I613831,I613780);
nand I_35961 (I613299,I613814,I613698);
not I_35962 (I613903,I2514);
DFFARX1 I_35963 (I295651,I2507,I613903,I613929,);
and I_35964 (I613937,I613929,I295666);
DFFARX1 I_35965 (I613937,I2507,I613903,I613886,);
DFFARX1 I_35966 (I295657,I2507,I613903,I613977,);
not I_35967 (I613985,I295651);
not I_35968 (I614002,I295669);
nand I_35969 (I614019,I614002,I613985);
nor I_35970 (I613874,I613977,I614019);
DFFARX1 I_35971 (I614019,I2507,I613903,I614059,);
not I_35972 (I613895,I614059);
not I_35973 (I614081,I295660);
nand I_35974 (I614098,I614002,I614081);
DFFARX1 I_35975 (I614098,I2507,I613903,I614124,);
not I_35976 (I614132,I614124);
not I_35977 (I614149,I295672);
nand I_35978 (I614166,I614149,I295648);
and I_35979 (I614183,I613985,I614166);
nor I_35980 (I614200,I614098,I614183);
DFFARX1 I_35981 (I614200,I2507,I613903,I613871,);
DFFARX1 I_35982 (I614183,I2507,I613903,I613892,);
nor I_35983 (I614245,I295672,I295648);
nor I_35984 (I613883,I614098,I614245);
or I_35985 (I614276,I295672,I295648);
nor I_35986 (I614293,I295654,I295663);
DFFARX1 I_35987 (I614293,I2507,I613903,I614319,);
not I_35988 (I614327,I614319);
nor I_35989 (I613889,I614327,I614132);
nand I_35990 (I614358,I614327,I613977);
not I_35991 (I614375,I295654);
nand I_35992 (I614392,I614375,I614081);
nand I_35993 (I614409,I614327,I614392);
nand I_35994 (I613880,I614409,I614358);
nand I_35995 (I613877,I614392,I614276);
not I_35996 (I614481,I2514);
DFFARX1 I_35997 (I657786,I2507,I614481,I614507,);
and I_35998 (I614515,I614507,I657780);
DFFARX1 I_35999 (I614515,I2507,I614481,I614464,);
DFFARX1 I_36000 (I657765,I2507,I614481,I614555,);
not I_36001 (I614563,I657771);
not I_36002 (I614580,I657783);
nand I_36003 (I614597,I614580,I614563);
nor I_36004 (I614452,I614555,I614597);
DFFARX1 I_36005 (I614597,I2507,I614481,I614637,);
not I_36006 (I614473,I614637);
not I_36007 (I614659,I657765);
nand I_36008 (I614676,I614580,I614659);
DFFARX1 I_36009 (I614676,I2507,I614481,I614702,);
not I_36010 (I614710,I614702);
not I_36011 (I614727,I657789);
nand I_36012 (I614744,I614727,I657777);
and I_36013 (I614761,I614563,I614744);
nor I_36014 (I614778,I614676,I614761);
DFFARX1 I_36015 (I614778,I2507,I614481,I614449,);
DFFARX1 I_36016 (I614761,I2507,I614481,I614470,);
nor I_36017 (I614823,I657789,I657768);
nor I_36018 (I614461,I614676,I614823);
or I_36019 (I614854,I657789,I657768);
nor I_36020 (I614871,I657774,I657768);
DFFARX1 I_36021 (I614871,I2507,I614481,I614897,);
not I_36022 (I614905,I614897);
nor I_36023 (I614467,I614905,I614710);
nand I_36024 (I614936,I614905,I614555);
not I_36025 (I614953,I657774);
nand I_36026 (I614970,I614953,I614659);
nand I_36027 (I614987,I614905,I614970);
nand I_36028 (I614458,I614987,I614936);
nand I_36029 (I614455,I614970,I614854);
not I_36030 (I615059,I2514);
DFFARX1 I_36031 (I108019,I2507,I615059,I615085,);
and I_36032 (I615093,I615085,I108022);
DFFARX1 I_36033 (I615093,I2507,I615059,I615042,);
DFFARX1 I_36034 (I108022,I2507,I615059,I615133,);
not I_36035 (I615141,I108037);
not I_36036 (I615158,I108043);
nand I_36037 (I615175,I615158,I615141);
nor I_36038 (I615030,I615133,I615175);
DFFARX1 I_36039 (I615175,I2507,I615059,I615215,);
not I_36040 (I615051,I615215);
not I_36041 (I615237,I108031);
nand I_36042 (I615254,I615158,I615237);
DFFARX1 I_36043 (I615254,I2507,I615059,I615280,);
not I_36044 (I615288,I615280);
not I_36045 (I615305,I108028);
nand I_36046 (I615322,I615305,I108025);
and I_36047 (I615339,I615141,I615322);
nor I_36048 (I615356,I615254,I615339);
DFFARX1 I_36049 (I615356,I2507,I615059,I615027,);
DFFARX1 I_36050 (I615339,I2507,I615059,I615048,);
nor I_36051 (I615401,I108028,I108019);
nor I_36052 (I615039,I615254,I615401);
or I_36053 (I615432,I108028,I108019);
nor I_36054 (I615449,I108034,I108040);
DFFARX1 I_36055 (I615449,I2507,I615059,I615475,);
not I_36056 (I615483,I615475);
nor I_36057 (I615045,I615483,I615288);
nand I_36058 (I615514,I615483,I615133);
not I_36059 (I615531,I108034);
nand I_36060 (I615548,I615531,I615237);
nand I_36061 (I615565,I615483,I615548);
nand I_36062 (I615036,I615565,I615514);
nand I_36063 (I615033,I615548,I615432);
not I_36064 (I615637,I2514);
DFFARX1 I_36065 (I381360,I2507,I615637,I615663,);
and I_36066 (I615671,I615663,I381348);
DFFARX1 I_36067 (I615671,I2507,I615637,I615620,);
DFFARX1 I_36068 (I381351,I2507,I615637,I615711,);
not I_36069 (I615719,I381345);
not I_36070 (I615736,I381369);
nand I_36071 (I615753,I615736,I615719);
nor I_36072 (I615608,I615711,I615753);
DFFARX1 I_36073 (I615753,I2507,I615637,I615793,);
not I_36074 (I615629,I615793);
not I_36075 (I615815,I381357);
nand I_36076 (I615832,I615736,I615815);
DFFARX1 I_36077 (I615832,I2507,I615637,I615858,);
not I_36078 (I615866,I615858);
not I_36079 (I615883,I381366);
nand I_36080 (I615900,I615883,I381363);
and I_36081 (I615917,I615719,I615900);
nor I_36082 (I615934,I615832,I615917);
DFFARX1 I_36083 (I615934,I2507,I615637,I615605,);
DFFARX1 I_36084 (I615917,I2507,I615637,I615626,);
nor I_36085 (I615979,I381366,I381354);
nor I_36086 (I615617,I615832,I615979);
or I_36087 (I616010,I381366,I381354);
nor I_36088 (I616027,I381345,I381348);
DFFARX1 I_36089 (I616027,I2507,I615637,I616053,);
not I_36090 (I616061,I616053);
nor I_36091 (I615623,I616061,I615866);
nand I_36092 (I616092,I616061,I615711);
not I_36093 (I616109,I381345);
nand I_36094 (I616126,I616109,I615815);
nand I_36095 (I616143,I616061,I616126);
nand I_36096 (I615614,I616143,I616092);
nand I_36097 (I615611,I616126,I616010);
not I_36098 (I616215,I2514);
DFFARX1 I_36099 (I442344,I2507,I616215,I616241,);
and I_36100 (I616249,I616241,I442350);
DFFARX1 I_36101 (I616249,I2507,I616215,I616198,);
DFFARX1 I_36102 (I442356,I2507,I616215,I616289,);
not I_36103 (I616297,I442341);
not I_36104 (I616314,I442341);
nand I_36105 (I616331,I616314,I616297);
nor I_36106 (I616186,I616289,I616331);
DFFARX1 I_36107 (I616331,I2507,I616215,I616371,);
not I_36108 (I616207,I616371);
not I_36109 (I616393,I442359);
nand I_36110 (I616410,I616314,I616393);
DFFARX1 I_36111 (I616410,I2507,I616215,I616436,);
not I_36112 (I616444,I616436);
not I_36113 (I616461,I442353);
nand I_36114 (I616478,I616461,I442344);
and I_36115 (I616495,I616297,I616478);
nor I_36116 (I616512,I616410,I616495);
DFFARX1 I_36117 (I616512,I2507,I616215,I616183,);
DFFARX1 I_36118 (I616495,I2507,I616215,I616204,);
nor I_36119 (I616557,I442353,I442362);
nor I_36120 (I616195,I616410,I616557);
or I_36121 (I616588,I442353,I442362);
nor I_36122 (I616605,I442347,I442347);
DFFARX1 I_36123 (I616605,I2507,I616215,I616631,);
not I_36124 (I616639,I616631);
nor I_36125 (I616201,I616639,I616444);
nand I_36126 (I616670,I616639,I616289);
not I_36127 (I616687,I442347);
nand I_36128 (I616704,I616687,I616393);
nand I_36129 (I616721,I616639,I616704);
nand I_36130 (I616192,I616721,I616670);
nand I_36131 (I616189,I616704,I616588);
not I_36132 (I616793,I2514);
DFFARX1 I_36133 (I35164,I2507,I616793,I616819,);
and I_36134 (I616827,I616819,I35140);
DFFARX1 I_36135 (I616827,I2507,I616793,I616776,);
DFFARX1 I_36136 (I35158,I2507,I616793,I616867,);
not I_36137 (I616875,I35146);
not I_36138 (I616892,I35143);
nand I_36139 (I616909,I616892,I616875);
nor I_36140 (I616764,I616867,I616909);
DFFARX1 I_36141 (I616909,I2507,I616793,I616949,);
not I_36142 (I616785,I616949);
not I_36143 (I616971,I35152);
nand I_36144 (I616988,I616892,I616971);
DFFARX1 I_36145 (I616988,I2507,I616793,I617014,);
not I_36146 (I617022,I617014);
not I_36147 (I617039,I35143);
nand I_36148 (I617056,I617039,I35161);
and I_36149 (I617073,I616875,I617056);
nor I_36150 (I617090,I616988,I617073);
DFFARX1 I_36151 (I617090,I2507,I616793,I616761,);
DFFARX1 I_36152 (I617073,I2507,I616793,I616782,);
nor I_36153 (I617135,I35143,I35155);
nor I_36154 (I616773,I616988,I617135);
or I_36155 (I617166,I35143,I35155);
nor I_36156 (I617183,I35149,I35140);
DFFARX1 I_36157 (I617183,I2507,I616793,I617209,);
not I_36158 (I617217,I617209);
nor I_36159 (I616779,I617217,I617022);
nand I_36160 (I617248,I617217,I616867);
not I_36161 (I617265,I35149);
nand I_36162 (I617282,I617265,I616971);
nand I_36163 (I617299,I617217,I617282);
nand I_36164 (I616770,I617299,I617248);
nand I_36165 (I616767,I617282,I617166);
not I_36166 (I617371,I2514);
DFFARX1 I_36167 (I184325,I2507,I617371,I617397,);
and I_36168 (I617405,I617397,I184310);
DFFARX1 I_36169 (I617405,I2507,I617371,I617354,);
DFFARX1 I_36170 (I184316,I2507,I617371,I617445,);
not I_36171 (I617453,I184298);
not I_36172 (I617470,I184319);
nand I_36173 (I617487,I617470,I617453);
nor I_36174 (I617342,I617445,I617487);
DFFARX1 I_36175 (I617487,I2507,I617371,I617527,);
not I_36176 (I617363,I617527);
not I_36177 (I617549,I184322);
nand I_36178 (I617566,I617470,I617549);
DFFARX1 I_36179 (I617566,I2507,I617371,I617592,);
not I_36180 (I617600,I617592);
not I_36181 (I617617,I184313);
nand I_36182 (I617634,I617617,I184301);
and I_36183 (I617651,I617453,I617634);
nor I_36184 (I617668,I617566,I617651);
DFFARX1 I_36185 (I617668,I2507,I617371,I617339,);
DFFARX1 I_36186 (I617651,I2507,I617371,I617360,);
nor I_36187 (I617713,I184313,I184307);
nor I_36188 (I617351,I617566,I617713);
or I_36189 (I617744,I184313,I184307);
nor I_36190 (I617761,I184304,I184298);
DFFARX1 I_36191 (I617761,I2507,I617371,I617787,);
not I_36192 (I617795,I617787);
nor I_36193 (I617357,I617795,I617600);
nand I_36194 (I617826,I617795,I617445);
not I_36195 (I617843,I184304);
nand I_36196 (I617860,I617843,I617549);
nand I_36197 (I617877,I617795,I617860);
nand I_36198 (I617348,I617877,I617826);
nand I_36199 (I617345,I617860,I617744);
not I_36200 (I617949,I2514);
DFFARX1 I_36201 (I326450,I2507,I617949,I617975,);
and I_36202 (I617983,I617975,I326438);
DFFARX1 I_36203 (I617983,I2507,I617949,I617932,);
DFFARX1 I_36204 (I326453,I2507,I617949,I618023,);
not I_36205 (I618031,I326444);
not I_36206 (I618048,I326435);
nand I_36207 (I618065,I618048,I618031);
nor I_36208 (I617920,I618023,I618065);
DFFARX1 I_36209 (I618065,I2507,I617949,I618105,);
not I_36210 (I617941,I618105);
not I_36211 (I618127,I326441);
nand I_36212 (I618144,I618048,I618127);
DFFARX1 I_36213 (I618144,I2507,I617949,I618170,);
not I_36214 (I618178,I618170);
not I_36215 (I618195,I326456);
nand I_36216 (I618212,I618195,I326459);
and I_36217 (I618229,I618031,I618212);
nor I_36218 (I618246,I618144,I618229);
DFFARX1 I_36219 (I618246,I2507,I617949,I617917,);
DFFARX1 I_36220 (I618229,I2507,I617949,I617938,);
nor I_36221 (I618291,I326456,I326435);
nor I_36222 (I617929,I618144,I618291);
or I_36223 (I618322,I326456,I326435);
nor I_36224 (I618339,I326447,I326438);
DFFARX1 I_36225 (I618339,I2507,I617949,I618365,);
not I_36226 (I618373,I618365);
nor I_36227 (I617935,I618373,I618178);
nand I_36228 (I618404,I618373,I618023);
not I_36229 (I618421,I326447);
nand I_36230 (I618438,I618421,I618127);
nand I_36231 (I618455,I618373,I618438);
nand I_36232 (I617926,I618455,I618404);
nand I_36233 (I617923,I618438,I618322);
not I_36234 (I618527,I2514);
DFFARX1 I_36235 (I644186,I2507,I618527,I618553,);
and I_36236 (I618561,I618553,I644180);
DFFARX1 I_36237 (I618561,I2507,I618527,I618510,);
DFFARX1 I_36238 (I644165,I2507,I618527,I618601,);
not I_36239 (I618609,I644171);
not I_36240 (I618626,I644183);
nand I_36241 (I618643,I618626,I618609);
nor I_36242 (I618498,I618601,I618643);
DFFARX1 I_36243 (I618643,I2507,I618527,I618683,);
not I_36244 (I618519,I618683);
not I_36245 (I618705,I644165);
nand I_36246 (I618722,I618626,I618705);
DFFARX1 I_36247 (I618722,I2507,I618527,I618748,);
not I_36248 (I618756,I618748);
not I_36249 (I618773,I644189);
nand I_36250 (I618790,I618773,I644177);
and I_36251 (I618807,I618609,I618790);
nor I_36252 (I618824,I618722,I618807);
DFFARX1 I_36253 (I618824,I2507,I618527,I618495,);
DFFARX1 I_36254 (I618807,I2507,I618527,I618516,);
nor I_36255 (I618869,I644189,I644168);
nor I_36256 (I618507,I618722,I618869);
or I_36257 (I618900,I644189,I644168);
nor I_36258 (I618917,I644174,I644168);
DFFARX1 I_36259 (I618917,I2507,I618527,I618943,);
not I_36260 (I618951,I618943);
nor I_36261 (I618513,I618951,I618756);
nand I_36262 (I618982,I618951,I618601);
not I_36263 (I618999,I644174);
nand I_36264 (I619016,I618999,I618705);
nand I_36265 (I619033,I618951,I619016);
nand I_36266 (I618504,I619033,I618982);
nand I_36267 (I618501,I619016,I618900);
not I_36268 (I619105,I2514);
DFFARX1 I_36269 (I26708,I2507,I619105,I619131,);
and I_36270 (I619139,I619131,I26711);
DFFARX1 I_36271 (I619139,I2507,I619105,I619088,);
DFFARX1 I_36272 (I26711,I2507,I619105,I619179,);
not I_36273 (I619187,I26714);
not I_36274 (I619204,I26729);
nand I_36275 (I619221,I619204,I619187);
nor I_36276 (I619076,I619179,I619221);
DFFARX1 I_36277 (I619221,I2507,I619105,I619261,);
not I_36278 (I619097,I619261);
not I_36279 (I619283,I26723);
nand I_36280 (I619300,I619204,I619283);
DFFARX1 I_36281 (I619300,I2507,I619105,I619326,);
not I_36282 (I619334,I619326);
not I_36283 (I619351,I26726);
nand I_36284 (I619368,I619351,I26708);
and I_36285 (I619385,I619187,I619368);
nor I_36286 (I619402,I619300,I619385);
DFFARX1 I_36287 (I619402,I2507,I619105,I619073,);
DFFARX1 I_36288 (I619385,I2507,I619105,I619094,);
nor I_36289 (I619447,I26726,I26720);
nor I_36290 (I619085,I619300,I619447);
or I_36291 (I619478,I26726,I26720);
nor I_36292 (I619495,I26717,I26732);
DFFARX1 I_36293 (I619495,I2507,I619105,I619521,);
not I_36294 (I619529,I619521);
nor I_36295 (I619091,I619529,I619334);
nand I_36296 (I619560,I619529,I619179);
not I_36297 (I619577,I26717);
nand I_36298 (I619594,I619577,I619283);
nand I_36299 (I619611,I619529,I619594);
nand I_36300 (I619082,I619611,I619560);
nand I_36301 (I619079,I619594,I619478);
not I_36302 (I619683,I2514);
DFFARX1 I_36303 (I513832,I2507,I619683,I619709,);
and I_36304 (I619717,I619709,I513826);
DFFARX1 I_36305 (I619717,I2507,I619683,I619666,);
DFFARX1 I_36306 (I513844,I2507,I619683,I619757,);
not I_36307 (I619765,I513835);
not I_36308 (I619782,I513847);
nand I_36309 (I619799,I619782,I619765);
nor I_36310 (I619654,I619757,I619799);
DFFARX1 I_36311 (I619799,I2507,I619683,I619839,);
not I_36312 (I619675,I619839);
not I_36313 (I619861,I513853);
nand I_36314 (I619878,I619782,I619861);
DFFARX1 I_36315 (I619878,I2507,I619683,I619904,);
not I_36316 (I619912,I619904);
not I_36317 (I619929,I513829);
nand I_36318 (I619946,I619929,I513850);
and I_36319 (I619963,I619765,I619946);
nor I_36320 (I619980,I619878,I619963);
DFFARX1 I_36321 (I619980,I2507,I619683,I619651,);
DFFARX1 I_36322 (I619963,I2507,I619683,I619672,);
nor I_36323 (I620025,I513829,I513841);
nor I_36324 (I619663,I619878,I620025);
or I_36325 (I620056,I513829,I513841);
nor I_36326 (I620073,I513826,I513838);
DFFARX1 I_36327 (I620073,I2507,I619683,I620099,);
not I_36328 (I620107,I620099);
nor I_36329 (I619669,I620107,I619912);
nand I_36330 (I620138,I620107,I619757);
not I_36331 (I620155,I513826);
nand I_36332 (I620172,I620155,I619861);
nand I_36333 (I620189,I620107,I620172);
nand I_36334 (I619660,I620189,I620138);
nand I_36335 (I619657,I620172,I620056);
not I_36336 (I620261,I2514);
DFFARX1 I_36337 (I461316,I2507,I620261,I620287,);
and I_36338 (I620295,I620287,I461322);
DFFARX1 I_36339 (I620295,I2507,I620261,I620244,);
DFFARX1 I_36340 (I461328,I2507,I620261,I620335,);
not I_36341 (I620343,I461313);
not I_36342 (I620360,I461313);
nand I_36343 (I620377,I620360,I620343);
nor I_36344 (I620232,I620335,I620377);
DFFARX1 I_36345 (I620377,I2507,I620261,I620417,);
not I_36346 (I620253,I620417);
not I_36347 (I620439,I461331);
nand I_36348 (I620456,I620360,I620439);
DFFARX1 I_36349 (I620456,I2507,I620261,I620482,);
not I_36350 (I620490,I620482);
not I_36351 (I620507,I461325);
nand I_36352 (I620524,I620507,I461316);
and I_36353 (I620541,I620343,I620524);
nor I_36354 (I620558,I620456,I620541);
DFFARX1 I_36355 (I620558,I2507,I620261,I620229,);
DFFARX1 I_36356 (I620541,I2507,I620261,I620250,);
nor I_36357 (I620603,I461325,I461334);
nor I_36358 (I620241,I620456,I620603);
or I_36359 (I620634,I461325,I461334);
nor I_36360 (I620651,I461319,I461319);
DFFARX1 I_36361 (I620651,I2507,I620261,I620677,);
not I_36362 (I620685,I620677);
nor I_36363 (I620247,I620685,I620490);
nand I_36364 (I620716,I620685,I620335);
not I_36365 (I620733,I461319);
nand I_36366 (I620750,I620733,I620439);
nand I_36367 (I620767,I620685,I620750);
nand I_36368 (I620238,I620767,I620716);
nand I_36369 (I620235,I620750,I620634);
not I_36370 (I620839,I2514);
DFFARX1 I_36371 (I322404,I2507,I620839,I620865,);
and I_36372 (I620873,I620865,I322392);
DFFARX1 I_36373 (I620873,I2507,I620839,I620822,);
DFFARX1 I_36374 (I322407,I2507,I620839,I620913,);
not I_36375 (I620921,I322398);
not I_36376 (I620938,I322389);
nand I_36377 (I620955,I620938,I620921);
nor I_36378 (I620810,I620913,I620955);
DFFARX1 I_36379 (I620955,I2507,I620839,I620995,);
not I_36380 (I620831,I620995);
not I_36381 (I621017,I322395);
nand I_36382 (I621034,I620938,I621017);
DFFARX1 I_36383 (I621034,I2507,I620839,I621060,);
not I_36384 (I621068,I621060);
not I_36385 (I621085,I322410);
nand I_36386 (I621102,I621085,I322413);
and I_36387 (I621119,I620921,I621102);
nor I_36388 (I621136,I621034,I621119);
DFFARX1 I_36389 (I621136,I2507,I620839,I620807,);
DFFARX1 I_36390 (I621119,I2507,I620839,I620828,);
nor I_36391 (I621181,I322410,I322389);
nor I_36392 (I620819,I621034,I621181);
or I_36393 (I621212,I322410,I322389);
nor I_36394 (I621229,I322401,I322392);
DFFARX1 I_36395 (I621229,I2507,I620839,I621255,);
not I_36396 (I621263,I621255);
nor I_36397 (I620825,I621263,I621068);
nand I_36398 (I621294,I621263,I620913);
not I_36399 (I621311,I322401);
nand I_36400 (I621328,I621311,I621017);
nand I_36401 (I621345,I621263,I621328);
nand I_36402 (I620816,I621345,I621294);
nand I_36403 (I620813,I621328,I621212);
not I_36404 (I621417,I2514);
DFFARX1 I_36405 (I701975,I2507,I621417,I621443,);
and I_36406 (I621451,I621443,I701957);
DFFARX1 I_36407 (I621451,I2507,I621417,I621400,);
DFFARX1 I_36408 (I701948,I2507,I621417,I621491,);
not I_36409 (I621499,I701963);
not I_36410 (I621516,I701951);
nand I_36411 (I621533,I621516,I621499);
nor I_36412 (I621388,I621491,I621533);
DFFARX1 I_36413 (I621533,I2507,I621417,I621573,);
not I_36414 (I621409,I621573);
not I_36415 (I621595,I701960);
nand I_36416 (I621612,I621516,I621595);
DFFARX1 I_36417 (I621612,I2507,I621417,I621638,);
not I_36418 (I621646,I621638);
not I_36419 (I621663,I701969);
nand I_36420 (I621680,I621663,I701948);
and I_36421 (I621697,I621499,I621680);
nor I_36422 (I621714,I621612,I621697);
DFFARX1 I_36423 (I621714,I2507,I621417,I621385,);
DFFARX1 I_36424 (I621697,I2507,I621417,I621406,);
nor I_36425 (I621759,I701969,I701972);
nor I_36426 (I621397,I621612,I621759);
or I_36427 (I621790,I701969,I701972);
nor I_36428 (I621807,I701966,I701954);
DFFARX1 I_36429 (I621807,I2507,I621417,I621833,);
not I_36430 (I621841,I621833);
nor I_36431 (I621403,I621841,I621646);
nand I_36432 (I621872,I621841,I621491);
not I_36433 (I621889,I701966);
nand I_36434 (I621906,I621889,I621595);
nand I_36435 (I621923,I621841,I621906);
nand I_36436 (I621394,I621923,I621872);
nand I_36437 (I621391,I621906,I621790);
not I_36438 (I621995,I2514);
DFFARX1 I_36439 (I21438,I2507,I621995,I622021,);
and I_36440 (I622029,I622021,I21441);
DFFARX1 I_36441 (I622029,I2507,I621995,I621978,);
DFFARX1 I_36442 (I21441,I2507,I621995,I622069,);
not I_36443 (I622077,I21444);
not I_36444 (I622094,I21459);
nand I_36445 (I622111,I622094,I622077);
nor I_36446 (I621966,I622069,I622111);
DFFARX1 I_36447 (I622111,I2507,I621995,I622151,);
not I_36448 (I621987,I622151);
not I_36449 (I622173,I21453);
nand I_36450 (I622190,I622094,I622173);
DFFARX1 I_36451 (I622190,I2507,I621995,I622216,);
not I_36452 (I622224,I622216);
not I_36453 (I622241,I21456);
nand I_36454 (I622258,I622241,I21438);
and I_36455 (I622275,I622077,I622258);
nor I_36456 (I622292,I622190,I622275);
DFFARX1 I_36457 (I622292,I2507,I621995,I621963,);
DFFARX1 I_36458 (I622275,I2507,I621995,I621984,);
nor I_36459 (I622337,I21456,I21450);
nor I_36460 (I621975,I622190,I622337);
or I_36461 (I622368,I21456,I21450);
nor I_36462 (I622385,I21447,I21462);
DFFARX1 I_36463 (I622385,I2507,I621995,I622411,);
not I_36464 (I622419,I622411);
nor I_36465 (I621981,I622419,I622224);
nand I_36466 (I622450,I622419,I622069);
not I_36467 (I622467,I21447);
nand I_36468 (I622484,I622467,I622173);
nand I_36469 (I622501,I622419,I622484);
nand I_36470 (I621972,I622501,I622450);
nand I_36471 (I621969,I622484,I622368);
not I_36472 (I622573,I2514);
DFFARX1 I_36473 (I4912,I2507,I622573,I622599,);
and I_36474 (I622607,I622599,I4918);
DFFARX1 I_36475 (I622607,I2507,I622573,I622556,);
DFFARX1 I_36476 (I4897,I2507,I622573,I622647,);
not I_36477 (I622655,I4903);
not I_36478 (I622672,I4909);
nand I_36479 (I622689,I622672,I622655);
nor I_36480 (I622544,I622647,I622689);
DFFARX1 I_36481 (I622689,I2507,I622573,I622729,);
not I_36482 (I622565,I622729);
not I_36483 (I622751,I4900);
nand I_36484 (I622768,I622672,I622751);
DFFARX1 I_36485 (I622768,I2507,I622573,I622794,);
not I_36486 (I622802,I622794);
not I_36487 (I622819,I4915);
nand I_36488 (I622836,I622819,I4900);
and I_36489 (I622853,I622655,I622836);
nor I_36490 (I622870,I622768,I622853);
DFFARX1 I_36491 (I622870,I2507,I622573,I622541,);
DFFARX1 I_36492 (I622853,I2507,I622573,I622562,);
nor I_36493 (I622915,I4915,I4903);
nor I_36494 (I622553,I622768,I622915);
or I_36495 (I622946,I4915,I4903);
nor I_36496 (I622963,I4906,I4897);
DFFARX1 I_36497 (I622963,I2507,I622573,I622989,);
not I_36498 (I622997,I622989);
nor I_36499 (I622559,I622997,I622802);
nand I_36500 (I623028,I622997,I622647);
not I_36501 (I623045,I4906);
nand I_36502 (I623062,I623045,I622751);
nand I_36503 (I623079,I622997,I623062);
nand I_36504 (I622550,I623079,I623028);
nand I_36505 (I622547,I623062,I622946);
not I_36506 (I623151,I2514);
DFFARX1 I_36507 (I563231,I2507,I623151,I623177,);
and I_36508 (I623185,I623177,I563228);
DFFARX1 I_36509 (I623185,I2507,I623151,I623134,);
DFFARX1 I_36510 (I563234,I2507,I623151,I623225,);
not I_36511 (I623233,I563237);
not I_36512 (I623250,I563231);
nand I_36513 (I623267,I623250,I623233);
nor I_36514 (I623122,I623225,I623267);
DFFARX1 I_36515 (I623267,I2507,I623151,I623307,);
not I_36516 (I623143,I623307);
not I_36517 (I623329,I563246);
nand I_36518 (I623346,I623250,I623329);
DFFARX1 I_36519 (I623346,I2507,I623151,I623372,);
not I_36520 (I623380,I623372);
not I_36521 (I623397,I563243);
nand I_36522 (I623414,I623397,I563249);
and I_36523 (I623431,I623233,I623414);
nor I_36524 (I623448,I623346,I623431);
DFFARX1 I_36525 (I623448,I2507,I623151,I623119,);
DFFARX1 I_36526 (I623431,I2507,I623151,I623140,);
nor I_36527 (I623493,I563243,I563228);
nor I_36528 (I623131,I623346,I623493);
or I_36529 (I623524,I563243,I563228);
nor I_36530 (I623541,I563240,I563234);
DFFARX1 I_36531 (I623541,I2507,I623151,I623567,);
not I_36532 (I623575,I623567);
nor I_36533 (I623137,I623575,I623380);
nand I_36534 (I623606,I623575,I623225);
not I_36535 (I623623,I563240);
nand I_36536 (I623640,I623623,I623329);
nand I_36537 (I623657,I623575,I623640);
nand I_36538 (I623128,I623657,I623606);
nand I_36539 (I623125,I623640,I623524);
not I_36540 (I623729,I2514);
DFFARX1 I_36541 (I728155,I2507,I623729,I623755,);
and I_36542 (I623763,I623755,I728137);
DFFARX1 I_36543 (I623763,I2507,I623729,I623712,);
DFFARX1 I_36544 (I728128,I2507,I623729,I623803,);
not I_36545 (I623811,I728143);
not I_36546 (I623828,I728131);
nand I_36547 (I623845,I623828,I623811);
nor I_36548 (I623700,I623803,I623845);
DFFARX1 I_36549 (I623845,I2507,I623729,I623885,);
not I_36550 (I623721,I623885);
not I_36551 (I623907,I728140);
nand I_36552 (I623924,I623828,I623907);
DFFARX1 I_36553 (I623924,I2507,I623729,I623950,);
not I_36554 (I623958,I623950);
not I_36555 (I623975,I728149);
nand I_36556 (I623992,I623975,I728128);
and I_36557 (I624009,I623811,I623992);
nor I_36558 (I624026,I623924,I624009);
DFFARX1 I_36559 (I624026,I2507,I623729,I623697,);
DFFARX1 I_36560 (I624009,I2507,I623729,I623718,);
nor I_36561 (I624071,I728149,I728152);
nor I_36562 (I623709,I623924,I624071);
or I_36563 (I624102,I728149,I728152);
nor I_36564 (I624119,I728146,I728134);
DFFARX1 I_36565 (I624119,I2507,I623729,I624145,);
not I_36566 (I624153,I624145);
nor I_36567 (I623715,I624153,I623958);
nand I_36568 (I624184,I624153,I623803);
not I_36569 (I624201,I728146);
nand I_36570 (I624218,I624201,I623907);
nand I_36571 (I624235,I624153,I624218);
nand I_36572 (I623706,I624235,I624184);
nand I_36573 (I623703,I624218,I624102);
not I_36574 (I624307,I2514);
DFFARX1 I_36575 (I475545,I2507,I624307,I624333,);
and I_36576 (I624341,I624333,I475551);
DFFARX1 I_36577 (I624341,I2507,I624307,I624290,);
DFFARX1 I_36578 (I475557,I2507,I624307,I624381,);
not I_36579 (I624389,I475542);
not I_36580 (I624406,I475542);
nand I_36581 (I624423,I624406,I624389);
nor I_36582 (I624278,I624381,I624423);
DFFARX1 I_36583 (I624423,I2507,I624307,I624463,);
not I_36584 (I624299,I624463);
not I_36585 (I624485,I475560);
nand I_36586 (I624502,I624406,I624485);
DFFARX1 I_36587 (I624502,I2507,I624307,I624528,);
not I_36588 (I624536,I624528);
not I_36589 (I624553,I475554);
nand I_36590 (I624570,I624553,I475545);
and I_36591 (I624587,I624389,I624570);
nor I_36592 (I624604,I624502,I624587);
DFFARX1 I_36593 (I624604,I2507,I624307,I624275,);
DFFARX1 I_36594 (I624587,I2507,I624307,I624296,);
nor I_36595 (I624649,I475554,I475563);
nor I_36596 (I624287,I624502,I624649);
or I_36597 (I624680,I475554,I475563);
nor I_36598 (I624697,I475548,I475548);
DFFARX1 I_36599 (I624697,I2507,I624307,I624723,);
not I_36600 (I624731,I624723);
nor I_36601 (I624293,I624731,I624536);
nand I_36602 (I624762,I624731,I624381);
not I_36603 (I624779,I475548);
nand I_36604 (I624796,I624779,I624485);
nand I_36605 (I624813,I624731,I624796);
nand I_36606 (I624284,I624813,I624762);
nand I_36607 (I624281,I624796,I624680);
not I_36608 (I624885,I2514);
DFFARX1 I_36609 (I274840,I2507,I624885,I624911,);
and I_36610 (I624919,I624911,I274855);
DFFARX1 I_36611 (I624919,I2507,I624885,I624868,);
DFFARX1 I_36612 (I274858,I2507,I624885,I624959,);
not I_36613 (I624967,I274852);
not I_36614 (I624984,I274867);
nand I_36615 (I625001,I624984,I624967);
nor I_36616 (I624856,I624959,I625001);
DFFARX1 I_36617 (I625001,I2507,I624885,I625041,);
not I_36618 (I624877,I625041);
not I_36619 (I625063,I274843);
nand I_36620 (I625080,I624984,I625063);
DFFARX1 I_36621 (I625080,I2507,I624885,I625106,);
not I_36622 (I625114,I625106);
not I_36623 (I625131,I274846);
nand I_36624 (I625148,I625131,I274840);
and I_36625 (I625165,I624967,I625148);
nor I_36626 (I625182,I625080,I625165);
DFFARX1 I_36627 (I625182,I2507,I624885,I624853,);
DFFARX1 I_36628 (I625165,I2507,I624885,I624874,);
nor I_36629 (I625227,I274846,I274849);
nor I_36630 (I624865,I625080,I625227);
or I_36631 (I625258,I274846,I274849);
nor I_36632 (I625275,I274864,I274861);
DFFARX1 I_36633 (I625275,I2507,I624885,I625301,);
not I_36634 (I625309,I625301);
nor I_36635 (I624871,I625309,I625114);
nand I_36636 (I625340,I625309,I624959);
not I_36637 (I625357,I274864);
nand I_36638 (I625374,I625357,I625063);
nand I_36639 (I625391,I625309,I625374);
nand I_36640 (I624862,I625391,I625340);
nand I_36641 (I624859,I625374,I625258);
not I_36642 (I625463,I2514);
DFFARX1 I_36643 (I303330,I2507,I625463,I625489,);
and I_36644 (I625497,I625489,I303318);
DFFARX1 I_36645 (I625497,I2507,I625463,I625446,);
DFFARX1 I_36646 (I303333,I2507,I625463,I625537,);
not I_36647 (I625545,I303324);
not I_36648 (I625562,I303315);
nand I_36649 (I625579,I625562,I625545);
nor I_36650 (I625434,I625537,I625579);
DFFARX1 I_36651 (I625579,I2507,I625463,I625619,);
not I_36652 (I625455,I625619);
not I_36653 (I625641,I303321);
nand I_36654 (I625658,I625562,I625641);
DFFARX1 I_36655 (I625658,I2507,I625463,I625684,);
not I_36656 (I625692,I625684);
not I_36657 (I625709,I303336);
nand I_36658 (I625726,I625709,I303339);
and I_36659 (I625743,I625545,I625726);
nor I_36660 (I625760,I625658,I625743);
DFFARX1 I_36661 (I625760,I2507,I625463,I625431,);
DFFARX1 I_36662 (I625743,I2507,I625463,I625452,);
nor I_36663 (I625805,I303336,I303315);
nor I_36664 (I625443,I625658,I625805);
or I_36665 (I625836,I303336,I303315);
nor I_36666 (I625853,I303327,I303318);
DFFARX1 I_36667 (I625853,I2507,I625463,I625879,);
not I_36668 (I625887,I625879);
nor I_36669 (I625449,I625887,I625692);
nand I_36670 (I625918,I625887,I625537);
not I_36671 (I625935,I303327);
nand I_36672 (I625952,I625935,I625641);
nand I_36673 (I625969,I625887,I625952);
nand I_36674 (I625440,I625969,I625918);
nand I_36675 (I625437,I625952,I625836);
not I_36676 (I626041,I2514);
DFFARX1 I_36677 (I75743,I2507,I626041,I626067,);
and I_36678 (I626075,I626067,I75719);
DFFARX1 I_36679 (I626075,I2507,I626041,I626024,);
DFFARX1 I_36680 (I75737,I2507,I626041,I626115,);
not I_36681 (I626123,I75725);
not I_36682 (I626140,I75722);
nand I_36683 (I626157,I626140,I626123);
nor I_36684 (I626012,I626115,I626157);
DFFARX1 I_36685 (I626157,I2507,I626041,I626197,);
not I_36686 (I626033,I626197);
not I_36687 (I626219,I75731);
nand I_36688 (I626236,I626140,I626219);
DFFARX1 I_36689 (I626236,I2507,I626041,I626262,);
not I_36690 (I626270,I626262);
not I_36691 (I626287,I75722);
nand I_36692 (I626304,I626287,I75740);
and I_36693 (I626321,I626123,I626304);
nor I_36694 (I626338,I626236,I626321);
DFFARX1 I_36695 (I626338,I2507,I626041,I626009,);
DFFARX1 I_36696 (I626321,I2507,I626041,I626030,);
nor I_36697 (I626383,I75722,I75734);
nor I_36698 (I626021,I626236,I626383);
or I_36699 (I626414,I75722,I75734);
nor I_36700 (I626431,I75728,I75719);
DFFARX1 I_36701 (I626431,I2507,I626041,I626457,);
not I_36702 (I626465,I626457);
nor I_36703 (I626027,I626465,I626270);
nand I_36704 (I626496,I626465,I626115);
not I_36705 (I626513,I75728);
nand I_36706 (I626530,I626513,I626219);
nand I_36707 (I626547,I626465,I626530);
nand I_36708 (I626018,I626547,I626496);
nand I_36709 (I626015,I626530,I626414);
not I_36710 (I626619,I2514);
DFFARX1 I_36711 (I40961,I2507,I626619,I626645,);
and I_36712 (I626653,I626645,I40937);
DFFARX1 I_36713 (I626653,I2507,I626619,I626602,);
DFFARX1 I_36714 (I40955,I2507,I626619,I626693,);
not I_36715 (I626701,I40943);
not I_36716 (I626718,I40940);
nand I_36717 (I626735,I626718,I626701);
nor I_36718 (I626590,I626693,I626735);
DFFARX1 I_36719 (I626735,I2507,I626619,I626775,);
not I_36720 (I626611,I626775);
not I_36721 (I626797,I40949);
nand I_36722 (I626814,I626718,I626797);
DFFARX1 I_36723 (I626814,I2507,I626619,I626840,);
not I_36724 (I626848,I626840);
not I_36725 (I626865,I40940);
nand I_36726 (I626882,I626865,I40958);
and I_36727 (I626899,I626701,I626882);
nor I_36728 (I626916,I626814,I626899);
DFFARX1 I_36729 (I626916,I2507,I626619,I626587,);
DFFARX1 I_36730 (I626899,I2507,I626619,I626608,);
nor I_36731 (I626961,I40940,I40952);
nor I_36732 (I626599,I626814,I626961);
or I_36733 (I626992,I40940,I40952);
nor I_36734 (I627009,I40946,I40937);
DFFARX1 I_36735 (I627009,I2507,I626619,I627035,);
not I_36736 (I627043,I627035);
nor I_36737 (I626605,I627043,I626848);
nand I_36738 (I627074,I627043,I626693);
not I_36739 (I627091,I40946);
nand I_36740 (I627108,I627091,I626797);
nand I_36741 (I627125,I627043,I627108);
nand I_36742 (I626596,I627125,I627074);
nand I_36743 (I626593,I627108,I626992);
not I_36744 (I627197,I2514);
DFFARX1 I_36745 (I453411,I2507,I627197,I627223,);
and I_36746 (I627231,I627223,I453417);
DFFARX1 I_36747 (I627231,I2507,I627197,I627180,);
DFFARX1 I_36748 (I453423,I2507,I627197,I627271,);
not I_36749 (I627279,I453408);
not I_36750 (I627296,I453408);
nand I_36751 (I627313,I627296,I627279);
nor I_36752 (I627168,I627271,I627313);
DFFARX1 I_36753 (I627313,I2507,I627197,I627353,);
not I_36754 (I627189,I627353);
not I_36755 (I627375,I453426);
nand I_36756 (I627392,I627296,I627375);
DFFARX1 I_36757 (I627392,I2507,I627197,I627418,);
not I_36758 (I627426,I627418);
not I_36759 (I627443,I453420);
nand I_36760 (I627460,I627443,I453411);
and I_36761 (I627477,I627279,I627460);
nor I_36762 (I627494,I627392,I627477);
DFFARX1 I_36763 (I627494,I2507,I627197,I627165,);
DFFARX1 I_36764 (I627477,I2507,I627197,I627186,);
nor I_36765 (I627539,I453420,I453429);
nor I_36766 (I627177,I627392,I627539);
or I_36767 (I627570,I453420,I453429);
nor I_36768 (I627587,I453414,I453414);
DFFARX1 I_36769 (I627587,I2507,I627197,I627613,);
not I_36770 (I627621,I627613);
nor I_36771 (I627183,I627621,I627426);
nand I_36772 (I627652,I627621,I627271);
not I_36773 (I627669,I453414);
nand I_36774 (I627686,I627669,I627375);
nand I_36775 (I627703,I627621,I627686);
nand I_36776 (I627174,I627703,I627652);
nand I_36777 (I627171,I627686,I627570);
not I_36778 (I627775,I2514);
DFFARX1 I_36779 (I91359,I2507,I627775,I627801,);
and I_36780 (I627809,I627801,I91362);
DFFARX1 I_36781 (I627809,I2507,I627775,I627758,);
DFFARX1 I_36782 (I91362,I2507,I627775,I627849,);
not I_36783 (I627857,I91377);
not I_36784 (I627874,I91383);
nand I_36785 (I627891,I627874,I627857);
nor I_36786 (I627746,I627849,I627891);
DFFARX1 I_36787 (I627891,I2507,I627775,I627931,);
not I_36788 (I627767,I627931);
not I_36789 (I627953,I91371);
nand I_36790 (I627970,I627874,I627953);
DFFARX1 I_36791 (I627970,I2507,I627775,I627996,);
not I_36792 (I628004,I627996);
not I_36793 (I628021,I91368);
nand I_36794 (I628038,I628021,I91365);
and I_36795 (I628055,I627857,I628038);
nor I_36796 (I628072,I627970,I628055);
DFFARX1 I_36797 (I628072,I2507,I627775,I627743,);
DFFARX1 I_36798 (I628055,I2507,I627775,I627764,);
nor I_36799 (I628117,I91368,I91359);
nor I_36800 (I627755,I627970,I628117);
or I_36801 (I628148,I91368,I91359);
nor I_36802 (I628165,I91374,I91380);
DFFARX1 I_36803 (I628165,I2507,I627775,I628191,);
not I_36804 (I628199,I628191);
nor I_36805 (I627761,I628199,I628004);
nand I_36806 (I628230,I628199,I627849);
not I_36807 (I628247,I91374);
nand I_36808 (I628264,I628247,I627953);
nand I_36809 (I628281,I628199,I628264);
nand I_36810 (I627752,I628281,I628230);
nand I_36811 (I627749,I628264,I628148);
not I_36812 (I628353,I2514);
DFFARX1 I_36813 (I66257,I2507,I628353,I628379,);
and I_36814 (I628387,I628379,I66233);
DFFARX1 I_36815 (I628387,I2507,I628353,I628336,);
DFFARX1 I_36816 (I66251,I2507,I628353,I628427,);
not I_36817 (I628435,I66239);
not I_36818 (I628452,I66236);
nand I_36819 (I628469,I628452,I628435);
nor I_36820 (I628324,I628427,I628469);
DFFARX1 I_36821 (I628469,I2507,I628353,I628509,);
not I_36822 (I628345,I628509);
not I_36823 (I628531,I66245);
nand I_36824 (I628548,I628452,I628531);
DFFARX1 I_36825 (I628548,I2507,I628353,I628574,);
not I_36826 (I628582,I628574);
not I_36827 (I628599,I66236);
nand I_36828 (I628616,I628599,I66254);
and I_36829 (I628633,I628435,I628616);
nor I_36830 (I628650,I628548,I628633);
DFFARX1 I_36831 (I628650,I2507,I628353,I628321,);
DFFARX1 I_36832 (I628633,I2507,I628353,I628342,);
nor I_36833 (I628695,I66236,I66248);
nor I_36834 (I628333,I628548,I628695);
or I_36835 (I628726,I66236,I66248);
nor I_36836 (I628743,I66242,I66233);
DFFARX1 I_36837 (I628743,I2507,I628353,I628769,);
not I_36838 (I628777,I628769);
nor I_36839 (I628339,I628777,I628582);
nand I_36840 (I628808,I628777,I628427);
not I_36841 (I628825,I66242);
nand I_36842 (I628842,I628825,I628531);
nand I_36843 (I628859,I628777,I628842);
nand I_36844 (I628330,I628859,I628808);
nand I_36845 (I628327,I628842,I628726);
not I_36846 (I628931,I2514);
DFFARX1 I_36847 (I297436,I2507,I628931,I628957,);
and I_36848 (I628965,I628957,I297451);
DFFARX1 I_36849 (I628965,I2507,I628931,I628914,);
DFFARX1 I_36850 (I297442,I2507,I628931,I629005,);
not I_36851 (I629013,I297436);
not I_36852 (I629030,I297454);
nand I_36853 (I629047,I629030,I629013);
nor I_36854 (I628902,I629005,I629047);
DFFARX1 I_36855 (I629047,I2507,I628931,I629087,);
not I_36856 (I628923,I629087);
not I_36857 (I629109,I297445);
nand I_36858 (I629126,I629030,I629109);
DFFARX1 I_36859 (I629126,I2507,I628931,I629152,);
not I_36860 (I629160,I629152);
not I_36861 (I629177,I297457);
nand I_36862 (I629194,I629177,I297433);
and I_36863 (I629211,I629013,I629194);
nor I_36864 (I629228,I629126,I629211);
DFFARX1 I_36865 (I629228,I2507,I628931,I628899,);
DFFARX1 I_36866 (I629211,I2507,I628931,I628920,);
nor I_36867 (I629273,I297457,I297433);
nor I_36868 (I628911,I629126,I629273);
or I_36869 (I629304,I297457,I297433);
nor I_36870 (I629321,I297439,I297448);
DFFARX1 I_36871 (I629321,I2507,I628931,I629347,);
not I_36872 (I629355,I629347);
nor I_36873 (I628917,I629355,I629160);
nand I_36874 (I629386,I629355,I629005);
not I_36875 (I629403,I297439);
nand I_36876 (I629420,I629403,I629109);
nand I_36877 (I629437,I629355,I629420);
nand I_36878 (I628908,I629437,I629386);
nand I_36879 (I628905,I629420,I629304);
not I_36880 (I629509,I2514);
DFFARX1 I_36881 (I511894,I2507,I629509,I629535,);
and I_36882 (I629543,I629535,I511888);
DFFARX1 I_36883 (I629543,I2507,I629509,I629492,);
DFFARX1 I_36884 (I511906,I2507,I629509,I629583,);
not I_36885 (I629591,I511897);
not I_36886 (I629608,I511909);
nand I_36887 (I629625,I629608,I629591);
nor I_36888 (I629480,I629583,I629625);
DFFARX1 I_36889 (I629625,I2507,I629509,I629665,);
not I_36890 (I629501,I629665);
not I_36891 (I629687,I511915);
nand I_36892 (I629704,I629608,I629687);
DFFARX1 I_36893 (I629704,I2507,I629509,I629730,);
not I_36894 (I629738,I629730);
not I_36895 (I629755,I511891);
nand I_36896 (I629772,I629755,I511912);
and I_36897 (I629789,I629591,I629772);
nor I_36898 (I629806,I629704,I629789);
DFFARX1 I_36899 (I629806,I2507,I629509,I629477,);
DFFARX1 I_36900 (I629789,I2507,I629509,I629498,);
nor I_36901 (I629851,I511891,I511903);
nor I_36902 (I629489,I629704,I629851);
or I_36903 (I629882,I511891,I511903);
nor I_36904 (I629899,I511888,I511900);
DFFARX1 I_36905 (I629899,I2507,I629509,I629925,);
not I_36906 (I629933,I629925);
nor I_36907 (I629495,I629933,I629738);
nand I_36908 (I629964,I629933,I629583);
not I_36909 (I629981,I511888);
nand I_36910 (I629998,I629981,I629687);
nand I_36911 (I630015,I629933,I629998);
nand I_36912 (I629486,I630015,I629964);
nand I_36913 (I629483,I629998,I629882);
not I_36914 (I630087,I2514);
DFFARX1 I_36915 (I257432,I2507,I630087,I630113,);
and I_36916 (I630121,I630113,I257447);
DFFARX1 I_36917 (I630121,I2507,I630087,I630070,);
DFFARX1 I_36918 (I257450,I2507,I630087,I630161,);
not I_36919 (I630169,I257444);
not I_36920 (I630186,I257459);
nand I_36921 (I630203,I630186,I630169);
nor I_36922 (I630058,I630161,I630203);
DFFARX1 I_36923 (I630203,I2507,I630087,I630243,);
not I_36924 (I630079,I630243);
not I_36925 (I630265,I257435);
nand I_36926 (I630282,I630186,I630265);
DFFARX1 I_36927 (I630282,I2507,I630087,I630308,);
not I_36928 (I630316,I630308);
not I_36929 (I630333,I257438);
nand I_36930 (I630350,I630333,I257432);
and I_36931 (I630367,I630169,I630350);
nor I_36932 (I630384,I630282,I630367);
DFFARX1 I_36933 (I630384,I2507,I630087,I630055,);
DFFARX1 I_36934 (I630367,I2507,I630087,I630076,);
nor I_36935 (I630429,I257438,I257441);
nor I_36936 (I630067,I630282,I630429);
or I_36937 (I630460,I257438,I257441);
nor I_36938 (I630477,I257456,I257453);
DFFARX1 I_36939 (I630477,I2507,I630087,I630503,);
not I_36940 (I630511,I630503);
nor I_36941 (I630073,I630511,I630316);
nand I_36942 (I630542,I630511,I630161);
not I_36943 (I630559,I257456);
nand I_36944 (I630576,I630559,I630265);
nand I_36945 (I630593,I630511,I630576);
nand I_36946 (I630064,I630593,I630542);
nand I_36947 (I630061,I630576,I630460);
not I_36948 (I630665,I2514);
DFFARX1 I_36949 (I467113,I2507,I630665,I630691,);
and I_36950 (I630699,I630691,I467119);
DFFARX1 I_36951 (I630699,I2507,I630665,I630648,);
DFFARX1 I_36952 (I467125,I2507,I630665,I630739,);
not I_36953 (I630747,I467110);
not I_36954 (I630764,I467110);
nand I_36955 (I630781,I630764,I630747);
nor I_36956 (I630636,I630739,I630781);
DFFARX1 I_36957 (I630781,I2507,I630665,I630821,);
not I_36958 (I630657,I630821);
not I_36959 (I630843,I467128);
nand I_36960 (I630860,I630764,I630843);
DFFARX1 I_36961 (I630860,I2507,I630665,I630886,);
not I_36962 (I630894,I630886);
not I_36963 (I630911,I467122);
nand I_36964 (I630928,I630911,I467113);
and I_36965 (I630945,I630747,I630928);
nor I_36966 (I630962,I630860,I630945);
DFFARX1 I_36967 (I630962,I2507,I630665,I630633,);
DFFARX1 I_36968 (I630945,I2507,I630665,I630654,);
nor I_36969 (I631007,I467122,I467131);
nor I_36970 (I630645,I630860,I631007);
or I_36971 (I631038,I467122,I467131);
nor I_36972 (I631055,I467116,I467116);
DFFARX1 I_36973 (I631055,I2507,I630665,I631081,);
not I_36974 (I631089,I631081);
nor I_36975 (I630651,I631089,I630894);
nand I_36976 (I631120,I631089,I630739);
not I_36977 (I631137,I467116);
nand I_36978 (I631154,I631137,I630843);
nand I_36979 (I631171,I631089,I631154);
nand I_36980 (I630642,I631171,I631120);
nand I_36981 (I630639,I631154,I631038);
not I_36982 (I631243,I2514);
DFFARX1 I_36983 (I376158,I2507,I631243,I631269,);
and I_36984 (I631277,I631269,I376146);
DFFARX1 I_36985 (I631277,I2507,I631243,I631226,);
DFFARX1 I_36986 (I376149,I2507,I631243,I631317,);
not I_36987 (I631325,I376143);
not I_36988 (I631342,I376167);
nand I_36989 (I631359,I631342,I631325);
nor I_36990 (I631214,I631317,I631359);
DFFARX1 I_36991 (I631359,I2507,I631243,I631399,);
not I_36992 (I631235,I631399);
not I_36993 (I631421,I376155);
nand I_36994 (I631438,I631342,I631421);
DFFARX1 I_36995 (I631438,I2507,I631243,I631464,);
not I_36996 (I631472,I631464);
not I_36997 (I631489,I376164);
nand I_36998 (I631506,I631489,I376161);
and I_36999 (I631523,I631325,I631506);
nor I_37000 (I631540,I631438,I631523);
DFFARX1 I_37001 (I631540,I2507,I631243,I631211,);
DFFARX1 I_37002 (I631523,I2507,I631243,I631232,);
nor I_37003 (I631585,I376164,I376152);
nor I_37004 (I631223,I631438,I631585);
or I_37005 (I631616,I376164,I376152);
nor I_37006 (I631633,I376143,I376146);
DFFARX1 I_37007 (I631633,I2507,I631243,I631659,);
not I_37008 (I631667,I631659);
nor I_37009 (I631229,I631667,I631472);
nand I_37010 (I631698,I631667,I631317);
not I_37011 (I631715,I376143);
nand I_37012 (I631732,I631715,I631421);
nand I_37013 (I631749,I631667,I631732);
nand I_37014 (I631220,I631749,I631698);
nand I_37015 (I631217,I631732,I631616);
not I_37016 (I631821,I2514);
DFFARX1 I_37017 (I186433,I2507,I631821,I631847,);
and I_37018 (I631855,I631847,I186418);
DFFARX1 I_37019 (I631855,I2507,I631821,I631804,);
DFFARX1 I_37020 (I186424,I2507,I631821,I631895,);
not I_37021 (I631903,I186406);
not I_37022 (I631920,I186427);
nand I_37023 (I631937,I631920,I631903);
nor I_37024 (I631792,I631895,I631937);
DFFARX1 I_37025 (I631937,I2507,I631821,I631977,);
not I_37026 (I631813,I631977);
not I_37027 (I631999,I186430);
nand I_37028 (I632016,I631920,I631999);
DFFARX1 I_37029 (I632016,I2507,I631821,I632042,);
not I_37030 (I632050,I632042);
not I_37031 (I632067,I186421);
nand I_37032 (I632084,I632067,I186409);
and I_37033 (I632101,I631903,I632084);
nor I_37034 (I632118,I632016,I632101);
DFFARX1 I_37035 (I632118,I2507,I631821,I631789,);
DFFARX1 I_37036 (I632101,I2507,I631821,I631810,);
nor I_37037 (I632163,I186421,I186415);
nor I_37038 (I631801,I632016,I632163);
or I_37039 (I632194,I186421,I186415);
nor I_37040 (I632211,I186412,I186406);
DFFARX1 I_37041 (I632211,I2507,I631821,I632237,);
not I_37042 (I632245,I632237);
nor I_37043 (I631807,I632245,I632050);
nand I_37044 (I632276,I632245,I631895);
not I_37045 (I632293,I186412);
nand I_37046 (I632310,I632293,I631999);
nand I_37047 (I632327,I632245,I632310);
nand I_37048 (I631798,I632327,I632276);
nand I_37049 (I631795,I632310,I632194);
not I_37050 (I632399,I2514);
DFFARX1 I_37051 (I49920,I2507,I632399,I632425,);
and I_37052 (I632433,I632425,I49896);
DFFARX1 I_37053 (I632433,I2507,I632399,I632382,);
DFFARX1 I_37054 (I49914,I2507,I632399,I632473,);
not I_37055 (I632481,I49902);
not I_37056 (I632498,I49899);
nand I_37057 (I632515,I632498,I632481);
nor I_37058 (I632370,I632473,I632515);
DFFARX1 I_37059 (I632515,I2507,I632399,I632555,);
not I_37060 (I632391,I632555);
not I_37061 (I632577,I49908);
nand I_37062 (I632594,I632498,I632577);
DFFARX1 I_37063 (I632594,I2507,I632399,I632620,);
not I_37064 (I632628,I632620);
not I_37065 (I632645,I49899);
nand I_37066 (I632662,I632645,I49917);
and I_37067 (I632679,I632481,I632662);
nor I_37068 (I632696,I632594,I632679);
DFFARX1 I_37069 (I632696,I2507,I632399,I632367,);
DFFARX1 I_37070 (I632679,I2507,I632399,I632388,);
nor I_37071 (I632741,I49899,I49911);
nor I_37072 (I632379,I632594,I632741);
or I_37073 (I632772,I49899,I49911);
nor I_37074 (I632789,I49905,I49896);
DFFARX1 I_37075 (I632789,I2507,I632399,I632815,);
not I_37076 (I632823,I632815);
nor I_37077 (I632385,I632823,I632628);
nand I_37078 (I632854,I632823,I632473);
not I_37079 (I632871,I49905);
nand I_37080 (I632888,I632871,I632577);
nand I_37081 (I632905,I632823,I632888);
nand I_37082 (I632376,I632905,I632854);
nand I_37083 (I632373,I632888,I632772);
not I_37084 (I632977,I2514);
DFFARX1 I_37085 (I417774,I2507,I632977,I633003,);
and I_37086 (I633011,I633003,I417762);
DFFARX1 I_37087 (I633011,I2507,I632977,I632960,);
DFFARX1 I_37088 (I417765,I2507,I632977,I633051,);
not I_37089 (I633059,I417759);
not I_37090 (I633076,I417783);
nand I_37091 (I633093,I633076,I633059);
nor I_37092 (I632948,I633051,I633093);
DFFARX1 I_37093 (I633093,I2507,I632977,I633133,);
not I_37094 (I632969,I633133);
not I_37095 (I633155,I417771);
nand I_37096 (I633172,I633076,I633155);
DFFARX1 I_37097 (I633172,I2507,I632977,I633198,);
not I_37098 (I633206,I633198);
not I_37099 (I633223,I417780);
nand I_37100 (I633240,I633223,I417777);
and I_37101 (I633257,I633059,I633240);
nor I_37102 (I633274,I633172,I633257);
DFFARX1 I_37103 (I633274,I2507,I632977,I632945,);
DFFARX1 I_37104 (I633257,I2507,I632977,I632966,);
nor I_37105 (I633319,I417780,I417768);
nor I_37106 (I632957,I633172,I633319);
or I_37107 (I633350,I417780,I417768);
nor I_37108 (I633367,I417759,I417762);
DFFARX1 I_37109 (I633367,I2507,I632977,I633393,);
not I_37110 (I633401,I633393);
nor I_37111 (I632963,I633401,I633206);
nand I_37112 (I633432,I633401,I633051);
not I_37113 (I633449,I417759);
nand I_37114 (I633466,I633449,I633155);
nand I_37115 (I633483,I633401,I633466);
nand I_37116 (I632954,I633483,I633432);
nand I_37117 (I632951,I633466,I633350);
not I_37118 (I633555,I2514);
DFFARX1 I_37119 (I660506,I2507,I633555,I633581,);
and I_37120 (I633589,I633581,I660500);
DFFARX1 I_37121 (I633589,I2507,I633555,I633538,);
DFFARX1 I_37122 (I660485,I2507,I633555,I633629,);
not I_37123 (I633637,I660491);
not I_37124 (I633654,I660503);
nand I_37125 (I633671,I633654,I633637);
nor I_37126 (I633526,I633629,I633671);
DFFARX1 I_37127 (I633671,I2507,I633555,I633711,);
not I_37128 (I633547,I633711);
not I_37129 (I633733,I660485);
nand I_37130 (I633750,I633654,I633733);
DFFARX1 I_37131 (I633750,I2507,I633555,I633776,);
not I_37132 (I633784,I633776);
not I_37133 (I633801,I660509);
nand I_37134 (I633818,I633801,I660497);
and I_37135 (I633835,I633637,I633818);
nor I_37136 (I633852,I633750,I633835);
DFFARX1 I_37137 (I633852,I2507,I633555,I633523,);
DFFARX1 I_37138 (I633835,I2507,I633555,I633544,);
nor I_37139 (I633897,I660509,I660488);
nor I_37140 (I633535,I633750,I633897);
or I_37141 (I633928,I660509,I660488);
nor I_37142 (I633945,I660494,I660488);
DFFARX1 I_37143 (I633945,I2507,I633555,I633971,);
not I_37144 (I633979,I633971);
nor I_37145 (I633541,I633979,I633784);
nand I_37146 (I634010,I633979,I633629);
not I_37147 (I634027,I660494);
nand I_37148 (I634044,I634027,I633733);
nand I_37149 (I634061,I633979,I634044);
nand I_37150 (I633532,I634061,I634010);
nand I_37151 (I633529,I634044,I633928);
not I_37152 (I634133,I2514);
DFFARX1 I_37153 (I408526,I2507,I634133,I634159,);
and I_37154 (I634167,I634159,I408514);
DFFARX1 I_37155 (I634167,I2507,I634133,I634116,);
DFFARX1 I_37156 (I408517,I2507,I634133,I634207,);
not I_37157 (I634215,I408511);
not I_37158 (I634232,I408535);
nand I_37159 (I634249,I634232,I634215);
nor I_37160 (I634104,I634207,I634249);
DFFARX1 I_37161 (I634249,I2507,I634133,I634289,);
not I_37162 (I634125,I634289);
not I_37163 (I634311,I408523);
nand I_37164 (I634328,I634232,I634311);
DFFARX1 I_37165 (I634328,I2507,I634133,I634354,);
not I_37166 (I634362,I634354);
not I_37167 (I634379,I408532);
nand I_37168 (I634396,I634379,I408529);
and I_37169 (I634413,I634215,I634396);
nor I_37170 (I634430,I634328,I634413);
DFFARX1 I_37171 (I634430,I2507,I634133,I634101,);
DFFARX1 I_37172 (I634413,I2507,I634133,I634122,);
nor I_37173 (I634475,I408532,I408520);
nor I_37174 (I634113,I634328,I634475);
or I_37175 (I634506,I408532,I408520);
nor I_37176 (I634523,I408511,I408514);
DFFARX1 I_37177 (I634523,I2507,I634133,I634549,);
not I_37178 (I634557,I634549);
nor I_37179 (I634119,I634557,I634362);
nand I_37180 (I634588,I634557,I634207);
not I_37181 (I634605,I408511);
nand I_37182 (I634622,I634605,I634311);
nand I_37183 (I634639,I634557,I634622);
nand I_37184 (I634110,I634639,I634588);
nand I_37185 (I634107,I634622,I634506);
not I_37186 (I634711,I2514);
DFFARX1 I_37187 (I92549,I2507,I634711,I634737,);
and I_37188 (I634745,I634737,I92552);
DFFARX1 I_37189 (I634745,I2507,I634711,I634694,);
DFFARX1 I_37190 (I92552,I2507,I634711,I634785,);
not I_37191 (I634793,I92567);
not I_37192 (I634810,I92573);
nand I_37193 (I634827,I634810,I634793);
nor I_37194 (I634682,I634785,I634827);
DFFARX1 I_37195 (I634827,I2507,I634711,I634867,);
not I_37196 (I634703,I634867);
not I_37197 (I634889,I92561);
nand I_37198 (I634906,I634810,I634889);
DFFARX1 I_37199 (I634906,I2507,I634711,I634932,);
not I_37200 (I634940,I634932);
not I_37201 (I634957,I92558);
nand I_37202 (I634974,I634957,I92555);
and I_37203 (I634991,I634793,I634974);
nor I_37204 (I635008,I634906,I634991);
DFFARX1 I_37205 (I635008,I2507,I634711,I634679,);
DFFARX1 I_37206 (I634991,I2507,I634711,I634700,);
nor I_37207 (I635053,I92558,I92549);
nor I_37208 (I634691,I634906,I635053);
or I_37209 (I635084,I92558,I92549);
nor I_37210 (I635101,I92564,I92570);
DFFARX1 I_37211 (I635101,I2507,I634711,I635127,);
not I_37212 (I635135,I635127);
nor I_37213 (I634697,I635135,I634940);
nand I_37214 (I635166,I635135,I634785);
not I_37215 (I635183,I92564);
nand I_37216 (I635200,I635183,I634889);
nand I_37217 (I635217,I635135,I635200);
nand I_37218 (I634688,I635217,I635166);
nand I_37219 (I634685,I635200,I635084);
not I_37220 (I635289,I2514);
DFFARX1 I_37221 (I100879,I2507,I635289,I635315,);
and I_37222 (I635323,I635315,I100882);
DFFARX1 I_37223 (I635323,I2507,I635289,I635272,);
DFFARX1 I_37224 (I100882,I2507,I635289,I635363,);
not I_37225 (I635371,I100897);
not I_37226 (I635388,I100903);
nand I_37227 (I635405,I635388,I635371);
nor I_37228 (I635260,I635363,I635405);
DFFARX1 I_37229 (I635405,I2507,I635289,I635445,);
not I_37230 (I635281,I635445);
not I_37231 (I635467,I100891);
nand I_37232 (I635484,I635388,I635467);
DFFARX1 I_37233 (I635484,I2507,I635289,I635510,);
not I_37234 (I635518,I635510);
not I_37235 (I635535,I100888);
nand I_37236 (I635552,I635535,I100885);
and I_37237 (I635569,I635371,I635552);
nor I_37238 (I635586,I635484,I635569);
DFFARX1 I_37239 (I635586,I2507,I635289,I635257,);
DFFARX1 I_37240 (I635569,I2507,I635289,I635278,);
nor I_37241 (I635631,I100888,I100879);
nor I_37242 (I635269,I635484,I635631);
or I_37243 (I635662,I100888,I100879);
nor I_37244 (I635679,I100894,I100900);
DFFARX1 I_37245 (I635679,I2507,I635289,I635705,);
not I_37246 (I635713,I635705);
nor I_37247 (I635275,I635713,I635518);
nand I_37248 (I635744,I635713,I635363);
not I_37249 (I635761,I100894);
nand I_37250 (I635778,I635761,I635467);
nand I_37251 (I635795,I635713,I635778);
nand I_37252 (I635266,I635795,I635744);
nand I_37253 (I635263,I635778,I635662);
not I_37254 (I635867,I2514);
DFFARX1 I_37255 (I539026,I2507,I635867,I635893,);
and I_37256 (I635901,I635893,I539020);
DFFARX1 I_37257 (I635901,I2507,I635867,I635850,);
DFFARX1 I_37258 (I539038,I2507,I635867,I635941,);
not I_37259 (I635949,I539029);
not I_37260 (I635966,I539041);
nand I_37261 (I635983,I635966,I635949);
nor I_37262 (I635838,I635941,I635983);
DFFARX1 I_37263 (I635983,I2507,I635867,I636023,);
not I_37264 (I635859,I636023);
not I_37265 (I636045,I539047);
nand I_37266 (I636062,I635966,I636045);
DFFARX1 I_37267 (I636062,I2507,I635867,I636088,);
not I_37268 (I636096,I636088);
not I_37269 (I636113,I539023);
nand I_37270 (I636130,I636113,I539044);
and I_37271 (I636147,I635949,I636130);
nor I_37272 (I636164,I636062,I636147);
DFFARX1 I_37273 (I636164,I2507,I635867,I635835,);
DFFARX1 I_37274 (I636147,I2507,I635867,I635856,);
nor I_37275 (I636209,I539023,I539035);
nor I_37276 (I635847,I636062,I636209);
or I_37277 (I636240,I539023,I539035);
nor I_37278 (I636257,I539020,I539032);
DFFARX1 I_37279 (I636257,I2507,I635867,I636283,);
not I_37280 (I636291,I636283);
nor I_37281 (I635853,I636291,I636096);
nand I_37282 (I636322,I636291,I635941);
not I_37283 (I636339,I539020);
nand I_37284 (I636356,I636339,I636045);
nand I_37285 (I636373,I636291,I636356);
nand I_37286 (I635844,I636373,I636322);
nand I_37287 (I635841,I636356,I636240);
not I_37288 (I636445,I2514);
DFFARX1 I_37289 (I60987,I2507,I636445,I636471,);
and I_37290 (I636479,I636471,I60963);
DFFARX1 I_37291 (I636479,I2507,I636445,I636428,);
DFFARX1 I_37292 (I60981,I2507,I636445,I636519,);
not I_37293 (I636527,I60969);
not I_37294 (I636544,I60966);
nand I_37295 (I636561,I636544,I636527);
nor I_37296 (I636416,I636519,I636561);
DFFARX1 I_37297 (I636561,I2507,I636445,I636601,);
not I_37298 (I636437,I636601);
not I_37299 (I636623,I60975);
nand I_37300 (I636640,I636544,I636623);
DFFARX1 I_37301 (I636640,I2507,I636445,I636666,);
not I_37302 (I636674,I636666);
not I_37303 (I636691,I60966);
nand I_37304 (I636708,I636691,I60984);
and I_37305 (I636725,I636527,I636708);
nor I_37306 (I636742,I636640,I636725);
DFFARX1 I_37307 (I636742,I2507,I636445,I636413,);
DFFARX1 I_37308 (I636725,I2507,I636445,I636434,);
nor I_37309 (I636787,I60966,I60978);
nor I_37310 (I636425,I636640,I636787);
or I_37311 (I636818,I60966,I60978);
nor I_37312 (I636835,I60972,I60963);
DFFARX1 I_37313 (I636835,I2507,I636445,I636861,);
not I_37314 (I636869,I636861);
nor I_37315 (I636431,I636869,I636674);
nand I_37316 (I636900,I636869,I636519);
not I_37317 (I636917,I60972);
nand I_37318 (I636934,I636917,I636623);
nand I_37319 (I636951,I636869,I636934);
nand I_37320 (I636422,I636951,I636900);
nand I_37321 (I636419,I636934,I636818);
not I_37322 (I637023,I2514);
DFFARX1 I_37323 (I194338,I2507,I637023,I637049,);
and I_37324 (I637057,I637049,I194323);
DFFARX1 I_37325 (I637057,I2507,I637023,I637006,);
DFFARX1 I_37326 (I194329,I2507,I637023,I637097,);
not I_37327 (I637105,I194311);
not I_37328 (I637122,I194332);
nand I_37329 (I637139,I637122,I637105);
nor I_37330 (I636994,I637097,I637139);
DFFARX1 I_37331 (I637139,I2507,I637023,I637179,);
not I_37332 (I637015,I637179);
not I_37333 (I637201,I194335);
nand I_37334 (I637218,I637122,I637201);
DFFARX1 I_37335 (I637218,I2507,I637023,I637244,);
not I_37336 (I637252,I637244);
not I_37337 (I637269,I194326);
nand I_37338 (I637286,I637269,I194314);
and I_37339 (I637303,I637105,I637286);
nor I_37340 (I637320,I637218,I637303);
DFFARX1 I_37341 (I637320,I2507,I637023,I636991,);
DFFARX1 I_37342 (I637303,I2507,I637023,I637012,);
nor I_37343 (I637365,I194326,I194320);
nor I_37344 (I637003,I637218,I637365);
or I_37345 (I637396,I194326,I194320);
nor I_37346 (I637413,I194317,I194311);
DFFARX1 I_37347 (I637413,I2507,I637023,I637439,);
not I_37348 (I637447,I637439);
nor I_37349 (I637009,I637447,I637252);
nand I_37350 (I637478,I637447,I637097);
not I_37351 (I637495,I194317);
nand I_37352 (I637512,I637495,I637201);
nand I_37353 (I637529,I637447,I637512);
nand I_37354 (I637000,I637529,I637478);
nand I_37355 (I636997,I637512,I637396);
not I_37356 (I637601,I2514);
DFFARX1 I_37357 (I463951,I2507,I637601,I637627,);
and I_37358 (I637635,I637627,I463957);
DFFARX1 I_37359 (I637635,I2507,I637601,I637584,);
DFFARX1 I_37360 (I463963,I2507,I637601,I637675,);
not I_37361 (I637683,I463948);
not I_37362 (I637700,I463948);
nand I_37363 (I637717,I637700,I637683);
nor I_37364 (I637572,I637675,I637717);
DFFARX1 I_37365 (I637717,I2507,I637601,I637757,);
not I_37366 (I637593,I637757);
not I_37367 (I637779,I463966);
nand I_37368 (I637796,I637700,I637779);
DFFARX1 I_37369 (I637796,I2507,I637601,I637822,);
not I_37370 (I637830,I637822);
not I_37371 (I637847,I463960);
nand I_37372 (I637864,I637847,I463951);
and I_37373 (I637881,I637683,I637864);
nor I_37374 (I637898,I637796,I637881);
DFFARX1 I_37375 (I637898,I2507,I637601,I637569,);
DFFARX1 I_37376 (I637881,I2507,I637601,I637590,);
nor I_37377 (I637943,I463960,I463969);
nor I_37378 (I637581,I637796,I637943);
or I_37379 (I637974,I463960,I463969);
nor I_37380 (I637991,I463954,I463954);
DFFARX1 I_37381 (I637991,I2507,I637601,I638017,);
not I_37382 (I638025,I638017);
nor I_37383 (I637587,I638025,I637830);
nand I_37384 (I638056,I638025,I637675);
not I_37385 (I638073,I463954);
nand I_37386 (I638090,I638073,I637779);
nand I_37387 (I638107,I638025,I638090);
nand I_37388 (I637578,I638107,I638056);
nand I_37389 (I637575,I638090,I637974);
not I_37390 (I638179,I2514);
DFFARX1 I_37391 (I236760,I2507,I638179,I638205,);
and I_37392 (I638213,I638205,I236775);
DFFARX1 I_37393 (I638213,I2507,I638179,I638162,);
DFFARX1 I_37394 (I236778,I2507,I638179,I638253,);
not I_37395 (I638261,I236772);
not I_37396 (I638278,I236787);
nand I_37397 (I638295,I638278,I638261);
nor I_37398 (I638150,I638253,I638295);
DFFARX1 I_37399 (I638295,I2507,I638179,I638335,);
not I_37400 (I638171,I638335);
not I_37401 (I638357,I236763);
nand I_37402 (I638374,I638278,I638357);
DFFARX1 I_37403 (I638374,I2507,I638179,I638400,);
not I_37404 (I638408,I638400);
not I_37405 (I638425,I236766);
nand I_37406 (I638442,I638425,I236760);
and I_37407 (I638459,I638261,I638442);
nor I_37408 (I638476,I638374,I638459);
DFFARX1 I_37409 (I638476,I2507,I638179,I638147,);
DFFARX1 I_37410 (I638459,I2507,I638179,I638168,);
nor I_37411 (I638521,I236766,I236769);
nor I_37412 (I638159,I638374,I638521);
or I_37413 (I638552,I236766,I236769);
nor I_37414 (I638569,I236784,I236781);
DFFARX1 I_37415 (I638569,I2507,I638179,I638595,);
not I_37416 (I638603,I638595);
nor I_37417 (I638165,I638603,I638408);
nand I_37418 (I638634,I638603,I638253);
not I_37419 (I638651,I236784);
nand I_37420 (I638668,I638651,I638357);
nand I_37421 (I638685,I638603,I638668);
nand I_37422 (I638156,I638685,I638634);
nand I_37423 (I638153,I638668,I638552);
not I_37424 (I638757,I2514);
DFFARX1 I_37425 (I455522,I2507,I638757,I638783,);
nand I_37426 (I638791,I638783,I455516);
DFFARX1 I_37427 (I455519,I2507,I638757,I638817,);
DFFARX1 I_37428 (I638817,I2507,I638757,I638834,);
not I_37429 (I638749,I638834);
not I_37430 (I638856,I455525);
nor I_37431 (I638873,I455525,I455519);
not I_37432 (I638890,I455528);
nand I_37433 (I638907,I638856,I638890);
nor I_37434 (I638924,I455528,I455525);
and I_37435 (I638728,I638924,I638791);
not I_37436 (I638955,I455537);
nand I_37437 (I638972,I638955,I455531);
nor I_37438 (I638989,I455537,I455534);
not I_37439 (I639006,I638989);
nand I_37440 (I638731,I638873,I639006);
DFFARX1 I_37441 (I638989,I2507,I638757,I638746,);
nor I_37442 (I639051,I455516,I455528);
nor I_37443 (I639068,I639051,I455519);
and I_37444 (I639085,I639068,I638972);
DFFARX1 I_37445 (I639085,I2507,I638757,I638743,);
nor I_37446 (I638740,I639051,I638907);
or I_37447 (I638737,I638989,I639051);
nor I_37448 (I639144,I455516,I455522);
DFFARX1 I_37449 (I639144,I2507,I638757,I639170,);
not I_37450 (I639178,I639170);
nand I_37451 (I639195,I639178,I638856);
nor I_37452 (I639212,I639195,I455519);
DFFARX1 I_37453 (I639212,I2507,I638757,I638725,);
nor I_37454 (I639243,I639178,I638907);
nor I_37455 (I638734,I639051,I639243);
not I_37456 (I639301,I2514);
DFFARX1 I_37457 (I570545,I2507,I639301,I639327,);
nand I_37458 (I639335,I639327,I570524);
DFFARX1 I_37459 (I570521,I2507,I639301,I639361,);
DFFARX1 I_37460 (I639361,I2507,I639301,I639378,);
not I_37461 (I639293,I639378);
not I_37462 (I639400,I570533);
nor I_37463 (I639417,I570533,I570542);
not I_37464 (I639434,I570530);
nand I_37465 (I639451,I639400,I639434);
nor I_37466 (I639468,I570530,I570533);
and I_37467 (I639272,I639468,I639335);
not I_37468 (I639499,I570539);
nand I_37469 (I639516,I639499,I570536);
nor I_37470 (I639533,I570539,I570521);
not I_37471 (I639550,I639533);
nand I_37472 (I639275,I639417,I639550);
DFFARX1 I_37473 (I639533,I2507,I639301,I639290,);
nor I_37474 (I639595,I570524,I570530);
nor I_37475 (I639612,I639595,I570542);
and I_37476 (I639629,I639612,I639516);
DFFARX1 I_37477 (I639629,I2507,I639301,I639287,);
nor I_37478 (I639284,I639595,I639451);
or I_37479 (I639281,I639533,I639595);
nor I_37480 (I639688,I570524,I570527);
DFFARX1 I_37481 (I639688,I2507,I639301,I639714,);
not I_37482 (I639722,I639714);
nand I_37483 (I639739,I639722,I639400);
nor I_37484 (I639756,I639739,I570542);
DFFARX1 I_37485 (I639756,I2507,I639301,I639269,);
nor I_37486 (I639787,I639722,I639451);
nor I_37487 (I639278,I639595,I639787);
not I_37488 (I639845,I2514);
DFFARX1 I_37489 (I506074,I2507,I639845,I639871,);
nand I_37490 (I639879,I639871,I506074);
DFFARX1 I_37491 (I506086,I2507,I639845,I639905,);
DFFARX1 I_37492 (I639905,I2507,I639845,I639922,);
not I_37493 (I639837,I639922);
not I_37494 (I639944,I506080);
nor I_37495 (I639961,I506080,I506101);
not I_37496 (I639978,I506089);
nand I_37497 (I639995,I639944,I639978);
nor I_37498 (I640012,I506089,I506080);
and I_37499 (I639816,I640012,I639879);
not I_37500 (I640043,I506083);
nand I_37501 (I640060,I640043,I506098);
nor I_37502 (I640077,I506083,I506092);
not I_37503 (I640094,I640077);
nand I_37504 (I639819,I639961,I640094);
DFFARX1 I_37505 (I640077,I2507,I639845,I639834,);
nor I_37506 (I640139,I506095,I506089);
nor I_37507 (I640156,I640139,I506101);
and I_37508 (I640173,I640156,I640060);
DFFARX1 I_37509 (I640173,I2507,I639845,I639831,);
nor I_37510 (I639828,I640139,I639995);
or I_37511 (I639825,I640077,I640139);
nor I_37512 (I640232,I506095,I506077);
DFFARX1 I_37513 (I640232,I2507,I639845,I640258,);
not I_37514 (I640266,I640258);
nand I_37515 (I640283,I640266,I639944);
nor I_37516 (I640300,I640283,I506101);
DFFARX1 I_37517 (I640300,I2507,I639845,I639813,);
nor I_37518 (I640331,I640266,I639995);
nor I_37519 (I639822,I640139,I640331);
not I_37520 (I640389,I2514);
DFFARX1 I_37521 (I40431,I2507,I640389,I640415,);
nand I_37522 (I640423,I640415,I40413);
DFFARX1 I_37523 (I40410,I2507,I640389,I640449,);
DFFARX1 I_37524 (I640449,I2507,I640389,I640466,);
not I_37525 (I640381,I640466);
not I_37526 (I640488,I40428);
nor I_37527 (I640505,I40428,I40422);
not I_37528 (I640522,I40410);
nand I_37529 (I640539,I640488,I640522);
nor I_37530 (I640556,I40410,I40428);
and I_37531 (I640360,I640556,I640423);
not I_37532 (I640587,I40419);
nand I_37533 (I640604,I640587,I40425);
nor I_37534 (I640621,I40419,I40413);
not I_37535 (I640638,I640621);
nand I_37536 (I640363,I640505,I640638);
DFFARX1 I_37537 (I640621,I2507,I640389,I640378,);
nor I_37538 (I640683,I40416,I40410);
nor I_37539 (I640700,I640683,I40422);
and I_37540 (I640717,I640700,I640604);
DFFARX1 I_37541 (I640717,I2507,I640389,I640375,);
nor I_37542 (I640372,I640683,I640539);
or I_37543 (I640369,I640621,I640683);
nor I_37544 (I640776,I40416,I40434);
DFFARX1 I_37545 (I640776,I2507,I640389,I640802,);
not I_37546 (I640810,I640802);
nand I_37547 (I640827,I640810,I640488);
nor I_37548 (I640844,I640827,I40422);
DFFARX1 I_37549 (I640844,I2507,I640389,I640357,);
nor I_37550 (I640875,I640810,I640539);
nor I_37551 (I640366,I640683,I640875);
not I_37552 (I640933,I2514);
DFFARX1 I_37553 (I325878,I2507,I640933,I640959,);
nand I_37554 (I640967,I640959,I325866);
DFFARX1 I_37555 (I325872,I2507,I640933,I640993,);
DFFARX1 I_37556 (I640993,I2507,I640933,I641010,);
not I_37557 (I640925,I641010);
not I_37558 (I641032,I325857);
nor I_37559 (I641049,I325857,I325869);
not I_37560 (I641066,I325860);
nand I_37561 (I641083,I641032,I641066);
nor I_37562 (I641100,I325860,I325857);
and I_37563 (I640904,I641100,I640967);
not I_37564 (I641131,I325875);
nand I_37565 (I641148,I641131,I325857);
nor I_37566 (I641165,I325875,I325881);
not I_37567 (I641182,I641165);
nand I_37568 (I640907,I641049,I641182);
DFFARX1 I_37569 (I641165,I2507,I640933,I640922,);
nor I_37570 (I641227,I325863,I325860);
nor I_37571 (I641244,I641227,I325869);
and I_37572 (I641261,I641244,I641148);
DFFARX1 I_37573 (I641261,I2507,I640933,I640919,);
nor I_37574 (I640916,I641227,I641083);
or I_37575 (I640913,I641165,I641227);
nor I_37576 (I641320,I325863,I325860);
DFFARX1 I_37577 (I641320,I2507,I640933,I641346,);
not I_37578 (I641354,I641346);
nand I_37579 (I641371,I641354,I641032);
nor I_37580 (I641388,I641371,I325869);
DFFARX1 I_37581 (I641388,I2507,I640933,I640901,);
nor I_37582 (I641419,I641354,I641083);
nor I_37583 (I640910,I641227,I641419);
not I_37584 (I641477,I2514);
DFFARX1 I_37585 (I564368,I2507,I641477,I641503,);
nand I_37586 (I641511,I641503,I564356);
DFFARX1 I_37587 (I564350,I2507,I641477,I641537,);
DFFARX1 I_37588 (I641537,I2507,I641477,I641554,);
not I_37589 (I641469,I641554);
not I_37590 (I641576,I564350);
nor I_37591 (I641593,I564350,I564362);
not I_37592 (I641610,I564359);
nand I_37593 (I641627,I641576,I641610);
nor I_37594 (I641644,I564359,I564350);
and I_37595 (I641448,I641644,I641511);
not I_37596 (I641675,I564353);
nand I_37597 (I641692,I641675,I564365);
nor I_37598 (I641709,I564353,I564371);
not I_37599 (I641726,I641709);
nand I_37600 (I641451,I641593,I641726);
DFFARX1 I_37601 (I641709,I2507,I641477,I641466,);
nor I_37602 (I641771,I564356,I564359);
nor I_37603 (I641788,I641771,I564362);
and I_37604 (I641805,I641788,I641692);
DFFARX1 I_37605 (I641805,I2507,I641477,I641463,);
nor I_37606 (I641460,I641771,I641627);
or I_37607 (I641457,I641709,I641771);
nor I_37608 (I641864,I564356,I564353);
DFFARX1 I_37609 (I641864,I2507,I641477,I641890,);
not I_37610 (I641898,I641890);
nand I_37611 (I641915,I641898,I641576);
nor I_37612 (I641932,I641915,I564362);
DFFARX1 I_37613 (I641932,I2507,I641477,I641445,);
nor I_37614 (I641963,I641898,I641627);
nor I_37615 (I641454,I641771,I641963);
not I_37616 (I642021,I2514);
DFFARX1 I_37617 (I67835,I2507,I642021,I642047,);
nand I_37618 (I642055,I642047,I67817);
DFFARX1 I_37619 (I67814,I2507,I642021,I642081,);
DFFARX1 I_37620 (I642081,I2507,I642021,I642098,);
not I_37621 (I642013,I642098);
not I_37622 (I642120,I67832);
nor I_37623 (I642137,I67832,I67826);
not I_37624 (I642154,I67814);
nand I_37625 (I642171,I642120,I642154);
nor I_37626 (I642188,I67814,I67832);
and I_37627 (I641992,I642188,I642055);
not I_37628 (I642219,I67823);
nand I_37629 (I642236,I642219,I67829);
nor I_37630 (I642253,I67823,I67817);
not I_37631 (I642270,I642253);
nand I_37632 (I641995,I642137,I642270);
DFFARX1 I_37633 (I642253,I2507,I642021,I642010,);
nor I_37634 (I642315,I67820,I67814);
nor I_37635 (I642332,I642315,I67826);
and I_37636 (I642349,I642332,I642236);
DFFARX1 I_37637 (I642349,I2507,I642021,I642007,);
nor I_37638 (I642004,I642315,I642171);
or I_37639 (I642001,I642253,I642315);
nor I_37640 (I642408,I67820,I67838);
DFFARX1 I_37641 (I642408,I2507,I642021,I642434,);
not I_37642 (I642442,I642434);
nand I_37643 (I642459,I642442,I642120);
nor I_37644 (I642476,I642459,I67826);
DFFARX1 I_37645 (I642476,I2507,I642021,I641989,);
nor I_37646 (I642507,I642442,I642171);
nor I_37647 (I641998,I642315,I642507);
not I_37648 (I642565,I2514);
DFFARX1 I_37649 (I208552,I2507,I642565,I642591,);
nand I_37650 (I642599,I642591,I208555);
DFFARX1 I_37651 (I208549,I2507,I642565,I642625,);
DFFARX1 I_37652 (I642625,I2507,I642565,I642642,);
not I_37653 (I642557,I642642);
not I_37654 (I642664,I208558);
nor I_37655 (I642681,I208558,I208543);
not I_37656 (I642698,I208567);
nand I_37657 (I642715,I642664,I642698);
nor I_37658 (I642732,I208567,I208558);
and I_37659 (I642536,I642732,I642599);
not I_37660 (I642763,I208546);
nand I_37661 (I642780,I642763,I208564);
nor I_37662 (I642797,I208546,I208540);
not I_37663 (I642814,I642797);
nand I_37664 (I642539,I642681,I642814);
DFFARX1 I_37665 (I642797,I2507,I642565,I642554,);
nor I_37666 (I642859,I208561,I208567);
nor I_37667 (I642876,I642859,I208543);
and I_37668 (I642893,I642876,I642780);
DFFARX1 I_37669 (I642893,I2507,I642565,I642551,);
nor I_37670 (I642548,I642859,I642715);
or I_37671 (I642545,I642797,I642859);
nor I_37672 (I642952,I208561,I208540);
DFFARX1 I_37673 (I642952,I2507,I642565,I642978,);
not I_37674 (I642986,I642978);
nand I_37675 (I643003,I642986,I642664);
nor I_37676 (I643020,I643003,I208543);
DFFARX1 I_37677 (I643020,I2507,I642565,I642533,);
nor I_37678 (I643051,I642986,I642715);
nor I_37679 (I642542,I642859,I643051);
not I_37680 (I643109,I2514);
DFFARX1 I_37681 (I417184,I2507,I643109,I643135,);
nand I_37682 (I643143,I643135,I417199);
DFFARX1 I_37683 (I417193,I2507,I643109,I643169,);
DFFARX1 I_37684 (I643169,I2507,I643109,I643186,);
not I_37685 (I643101,I643186);
not I_37686 (I643208,I417196);
nor I_37687 (I643225,I417196,I417202);
not I_37688 (I643242,I417184);
nand I_37689 (I643259,I643208,I643242);
nor I_37690 (I643276,I417184,I417196);
and I_37691 (I643080,I643276,I643143);
not I_37692 (I643307,I417181);
nand I_37693 (I643324,I643307,I417187);
nor I_37694 (I643341,I417181,I417181);
not I_37695 (I643358,I643341);
nand I_37696 (I643083,I643225,I643358);
DFFARX1 I_37697 (I643341,I2507,I643109,I643098,);
nor I_37698 (I643403,I417190,I417184);
nor I_37699 (I643420,I643403,I417202);
and I_37700 (I643437,I643420,I643324);
DFFARX1 I_37701 (I643437,I2507,I643109,I643095,);
nor I_37702 (I643092,I643403,I643259);
or I_37703 (I643089,I643341,I643403);
nor I_37704 (I643496,I417190,I417205);
DFFARX1 I_37705 (I643496,I2507,I643109,I643522,);
not I_37706 (I643530,I643522);
nand I_37707 (I643547,I643530,I643208);
nor I_37708 (I643564,I643547,I417202);
DFFARX1 I_37709 (I643564,I2507,I643109,I643077,);
nor I_37710 (I643595,I643530,I643259);
nor I_37711 (I643086,I643403,I643595);
not I_37712 (I643653,I2514);
DFFARX1 I_37713 (I34634,I2507,I643653,I643679,);
nand I_37714 (I643687,I643679,I34616);
DFFARX1 I_37715 (I34613,I2507,I643653,I643713,);
DFFARX1 I_37716 (I643713,I2507,I643653,I643730,);
not I_37717 (I643645,I643730);
not I_37718 (I643752,I34631);
nor I_37719 (I643769,I34631,I34625);
not I_37720 (I643786,I34613);
nand I_37721 (I643803,I643752,I643786);
nor I_37722 (I643820,I34613,I34631);
and I_37723 (I643624,I643820,I643687);
not I_37724 (I643851,I34622);
nand I_37725 (I643868,I643851,I34628);
nor I_37726 (I643885,I34622,I34616);
not I_37727 (I643902,I643885);
nand I_37728 (I643627,I643769,I643902);
DFFARX1 I_37729 (I643885,I2507,I643653,I643642,);
nor I_37730 (I643947,I34619,I34613);
nor I_37731 (I643964,I643947,I34625);
and I_37732 (I643981,I643964,I643868);
DFFARX1 I_37733 (I643981,I2507,I643653,I643639,);
nor I_37734 (I643636,I643947,I643803);
or I_37735 (I643633,I643885,I643947);
nor I_37736 (I644040,I34619,I34637);
DFFARX1 I_37737 (I644040,I2507,I643653,I644066,);
not I_37738 (I644074,I644066);
nand I_37739 (I644091,I644074,I643752);
nor I_37740 (I644108,I644091,I34625);
DFFARX1 I_37741 (I644108,I2507,I643653,I643621,);
nor I_37742 (I644139,I644074,I643803);
nor I_37743 (I643630,I643947,I644139);
not I_37744 (I644197,I2514);
DFFARX1 I_37745 (I722205,I2507,I644197,I644223,);
nand I_37746 (I644231,I644223,I722190);
DFFARX1 I_37747 (I722184,I2507,I644197,I644257,);
DFFARX1 I_37748 (I644257,I2507,I644197,I644274,);
not I_37749 (I644189,I644274);
not I_37750 (I644296,I722178);
nor I_37751 (I644313,I722178,I722199);
not I_37752 (I644330,I722187);
nand I_37753 (I644347,I644296,I644330);
nor I_37754 (I644364,I722187,I722178);
and I_37755 (I644168,I644364,I644231);
not I_37756 (I644395,I722196);
nand I_37757 (I644412,I644395,I722202);
nor I_37758 (I644429,I722196,I722193);
not I_37759 (I644446,I644429);
nand I_37760 (I644171,I644313,I644446);
DFFARX1 I_37761 (I644429,I2507,I644197,I644186,);
nor I_37762 (I644491,I722181,I722187);
nor I_37763 (I644508,I644491,I722199);
and I_37764 (I644525,I644508,I644412);
DFFARX1 I_37765 (I644525,I2507,I644197,I644183,);
nor I_37766 (I644180,I644491,I644347);
or I_37767 (I644177,I644429,I644491);
nor I_37768 (I644584,I722181,I722178);
DFFARX1 I_37769 (I644584,I2507,I644197,I644610,);
not I_37770 (I644618,I644610);
nand I_37771 (I644635,I644618,I644296);
nor I_37772 (I644652,I644635,I722199);
DFFARX1 I_37773 (I644652,I2507,I644197,I644165,);
nor I_37774 (I644683,I644618,I644347);
nor I_37775 (I644174,I644491,I644683);
not I_37776 (I644741,I2514);
DFFARX1 I_37777 (I219619,I2507,I644741,I644767,);
nand I_37778 (I644775,I644767,I219622);
DFFARX1 I_37779 (I219616,I2507,I644741,I644801,);
DFFARX1 I_37780 (I644801,I2507,I644741,I644818,);
not I_37781 (I644733,I644818);
not I_37782 (I644840,I219625);
nor I_37783 (I644857,I219625,I219610);
not I_37784 (I644874,I219634);
nand I_37785 (I644891,I644840,I644874);
nor I_37786 (I644908,I219634,I219625);
and I_37787 (I644712,I644908,I644775);
not I_37788 (I644939,I219613);
nand I_37789 (I644956,I644939,I219631);
nor I_37790 (I644973,I219613,I219607);
not I_37791 (I644990,I644973);
nand I_37792 (I644715,I644857,I644990);
DFFARX1 I_37793 (I644973,I2507,I644741,I644730,);
nor I_37794 (I645035,I219628,I219634);
nor I_37795 (I645052,I645035,I219610);
and I_37796 (I645069,I645052,I644956);
DFFARX1 I_37797 (I645069,I2507,I644741,I644727,);
nor I_37798 (I644724,I645035,I644891);
or I_37799 (I644721,I644973,I645035);
nor I_37800 (I645128,I219628,I219607);
DFFARX1 I_37801 (I645128,I2507,I644741,I645154,);
not I_37802 (I645162,I645154);
nand I_37803 (I645179,I645162,I644840);
nor I_37804 (I645196,I645179,I219610);
DFFARX1 I_37805 (I645196,I2507,I644741,I644709,);
nor I_37806 (I645227,I645162,I644891);
nor I_37807 (I644718,I645035,I645227);
not I_37808 (I645285,I2514);
DFFARX1 I_37809 (I554831,I2507,I645285,I645311,);
nand I_37810 (I645319,I645311,I554819);
DFFARX1 I_37811 (I554813,I2507,I645285,I645345,);
DFFARX1 I_37812 (I645345,I2507,I645285,I645362,);
not I_37813 (I645277,I645362);
not I_37814 (I645384,I554813);
nor I_37815 (I645401,I554813,I554825);
not I_37816 (I645418,I554822);
nand I_37817 (I645435,I645384,I645418);
nor I_37818 (I645452,I554822,I554813);
and I_37819 (I645256,I645452,I645319);
not I_37820 (I645483,I554816);
nand I_37821 (I645500,I645483,I554828);
nor I_37822 (I645517,I554816,I554834);
not I_37823 (I645534,I645517);
nand I_37824 (I645259,I645401,I645534);
DFFARX1 I_37825 (I645517,I2507,I645285,I645274,);
nor I_37826 (I645579,I554819,I554822);
nor I_37827 (I645596,I645579,I554825);
and I_37828 (I645613,I645596,I645500);
DFFARX1 I_37829 (I645613,I2507,I645285,I645271,);
nor I_37830 (I645268,I645579,I645435);
or I_37831 (I645265,I645517,I645579);
nor I_37832 (I645672,I554819,I554816);
DFFARX1 I_37833 (I645672,I2507,I645285,I645698,);
not I_37834 (I645706,I645698);
nand I_37835 (I645723,I645706,I645384);
nor I_37836 (I645740,I645723,I554825);
DFFARX1 I_37837 (I645740,I2507,I645285,I645253,);
nor I_37838 (I645771,I645706,I645435);
nor I_37839 (I645262,I645579,I645771);
not I_37840 (I645829,I2514);
DFFARX1 I_37841 (I57822,I2507,I645829,I645855,);
nand I_37842 (I645863,I645855,I57804);
DFFARX1 I_37843 (I57801,I2507,I645829,I645889,);
DFFARX1 I_37844 (I645889,I2507,I645829,I645906,);
not I_37845 (I645821,I645906);
not I_37846 (I645928,I57819);
nor I_37847 (I645945,I57819,I57813);
not I_37848 (I645962,I57801);
nand I_37849 (I645979,I645928,I645962);
nor I_37850 (I645996,I57801,I57819);
and I_37851 (I645800,I645996,I645863);
not I_37852 (I646027,I57810);
nand I_37853 (I646044,I646027,I57816);
nor I_37854 (I646061,I57810,I57804);
not I_37855 (I646078,I646061);
nand I_37856 (I645803,I645945,I646078);
DFFARX1 I_37857 (I646061,I2507,I645829,I645818,);
nor I_37858 (I646123,I57807,I57801);
nor I_37859 (I646140,I646123,I57813);
and I_37860 (I646157,I646140,I646044);
DFFARX1 I_37861 (I646157,I2507,I645829,I645815,);
nor I_37862 (I645812,I646123,I645979);
or I_37863 (I645809,I646061,I646123);
nor I_37864 (I646216,I57807,I57825);
DFFARX1 I_37865 (I646216,I2507,I645829,I646242,);
not I_37866 (I646250,I646242);
nand I_37867 (I646267,I646250,I645928);
nor I_37868 (I646284,I646267,I57813);
DFFARX1 I_37869 (I646284,I2507,I645829,I645797,);
nor I_37870 (I646315,I646250,I645979);
nor I_37871 (I645806,I646123,I646315);
not I_37872 (I646373,I2514);
DFFARX1 I_37873 (I600023,I2507,I646373,I646399,);
nand I_37874 (I646407,I646399,I600002);
DFFARX1 I_37875 (I599999,I2507,I646373,I646433,);
DFFARX1 I_37876 (I646433,I2507,I646373,I646450,);
not I_37877 (I646365,I646450);
not I_37878 (I646472,I600011);
nor I_37879 (I646489,I600011,I600020);
not I_37880 (I646506,I600008);
nand I_37881 (I646523,I646472,I646506);
nor I_37882 (I646540,I600008,I600011);
and I_37883 (I646344,I646540,I646407);
not I_37884 (I646571,I600017);
nand I_37885 (I646588,I646571,I600014);
nor I_37886 (I646605,I600017,I599999);
not I_37887 (I646622,I646605);
nand I_37888 (I646347,I646489,I646622);
DFFARX1 I_37889 (I646605,I2507,I646373,I646362,);
nor I_37890 (I646667,I600002,I600008);
nor I_37891 (I646684,I646667,I600020);
and I_37892 (I646701,I646684,I646588);
DFFARX1 I_37893 (I646701,I2507,I646373,I646359,);
nor I_37894 (I646356,I646667,I646523);
or I_37895 (I646353,I646605,I646667);
nor I_37896 (I646760,I600002,I600005);
DFFARX1 I_37897 (I646760,I2507,I646373,I646786,);
not I_37898 (I646794,I646786);
nand I_37899 (I646811,I646794,I646472);
nor I_37900 (I646828,I646811,I600020);
DFFARX1 I_37901 (I646828,I2507,I646373,I646341,);
nor I_37902 (I646859,I646794,I646523);
nor I_37903 (I646350,I646667,I646859);
not I_37904 (I646917,I2514);
DFFARX1 I_37905 (I354760,I2507,I646917,I646943,);
nand I_37906 (I646951,I646943,I354775);
DFFARX1 I_37907 (I354769,I2507,I646917,I646977,);
DFFARX1 I_37908 (I646977,I2507,I646917,I646994,);
not I_37909 (I646909,I646994);
not I_37910 (I647016,I354772);
nor I_37911 (I647033,I354772,I354778);
not I_37912 (I647050,I354760);
nand I_37913 (I647067,I647016,I647050);
nor I_37914 (I647084,I354760,I354772);
and I_37915 (I646888,I647084,I646951);
not I_37916 (I647115,I354757);
nand I_37917 (I647132,I647115,I354763);
nor I_37918 (I647149,I354757,I354757);
not I_37919 (I647166,I647149);
nand I_37920 (I646891,I647033,I647166);
DFFARX1 I_37921 (I647149,I2507,I646917,I646906,);
nor I_37922 (I647211,I354766,I354760);
nor I_37923 (I647228,I647211,I354778);
and I_37924 (I647245,I647228,I647132);
DFFARX1 I_37925 (I647245,I2507,I646917,I646903,);
nor I_37926 (I646900,I647211,I647067);
or I_37927 (I646897,I647149,I647211);
nor I_37928 (I647304,I354766,I354781);
DFFARX1 I_37929 (I647304,I2507,I646917,I647330,);
not I_37930 (I647338,I647330);
nand I_37931 (I647355,I647338,I647016);
nor I_37932 (I647372,I647355,I354778);
DFFARX1 I_37933 (I647372,I2507,I646917,I646885,);
nor I_37934 (I647403,I647338,I647067);
nor I_37935 (I646894,I647211,I647403);
not I_37936 (I647461,I2514);
DFFARX1 I_37937 (I601757,I2507,I647461,I647487,);
nand I_37938 (I647495,I647487,I601736);
DFFARX1 I_37939 (I601733,I2507,I647461,I647521,);
DFFARX1 I_37940 (I647521,I2507,I647461,I647538,);
not I_37941 (I647453,I647538);
not I_37942 (I647560,I601745);
nor I_37943 (I647577,I601745,I601754);
not I_37944 (I647594,I601742);
nand I_37945 (I647611,I647560,I647594);
nor I_37946 (I647628,I601742,I601745);
and I_37947 (I647432,I647628,I647495);
not I_37948 (I647659,I601751);
nand I_37949 (I647676,I647659,I601748);
nor I_37950 (I647693,I601751,I601733);
not I_37951 (I647710,I647693);
nand I_37952 (I647435,I647577,I647710);
DFFARX1 I_37953 (I647693,I2507,I647461,I647450,);
nor I_37954 (I647755,I601736,I601742);
nor I_37955 (I647772,I647755,I601754);
and I_37956 (I647789,I647772,I647676);
DFFARX1 I_37957 (I647789,I2507,I647461,I647447,);
nor I_37958 (I647444,I647755,I647611);
or I_37959 (I647441,I647693,I647755);
nor I_37960 (I647848,I601736,I601739);
DFFARX1 I_37961 (I647848,I2507,I647461,I647874,);
not I_37962 (I647882,I647874);
nand I_37963 (I647899,I647882,I647560);
nor I_37964 (I647916,I647899,I601754);
DFFARX1 I_37965 (I647916,I2507,I647461,I647429,);
nor I_37966 (I647947,I647882,I647611);
nor I_37967 (I647438,I647755,I647947);
not I_37968 (I648005,I2514);
DFFARX1 I_37969 (I160983,I2507,I648005,I648031,);
nand I_37970 (I648039,I648031,I160998);
DFFARX1 I_37971 (I160995,I2507,I648005,I648065,);
DFFARX1 I_37972 (I648065,I2507,I648005,I648082,);
not I_37973 (I647997,I648082);
not I_37974 (I648104,I160974);
nor I_37975 (I648121,I160974,I160980);
not I_37976 (I648138,I160986);
nand I_37977 (I648155,I648104,I648138);
nor I_37978 (I648172,I160986,I160974);
and I_37979 (I647976,I648172,I648039);
not I_37980 (I648203,I160992);
nand I_37981 (I648220,I648203,I160974);
nor I_37982 (I648237,I160992,I160977);
not I_37983 (I648254,I648237);
nand I_37984 (I647979,I648121,I648254);
DFFARX1 I_37985 (I648237,I2507,I648005,I647994,);
nor I_37986 (I648299,I160977,I160986);
nor I_37987 (I648316,I648299,I160980);
and I_37988 (I648333,I648316,I648220);
DFFARX1 I_37989 (I648333,I2507,I648005,I647991,);
nor I_37990 (I647988,I648299,I648155);
or I_37991 (I647985,I648237,I648299);
nor I_37992 (I648392,I160977,I160989);
DFFARX1 I_37993 (I648392,I2507,I648005,I648418,);
not I_37994 (I648426,I648418);
nand I_37995 (I648443,I648426,I648104);
nor I_37996 (I648460,I648443,I160980);
DFFARX1 I_37997 (I648460,I2507,I648005,I647973,);
nor I_37998 (I648491,I648426,I648155);
nor I_37999 (I647982,I648299,I648491);
not I_38000 (I648549,I2514);
DFFARX1 I_38001 (I579215,I2507,I648549,I648575,);
nand I_38002 (I648583,I648575,I579194);
DFFARX1 I_38003 (I579191,I2507,I648549,I648609,);
DFFARX1 I_38004 (I648609,I2507,I648549,I648626,);
not I_38005 (I648541,I648626);
not I_38006 (I648648,I579203);
nor I_38007 (I648665,I579203,I579212);
not I_38008 (I648682,I579200);
nand I_38009 (I648699,I648648,I648682);
nor I_38010 (I648716,I579200,I579203);
and I_38011 (I648520,I648716,I648583);
not I_38012 (I648747,I579209);
nand I_38013 (I648764,I648747,I579206);
nor I_38014 (I648781,I579209,I579191);
not I_38015 (I648798,I648781);
nand I_38016 (I648523,I648665,I648798);
DFFARX1 I_38017 (I648781,I2507,I648549,I648538,);
nor I_38018 (I648843,I579194,I579200);
nor I_38019 (I648860,I648843,I579212);
and I_38020 (I648877,I648860,I648764);
DFFARX1 I_38021 (I648877,I2507,I648549,I648535,);
nor I_38022 (I648532,I648843,I648699);
or I_38023 (I648529,I648781,I648843);
nor I_38024 (I648936,I579194,I579197);
DFFARX1 I_38025 (I648936,I2507,I648549,I648962,);
not I_38026 (I648970,I648962);
nand I_38027 (I648987,I648970,I648648);
nor I_38028 (I649004,I648987,I579212);
DFFARX1 I_38029 (I649004,I2507,I648549,I648517,);
nor I_38030 (I649035,I648970,I648699);
nor I_38031 (I648526,I648843,I649035);
not I_38032 (I649093,I2514);
DFFARX1 I_38033 (I459211,I2507,I649093,I649119,);
nand I_38034 (I649127,I649119,I459205);
DFFARX1 I_38035 (I459208,I2507,I649093,I649153,);
DFFARX1 I_38036 (I649153,I2507,I649093,I649170,);
not I_38037 (I649085,I649170);
not I_38038 (I649192,I459214);
nor I_38039 (I649209,I459214,I459208);
not I_38040 (I649226,I459217);
nand I_38041 (I649243,I649192,I649226);
nor I_38042 (I649260,I459217,I459214);
and I_38043 (I649064,I649260,I649127);
not I_38044 (I649291,I459226);
nand I_38045 (I649308,I649291,I459220);
nor I_38046 (I649325,I459226,I459223);
not I_38047 (I649342,I649325);
nand I_38048 (I649067,I649209,I649342);
DFFARX1 I_38049 (I649325,I2507,I649093,I649082,);
nor I_38050 (I649387,I459205,I459217);
nor I_38051 (I649404,I649387,I459208);
and I_38052 (I649421,I649404,I649308);
DFFARX1 I_38053 (I649421,I2507,I649093,I649079,);
nor I_38054 (I649076,I649387,I649243);
or I_38055 (I649073,I649325,I649387);
nor I_38056 (I649480,I459205,I459211);
DFFARX1 I_38057 (I649480,I2507,I649093,I649506,);
not I_38058 (I649514,I649506);
nand I_38059 (I649531,I649514,I649192);
nor I_38060 (I649548,I649531,I459208);
DFFARX1 I_38061 (I649548,I2507,I649093,I649061,);
nor I_38062 (I649579,I649514,I649243);
nor I_38063 (I649070,I649387,I649579);
not I_38064 (I649637,I2514);
DFFARX1 I_38065 (I33041,I2507,I649637,I649663,);
nand I_38066 (I649671,I649663,I33035);
DFFARX1 I_38067 (I33056,I2507,I649637,I649697,);
DFFARX1 I_38068 (I649697,I2507,I649637,I649714,);
not I_38069 (I649629,I649714);
not I_38070 (I649736,I33044);
nor I_38071 (I649753,I33044,I33053);
not I_38072 (I649770,I33032);
nand I_38073 (I649787,I649736,I649770);
nor I_38074 (I649804,I33032,I33044);
and I_38075 (I649608,I649804,I649671);
not I_38076 (I649835,I33050);
nand I_38077 (I649852,I649835,I33038);
nor I_38078 (I649869,I33050,I33032);
not I_38079 (I649886,I649869);
nand I_38080 (I649611,I649753,I649886);
DFFARX1 I_38081 (I649869,I2507,I649637,I649626,);
nor I_38082 (I649931,I33035,I33032);
nor I_38083 (I649948,I649931,I33053);
and I_38084 (I649965,I649948,I649852);
DFFARX1 I_38085 (I649965,I2507,I649637,I649623,);
nor I_38086 (I649620,I649931,I649787);
or I_38087 (I649617,I649869,I649931);
nor I_38088 (I650024,I33035,I33047);
DFFARX1 I_38089 (I650024,I2507,I649637,I650050,);
not I_38090 (I650058,I650050);
nand I_38091 (I650075,I650058,I649736);
nor I_38092 (I650092,I650075,I33053);
DFFARX1 I_38093 (I650092,I2507,I649637,I649605,);
nor I_38094 (I650123,I650058,I649787);
nor I_38095 (I649614,I649931,I650123);
not I_38096 (I650181,I2514);
DFFARX1 I_38097 (I316630,I2507,I650181,I650207,);
nand I_38098 (I650215,I650207,I316618);
DFFARX1 I_38099 (I316624,I2507,I650181,I650241,);
DFFARX1 I_38100 (I650241,I2507,I650181,I650258,);
not I_38101 (I650173,I650258);
not I_38102 (I650280,I316609);
nor I_38103 (I650297,I316609,I316621);
not I_38104 (I650314,I316612);
nand I_38105 (I650331,I650280,I650314);
nor I_38106 (I650348,I316612,I316609);
and I_38107 (I650152,I650348,I650215);
not I_38108 (I650379,I316627);
nand I_38109 (I650396,I650379,I316609);
nor I_38110 (I650413,I316627,I316633);
not I_38111 (I650430,I650413);
nand I_38112 (I650155,I650297,I650430);
DFFARX1 I_38113 (I650413,I2507,I650181,I650170,);
nor I_38114 (I650475,I316615,I316612);
nor I_38115 (I650492,I650475,I316621);
and I_38116 (I650509,I650492,I650396);
DFFARX1 I_38117 (I650509,I2507,I650181,I650167,);
nor I_38118 (I650164,I650475,I650331);
or I_38119 (I650161,I650413,I650475);
nor I_38120 (I650568,I316615,I316612);
DFFARX1 I_38121 (I650568,I2507,I650181,I650594,);
not I_38122 (I650602,I650594);
nand I_38123 (I650619,I650602,I650280);
nor I_38124 (I650636,I650619,I316621);
DFFARX1 I_38125 (I650636,I2507,I650181,I650149,);
nor I_38126 (I650667,I650602,I650331);
nor I_38127 (I650158,I650475,I650667);
not I_38128 (I650725,I2514);
DFFARX1 I_38129 (I374990,I2507,I650725,I650751,);
nand I_38130 (I650759,I650751,I375005);
DFFARX1 I_38131 (I374999,I2507,I650725,I650785,);
DFFARX1 I_38132 (I650785,I2507,I650725,I650802,);
not I_38133 (I650717,I650802);
not I_38134 (I650824,I375002);
nor I_38135 (I650841,I375002,I375008);
not I_38136 (I650858,I374990);
nand I_38137 (I650875,I650824,I650858);
nor I_38138 (I650892,I374990,I375002);
and I_38139 (I650696,I650892,I650759);
not I_38140 (I650923,I374987);
nand I_38141 (I650940,I650923,I374993);
nor I_38142 (I650957,I374987,I374987);
not I_38143 (I650974,I650957);
nand I_38144 (I650699,I650841,I650974);
DFFARX1 I_38145 (I650957,I2507,I650725,I650714,);
nor I_38146 (I651019,I374996,I374990);
nor I_38147 (I651036,I651019,I375008);
and I_38148 (I651053,I651036,I650940);
DFFARX1 I_38149 (I651053,I2507,I650725,I650711,);
nor I_38150 (I650708,I651019,I650875);
or I_38151 (I650705,I650957,I651019);
nor I_38152 (I651112,I374996,I375011);
DFFARX1 I_38153 (I651112,I2507,I650725,I651138,);
not I_38154 (I651146,I651138);
nand I_38155 (I651163,I651146,I650824);
nor I_38156 (I651180,I651163,I375008);
DFFARX1 I_38157 (I651180,I2507,I650725,I650693,);
nor I_38158 (I651211,I651146,I650875);
nor I_38159 (I650702,I651019,I651211);
not I_38160 (I651269,I2514);
DFFARX1 I_38161 (I731725,I2507,I651269,I651295,);
nand I_38162 (I651303,I651295,I731710);
DFFARX1 I_38163 (I731704,I2507,I651269,I651329,);
DFFARX1 I_38164 (I651329,I2507,I651269,I651346,);
not I_38165 (I651261,I651346);
not I_38166 (I651368,I731698);
nor I_38167 (I651385,I731698,I731719);
not I_38168 (I651402,I731707);
nand I_38169 (I651419,I651368,I651402);
nor I_38170 (I651436,I731707,I731698);
and I_38171 (I651240,I651436,I651303);
not I_38172 (I651467,I731716);
nand I_38173 (I651484,I651467,I731722);
nor I_38174 (I651501,I731716,I731713);
not I_38175 (I651518,I651501);
nand I_38176 (I651243,I651385,I651518);
DFFARX1 I_38177 (I651501,I2507,I651269,I651258,);
nor I_38178 (I651563,I731701,I731707);
nor I_38179 (I651580,I651563,I731719);
and I_38180 (I651597,I651580,I651484);
DFFARX1 I_38181 (I651597,I2507,I651269,I651255,);
nor I_38182 (I651252,I651563,I651419);
or I_38183 (I651249,I651501,I651563);
nor I_38184 (I651656,I731701,I731698);
DFFARX1 I_38185 (I651656,I2507,I651269,I651682,);
not I_38186 (I651690,I651682);
nand I_38187 (I651707,I651690,I651368);
nor I_38188 (I651724,I651707,I731719);
DFFARX1 I_38189 (I651724,I2507,I651269,I651237,);
nor I_38190 (I651755,I651690,I651419);
nor I_38191 (I651246,I651563,I651755);
not I_38192 (I651813,I2514);
DFFARX1 I_38193 (I219092,I2507,I651813,I651839,);
nand I_38194 (I651847,I651839,I219095);
DFFARX1 I_38195 (I219089,I2507,I651813,I651873,);
DFFARX1 I_38196 (I651873,I2507,I651813,I651890,);
not I_38197 (I651805,I651890);
not I_38198 (I651912,I219098);
nor I_38199 (I651929,I219098,I219083);
not I_38200 (I651946,I219107);
nand I_38201 (I651963,I651912,I651946);
nor I_38202 (I651980,I219107,I219098);
and I_38203 (I651784,I651980,I651847);
not I_38204 (I652011,I219086);
nand I_38205 (I652028,I652011,I219104);
nor I_38206 (I652045,I219086,I219080);
not I_38207 (I652062,I652045);
nand I_38208 (I651787,I651929,I652062);
DFFARX1 I_38209 (I652045,I2507,I651813,I651802,);
nor I_38210 (I652107,I219101,I219107);
nor I_38211 (I652124,I652107,I219083);
and I_38212 (I652141,I652124,I652028);
DFFARX1 I_38213 (I652141,I2507,I651813,I651799,);
nor I_38214 (I651796,I652107,I651963);
or I_38215 (I651793,I652045,I652107);
nor I_38216 (I652200,I219101,I219080);
DFFARX1 I_38217 (I652200,I2507,I651813,I652226,);
not I_38218 (I652234,I652226);
nand I_38219 (I652251,I652234,I651912);
nor I_38220 (I652268,I652251,I219083);
DFFARX1 I_38221 (I652268,I2507,I651813,I651781,);
nor I_38222 (I652299,I652234,I651963);
nor I_38223 (I651790,I652107,I652299);
not I_38224 (I652357,I2514);
DFFARX1 I_38225 (I488632,I2507,I652357,I652383,);
nand I_38226 (I652391,I652383,I488632);
DFFARX1 I_38227 (I488644,I2507,I652357,I652417,);
DFFARX1 I_38228 (I652417,I2507,I652357,I652434,);
not I_38229 (I652349,I652434);
not I_38230 (I652456,I488638);
nor I_38231 (I652473,I488638,I488659);
not I_38232 (I652490,I488647);
nand I_38233 (I652507,I652456,I652490);
nor I_38234 (I652524,I488647,I488638);
and I_38235 (I652328,I652524,I652391);
not I_38236 (I652555,I488641);
nand I_38237 (I652572,I652555,I488656);
nor I_38238 (I652589,I488641,I488650);
not I_38239 (I652606,I652589);
nand I_38240 (I652331,I652473,I652606);
DFFARX1 I_38241 (I652589,I2507,I652357,I652346,);
nor I_38242 (I652651,I488653,I488647);
nor I_38243 (I652668,I652651,I488659);
and I_38244 (I652685,I652668,I652572);
DFFARX1 I_38245 (I652685,I2507,I652357,I652343,);
nor I_38246 (I652340,I652651,I652507);
or I_38247 (I652337,I652589,I652651);
nor I_38248 (I652744,I488653,I488635);
DFFARX1 I_38249 (I652744,I2507,I652357,I652770,);
not I_38250 (I652778,I652770);
nand I_38251 (I652795,I652778,I652456);
nor I_38252 (I652812,I652795,I488659);
DFFARX1 I_38253 (I652812,I2507,I652357,I652325,);
nor I_38254 (I652843,I652778,I652507);
nor I_38255 (I652334,I652651,I652843);
not I_38256 (I652901,I2514);
DFFARX1 I_38257 (I159198,I2507,I652901,I652927,);
nand I_38258 (I652935,I652927,I159213);
DFFARX1 I_38259 (I159210,I2507,I652901,I652961,);
DFFARX1 I_38260 (I652961,I2507,I652901,I652978,);
not I_38261 (I652893,I652978);
not I_38262 (I653000,I159189);
nor I_38263 (I653017,I159189,I159195);
not I_38264 (I653034,I159201);
nand I_38265 (I653051,I653000,I653034);
nor I_38266 (I653068,I159201,I159189);
and I_38267 (I652872,I653068,I652935);
not I_38268 (I653099,I159207);
nand I_38269 (I653116,I653099,I159189);
nor I_38270 (I653133,I159207,I159192);
not I_38271 (I653150,I653133);
nand I_38272 (I652875,I653017,I653150);
DFFARX1 I_38273 (I653133,I2507,I652901,I652890,);
nor I_38274 (I653195,I159192,I159201);
nor I_38275 (I653212,I653195,I159195);
and I_38276 (I653229,I653212,I653116);
DFFARX1 I_38277 (I653229,I2507,I652901,I652887,);
nor I_38278 (I652884,I653195,I653051);
or I_38279 (I652881,I653133,I653195);
nor I_38280 (I653288,I159192,I159204);
DFFARX1 I_38281 (I653288,I2507,I652901,I653314,);
not I_38282 (I653322,I653314);
nand I_38283 (I653339,I653322,I653000);
nor I_38284 (I653356,I653339,I159195);
DFFARX1 I_38285 (I653356,I2507,I652901,I652869,);
nor I_38286 (I653387,I653322,I653051);
nor I_38287 (I652878,I653195,I653387);
not I_38288 (I653445,I2514);
DFFARX1 I_38289 (I306804,I2507,I653445,I653471,);
nand I_38290 (I653479,I653471,I306792);
DFFARX1 I_38291 (I306798,I2507,I653445,I653505,);
DFFARX1 I_38292 (I653505,I2507,I653445,I653522,);
not I_38293 (I653437,I653522);
not I_38294 (I653544,I306783);
nor I_38295 (I653561,I306783,I306795);
not I_38296 (I653578,I306786);
nand I_38297 (I653595,I653544,I653578);
nor I_38298 (I653612,I306786,I306783);
and I_38299 (I653416,I653612,I653479);
not I_38300 (I653643,I306801);
nand I_38301 (I653660,I653643,I306783);
nor I_38302 (I653677,I306801,I306807);
not I_38303 (I653694,I653677);
nand I_38304 (I653419,I653561,I653694);
DFFARX1 I_38305 (I653677,I2507,I653445,I653434,);
nor I_38306 (I653739,I306789,I306786);
nor I_38307 (I653756,I653739,I306795);
and I_38308 (I653773,I653756,I653660);
DFFARX1 I_38309 (I653773,I2507,I653445,I653431,);
nor I_38310 (I653428,I653739,I653595);
or I_38311 (I653425,I653677,I653739);
nor I_38312 (I653832,I306789,I306786);
DFFARX1 I_38313 (I653832,I2507,I653445,I653858,);
not I_38314 (I653866,I653858);
nand I_38315 (I653883,I653866,I653544);
nor I_38316 (I653900,I653883,I306795);
DFFARX1 I_38317 (I653900,I2507,I653445,I653413,);
nor I_38318 (I653931,I653866,I653595);
nor I_38319 (I653422,I653739,I653931);
not I_38320 (I653989,I2514);
DFFARX1 I_38321 (I180621,I2507,I653989,I654015,);
nand I_38322 (I654023,I654015,I180624);
DFFARX1 I_38323 (I180618,I2507,I653989,I654049,);
DFFARX1 I_38324 (I654049,I2507,I653989,I654066,);
not I_38325 (I653981,I654066);
not I_38326 (I654088,I180627);
nor I_38327 (I654105,I180627,I180612);
not I_38328 (I654122,I180636);
nand I_38329 (I654139,I654088,I654122);
nor I_38330 (I654156,I180636,I180627);
and I_38331 (I653960,I654156,I654023);
not I_38332 (I654187,I180615);
nand I_38333 (I654204,I654187,I180633);
nor I_38334 (I654221,I180615,I180609);
not I_38335 (I654238,I654221);
nand I_38336 (I653963,I654105,I654238);
DFFARX1 I_38337 (I654221,I2507,I653989,I653978,);
nor I_38338 (I654283,I180630,I180636);
nor I_38339 (I654300,I654283,I180612);
and I_38340 (I654317,I654300,I654204);
DFFARX1 I_38341 (I654317,I2507,I653989,I653975,);
nor I_38342 (I653972,I654283,I654139);
or I_38343 (I653969,I654221,I654283);
nor I_38344 (I654376,I180630,I180609);
DFFARX1 I_38345 (I654376,I2507,I653989,I654402,);
not I_38346 (I654410,I654402);
nand I_38347 (I654427,I654410,I654088);
nor I_38348 (I654444,I654427,I180612);
DFFARX1 I_38349 (I654444,I2507,I653989,I653957,);
nor I_38350 (I654475,I654410,I654139);
nor I_38351 (I653966,I654283,I654475);
not I_38352 (I654533,I2514);
DFFARX1 I_38353 (I28825,I2507,I654533,I654559,);
nand I_38354 (I654567,I654559,I28819);
DFFARX1 I_38355 (I28840,I2507,I654533,I654593,);
DFFARX1 I_38356 (I654593,I2507,I654533,I654610,);
not I_38357 (I654525,I654610);
not I_38358 (I654632,I28828);
nor I_38359 (I654649,I28828,I28837);
not I_38360 (I654666,I28816);
nand I_38361 (I654683,I654632,I654666);
nor I_38362 (I654700,I28816,I28828);
and I_38363 (I654504,I654700,I654567);
not I_38364 (I654731,I28834);
nand I_38365 (I654748,I654731,I28822);
nor I_38366 (I654765,I28834,I28816);
not I_38367 (I654782,I654765);
nand I_38368 (I654507,I654649,I654782);
DFFARX1 I_38369 (I654765,I2507,I654533,I654522,);
nor I_38370 (I654827,I28819,I28816);
nor I_38371 (I654844,I654827,I28837);
and I_38372 (I654861,I654844,I654748);
DFFARX1 I_38373 (I654861,I2507,I654533,I654519,);
nor I_38374 (I654516,I654827,I654683);
or I_38375 (I654513,I654765,I654827);
nor I_38376 (I654920,I28819,I28831);
DFFARX1 I_38377 (I654920,I2507,I654533,I654946,);
not I_38378 (I654954,I654946);
nand I_38379 (I654971,I654954,I654632);
nor I_38380 (I654988,I654971,I28837);
DFFARX1 I_38381 (I654988,I2507,I654533,I654501,);
nor I_38382 (I655019,I654954,I654683);
nor I_38383 (I654510,I654827,I655019);
not I_38384 (I655077,I2514);
DFFARX1 I_38385 (I533206,I2507,I655077,I655103,);
nand I_38386 (I655111,I655103,I533206);
DFFARX1 I_38387 (I533218,I2507,I655077,I655137,);
DFFARX1 I_38388 (I655137,I2507,I655077,I655154,);
not I_38389 (I655069,I655154);
not I_38390 (I655176,I533212);
nor I_38391 (I655193,I533212,I533233);
not I_38392 (I655210,I533221);
nand I_38393 (I655227,I655176,I655210);
nor I_38394 (I655244,I533221,I533212);
and I_38395 (I655048,I655244,I655111);
not I_38396 (I655275,I533215);
nand I_38397 (I655292,I655275,I533230);
nor I_38398 (I655309,I533215,I533224);
not I_38399 (I655326,I655309);
nand I_38400 (I655051,I655193,I655326);
DFFARX1 I_38401 (I655309,I2507,I655077,I655066,);
nor I_38402 (I655371,I533227,I533221);
nor I_38403 (I655388,I655371,I533233);
and I_38404 (I655405,I655388,I655292);
DFFARX1 I_38405 (I655405,I2507,I655077,I655063,);
nor I_38406 (I655060,I655371,I655227);
or I_38407 (I655057,I655309,I655371);
nor I_38408 (I655464,I533227,I533209);
DFFARX1 I_38409 (I655464,I2507,I655077,I655490,);
not I_38410 (I655498,I655490);
nand I_38411 (I655515,I655498,I655176);
nor I_38412 (I655532,I655515,I533233);
DFFARX1 I_38413 (I655532,I2507,I655077,I655045,);
nor I_38414 (I655563,I655498,I655227);
nor I_38415 (I655054,I655371,I655563);
not I_38416 (I655621,I2514);
DFFARX1 I_38417 (I286723,I2507,I655621,I655647,);
nand I_38418 (I655655,I655647,I286747);
DFFARX1 I_38419 (I286726,I2507,I655621,I655681,);
DFFARX1 I_38420 (I655681,I2507,I655621,I655698,);
not I_38421 (I655613,I655698);
not I_38422 (I655720,I286729);
nor I_38423 (I655737,I286729,I286744);
not I_38424 (I655754,I286735);
nand I_38425 (I655771,I655720,I655754);
nor I_38426 (I655788,I286735,I286729);
and I_38427 (I655592,I655788,I655655);
not I_38428 (I655819,I286732);
nand I_38429 (I655836,I655819,I286726);
nor I_38430 (I655853,I286732,I286741);
not I_38431 (I655870,I655853);
nand I_38432 (I655595,I655737,I655870);
DFFARX1 I_38433 (I655853,I2507,I655621,I655610,);
nor I_38434 (I655915,I286738,I286735);
nor I_38435 (I655932,I655915,I286744);
and I_38436 (I655949,I655932,I655836);
DFFARX1 I_38437 (I655949,I2507,I655621,I655607,);
nor I_38438 (I655604,I655915,I655771);
or I_38439 (I655601,I655853,I655915);
nor I_38440 (I656008,I286738,I286723);
DFFARX1 I_38441 (I656008,I2507,I655621,I656034,);
not I_38442 (I656042,I656034);
nand I_38443 (I656059,I656042,I655720);
nor I_38444 (I656076,I656059,I286744);
DFFARX1 I_38445 (I656076,I2507,I655621,I655589,);
nor I_38446 (I656107,I656042,I655771);
nor I_38447 (I655598,I655915,I656107);
not I_38448 (I656165,I2514);
DFFARX1 I_38449 (I551465,I2507,I656165,I656191,);
nand I_38450 (I656199,I656191,I551453);
DFFARX1 I_38451 (I551447,I2507,I656165,I656225,);
DFFARX1 I_38452 (I656225,I2507,I656165,I656242,);
not I_38453 (I656157,I656242);
not I_38454 (I656264,I551447);
nor I_38455 (I656281,I551447,I551459);
not I_38456 (I656298,I551456);
nand I_38457 (I656315,I656264,I656298);
nor I_38458 (I656332,I551456,I551447);
and I_38459 (I656136,I656332,I656199);
not I_38460 (I656363,I551450);
nand I_38461 (I656380,I656363,I551462);
nor I_38462 (I656397,I551450,I551468);
not I_38463 (I656414,I656397);
nand I_38464 (I656139,I656281,I656414);
DFFARX1 I_38465 (I656397,I2507,I656165,I656154,);
nor I_38466 (I656459,I551453,I551456);
nor I_38467 (I656476,I656459,I551459);
and I_38468 (I656493,I656476,I656380);
DFFARX1 I_38469 (I656493,I2507,I656165,I656151,);
nor I_38470 (I656148,I656459,I656315);
or I_38471 (I656145,I656397,I656459);
nor I_38472 (I656552,I551453,I551450);
DFFARX1 I_38473 (I656552,I2507,I656165,I656578,);
not I_38474 (I656586,I656578);
nand I_38475 (I656603,I656586,I656264);
nor I_38476 (I656620,I656603,I551459);
DFFARX1 I_38477 (I656620,I2507,I656165,I656133,);
nor I_38478 (I656651,I656586,I656315);
nor I_38479 (I656142,I656459,I656651);
not I_38480 (I656709,I2514);
DFFARX1 I_38481 (I508012,I2507,I656709,I656735,);
nand I_38482 (I656743,I656735,I508012);
DFFARX1 I_38483 (I508024,I2507,I656709,I656769,);
DFFARX1 I_38484 (I656769,I2507,I656709,I656786,);
not I_38485 (I656701,I656786);
not I_38486 (I656808,I508018);
nor I_38487 (I656825,I508018,I508039);
not I_38488 (I656842,I508027);
nand I_38489 (I656859,I656808,I656842);
nor I_38490 (I656876,I508027,I508018);
and I_38491 (I656680,I656876,I656743);
not I_38492 (I656907,I508021);
nand I_38493 (I656924,I656907,I508036);
nor I_38494 (I656941,I508021,I508030);
not I_38495 (I656958,I656941);
nand I_38496 (I656683,I656825,I656958);
DFFARX1 I_38497 (I656941,I2507,I656709,I656698,);
nor I_38498 (I657003,I508033,I508027);
nor I_38499 (I657020,I657003,I508039);
and I_38500 (I657037,I657020,I656924);
DFFARX1 I_38501 (I657037,I2507,I656709,I656695,);
nor I_38502 (I656692,I657003,I656859);
or I_38503 (I656689,I656941,I657003);
nor I_38504 (I657096,I508033,I508015);
DFFARX1 I_38505 (I657096,I2507,I656709,I657122,);
not I_38506 (I657130,I657122);
nand I_38507 (I657147,I657130,I656808);
nor I_38508 (I657164,I657147,I508039);
DFFARX1 I_38509 (I657164,I2507,I656709,I656677,);
nor I_38510 (I657195,I657130,I656859);
nor I_38511 (I656686,I657003,I657195);
not I_38512 (I657253,I2514);
DFFARX1 I_38513 (I14596,I2507,I657253,I657279,);
nand I_38514 (I657287,I657279,I14590);
DFFARX1 I_38515 (I14611,I2507,I657253,I657313,);
DFFARX1 I_38516 (I657313,I2507,I657253,I657330,);
not I_38517 (I657245,I657330);
not I_38518 (I657352,I14599);
nor I_38519 (I657369,I14599,I14608);
not I_38520 (I657386,I14587);
nand I_38521 (I657403,I657352,I657386);
nor I_38522 (I657420,I14587,I14599);
and I_38523 (I657224,I657420,I657287);
not I_38524 (I657451,I14605);
nand I_38525 (I657468,I657451,I14593);
nor I_38526 (I657485,I14605,I14587);
not I_38527 (I657502,I657485);
nand I_38528 (I657227,I657369,I657502);
DFFARX1 I_38529 (I657485,I2507,I657253,I657242,);
nor I_38530 (I657547,I14590,I14587);
nor I_38531 (I657564,I657547,I14608);
and I_38532 (I657581,I657564,I657468);
DFFARX1 I_38533 (I657581,I2507,I657253,I657239,);
nor I_38534 (I657236,I657547,I657403);
or I_38535 (I657233,I657485,I657547);
nor I_38536 (I657640,I14590,I14602);
DFFARX1 I_38537 (I657640,I2507,I657253,I657666,);
not I_38538 (I657674,I657666);
nand I_38539 (I657691,I657674,I657352);
nor I_38540 (I657708,I657691,I14608);
DFFARX1 I_38541 (I657708,I2507,I657253,I657221,);
nor I_38542 (I657739,I657674,I657403);
nor I_38543 (I657230,I657547,I657739);
not I_38544 (I657797,I2514);
DFFARX1 I_38545 (I121118,I2507,I657797,I657823,);
nand I_38546 (I657831,I657823,I121133);
DFFARX1 I_38547 (I121130,I2507,I657797,I657857,);
DFFARX1 I_38548 (I657857,I2507,I657797,I657874,);
not I_38549 (I657789,I657874);
not I_38550 (I657896,I121109);
nor I_38551 (I657913,I121109,I121115);
not I_38552 (I657930,I121121);
nand I_38553 (I657947,I657896,I657930);
nor I_38554 (I657964,I121121,I121109);
and I_38555 (I657768,I657964,I657831);
not I_38556 (I657995,I121127);
nand I_38557 (I658012,I657995,I121109);
nor I_38558 (I658029,I121127,I121112);
not I_38559 (I658046,I658029);
nand I_38560 (I657771,I657913,I658046);
DFFARX1 I_38561 (I658029,I2507,I657797,I657786,);
nor I_38562 (I658091,I121112,I121121);
nor I_38563 (I658108,I658091,I121115);
and I_38564 (I658125,I658108,I658012);
DFFARX1 I_38565 (I658125,I2507,I657797,I657783,);
nor I_38566 (I657780,I658091,I657947);
or I_38567 (I657777,I658029,I658091);
nor I_38568 (I658184,I121112,I121124);
DFFARX1 I_38569 (I658184,I2507,I657797,I658210,);
not I_38570 (I658218,I658210);
nand I_38571 (I658235,I658218,I657896);
nor I_38572 (I658252,I658235,I121115);
DFFARX1 I_38573 (I658252,I2507,I657797,I657765,);
nor I_38574 (I658283,I658218,I657947);
nor I_38575 (I657774,I658091,I658283);
not I_38576 (I658341,I2514);
DFFARX1 I_38577 (I561563,I2507,I658341,I658367,);
nand I_38578 (I658375,I658367,I561551);
DFFARX1 I_38579 (I561545,I2507,I658341,I658401,);
DFFARX1 I_38580 (I658401,I2507,I658341,I658418,);
not I_38581 (I658333,I658418);
not I_38582 (I658440,I561545);
nor I_38583 (I658457,I561545,I561557);
not I_38584 (I658474,I561554);
nand I_38585 (I658491,I658440,I658474);
nor I_38586 (I658508,I561554,I561545);
and I_38587 (I658312,I658508,I658375);
not I_38588 (I658539,I561548);
nand I_38589 (I658556,I658539,I561560);
nor I_38590 (I658573,I561548,I561566);
not I_38591 (I658590,I658573);
nand I_38592 (I658315,I658457,I658590);
DFFARX1 I_38593 (I658573,I2507,I658341,I658330,);
nor I_38594 (I658635,I561551,I561554);
nor I_38595 (I658652,I658635,I561557);
and I_38596 (I658669,I658652,I658556);
DFFARX1 I_38597 (I658669,I2507,I658341,I658327,);
nor I_38598 (I658324,I658635,I658491);
or I_38599 (I658321,I658573,I658635);
nor I_38600 (I658728,I561551,I561548);
DFFARX1 I_38601 (I658728,I2507,I658341,I658754,);
not I_38602 (I658762,I658754);
nand I_38603 (I658779,I658762,I658440);
nor I_38604 (I658796,I658779,I561557);
DFFARX1 I_38605 (I658796,I2507,I658341,I658309,);
nor I_38606 (I658827,I658762,I658491);
nor I_38607 (I658318,I658635,I658827);
not I_38608 (I658885,I2514);
DFFARX1 I_38609 (I424698,I2507,I658885,I658911,);
nand I_38610 (I658919,I658911,I424713);
DFFARX1 I_38611 (I424707,I2507,I658885,I658945,);
DFFARX1 I_38612 (I658945,I2507,I658885,I658962,);
not I_38613 (I658877,I658962);
not I_38614 (I658984,I424710);
nor I_38615 (I659001,I424710,I424716);
not I_38616 (I659018,I424698);
nand I_38617 (I659035,I658984,I659018);
nor I_38618 (I659052,I424698,I424710);
and I_38619 (I658856,I659052,I658919);
not I_38620 (I659083,I424695);
nand I_38621 (I659100,I659083,I424701);
nor I_38622 (I659117,I424695,I424695);
not I_38623 (I659134,I659117);
nand I_38624 (I658859,I659001,I659134);
DFFARX1 I_38625 (I659117,I2507,I658885,I658874,);
nor I_38626 (I659179,I424704,I424698);
nor I_38627 (I659196,I659179,I424716);
and I_38628 (I659213,I659196,I659100);
DFFARX1 I_38629 (I659213,I2507,I658885,I658871,);
nor I_38630 (I658868,I659179,I659035);
or I_38631 (I658865,I659117,I659179);
nor I_38632 (I659272,I424704,I424719);
DFFARX1 I_38633 (I659272,I2507,I658885,I659298,);
not I_38634 (I659306,I659298);
nand I_38635 (I659323,I659306,I658984);
nor I_38636 (I659340,I659323,I424716);
DFFARX1 I_38637 (I659340,I2507,I658885,I658853,);
nor I_38638 (I659371,I659306,I659035);
nor I_38639 (I658862,I659179,I659371);
not I_38640 (I659429,I2514);
DFFARX1 I_38641 (I498322,I2507,I659429,I659455,);
nand I_38642 (I659463,I659455,I498322);
DFFARX1 I_38643 (I498334,I2507,I659429,I659489,);
DFFARX1 I_38644 (I659489,I2507,I659429,I659506,);
not I_38645 (I659421,I659506);
not I_38646 (I659528,I498328);
nor I_38647 (I659545,I498328,I498349);
not I_38648 (I659562,I498337);
nand I_38649 (I659579,I659528,I659562);
nor I_38650 (I659596,I498337,I498328);
and I_38651 (I659400,I659596,I659463);
not I_38652 (I659627,I498331);
nand I_38653 (I659644,I659627,I498346);
nor I_38654 (I659661,I498331,I498340);
not I_38655 (I659678,I659661);
nand I_38656 (I659403,I659545,I659678);
DFFARX1 I_38657 (I659661,I2507,I659429,I659418,);
nor I_38658 (I659723,I498343,I498337);
nor I_38659 (I659740,I659723,I498349);
and I_38660 (I659757,I659740,I659644);
DFFARX1 I_38661 (I659757,I2507,I659429,I659415,);
nor I_38662 (I659412,I659723,I659579);
or I_38663 (I659409,I659661,I659723);
nor I_38664 (I659816,I498343,I498325);
DFFARX1 I_38665 (I659816,I2507,I659429,I659842,);
not I_38666 (I659850,I659842);
nand I_38667 (I659867,I659850,I659528);
nor I_38668 (I659884,I659867,I498349);
DFFARX1 I_38669 (I659884,I2507,I659429,I659397,);
nor I_38670 (I659915,I659850,I659579);
nor I_38671 (I659406,I659723,I659915);
not I_38672 (I659973,I2514);
DFFARX1 I_38673 (I537082,I2507,I659973,I659999,);
nand I_38674 (I660007,I659999,I537082);
DFFARX1 I_38675 (I537094,I2507,I659973,I660033,);
DFFARX1 I_38676 (I660033,I2507,I659973,I660050,);
not I_38677 (I659965,I660050);
not I_38678 (I660072,I537088);
nor I_38679 (I660089,I537088,I537109);
not I_38680 (I660106,I537097);
nand I_38681 (I660123,I660072,I660106);
nor I_38682 (I660140,I537097,I537088);
and I_38683 (I659944,I660140,I660007);
not I_38684 (I660171,I537091);
nand I_38685 (I660188,I660171,I537106);
nor I_38686 (I660205,I537091,I537100);
not I_38687 (I660222,I660205);
nand I_38688 (I659947,I660089,I660222);
DFFARX1 I_38689 (I660205,I2507,I659973,I659962,);
nor I_38690 (I660267,I537103,I537097);
nor I_38691 (I660284,I660267,I537109);
and I_38692 (I660301,I660284,I660188);
DFFARX1 I_38693 (I660301,I2507,I659973,I659959,);
nor I_38694 (I659956,I660267,I660123);
or I_38695 (I659953,I660205,I660267);
nor I_38696 (I660360,I537103,I537085);
DFFARX1 I_38697 (I660360,I2507,I659973,I660386,);
not I_38698 (I660394,I660386);
nand I_38699 (I660411,I660394,I660072);
nor I_38700 (I660428,I660411,I537109);
DFFARX1 I_38701 (I660428,I2507,I659973,I659941,);
nor I_38702 (I660459,I660394,I660123);
nor I_38703 (I659950,I660267,I660459);
not I_38704 (I660517,I2514);
DFFARX1 I_38705 (I254192,I2507,I660517,I660543,);
nand I_38706 (I660551,I660543,I254189);
DFFARX1 I_38707 (I254168,I2507,I660517,I660577,);
DFFARX1 I_38708 (I660577,I2507,I660517,I660594,);
not I_38709 (I660509,I660594);
not I_38710 (I660616,I254183);
nor I_38711 (I660633,I254183,I254186);
not I_38712 (I660650,I254177);
nand I_38713 (I660667,I660616,I660650);
nor I_38714 (I660684,I254177,I254183);
and I_38715 (I660488,I660684,I660551);
not I_38716 (I660715,I254174);
nand I_38717 (I660732,I660715,I254195);
nor I_38718 (I660749,I254174,I254171);
not I_38719 (I660766,I660749);
nand I_38720 (I660491,I660633,I660766);
DFFARX1 I_38721 (I660749,I2507,I660517,I660506,);
nor I_38722 (I660811,I254180,I254177);
nor I_38723 (I660828,I660811,I254186);
and I_38724 (I660845,I660828,I660732);
DFFARX1 I_38725 (I660845,I2507,I660517,I660503,);
nor I_38726 (I660500,I660811,I660667);
or I_38727 (I660497,I660749,I660811);
nor I_38728 (I660904,I254180,I254168);
DFFARX1 I_38729 (I660904,I2507,I660517,I660930,);
not I_38730 (I660938,I660930);
nand I_38731 (I660955,I660938,I660616);
nor I_38732 (I660972,I660955,I254186);
DFFARX1 I_38733 (I660972,I2507,I660517,I660485,);
nor I_38734 (I661003,I660938,I660667);
nor I_38735 (I660494,I660811,I661003);
not I_38736 (I661061,I2514);
DFFARX1 I_38737 (I611005,I2507,I661061,I661087,);
nand I_38738 (I661095,I661087,I610984);
DFFARX1 I_38739 (I610981,I2507,I661061,I661121,);
DFFARX1 I_38740 (I661121,I2507,I661061,I661138,);
not I_38741 (I661053,I661138);
not I_38742 (I661160,I610993);
nor I_38743 (I661177,I610993,I611002);
not I_38744 (I661194,I610990);
nand I_38745 (I661211,I661160,I661194);
nor I_38746 (I661228,I610990,I610993);
and I_38747 (I661032,I661228,I661095);
not I_38748 (I661259,I610999);
nand I_38749 (I661276,I661259,I610996);
nor I_38750 (I661293,I610999,I610981);
not I_38751 (I661310,I661293);
nand I_38752 (I661035,I661177,I661310);
DFFARX1 I_38753 (I661293,I2507,I661061,I661050,);
nor I_38754 (I661355,I610984,I610990);
nor I_38755 (I661372,I661355,I611002);
and I_38756 (I661389,I661372,I661276);
DFFARX1 I_38757 (I661389,I2507,I661061,I661047,);
nor I_38758 (I661044,I661355,I661211);
or I_38759 (I661041,I661293,I661355);
nor I_38760 (I661448,I610984,I610987);
DFFARX1 I_38761 (I661448,I2507,I661061,I661474,);
not I_38762 (I661482,I661474);
nand I_38763 (I661499,I661482,I661160);
nor I_38764 (I661516,I661499,I611002);
DFFARX1 I_38765 (I661516,I2507,I661061,I661029,);
nor I_38766 (I661547,I661482,I661211);
nor I_38767 (I661038,I661355,I661547);
not I_38768 (I661605,I2514);
DFFARX1 I_38769 (I731130,I2507,I661605,I661631,);
nand I_38770 (I661639,I661631,I731115);
DFFARX1 I_38771 (I731109,I2507,I661605,I661665,);
DFFARX1 I_38772 (I661665,I2507,I661605,I661682,);
not I_38773 (I661597,I661682);
not I_38774 (I661704,I731103);
nor I_38775 (I661721,I731103,I731124);
not I_38776 (I661738,I731112);
nand I_38777 (I661755,I661704,I661738);
nor I_38778 (I661772,I731112,I731103);
and I_38779 (I661576,I661772,I661639);
not I_38780 (I661803,I731121);
nand I_38781 (I661820,I661803,I731127);
nor I_38782 (I661837,I731121,I731118);
not I_38783 (I661854,I661837);
nand I_38784 (I661579,I661721,I661854);
DFFARX1 I_38785 (I661837,I2507,I661605,I661594,);
nor I_38786 (I661899,I731106,I731112);
nor I_38787 (I661916,I661899,I731124);
and I_38788 (I661933,I661916,I661820);
DFFARX1 I_38789 (I661933,I2507,I661605,I661591,);
nor I_38790 (I661588,I661899,I661755);
or I_38791 (I661585,I661837,I661899);
nor I_38792 (I661992,I731106,I731103);
DFFARX1 I_38793 (I661992,I2507,I661605,I662018,);
not I_38794 (I662026,I662018);
nand I_38795 (I662043,I662026,I661704);
nor I_38796 (I662060,I662043,I731124);
DFFARX1 I_38797 (I662060,I2507,I661605,I661573,);
nor I_38798 (I662091,I662026,I661755);
nor I_38799 (I661582,I661899,I662091);
not I_38800 (I662149,I2514);
DFFARX1 I_38801 (I723990,I2507,I662149,I662175,);
nand I_38802 (I662183,I662175,I723975);
DFFARX1 I_38803 (I723969,I2507,I662149,I662209,);
DFFARX1 I_38804 (I662209,I2507,I662149,I662226,);
not I_38805 (I662141,I662226);
not I_38806 (I662248,I723963);
nor I_38807 (I662265,I723963,I723984);
not I_38808 (I662282,I723972);
nand I_38809 (I662299,I662248,I662282);
nor I_38810 (I662316,I723972,I723963);
and I_38811 (I662120,I662316,I662183);
not I_38812 (I662347,I723981);
nand I_38813 (I662364,I662347,I723987);
nor I_38814 (I662381,I723981,I723978);
not I_38815 (I662398,I662381);
nand I_38816 (I662123,I662265,I662398);
DFFARX1 I_38817 (I662381,I2507,I662149,I662138,);
nor I_38818 (I662443,I723966,I723972);
nor I_38819 (I662460,I662443,I723984);
and I_38820 (I662477,I662460,I662364);
DFFARX1 I_38821 (I662477,I2507,I662149,I662135,);
nor I_38822 (I662132,I662443,I662299);
or I_38823 (I662129,I662381,I662443);
nor I_38824 (I662536,I723966,I723963);
DFFARX1 I_38825 (I662536,I2507,I662149,I662562,);
not I_38826 (I662570,I662562);
nand I_38827 (I662587,I662570,I662248);
nor I_38828 (I662604,I662587,I723984);
DFFARX1 I_38829 (I662604,I2507,I662149,I662117,);
nor I_38830 (I662635,I662570,I662299);
nor I_38831 (I662126,I662443,I662635);
not I_38832 (I662693,I2514);
DFFARX1 I_38833 (I241136,I2507,I662693,I662719,);
nand I_38834 (I662727,I662719,I241133);
DFFARX1 I_38835 (I241112,I2507,I662693,I662753,);
DFFARX1 I_38836 (I662753,I2507,I662693,I662770,);
not I_38837 (I662685,I662770);
not I_38838 (I662792,I241127);
nor I_38839 (I662809,I241127,I241130);
not I_38840 (I662826,I241121);
nand I_38841 (I662843,I662792,I662826);
nor I_38842 (I662860,I241121,I241127);
and I_38843 (I662664,I662860,I662727);
not I_38844 (I662891,I241118);
nand I_38845 (I662908,I662891,I241139);
nor I_38846 (I662925,I241118,I241115);
not I_38847 (I662942,I662925);
nand I_38848 (I662667,I662809,I662942);
DFFARX1 I_38849 (I662925,I2507,I662693,I662682,);
nor I_38850 (I662987,I241124,I241121);
nor I_38851 (I663004,I662987,I241130);
and I_38852 (I663021,I663004,I662908);
DFFARX1 I_38853 (I663021,I2507,I662693,I662679,);
nor I_38854 (I662676,I662987,I662843);
or I_38855 (I662673,I662925,I662987);
nor I_38856 (I663080,I241124,I241112);
DFFARX1 I_38857 (I663080,I2507,I662693,I663106,);
not I_38858 (I663114,I663106);
nand I_38859 (I663131,I663114,I662792);
nor I_38860 (I663148,I663131,I241130);
DFFARX1 I_38861 (I663148,I2507,I662693,I662661,);
nor I_38862 (I663179,I663114,I662843);
nor I_38863 (I662670,I662987,I663179);
not I_38864 (I663237,I2514);
DFFARX1 I_38865 (I413138,I2507,I663237,I663263,);
nand I_38866 (I663271,I663263,I413153);
DFFARX1 I_38867 (I413147,I2507,I663237,I663297,);
DFFARX1 I_38868 (I663297,I2507,I663237,I663314,);
not I_38869 (I663229,I663314);
not I_38870 (I663336,I413150);
nor I_38871 (I663353,I413150,I413156);
not I_38872 (I663370,I413138);
nand I_38873 (I663387,I663336,I663370);
nor I_38874 (I663404,I413138,I413150);
and I_38875 (I663208,I663404,I663271);
not I_38876 (I663435,I413135);
nand I_38877 (I663452,I663435,I413141);
nor I_38878 (I663469,I413135,I413135);
not I_38879 (I663486,I663469);
nand I_38880 (I663211,I663353,I663486);
DFFARX1 I_38881 (I663469,I2507,I663237,I663226,);
nor I_38882 (I663531,I413144,I413138);
nor I_38883 (I663548,I663531,I413156);
and I_38884 (I663565,I663548,I663452);
DFFARX1 I_38885 (I663565,I2507,I663237,I663223,);
nor I_38886 (I663220,I663531,I663387);
or I_38887 (I663217,I663469,I663531);
nor I_38888 (I663624,I413144,I413159);
DFFARX1 I_38889 (I663624,I2507,I663237,I663650,);
not I_38890 (I663658,I663650);
nand I_38891 (I663675,I663658,I663336);
nor I_38892 (I663692,I663675,I413156);
DFFARX1 I_38893 (I663692,I2507,I663237,I663205,);
nor I_38894 (I663723,I663658,I663387);
nor I_38895 (I663214,I663531,I663723);
not I_38896 (I663781,I2514);
DFFARX1 I_38897 (I10907,I2507,I663781,I663807,);
nand I_38898 (I663815,I663807,I10901);
DFFARX1 I_38899 (I10922,I2507,I663781,I663841,);
DFFARX1 I_38900 (I663841,I2507,I663781,I663858,);
not I_38901 (I663773,I663858);
not I_38902 (I663880,I10910);
nor I_38903 (I663897,I10910,I10919);
not I_38904 (I663914,I10898);
nand I_38905 (I663931,I663880,I663914);
nor I_38906 (I663948,I10898,I10910);
and I_38907 (I663752,I663948,I663815);
not I_38908 (I663979,I10916);
nand I_38909 (I663996,I663979,I10904);
nor I_38910 (I664013,I10916,I10898);
not I_38911 (I664030,I664013);
nand I_38912 (I663755,I663897,I664030);
DFFARX1 I_38913 (I664013,I2507,I663781,I663770,);
nor I_38914 (I664075,I10901,I10898);
nor I_38915 (I664092,I664075,I10919);
and I_38916 (I664109,I664092,I663996);
DFFARX1 I_38917 (I664109,I2507,I663781,I663767,);
nor I_38918 (I663764,I664075,I663931);
or I_38919 (I663761,I664013,I664075);
nor I_38920 (I664168,I10901,I10913);
DFFARX1 I_38921 (I664168,I2507,I663781,I664194,);
not I_38922 (I664202,I664194);
nand I_38923 (I664219,I664202,I663880);
nor I_38924 (I664236,I664219,I10919);
DFFARX1 I_38925 (I664236,I2507,I663781,I663749,);
nor I_38926 (I664267,I664202,I663931);
nor I_38927 (I663758,I664075,I664267);
not I_38928 (I664325,I2514);
DFFARX1 I_38929 (I550343,I2507,I664325,I664351,);
nand I_38930 (I664359,I664351,I550331);
DFFARX1 I_38931 (I550325,I2507,I664325,I664385,);
DFFARX1 I_38932 (I664385,I2507,I664325,I664402,);
not I_38933 (I664317,I664402);
not I_38934 (I664424,I550325);
nor I_38935 (I664441,I550325,I550337);
not I_38936 (I664458,I550334);
nand I_38937 (I664475,I664424,I664458);
nor I_38938 (I664492,I550334,I550325);
and I_38939 (I664296,I664492,I664359);
not I_38940 (I664523,I550328);
nand I_38941 (I664540,I664523,I550340);
nor I_38942 (I664557,I550328,I550346);
not I_38943 (I664574,I664557);
nand I_38944 (I664299,I664441,I664574);
DFFARX1 I_38945 (I664557,I2507,I664325,I664314,);
nor I_38946 (I664619,I550331,I550334);
nor I_38947 (I664636,I664619,I550337);
and I_38948 (I664653,I664636,I664540);
DFFARX1 I_38949 (I664653,I2507,I664325,I664311,);
nor I_38950 (I664308,I664619,I664475);
or I_38951 (I664305,I664557,I664619);
nor I_38952 (I664712,I550331,I550328);
DFFARX1 I_38953 (I664712,I2507,I664325,I664738,);
not I_38954 (I664746,I664738);
nand I_38955 (I664763,I664746,I664424);
nor I_38956 (I664780,I664763,I550337);
DFFARX1 I_38957 (I664780,I2507,I664325,I664293,);
nor I_38958 (I664811,I664746,I664475);
nor I_38959 (I664302,I664619,I664811);
not I_38960 (I664869,I2514);
DFFARX1 I_38961 (I105648,I2507,I664869,I664895,);
nand I_38962 (I664903,I664895,I105663);
DFFARX1 I_38963 (I105660,I2507,I664869,I664929,);
DFFARX1 I_38964 (I664929,I2507,I664869,I664946,);
not I_38965 (I664861,I664946);
not I_38966 (I664968,I105639);
nor I_38967 (I664985,I105639,I105645);
not I_38968 (I665002,I105651);
nand I_38969 (I665019,I664968,I665002);
nor I_38970 (I665036,I105651,I105639);
and I_38971 (I664840,I665036,I664903);
not I_38972 (I665067,I105657);
nand I_38973 (I665084,I665067,I105639);
nor I_38974 (I665101,I105657,I105642);
not I_38975 (I665118,I665101);
nand I_38976 (I664843,I664985,I665118);
DFFARX1 I_38977 (I665101,I2507,I664869,I664858,);
nor I_38978 (I665163,I105642,I105651);
nor I_38979 (I665180,I665163,I105645);
and I_38980 (I665197,I665180,I665084);
DFFARX1 I_38981 (I665197,I2507,I664869,I664855,);
nor I_38982 (I664852,I665163,I665019);
or I_38983 (I664849,I665101,I665163);
nor I_38984 (I665256,I105642,I105654);
DFFARX1 I_38985 (I665256,I2507,I664869,I665282,);
not I_38986 (I665290,I665282);
nand I_38987 (I665307,I665290,I664968);
nor I_38988 (I665324,I665307,I105645);
DFFARX1 I_38989 (I665324,I2507,I664869,I664837,);
nor I_38990 (I665355,I665290,I665019);
nor I_38991 (I664846,I665163,I665355);
not I_38992 (I665413,I2514);
DFFARX1 I_38993 (I58349,I2507,I665413,I665439,);
nand I_38994 (I665447,I665439,I58331);
DFFARX1 I_38995 (I58328,I2507,I665413,I665473,);
DFFARX1 I_38996 (I665473,I2507,I665413,I665490,);
not I_38997 (I665405,I665490);
not I_38998 (I665512,I58346);
nor I_38999 (I665529,I58346,I58340);
not I_39000 (I665546,I58328);
nand I_39001 (I665563,I665512,I665546);
nor I_39002 (I665580,I58328,I58346);
and I_39003 (I665384,I665580,I665447);
not I_39004 (I665611,I58337);
nand I_39005 (I665628,I665611,I58343);
nor I_39006 (I665645,I58337,I58331);
not I_39007 (I665662,I665645);
nand I_39008 (I665387,I665529,I665662);
DFFARX1 I_39009 (I665645,I2507,I665413,I665402,);
nor I_39010 (I665707,I58334,I58328);
nor I_39011 (I665724,I665707,I58340);
and I_39012 (I665741,I665724,I665628);
DFFARX1 I_39013 (I665741,I2507,I665413,I665399,);
nor I_39014 (I665396,I665707,I665563);
or I_39015 (I665393,I665645,I665707);
nor I_39016 (I665800,I58334,I58352);
DFFARX1 I_39017 (I665800,I2507,I665413,I665826,);
not I_39018 (I665834,I665826);
nand I_39019 (I665851,I665834,I665512);
nor I_39020 (I665868,I665851,I58340);
DFFARX1 I_39021 (I665868,I2507,I665413,I665381,);
nor I_39022 (I665899,I665834,I665563);
nor I_39023 (I665390,I665707,I665899);
not I_39024 (I665957,I2514);
DFFARX1 I_39025 (I410823,I2507,I665957,I665983,);
nand I_39026 (I665991,I665983,I410826);
not I_39027 (I666008,I665991);
DFFARX1 I_39028 (I410838,I2507,I665957,I666034,);
not I_39029 (I666042,I666034);
not I_39030 (I666059,I410823);
or I_39031 (I666076,I410832,I410823);
nor I_39032 (I666093,I410832,I410823);
or I_39033 (I666110,I410841,I410832);
DFFARX1 I_39034 (I666110,I2507,I665957,I665949,);
not I_39035 (I666141,I410844);
nand I_39036 (I666158,I666141,I410826);
nand I_39037 (I666175,I666059,I666158);
and I_39038 (I665928,I666042,I666175);
nor I_39039 (I666206,I410844,I410829);
and I_39040 (I666223,I666042,I666206);
nor I_39041 (I665934,I666008,I666223);
DFFARX1 I_39042 (I666206,I2507,I665957,I666263,);
not I_39043 (I666271,I666263);
nor I_39044 (I665943,I666042,I666271);
or I_39045 (I666302,I666110,I410835);
nor I_39046 (I666319,I410835,I410841);
nand I_39047 (I666336,I666175,I666319);
nand I_39048 (I666353,I666302,I666336);
DFFARX1 I_39049 (I666353,I2507,I665957,I665946,);
nor I_39050 (I666384,I666319,I666076);
DFFARX1 I_39051 (I666384,I2507,I665957,I665925,);
nor I_39052 (I666415,I410835,I410847);
DFFARX1 I_39053 (I666415,I2507,I665957,I666441,);
DFFARX1 I_39054 (I666441,I2507,I665957,I665940,);
not I_39055 (I666463,I666441);
nand I_39056 (I665937,I666463,I665991);
nand I_39057 (I665931,I666463,I666093);
not I_39058 (I666535,I2514);
DFFARX1 I_39059 (I448141,I2507,I666535,I666561,);
nand I_39060 (I666569,I666561,I448141);
not I_39061 (I666586,I666569);
DFFARX1 I_39062 (I448147,I2507,I666535,I666612,);
not I_39063 (I666620,I666612);
not I_39064 (I666637,I448159);
or I_39065 (I666654,I448144,I448159);
nor I_39066 (I666671,I448144,I448159);
or I_39067 (I666688,I448138,I448144);
DFFARX1 I_39068 (I666688,I2507,I666535,I666527,);
not I_39069 (I666719,I448156);
nand I_39070 (I666736,I666719,I448150);
nand I_39071 (I666753,I666637,I666736);
and I_39072 (I666506,I666620,I666753);
nor I_39073 (I666784,I448156,I448138);
and I_39074 (I666801,I666620,I666784);
nor I_39075 (I666512,I666586,I666801);
DFFARX1 I_39076 (I666784,I2507,I666535,I666841,);
not I_39077 (I666849,I666841);
nor I_39078 (I666521,I666620,I666849);
or I_39079 (I666880,I666688,I448153);
nor I_39080 (I666897,I448153,I448138);
nand I_39081 (I666914,I666753,I666897);
nand I_39082 (I666931,I666880,I666914);
DFFARX1 I_39083 (I666931,I2507,I666535,I666524,);
nor I_39084 (I666962,I666897,I666654);
DFFARX1 I_39085 (I666962,I2507,I666535,I666503,);
nor I_39086 (I666993,I448153,I448144);
DFFARX1 I_39087 (I666993,I2507,I666535,I667019,);
DFFARX1 I_39088 (I667019,I2507,I666535,I666518,);
not I_39089 (I667041,I667019);
nand I_39090 (I666515,I667041,I666569);
nand I_39091 (I666509,I667041,I666671);
not I_39092 (I667113,I2514);
DFFARX1 I_39093 (I174818,I2507,I667113,I667139,);
nand I_39094 (I667147,I667139,I174839);
not I_39095 (I667164,I667147);
DFFARX1 I_39096 (I174833,I2507,I667113,I667190,);
not I_39097 (I667198,I667190);
not I_39098 (I667215,I174821);
or I_39099 (I667232,I174836,I174821);
nor I_39100 (I667249,I174836,I174821);
or I_39101 (I667266,I174827,I174836);
DFFARX1 I_39102 (I667266,I2507,I667113,I667105,);
not I_39103 (I667297,I174815);
nand I_39104 (I667314,I667297,I174812);
nand I_39105 (I667331,I667215,I667314);
and I_39106 (I667084,I667198,I667331);
nor I_39107 (I667362,I174815,I174824);
and I_39108 (I667379,I667198,I667362);
nor I_39109 (I667090,I667164,I667379);
DFFARX1 I_39110 (I667362,I2507,I667113,I667419,);
not I_39111 (I667427,I667419);
nor I_39112 (I667099,I667198,I667427);
or I_39113 (I667458,I667266,I174830);
nor I_39114 (I667475,I174830,I174827);
nand I_39115 (I667492,I667331,I667475);
nand I_39116 (I667509,I667458,I667492);
DFFARX1 I_39117 (I667509,I2507,I667113,I667102,);
nor I_39118 (I667540,I667475,I667232);
DFFARX1 I_39119 (I667540,I2507,I667113,I667081,);
nor I_39120 (I667571,I174830,I174812);
DFFARX1 I_39121 (I667571,I2507,I667113,I667597,);
DFFARX1 I_39122 (I667597,I2507,I667113,I667096,);
not I_39123 (I667619,I667597);
nand I_39124 (I667093,I667619,I667147);
nand I_39125 (I667087,I667619,I667249);
not I_39126 (I667691,I2514);
DFFARX1 I_39127 (I348977,I2507,I667691,I667717,);
nand I_39128 (I667725,I667717,I348980);
not I_39129 (I667742,I667725);
DFFARX1 I_39130 (I348992,I2507,I667691,I667768,);
not I_39131 (I667776,I667768);
not I_39132 (I667793,I348977);
or I_39133 (I667810,I348986,I348977);
nor I_39134 (I667827,I348986,I348977);
or I_39135 (I667844,I348995,I348986);
DFFARX1 I_39136 (I667844,I2507,I667691,I667683,);
not I_39137 (I667875,I348998);
nand I_39138 (I667892,I667875,I348980);
nand I_39139 (I667909,I667793,I667892);
and I_39140 (I667662,I667776,I667909);
nor I_39141 (I667940,I348998,I348983);
and I_39142 (I667957,I667776,I667940);
nor I_39143 (I667668,I667742,I667957);
DFFARX1 I_39144 (I667940,I2507,I667691,I667997,);
not I_39145 (I668005,I667997);
nor I_39146 (I667677,I667776,I668005);
or I_39147 (I668036,I667844,I348989);
nor I_39148 (I668053,I348989,I348995);
nand I_39149 (I668070,I667909,I668053);
nand I_39150 (I668087,I668036,I668070);
DFFARX1 I_39151 (I668087,I2507,I667691,I667680,);
nor I_39152 (I668118,I668053,I667810);
DFFARX1 I_39153 (I668118,I2507,I667691,I667659,);
nor I_39154 (I668149,I348989,I349001);
DFFARX1 I_39155 (I668149,I2507,I667691,I668175,);
DFFARX1 I_39156 (I668175,I2507,I667691,I667674,);
not I_39157 (I668197,I668175);
nand I_39158 (I667671,I668197,I667725);
nand I_39159 (I667665,I668197,I667827);
not I_39160 (I668269,I2514);
DFFARX1 I_39161 (I70461,I2507,I668269,I668295,);
nand I_39162 (I668303,I668295,I70452);
not I_39163 (I668320,I668303);
DFFARX1 I_39164 (I70449,I2507,I668269,I668346,);
not I_39165 (I668354,I668346);
not I_39166 (I668371,I70458);
or I_39167 (I668388,I70449,I70458);
nor I_39168 (I668405,I70449,I70458);
or I_39169 (I668422,I70455,I70449);
DFFARX1 I_39170 (I668422,I2507,I668269,I668261,);
not I_39171 (I668453,I70464);
nand I_39172 (I668470,I668453,I70473);
nand I_39173 (I668487,I668371,I668470);
and I_39174 (I668240,I668354,I668487);
nor I_39175 (I668518,I70464,I70467);
and I_39176 (I668535,I668354,I668518);
nor I_39177 (I668246,I668320,I668535);
DFFARX1 I_39178 (I668518,I2507,I668269,I668575,);
not I_39179 (I668583,I668575);
nor I_39180 (I668255,I668354,I668583);
or I_39181 (I668614,I668422,I70452);
nor I_39182 (I668631,I70452,I70455);
nand I_39183 (I668648,I668487,I668631);
nand I_39184 (I668665,I668614,I668648);
DFFARX1 I_39185 (I668665,I2507,I668269,I668258,);
nor I_39186 (I668696,I668631,I668388);
DFFARX1 I_39187 (I668696,I2507,I668269,I668237,);
nor I_39188 (I668727,I70452,I70470);
DFFARX1 I_39189 (I668727,I2507,I668269,I668753,);
DFFARX1 I_39190 (I668753,I2507,I668269,I668252,);
not I_39191 (I668775,I668753);
nand I_39192 (I668249,I668775,I668303);
nand I_39193 (I668243,I668775,I668405);
not I_39194 (I668847,I2514);
DFFARX1 I_39195 (I553700,I2507,I668847,I668873,);
nand I_39196 (I668881,I668873,I553697);
not I_39197 (I668898,I668881);
DFFARX1 I_39198 (I553697,I2507,I668847,I668924,);
not I_39199 (I668932,I668924);
not I_39200 (I668949,I553694);
or I_39201 (I668966,I553703,I553694);
nor I_39202 (I668983,I553703,I553694);
or I_39203 (I669000,I553706,I553703);
DFFARX1 I_39204 (I669000,I2507,I668847,I668839,);
not I_39205 (I669031,I553694);
nand I_39206 (I669048,I669031,I553691);
nand I_39207 (I669065,I668949,I669048);
and I_39208 (I668818,I668932,I669065);
nor I_39209 (I669096,I553694,I553709);
and I_39210 (I669113,I668932,I669096);
nor I_39211 (I668824,I668898,I669113);
DFFARX1 I_39212 (I669096,I2507,I668847,I669153,);
not I_39213 (I669161,I669153);
nor I_39214 (I668833,I668932,I669161);
or I_39215 (I669192,I669000,I553712);
nor I_39216 (I669209,I553712,I553706);
nand I_39217 (I669226,I669065,I669209);
nand I_39218 (I669243,I669192,I669226);
DFFARX1 I_39219 (I669243,I2507,I668847,I668836,);
nor I_39220 (I669274,I669209,I668966);
DFFARX1 I_39221 (I669274,I2507,I668847,I668815,);
nor I_39222 (I669305,I553712,I553691);
DFFARX1 I_39223 (I669305,I2507,I668847,I669331,);
DFFARX1 I_39224 (I669331,I2507,I668847,I668830,);
not I_39225 (I669353,I669331);
nand I_39226 (I668827,I669353,I668881);
nand I_39227 (I668821,I669353,I668983);
not I_39228 (I669425,I2514);
DFFARX1 I_39229 (I110399,I2507,I669425,I669451,);
nand I_39230 (I669459,I669451,I110402);
not I_39231 (I669476,I669459);
DFFARX1 I_39232 (I110411,I2507,I669425,I669502,);
not I_39233 (I669510,I669502);
not I_39234 (I669527,I110414);
or I_39235 (I669544,I110405,I110414);
nor I_39236 (I669561,I110405,I110414);
or I_39237 (I669578,I110417,I110405);
DFFARX1 I_39238 (I669578,I2507,I669425,I669417,);
not I_39239 (I669609,I110402);
nand I_39240 (I669626,I669609,I110408);
nand I_39241 (I669643,I669527,I669626);
and I_39242 (I669396,I669510,I669643);
nor I_39243 (I669674,I110402,I110420);
and I_39244 (I669691,I669510,I669674);
nor I_39245 (I669402,I669476,I669691);
DFFARX1 I_39246 (I669674,I2507,I669425,I669731,);
not I_39247 (I669739,I669731);
nor I_39248 (I669411,I669510,I669739);
or I_39249 (I669770,I669578,I110399);
nor I_39250 (I669787,I110399,I110417);
nand I_39251 (I669804,I669643,I669787);
nand I_39252 (I669821,I669770,I669804);
DFFARX1 I_39253 (I669821,I2507,I669425,I669414,);
nor I_39254 (I669852,I669787,I669544);
DFFARX1 I_39255 (I669852,I2507,I669425,I669393,);
nor I_39256 (I669883,I110399,I110423);
DFFARX1 I_39257 (I669883,I2507,I669425,I669909,);
DFFARX1 I_39258 (I669909,I2507,I669425,I669408,);
not I_39259 (I669931,I669909);
nand I_39260 (I669405,I669931,I669459);
nand I_39261 (I669399,I669931,I669561);
not I_39262 (I670003,I2514);
DFFARX1 I_39263 (I91954,I2507,I670003,I670029,);
nand I_39264 (I670037,I670029,I91957);
not I_39265 (I670054,I670037);
DFFARX1 I_39266 (I91966,I2507,I670003,I670080,);
not I_39267 (I670088,I670080);
not I_39268 (I670105,I91969);
or I_39269 (I670122,I91960,I91969);
nor I_39270 (I670139,I91960,I91969);
or I_39271 (I670156,I91972,I91960);
DFFARX1 I_39272 (I670156,I2507,I670003,I669995,);
not I_39273 (I670187,I91957);
nand I_39274 (I670204,I670187,I91963);
nand I_39275 (I670221,I670105,I670204);
and I_39276 (I669974,I670088,I670221);
nor I_39277 (I670252,I91957,I91975);
and I_39278 (I670269,I670088,I670252);
nor I_39279 (I669980,I670054,I670269);
DFFARX1 I_39280 (I670252,I2507,I670003,I670309,);
not I_39281 (I670317,I670309);
nor I_39282 (I669989,I670088,I670317);
or I_39283 (I670348,I670156,I91954);
nor I_39284 (I670365,I91954,I91972);
nand I_39285 (I670382,I670221,I670365);
nand I_39286 (I670399,I670348,I670382);
DFFARX1 I_39287 (I670399,I2507,I670003,I669992,);
nor I_39288 (I670430,I670365,I670122);
DFFARX1 I_39289 (I670430,I2507,I670003,I669971,);
nor I_39290 (I670461,I91954,I91978);
DFFARX1 I_39291 (I670461,I2507,I670003,I670487,);
DFFARX1 I_39292 (I670487,I2507,I670003,I669986,);
not I_39293 (I670509,I670487);
nand I_39294 (I669983,I670509,I670037);
nand I_39295 (I669977,I670509,I670139);
not I_39296 (I670581,I2514);
DFFARX1 I_39297 (I381923,I2507,I670581,I670607,);
nand I_39298 (I670615,I670607,I381926);
not I_39299 (I670632,I670615);
DFFARX1 I_39300 (I381938,I2507,I670581,I670658,);
not I_39301 (I670666,I670658);
not I_39302 (I670683,I381923);
or I_39303 (I670700,I381932,I381923);
nor I_39304 (I670717,I381932,I381923);
or I_39305 (I670734,I381941,I381932);
DFFARX1 I_39306 (I670734,I2507,I670581,I670573,);
not I_39307 (I670765,I381944);
nand I_39308 (I670782,I670765,I381926);
nand I_39309 (I670799,I670683,I670782);
and I_39310 (I670552,I670666,I670799);
nor I_39311 (I670830,I381944,I381929);
and I_39312 (I670847,I670666,I670830);
nor I_39313 (I670558,I670632,I670847);
DFFARX1 I_39314 (I670830,I2507,I670581,I670887,);
not I_39315 (I670895,I670887);
nor I_39316 (I670567,I670666,I670895);
or I_39317 (I670926,I670734,I381935);
nor I_39318 (I670943,I381935,I381941);
nand I_39319 (I670960,I670799,I670943);
nand I_39320 (I670977,I670926,I670960);
DFFARX1 I_39321 (I670977,I2507,I670581,I670570,);
nor I_39322 (I671008,I670943,I670700);
DFFARX1 I_39323 (I671008,I2507,I670581,I670549,);
nor I_39324 (I671039,I381935,I381947);
DFFARX1 I_39325 (I671039,I2507,I670581,I671065,);
DFFARX1 I_39326 (I671065,I2507,I670581,I670564,);
not I_39327 (I671087,I671065);
nand I_39328 (I670561,I671087,I670615);
nand I_39329 (I670555,I671087,I670717);
not I_39330 (I671159,I2514);
DFFARX1 I_39331 (I424117,I2507,I671159,I671185,);
nand I_39332 (I671193,I671185,I424120);
not I_39333 (I671210,I671193);
DFFARX1 I_39334 (I424132,I2507,I671159,I671236,);
not I_39335 (I671244,I671236);
not I_39336 (I671261,I424117);
or I_39337 (I671278,I424126,I424117);
nor I_39338 (I671295,I424126,I424117);
or I_39339 (I671312,I424135,I424126);
DFFARX1 I_39340 (I671312,I2507,I671159,I671151,);
not I_39341 (I671343,I424138);
nand I_39342 (I671360,I671343,I424120);
nand I_39343 (I671377,I671261,I671360);
and I_39344 (I671130,I671244,I671377);
nor I_39345 (I671408,I424138,I424123);
and I_39346 (I671425,I671244,I671408);
nor I_39347 (I671136,I671210,I671425);
DFFARX1 I_39348 (I671408,I2507,I671159,I671465,);
not I_39349 (I671473,I671465);
nor I_39350 (I671145,I671244,I671473);
or I_39351 (I671504,I671312,I424129);
nor I_39352 (I671521,I424129,I424135);
nand I_39353 (I671538,I671377,I671521);
nand I_39354 (I671555,I671504,I671538);
DFFARX1 I_39355 (I671555,I2507,I671159,I671148,);
nor I_39356 (I671586,I671521,I671278);
DFFARX1 I_39357 (I671586,I2507,I671159,I671127,);
nor I_39358 (I671617,I424129,I424141);
DFFARX1 I_39359 (I671617,I2507,I671159,I671643,);
DFFARX1 I_39360 (I671643,I2507,I671159,I671142,);
not I_39361 (I671665,I671643);
nand I_39362 (I671139,I671665,I671193);
nand I_39363 (I671133,I671665,I671295);
not I_39364 (I671737,I2514);
DFFARX1 I_39365 (I407933,I2507,I671737,I671763,);
nand I_39366 (I671771,I671763,I407936);
not I_39367 (I671788,I671771);
DFFARX1 I_39368 (I407948,I2507,I671737,I671814,);
not I_39369 (I671822,I671814);
not I_39370 (I671839,I407933);
or I_39371 (I671856,I407942,I407933);
nor I_39372 (I671873,I407942,I407933);
or I_39373 (I671890,I407951,I407942);
DFFARX1 I_39374 (I671890,I2507,I671737,I671729,);
not I_39375 (I671921,I407954);
nand I_39376 (I671938,I671921,I407936);
nand I_39377 (I671955,I671839,I671938);
and I_39378 (I671708,I671822,I671955);
nor I_39379 (I671986,I407954,I407939);
and I_39380 (I672003,I671822,I671986);
nor I_39381 (I671714,I671788,I672003);
DFFARX1 I_39382 (I671986,I2507,I671737,I672043,);
not I_39383 (I672051,I672043);
nor I_39384 (I671723,I671822,I672051);
or I_39385 (I672082,I671890,I407945);
nor I_39386 (I672099,I407945,I407951);
nand I_39387 (I672116,I671955,I672099);
nand I_39388 (I672133,I672082,I672116);
DFFARX1 I_39389 (I672133,I2507,I671737,I671726,);
nor I_39390 (I672164,I672099,I671856);
DFFARX1 I_39391 (I672164,I2507,I671737,I671705,);
nor I_39392 (I672195,I407945,I407957);
DFFARX1 I_39393 (I672195,I2507,I671737,I672221,);
DFFARX1 I_39394 (I672221,I2507,I671737,I671720,);
not I_39395 (I672243,I672221);
nand I_39396 (I671717,I672243,I671771);
nand I_39397 (I671711,I672243,I671873);
not I_39398 (I672315,I2514);
DFFARX1 I_39399 (I481532,I2507,I672315,I672341,);
nand I_39400 (I672349,I672341,I481553);
not I_39401 (I672366,I672349);
DFFARX1 I_39402 (I481526,I2507,I672315,I672392,);
not I_39403 (I672400,I672392);
not I_39404 (I672417,I481547);
or I_39405 (I672434,I481538,I481547);
nor I_39406 (I672451,I481538,I481547);
or I_39407 (I672468,I481541,I481538);
DFFARX1 I_39408 (I672468,I2507,I672315,I672307,);
not I_39409 (I672499,I481529);
nand I_39410 (I672516,I672499,I481544);
nand I_39411 (I672533,I672417,I672516);
and I_39412 (I672286,I672400,I672533);
nor I_39413 (I672564,I481529,I481526);
and I_39414 (I672581,I672400,I672564);
nor I_39415 (I672292,I672366,I672581);
DFFARX1 I_39416 (I672564,I2507,I672315,I672621,);
not I_39417 (I672629,I672621);
nor I_39418 (I672301,I672400,I672629);
or I_39419 (I672660,I672468,I481550);
nor I_39420 (I672677,I481550,I481541);
nand I_39421 (I672694,I672533,I672677);
nand I_39422 (I672711,I672660,I672694);
DFFARX1 I_39423 (I672711,I2507,I672315,I672304,);
nor I_39424 (I672742,I672677,I672434);
DFFARX1 I_39425 (I672742,I2507,I672315,I672283,);
nor I_39426 (I672773,I481550,I481535);
DFFARX1 I_39427 (I672773,I2507,I672315,I672799,);
DFFARX1 I_39428 (I672799,I2507,I672315,I672298,);
not I_39429 (I672821,I672799);
nand I_39430 (I672295,I672821,I672349);
nand I_39431 (I672289,I672821,I672451);
not I_39432 (I672893,I2514);
DFFARX1 I_39433 (I278107,I2507,I672893,I672919,);
nand I_39434 (I672927,I672919,I278116);
not I_39435 (I672944,I672927);
DFFARX1 I_39436 (I278104,I2507,I672893,I672970,);
not I_39437 (I672978,I672970);
not I_39438 (I672995,I278110);
or I_39439 (I673012,I278104,I278110);
nor I_39440 (I673029,I278104,I278110);
or I_39441 (I673046,I278119,I278104);
DFFARX1 I_39442 (I673046,I2507,I672893,I672885,);
not I_39443 (I673077,I278113);
nand I_39444 (I673094,I673077,I278128);
nand I_39445 (I673111,I672995,I673094);
and I_39446 (I672864,I672978,I673111);
nor I_39447 (I673142,I278113,I278131);
and I_39448 (I673159,I672978,I673142);
nor I_39449 (I672870,I672944,I673159);
DFFARX1 I_39450 (I673142,I2507,I672893,I673199,);
not I_39451 (I673207,I673199);
nor I_39452 (I672879,I672978,I673207);
or I_39453 (I673238,I673046,I278122);
nor I_39454 (I673255,I278122,I278119);
nand I_39455 (I673272,I673111,I673255);
nand I_39456 (I673289,I673238,I673272);
DFFARX1 I_39457 (I673289,I2507,I672893,I672882,);
nor I_39458 (I673320,I673255,I673012);
DFFARX1 I_39459 (I673320,I2507,I672893,I672861,);
nor I_39460 (I673351,I278122,I278125);
DFFARX1 I_39461 (I673351,I2507,I672893,I673377,);
DFFARX1 I_39462 (I673377,I2507,I672893,I672876,);
not I_39463 (I673399,I673377);
nand I_39464 (I672873,I673399,I672927);
nand I_39465 (I672867,I673399,I673029);
not I_39466 (I673471,I2514);
DFFARX1 I_39467 (I130034,I2507,I673471,I673497,);
nand I_39468 (I673505,I673497,I130037);
not I_39469 (I673522,I673505);
DFFARX1 I_39470 (I130046,I2507,I673471,I673548,);
not I_39471 (I673556,I673548);
not I_39472 (I673573,I130049);
or I_39473 (I673590,I130040,I130049);
nor I_39474 (I673607,I130040,I130049);
or I_39475 (I673624,I130052,I130040);
DFFARX1 I_39476 (I673624,I2507,I673471,I673463,);
not I_39477 (I673655,I130037);
nand I_39478 (I673672,I673655,I130043);
nand I_39479 (I673689,I673573,I673672);
and I_39480 (I673442,I673556,I673689);
nor I_39481 (I673720,I130037,I130055);
and I_39482 (I673737,I673556,I673720);
nor I_39483 (I673448,I673522,I673737);
DFFARX1 I_39484 (I673720,I2507,I673471,I673777,);
not I_39485 (I673785,I673777);
nor I_39486 (I673457,I673556,I673785);
or I_39487 (I673816,I673624,I130034);
nor I_39488 (I673833,I130034,I130052);
nand I_39489 (I673850,I673689,I673833);
nand I_39490 (I673867,I673816,I673850);
DFFARX1 I_39491 (I673867,I2507,I673471,I673460,);
nor I_39492 (I673898,I673833,I673590);
DFFARX1 I_39493 (I673898,I2507,I673471,I673439,);
nor I_39494 (I673929,I130034,I130058);
DFFARX1 I_39495 (I673929,I2507,I673471,I673955,);
DFFARX1 I_39496 (I673955,I2507,I673471,I673454,);
not I_39497 (I673977,I673955);
nand I_39498 (I673451,I673977,I673505);
nand I_39499 (I673445,I673977,I673607);
not I_39500 (I674049,I2514);
DFFARX1 I_39501 (I250907,I2507,I674049,I674075,);
nand I_39502 (I674083,I674075,I250916);
not I_39503 (I674100,I674083);
DFFARX1 I_39504 (I250904,I2507,I674049,I674126,);
not I_39505 (I674134,I674126);
not I_39506 (I674151,I250910);
or I_39507 (I674168,I250904,I250910);
nor I_39508 (I674185,I250904,I250910);
or I_39509 (I674202,I250919,I250904);
DFFARX1 I_39510 (I674202,I2507,I674049,I674041,);
not I_39511 (I674233,I250913);
nand I_39512 (I674250,I674233,I250928);
nand I_39513 (I674267,I674151,I674250);
and I_39514 (I674020,I674134,I674267);
nor I_39515 (I674298,I250913,I250931);
and I_39516 (I674315,I674134,I674298);
nor I_39517 (I674026,I674100,I674315);
DFFARX1 I_39518 (I674298,I2507,I674049,I674355,);
not I_39519 (I674363,I674355);
nor I_39520 (I674035,I674134,I674363);
or I_39521 (I674394,I674202,I250922);
nor I_39522 (I674411,I250922,I250919);
nand I_39523 (I674428,I674267,I674411);
nand I_39524 (I674445,I674394,I674428);
DFFARX1 I_39525 (I674445,I2507,I674049,I674038,);
nor I_39526 (I674476,I674411,I674168);
DFFARX1 I_39527 (I674476,I2507,I674049,I674017,);
nor I_39528 (I674507,I250922,I250925);
DFFARX1 I_39529 (I674507,I2507,I674049,I674533,);
DFFARX1 I_39530 (I674533,I2507,I674049,I674032,);
not I_39531 (I674555,I674533);
nand I_39532 (I674029,I674555,I674083);
nand I_39533 (I674023,I674555,I674185);
not I_39534 (I674627,I2514);
DFFARX1 I_39535 (I11958,I2507,I674627,I674653,);
nand I_39536 (I674661,I674653,I11952);
not I_39537 (I674678,I674661);
DFFARX1 I_39538 (I11970,I2507,I674627,I674704,);
not I_39539 (I674712,I674704);
not I_39540 (I674729,I11973);
or I_39541 (I674746,I11976,I11973);
nor I_39542 (I674763,I11976,I11973);
or I_39543 (I674780,I11961,I11976);
DFFARX1 I_39544 (I674780,I2507,I674627,I674619,);
not I_39545 (I674811,I11964);
nand I_39546 (I674828,I674811,I11967);
nand I_39547 (I674845,I674729,I674828);
and I_39548 (I674598,I674712,I674845);
nor I_39549 (I674876,I11964,I11955);
and I_39550 (I674893,I674712,I674876);
nor I_39551 (I674604,I674678,I674893);
DFFARX1 I_39552 (I674876,I2507,I674627,I674933,);
not I_39553 (I674941,I674933);
nor I_39554 (I674613,I674712,I674941);
or I_39555 (I674972,I674780,I11955);
nor I_39556 (I674989,I11955,I11961);
nand I_39557 (I675006,I674845,I674989);
nand I_39558 (I675023,I674972,I675006);
DFFARX1 I_39559 (I675023,I2507,I674627,I674616,);
nor I_39560 (I675054,I674989,I674746);
DFFARX1 I_39561 (I675054,I2507,I674627,I674595,);
nor I_39562 (I675085,I11955,I11952);
DFFARX1 I_39563 (I675085,I2507,I674627,I675111,);
DFFARX1 I_39564 (I675111,I2507,I674627,I674610,);
not I_39565 (I675133,I675111);
nand I_39566 (I674607,I675133,I674661);
nand I_39567 (I674601,I675133,I674763);
not I_39568 (I675205,I2514);
DFFARX1 I_39569 (I394061,I2507,I675205,I675231,);
nand I_39570 (I675239,I675231,I394064);
not I_39571 (I675256,I675239);
DFFARX1 I_39572 (I394076,I2507,I675205,I675282,);
not I_39573 (I675290,I675282);
not I_39574 (I675307,I394061);
or I_39575 (I675324,I394070,I394061);
nor I_39576 (I675341,I394070,I394061);
or I_39577 (I675358,I394079,I394070);
DFFARX1 I_39578 (I675358,I2507,I675205,I675197,);
not I_39579 (I675389,I394082);
nand I_39580 (I675406,I675389,I394064);
nand I_39581 (I675423,I675307,I675406);
and I_39582 (I675176,I675290,I675423);
nor I_39583 (I675454,I394082,I394067);
and I_39584 (I675471,I675290,I675454);
nor I_39585 (I675182,I675256,I675471);
DFFARX1 I_39586 (I675454,I2507,I675205,I675511,);
not I_39587 (I675519,I675511);
nor I_39588 (I675191,I675290,I675519);
or I_39589 (I675550,I675358,I394073);
nor I_39590 (I675567,I394073,I394079);
nand I_39591 (I675584,I675423,I675567);
nand I_39592 (I675601,I675550,I675584);
DFFARX1 I_39593 (I675601,I2507,I675205,I675194,);
nor I_39594 (I675632,I675567,I675324);
DFFARX1 I_39595 (I675632,I2507,I675205,I675173,);
nor I_39596 (I675663,I394073,I394085);
DFFARX1 I_39597 (I675663,I2507,I675205,I675689,);
DFFARX1 I_39598 (I675689,I2507,I675205,I675188,);
not I_39599 (I675711,I675689);
nand I_39600 (I675185,I675711,I675239);
nand I_39601 (I675179,I675711,I675341);
not I_39602 (I675783,I2514);
DFFARX1 I_39603 (I55178,I2507,I675783,I675809,);
nand I_39604 (I675817,I675809,I55169);
not I_39605 (I675834,I675817);
DFFARX1 I_39606 (I55166,I2507,I675783,I675860,);
not I_39607 (I675868,I675860);
not I_39608 (I675885,I55175);
or I_39609 (I675902,I55166,I55175);
nor I_39610 (I675919,I55166,I55175);
or I_39611 (I675936,I55172,I55166);
DFFARX1 I_39612 (I675936,I2507,I675783,I675775,);
not I_39613 (I675967,I55181);
nand I_39614 (I675984,I675967,I55190);
nand I_39615 (I676001,I675885,I675984);
and I_39616 (I675754,I675868,I676001);
nor I_39617 (I676032,I55181,I55184);
and I_39618 (I676049,I675868,I676032);
nor I_39619 (I675760,I675834,I676049);
DFFARX1 I_39620 (I676032,I2507,I675783,I676089,);
not I_39621 (I676097,I676089);
nor I_39622 (I675769,I675868,I676097);
or I_39623 (I676128,I675936,I55169);
nor I_39624 (I676145,I55169,I55172);
nand I_39625 (I676162,I676001,I676145);
nand I_39626 (I676179,I676128,I676162);
DFFARX1 I_39627 (I676179,I2507,I675783,I675772,);
nor I_39628 (I676210,I676145,I675902);
DFFARX1 I_39629 (I676210,I2507,I675783,I675751,);
nor I_39630 (I676241,I55169,I55187);
DFFARX1 I_39631 (I676241,I2507,I675783,I676267,);
DFFARX1 I_39632 (I676267,I2507,I675783,I675766,);
not I_39633 (I676289,I676267);
nand I_39634 (I675763,I676289,I675817);
nand I_39635 (I675757,I676289,I675919);
not I_39636 (I676361,I2514);
DFFARX1 I_39637 (I533858,I2507,I676361,I676387,);
nand I_39638 (I676395,I676387,I533879);
not I_39639 (I676412,I676395);
DFFARX1 I_39640 (I533852,I2507,I676361,I676438,);
not I_39641 (I676446,I676438);
not I_39642 (I676463,I533873);
or I_39643 (I676480,I533864,I533873);
nor I_39644 (I676497,I533864,I533873);
or I_39645 (I676514,I533867,I533864);
DFFARX1 I_39646 (I676514,I2507,I676361,I676353,);
not I_39647 (I676545,I533855);
nand I_39648 (I676562,I676545,I533870);
nand I_39649 (I676579,I676463,I676562);
and I_39650 (I676332,I676446,I676579);
nor I_39651 (I676610,I533855,I533852);
and I_39652 (I676627,I676446,I676610);
nor I_39653 (I676338,I676412,I676627);
DFFARX1 I_39654 (I676610,I2507,I676361,I676667,);
not I_39655 (I676675,I676667);
nor I_39656 (I676347,I676446,I676675);
or I_39657 (I676706,I676514,I533876);
nor I_39658 (I676723,I533876,I533867);
nand I_39659 (I676740,I676579,I676723);
nand I_39660 (I676757,I676706,I676740);
DFFARX1 I_39661 (I676757,I2507,I676361,I676350,);
nor I_39662 (I676788,I676723,I676480);
DFFARX1 I_39663 (I676788,I2507,I676361,I676329,);
nor I_39664 (I676819,I533876,I533861);
DFFARX1 I_39665 (I676819,I2507,I676361,I676845,);
DFFARX1 I_39666 (I676845,I2507,I676361,I676344,);
not I_39667 (I676867,I676845);
nand I_39668 (I676341,I676867,I676395);
nand I_39669 (I676335,I676867,I676497);
not I_39670 (I676939,I2514);
DFFARX1 I_39671 (I244379,I2507,I676939,I676965,);
nand I_39672 (I676973,I676965,I244388);
not I_39673 (I676990,I676973);
DFFARX1 I_39674 (I244376,I2507,I676939,I677016,);
not I_39675 (I677024,I677016);
not I_39676 (I677041,I244382);
or I_39677 (I677058,I244376,I244382);
nor I_39678 (I677075,I244376,I244382);
or I_39679 (I677092,I244391,I244376);
DFFARX1 I_39680 (I677092,I2507,I676939,I676931,);
not I_39681 (I677123,I244385);
nand I_39682 (I677140,I677123,I244400);
nand I_39683 (I677157,I677041,I677140);
and I_39684 (I676910,I677024,I677157);
nor I_39685 (I677188,I244385,I244403);
and I_39686 (I677205,I677024,I677188);
nor I_39687 (I676916,I676990,I677205);
DFFARX1 I_39688 (I677188,I2507,I676939,I677245,);
not I_39689 (I677253,I677245);
nor I_39690 (I676925,I677024,I677253);
or I_39691 (I677284,I677092,I244394);
nor I_39692 (I677301,I244394,I244391);
nand I_39693 (I677318,I677157,I677301);
nand I_39694 (I677335,I677284,I677318);
DFFARX1 I_39695 (I677335,I2507,I676939,I676928,);
nor I_39696 (I677366,I677301,I677058);
DFFARX1 I_39697 (I677366,I2507,I676939,I676907,);
nor I_39698 (I677397,I244394,I244397);
DFFARX1 I_39699 (I677397,I2507,I676939,I677423,);
DFFARX1 I_39700 (I677423,I2507,I676939,I676922,);
not I_39701 (I677445,I677423);
nand I_39702 (I676919,I677445,I676973);
nand I_39703 (I676913,I677445,I677075);
not I_39704 (I677517,I2514);
DFFARX1 I_39705 (I445506,I2507,I677517,I677543,);
nand I_39706 (I677551,I677543,I445506);
not I_39707 (I677568,I677551);
DFFARX1 I_39708 (I445512,I2507,I677517,I677594,);
not I_39709 (I677602,I677594);
not I_39710 (I677619,I445524);
or I_39711 (I677636,I445509,I445524);
nor I_39712 (I677653,I445509,I445524);
or I_39713 (I677670,I445503,I445509);
DFFARX1 I_39714 (I677670,I2507,I677517,I677509,);
not I_39715 (I677701,I445521);
nand I_39716 (I677718,I677701,I445515);
nand I_39717 (I677735,I677619,I677718);
and I_39718 (I677488,I677602,I677735);
nor I_39719 (I677766,I445521,I445503);
and I_39720 (I677783,I677602,I677766);
nor I_39721 (I677494,I677568,I677783);
DFFARX1 I_39722 (I677766,I2507,I677517,I677823,);
not I_39723 (I677831,I677823);
nor I_39724 (I677503,I677602,I677831);
or I_39725 (I677862,I677670,I445518);
nor I_39726 (I677879,I445518,I445503);
nand I_39727 (I677896,I677735,I677879);
nand I_39728 (I677913,I677862,I677896);
DFFARX1 I_39729 (I677913,I2507,I677517,I677506,);
nor I_39730 (I677944,I677879,I677636);
DFFARX1 I_39731 (I677944,I2507,I677517,I677485,);
nor I_39732 (I677975,I445518,I445509);
DFFARX1 I_39733 (I677975,I2507,I677517,I678001,);
DFFARX1 I_39734 (I678001,I2507,I677517,I677500,);
not I_39735 (I678023,I678001);
nand I_39736 (I677497,I678023,I677551);
nand I_39737 (I677491,I678023,I677653);
not I_39738 (I678095,I2514);
DFFARX1 I_39739 (I613889,I2507,I678095,I678121,);
nand I_39740 (I678129,I678121,I613874);
not I_39741 (I678146,I678129);
DFFARX1 I_39742 (I613877,I2507,I678095,I678172,);
not I_39743 (I678180,I678172);
not I_39744 (I678197,I613892);
or I_39745 (I678214,I613895,I613892);
nor I_39746 (I678231,I613895,I613892);
or I_39747 (I678248,I613871,I613895);
DFFARX1 I_39748 (I678248,I2507,I678095,I678087,);
not I_39749 (I678279,I613883);
nand I_39750 (I678296,I678279,I613886);
nand I_39751 (I678313,I678197,I678296);
and I_39752 (I678066,I678180,I678313);
nor I_39753 (I678344,I613883,I613880);
and I_39754 (I678361,I678180,I678344);
nor I_39755 (I678072,I678146,I678361);
DFFARX1 I_39756 (I678344,I2507,I678095,I678401,);
not I_39757 (I678409,I678401);
nor I_39758 (I678081,I678180,I678409);
or I_39759 (I678440,I678248,I613871);
nor I_39760 (I678457,I613871,I613871);
nand I_39761 (I678474,I678313,I678457);
nand I_39762 (I678491,I678440,I678474);
DFFARX1 I_39763 (I678491,I2507,I678095,I678084,);
nor I_39764 (I678522,I678457,I678214);
DFFARX1 I_39765 (I678522,I2507,I678095,I678063,);
nor I_39766 (I678553,I613871,I613874);
DFFARX1 I_39767 (I678553,I2507,I678095,I678579,);
DFFARX1 I_39768 (I678579,I2507,I678095,I678078,);
not I_39769 (I678601,I678579);
nand I_39770 (I678075,I678601,I678129);
nand I_39771 (I678069,I678601,I678231);
not I_39772 (I678673,I2514);
DFFARX1 I_39773 (I725177,I2507,I678673,I678699,);
nand I_39774 (I678707,I678699,I725168);
not I_39775 (I678724,I678707);
DFFARX1 I_39776 (I725153,I2507,I678673,I678750,);
not I_39777 (I678758,I678750);
not I_39778 (I678775,I725156);
or I_39779 (I678792,I725165,I725156);
nor I_39780 (I678809,I725165,I725156);
or I_39781 (I678826,I725162,I725165);
DFFARX1 I_39782 (I678826,I2507,I678673,I678665,);
not I_39783 (I678857,I725174);
nand I_39784 (I678874,I678857,I725153);
nand I_39785 (I678891,I678775,I678874);
and I_39786 (I678644,I678758,I678891);
nor I_39787 (I678922,I725174,I725159);
and I_39788 (I678939,I678758,I678922);
nor I_39789 (I678650,I678724,I678939);
DFFARX1 I_39790 (I678922,I2507,I678673,I678979,);
not I_39791 (I678987,I678979);
nor I_39792 (I678659,I678758,I678987);
or I_39793 (I679018,I678826,I725180);
nor I_39794 (I679035,I725180,I725162);
nand I_39795 (I679052,I678891,I679035);
nand I_39796 (I679069,I679018,I679052);
DFFARX1 I_39797 (I679069,I2507,I678673,I678662,);
nor I_39798 (I679100,I679035,I678792);
DFFARX1 I_39799 (I679100,I2507,I678673,I678641,);
nor I_39800 (I679131,I725180,I725171);
DFFARX1 I_39801 (I679131,I2507,I678673,I679157,);
DFFARX1 I_39802 (I679157,I2507,I678673,I678656,);
not I_39803 (I679179,I679157);
nand I_39804 (I678653,I679179,I678707);
nand I_39805 (I678647,I679179,I678809);
not I_39806 (I679251,I2514);
DFFARX1 I_39807 (I318924,I2507,I679251,I679277,);
nand I_39808 (I679285,I679277,I318939);
not I_39809 (I679302,I679285);
DFFARX1 I_39810 (I318921,I2507,I679251,I679328,);
not I_39811 (I679336,I679328);
not I_39812 (I679353,I318930);
or I_39813 (I679370,I318924,I318930);
nor I_39814 (I679387,I318924,I318930);
or I_39815 (I679404,I318921,I318924);
DFFARX1 I_39816 (I679404,I2507,I679251,I679243,);
not I_39817 (I679435,I318942);
nand I_39818 (I679452,I679435,I318945);
nand I_39819 (I679469,I679353,I679452);
and I_39820 (I679222,I679336,I679469);
nor I_39821 (I679500,I318942,I318927);
and I_39822 (I679517,I679336,I679500);
nor I_39823 (I679228,I679302,I679517);
DFFARX1 I_39824 (I679500,I2507,I679251,I679557,);
not I_39825 (I679565,I679557);
nor I_39826 (I679237,I679336,I679565);
or I_39827 (I679596,I679404,I318933);
nor I_39828 (I679613,I318933,I318921);
nand I_39829 (I679630,I679469,I679613);
nand I_39830 (I679647,I679596,I679630);
DFFARX1 I_39831 (I679647,I2507,I679251,I679240,);
nor I_39832 (I679678,I679613,I679370);
DFFARX1 I_39833 (I679678,I2507,I679251,I679219,);
nor I_39834 (I679709,I318933,I318936);
DFFARX1 I_39835 (I679709,I2507,I679251,I679735,);
DFFARX1 I_39836 (I679735,I2507,I679251,I679234,);
not I_39837 (I679757,I679735);
nand I_39838 (I679231,I679757,I679285);
nand I_39839 (I679225,I679757,I679387);
not I_39840 (I679829,I2514);
DFFARX1 I_39841 (I170602,I2507,I679829,I679855,);
nand I_39842 (I679863,I679855,I170623);
not I_39843 (I679880,I679863);
DFFARX1 I_39844 (I170617,I2507,I679829,I679906,);
not I_39845 (I679914,I679906);
not I_39846 (I679931,I170605);
or I_39847 (I679948,I170620,I170605);
nor I_39848 (I679965,I170620,I170605);
or I_39849 (I679982,I170611,I170620);
DFFARX1 I_39850 (I679982,I2507,I679829,I679821,);
not I_39851 (I680013,I170599);
nand I_39852 (I680030,I680013,I170596);
nand I_39853 (I680047,I679931,I680030);
and I_39854 (I679800,I679914,I680047);
nor I_39855 (I680078,I170599,I170608);
and I_39856 (I680095,I679914,I680078);
nor I_39857 (I679806,I679880,I680095);
DFFARX1 I_39858 (I680078,I2507,I679829,I680135,);
not I_39859 (I680143,I680135);
nor I_39860 (I679815,I679914,I680143);
or I_39861 (I680174,I679982,I170614);
nor I_39862 (I680191,I170614,I170611);
nand I_39863 (I680208,I680047,I680191);
nand I_39864 (I680225,I680174,I680208);
DFFARX1 I_39865 (I680225,I2507,I679829,I679818,);
nor I_39866 (I680256,I680191,I679948);
DFFARX1 I_39867 (I680256,I2507,I679829,I679797,);
nor I_39868 (I680287,I170614,I170596);
DFFARX1 I_39869 (I680287,I2507,I679829,I680313,);
DFFARX1 I_39870 (I680313,I2507,I679829,I679812,);
not I_39871 (I680335,I680313);
nand I_39872 (I679809,I680335,I679863);
nand I_39873 (I679803,I680335,I679965);
not I_39874 (I680407,I2514);
DFFARX1 I_39875 (I490576,I2507,I680407,I680433,);
nand I_39876 (I680441,I680433,I490597);
not I_39877 (I680458,I680441);
DFFARX1 I_39878 (I490570,I2507,I680407,I680484,);
not I_39879 (I680492,I680484);
not I_39880 (I680509,I490591);
or I_39881 (I680526,I490582,I490591);
nor I_39882 (I680543,I490582,I490591);
or I_39883 (I680560,I490585,I490582);
DFFARX1 I_39884 (I680560,I2507,I680407,I680399,);
not I_39885 (I680591,I490573);
nand I_39886 (I680608,I680591,I490588);
nand I_39887 (I680625,I680509,I680608);
and I_39888 (I680378,I680492,I680625);
nor I_39889 (I680656,I490573,I490570);
and I_39890 (I680673,I680492,I680656);
nor I_39891 (I680384,I680458,I680673);
DFFARX1 I_39892 (I680656,I2507,I680407,I680713,);
not I_39893 (I680721,I680713);
nor I_39894 (I680393,I680492,I680721);
or I_39895 (I680752,I680560,I490594);
nor I_39896 (I680769,I490594,I490585);
nand I_39897 (I680786,I680625,I680769);
nand I_39898 (I680803,I680752,I680786);
DFFARX1 I_39899 (I680803,I2507,I680407,I680396,);
nor I_39900 (I680834,I680769,I680526);
DFFARX1 I_39901 (I680834,I2507,I680407,I680375,);
nor I_39902 (I680865,I490594,I490579);
DFFARX1 I_39903 (I680865,I2507,I680407,I680891,);
DFFARX1 I_39904 (I680891,I2507,I680407,I680390,);
not I_39905 (I680913,I680891);
nand I_39906 (I680387,I680913,I680441);
nand I_39907 (I680381,I680913,I680543);
not I_39908 (I680985,I2514);
DFFARX1 I_39909 (I543041,I2507,I680985,I681011,);
nand I_39910 (I681019,I681011,I543038);
not I_39911 (I681036,I681019);
DFFARX1 I_39912 (I543038,I2507,I680985,I681062,);
not I_39913 (I681070,I681062);
not I_39914 (I681087,I543035);
or I_39915 (I681104,I543044,I543035);
nor I_39916 (I681121,I543044,I543035);
or I_39917 (I681138,I543047,I543044);
DFFARX1 I_39918 (I681138,I2507,I680985,I680977,);
not I_39919 (I681169,I543035);
nand I_39920 (I681186,I681169,I543032);
nand I_39921 (I681203,I681087,I681186);
and I_39922 (I680956,I681070,I681203);
nor I_39923 (I681234,I543035,I543050);
and I_39924 (I681251,I681070,I681234);
nor I_39925 (I680962,I681036,I681251);
DFFARX1 I_39926 (I681234,I2507,I680985,I681291,);
not I_39927 (I681299,I681291);
nor I_39928 (I680971,I681070,I681299);
or I_39929 (I681330,I681138,I543053);
nor I_39930 (I681347,I543053,I543047);
nand I_39931 (I681364,I681203,I681347);
nand I_39932 (I681381,I681330,I681364);
DFFARX1 I_39933 (I681381,I2507,I680985,I680974,);
nor I_39934 (I681412,I681347,I681104);
DFFARX1 I_39935 (I681412,I2507,I680985,I680953,);
nor I_39936 (I681443,I543053,I543032);
DFFARX1 I_39937 (I681443,I2507,I680985,I681469,);
DFFARX1 I_39938 (I681469,I2507,I680985,I680968,);
not I_39939 (I681491,I681469);
nand I_39940 (I680965,I681491,I681019);
nand I_39941 (I680959,I681491,I681121);
not I_39942 (I681563,I2514);
DFFARX1 I_39943 (I383079,I2507,I681563,I681589,);
nand I_39944 (I681597,I681589,I383082);
not I_39945 (I681614,I681597);
DFFARX1 I_39946 (I383094,I2507,I681563,I681640,);
not I_39947 (I681648,I681640);
not I_39948 (I681665,I383079);
or I_39949 (I681682,I383088,I383079);
nor I_39950 (I681699,I383088,I383079);
or I_39951 (I681716,I383097,I383088);
DFFARX1 I_39952 (I681716,I2507,I681563,I681555,);
not I_39953 (I681747,I383100);
nand I_39954 (I681764,I681747,I383082);
nand I_39955 (I681781,I681665,I681764);
and I_39956 (I681534,I681648,I681781);
nor I_39957 (I681812,I383100,I383085);
and I_39958 (I681829,I681648,I681812);
nor I_39959 (I681540,I681614,I681829);
DFFARX1 I_39960 (I681812,I2507,I681563,I681869,);
not I_39961 (I681877,I681869);
nor I_39962 (I681549,I681648,I681877);
or I_39963 (I681908,I681716,I383091);
nor I_39964 (I681925,I383091,I383097);
nand I_39965 (I681942,I681781,I681925);
nand I_39966 (I681959,I681908,I681942);
DFFARX1 I_39967 (I681959,I2507,I681563,I681552,);
nor I_39968 (I681990,I681925,I681682);
DFFARX1 I_39969 (I681990,I2507,I681563,I681531,);
nor I_39970 (I682021,I383091,I383103);
DFFARX1 I_39971 (I682021,I2507,I681563,I682047,);
DFFARX1 I_39972 (I682047,I2507,I681563,I681546,);
not I_39973 (I682069,I682047);
nand I_39974 (I681543,I682069,I681597);
nand I_39975 (I681537,I682069,I681699);
not I_39976 (I682141,I2514);
DFFARX1 I_39977 (I182196,I2507,I682141,I682167,);
nand I_39978 (I682175,I682167,I182217);
not I_39979 (I682192,I682175);
DFFARX1 I_39980 (I182211,I2507,I682141,I682218,);
not I_39981 (I682226,I682218);
not I_39982 (I682243,I182199);
or I_39983 (I682260,I182214,I182199);
nor I_39984 (I682277,I182214,I182199);
or I_39985 (I682294,I182205,I182214);
DFFARX1 I_39986 (I682294,I2507,I682141,I682133,);
not I_39987 (I682325,I182193);
nand I_39988 (I682342,I682325,I182190);
nand I_39989 (I682359,I682243,I682342);
and I_39990 (I682112,I682226,I682359);
nor I_39991 (I682390,I182193,I182202);
and I_39992 (I682407,I682226,I682390);
nor I_39993 (I682118,I682192,I682407);
DFFARX1 I_39994 (I682390,I2507,I682141,I682447,);
not I_39995 (I682455,I682447);
nor I_39996 (I682127,I682226,I682455);
or I_39997 (I682486,I682294,I182208);
nor I_39998 (I682503,I182208,I182205);
nand I_39999 (I682520,I682359,I682503);
nand I_40000 (I682537,I682486,I682520);
DFFARX1 I_40001 (I682537,I2507,I682141,I682130,);
nor I_40002 (I682568,I682503,I682260);
DFFARX1 I_40003 (I682568,I2507,I682141,I682109,);
nor I_40004 (I682599,I182208,I182190);
DFFARX1 I_40005 (I682599,I2507,I682141,I682625,);
DFFARX1 I_40006 (I682625,I2507,I682141,I682124,);
not I_40007 (I682647,I682625);
nand I_40008 (I682121,I682647,I682175);
nand I_40009 (I682115,I682647,I682277);
not I_40010 (I682719,I2514);
DFFARX1 I_40011 (I433912,I2507,I682719,I682745,);
nand I_40012 (I682753,I682745,I433912);
not I_40013 (I682770,I682753);
DFFARX1 I_40014 (I433918,I2507,I682719,I682796,);
not I_40015 (I682804,I682796);
not I_40016 (I682821,I433930);
or I_40017 (I682838,I433915,I433930);
nor I_40018 (I682855,I433915,I433930);
or I_40019 (I682872,I433909,I433915);
DFFARX1 I_40020 (I682872,I2507,I682719,I682711,);
not I_40021 (I682903,I433927);
nand I_40022 (I682920,I682903,I433921);
nand I_40023 (I682937,I682821,I682920);
and I_40024 (I682690,I682804,I682937);
nor I_40025 (I682968,I433927,I433909);
and I_40026 (I682985,I682804,I682968);
nor I_40027 (I682696,I682770,I682985);
DFFARX1 I_40028 (I682968,I2507,I682719,I683025,);
not I_40029 (I683033,I683025);
nor I_40030 (I682705,I682804,I683033);
or I_40031 (I683064,I682872,I433924);
nor I_40032 (I683081,I433924,I433909);
nand I_40033 (I683098,I682937,I683081);
nand I_40034 (I683115,I683064,I683098);
DFFARX1 I_40035 (I683115,I2507,I682719,I682708,);
nor I_40036 (I683146,I683081,I682838);
DFFARX1 I_40037 (I683146,I2507,I682719,I682687,);
nor I_40038 (I683177,I433924,I433915);
DFFARX1 I_40039 (I683177,I2507,I682719,I683203,);
DFFARX1 I_40040 (I683203,I2507,I682719,I682702,);
not I_40041 (I683225,I683203);
nand I_40042 (I682699,I683225,I682753);
nand I_40043 (I682693,I683225,I682855);
not I_40044 (I683297,I2514);
DFFARX1 I_40045 (I596549,I2507,I683297,I683323,);
nand I_40046 (I683331,I683323,I596534);
not I_40047 (I683348,I683331);
DFFARX1 I_40048 (I596537,I2507,I683297,I683374,);
not I_40049 (I683382,I683374);
not I_40050 (I683399,I596552);
or I_40051 (I683416,I596555,I596552);
nor I_40052 (I683433,I596555,I596552);
or I_40053 (I683450,I596531,I596555);
DFFARX1 I_40054 (I683450,I2507,I683297,I683289,);
not I_40055 (I683481,I596543);
nand I_40056 (I683498,I683481,I596546);
nand I_40057 (I683515,I683399,I683498);
and I_40058 (I683268,I683382,I683515);
nor I_40059 (I683546,I596543,I596540);
and I_40060 (I683563,I683382,I683546);
nor I_40061 (I683274,I683348,I683563);
DFFARX1 I_40062 (I683546,I2507,I683297,I683603,);
not I_40063 (I683611,I683603);
nor I_40064 (I683283,I683382,I683611);
or I_40065 (I683642,I683450,I596531);
nor I_40066 (I683659,I596531,I596531);
nand I_40067 (I683676,I683515,I683659);
nand I_40068 (I683693,I683642,I683676);
DFFARX1 I_40069 (I683693,I2507,I683297,I683286,);
nor I_40070 (I683724,I683659,I683416);
DFFARX1 I_40071 (I683724,I2507,I683297,I683265,);
nor I_40072 (I683755,I596531,I596534);
DFFARX1 I_40073 (I683755,I2507,I683297,I683781,);
DFFARX1 I_40074 (I683781,I2507,I683297,I683280,);
not I_40075 (I683803,I683781);
nand I_40076 (I683277,I683803,I683331);
nand I_40077 (I683271,I683803,I683433);
not I_40078 (I683878,I2514);
DFFARX1 I_40079 (I360555,I2507,I683878,I683904,);
nand I_40080 (I683912,I683904,I360540);
not I_40081 (I683929,I683912);
DFFARX1 I_40082 (I360558,I2507,I683878,I683955,);
not I_40083 (I683963,I683955);
nor I_40084 (I683980,I360537,I360552);
not I_40085 (I683997,I683980);
DFFARX1 I_40086 (I683997,I2507,I683878,I683864,);
or I_40087 (I684028,I360549,I360537);
DFFARX1 I_40088 (I684028,I2507,I683878,I683867,);
not I_40089 (I684059,I360537);
nor I_40090 (I684076,I684059,I360546);
nor I_40091 (I684093,I684076,I360552);
nor I_40092 (I684110,I360546,I360540);
nor I_40093 (I684127,I683963,I684110);
nor I_40094 (I683852,I683929,I684127);
not I_40095 (I684158,I684110);
nand I_40096 (I683855,I684158,I683912);
nand I_40097 (I683849,I684158,I683980);
nor I_40098 (I683846,I684110,I684093);
nor I_40099 (I684217,I360543,I360549);
not I_40100 (I684234,I684217);
DFFARX1 I_40101 (I684217,I2507,I683878,I684260,);
not I_40102 (I683870,I684260);
nor I_40103 (I684282,I360543,I360561);
DFFARX1 I_40104 (I684282,I2507,I683878,I684308,);
and I_40105 (I684316,I684308,I360537);
nor I_40106 (I684333,I684316,I684234);
DFFARX1 I_40107 (I684333,I2507,I683878,I683861,);
nor I_40108 (I684364,I684308,I684093);
DFFARX1 I_40109 (I684364,I2507,I683878,I683843,);
nor I_40110 (I683858,I684308,I683997);
not I_40111 (I684439,I2514);
DFFARX1 I_40112 (I133009,I2507,I684439,I684465,);
nand I_40113 (I684473,I684465,I133033);
not I_40114 (I684490,I684473);
DFFARX1 I_40115 (I133021,I2507,I684439,I684516,);
not I_40116 (I684524,I684516);
nor I_40117 (I684541,I133012,I133030);
not I_40118 (I684558,I684541);
DFFARX1 I_40119 (I684558,I2507,I684439,I684425,);
or I_40120 (I684589,I133024,I133012);
DFFARX1 I_40121 (I684589,I2507,I684439,I684428,);
not I_40122 (I684620,I133012);
nor I_40123 (I684637,I684620,I133027);
nor I_40124 (I684654,I684637,I133030);
nor I_40125 (I684671,I133027,I133018);
nor I_40126 (I684688,I684524,I684671);
nor I_40127 (I684413,I684490,I684688);
not I_40128 (I684719,I684671);
nand I_40129 (I684416,I684719,I684473);
nand I_40130 (I684410,I684719,I684541);
nor I_40131 (I684407,I684671,I684654);
nor I_40132 (I684778,I133015,I133024);
not I_40133 (I684795,I684778);
DFFARX1 I_40134 (I684778,I2507,I684439,I684821,);
not I_40135 (I684431,I684821);
nor I_40136 (I684843,I133015,I133009);
DFFARX1 I_40137 (I684843,I2507,I684439,I684869,);
and I_40138 (I684877,I684869,I133012);
nor I_40139 (I684894,I684877,I684795);
DFFARX1 I_40140 (I684894,I2507,I684439,I684422,);
nor I_40141 (I684925,I684869,I684654);
DFFARX1 I_40142 (I684925,I2507,I684439,I684404,);
nor I_40143 (I684419,I684869,I684558);
not I_40144 (I685000,I2514);
DFFARX1 I_40145 (I703153,I2507,I685000,I685026,);
nand I_40146 (I685034,I685026,I703147);
not I_40147 (I685051,I685034);
DFFARX1 I_40148 (I703165,I2507,I685000,I685077,);
not I_40149 (I685085,I685077);
nor I_40150 (I685102,I703150,I703141);
not I_40151 (I685119,I685102);
DFFARX1 I_40152 (I685119,I2507,I685000,I684986,);
or I_40153 (I685150,I703156,I703150);
DFFARX1 I_40154 (I685150,I2507,I685000,I684989,);
not I_40155 (I685181,I703159);
nor I_40156 (I685198,I685181,I703162);
nor I_40157 (I685215,I685198,I703141);
nor I_40158 (I685232,I703162,I703144);
nor I_40159 (I685249,I685085,I685232);
nor I_40160 (I684974,I685051,I685249);
not I_40161 (I685280,I685232);
nand I_40162 (I684977,I685280,I685034);
nand I_40163 (I684971,I685280,I685102);
nor I_40164 (I684968,I685232,I685215);
nor I_40165 (I685339,I703138,I703156);
not I_40166 (I685356,I685339);
DFFARX1 I_40167 (I685339,I2507,I685000,I685382,);
not I_40168 (I684992,I685382);
nor I_40169 (I685404,I703138,I703138);
DFFARX1 I_40170 (I685404,I2507,I685000,I685430,);
and I_40171 (I685438,I685430,I703150);
nor I_40172 (I685455,I685438,I685356);
DFFARX1 I_40173 (I685455,I2507,I685000,I684983,);
nor I_40174 (I685486,I685430,I685215);
DFFARX1 I_40175 (I685486,I2507,I685000,I684965,);
nor I_40176 (I684980,I685430,I685119);
not I_40177 (I685561,I2514);
DFFARX1 I_40178 (I302761,I2507,I685561,I685587,);
nand I_40179 (I685595,I685587,I302740);
not I_40180 (I685612,I685595);
DFFARX1 I_40181 (I302752,I2507,I685561,I685638,);
not I_40182 (I685646,I685638);
nor I_40183 (I685663,I302740,I302749);
not I_40184 (I685680,I685663);
DFFARX1 I_40185 (I685680,I2507,I685561,I685547,);
or I_40186 (I685711,I302743,I302740);
DFFARX1 I_40187 (I685711,I2507,I685561,I685550,);
not I_40188 (I685742,I302746);
nor I_40189 (I685759,I685742,I302737);
nor I_40190 (I685776,I685759,I302749);
nor I_40191 (I685793,I302737,I302755);
nor I_40192 (I685810,I685646,I685793);
nor I_40193 (I685535,I685612,I685810);
not I_40194 (I685841,I685793);
nand I_40195 (I685538,I685841,I685595);
nand I_40196 (I685532,I685841,I685663);
nor I_40197 (I685529,I685793,I685776);
nor I_40198 (I685900,I302758,I302743);
not I_40199 (I685917,I685900);
DFFARX1 I_40200 (I685900,I2507,I685561,I685943,);
not I_40201 (I685553,I685943);
nor I_40202 (I685965,I302758,I302737);
DFFARX1 I_40203 (I685965,I2507,I685561,I685991,);
and I_40204 (I685999,I685991,I302740);
nor I_40205 (I686016,I685999,I685917);
DFFARX1 I_40206 (I686016,I2507,I685561,I685544,);
nor I_40207 (I686047,I685991,I685776);
DFFARX1 I_40208 (I686047,I2507,I685561,I685526,);
nor I_40209 (I685541,I685991,I685680);
not I_40210 (I686122,I2514);
DFFARX1 I_40211 (I328771,I2507,I686122,I686148,);
nand I_40212 (I686156,I686148,I328750);
not I_40213 (I686173,I686156);
DFFARX1 I_40214 (I328762,I2507,I686122,I686199,);
not I_40215 (I686207,I686199);
nor I_40216 (I686224,I328750,I328759);
not I_40217 (I686241,I686224);
DFFARX1 I_40218 (I686241,I2507,I686122,I686108,);
or I_40219 (I686272,I328753,I328750);
DFFARX1 I_40220 (I686272,I2507,I686122,I686111,);
not I_40221 (I686303,I328756);
nor I_40222 (I686320,I686303,I328747);
nor I_40223 (I686337,I686320,I328759);
nor I_40224 (I686354,I328747,I328765);
nor I_40225 (I686371,I686207,I686354);
nor I_40226 (I686096,I686173,I686371);
not I_40227 (I686402,I686354);
nand I_40228 (I686099,I686402,I686156);
nand I_40229 (I686093,I686402,I686224);
nor I_40230 (I686090,I686354,I686337);
nor I_40231 (I686461,I328768,I328753);
not I_40232 (I686478,I686461);
DFFARX1 I_40233 (I686461,I2507,I686122,I686504,);
not I_40234 (I686114,I686504);
nor I_40235 (I686526,I328768,I328747);
DFFARX1 I_40236 (I686526,I2507,I686122,I686552,);
and I_40237 (I686560,I686552,I328750);
nor I_40238 (I686577,I686560,I686478);
DFFARX1 I_40239 (I686577,I2507,I686122,I686105,);
nor I_40240 (I686608,I686552,I686337);
DFFARX1 I_40241 (I686608,I2507,I686122,I686087,);
nor I_40242 (I686102,I686552,I686241);
not I_40243 (I686683,I2514);
DFFARX1 I_40244 (I345533,I2507,I686683,I686709,);
nand I_40245 (I686717,I686709,I345512);
not I_40246 (I686734,I686717);
DFFARX1 I_40247 (I345524,I2507,I686683,I686760,);
not I_40248 (I686768,I686760);
nor I_40249 (I686785,I345512,I345521);
not I_40250 (I686802,I686785);
DFFARX1 I_40251 (I686802,I2507,I686683,I686669,);
or I_40252 (I686833,I345515,I345512);
DFFARX1 I_40253 (I686833,I2507,I686683,I686672,);
not I_40254 (I686864,I345518);
nor I_40255 (I686881,I686864,I345509);
nor I_40256 (I686898,I686881,I345521);
nor I_40257 (I686915,I345509,I345527);
nor I_40258 (I686932,I686768,I686915);
nor I_40259 (I686657,I686734,I686932);
not I_40260 (I686963,I686915);
nand I_40261 (I686660,I686963,I686717);
nand I_40262 (I686654,I686963,I686785);
nor I_40263 (I686651,I686915,I686898);
nor I_40264 (I687022,I345530,I345515);
not I_40265 (I687039,I687022);
DFFARX1 I_40266 (I687022,I2507,I686683,I687065,);
not I_40267 (I686675,I687065);
nor I_40268 (I687087,I345530,I345509);
DFFARX1 I_40269 (I687087,I2507,I686683,I687113,);
and I_40270 (I687121,I687113,I345512);
nor I_40271 (I687138,I687121,I687039);
DFFARX1 I_40272 (I687138,I2507,I686683,I686666,);
nor I_40273 (I687169,I687113,I686898);
DFFARX1 I_40274 (I687169,I2507,I686683,I686648,);
nor I_40275 (I686663,I687113,I686802);
not I_40276 (I687244,I2514);
DFFARX1 I_40277 (I579772,I2507,I687244,I687270,);
nand I_40278 (I687278,I687270,I579769);
not I_40279 (I687295,I687278);
DFFARX1 I_40280 (I579772,I2507,I687244,I687321,);
not I_40281 (I687329,I687321);
nor I_40282 (I687346,I579790,I579784);
not I_40283 (I687363,I687346);
DFFARX1 I_40284 (I687363,I2507,I687244,I687230,);
or I_40285 (I687394,I579793,I579790);
DFFARX1 I_40286 (I687394,I2507,I687244,I687233,);
not I_40287 (I687425,I579781);
nor I_40288 (I687442,I687425,I579778);
nor I_40289 (I687459,I687442,I579784);
nor I_40290 (I687476,I579778,I579769);
nor I_40291 (I687493,I687329,I687476);
nor I_40292 (I687218,I687295,I687493);
not I_40293 (I687524,I687476);
nand I_40294 (I687221,I687524,I687278);
nand I_40295 (I687215,I687524,I687346);
nor I_40296 (I687212,I687476,I687459);
nor I_40297 (I687583,I579775,I579793);
not I_40298 (I687600,I687583);
DFFARX1 I_40299 (I687583,I2507,I687244,I687626,);
not I_40300 (I687236,I687626);
nor I_40301 (I687648,I579775,I579787);
DFFARX1 I_40302 (I687648,I2507,I687244,I687674,);
and I_40303 (I687682,I687674,I579790);
nor I_40304 (I687699,I687682,I687600);
DFFARX1 I_40305 (I687699,I2507,I687244,I687227,);
nor I_40306 (I687730,I687674,I687459);
DFFARX1 I_40307 (I687730,I2507,I687244,I687209,);
nor I_40308 (I687224,I687674,I687363);
not I_40309 (I687805,I2514);
DFFARX1 I_40310 (I509974,I2507,I687805,I687831,);
nand I_40311 (I687839,I687831,I509956);
not I_40312 (I687856,I687839);
DFFARX1 I_40313 (I509968,I2507,I687805,I687882,);
not I_40314 (I687890,I687882);
nor I_40315 (I687907,I509950,I509950);
not I_40316 (I687924,I687907);
DFFARX1 I_40317 (I687924,I2507,I687805,I687791,);
or I_40318 (I687955,I509962,I509950);
DFFARX1 I_40319 (I687955,I2507,I687805,I687794,);
not I_40320 (I687986,I509977);
nor I_40321 (I688003,I687986,I509965);
nor I_40322 (I688020,I688003,I509950);
nor I_40323 (I688037,I509965,I509953);
nor I_40324 (I688054,I687890,I688037);
nor I_40325 (I687779,I687856,I688054);
not I_40326 (I688085,I688037);
nand I_40327 (I687782,I688085,I687839);
nand I_40328 (I687776,I688085,I687907);
nor I_40329 (I687773,I688037,I688020);
nor I_40330 (I688144,I509959,I509962);
not I_40331 (I688161,I688144);
DFFARX1 I_40332 (I688144,I2507,I687805,I688187,);
not I_40333 (I687797,I688187);
nor I_40334 (I688209,I509959,I509971);
DFFARX1 I_40335 (I688209,I2507,I687805,I688235,);
and I_40336 (I688243,I688235,I509950);
nor I_40337 (I688260,I688243,I688161);
DFFARX1 I_40338 (I688260,I2507,I687805,I687788,);
nor I_40339 (I688291,I688235,I688020);
DFFARX1 I_40340 (I688291,I2507,I687805,I687770,);
nor I_40341 (I687785,I688235,I687924);
not I_40342 (I688366,I2514);
DFFARX1 I_40343 (I102069,I2507,I688366,I688392,);
nand I_40344 (I688400,I688392,I102093);
not I_40345 (I688417,I688400);
DFFARX1 I_40346 (I102081,I2507,I688366,I688443,);
not I_40347 (I688451,I688443);
nor I_40348 (I688468,I102072,I102090);
not I_40349 (I688485,I688468);
DFFARX1 I_40350 (I688485,I2507,I688366,I688352,);
or I_40351 (I688516,I102084,I102072);
DFFARX1 I_40352 (I688516,I2507,I688366,I688355,);
not I_40353 (I688547,I102072);
nor I_40354 (I688564,I688547,I102087);
nor I_40355 (I688581,I688564,I102090);
nor I_40356 (I688598,I102087,I102078);
nor I_40357 (I688615,I688451,I688598);
nor I_40358 (I688340,I688417,I688615);
not I_40359 (I688646,I688598);
nand I_40360 (I688343,I688646,I688400);
nand I_40361 (I688337,I688646,I688468);
nor I_40362 (I688334,I688598,I688581);
nor I_40363 (I688705,I102075,I102084);
not I_40364 (I688722,I688705);
DFFARX1 I_40365 (I688705,I2507,I688366,I688748,);
not I_40366 (I688358,I688748);
nor I_40367 (I688770,I102075,I102069);
DFFARX1 I_40368 (I688770,I2507,I688366,I688796,);
and I_40369 (I688804,I688796,I102072);
nor I_40370 (I688821,I688804,I688722);
DFFARX1 I_40371 (I688821,I2507,I688366,I688349,);
nor I_40372 (I688852,I688796,I688581);
DFFARX1 I_40373 (I688852,I2507,I688366,I688331,);
nor I_40374 (I688346,I688796,I688485);
not I_40375 (I688927,I2514);
DFFARX1 I_40376 (I88979,I2507,I688927,I688953,);
nand I_40377 (I688961,I688953,I89003);
not I_40378 (I688978,I688961);
DFFARX1 I_40379 (I88991,I2507,I688927,I689004,);
not I_40380 (I689012,I689004);
nor I_40381 (I689029,I88982,I89000);
not I_40382 (I689046,I689029);
DFFARX1 I_40383 (I689046,I2507,I688927,I688913,);
or I_40384 (I689077,I88994,I88982);
DFFARX1 I_40385 (I689077,I2507,I688927,I688916,);
not I_40386 (I689108,I88982);
nor I_40387 (I689125,I689108,I88997);
nor I_40388 (I689142,I689125,I89000);
nor I_40389 (I689159,I88997,I88988);
nor I_40390 (I689176,I689012,I689159);
nor I_40391 (I688901,I688978,I689176);
not I_40392 (I689207,I689159);
nand I_40393 (I688904,I689207,I688961);
nand I_40394 (I688898,I689207,I689029);
nor I_40395 (I688895,I689159,I689142);
nor I_40396 (I689266,I88985,I88994);
not I_40397 (I689283,I689266);
DFFARX1 I_40398 (I689266,I2507,I688927,I689309,);
not I_40399 (I688919,I689309);
nor I_40400 (I689331,I88985,I88979);
DFFARX1 I_40401 (I689331,I2507,I688927,I689357,);
and I_40402 (I689365,I689357,I88982);
nor I_40403 (I689382,I689365,I689283);
DFFARX1 I_40404 (I689382,I2507,I688927,I688910,);
nor I_40405 (I689413,I689357,I689142);
DFFARX1 I_40406 (I689413,I2507,I688927,I688892,);
nor I_40407 (I688907,I689357,I689046);
not I_40408 (I689488,I2514);
DFFARX1 I_40409 (I171671,I2507,I689488,I689514,);
DFFARX1 I_40410 (I171665,I2507,I689488,I689531,);
not I_40411 (I689539,I689531);
nor I_40412 (I689456,I689514,I689539);
DFFARX1 I_40413 (I689539,I2507,I689488,I689471,);
nor I_40414 (I689584,I171653,I171674);
and I_40415 (I689601,I689584,I171668);
nor I_40416 (I689618,I689601,I171653);
not I_40417 (I689635,I171653);
and I_40418 (I689652,I689635,I171650);
nand I_40419 (I689669,I689652,I171662);
nor I_40420 (I689686,I689635,I689669);
DFFARX1 I_40421 (I689686,I2507,I689488,I689453,);
not I_40422 (I689717,I689669);
nand I_40423 (I689734,I689539,I689717);
nand I_40424 (I689465,I689601,I689717);
DFFARX1 I_40425 (I689635,I2507,I689488,I689480,);
not I_40426 (I689779,I171677);
nor I_40427 (I689796,I689779,I171650);
nor I_40428 (I689813,I689796,I689618);
DFFARX1 I_40429 (I689813,I2507,I689488,I689477,);
not I_40430 (I689844,I689796);
DFFARX1 I_40431 (I689844,I2507,I689488,I689870,);
not I_40432 (I689878,I689870);
nor I_40433 (I689474,I689878,I689796);
nor I_40434 (I689909,I689779,I171659);
and I_40435 (I689926,I689909,I171656);
or I_40436 (I689943,I689926,I171650);
DFFARX1 I_40437 (I689943,I2507,I689488,I689969,);
not I_40438 (I689977,I689969);
nand I_40439 (I689994,I689977,I689717);
not I_40440 (I689468,I689994);
nand I_40441 (I689462,I689994,I689734);
nand I_40442 (I689459,I689977,I689601);
not I_40443 (I690083,I2514);
DFFARX1 I_40444 (I610406,I2507,I690083,I690109,);
DFFARX1 I_40445 (I610418,I2507,I690083,I690126,);
not I_40446 (I690134,I690126);
nor I_40447 (I690051,I690109,I690134);
DFFARX1 I_40448 (I690134,I2507,I690083,I690066,);
nor I_40449 (I690179,I610415,I610409);
and I_40450 (I690196,I690179,I610403);
nor I_40451 (I690213,I690196,I610415);
not I_40452 (I690230,I610415);
and I_40453 (I690247,I690230,I610412);
nand I_40454 (I690264,I690247,I610403);
nor I_40455 (I690281,I690230,I690264);
DFFARX1 I_40456 (I690281,I2507,I690083,I690048,);
not I_40457 (I690312,I690264);
nand I_40458 (I690329,I690134,I690312);
nand I_40459 (I690060,I690196,I690312);
DFFARX1 I_40460 (I690230,I2507,I690083,I690075,);
not I_40461 (I690374,I610427);
nor I_40462 (I690391,I690374,I610412);
nor I_40463 (I690408,I690391,I690213);
DFFARX1 I_40464 (I690408,I2507,I690083,I690072,);
not I_40465 (I690439,I690391);
DFFARX1 I_40466 (I690439,I2507,I690083,I690465,);
not I_40467 (I690473,I690465);
nor I_40468 (I690069,I690473,I690391);
nor I_40469 (I690504,I690374,I610421);
and I_40470 (I690521,I690504,I610424);
or I_40471 (I690538,I690521,I610406);
DFFARX1 I_40472 (I690538,I2507,I690083,I690564,);
not I_40473 (I690572,I690564);
nand I_40474 (I690589,I690572,I690312);
not I_40475 (I690063,I690589);
nand I_40476 (I690057,I690589,I690329);
nand I_40477 (I690054,I690572,I690196);
not I_40478 (I690678,I2514);
DFFARX1 I_40479 (I185373,I2507,I690678,I690704,);
DFFARX1 I_40480 (I185367,I2507,I690678,I690721,);
not I_40481 (I690729,I690721);
nor I_40482 (I690646,I690704,I690729);
DFFARX1 I_40483 (I690729,I2507,I690678,I690661,);
nor I_40484 (I690774,I185355,I185376);
and I_40485 (I690791,I690774,I185370);
nor I_40486 (I690808,I690791,I185355);
not I_40487 (I690825,I185355);
and I_40488 (I690842,I690825,I185352);
nand I_40489 (I690859,I690842,I185364);
nor I_40490 (I690876,I690825,I690859);
DFFARX1 I_40491 (I690876,I2507,I690678,I690643,);
not I_40492 (I690907,I690859);
nand I_40493 (I690924,I690729,I690907);
nand I_40494 (I690655,I690791,I690907);
DFFARX1 I_40495 (I690825,I2507,I690678,I690670,);
not I_40496 (I690969,I185379);
nor I_40497 (I690986,I690969,I185352);
nor I_40498 (I691003,I690986,I690808);
DFFARX1 I_40499 (I691003,I2507,I690678,I690667,);
not I_40500 (I691034,I690986);
DFFARX1 I_40501 (I691034,I2507,I690678,I691060,);
not I_40502 (I691068,I691060);
nor I_40503 (I690664,I691068,I690986);
nor I_40504 (I691099,I690969,I185361);
and I_40505 (I691116,I691099,I185358);
or I_40506 (I691133,I691116,I185352);
DFFARX1 I_40507 (I691133,I2507,I690678,I691159,);
not I_40508 (I691167,I691159);
nand I_40509 (I691184,I691167,I690907);
not I_40510 (I690658,I691184);
nand I_40511 (I690652,I691184,I690924);
nand I_40512 (I690649,I691167,I690791);
not I_40513 (I691273,I2514);
DFFARX1 I_40514 (I76794,I2507,I691273,I691299,);
DFFARX1 I_40515 (I76782,I2507,I691273,I691316,);
not I_40516 (I691324,I691316);
nor I_40517 (I691241,I691299,I691324);
DFFARX1 I_40518 (I691324,I2507,I691273,I691256,);
nor I_40519 (I691369,I76773,I76797);
and I_40520 (I691386,I691369,I76776);
nor I_40521 (I691403,I691386,I76773);
not I_40522 (I691420,I76773);
and I_40523 (I691437,I691420,I76779);
nand I_40524 (I691454,I691437,I76791);
nor I_40525 (I691471,I691420,I691454);
DFFARX1 I_40526 (I691471,I2507,I691273,I691238,);
not I_40527 (I691502,I691454);
nand I_40528 (I691519,I691324,I691502);
nand I_40529 (I691250,I691386,I691502);
DFFARX1 I_40530 (I691420,I2507,I691273,I691265,);
not I_40531 (I691564,I76773);
nor I_40532 (I691581,I691564,I76779);
nor I_40533 (I691598,I691581,I691403);
DFFARX1 I_40534 (I691598,I2507,I691273,I691262,);
not I_40535 (I691629,I691581);
DFFARX1 I_40536 (I691629,I2507,I691273,I691655,);
not I_40537 (I691663,I691655);
nor I_40538 (I691259,I691663,I691581);
nor I_40539 (I691694,I691564,I76776);
and I_40540 (I691711,I691694,I76785);
or I_40541 (I691728,I691711,I76788);
DFFARX1 I_40542 (I691728,I2507,I691273,I691754,);
not I_40543 (I691762,I691754);
nand I_40544 (I691779,I691762,I691502);
not I_40545 (I691253,I691779);
nand I_40546 (I691247,I691779,I691519);
nand I_40547 (I691244,I691762,I691386);
not I_40548 (I691868,I2514);
DFFARX1 I_40549 (I598268,I2507,I691868,I691894,);
DFFARX1 I_40550 (I598280,I2507,I691868,I691911,);
not I_40551 (I691919,I691911);
nor I_40552 (I691836,I691894,I691919);
DFFARX1 I_40553 (I691919,I2507,I691868,I691851,);
nor I_40554 (I691964,I598277,I598271);
and I_40555 (I691981,I691964,I598265);
nor I_40556 (I691998,I691981,I598277);
not I_40557 (I692015,I598277);
and I_40558 (I692032,I692015,I598274);
nand I_40559 (I692049,I692032,I598265);
nor I_40560 (I692066,I692015,I692049);
DFFARX1 I_40561 (I692066,I2507,I691868,I691833,);
not I_40562 (I692097,I692049);
nand I_40563 (I692114,I691919,I692097);
nand I_40564 (I691845,I691981,I692097);
DFFARX1 I_40565 (I692015,I2507,I691868,I691860,);
not I_40566 (I692159,I598289);
nor I_40567 (I692176,I692159,I598274);
nor I_40568 (I692193,I692176,I691998);
DFFARX1 I_40569 (I692193,I2507,I691868,I691857,);
not I_40570 (I692224,I692176);
DFFARX1 I_40571 (I692224,I2507,I691868,I692250,);
not I_40572 (I692258,I692250);
nor I_40573 (I691854,I692258,I692176);
nor I_40574 (I692289,I692159,I598283);
and I_40575 (I692306,I692289,I598286);
or I_40576 (I692323,I692306,I598268);
DFFARX1 I_40577 (I692323,I2507,I691868,I692349,);
not I_40578 (I692357,I692349);
nand I_40579 (I692374,I692357,I692097);
not I_40580 (I691848,I692374);
nand I_40581 (I691842,I692374,I692114);
nand I_40582 (I691839,I692357,I691981);
not I_40583 (I692463,I2514);
DFFARX1 I_40584 (I315474,I2507,I692463,I692489,);
DFFARX1 I_40585 (I315468,I2507,I692463,I692506,);
not I_40586 (I692514,I692506);
nor I_40587 (I692431,I692489,I692514);
DFFARX1 I_40588 (I692514,I2507,I692463,I692446,);
nor I_40589 (I692559,I315465,I315456);
and I_40590 (I692576,I692559,I315453);
nor I_40591 (I692593,I692576,I315465);
not I_40592 (I692610,I315465);
and I_40593 (I692627,I692610,I315459);
nand I_40594 (I692644,I692627,I315471);
nor I_40595 (I692661,I692610,I692644);
DFFARX1 I_40596 (I692661,I2507,I692463,I692428,);
not I_40597 (I692692,I692644);
nand I_40598 (I692709,I692514,I692692);
nand I_40599 (I692440,I692576,I692692);
DFFARX1 I_40600 (I692610,I2507,I692463,I692455,);
not I_40601 (I692754,I315477);
nor I_40602 (I692771,I692754,I315459);
nor I_40603 (I692788,I692771,I692593);
DFFARX1 I_40604 (I692788,I2507,I692463,I692452,);
not I_40605 (I692819,I692771);
DFFARX1 I_40606 (I692819,I2507,I692463,I692845,);
not I_40607 (I692853,I692845);
nor I_40608 (I692449,I692853,I692771);
nor I_40609 (I692884,I692754,I315456);
and I_40610 (I692901,I692884,I315462);
or I_40611 (I692918,I692901,I315453);
DFFARX1 I_40612 (I692918,I2507,I692463,I692944,);
not I_40613 (I692952,I692944);
nand I_40614 (I692969,I692952,I692692);
not I_40615 (I692443,I692969);
nand I_40616 (I692437,I692969,I692709);
nand I_40617 (I692434,I692952,I692576);
not I_40618 (I693058,I2514);
DFFARX1 I_40619 (I558752,I2507,I693058,I693084,);
DFFARX1 I_40620 (I558743,I2507,I693058,I693101,);
not I_40621 (I693109,I693101);
nor I_40622 (I693026,I693084,I693109);
DFFARX1 I_40623 (I693109,I2507,I693058,I693041,);
nor I_40624 (I693154,I558749,I558758);
and I_40625 (I693171,I693154,I558761);
nor I_40626 (I693188,I693171,I558749);
not I_40627 (I693205,I558749);
and I_40628 (I693222,I693205,I558740);
nand I_40629 (I693239,I693222,I558746);
nor I_40630 (I693256,I693205,I693239);
DFFARX1 I_40631 (I693256,I2507,I693058,I693023,);
not I_40632 (I693287,I693239);
nand I_40633 (I693304,I693109,I693287);
nand I_40634 (I693035,I693171,I693287);
DFFARX1 I_40635 (I693205,I2507,I693058,I693050,);
not I_40636 (I693349,I558755);
nor I_40637 (I693366,I693349,I558740);
nor I_40638 (I693383,I693366,I693188);
DFFARX1 I_40639 (I693383,I2507,I693058,I693047,);
not I_40640 (I693414,I693366);
DFFARX1 I_40641 (I693414,I2507,I693058,I693440,);
not I_40642 (I693448,I693440);
nor I_40643 (I693044,I693448,I693366);
nor I_40644 (I693479,I693349,I558740);
and I_40645 (I693496,I693479,I558743);
or I_40646 (I693513,I693496,I558746);
DFFARX1 I_40647 (I693513,I2507,I693058,I693539,);
not I_40648 (I693547,I693539);
nand I_40649 (I693564,I693547,I693287);
not I_40650 (I693038,I693564);
nand I_40651 (I693032,I693564,I693304);
nand I_40652 (I693029,I693547,I693171);
not I_40653 (I693653,I2514);
DFFARX1 I_40654 (I374430,I2507,I693653,I693679,);
DFFARX1 I_40655 (I374412,I2507,I693653,I693696,);
not I_40656 (I693704,I693696);
nor I_40657 (I693621,I693679,I693704);
DFFARX1 I_40658 (I693704,I2507,I693653,I693636,);
nor I_40659 (I693749,I374418,I374421);
and I_40660 (I693766,I693749,I374409);
nor I_40661 (I693783,I693766,I374418);
not I_40662 (I693800,I374418);
and I_40663 (I693817,I693800,I374427);
nand I_40664 (I693834,I693817,I374415);
nor I_40665 (I693851,I693800,I693834);
DFFARX1 I_40666 (I693851,I2507,I693653,I693618,);
not I_40667 (I693882,I693834);
nand I_40668 (I693899,I693704,I693882);
nand I_40669 (I693630,I693766,I693882);
DFFARX1 I_40670 (I693800,I2507,I693653,I693645,);
not I_40671 (I693944,I374412);
nor I_40672 (I693961,I693944,I374427);
nor I_40673 (I693978,I693961,I693783);
DFFARX1 I_40674 (I693978,I2507,I693653,I693642,);
not I_40675 (I694009,I693961);
DFFARX1 I_40676 (I694009,I2507,I693653,I694035,);
not I_40677 (I694043,I694035);
nor I_40678 (I693639,I694043,I693961);
nor I_40679 (I694074,I693944,I374424);
and I_40680 (I694091,I694074,I374433);
or I_40681 (I694108,I694091,I374409);
DFFARX1 I_40682 (I694108,I2507,I693653,I694134,);
not I_40683 (I694142,I694134);
nand I_40684 (I694159,I694142,I693882);
not I_40685 (I693633,I694159);
nand I_40686 (I693627,I694159,I693899);
nand I_40687 (I693624,I694142,I693766);
not I_40688 (I694248,I2514);
DFFARX1 I_40689 (I156809,I2507,I694248,I694274,);
DFFARX1 I_40690 (I156812,I2507,I694248,I694291,);
not I_40691 (I694299,I694291);
nor I_40692 (I694216,I694274,I694299);
DFFARX1 I_40693 (I694299,I2507,I694248,I694231,);
nor I_40694 (I694344,I156818,I156812);
and I_40695 (I694361,I694344,I156815);
nor I_40696 (I694378,I694361,I156818);
not I_40697 (I694395,I156818);
and I_40698 (I694412,I694395,I156809);
nand I_40699 (I694429,I694412,I156827);
nor I_40700 (I694446,I694395,I694429);
DFFARX1 I_40701 (I694446,I2507,I694248,I694213,);
not I_40702 (I694477,I694429);
nand I_40703 (I694494,I694299,I694477);
nand I_40704 (I694225,I694361,I694477);
DFFARX1 I_40705 (I694395,I2507,I694248,I694240,);
not I_40706 (I694539,I156821);
nor I_40707 (I694556,I694539,I156809);
nor I_40708 (I694573,I694556,I694378);
DFFARX1 I_40709 (I694573,I2507,I694248,I694237,);
not I_40710 (I694604,I694556);
DFFARX1 I_40711 (I694604,I2507,I694248,I694630,);
not I_40712 (I694638,I694630);
nor I_40713 (I694234,I694638,I694556);
nor I_40714 (I694669,I694539,I156824);
and I_40715 (I694686,I694669,I156830);
or I_40716 (I694703,I694686,I156833);
DFFARX1 I_40717 (I694703,I2507,I694248,I694729,);
not I_40718 (I694737,I694729);
nand I_40719 (I694754,I694737,I694477);
not I_40720 (I694228,I694754);
nand I_40721 (I694222,I694754,I694494);
nand I_40722 (I694219,I694737,I694361);
not I_40723 (I694843,I2514);
DFFARX1 I_40724 (I271032,I2507,I694843,I694869,);
DFFARX1 I_40725 (I271038,I2507,I694843,I694886,);
not I_40726 (I694894,I694886);
nor I_40727 (I694811,I694869,I694894);
DFFARX1 I_40728 (I694894,I2507,I694843,I694826,);
nor I_40729 (I694939,I271047,I271032);
and I_40730 (I694956,I694939,I271059);
nor I_40731 (I694973,I694956,I271047);
not I_40732 (I694990,I271047);
and I_40733 (I695007,I694990,I271035);
nand I_40734 (I695024,I695007,I271056);
nor I_40735 (I695041,I694990,I695024);
DFFARX1 I_40736 (I695041,I2507,I694843,I694808,);
not I_40737 (I695072,I695024);
nand I_40738 (I695089,I694894,I695072);
nand I_40739 (I694820,I694956,I695072);
DFFARX1 I_40740 (I694990,I2507,I694843,I694835,);
not I_40741 (I695134,I271044);
nor I_40742 (I695151,I695134,I271035);
nor I_40743 (I695168,I695151,I694973);
DFFARX1 I_40744 (I695168,I2507,I694843,I694832,);
not I_40745 (I695199,I695151);
DFFARX1 I_40746 (I695199,I2507,I694843,I695225,);
not I_40747 (I695233,I695225);
nor I_40748 (I694829,I695233,I695151);
nor I_40749 (I695264,I695134,I271041);
and I_40750 (I695281,I695264,I271053);
or I_40751 (I695298,I695281,I271050);
DFFARX1 I_40752 (I695298,I2507,I694843,I695324,);
not I_40753 (I695332,I695324);
nand I_40754 (I695349,I695332,I695072);
not I_40755 (I694823,I695349);
nand I_40756 (I694817,I695349,I695089);
nand I_40757 (I694814,I695332,I694956);
not I_40758 (I695438,I2514);
DFFARX1 I_40759 (I344952,I2507,I695438,I695464,);
DFFARX1 I_40760 (I344946,I2507,I695438,I695481,);
not I_40761 (I695489,I695481);
nor I_40762 (I695406,I695464,I695489);
DFFARX1 I_40763 (I695489,I2507,I695438,I695421,);
nor I_40764 (I695534,I344943,I344934);
and I_40765 (I695551,I695534,I344931);
nor I_40766 (I695568,I695551,I344943);
not I_40767 (I695585,I344943);
and I_40768 (I695602,I695585,I344937);
nand I_40769 (I695619,I695602,I344949);
nor I_40770 (I695636,I695585,I695619);
DFFARX1 I_40771 (I695636,I2507,I695438,I695403,);
not I_40772 (I695667,I695619);
nand I_40773 (I695684,I695489,I695667);
nand I_40774 (I695415,I695551,I695667);
DFFARX1 I_40775 (I695585,I2507,I695438,I695430,);
not I_40776 (I695729,I344955);
nor I_40777 (I695746,I695729,I344937);
nor I_40778 (I695763,I695746,I695568);
DFFARX1 I_40779 (I695763,I2507,I695438,I695427,);
not I_40780 (I695794,I695746);
DFFARX1 I_40781 (I695794,I2507,I695438,I695820,);
not I_40782 (I695828,I695820);
nor I_40783 (I695424,I695828,I695746);
nor I_40784 (I695859,I695729,I344934);
and I_40785 (I695876,I695859,I344940);
or I_40786 (I695893,I695876,I344931);
DFFARX1 I_40787 (I695893,I2507,I695438,I695919,);
not I_40788 (I695927,I695919);
nand I_40789 (I695944,I695927,I695667);
not I_40790 (I695418,I695944);
nand I_40791 (I695412,I695944,I695684);
nand I_40792 (I695409,I695927,I695551);
not I_40793 (I696033,I2514);
DFFARX1 I_40794 (I591332,I2507,I696033,I696059,);
DFFARX1 I_40795 (I591344,I2507,I696033,I696076,);
not I_40796 (I696084,I696076);
nor I_40797 (I696001,I696059,I696084);
DFFARX1 I_40798 (I696084,I2507,I696033,I696016,);
nor I_40799 (I696129,I591341,I591335);
and I_40800 (I696146,I696129,I591329);
nor I_40801 (I696163,I696146,I591341);
not I_40802 (I696180,I591341);
and I_40803 (I696197,I696180,I591338);
nand I_40804 (I696214,I696197,I591329);
nor I_40805 (I696231,I696180,I696214);
DFFARX1 I_40806 (I696231,I2507,I696033,I695998,);
not I_40807 (I696262,I696214);
nand I_40808 (I696279,I696084,I696262);
nand I_40809 (I696010,I696146,I696262);
DFFARX1 I_40810 (I696180,I2507,I696033,I696025,);
not I_40811 (I696324,I591353);
nor I_40812 (I696341,I696324,I591338);
nor I_40813 (I696358,I696341,I696163);
DFFARX1 I_40814 (I696358,I2507,I696033,I696022,);
not I_40815 (I696389,I696341);
DFFARX1 I_40816 (I696389,I2507,I696033,I696415,);
not I_40817 (I696423,I696415);
nor I_40818 (I696019,I696423,I696341);
nor I_40819 (I696454,I696324,I591347);
and I_40820 (I696471,I696454,I591350);
or I_40821 (I696488,I696471,I591332);
DFFARX1 I_40822 (I696488,I2507,I696033,I696514,);
not I_40823 (I696522,I696514);
nand I_40824 (I696539,I696522,I696262);
not I_40825 (I696013,I696539);
nand I_40826 (I696007,I696539,I696279);
nand I_40827 (I696004,I696522,I696146);
not I_40828 (I696628,I2514);
DFFARX1 I_40829 (I142529,I2507,I696628,I696654,);
DFFARX1 I_40830 (I142532,I2507,I696628,I696671,);
not I_40831 (I696679,I696671);
nor I_40832 (I696596,I696654,I696679);
DFFARX1 I_40833 (I696679,I2507,I696628,I696611,);
nor I_40834 (I696724,I142538,I142532);
and I_40835 (I696741,I696724,I142535);
nor I_40836 (I696758,I696741,I142538);
not I_40837 (I696775,I142538);
and I_40838 (I696792,I696775,I142529);
nand I_40839 (I696809,I696792,I142547);
nor I_40840 (I696826,I696775,I696809);
DFFARX1 I_40841 (I696826,I2507,I696628,I696593,);
not I_40842 (I696857,I696809);
nand I_40843 (I696874,I696679,I696857);
nand I_40844 (I696605,I696741,I696857);
DFFARX1 I_40845 (I696775,I2507,I696628,I696620,);
not I_40846 (I696919,I142541);
nor I_40847 (I696936,I696919,I142529);
nor I_40848 (I696953,I696936,I696758);
DFFARX1 I_40849 (I696953,I2507,I696628,I696617,);
not I_40850 (I696984,I696936);
DFFARX1 I_40851 (I696984,I2507,I696628,I697010,);
not I_40852 (I697018,I697010);
nor I_40853 (I696614,I697018,I696936);
nor I_40854 (I697049,I696919,I142544);
and I_40855 (I697066,I697049,I142550);
or I_40856 (I697083,I697066,I142553);
DFFARX1 I_40857 (I697083,I2507,I696628,I697109,);
not I_40858 (I697117,I697109);
nand I_40859 (I697134,I697117,I696857);
not I_40860 (I696608,I697134);
nand I_40861 (I696602,I697134,I696874);
nand I_40862 (I696599,I697117,I696741);
not I_40863 (I697223,I2514);
DFFARX1 I_40864 (I113969,I2507,I697223,I697249,);
DFFARX1 I_40865 (I113972,I2507,I697223,I697266,);
not I_40866 (I697274,I697266);
nor I_40867 (I697191,I697249,I697274);
DFFARX1 I_40868 (I697274,I2507,I697223,I697206,);
nor I_40869 (I697319,I113978,I113972);
and I_40870 (I697336,I697319,I113975);
nor I_40871 (I697353,I697336,I113978);
not I_40872 (I697370,I113978);
and I_40873 (I697387,I697370,I113969);
nand I_40874 (I697404,I697387,I113987);
nor I_40875 (I697421,I697370,I697404);
DFFARX1 I_40876 (I697421,I2507,I697223,I697188,);
not I_40877 (I697452,I697404);
nand I_40878 (I697469,I697274,I697452);
nand I_40879 (I697200,I697336,I697452);
DFFARX1 I_40880 (I697370,I2507,I697223,I697215,);
not I_40881 (I697514,I113981);
nor I_40882 (I697531,I697514,I113969);
nor I_40883 (I697548,I697531,I697353);
DFFARX1 I_40884 (I697548,I2507,I697223,I697212,);
not I_40885 (I697579,I697531);
DFFARX1 I_40886 (I697579,I2507,I697223,I697605,);
not I_40887 (I697613,I697605);
nor I_40888 (I697209,I697613,I697531);
nor I_40889 (I697644,I697514,I113984);
and I_40890 (I697661,I697644,I113990);
or I_40891 (I697678,I697661,I113993);
DFFARX1 I_40892 (I697678,I2507,I697223,I697704,);
not I_40893 (I697712,I697704);
nand I_40894 (I697729,I697712,I697452);
not I_40895 (I697203,I697729);
nand I_40896 (I697197,I697729,I697469);
nand I_40897 (I697194,I697712,I697336);
not I_40898 (I697818,I2514);
DFFARX1 I_40899 (I192751,I2507,I697818,I697844,);
DFFARX1 I_40900 (I192745,I2507,I697818,I697861,);
not I_40901 (I697869,I697861);
nor I_40902 (I697786,I697844,I697869);
DFFARX1 I_40903 (I697869,I2507,I697818,I697801,);
nor I_40904 (I697914,I192733,I192754);
and I_40905 (I697931,I697914,I192748);
nor I_40906 (I697948,I697931,I192733);
not I_40907 (I697965,I192733);
and I_40908 (I697982,I697965,I192730);
nand I_40909 (I697999,I697982,I192742);
nor I_40910 (I698016,I697965,I697999);
DFFARX1 I_40911 (I698016,I2507,I697818,I697783,);
not I_40912 (I698047,I697999);
nand I_40913 (I698064,I697869,I698047);
nand I_40914 (I697795,I697931,I698047);
DFFARX1 I_40915 (I697965,I2507,I697818,I697810,);
not I_40916 (I698109,I192757);
nor I_40917 (I698126,I698109,I192730);
nor I_40918 (I698143,I698126,I697948);
DFFARX1 I_40919 (I698143,I2507,I697818,I697807,);
not I_40920 (I698174,I698126);
DFFARX1 I_40921 (I698174,I2507,I697818,I698200,);
not I_40922 (I698208,I698200);
nor I_40923 (I697804,I698208,I698126);
nor I_40924 (I698239,I698109,I192739);
and I_40925 (I698256,I698239,I192736);
or I_40926 (I698273,I698256,I192730);
DFFARX1 I_40927 (I698273,I2507,I697818,I698299,);
not I_40928 (I698307,I698299);
nand I_40929 (I698324,I698307,I698047);
not I_40930 (I697798,I698324);
nand I_40931 (I697792,I698324,I698064);
nand I_40932 (I697789,I698307,I697931);
not I_40933 (I698413,I2514);
DFFARX1 I_40934 (I361136,I2507,I698413,I698439,);
DFFARX1 I_40935 (I361118,I2507,I698413,I698456,);
not I_40936 (I698464,I698456);
nor I_40937 (I698381,I698439,I698464);
DFFARX1 I_40938 (I698464,I2507,I698413,I698396,);
nor I_40939 (I698509,I361124,I361127);
and I_40940 (I698526,I698509,I361115);
nor I_40941 (I698543,I698526,I361124);
not I_40942 (I698560,I361124);
and I_40943 (I698577,I698560,I361133);
nand I_40944 (I698594,I698577,I361121);
nor I_40945 (I698611,I698560,I698594);
DFFARX1 I_40946 (I698611,I2507,I698413,I698378,);
not I_40947 (I698642,I698594);
nand I_40948 (I698659,I698464,I698642);
nand I_40949 (I698390,I698526,I698642);
DFFARX1 I_40950 (I698560,I2507,I698413,I698405,);
not I_40951 (I698704,I361118);
nor I_40952 (I698721,I698704,I361133);
nor I_40953 (I698738,I698721,I698543);
DFFARX1 I_40954 (I698738,I2507,I698413,I698402,);
not I_40955 (I698769,I698721);
DFFARX1 I_40956 (I698769,I2507,I698413,I698795,);
not I_40957 (I698803,I698795);
nor I_40958 (I698399,I698803,I698721);
nor I_40959 (I698834,I698704,I361130);
and I_40960 (I698851,I698834,I361139);
or I_40961 (I698868,I698851,I361115);
DFFARX1 I_40962 (I698868,I2507,I698413,I698894,);
not I_40963 (I698902,I698894);
nand I_40964 (I698919,I698902,I698642);
not I_40965 (I698393,I698919);
nand I_40966 (I698387,I698919,I698659);
nand I_40967 (I698384,I698902,I698526);
not I_40968 (I699008,I2514);
DFFARX1 I_40969 (I232408,I2507,I699008,I699034,);
DFFARX1 I_40970 (I232414,I2507,I699008,I699051,);
not I_40971 (I699059,I699051);
nor I_40972 (I698976,I699034,I699059);
DFFARX1 I_40973 (I699059,I2507,I699008,I698991,);
nor I_40974 (I699104,I232423,I232408);
and I_40975 (I699121,I699104,I232435);
nor I_40976 (I699138,I699121,I232423);
not I_40977 (I699155,I232423);
and I_40978 (I699172,I699155,I232411);
nand I_40979 (I699189,I699172,I232432);
nor I_40980 (I699206,I699155,I699189);
DFFARX1 I_40981 (I699206,I2507,I699008,I698973,);
not I_40982 (I699237,I699189);
nand I_40983 (I699254,I699059,I699237);
nand I_40984 (I698985,I699121,I699237);
DFFARX1 I_40985 (I699155,I2507,I699008,I699000,);
not I_40986 (I699299,I232420);
nor I_40987 (I699316,I699299,I232411);
nor I_40988 (I699333,I699316,I699138);
DFFARX1 I_40989 (I699333,I2507,I699008,I698997,);
not I_40990 (I699364,I699316);
DFFARX1 I_40991 (I699364,I2507,I699008,I699390,);
not I_40992 (I699398,I699390);
nor I_40993 (I698994,I699398,I699316);
nor I_40994 (I699429,I699299,I232417);
and I_40995 (I699446,I699429,I232429);
or I_40996 (I699463,I699446,I232426);
DFFARX1 I_40997 (I699463,I2507,I699008,I699489,);
not I_40998 (I699497,I699489);
nand I_40999 (I699514,I699497,I699237);
not I_41000 (I698988,I699514);
nand I_41001 (I698982,I699514,I699254);
nand I_41002 (I698979,I699497,I699121);
not I_41003 (I699603,I2514);
DFFARX1 I_41004 (I625434,I2507,I699603,I699629,);
DFFARX1 I_41005 (I625446,I2507,I699603,I699646,);
not I_41006 (I699654,I699646);
nor I_41007 (I699571,I699629,I699654);
DFFARX1 I_41008 (I699654,I2507,I699603,I699586,);
nor I_41009 (I699699,I625443,I625437);
and I_41010 (I699716,I699699,I625431);
nor I_41011 (I699733,I699716,I625443);
not I_41012 (I699750,I625443);
and I_41013 (I699767,I699750,I625440);
nand I_41014 (I699784,I699767,I625431);
nor I_41015 (I699801,I699750,I699784);
DFFARX1 I_41016 (I699801,I2507,I699603,I699568,);
not I_41017 (I699832,I699784);
nand I_41018 (I699849,I699654,I699832);
nand I_41019 (I699580,I699716,I699832);
DFFARX1 I_41020 (I699750,I2507,I699603,I699595,);
not I_41021 (I699894,I625455);
nor I_41022 (I699911,I699894,I625440);
nor I_41023 (I699928,I699911,I699733);
DFFARX1 I_41024 (I699928,I2507,I699603,I699592,);
not I_41025 (I699959,I699911);
DFFARX1 I_41026 (I699959,I2507,I699603,I699985,);
not I_41027 (I699993,I699985);
nor I_41028 (I699589,I699993,I699911);
nor I_41029 (I700024,I699894,I625449);
and I_41030 (I700041,I700024,I625452);
or I_41031 (I700058,I700041,I625434);
DFFARX1 I_41032 (I700058,I2507,I699603,I700084,);
not I_41033 (I700092,I700084);
nand I_41034 (I700109,I700092,I699832);
not I_41035 (I699583,I700109);
nand I_41036 (I699577,I700109,I699849);
nand I_41037 (I699574,I700092,I699716);
not I_41038 (I700198,I2514);
DFFARX1 I_41039 (I560996,I2507,I700198,I700224,);
DFFARX1 I_41040 (I560987,I2507,I700198,I700241,);
not I_41041 (I700249,I700241);
nor I_41042 (I700166,I700224,I700249);
DFFARX1 I_41043 (I700249,I2507,I700198,I700181,);
nor I_41044 (I700294,I560993,I561002);
and I_41045 (I700311,I700294,I561005);
nor I_41046 (I700328,I700311,I560993);
not I_41047 (I700345,I560993);
and I_41048 (I700362,I700345,I560984);
nand I_41049 (I700379,I700362,I560990);
nor I_41050 (I700396,I700345,I700379);
DFFARX1 I_41051 (I700396,I2507,I700198,I700163,);
not I_41052 (I700427,I700379);
nand I_41053 (I700444,I700249,I700427);
nand I_41054 (I700175,I700311,I700427);
DFFARX1 I_41055 (I700345,I2507,I700198,I700190,);
not I_41056 (I700489,I560999);
nor I_41057 (I700506,I700489,I560984);
nor I_41058 (I700523,I700506,I700328);
DFFARX1 I_41059 (I700523,I2507,I700198,I700187,);
not I_41060 (I700554,I700506);
DFFARX1 I_41061 (I700554,I2507,I700198,I700580,);
not I_41062 (I700588,I700580);
nor I_41063 (I700184,I700588,I700506);
nor I_41064 (I700619,I700489,I560984);
and I_41065 (I700636,I700619,I560987);
or I_41066 (I700653,I700636,I560990);
DFFARX1 I_41067 (I700653,I2507,I700198,I700679,);
not I_41068 (I700687,I700679);
nand I_41069 (I700704,I700687,I700427);
not I_41070 (I700178,I700704);
nand I_41071 (I700172,I700704,I700444);
nand I_41072 (I700169,I700687,I700311);
not I_41073 (I700793,I2514);
DFFARX1 I_41074 (I434445,I2507,I700793,I700819,);
DFFARX1 I_41075 (I434442,I2507,I700793,I700836,);
not I_41076 (I700844,I700836);
nor I_41077 (I700761,I700819,I700844);
DFFARX1 I_41078 (I700844,I2507,I700793,I700776,);
nor I_41079 (I700889,I434457,I434439);
and I_41080 (I700906,I700889,I434436);
nor I_41081 (I700923,I700906,I434457);
not I_41082 (I700940,I434457);
and I_41083 (I700957,I700940,I434442);
nand I_41084 (I700974,I700957,I434454);
nor I_41085 (I700991,I700940,I700974);
DFFARX1 I_41086 (I700991,I2507,I700793,I700758,);
not I_41087 (I701022,I700974);
nand I_41088 (I701039,I700844,I701022);
nand I_41089 (I700770,I700906,I701022);
DFFARX1 I_41090 (I700940,I2507,I700793,I700785,);
not I_41091 (I701084,I434448);
nor I_41092 (I701101,I701084,I434442);
nor I_41093 (I701118,I701101,I700923);
DFFARX1 I_41094 (I701118,I2507,I700793,I700782,);
not I_41095 (I701149,I701101);
DFFARX1 I_41096 (I701149,I2507,I700793,I701175,);
not I_41097 (I701183,I701175);
nor I_41098 (I700779,I701183,I701101);
nor I_41099 (I701214,I701084,I434436);
and I_41100 (I701231,I701214,I434451);
or I_41101 (I701248,I701231,I434439);
DFFARX1 I_41102 (I701248,I2507,I700793,I701274,);
not I_41103 (I701282,I701274);
nand I_41104 (I701299,I701282,I701022);
not I_41105 (I700773,I701299);
nand I_41106 (I700767,I701299,I701039);
nand I_41107 (I700764,I701282,I700906);
not I_41108 (I701388,I2514);
DFFARX1 I_41109 (I73105,I2507,I701388,I701414,);
DFFARX1 I_41110 (I73093,I2507,I701388,I701431,);
not I_41111 (I701439,I701431);
nor I_41112 (I701356,I701414,I701439);
DFFARX1 I_41113 (I701439,I2507,I701388,I701371,);
nor I_41114 (I701484,I73084,I73108);
and I_41115 (I701501,I701484,I73087);
nor I_41116 (I701518,I701501,I73084);
not I_41117 (I701535,I73084);
and I_41118 (I701552,I701535,I73090);
nand I_41119 (I701569,I701552,I73102);
nor I_41120 (I701586,I701535,I701569);
DFFARX1 I_41121 (I701586,I2507,I701388,I701353,);
not I_41122 (I701617,I701569);
nand I_41123 (I701634,I701439,I701617);
nand I_41124 (I701365,I701501,I701617);
DFFARX1 I_41125 (I701535,I2507,I701388,I701380,);
not I_41126 (I701679,I73084);
nor I_41127 (I701696,I701679,I73090);
nor I_41128 (I701713,I701696,I701518);
DFFARX1 I_41129 (I701713,I2507,I701388,I701377,);
not I_41130 (I701744,I701696);
DFFARX1 I_41131 (I701744,I2507,I701388,I701770,);
not I_41132 (I701778,I701770);
nor I_41133 (I701374,I701778,I701696);
nor I_41134 (I701809,I701679,I73087);
and I_41135 (I701826,I701809,I73096);
or I_41136 (I701843,I701826,I73099);
DFFARX1 I_41137 (I701843,I2507,I701388,I701869,);
not I_41138 (I701877,I701869);
nand I_41139 (I701894,I701877,I701617);
not I_41140 (I701368,I701894);
nand I_41141 (I701362,I701894,I701634);
nand I_41142 (I701359,I701877,I701501);
not I_41143 (I701983,I2514);
DFFARX1 I_41144 (I317786,I2507,I701983,I702009,);
DFFARX1 I_41145 (I317780,I2507,I701983,I702026,);
not I_41146 (I702034,I702026);
nor I_41147 (I701951,I702009,I702034);
DFFARX1 I_41148 (I702034,I2507,I701983,I701966,);
nor I_41149 (I702079,I317777,I317768);
and I_41150 (I702096,I702079,I317765);
nor I_41151 (I702113,I702096,I317777);
not I_41152 (I702130,I317777);
and I_41153 (I702147,I702130,I317771);
nand I_41154 (I702164,I702147,I317783);
nor I_41155 (I702181,I702130,I702164);
DFFARX1 I_41156 (I702181,I2507,I701983,I701948,);
not I_41157 (I702212,I702164);
nand I_41158 (I702229,I702034,I702212);
nand I_41159 (I701960,I702096,I702212);
DFFARX1 I_41160 (I702130,I2507,I701983,I701975,);
not I_41161 (I702274,I317789);
nor I_41162 (I702291,I702274,I317771);
nor I_41163 (I702308,I702291,I702113);
DFFARX1 I_41164 (I702308,I2507,I701983,I701972,);
not I_41165 (I702339,I702291);
DFFARX1 I_41166 (I702339,I2507,I701983,I702365,);
not I_41167 (I702373,I702365);
nor I_41168 (I701969,I702373,I702291);
nor I_41169 (I702404,I702274,I317768);
and I_41170 (I702421,I702404,I317774);
or I_41171 (I702438,I702421,I317765);
DFFARX1 I_41172 (I702438,I2507,I701983,I702464,);
not I_41173 (I702472,I702464);
nand I_41174 (I702489,I702472,I702212);
not I_41175 (I701963,I702489);
nand I_41176 (I701957,I702489,I702229);
nand I_41177 (I701954,I702472,I702096);
not I_41178 (I702578,I2514);
DFFARX1 I_41179 (I106829,I2507,I702578,I702604,);
DFFARX1 I_41180 (I106832,I2507,I702578,I702621,);
not I_41181 (I702629,I702621);
nor I_41182 (I702546,I702604,I702629);
DFFARX1 I_41183 (I702629,I2507,I702578,I702561,);
nor I_41184 (I702674,I106838,I106832);
and I_41185 (I702691,I702674,I106835);
nor I_41186 (I702708,I702691,I106838);
not I_41187 (I702725,I106838);
and I_41188 (I702742,I702725,I106829);
nand I_41189 (I702759,I702742,I106847);
nor I_41190 (I702776,I702725,I702759);
DFFARX1 I_41191 (I702776,I2507,I702578,I702543,);
not I_41192 (I702807,I702759);
nand I_41193 (I702824,I702629,I702807);
nand I_41194 (I702555,I702691,I702807);
DFFARX1 I_41195 (I702725,I2507,I702578,I702570,);
not I_41196 (I702869,I106841);
nor I_41197 (I702886,I702869,I106829);
nor I_41198 (I702903,I702886,I702708);
DFFARX1 I_41199 (I702903,I2507,I702578,I702567,);
not I_41200 (I702934,I702886);
DFFARX1 I_41201 (I702934,I2507,I702578,I702960,);
not I_41202 (I702968,I702960);
nor I_41203 (I702564,I702968,I702886);
nor I_41204 (I702999,I702869,I106844);
and I_41205 (I703016,I702999,I106850);
or I_41206 (I703033,I703016,I106853);
DFFARX1 I_41207 (I703033,I2507,I702578,I703059,);
not I_41208 (I703067,I703059);
nand I_41209 (I703084,I703067,I702807);
not I_41210 (I702558,I703084);
nand I_41211 (I702552,I703084,I702824);
nand I_41212 (I702549,I703067,I702691);
not I_41213 (I703173,I2514);
DFFARX1 I_41214 (I663749,I2507,I703173,I703199,);
DFFARX1 I_41215 (I663752,I2507,I703173,I703216,);
not I_41216 (I703224,I703216);
nor I_41217 (I703141,I703199,I703224);
DFFARX1 I_41218 (I703224,I2507,I703173,I703156,);
nor I_41219 (I703269,I663752,I663767);
and I_41220 (I703286,I703269,I663761);
nor I_41221 (I703303,I703286,I663752);
not I_41222 (I703320,I663752);
and I_41223 (I703337,I703320,I663770);
nand I_41224 (I703354,I703337,I663758);
nor I_41225 (I703371,I703320,I703354);
DFFARX1 I_41226 (I703371,I2507,I703173,I703138,);
not I_41227 (I703402,I703354);
nand I_41228 (I703419,I703224,I703402);
nand I_41229 (I703150,I703286,I703402);
DFFARX1 I_41230 (I703320,I2507,I703173,I703165,);
not I_41231 (I703464,I663764);
nor I_41232 (I703481,I703464,I663770);
nor I_41233 (I703498,I703481,I703303);
DFFARX1 I_41234 (I703498,I2507,I703173,I703162,);
not I_41235 (I703529,I703481);
DFFARX1 I_41236 (I703529,I2507,I703173,I703555,);
not I_41237 (I703563,I703555);
nor I_41238 (I703159,I703563,I703481);
nor I_41239 (I703594,I703464,I663749);
and I_41240 (I703611,I703594,I663773);
or I_41241 (I703628,I703611,I663755);
DFFARX1 I_41242 (I703628,I2507,I703173,I703654,);
not I_41243 (I703662,I703654);
nand I_41244 (I703679,I703662,I703402);
not I_41245 (I703153,I703679);
nand I_41246 (I703147,I703679,I703419);
nand I_41247 (I703144,I703662,I703286);
not I_41248 (I703768,I2514);
DFFARX1 I_41249 (I583240,I2507,I703768,I703794,);
DFFARX1 I_41250 (I583252,I2507,I703768,I703811,);
not I_41251 (I703819,I703811);
nor I_41252 (I703736,I703794,I703819);
DFFARX1 I_41253 (I703819,I2507,I703768,I703751,);
nor I_41254 (I703864,I583249,I583243);
and I_41255 (I703881,I703864,I583237);
nor I_41256 (I703898,I703881,I583249);
not I_41257 (I703915,I583249);
and I_41258 (I703932,I703915,I583246);
nand I_41259 (I703949,I703932,I583237);
nor I_41260 (I703966,I703915,I703949);
DFFARX1 I_41261 (I703966,I2507,I703768,I703733,);
not I_41262 (I703997,I703949);
nand I_41263 (I704014,I703819,I703997);
nand I_41264 (I703745,I703881,I703997);
DFFARX1 I_41265 (I703915,I2507,I703768,I703760,);
not I_41266 (I704059,I583261);
nor I_41267 (I704076,I704059,I583246);
nor I_41268 (I704093,I704076,I703898);
DFFARX1 I_41269 (I704093,I2507,I703768,I703757,);
not I_41270 (I704124,I704076);
DFFARX1 I_41271 (I704124,I2507,I703768,I704150,);
not I_41272 (I704158,I704150);
nor I_41273 (I703754,I704158,I704076);
nor I_41274 (I704189,I704059,I583255);
and I_41275 (I704206,I704189,I583258);
or I_41276 (I704223,I704206,I583240);
DFFARX1 I_41277 (I704223,I2507,I703768,I704249,);
not I_41278 (I704257,I704249);
nand I_41279 (I704274,I704257,I703997);
not I_41280 (I703748,I704274);
nand I_41281 (I703742,I704274,I704014);
nand I_41282 (I703739,I704257,I703881);
not I_41283 (I704363,I2514);
DFFARX1 I_41284 (I683870,I2507,I704363,I704389,);
DFFARX1 I_41285 (I683855,I2507,I704363,I704406,);
not I_41286 (I704414,I704406);
nor I_41287 (I704331,I704389,I704414);
DFFARX1 I_41288 (I704414,I2507,I704363,I704346,);
nor I_41289 (I704459,I683852,I683861);
and I_41290 (I704476,I704459,I683867);
nor I_41291 (I704493,I704476,I683852);
not I_41292 (I704510,I683852);
and I_41293 (I704527,I704510,I683849);
nand I_41294 (I704544,I704527,I683843);
nor I_41295 (I704561,I704510,I704544);
DFFARX1 I_41296 (I704561,I2507,I704363,I704328,);
not I_41297 (I704592,I704544);
nand I_41298 (I704609,I704414,I704592);
nand I_41299 (I704340,I704476,I704592);
DFFARX1 I_41300 (I704510,I2507,I704363,I704355,);
not I_41301 (I704654,I683843);
nor I_41302 (I704671,I704654,I683849);
nor I_41303 (I704688,I704671,I704493);
DFFARX1 I_41304 (I704688,I2507,I704363,I704352,);
not I_41305 (I704719,I704671);
DFFARX1 I_41306 (I704719,I2507,I704363,I704745,);
not I_41307 (I704753,I704745);
nor I_41308 (I704349,I704753,I704671);
nor I_41309 (I704784,I704654,I683858);
and I_41310 (I704801,I704784,I683864);
or I_41311 (I704818,I704801,I683846);
DFFARX1 I_41312 (I704818,I2507,I704363,I704844,);
not I_41313 (I704852,I704844);
nand I_41314 (I704869,I704852,I704592);
not I_41315 (I704343,I704869);
nand I_41316 (I704337,I704869,I704609);
nand I_41317 (I704334,I704852,I704476);
not I_41318 (I704958,I2514);
DFFARX1 I_41319 (I280280,I2507,I704958,I704984,);
DFFARX1 I_41320 (I280286,I2507,I704958,I705001,);
not I_41321 (I705009,I705001);
nor I_41322 (I704926,I704984,I705009);
DFFARX1 I_41323 (I705009,I2507,I704958,I704941,);
nor I_41324 (I705054,I280295,I280280);
and I_41325 (I705071,I705054,I280307);
nor I_41326 (I705088,I705071,I280295);
not I_41327 (I705105,I280295);
and I_41328 (I705122,I705105,I280283);
nand I_41329 (I705139,I705122,I280304);
nor I_41330 (I705156,I705105,I705139);
DFFARX1 I_41331 (I705156,I2507,I704958,I704923,);
not I_41332 (I705187,I705139);
nand I_41333 (I705204,I705009,I705187);
nand I_41334 (I704935,I705071,I705187);
DFFARX1 I_41335 (I705105,I2507,I704958,I704950,);
not I_41336 (I705249,I280292);
nor I_41337 (I705266,I705249,I280283);
nor I_41338 (I705283,I705266,I705088);
DFFARX1 I_41339 (I705283,I2507,I704958,I704947,);
not I_41340 (I705314,I705266);
DFFARX1 I_41341 (I705314,I2507,I704958,I705340,);
not I_41342 (I705348,I705340);
nor I_41343 (I704944,I705348,I705266);
nor I_41344 (I705379,I705249,I280289);
and I_41345 (I705396,I705379,I280301);
or I_41346 (I705413,I705396,I280298);
DFFARX1 I_41347 (I705413,I2507,I704958,I705439,);
not I_41348 (I705447,I705439);
nand I_41349 (I705464,I705447,I705187);
not I_41350 (I704938,I705464);
nand I_41351 (I704932,I705464,I705204);
nand I_41352 (I704929,I705447,I705071);
not I_41353 (I705553,I2514);
DFFARX1 I_41354 (I397550,I2507,I705553,I705579,);
DFFARX1 I_41355 (I397532,I2507,I705553,I705596,);
not I_41356 (I705604,I705596);
nor I_41357 (I705521,I705579,I705604);
DFFARX1 I_41358 (I705604,I2507,I705553,I705536,);
nor I_41359 (I705649,I397538,I397541);
and I_41360 (I705666,I705649,I397529);
nor I_41361 (I705683,I705666,I397538);
not I_41362 (I705700,I397538);
and I_41363 (I705717,I705700,I397547);
nand I_41364 (I705734,I705717,I397535);
nor I_41365 (I705751,I705700,I705734);
DFFARX1 I_41366 (I705751,I2507,I705553,I705518,);
not I_41367 (I705782,I705734);
nand I_41368 (I705799,I705604,I705782);
nand I_41369 (I705530,I705666,I705782);
DFFARX1 I_41370 (I705700,I2507,I705553,I705545,);
not I_41371 (I705844,I397532);
nor I_41372 (I705861,I705844,I397547);
nor I_41373 (I705878,I705861,I705683);
DFFARX1 I_41374 (I705878,I2507,I705553,I705542,);
not I_41375 (I705909,I705861);
DFFARX1 I_41376 (I705909,I2507,I705553,I705935,);
not I_41377 (I705943,I705935);
nor I_41378 (I705539,I705943,I705861);
nor I_41379 (I705974,I705844,I397544);
and I_41380 (I705991,I705974,I397553);
or I_41381 (I706008,I705991,I397529);
DFFARX1 I_41382 (I706008,I2507,I705553,I706034,);
not I_41383 (I706042,I706034);
nand I_41384 (I706059,I706042,I705782);
not I_41385 (I705533,I706059);
nand I_41386 (I705527,I706059,I705799);
nand I_41387 (I705524,I706042,I705666);
not I_41388 (I706148,I2514);
DFFARX1 I_41389 (I441296,I2507,I706148,I706174,);
DFFARX1 I_41390 (I441293,I2507,I706148,I706191,);
not I_41391 (I706199,I706191);
nor I_41392 (I706116,I706174,I706199);
DFFARX1 I_41393 (I706199,I2507,I706148,I706131,);
nor I_41394 (I706244,I441308,I441290);
and I_41395 (I706261,I706244,I441287);
nor I_41396 (I706278,I706261,I441308);
not I_41397 (I706295,I441308);
and I_41398 (I706312,I706295,I441293);
nand I_41399 (I706329,I706312,I441305);
nor I_41400 (I706346,I706295,I706329);
DFFARX1 I_41401 (I706346,I2507,I706148,I706113,);
not I_41402 (I706377,I706329);
nand I_41403 (I706394,I706199,I706377);
nand I_41404 (I706125,I706261,I706377);
DFFARX1 I_41405 (I706295,I2507,I706148,I706140,);
not I_41406 (I706439,I441299);
nor I_41407 (I706456,I706439,I441293);
nor I_41408 (I706473,I706456,I706278);
DFFARX1 I_41409 (I706473,I2507,I706148,I706137,);
not I_41410 (I706504,I706456);
DFFARX1 I_41411 (I706504,I2507,I706148,I706530,);
not I_41412 (I706538,I706530);
nor I_41413 (I706134,I706538,I706456);
nor I_41414 (I706569,I706439,I441287);
and I_41415 (I706586,I706569,I441302);
or I_41416 (I706603,I706586,I441290);
DFFARX1 I_41417 (I706603,I2507,I706148,I706629,);
not I_41418 (I706637,I706629);
nand I_41419 (I706654,I706637,I706377);
not I_41420 (I706128,I706654);
nand I_41421 (I706122,I706654,I706394);
nand I_41422 (I706119,I706637,I706261);
not I_41423 (I706743,I2514);
DFFARX1 I_41424 (I319520,I2507,I706743,I706769,);
DFFARX1 I_41425 (I319514,I2507,I706743,I706786,);
not I_41426 (I706794,I706786);
nor I_41427 (I706711,I706769,I706794);
DFFARX1 I_41428 (I706794,I2507,I706743,I706726,);
nor I_41429 (I706839,I319511,I319502);
and I_41430 (I706856,I706839,I319499);
nor I_41431 (I706873,I706856,I319511);
not I_41432 (I706890,I319511);
and I_41433 (I706907,I706890,I319505);
nand I_41434 (I706924,I706907,I319517);
nor I_41435 (I706941,I706890,I706924);
DFFARX1 I_41436 (I706941,I2507,I706743,I706708,);
not I_41437 (I706972,I706924);
nand I_41438 (I706989,I706794,I706972);
nand I_41439 (I706720,I706856,I706972);
DFFARX1 I_41440 (I706890,I2507,I706743,I706735,);
not I_41441 (I707034,I319523);
nor I_41442 (I707051,I707034,I319505);
nor I_41443 (I707068,I707051,I706873);
DFFARX1 I_41444 (I707068,I2507,I706743,I706732,);
not I_41445 (I707099,I707051);
DFFARX1 I_41446 (I707099,I2507,I706743,I707125,);
not I_41447 (I707133,I707125);
nor I_41448 (I706729,I707133,I707051);
nor I_41449 (I707164,I707034,I319502);
and I_41450 (I707181,I707164,I319508);
or I_41451 (I707198,I707181,I319499);
DFFARX1 I_41452 (I707198,I2507,I706743,I707224,);
not I_41453 (I707232,I707224);
nand I_41454 (I707249,I707232,I706972);
not I_41455 (I706723,I707249);
nand I_41456 (I706717,I707249,I706989);
nand I_41457 (I706714,I707232,I706856);
not I_41458 (I707338,I2514);
DFFARX1 I_41459 (I415468,I2507,I707338,I707364,);
DFFARX1 I_41460 (I415450,I2507,I707338,I707381,);
not I_41461 (I707389,I707381);
nor I_41462 (I707306,I707364,I707389);
DFFARX1 I_41463 (I707389,I2507,I707338,I707321,);
nor I_41464 (I707434,I415456,I415459);
and I_41465 (I707451,I707434,I415447);
nor I_41466 (I707468,I707451,I415456);
not I_41467 (I707485,I415456);
and I_41468 (I707502,I707485,I415465);
nand I_41469 (I707519,I707502,I415453);
nor I_41470 (I707536,I707485,I707519);
DFFARX1 I_41471 (I707536,I2507,I707338,I707303,);
not I_41472 (I707567,I707519);
nand I_41473 (I707584,I707389,I707567);
nand I_41474 (I707315,I707451,I707567);
DFFARX1 I_41475 (I707485,I2507,I707338,I707330,);
not I_41476 (I707629,I415450);
nor I_41477 (I707646,I707629,I415465);
nor I_41478 (I707663,I707646,I707468);
DFFARX1 I_41479 (I707663,I2507,I707338,I707327,);
not I_41480 (I707694,I707646);
DFFARX1 I_41481 (I707694,I2507,I707338,I707720,);
not I_41482 (I707728,I707720);
nor I_41483 (I707324,I707728,I707646);
nor I_41484 (I707759,I707629,I415462);
and I_41485 (I707776,I707759,I415471);
or I_41486 (I707793,I707776,I415447);
DFFARX1 I_41487 (I707793,I2507,I707338,I707819,);
not I_41488 (I707827,I707819);
nand I_41489 (I707844,I707827,I707567);
not I_41490 (I707318,I707844);
nand I_41491 (I707312,I707844,I707584);
nand I_41492 (I707309,I707827,I707451);
not I_41493 (I707933,I2514);
DFFARX1 I_41494 (I466065,I2507,I707933,I707959,);
DFFARX1 I_41495 (I466062,I2507,I707933,I707976,);
not I_41496 (I707984,I707976);
nor I_41497 (I707901,I707959,I707984);
DFFARX1 I_41498 (I707984,I2507,I707933,I707916,);
nor I_41499 (I708029,I466077,I466059);
and I_41500 (I708046,I708029,I466056);
nor I_41501 (I708063,I708046,I466077);
not I_41502 (I708080,I466077);
and I_41503 (I708097,I708080,I466062);
nand I_41504 (I708114,I708097,I466074);
nor I_41505 (I708131,I708080,I708114);
DFFARX1 I_41506 (I708131,I2507,I707933,I707898,);
not I_41507 (I708162,I708114);
nand I_41508 (I708179,I707984,I708162);
nand I_41509 (I707910,I708046,I708162);
DFFARX1 I_41510 (I708080,I2507,I707933,I707925,);
not I_41511 (I708224,I466068);
nor I_41512 (I708241,I708224,I466062);
nor I_41513 (I708258,I708241,I708063);
DFFARX1 I_41514 (I708258,I2507,I707933,I707922,);
not I_41515 (I708289,I708241);
DFFARX1 I_41516 (I708289,I2507,I707933,I708315,);
not I_41517 (I708323,I708315);
nor I_41518 (I707919,I708323,I708241);
nor I_41519 (I708354,I708224,I466056);
and I_41520 (I708371,I708354,I466071);
or I_41521 (I708388,I708371,I466059);
DFFARX1 I_41522 (I708388,I2507,I707933,I708414,);
not I_41523 (I708422,I708414);
nand I_41524 (I708439,I708422,I708162);
not I_41525 (I707913,I708439);
nand I_41526 (I707907,I708439,I708179);
nand I_41527 (I707904,I708422,I708046);
not I_41528 (I708528,I2514);
DFFARX1 I_41529 (I433391,I2507,I708528,I708554,);
DFFARX1 I_41530 (I433388,I2507,I708528,I708571,);
not I_41531 (I708579,I708571);
nor I_41532 (I708496,I708554,I708579);
DFFARX1 I_41533 (I708579,I2507,I708528,I708511,);
nor I_41534 (I708624,I433403,I433385);
and I_41535 (I708641,I708624,I433382);
nor I_41536 (I708658,I708641,I433403);
not I_41537 (I708675,I433403);
and I_41538 (I708692,I708675,I433388);
nand I_41539 (I708709,I708692,I433400);
nor I_41540 (I708726,I708675,I708709);
DFFARX1 I_41541 (I708726,I2507,I708528,I708493,);
not I_41542 (I708757,I708709);
nand I_41543 (I708774,I708579,I708757);
nand I_41544 (I708505,I708641,I708757);
DFFARX1 I_41545 (I708675,I2507,I708528,I708520,);
not I_41546 (I708819,I433394);
nor I_41547 (I708836,I708819,I433388);
nor I_41548 (I708853,I708836,I708658);
DFFARX1 I_41549 (I708853,I2507,I708528,I708517,);
not I_41550 (I708884,I708836);
DFFARX1 I_41551 (I708884,I2507,I708528,I708910,);
not I_41552 (I708918,I708910);
nor I_41553 (I708514,I708918,I708836);
nor I_41554 (I708949,I708819,I433382);
and I_41555 (I708966,I708949,I433397);
or I_41556 (I708983,I708966,I433385);
DFFARX1 I_41557 (I708983,I2507,I708528,I709009,);
not I_41558 (I709017,I709009);
nand I_41559 (I709034,I709017,I708757);
not I_41560 (I708508,I709034);
nand I_41561 (I708502,I709034,I708774);
nand I_41562 (I708499,I709017,I708641);
not I_41563 (I709123,I2514);
DFFARX1 I_41564 (I566606,I2507,I709123,I709149,);
DFFARX1 I_41565 (I566597,I2507,I709123,I709166,);
not I_41566 (I709174,I709166);
nor I_41567 (I709091,I709149,I709174);
DFFARX1 I_41568 (I709174,I2507,I709123,I709106,);
nor I_41569 (I709219,I566603,I566612);
and I_41570 (I709236,I709219,I566615);
nor I_41571 (I709253,I709236,I566603);
not I_41572 (I709270,I566603);
and I_41573 (I709287,I709270,I566594);
nand I_41574 (I709304,I709287,I566600);
nor I_41575 (I709321,I709270,I709304);
DFFARX1 I_41576 (I709321,I2507,I709123,I709088,);
not I_41577 (I709352,I709304);
nand I_41578 (I709369,I709174,I709352);
nand I_41579 (I709100,I709236,I709352);
DFFARX1 I_41580 (I709270,I2507,I709123,I709115,);
not I_41581 (I709414,I566609);
nor I_41582 (I709431,I709414,I566594);
nor I_41583 (I709448,I709431,I709253);
DFFARX1 I_41584 (I709448,I2507,I709123,I709112,);
not I_41585 (I709479,I709431);
DFFARX1 I_41586 (I709479,I2507,I709123,I709505,);
not I_41587 (I709513,I709505);
nor I_41588 (I709109,I709513,I709431);
nor I_41589 (I709544,I709414,I566594);
and I_41590 (I709561,I709544,I566597);
or I_41591 (I709578,I709561,I566600);
DFFARX1 I_41592 (I709578,I2507,I709123,I709604,);
not I_41593 (I709612,I709604);
nand I_41594 (I709629,I709612,I709352);
not I_41595 (I709103,I709629);
nand I_41596 (I709097,I709629,I709369);
nand I_41597 (I709094,I709612,I709236);
not I_41598 (I709718,I2514);
DFFARX1 I_41599 (I688919,I2507,I709718,I709744,);
DFFARX1 I_41600 (I688904,I2507,I709718,I709761,);
not I_41601 (I709769,I709761);
nor I_41602 (I709686,I709744,I709769);
DFFARX1 I_41603 (I709769,I2507,I709718,I709701,);
nor I_41604 (I709814,I688901,I688910);
and I_41605 (I709831,I709814,I688916);
nor I_41606 (I709848,I709831,I688901);
not I_41607 (I709865,I688901);
and I_41608 (I709882,I709865,I688898);
nand I_41609 (I709899,I709882,I688892);
nor I_41610 (I709916,I709865,I709899);
DFFARX1 I_41611 (I709916,I2507,I709718,I709683,);
not I_41612 (I709947,I709899);
nand I_41613 (I709964,I709769,I709947);
nand I_41614 (I709695,I709831,I709947);
DFFARX1 I_41615 (I709865,I2507,I709718,I709710,);
not I_41616 (I710009,I688892);
nor I_41617 (I710026,I710009,I688898);
nor I_41618 (I710043,I710026,I709848);
DFFARX1 I_41619 (I710043,I2507,I709718,I709707,);
not I_41620 (I710074,I710026);
DFFARX1 I_41621 (I710074,I2507,I709718,I710100,);
not I_41622 (I710108,I710100);
nor I_41623 (I709704,I710108,I710026);
nor I_41624 (I710139,I710009,I688907);
and I_41625 (I710156,I710139,I688913);
or I_41626 (I710173,I710156,I688895);
DFFARX1 I_41627 (I710173,I2507,I709718,I710199,);
not I_41628 (I710207,I710199);
nand I_41629 (I710224,I710207,I709947);
not I_41630 (I709698,I710224);
nand I_41631 (I709692,I710224,I709964);
nand I_41632 (I709689,I710207,I709831);
not I_41633 (I710313,I2514);
DFFARX1 I_41634 (I190116,I2507,I710313,I710339,);
DFFARX1 I_41635 (I190110,I2507,I710313,I710356,);
not I_41636 (I710364,I710356);
nor I_41637 (I710281,I710339,I710364);
DFFARX1 I_41638 (I710364,I2507,I710313,I710296,);
nor I_41639 (I710409,I190098,I190119);
and I_41640 (I710426,I710409,I190113);
nor I_41641 (I710443,I710426,I190098);
not I_41642 (I710460,I190098);
and I_41643 (I710477,I710460,I190095);
nand I_41644 (I710494,I710477,I190107);
nor I_41645 (I710511,I710460,I710494);
DFFARX1 I_41646 (I710511,I2507,I710313,I710278,);
not I_41647 (I710542,I710494);
nand I_41648 (I710559,I710364,I710542);
nand I_41649 (I710290,I710426,I710542);
DFFARX1 I_41650 (I710460,I2507,I710313,I710305,);
not I_41651 (I710604,I190122);
nor I_41652 (I710621,I710604,I190095);
nor I_41653 (I710638,I710621,I710443);
DFFARX1 I_41654 (I710638,I2507,I710313,I710302,);
not I_41655 (I710669,I710621);
DFFARX1 I_41656 (I710669,I2507,I710313,I710695,);
not I_41657 (I710703,I710695);
nor I_41658 (I710299,I710703,I710621);
nor I_41659 (I710734,I710604,I190104);
and I_41660 (I710751,I710734,I190101);
or I_41661 (I710768,I710751,I190095);
DFFARX1 I_41662 (I710768,I2507,I710313,I710794,);
not I_41663 (I710802,I710794);
nand I_41664 (I710819,I710802,I710542);
not I_41665 (I710293,I710819);
nand I_41666 (I710287,I710819,I710559);
nand I_41667 (I710284,I710802,I710426);
not I_41668 (I710908,I2514);
DFFARX1 I_41669 (I98499,I2507,I710908,I710934,);
DFFARX1 I_41670 (I98502,I2507,I710908,I710951,);
not I_41671 (I710959,I710951);
nor I_41672 (I710876,I710934,I710959);
DFFARX1 I_41673 (I710959,I2507,I710908,I710891,);
nor I_41674 (I711004,I98508,I98502);
and I_41675 (I711021,I711004,I98505);
nor I_41676 (I711038,I711021,I98508);
not I_41677 (I711055,I98508);
and I_41678 (I711072,I711055,I98499);
nand I_41679 (I711089,I711072,I98517);
nor I_41680 (I711106,I711055,I711089);
DFFARX1 I_41681 (I711106,I2507,I710908,I710873,);
not I_41682 (I711137,I711089);
nand I_41683 (I711154,I710959,I711137);
nand I_41684 (I710885,I711021,I711137);
DFFARX1 I_41685 (I711055,I2507,I710908,I710900,);
not I_41686 (I711199,I98511);
nor I_41687 (I711216,I711199,I98499);
nor I_41688 (I711233,I711216,I711038);
DFFARX1 I_41689 (I711233,I2507,I710908,I710897,);
not I_41690 (I711264,I711216);
DFFARX1 I_41691 (I711264,I2507,I710908,I711290,);
not I_41692 (I711298,I711290);
nor I_41693 (I710894,I711298,I711216);
nor I_41694 (I711329,I711199,I98514);
and I_41695 (I711346,I711329,I98520);
or I_41696 (I711363,I711346,I98523);
DFFARX1 I_41697 (I711363,I2507,I710908,I711389,);
not I_41698 (I711397,I711389);
nand I_41699 (I711414,I711397,I711137);
not I_41700 (I710888,I711414);
nand I_41701 (I710882,I711414,I711154);
nand I_41702 (I710879,I711397,I711021);
not I_41703 (I711503,I2514);
DFFARX1 I_41704 (I118134,I2507,I711503,I711529,);
DFFARX1 I_41705 (I118137,I2507,I711503,I711546,);
not I_41706 (I711554,I711546);
nor I_41707 (I711471,I711529,I711554);
DFFARX1 I_41708 (I711554,I2507,I711503,I711486,);
nor I_41709 (I711599,I118143,I118137);
and I_41710 (I711616,I711599,I118140);
nor I_41711 (I711633,I711616,I118143);
not I_41712 (I711650,I118143);
and I_41713 (I711667,I711650,I118134);
nand I_41714 (I711684,I711667,I118152);
nor I_41715 (I711701,I711650,I711684);
DFFARX1 I_41716 (I711701,I2507,I711503,I711468,);
not I_41717 (I711732,I711684);
nand I_41718 (I711749,I711554,I711732);
nand I_41719 (I711480,I711616,I711732);
DFFARX1 I_41720 (I711650,I2507,I711503,I711495,);
not I_41721 (I711794,I118146);
nor I_41722 (I711811,I711794,I118134);
nor I_41723 (I711828,I711811,I711633);
DFFARX1 I_41724 (I711828,I2507,I711503,I711492,);
not I_41725 (I711859,I711811);
DFFARX1 I_41726 (I711859,I2507,I711503,I711885,);
not I_41727 (I711893,I711885);
nor I_41728 (I711489,I711893,I711811);
nor I_41729 (I711924,I711794,I118149);
and I_41730 (I711941,I711924,I118155);
or I_41731 (I711958,I711941,I118158);
DFFARX1 I_41732 (I711958,I2507,I711503,I711984,);
not I_41733 (I711992,I711984);
nand I_41734 (I712009,I711992,I711732);
not I_41735 (I711483,I712009);
nand I_41736 (I711477,I712009,I711749);
nand I_41737 (I711474,I711992,I711616);
not I_41738 (I712098,I2514);
DFFARX1 I_41739 (I362870,I2507,I712098,I712124,);
DFFARX1 I_41740 (I362852,I2507,I712098,I712141,);
not I_41741 (I712149,I712141);
nor I_41742 (I712066,I712124,I712149);
DFFARX1 I_41743 (I712149,I2507,I712098,I712081,);
nor I_41744 (I712194,I362858,I362861);
and I_41745 (I712211,I712194,I362849);
nor I_41746 (I712228,I712211,I362858);
not I_41747 (I712245,I362858);
and I_41748 (I712262,I712245,I362867);
nand I_41749 (I712279,I712262,I362855);
nor I_41750 (I712296,I712245,I712279);
DFFARX1 I_41751 (I712296,I2507,I712098,I712063,);
not I_41752 (I712327,I712279);
nand I_41753 (I712344,I712149,I712327);
nand I_41754 (I712075,I712211,I712327);
DFFARX1 I_41755 (I712245,I2507,I712098,I712090,);
not I_41756 (I712389,I362852);
nor I_41757 (I712406,I712389,I362867);
nor I_41758 (I712423,I712406,I712228);
DFFARX1 I_41759 (I712423,I2507,I712098,I712087,);
not I_41760 (I712454,I712406);
DFFARX1 I_41761 (I712454,I2507,I712098,I712480,);
not I_41762 (I712488,I712480);
nor I_41763 (I712084,I712488,I712406);
nor I_41764 (I712519,I712389,I362864);
and I_41765 (I712536,I712519,I362873);
or I_41766 (I712553,I712536,I362849);
DFFARX1 I_41767 (I712553,I2507,I712098,I712579,);
not I_41768 (I712587,I712579);
nand I_41769 (I712604,I712587,I712327);
not I_41770 (I712078,I712604);
nand I_41771 (I712072,I712604,I712344);
nand I_41772 (I712069,I712587,I712211);
not I_41773 (I712693,I2514);
DFFARX1 I_41774 (I634682,I2507,I712693,I712719,);
DFFARX1 I_41775 (I634694,I2507,I712693,I712736,);
not I_41776 (I712744,I712736);
nor I_41777 (I712661,I712719,I712744);
DFFARX1 I_41778 (I712744,I2507,I712693,I712676,);
nor I_41779 (I712789,I634691,I634685);
and I_41780 (I712806,I712789,I634679);
nor I_41781 (I712823,I712806,I634691);
not I_41782 (I712840,I634691);
and I_41783 (I712857,I712840,I634688);
nand I_41784 (I712874,I712857,I634679);
nor I_41785 (I712891,I712840,I712874);
DFFARX1 I_41786 (I712891,I2507,I712693,I712658,);
not I_41787 (I712922,I712874);
nand I_41788 (I712939,I712744,I712922);
nand I_41789 (I712670,I712806,I712922);
DFFARX1 I_41790 (I712840,I2507,I712693,I712685,);
not I_41791 (I712984,I634703);
nor I_41792 (I713001,I712984,I634688);
nor I_41793 (I713018,I713001,I712823);
DFFARX1 I_41794 (I713018,I2507,I712693,I712682,);
not I_41795 (I713049,I713001);
DFFARX1 I_41796 (I713049,I2507,I712693,I713075,);
not I_41797 (I713083,I713075);
nor I_41798 (I712679,I713083,I713001);
nor I_41799 (I713114,I712984,I634697);
and I_41800 (I713131,I713114,I634700);
or I_41801 (I713148,I713131,I634682);
DFFARX1 I_41802 (I713148,I2507,I712693,I713174,);
not I_41803 (I713182,I713174);
nand I_41804 (I713199,I713182,I712922);
not I_41805 (I712673,I713199);
nand I_41806 (I712667,I713199,I712939);
nand I_41807 (I712664,I713182,I712806);
not I_41808 (I713288,I2514);
DFFARX1 I_41809 (I244920,I2507,I713288,I713314,);
DFFARX1 I_41810 (I244926,I2507,I713288,I713331,);
not I_41811 (I713339,I713331);
nor I_41812 (I713256,I713314,I713339);
DFFARX1 I_41813 (I713339,I2507,I713288,I713271,);
nor I_41814 (I713384,I244935,I244920);
and I_41815 (I713401,I713384,I244947);
nor I_41816 (I713418,I713401,I244935);
not I_41817 (I713435,I244935);
and I_41818 (I713452,I713435,I244923);
nand I_41819 (I713469,I713452,I244944);
nor I_41820 (I713486,I713435,I713469);
DFFARX1 I_41821 (I713486,I2507,I713288,I713253,);
not I_41822 (I713517,I713469);
nand I_41823 (I713534,I713339,I713517);
nand I_41824 (I713265,I713401,I713517);
DFFARX1 I_41825 (I713435,I2507,I713288,I713280,);
not I_41826 (I713579,I244932);
nor I_41827 (I713596,I713579,I244923);
nor I_41828 (I713613,I713596,I713418);
DFFARX1 I_41829 (I713613,I2507,I713288,I713277,);
not I_41830 (I713644,I713596);
DFFARX1 I_41831 (I713644,I2507,I713288,I713670,);
not I_41832 (I713678,I713670);
nor I_41833 (I713274,I713678,I713596);
nor I_41834 (I713709,I713579,I244929);
and I_41835 (I713726,I713709,I244941);
or I_41836 (I713743,I713726,I244938);
DFFARX1 I_41837 (I713743,I2507,I713288,I713769,);
not I_41838 (I713777,I713769);
nand I_41839 (I713794,I713777,I713517);
not I_41840 (I713268,I713794);
nand I_41841 (I713262,I713794,I713534);
nand I_41842 (I713259,I713777,I713401);
not I_41843 (I713883,I2514);
DFFARX1 I_41844 (I446039,I2507,I713883,I713909,);
DFFARX1 I_41845 (I446036,I2507,I713883,I713926,);
not I_41846 (I713934,I713926);
nor I_41847 (I713851,I713909,I713934);
DFFARX1 I_41848 (I713934,I2507,I713883,I713866,);
nor I_41849 (I713979,I446051,I446033);
and I_41850 (I713996,I713979,I446030);
nor I_41851 (I714013,I713996,I446051);
not I_41852 (I714030,I446051);
and I_41853 (I714047,I714030,I446036);
nand I_41854 (I714064,I714047,I446048);
nor I_41855 (I714081,I714030,I714064);
DFFARX1 I_41856 (I714081,I2507,I713883,I713848,);
not I_41857 (I714112,I714064);
nand I_41858 (I714129,I713934,I714112);
nand I_41859 (I713860,I713996,I714112);
DFFARX1 I_41860 (I714030,I2507,I713883,I713875,);
not I_41861 (I714174,I446042);
nor I_41862 (I714191,I714174,I446036);
nor I_41863 (I714208,I714191,I714013);
DFFARX1 I_41864 (I714208,I2507,I713883,I713872,);
not I_41865 (I714239,I714191);
DFFARX1 I_41866 (I714239,I2507,I713883,I714265,);
not I_41867 (I714273,I714265);
nor I_41868 (I713869,I714273,I714191);
nor I_41869 (I714304,I714174,I446030);
and I_41870 (I714321,I714304,I446045);
or I_41871 (I714338,I714321,I446033);
DFFARX1 I_41872 (I714338,I2507,I713883,I714364,);
not I_41873 (I714372,I714364);
nand I_41874 (I714389,I714372,I714112);
not I_41875 (I713863,I714389);
nand I_41876 (I713857,I714389,I714129);
nand I_41877 (I713854,I714372,I713996);
not I_41878 (I714478,I2514);
DFFARX1 I_41879 (I456579,I2507,I714478,I714504,);
DFFARX1 I_41880 (I456576,I2507,I714478,I714521,);
not I_41881 (I714529,I714521);
nor I_41882 (I714446,I714504,I714529);
DFFARX1 I_41883 (I714529,I2507,I714478,I714461,);
nor I_41884 (I714574,I456591,I456573);
and I_41885 (I714591,I714574,I456570);
nor I_41886 (I714608,I714591,I456591);
not I_41887 (I714625,I456591);
and I_41888 (I714642,I714625,I456576);
nand I_41889 (I714659,I714642,I456588);
nor I_41890 (I714676,I714625,I714659);
DFFARX1 I_41891 (I714676,I2507,I714478,I714443,);
not I_41892 (I714707,I714659);
nand I_41893 (I714724,I714529,I714707);
nand I_41894 (I714455,I714591,I714707);
DFFARX1 I_41895 (I714625,I2507,I714478,I714470,);
not I_41896 (I714769,I456582);
nor I_41897 (I714786,I714769,I456576);
nor I_41898 (I714803,I714786,I714608);
DFFARX1 I_41899 (I714803,I2507,I714478,I714467,);
not I_41900 (I714834,I714786);
DFFARX1 I_41901 (I714834,I2507,I714478,I714860,);
not I_41902 (I714868,I714860);
nor I_41903 (I714464,I714868,I714786);
nor I_41904 (I714899,I714769,I456570);
and I_41905 (I714916,I714899,I456585);
or I_41906 (I714933,I714916,I456573);
DFFARX1 I_41907 (I714933,I2507,I714478,I714959,);
not I_41908 (I714967,I714959);
nand I_41909 (I714984,I714967,I714707);
not I_41910 (I714458,I714984);
nand I_41911 (I714452,I714984,I714724);
nand I_41912 (I714449,I714967,I714591);
not I_41913 (I715073,I2514);
DFFARX1 I_41914 (I161569,I2507,I715073,I715099,);
DFFARX1 I_41915 (I161572,I2507,I715073,I715116,);
not I_41916 (I715124,I715116);
nor I_41917 (I715041,I715099,I715124);
DFFARX1 I_41918 (I715124,I2507,I715073,I715056,);
nor I_41919 (I715169,I161578,I161572);
and I_41920 (I715186,I715169,I161575);
nor I_41921 (I715203,I715186,I161578);
not I_41922 (I715220,I161578);
and I_41923 (I715237,I715220,I161569);
nand I_41924 (I715254,I715237,I161587);
nor I_41925 (I715271,I715220,I715254);
DFFARX1 I_41926 (I715271,I2507,I715073,I715038,);
not I_41927 (I715302,I715254);
nand I_41928 (I715319,I715124,I715302);
nand I_41929 (I715050,I715186,I715302);
DFFARX1 I_41930 (I715220,I2507,I715073,I715065,);
not I_41931 (I715364,I161581);
nor I_41932 (I715381,I715364,I161569);
nor I_41933 (I715398,I715381,I715203);
DFFARX1 I_41934 (I715398,I2507,I715073,I715062,);
not I_41935 (I715429,I715381);
DFFARX1 I_41936 (I715429,I2507,I715073,I715455,);
not I_41937 (I715463,I715455);
nor I_41938 (I715059,I715463,I715381);
nor I_41939 (I715494,I715364,I161584);
and I_41940 (I715511,I715494,I161590);
or I_41941 (I715528,I715511,I161593);
DFFARX1 I_41942 (I715528,I2507,I715073,I715554,);
not I_41943 (I715562,I715554);
nand I_41944 (I715579,I715562,I715302);
not I_41945 (I715053,I715579);
nand I_41946 (I715047,I715579,I715319);
nand I_41947 (I715044,I715562,I715186);
not I_41948 (I715668,I2514);
DFFARX1 I_41949 (I172725,I2507,I715668,I715694,);
DFFARX1 I_41950 (I172719,I2507,I715668,I715711,);
not I_41951 (I715719,I715711);
nor I_41952 (I715636,I715694,I715719);
DFFARX1 I_41953 (I715719,I2507,I715668,I715651,);
nor I_41954 (I715764,I172707,I172728);
and I_41955 (I715781,I715764,I172722);
nor I_41956 (I715798,I715781,I172707);
not I_41957 (I715815,I172707);
and I_41958 (I715832,I715815,I172704);
nand I_41959 (I715849,I715832,I172716);
nor I_41960 (I715866,I715815,I715849);
DFFARX1 I_41961 (I715866,I2507,I715668,I715633,);
not I_41962 (I715897,I715849);
nand I_41963 (I715914,I715719,I715897);
nand I_41964 (I715645,I715781,I715897);
DFFARX1 I_41965 (I715815,I2507,I715668,I715660,);
not I_41966 (I715959,I172731);
nor I_41967 (I715976,I715959,I172704);
nor I_41968 (I715993,I715976,I715798);
DFFARX1 I_41969 (I715993,I2507,I715668,I715657,);
not I_41970 (I716024,I715976);
DFFARX1 I_41971 (I716024,I2507,I715668,I716050,);
not I_41972 (I716058,I716050);
nor I_41973 (I715654,I716058,I715976);
nor I_41974 (I716089,I715959,I172713);
and I_41975 (I716106,I716089,I172710);
or I_41976 (I716123,I716106,I172704);
DFFARX1 I_41977 (I716123,I2507,I715668,I716149,);
not I_41978 (I716157,I716149);
nand I_41979 (I716174,I716157,I715897);
not I_41980 (I715648,I716174);
nand I_41981 (I715642,I716174,I715914);
nand I_41982 (I715639,I716157,I715781);
not I_41983 (I716263,I2514);
DFFARX1 I_41984 (I582084,I2507,I716263,I716289,);
DFFARX1 I_41985 (I582096,I2507,I716263,I716306,);
not I_41986 (I716314,I716306);
nor I_41987 (I716231,I716289,I716314);
DFFARX1 I_41988 (I716314,I2507,I716263,I716246,);
nor I_41989 (I716359,I582093,I582087);
and I_41990 (I716376,I716359,I582081);
nor I_41991 (I716393,I716376,I582093);
not I_41992 (I716410,I582093);
and I_41993 (I716427,I716410,I582090);
nand I_41994 (I716444,I716427,I582081);
nor I_41995 (I716461,I716410,I716444);
DFFARX1 I_41996 (I716461,I2507,I716263,I716228,);
not I_41997 (I716492,I716444);
nand I_41998 (I716509,I716314,I716492);
nand I_41999 (I716240,I716376,I716492);
DFFARX1 I_42000 (I716410,I2507,I716263,I716255,);
not I_42001 (I716554,I582105);
nor I_42002 (I716571,I716554,I582090);
nor I_42003 (I716588,I716571,I716393);
DFFARX1 I_42004 (I716588,I2507,I716263,I716252,);
not I_42005 (I716619,I716571);
DFFARX1 I_42006 (I716619,I2507,I716263,I716645,);
not I_42007 (I716653,I716645);
nor I_42008 (I716249,I716653,I716571);
nor I_42009 (I716684,I716554,I582099);
and I_42010 (I716701,I716684,I582102);
or I_42011 (I716718,I716701,I582084);
DFFARX1 I_42012 (I716718,I2507,I716263,I716744,);
not I_42013 (I716752,I716744);
nand I_42014 (I716769,I716752,I716492);
not I_42015 (I716243,I716769);
nand I_42016 (I716237,I716769,I716509);
nand I_42017 (I716234,I716752,I716376);
not I_42018 (I716858,I2514);
DFFARX1 I_42019 (I559874,I2507,I716858,I716884,);
DFFARX1 I_42020 (I559865,I2507,I716858,I716901,);
not I_42021 (I716909,I716901);
nor I_42022 (I716826,I716884,I716909);
DFFARX1 I_42023 (I716909,I2507,I716858,I716841,);
nor I_42024 (I716954,I559871,I559880);
and I_42025 (I716971,I716954,I559883);
nor I_42026 (I716988,I716971,I559871);
not I_42027 (I717005,I559871);
and I_42028 (I717022,I717005,I559862);
nand I_42029 (I717039,I717022,I559868);
nor I_42030 (I717056,I717005,I717039);
DFFARX1 I_42031 (I717056,I2507,I716858,I716823,);
not I_42032 (I717087,I717039);
nand I_42033 (I717104,I716909,I717087);
nand I_42034 (I716835,I716971,I717087);
DFFARX1 I_42035 (I717005,I2507,I716858,I716850,);
not I_42036 (I717149,I559877);
nor I_42037 (I717166,I717149,I559862);
nor I_42038 (I717183,I717166,I716988);
DFFARX1 I_42039 (I717183,I2507,I716858,I716847,);
not I_42040 (I717214,I717166);
DFFARX1 I_42041 (I717214,I2507,I716858,I717240,);
not I_42042 (I717248,I717240);
nor I_42043 (I716844,I717248,I717166);
nor I_42044 (I717279,I717149,I559862);
and I_42045 (I717296,I717279,I559865);
or I_42046 (I717313,I717296,I559868);
DFFARX1 I_42047 (I717313,I2507,I716858,I717339,);
not I_42048 (I717347,I717339);
nand I_42049 (I717364,I717347,I717087);
not I_42050 (I716838,I717364);
nand I_42051 (I716832,I717364,I717104);
nand I_42052 (I716829,I717347,I716971);
not I_42053 (I717453,I2514);
DFFARX1 I_42054 (I522876,I2507,I717453,I717479,);
DFFARX1 I_42055 (I522894,I2507,I717453,I717496,);
not I_42056 (I717504,I717496);
nor I_42057 (I717421,I717479,I717504);
DFFARX1 I_42058 (I717504,I2507,I717453,I717436,);
nor I_42059 (I717549,I522873,I522885);
and I_42060 (I717566,I717549,I522870);
nor I_42061 (I717583,I717566,I522873);
not I_42062 (I717600,I522873);
and I_42063 (I717617,I717600,I522879);
nand I_42064 (I717634,I717617,I522891);
nor I_42065 (I717651,I717600,I717634);
DFFARX1 I_42066 (I717651,I2507,I717453,I717418,);
not I_42067 (I717682,I717634);
nand I_42068 (I717699,I717504,I717682);
nand I_42069 (I717430,I717566,I717682);
DFFARX1 I_42070 (I717600,I2507,I717453,I717445,);
not I_42071 (I717744,I522882);
nor I_42072 (I717761,I717744,I522879);
nor I_42073 (I717778,I717761,I717583);
DFFARX1 I_42074 (I717778,I2507,I717453,I717442,);
not I_42075 (I717809,I717761);
DFFARX1 I_42076 (I717809,I2507,I717453,I717835,);
not I_42077 (I717843,I717835);
nor I_42078 (I717439,I717843,I717761);
nor I_42079 (I717874,I717744,I522870);
and I_42080 (I717891,I717874,I522897);
or I_42081 (I717908,I717891,I522888);
DFFARX1 I_42082 (I717908,I2507,I717453,I717934,);
not I_42083 (I717942,I717934);
nand I_42084 (I717959,I717942,I717682);
not I_42085 (I717433,I717959);
nand I_42086 (I717427,I717959,I717699);
nand I_42087 (I717424,I717942,I717566);
not I_42088 (I718048,I2514);
DFFARX1 I_42089 (I609250,I2507,I718048,I718074,);
DFFARX1 I_42090 (I609262,I2507,I718048,I718091,);
not I_42091 (I718099,I718091);
nor I_42092 (I718016,I718074,I718099);
DFFARX1 I_42093 (I718099,I2507,I718048,I718031,);
nor I_42094 (I718144,I609259,I609253);
and I_42095 (I718161,I718144,I609247);
nor I_42096 (I718178,I718161,I609259);
not I_42097 (I718195,I609259);
and I_42098 (I718212,I718195,I609256);
nand I_42099 (I718229,I718212,I609247);
nor I_42100 (I718246,I718195,I718229);
DFFARX1 I_42101 (I718246,I2507,I718048,I718013,);
not I_42102 (I718277,I718229);
nand I_42103 (I718294,I718099,I718277);
nand I_42104 (I718025,I718161,I718277);
DFFARX1 I_42105 (I718195,I2507,I718048,I718040,);
not I_42106 (I718339,I609271);
nor I_42107 (I718356,I718339,I609256);
nor I_42108 (I718373,I718356,I718178);
DFFARX1 I_42109 (I718373,I2507,I718048,I718037,);
not I_42110 (I718404,I718356);
DFFARX1 I_42111 (I718404,I2507,I718048,I718430,);
not I_42112 (I718438,I718430);
nor I_42113 (I718034,I718438,I718356);
nor I_42114 (I718469,I718339,I609265);
and I_42115 (I718486,I718469,I609268);
or I_42116 (I718503,I718486,I609250);
DFFARX1 I_42117 (I718503,I2507,I718048,I718529,);
not I_42118 (I718537,I718529);
nand I_42119 (I718554,I718537,I718277);
not I_42120 (I718028,I718554);
nand I_42121 (I718022,I718554,I718294);
nand I_42122 (I718019,I718537,I718161);
not I_42123 (I718643,I2514);
DFFARX1 I_42124 (I495098,I2507,I718643,I718669,);
DFFARX1 I_42125 (I495116,I2507,I718643,I718686,);
not I_42126 (I718694,I718686);
nor I_42127 (I718611,I718669,I718694);
DFFARX1 I_42128 (I718694,I2507,I718643,I718626,);
nor I_42129 (I718739,I495095,I495107);
and I_42130 (I718756,I718739,I495092);
nor I_42131 (I718773,I718756,I495095);
not I_42132 (I718790,I495095);
and I_42133 (I718807,I718790,I495101);
nand I_42134 (I718824,I718807,I495113);
nor I_42135 (I718841,I718790,I718824);
DFFARX1 I_42136 (I718841,I2507,I718643,I718608,);
not I_42137 (I718872,I718824);
nand I_42138 (I718889,I718694,I718872);
nand I_42139 (I718620,I718756,I718872);
DFFARX1 I_42140 (I718790,I2507,I718643,I718635,);
not I_42141 (I718934,I495104);
nor I_42142 (I718951,I718934,I495101);
nor I_42143 (I718968,I718951,I718773);
DFFARX1 I_42144 (I718968,I2507,I718643,I718632,);
not I_42145 (I718999,I718951);
DFFARX1 I_42146 (I718999,I2507,I718643,I719025,);
not I_42147 (I719033,I719025);
nor I_42148 (I718629,I719033,I718951);
nor I_42149 (I719064,I718934,I495092);
and I_42150 (I719081,I719064,I495119);
or I_42151 (I719098,I719081,I495110);
DFFARX1 I_42152 (I719098,I2507,I718643,I719124,);
not I_42153 (I719132,I719124);
nand I_42154 (I719149,I719132,I718872);
not I_42155 (I718623,I719149);
nand I_42156 (I718617,I719149,I718889);
nand I_42157 (I718614,I719132,I718756);
not I_42158 (I719238,I2514);
DFFARX1 I_42159 (I487346,I2507,I719238,I719264,);
DFFARX1 I_42160 (I487364,I2507,I719238,I719281,);
not I_42161 (I719289,I719281);
nor I_42162 (I719206,I719264,I719289);
DFFARX1 I_42163 (I719289,I2507,I719238,I719221,);
nor I_42164 (I719334,I487343,I487355);
and I_42165 (I719351,I719334,I487340);
nor I_42166 (I719368,I719351,I487343);
not I_42167 (I719385,I487343);
and I_42168 (I719402,I719385,I487349);
nand I_42169 (I719419,I719402,I487361);
nor I_42170 (I719436,I719385,I719419);
DFFARX1 I_42171 (I719436,I2507,I719238,I719203,);
not I_42172 (I719467,I719419);
nand I_42173 (I719484,I719289,I719467);
nand I_42174 (I719215,I719351,I719467);
DFFARX1 I_42175 (I719385,I2507,I719238,I719230,);
not I_42176 (I719529,I487352);
nor I_42177 (I719546,I719529,I487349);
nor I_42178 (I719563,I719546,I719368);
DFFARX1 I_42179 (I719563,I2507,I719238,I719227,);
not I_42180 (I719594,I719546);
DFFARX1 I_42181 (I719594,I2507,I719238,I719620,);
not I_42182 (I719628,I719620);
nor I_42183 (I719224,I719628,I719546);
nor I_42184 (I719659,I719529,I487340);
and I_42185 (I719676,I719659,I487367);
or I_42186 (I719693,I719676,I487358);
DFFARX1 I_42187 (I719693,I2507,I719238,I719719,);
not I_42188 (I719727,I719719);
nand I_42189 (I719744,I719727,I719467);
not I_42190 (I719218,I719744);
nand I_42191 (I719212,I719744,I719484);
nand I_42192 (I719209,I719727,I719351);
not I_42193 (I719833,I2514);
DFFARX1 I_42194 (I674613,I2507,I719833,I719859,);
DFFARX1 I_42195 (I674604,I2507,I719833,I719876,);
not I_42196 (I719884,I719876);
nor I_42197 (I719801,I719859,I719884);
DFFARX1 I_42198 (I719884,I2507,I719833,I719816,);
nor I_42199 (I719929,I674595,I674610);
and I_42200 (I719946,I719929,I674598);
nor I_42201 (I719963,I719946,I674595);
not I_42202 (I719980,I674595);
and I_42203 (I719997,I719980,I674601);
nand I_42204 (I720014,I719997,I674619);
nor I_42205 (I720031,I719980,I720014);
DFFARX1 I_42206 (I720031,I2507,I719833,I719798,);
not I_42207 (I720062,I720014);
nand I_42208 (I720079,I719884,I720062);
nand I_42209 (I719810,I719946,I720062);
DFFARX1 I_42210 (I719980,I2507,I719833,I719825,);
not I_42211 (I720124,I674595);
nor I_42212 (I720141,I720124,I674601);
nor I_42213 (I720158,I720141,I719963);
DFFARX1 I_42214 (I720158,I2507,I719833,I719822,);
not I_42215 (I720189,I720141);
DFFARX1 I_42216 (I720189,I2507,I719833,I720215,);
not I_42217 (I720223,I720215);
nor I_42218 (I719819,I720223,I720141);
nor I_42219 (I720254,I720124,I674598);
and I_42220 (I720271,I720254,I674607);
or I_42221 (I720288,I720271,I674616);
DFFARX1 I_42222 (I720288,I2507,I719833,I720314,);
not I_42223 (I720322,I720314);
nand I_42224 (I720339,I720322,I720062);
not I_42225 (I719813,I720339);
nand I_42226 (I719807,I720339,I720079);
nand I_42227 (I719804,I720322,I719946);
not I_42228 (I720428,I2514);
DFFARX1 I_42229 (I467646,I2507,I720428,I720454,);
DFFARX1 I_42230 (I467643,I2507,I720428,I720471,);
not I_42231 (I720479,I720471);
nor I_42232 (I720396,I720454,I720479);
DFFARX1 I_42233 (I720479,I2507,I720428,I720411,);
nor I_42234 (I720524,I467658,I467640);
and I_42235 (I720541,I720524,I467637);
nor I_42236 (I720558,I720541,I467658);
not I_42237 (I720575,I467658);
and I_42238 (I720592,I720575,I467643);
nand I_42239 (I720609,I720592,I467655);
nor I_42240 (I720626,I720575,I720609);
DFFARX1 I_42241 (I720626,I2507,I720428,I720393,);
not I_42242 (I720657,I720609);
nand I_42243 (I720674,I720479,I720657);
nand I_42244 (I720405,I720541,I720657);
DFFARX1 I_42245 (I720575,I2507,I720428,I720420,);
not I_42246 (I720719,I467649);
nor I_42247 (I720736,I720719,I467643);
nor I_42248 (I720753,I720736,I720558);
DFFARX1 I_42249 (I720753,I2507,I720428,I720417,);
not I_42250 (I720784,I720736);
DFFARX1 I_42251 (I720784,I2507,I720428,I720810,);
not I_42252 (I720818,I720810);
nor I_42253 (I720414,I720818,I720736);
nor I_42254 (I720849,I720719,I467637);
and I_42255 (I720866,I720849,I467652);
or I_42256 (I720883,I720866,I467640);
DFFARX1 I_42257 (I720883,I2507,I720428,I720909,);
not I_42258 (I720917,I720909);
nand I_42259 (I720934,I720917,I720657);
not I_42260 (I720408,I720934);
nand I_42261 (I720402,I720934,I720674);
nand I_42262 (I720399,I720917,I720541);
not I_42263 (I721023,I2514);
DFFARX1 I_42264 (I431283,I2507,I721023,I721049,);
DFFARX1 I_42265 (I431280,I2507,I721023,I721066,);
not I_42266 (I721074,I721066);
nor I_42267 (I720991,I721049,I721074);
DFFARX1 I_42268 (I721074,I2507,I721023,I721006,);
nor I_42269 (I721119,I431295,I431277);
and I_42270 (I721136,I721119,I431274);
nor I_42271 (I721153,I721136,I431295);
not I_42272 (I721170,I431295);
and I_42273 (I721187,I721170,I431280);
nand I_42274 (I721204,I721187,I431292);
nor I_42275 (I721221,I721170,I721204);
DFFARX1 I_42276 (I721221,I2507,I721023,I720988,);
not I_42277 (I721252,I721204);
nand I_42278 (I721269,I721074,I721252);
nand I_42279 (I721000,I721136,I721252);
DFFARX1 I_42280 (I721170,I2507,I721023,I721015,);
not I_42281 (I721314,I431286);
nor I_42282 (I721331,I721314,I431280);
nor I_42283 (I721348,I721331,I721153);
DFFARX1 I_42284 (I721348,I2507,I721023,I721012,);
not I_42285 (I721379,I721331);
DFFARX1 I_42286 (I721379,I2507,I721023,I721405,);
not I_42287 (I721413,I721405);
nor I_42288 (I721009,I721413,I721331);
nor I_42289 (I721444,I721314,I431274);
and I_42290 (I721461,I721444,I431289);
or I_42291 (I721478,I721461,I431277);
DFFARX1 I_42292 (I721478,I2507,I721023,I721504,);
not I_42293 (I721512,I721504);
nand I_42294 (I721529,I721512,I721252);
not I_42295 (I721003,I721529);
nand I_42296 (I720997,I721529,I721269);
nand I_42297 (I720994,I721512,I721136);
not I_42298 (I721618,I2514);
DFFARX1 I_42299 (I137769,I2507,I721618,I721644,);
DFFARX1 I_42300 (I137772,I2507,I721618,I721661,);
not I_42301 (I721669,I721661);
nor I_42302 (I721586,I721644,I721669);
DFFARX1 I_42303 (I721669,I2507,I721618,I721601,);
nor I_42304 (I721714,I137778,I137772);
and I_42305 (I721731,I721714,I137775);
nor I_42306 (I721748,I721731,I137778);
not I_42307 (I721765,I137778);
and I_42308 (I721782,I721765,I137769);
nand I_42309 (I721799,I721782,I137787);
nor I_42310 (I721816,I721765,I721799);
DFFARX1 I_42311 (I721816,I2507,I721618,I721583,);
not I_42312 (I721847,I721799);
nand I_42313 (I721864,I721669,I721847);
nand I_42314 (I721595,I721731,I721847);
DFFARX1 I_42315 (I721765,I2507,I721618,I721610,);
not I_42316 (I721909,I137781);
nor I_42317 (I721926,I721909,I137769);
nor I_42318 (I721943,I721926,I721748);
DFFARX1 I_42319 (I721943,I2507,I721618,I721607,);
not I_42320 (I721974,I721926);
DFFARX1 I_42321 (I721974,I2507,I721618,I722000,);
not I_42322 (I722008,I722000);
nor I_42323 (I721604,I722008,I721926);
nor I_42324 (I722039,I721909,I137784);
and I_42325 (I722056,I722039,I137790);
or I_42326 (I722073,I722056,I137793);
DFFARX1 I_42327 (I722073,I2507,I721618,I722099,);
not I_42328 (I722107,I722099);
nand I_42329 (I722124,I722107,I721847);
not I_42330 (I721598,I722124);
nand I_42331 (I721592,I722124,I721864);
nand I_42332 (I721589,I722107,I721731);
not I_42333 (I722213,I2514);
DFFARX1 I_42334 (I602892,I2507,I722213,I722239,);
DFFARX1 I_42335 (I602904,I2507,I722213,I722256,);
not I_42336 (I722264,I722256);
nor I_42337 (I722181,I722239,I722264);
DFFARX1 I_42338 (I722264,I2507,I722213,I722196,);
nor I_42339 (I722309,I602901,I602895);
and I_42340 (I722326,I722309,I602889);
nor I_42341 (I722343,I722326,I602901);
not I_42342 (I722360,I602901);
and I_42343 (I722377,I722360,I602898);
nand I_42344 (I722394,I722377,I602889);
nor I_42345 (I722411,I722360,I722394);
DFFARX1 I_42346 (I722411,I2507,I722213,I722178,);
not I_42347 (I722442,I722394);
nand I_42348 (I722459,I722264,I722442);
nand I_42349 (I722190,I722326,I722442);
DFFARX1 I_42350 (I722360,I2507,I722213,I722205,);
not I_42351 (I722504,I602913);
nor I_42352 (I722521,I722504,I602898);
nor I_42353 (I722538,I722521,I722343);
DFFARX1 I_42354 (I722538,I2507,I722213,I722202,);
not I_42355 (I722569,I722521);
DFFARX1 I_42356 (I722569,I2507,I722213,I722595,);
not I_42357 (I722603,I722595);
nor I_42358 (I722199,I722603,I722521);
nor I_42359 (I722634,I722504,I602907);
and I_42360 (I722651,I722634,I602910);
or I_42361 (I722668,I722651,I602892);
DFFARX1 I_42362 (I722668,I2507,I722213,I722694,);
not I_42363 (I722702,I722694);
nand I_42364 (I722719,I722702,I722442);
not I_42365 (I722193,I722719);
nand I_42366 (I722187,I722719,I722459);
nand I_42367 (I722184,I722702,I722326);
not I_42368 (I722808,I2514);
DFFARX1 I_42369 (I124084,I2507,I722808,I722834,);
DFFARX1 I_42370 (I124087,I2507,I722808,I722851,);
not I_42371 (I722859,I722851);
nor I_42372 (I722776,I722834,I722859);
DFFARX1 I_42373 (I722859,I2507,I722808,I722791,);
nor I_42374 (I722904,I124093,I124087);
and I_42375 (I722921,I722904,I124090);
nor I_42376 (I722938,I722921,I124093);
not I_42377 (I722955,I124093);
and I_42378 (I722972,I722955,I124084);
nand I_42379 (I722989,I722972,I124102);
nor I_42380 (I723006,I722955,I722989);
DFFARX1 I_42381 (I723006,I2507,I722808,I722773,);
not I_42382 (I723037,I722989);
nand I_42383 (I723054,I722859,I723037);
nand I_42384 (I722785,I722921,I723037);
DFFARX1 I_42385 (I722955,I2507,I722808,I722800,);
not I_42386 (I723099,I124096);
nor I_42387 (I723116,I723099,I124084);
nor I_42388 (I723133,I723116,I722938);
DFFARX1 I_42389 (I723133,I2507,I722808,I722797,);
not I_42390 (I723164,I723116);
DFFARX1 I_42391 (I723164,I2507,I722808,I723190,);
not I_42392 (I723198,I723190);
nor I_42393 (I722794,I723198,I723116);
nor I_42394 (I723229,I723099,I124099);
and I_42395 (I723246,I723229,I124105);
or I_42396 (I723263,I723246,I124108);
DFFARX1 I_42397 (I723263,I2507,I722808,I723289,);
not I_42398 (I723297,I723289);
nand I_42399 (I723314,I723297,I723037);
not I_42400 (I722788,I723314);
nand I_42401 (I722782,I723314,I723054);
nand I_42402 (I722779,I723297,I722921);
not I_42403 (I723403,I2514);
DFFARX1 I_42404 (I402752,I2507,I723403,I723429,);
DFFARX1 I_42405 (I402734,I2507,I723403,I723446,);
not I_42406 (I723454,I723446);
nor I_42407 (I723371,I723429,I723454);
DFFARX1 I_42408 (I723454,I2507,I723403,I723386,);
nor I_42409 (I723499,I402740,I402743);
and I_42410 (I723516,I723499,I402731);
nor I_42411 (I723533,I723516,I402740);
not I_42412 (I723550,I402740);
and I_42413 (I723567,I723550,I402749);
nand I_42414 (I723584,I723567,I402737);
nor I_42415 (I723601,I723550,I723584);
DFFARX1 I_42416 (I723601,I2507,I723403,I723368,);
not I_42417 (I723632,I723584);
nand I_42418 (I723649,I723454,I723632);
nand I_42419 (I723380,I723516,I723632);
DFFARX1 I_42420 (I723550,I2507,I723403,I723395,);
not I_42421 (I723694,I402734);
nor I_42422 (I723711,I723694,I402749);
nor I_42423 (I723728,I723711,I723533);
DFFARX1 I_42424 (I723728,I2507,I723403,I723392,);
not I_42425 (I723759,I723711);
DFFARX1 I_42426 (I723759,I2507,I723403,I723785,);
not I_42427 (I723793,I723785);
nor I_42428 (I723389,I723793,I723711);
nor I_42429 (I723824,I723694,I402746);
and I_42430 (I723841,I723824,I402755);
or I_42431 (I723858,I723841,I402731);
DFFARX1 I_42432 (I723858,I2507,I723403,I723884,);
not I_42433 (I723892,I723884);
nand I_42434 (I723909,I723892,I723632);
not I_42435 (I723383,I723909);
nand I_42436 (I723377,I723909,I723649);
nand I_42437 (I723374,I723892,I723516);
not I_42438 (I723998,I2514);
DFFARX1 I_42439 (I440242,I2507,I723998,I724024,);
DFFARX1 I_42440 (I440239,I2507,I723998,I724041,);
not I_42441 (I724049,I724041);
nor I_42442 (I723966,I724024,I724049);
DFFARX1 I_42443 (I724049,I2507,I723998,I723981,);
nor I_42444 (I724094,I440254,I440236);
and I_42445 (I724111,I724094,I440233);
nor I_42446 (I724128,I724111,I440254);
not I_42447 (I724145,I440254);
and I_42448 (I724162,I724145,I440239);
nand I_42449 (I724179,I724162,I440251);
nor I_42450 (I724196,I724145,I724179);
DFFARX1 I_42451 (I724196,I2507,I723998,I723963,);
not I_42452 (I724227,I724179);
nand I_42453 (I724244,I724049,I724227);
nand I_42454 (I723975,I724111,I724227);
DFFARX1 I_42455 (I724145,I2507,I723998,I723990,);
not I_42456 (I724289,I440245);
nor I_42457 (I724306,I724289,I440239);
nor I_42458 (I724323,I724306,I724128);
DFFARX1 I_42459 (I724323,I2507,I723998,I723987,);
not I_42460 (I724354,I724306);
DFFARX1 I_42461 (I724354,I2507,I723998,I724380,);
not I_42462 (I724388,I724380);
nor I_42463 (I723984,I724388,I724306);
nor I_42464 (I724419,I724289,I440233);
and I_42465 (I724436,I724419,I440248);
or I_42466 (I724453,I724436,I440236);
DFFARX1 I_42467 (I724453,I2507,I723998,I724479,);
not I_42468 (I724487,I724479);
nand I_42469 (I724504,I724487,I724227);
not I_42470 (I723978,I724504);
nand I_42471 (I723972,I724504,I724244);
nand I_42472 (I723969,I724487,I724111);
not I_42473 (I724593,I2514);
DFFARX1 I_42474 (I548093,I2507,I724593,I724619,);
DFFARX1 I_42475 (I548084,I2507,I724593,I724636,);
not I_42476 (I724644,I724636);
nor I_42477 (I724561,I724619,I724644);
DFFARX1 I_42478 (I724644,I2507,I724593,I724576,);
nor I_42479 (I724689,I548090,I548099);
and I_42480 (I724706,I724689,I548102);
nor I_42481 (I724723,I724706,I548090);
not I_42482 (I724740,I548090);
and I_42483 (I724757,I724740,I548081);
nand I_42484 (I724774,I724757,I548087);
nor I_42485 (I724791,I724740,I724774);
DFFARX1 I_42486 (I724791,I2507,I724593,I724558,);
not I_42487 (I724822,I724774);
nand I_42488 (I724839,I724644,I724822);
nand I_42489 (I724570,I724706,I724822);
DFFARX1 I_42490 (I724740,I2507,I724593,I724585,);
not I_42491 (I724884,I548096);
nor I_42492 (I724901,I724884,I548081);
nor I_42493 (I724918,I724901,I724723);
DFFARX1 I_42494 (I724918,I2507,I724593,I724582,);
not I_42495 (I724949,I724901);
DFFARX1 I_42496 (I724949,I2507,I724593,I724975,);
not I_42497 (I724983,I724975);
nor I_42498 (I724579,I724983,I724901);
nor I_42499 (I725014,I724884,I548081);
and I_42500 (I725031,I725014,I548084);
or I_42501 (I725048,I725031,I548087);
DFFARX1 I_42502 (I725048,I2507,I724593,I725074,);
not I_42503 (I725082,I725074);
nand I_42504 (I725099,I725082,I724822);
not I_42505 (I724573,I725099);
nand I_42506 (I724567,I725099,I724839);
nand I_42507 (I724564,I725082,I724706);
not I_42508 (I725188,I2514);
DFFARX1 I_42509 (I414890,I2507,I725188,I725214,);
DFFARX1 I_42510 (I414872,I2507,I725188,I725231,);
not I_42511 (I725239,I725231);
nor I_42512 (I725156,I725214,I725239);
DFFARX1 I_42513 (I725239,I2507,I725188,I725171,);
nor I_42514 (I725284,I414878,I414881);
and I_42515 (I725301,I725284,I414869);
nor I_42516 (I725318,I725301,I414878);
not I_42517 (I725335,I414878);
and I_42518 (I725352,I725335,I414887);
nand I_42519 (I725369,I725352,I414875);
nor I_42520 (I725386,I725335,I725369);
DFFARX1 I_42521 (I725386,I2507,I725188,I725153,);
not I_42522 (I725417,I725369);
nand I_42523 (I725434,I725239,I725417);
nand I_42524 (I725165,I725301,I725417);
DFFARX1 I_42525 (I725335,I2507,I725188,I725180,);
not I_42526 (I725479,I414872);
nor I_42527 (I725496,I725479,I414887);
nor I_42528 (I725513,I725496,I725318);
DFFARX1 I_42529 (I725513,I2507,I725188,I725177,);
not I_42530 (I725544,I725496);
DFFARX1 I_42531 (I725544,I2507,I725188,I725570,);
not I_42532 (I725578,I725570);
nor I_42533 (I725174,I725578,I725496);
nor I_42534 (I725609,I725479,I414884);
and I_42535 (I725626,I725609,I414893);
or I_42536 (I725643,I725626,I414869);
DFFARX1 I_42537 (I725643,I2507,I725188,I725669,);
not I_42538 (I725677,I725669);
nand I_42539 (I725694,I725677,I725417);
not I_42540 (I725168,I725694);
nand I_42541 (I725162,I725694,I725434);
nand I_42542 (I725159,I725677,I725301);
not I_42543 (I725783,I2514);
DFFARX1 I_42544 (I453944,I2507,I725783,I725809,);
DFFARX1 I_42545 (I453941,I2507,I725783,I725826,);
not I_42546 (I725834,I725826);
nor I_42547 (I725751,I725809,I725834);
DFFARX1 I_42548 (I725834,I2507,I725783,I725766,);
nor I_42549 (I725879,I453956,I453938);
and I_42550 (I725896,I725879,I453935);
nor I_42551 (I725913,I725896,I453956);
not I_42552 (I725930,I453956);
and I_42553 (I725947,I725930,I453941);
nand I_42554 (I725964,I725947,I453953);
nor I_42555 (I725981,I725930,I725964);
DFFARX1 I_42556 (I725981,I2507,I725783,I725748,);
not I_42557 (I726012,I725964);
nand I_42558 (I726029,I725834,I726012);
nand I_42559 (I725760,I725896,I726012);
DFFARX1 I_42560 (I725930,I2507,I725783,I725775,);
not I_42561 (I726074,I453947);
nor I_42562 (I726091,I726074,I453941);
nor I_42563 (I726108,I726091,I725913);
DFFARX1 I_42564 (I726108,I2507,I725783,I725772,);
not I_42565 (I726139,I726091);
DFFARX1 I_42566 (I726139,I2507,I725783,I726165,);
not I_42567 (I726173,I726165);
nor I_42568 (I725769,I726173,I726091);
nor I_42569 (I726204,I726074,I453935);
and I_42570 (I726221,I726204,I453950);
or I_42571 (I726238,I726221,I453938);
DFFARX1 I_42572 (I726238,I2507,I725783,I726264,);
not I_42573 (I726272,I726264);
nand I_42574 (I726289,I726272,I726012);
not I_42575 (I725763,I726289);
nand I_42576 (I725757,I726289,I726029);
nand I_42577 (I725754,I726272,I725896);
not I_42578 (I726378,I2514);
DFFARX1 I_42579 (I682705,I2507,I726378,I726404,);
DFFARX1 I_42580 (I682696,I2507,I726378,I726421,);
not I_42581 (I726429,I726421);
nor I_42582 (I726346,I726404,I726429);
DFFARX1 I_42583 (I726429,I2507,I726378,I726361,);
nor I_42584 (I726474,I682687,I682702);
and I_42585 (I726491,I726474,I682690);
nor I_42586 (I726508,I726491,I682687);
not I_42587 (I726525,I682687);
and I_42588 (I726542,I726525,I682693);
nand I_42589 (I726559,I726542,I682711);
nor I_42590 (I726576,I726525,I726559);
DFFARX1 I_42591 (I726576,I2507,I726378,I726343,);
not I_42592 (I726607,I726559);
nand I_42593 (I726624,I726429,I726607);
nand I_42594 (I726355,I726491,I726607);
DFFARX1 I_42595 (I726525,I2507,I726378,I726370,);
not I_42596 (I726669,I682687);
nor I_42597 (I726686,I726669,I682693);
nor I_42598 (I726703,I726686,I726508);
DFFARX1 I_42599 (I726703,I2507,I726378,I726367,);
not I_42600 (I726734,I726686);
DFFARX1 I_42601 (I726734,I2507,I726378,I726760,);
not I_42602 (I726768,I726760);
nor I_42603 (I726364,I726768,I726686);
nor I_42604 (I726799,I726669,I682690);
and I_42605 (I726816,I726799,I682699);
or I_42606 (I726833,I726816,I682708);
DFFARX1 I_42607 (I726833,I2507,I726378,I726859,);
not I_42608 (I726867,I726859);
nand I_42609 (I726884,I726867,I726607);
not I_42610 (I726358,I726884);
nand I_42611 (I726352,I726884,I726624);
nand I_42612 (I726349,I726867,I726491);
not I_42613 (I726973,I2514);
DFFARX1 I_42614 (I43593,I2507,I726973,I726999,);
DFFARX1 I_42615 (I43581,I2507,I726973,I727016,);
not I_42616 (I727024,I727016);
nor I_42617 (I726941,I726999,I727024);
DFFARX1 I_42618 (I727024,I2507,I726973,I726956,);
nor I_42619 (I727069,I43572,I43596);
and I_42620 (I727086,I727069,I43575);
nor I_42621 (I727103,I727086,I43572);
not I_42622 (I727120,I43572);
and I_42623 (I727137,I727120,I43578);
nand I_42624 (I727154,I727137,I43590);
nor I_42625 (I727171,I727120,I727154);
DFFARX1 I_42626 (I727171,I2507,I726973,I726938,);
not I_42627 (I727202,I727154);
nand I_42628 (I727219,I727024,I727202);
nand I_42629 (I726950,I727086,I727202);
DFFARX1 I_42630 (I727120,I2507,I726973,I726965,);
not I_42631 (I727264,I43572);
nor I_42632 (I727281,I727264,I43578);
nor I_42633 (I727298,I727281,I727103);
DFFARX1 I_42634 (I727298,I2507,I726973,I726962,);
not I_42635 (I727329,I727281);
DFFARX1 I_42636 (I727329,I2507,I726973,I727355,);
not I_42637 (I727363,I727355);
nor I_42638 (I726959,I727363,I727281);
nor I_42639 (I727394,I727264,I43575);
and I_42640 (I727411,I727394,I43584);
or I_42641 (I727428,I727411,I43587);
DFFARX1 I_42642 (I727428,I2507,I726973,I727454,);
not I_42643 (I727462,I727454);
nand I_42644 (I727479,I727462,I727202);
not I_42645 (I726953,I727479);
nand I_42646 (I726947,I727479,I727219);
nand I_42647 (I726944,I727462,I727086);
not I_42648 (I727568,I2514);
DFFARX1 I_42649 (I524168,I2507,I727568,I727594,);
DFFARX1 I_42650 (I524186,I2507,I727568,I727611,);
not I_42651 (I727619,I727611);
nor I_42652 (I727536,I727594,I727619);
DFFARX1 I_42653 (I727619,I2507,I727568,I727551,);
nor I_42654 (I727664,I524165,I524177);
and I_42655 (I727681,I727664,I524162);
nor I_42656 (I727698,I727681,I524165);
not I_42657 (I727715,I524165);
and I_42658 (I727732,I727715,I524171);
nand I_42659 (I727749,I727732,I524183);
nor I_42660 (I727766,I727715,I727749);
DFFARX1 I_42661 (I727766,I2507,I727568,I727533,);
not I_42662 (I727797,I727749);
nand I_42663 (I727814,I727619,I727797);
nand I_42664 (I727545,I727681,I727797);
DFFARX1 I_42665 (I727715,I2507,I727568,I727560,);
not I_42666 (I727859,I524174);
nor I_42667 (I727876,I727859,I524171);
nor I_42668 (I727893,I727876,I727698);
DFFARX1 I_42669 (I727893,I2507,I727568,I727557,);
not I_42670 (I727924,I727876);
DFFARX1 I_42671 (I727924,I2507,I727568,I727950,);
not I_42672 (I727958,I727950);
nor I_42673 (I727554,I727958,I727876);
nor I_42674 (I727989,I727859,I524162);
and I_42675 (I728006,I727989,I524189);
or I_42676 (I728023,I728006,I524180);
DFFARX1 I_42677 (I728023,I2507,I727568,I728049,);
not I_42678 (I728057,I728049);
nand I_42679 (I728074,I728057,I727797);
not I_42680 (I727548,I728074);
nand I_42681 (I727542,I728074,I727814);
nand I_42682 (I727539,I728057,I727681);
not I_42683 (I728163,I2514);
DFFARX1 I_42684 (I203291,I2507,I728163,I728189,);
DFFARX1 I_42685 (I203285,I2507,I728163,I728206,);
not I_42686 (I728214,I728206);
nor I_42687 (I728131,I728189,I728214);
DFFARX1 I_42688 (I728214,I2507,I728163,I728146,);
nor I_42689 (I728259,I203273,I203294);
and I_42690 (I728276,I728259,I203288);
nor I_42691 (I728293,I728276,I203273);
not I_42692 (I728310,I203273);
and I_42693 (I728327,I728310,I203270);
nand I_42694 (I728344,I728327,I203282);
nor I_42695 (I728361,I728310,I728344);
DFFARX1 I_42696 (I728361,I2507,I728163,I728128,);
not I_42697 (I728392,I728344);
nand I_42698 (I728409,I728214,I728392);
nand I_42699 (I728140,I728276,I728392);
DFFARX1 I_42700 (I728310,I2507,I728163,I728155,);
not I_42701 (I728454,I203297);
nor I_42702 (I728471,I728454,I203270);
nor I_42703 (I728488,I728471,I728293);
DFFARX1 I_42704 (I728488,I2507,I728163,I728152,);
not I_42705 (I728519,I728471);
DFFARX1 I_42706 (I728519,I2507,I728163,I728545,);
not I_42707 (I728553,I728545);
nor I_42708 (I728149,I728553,I728471);
nor I_42709 (I728584,I728454,I203279);
and I_42710 (I728601,I728584,I203276);
or I_42711 (I728618,I728601,I203270);
DFFARX1 I_42712 (I728618,I2507,I728163,I728644,);
not I_42713 (I728652,I728644);
nand I_42714 (I728669,I728652,I728392);
not I_42715 (I728143,I728669);
nand I_42716 (I728137,I728669,I728409);
nand I_42717 (I728134,I728652,I728276);
not I_42718 (I728758,I2514);
DFFARX1 I_42719 (I553142,I2507,I728758,I728784,);
DFFARX1 I_42720 (I553133,I2507,I728758,I728801,);
not I_42721 (I728809,I728801);
nor I_42722 (I728726,I728784,I728809);
DFFARX1 I_42723 (I728809,I2507,I728758,I728741,);
nor I_42724 (I728854,I553139,I553148);
and I_42725 (I728871,I728854,I553151);
nor I_42726 (I728888,I728871,I553139);
not I_42727 (I728905,I553139);
and I_42728 (I728922,I728905,I553130);
nand I_42729 (I728939,I728922,I553136);
nor I_42730 (I728956,I728905,I728939);
DFFARX1 I_42731 (I728956,I2507,I728758,I728723,);
not I_42732 (I728987,I728939);
nand I_42733 (I729004,I728809,I728987);
nand I_42734 (I728735,I728871,I728987);
DFFARX1 I_42735 (I728905,I2507,I728758,I728750,);
not I_42736 (I729049,I553145);
nor I_42737 (I729066,I729049,I553130);
nor I_42738 (I729083,I729066,I728888);
DFFARX1 I_42739 (I729083,I2507,I728758,I728747,);
not I_42740 (I729114,I729066);
DFFARX1 I_42741 (I729114,I2507,I728758,I729140,);
not I_42742 (I729148,I729140);
nor I_42743 (I728744,I729148,I729066);
nor I_42744 (I729179,I729049,I553130);
and I_42745 (I729196,I729179,I553133);
or I_42746 (I729213,I729196,I553136);
DFFARX1 I_42747 (I729213,I2507,I728758,I729239,);
not I_42748 (I729247,I729239);
nand I_42749 (I729264,I729247,I728987);
not I_42750 (I728738,I729264);
nand I_42751 (I728732,I729264,I729004);
nand I_42752 (I728729,I729247,I728871);
not I_42753 (I729353,I2514);
DFFARX1 I_42754 (I115754,I2507,I729353,I729379,);
DFFARX1 I_42755 (I115757,I2507,I729353,I729396,);
not I_42756 (I729404,I729396);
nor I_42757 (I729321,I729379,I729404);
DFFARX1 I_42758 (I729404,I2507,I729353,I729336,);
nor I_42759 (I729449,I115763,I115757);
and I_42760 (I729466,I729449,I115760);
nor I_42761 (I729483,I729466,I115763);
not I_42762 (I729500,I115763);
and I_42763 (I729517,I729500,I115754);
nand I_42764 (I729534,I729517,I115772);
nor I_42765 (I729551,I729500,I729534);
DFFARX1 I_42766 (I729551,I2507,I729353,I729318,);
not I_42767 (I729582,I729534);
nand I_42768 (I729599,I729404,I729582);
nand I_42769 (I729330,I729466,I729582);
DFFARX1 I_42770 (I729500,I2507,I729353,I729345,);
not I_42771 (I729644,I115766);
nor I_42772 (I729661,I729644,I115754);
nor I_42773 (I729678,I729661,I729483);
DFFARX1 I_42774 (I729678,I2507,I729353,I729342,);
not I_42775 (I729709,I729661);
DFFARX1 I_42776 (I729709,I2507,I729353,I729735,);
not I_42777 (I729743,I729735);
nor I_42778 (I729339,I729743,I729661);
nor I_42779 (I729774,I729644,I115769);
and I_42780 (I729791,I729774,I115775);
or I_42781 (I729808,I729791,I115778);
DFFARX1 I_42782 (I729808,I2507,I729353,I729834,);
not I_42783 (I729842,I729834);
nand I_42784 (I729859,I729842,I729582);
not I_42785 (I729333,I729859);
nand I_42786 (I729327,I729859,I729599);
nand I_42787 (I729324,I729842,I729466);
not I_42788 (I729948,I2514);
DFFARX1 I_42789 (I101474,I2507,I729948,I729974,);
DFFARX1 I_42790 (I101477,I2507,I729948,I729991,);
not I_42791 (I729999,I729991);
nor I_42792 (I729916,I729974,I729999);
DFFARX1 I_42793 (I729999,I2507,I729948,I729931,);
nor I_42794 (I730044,I101483,I101477);
and I_42795 (I730061,I730044,I101480);
nor I_42796 (I730078,I730061,I101483);
not I_42797 (I730095,I101483);
and I_42798 (I730112,I730095,I101474);
nand I_42799 (I730129,I730112,I101492);
nor I_42800 (I730146,I730095,I730129);
DFFARX1 I_42801 (I730146,I2507,I729948,I729913,);
not I_42802 (I730177,I730129);
nand I_42803 (I730194,I729999,I730177);
nand I_42804 (I729925,I730061,I730177);
DFFARX1 I_42805 (I730095,I2507,I729948,I729940,);
not I_42806 (I730239,I101486);
nor I_42807 (I730256,I730239,I101474);
nor I_42808 (I730273,I730256,I730078);
DFFARX1 I_42809 (I730273,I2507,I729948,I729937,);
not I_42810 (I730304,I730256);
DFFARX1 I_42811 (I730304,I2507,I729948,I730330,);
not I_42812 (I730338,I730330);
nor I_42813 (I729934,I730338,I730256);
nor I_42814 (I730369,I730239,I101489);
and I_42815 (I730386,I730369,I101495);
or I_42816 (I730403,I730386,I101498);
DFFARX1 I_42817 (I730403,I2507,I729948,I730429,);
not I_42818 (I730437,I730429);
nand I_42819 (I730454,I730437,I730177);
not I_42820 (I729928,I730454);
nand I_42821 (I729922,I730454,I730194);
nand I_42822 (I729919,I730437,I730061);
not I_42823 (I730543,I2514);
DFFARX1 I_42824 (I212777,I2507,I730543,I730569,);
DFFARX1 I_42825 (I212771,I2507,I730543,I730586,);
not I_42826 (I730594,I730586);
nor I_42827 (I730511,I730569,I730594);
DFFARX1 I_42828 (I730594,I2507,I730543,I730526,);
nor I_42829 (I730639,I212759,I212780);
and I_42830 (I730656,I730639,I212774);
nor I_42831 (I730673,I730656,I212759);
not I_42832 (I730690,I212759);
and I_42833 (I730707,I730690,I212756);
nand I_42834 (I730724,I730707,I212768);
nor I_42835 (I730741,I730690,I730724);
DFFARX1 I_42836 (I730741,I2507,I730543,I730508,);
not I_42837 (I730772,I730724);
nand I_42838 (I730789,I730594,I730772);
nand I_42839 (I730520,I730656,I730772);
DFFARX1 I_42840 (I730690,I2507,I730543,I730535,);
not I_42841 (I730834,I212783);
nor I_42842 (I730851,I730834,I212756);
nor I_42843 (I730868,I730851,I730673);
DFFARX1 I_42844 (I730868,I2507,I730543,I730532,);
not I_42845 (I730899,I730851);
DFFARX1 I_42846 (I730899,I2507,I730543,I730925,);
not I_42847 (I730933,I730925);
nor I_42848 (I730529,I730933,I730851);
nor I_42849 (I730964,I730834,I212765);
and I_42850 (I730981,I730964,I212762);
or I_42851 (I730998,I730981,I212756);
DFFARX1 I_42852 (I730998,I2507,I730543,I731024,);
not I_42853 (I731032,I731024);
nand I_42854 (I731049,I731032,I730772);
not I_42855 (I730523,I731049);
nand I_42856 (I730517,I731049,I730789);
nand I_42857 (I730514,I731032,I730656);
not I_42858 (I731138,I2514);
DFFARX1 I_42859 (I145504,I2507,I731138,I731164,);
DFFARX1 I_42860 (I145507,I2507,I731138,I731181,);
not I_42861 (I731189,I731181);
nor I_42862 (I731106,I731164,I731189);
DFFARX1 I_42863 (I731189,I2507,I731138,I731121,);
nor I_42864 (I731234,I145513,I145507);
and I_42865 (I731251,I731234,I145510);
nor I_42866 (I731268,I731251,I145513);
not I_42867 (I731285,I145513);
and I_42868 (I731302,I731285,I145504);
nand I_42869 (I731319,I731302,I145522);
nor I_42870 (I731336,I731285,I731319);
DFFARX1 I_42871 (I731336,I2507,I731138,I731103,);
not I_42872 (I731367,I731319);
nand I_42873 (I731384,I731189,I731367);
nand I_42874 (I731115,I731251,I731367);
DFFARX1 I_42875 (I731285,I2507,I731138,I731130,);
not I_42876 (I731429,I145516);
nor I_42877 (I731446,I731429,I145504);
nor I_42878 (I731463,I731446,I731268);
DFFARX1 I_42879 (I731463,I2507,I731138,I731127,);
not I_42880 (I731494,I731446);
DFFARX1 I_42881 (I731494,I2507,I731138,I731520,);
not I_42882 (I731528,I731520);
nor I_42883 (I731124,I731528,I731446);
nor I_42884 (I731559,I731429,I145519);
and I_42885 (I731576,I731559,I145525);
or I_42886 (I731593,I731576,I145528);
DFFARX1 I_42887 (I731593,I2507,I731138,I731619,);
not I_42888 (I731627,I731619);
nand I_42889 (I731644,I731627,I731367);
not I_42890 (I731118,I731644);
nand I_42891 (I731112,I731644,I731384);
nand I_42892 (I731109,I731627,I731251);
not I_42893 (I731733,I2514);
DFFARX1 I_42894 (I511248,I2507,I731733,I731759,);
DFFARX1 I_42895 (I511266,I2507,I731733,I731776,);
not I_42896 (I731784,I731776);
nor I_42897 (I731701,I731759,I731784);
DFFARX1 I_42898 (I731784,I2507,I731733,I731716,);
nor I_42899 (I731829,I511245,I511257);
and I_42900 (I731846,I731829,I511242);
nor I_42901 (I731863,I731846,I511245);
not I_42902 (I731880,I511245);
and I_42903 (I731897,I731880,I511251);
nand I_42904 (I731914,I731897,I511263);
nor I_42905 (I731931,I731880,I731914);
DFFARX1 I_42906 (I731931,I2507,I731733,I731698,);
not I_42907 (I731962,I731914);
nand I_42908 (I731979,I731784,I731962);
nand I_42909 (I731710,I731846,I731962);
DFFARX1 I_42910 (I731880,I2507,I731733,I731725,);
not I_42911 (I732024,I511254);
nor I_42912 (I732041,I732024,I511251);
nor I_42913 (I732058,I732041,I731863);
DFFARX1 I_42914 (I732058,I2507,I731733,I731722,);
not I_42915 (I732089,I732041);
DFFARX1 I_42916 (I732089,I2507,I731733,I732115,);
not I_42917 (I732123,I732115);
nor I_42918 (I731719,I732123,I732041);
nor I_42919 (I732154,I732024,I511242);
and I_42920 (I732171,I732154,I511269);
or I_42921 (I732188,I732171,I511260);
DFFARX1 I_42922 (I732188,I2507,I731733,I732214,);
not I_42923 (I732222,I732214);
nand I_42924 (I732239,I732222,I731962);
not I_42925 (I731713,I732239);
nand I_42926 (I731707,I732239,I731979);
nand I_42927 (I731704,I732222,I731846);
endmodule


