// Verilog
// c2670
// Ninputs 157
// Noutputs 64
// NtotalGates 1193

module c2670(G1,G10,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G11,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G12,G120,G121,G122,G123,G124,G125,G126,G127,G128,G129,G13,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G14,G140,G141,G142,G143,G144,G145,G146,G147,G148,G149,G15,G150,G151,G152,G153,G154,G155,G156,G157,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,G2541,G2542,G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,G2555,G2556,G2557,G2558,G2559,G2560,G2561,G2562,G2563,G2564,G2565,G2566,G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,G2579,G2580,G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,G2591,G2592,G2593,G2594,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G5,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G6,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G7,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G8,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,G9,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G120,G121,G122,G123,G124,G125,G126,G127,G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,G141,G142,G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157;
output G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,G2541,G2542,G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,G2555,G2556,G2557,G2558,G2559,G2560,G2561,G2562,G2563,G2564,G2565,G2566,G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,G2579,G2580,G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,G2591,G2592,G2593,G2594;

wire G282,G283,G284,G285,G286,G287,G288,G291,G292,G295,G298,G301,G313,G325,G329,G335,G336,G339,G342,G354,G366,G370,G374,G386,G398,G399,G400,G401,G402,G403,G404,G405,G417,G429,G435,G442,G443,G447,G451,G455,G459,G463,G467,G471,G475,G479,G485,G491,G497,G503,G507,G511,G515,G519,G522,G525,G526,G527,G530,G533,G536,G539,G542,G545,G548,G551,G554,G557,G560,G563,G566,G569,G572,G575,G578,G581,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G598,G603,G614,G625,G626,G627,G628,G629,G630,G631,G636,G647,G658,G659,G660,G661,G662,G663,G674,G685,G686,G687,G688,G689,G690,G694,G698,G701,G702,G703,G704,G705,G706,G707,G718,G729,G730,G731,G732,G733,G734,G739,G745,G746,G747,G748,G749,G750,G751,G756,G761,G766,G771,G772,G773,G774,G775,G776,G777,G780,G783,G786,G789,G792,G795,G798,G801,G804,G807,G810,G811,G812,G815,G818,G821,G824,G827,G830,G831,G832,G833,G834,G835,G836,G837,G838,G839,G840,G841,G842,G843,G844,G845,G846,G847,G848,G849,G850,G851,G852,G853,G854,G855,G856,G857,G858,G859,G860,G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,G874,G875,G876,G877,G878,G879,G880,G881,G882,G883,G884,G885,G886,G887,G888,G889,G890,G891,G892,G893,G894,G895,G896,G897,G898,G901,G904,G908,G912,G915,G918,G921,G922,G923,G924,G925,G926,G927,G928,G929,G930,G931,G932,G933,G934,G935,G936,G937,G938,G939,G940,G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,G959,G963,G966,G967,G968,G969,G970,G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,G983,G984,G987,G990,G993,G998,G1002,G1008,G1014,G1017,G1021,G1026,G1030,G1033,G1036,G1039,G1044,G1049,G1053,G1058,G1062,G1067,G1072,G1076,G1079,G1082,G1085,G1088,G1089,G1090,G1093,G1096,G1097,G1098,G1101,G1104,G1107,G1110,G1111,G1112,G1113,G1114,G1115,G1116,G1117,G1118,G1119,G1120,G1123,G1126,G1127,G1128,G1129,G1132,G1137,G1144,G1148,G1152,G1159,G1166,G1171,G1176,G1181,G1184,G1187,G1190,G1193,G1196,G1197,G1198,G1199,G1200,G1201,G1202,G1203,G1204,G1205,G1206,G1207,G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1219,G1220,G1221,G1222,G1225,G1228,G1231,G1234,G1237,G1240,G1243,G1246,G1249,G1250,G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,G1263,G1266,G1269,G1272,G1275,G1278,G1281,G1284,G1287,G1290,G1293,G1296,G1299,G1302,G1305,G1308,G1311,G1314,G1320,G1321,G1326,G1327,G1328,G1329,G1336,G1342,G1345,G1348,G1351,G1354,G1355,G1356,G1357,G1358,G1359,G1360,G1361,G1362,G1363,G1364,G1365,G1366,G1367,G1368,G1371,G1374,G1377,G1380,G1383,G1384,G1387,G1390,G1393,G1396,G1399,G1402,G1405,G1406,G1407,G1408,G1409,G1412,G1415,G1418,G1421,G1424,G1425,G1426,G1427,G1428,G1429,G1430,G1431,G1432,G1433,G1434,G1435,G1436,G1437,G1438,G1439,G1440,G1441,G1442,G1443,G1444,G1445,G1446,G1447,G1448,G1449,G1450,G1451,G1452,G1453,G1454,G1455,G1456,G1457,G1458,G1459,G1460,G1461,G1462,G1463,G1464,G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1475,G1476,G1477,G1478,G1479,G1483,G1484,G1485,G1486,G1487,G1488,G1493,G1497,G1498,G1502,G1507,G1508,G1509,G1510,G1511,G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,G1524,G1528,G1531,G1532,G1533,G1534,G1535,G1536,G1537,G1540,G1543,G1546,G1549,G1552,G1555,G1556,G1557,G1560,G1563,G1566,G1569,G1572,G1575,G1578,G1581,G1584,G1587,G1590,G1593,G1596,G1599,G1600,G1601,G1602,G1603,G1606,G1607,G1610,G1613,G1616,G1619,G1620,G1621,G1622,G1623,G1624,G1625,G1626,G1627,G1628,G1629,G1630,G1631,G1632,G1633,G1634,G1635,G1636,G1640,G1641,G1642,G1643,G1644,G1645,G1646,G1650,G1651,G1652,G1653,G1654,G1657,G1661,G1662,G1663,G1664,G1665,G1666,G1667,G1668,G1669,G1670,G1675,G1676,G1681,G1682,G1683,G1684,G1688,G1689,G1690,G1691,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1700,G1701,G1702,G1703,G1704,G1705,G1706,G1709,G1712,G1715,G1718,G1719,G1720,G1721,G1722,G1723,G1724,G1725,G1726,G1727,G1728,G1731,G1732,G1733,G1734,G1735,G1736,G1737,G1738,G1739,G1744,G1749,G1750,G1751,G1752,G1753,G1754,G1755,G1756,G1761,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,G1774,G1775,G1776,G1777,G1778,G1779,G1780,G1781,G1782,G1785,G1789,G1792,G1795,G1798,G1799,G1800,G1801,G1802,G1805,G1811,G1814,G1815,G1816,G1822,G1823,G1824,G1825,G1826,G1829,G1835,G1840,G1846,G1851,G1854,G1857,G1858,G1859,G1862,G1865,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1878,G1879,G1880,G1881,G1882,G1883,G1884,G1887,G1888,G1889,G1890,G1893,G1896,G1899,G1902,G1903,G1904,G1907,G1910,G1913,G1916,G1919,G1922,G1925,G1926,G1927,G1928,G1931,G1934,G1937,G1940,G1943,G1946,G1947,G1948,G1953,G1954,G1955,G1956,G1961,G1962,G1963,G1964,G1965,G1966,G1967,G1970,G1971,G1972,G1973,G1974,G1975,G1976,G1977,G1978,G1981,G1982,G1983,G1984,G1985,G1986,G1987,G1988,G1989,G1990,G1991,G1992,G1993,G1996,G1999,G2002,G2005,G2008,G2011,G2014,G2017,G2020,G2023,G2026,G2029,G2032,G2035,G2038,G2041,G2044,G2045,G2046,G2047,G2048,G2051,G2052,G2053,G2054,G2055,G2056,G2057,G2058,G2059,G2060,G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071,G2072,G2073,G2076,G2079,G2082,G2085,G2088,G2091,G2094,G2097,G2100,G2103,G2106,G2109,G2112,G2115,G2116,G2117,G2118,G2119,G2120,G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,G2133,G2134,G2135,G2138,G2141,G2144,G2147,G2150,G2153,G2154,G2155,G2156,G2157,G2158,G2161,G2164,G2167,G2170,G2173,G2176,G2179,G2182,G2185,G2188,G2191,G2194,G2197,G2200,G2203,G2206,G2207,G2208,G2209,G2210,G2211,G2212,G2213,G2214,G2215,G2216,G2217,G2218,G2219,G2220,G2221,G2222,G2223,G2224,G2225,G2226,G2227,G2228,G2231,G2234,G2237,G2240,G2241,G2242,G2243,G2244,G2245,G2246,G2247,G2248,G2249,G2250,G2251,G2252,G2253,G2254,G2255,G2256,G2257,G2258,G2259,G2260,G2261,G2262,G2263,G2264,G2265,G2266,G2267,G2268,G2269,G2270,G2271,G2272,G2273,G2274,G2275,G2276,G2279,G2282,G2285,G2288,G2291,G2294,G2297,G2300,G2301,G2302,G2303,G2304,G2305,G2306,G2307,G2308,G2309,G2310,G2311,G2312,G2313,G2314,G2315,G2316,G2317,G2320,G2323,G2326,G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2340,G2345,G2349,G2352,G2353,G2359,G2364,G2365,G2366,G2367,G2368,G2369,G2370,G2375,G2379,G2382,G2383,G2389,G2394,G2395,G2396,G2397,G2398,G2399,G2400,G2401,G2402,G2403,G2404,G2405,G2406,G2407,G2408,G2409,G2410,G2411,G2412,G2413,G2414,G2417,G2418,G2419,G2420,G2421,G2422,G2423,G2424,G2425,G2426,G2427,G2428,G2431,G2432,G2433,G2434,G2435,G2436,G2437,G2438,G2439,G2440,G2441,G2442,G2443,G2447,G2450,G2451,G2454,G2458,G2461,G2462,G2465,G2466,G2467,G2470,G2473,G2474,G2475,G2476,G2477,G2478,G2479,G2480,G2481,G2482,G2483,G2484,G2485,G2486,G2487,G2488,G2489,G2490,G2491,G2492,G2495,G2496,G2499,G2500,G2501,G2502,G2503,G2504,G2505,G2508,G2512,G2515,G2516,G2517,G2520,G2523,G2524,G2527,G2528;

and AND2_0(G282,G1,G3);
not NOT_0(G283,G118);
not NOT_1(G284,G127);
and AND4_0(G285,G142,G141,G140,G139);
not NOT_2(G286,G282);
and AND3_0(G287,G2,G11,G121);
not NOT_3(G288,G121);
and AND2_1(G291,G29,G29);
not NOT_4(G292,G115);
not NOT_5(G295,G8);
not NOT_6(G298,G8);
not NOT_7(G301,G117);
not NOT_8(G313,G120);
not NOT_9(G325,G122);
not NOT_10(G329,G123);
and AND2_2(G335,G9,G123);
and AND4_1(G336,G106,G64,G76,G32);
and AND4_2(G339,G96,G43,G86,G53);
not NOT_11(G342,G117);
not NOT_12(G354,G120);
not NOT_13(G366,G125);
not NOT_14(G370,G126);
not NOT_15(G374,G145);
not NOT_16(G386,G146);
not NOT_17(G398,G148);
not NOT_18(G399,G149);
not NOT_19(G400,G150);
not NOT_20(G401,G151);
not NOT_21(G402,G152);
not NOT_22(G403,G153);
not NOT_23(G404,G156);
not NOT_24(G405,G145);
not NOT_25(G417,G146);
not NOT_26(G429,G12);
not NOT_27(G435,G12);
not NOT_28(G442,G157);
and AND2_3(G443,G7,G121);
not NOT_29(G447,G128);
not NOT_30(G451,G129);
not NOT_31(G455,G130);
not NOT_32(G459,G131);
not NOT_33(G463,G132);
not NOT_34(G467,G133);
not NOT_35(G471,G134);
not NOT_36(G475,G135);
not NOT_37(G479,G136);
not NOT_38(G485,G23);
not NOT_39(G491,G23);
not NOT_40(G497,G138);
not NOT_41(G503,G139);
not NOT_42(G507,G140);
not NOT_43(G511,G141);
not NOT_44(G515,G142);
not NOT_45(G519,G143);
not NOT_46(G522,G144);
not NOT_47(G525,G154);
not NOT_48(G526,G155);
not NOT_49(G527,G126);
not NOT_50(G530,G125);
not NOT_51(G533,G128);
not NOT_52(G536,G130);
not NOT_53(G539,G129);
not NOT_54(G542,G132);
not NOT_55(G545,G131);
not NOT_56(G548,G134);
not NOT_57(G551,G133);
not NOT_58(G554,G136);
not NOT_59(G557,G135);
not NOT_60(G560,G138);
not NOT_61(G563,G140);
not NOT_62(G566,G139);
not NOT_63(G569,G142);
not NOT_64(G572,G141);
not NOT_65(G575,G144);
not NOT_66(G578,G143);
not NOT_67(G581,G291);
nand NAND2_0(G584,G149,G398);
nand NAND2_1(G585,G148,G399);
nand NAND2_2(G586,G151,G400);
nand NAND2_3(G587,G150,G401);
nand NAND2_4(G588,G153,G402);
nand NAND2_5(G589,G152,G403);
nand NAND2_6(G590,G155,G525);
nand NAND2_7(G591,G154,G526);
and AND2_4(G592,G147,G443);
not NOT_68(G593,G336);
not NOT_69(G594,G339);
and AND2_5(G595,G339,G336);
not NOT_70(G598,G295);
not NOT_71(G603,G301);
not NOT_72(G614,G313);
and AND3_1(G625,G62,G301,G313);
and AND3_2(G626,G52,G301,G313);
and AND3_3(G627,G61,G301,G313);
and AND3_4(G628,G60,G301,G313);
and AND3_5(G629,G59,G301,G313);
and AND2_6(G630,G9,G329);
not NOT_73(G631,G295);
not NOT_74(G636,G342);
not NOT_75(G647,G354);
and AND3_6(G658,G58,G342,G354);
and AND3_7(G659,G57,G342,G354);
and AND3_8(G660,G56,G342,G354);
and AND3_9(G661,G55,G342,G354);
and AND3_10(G662,G54,G342,G354);
not NOT_76(G663,G374);
not NOT_77(G674,G386);
and AND3_11(G685,G90,G374,G386);
and AND3_12(G686,G89,G374,G386);
and AND3_13(G687,G88,G374,G386);
and AND3_14(G688,G87,G374,G386);
and AND2_7(G689,G374,G386);
nand NAND2_8(G690,G584,G585);
nand NAND2_9(G694,G586,G587);
nand NAND2_10(G698,G588,G589);
not NOT_78(G701,G533);
nand NAND2_11(G702,G533,G404);
not NOT_79(G703,G536);
not NOT_80(G704,G539);
not NOT_81(G705,G542);
not NOT_82(G706,G545);
not NOT_83(G707,G405);
not NOT_84(G718,G417);
and AND3_15(G729,G94,G405,G417);
and AND3_16(G730,G85,G405,G417);
and AND3_17(G731,G93,G405,G417);
and AND3_18(G732,G92,G405,G417);
and AND3_19(G733,G91,G405,G417);
not NOT_85(G734,G429);
not NOT_86(G739,G435);
not NOT_87(G745,G560);
nand NAND2_12(G746,G560,G442);
not NOT_88(G747,G563);
not NOT_89(G748,G566);
not NOT_90(G749,G569);
not NOT_91(G750,G572);
not NOT_92(G751,G298);
not NOT_93(G756,G298);
not NOT_94(G761,G485);
not NOT_95(G766,G491);
not NOT_96(G771,G527);
not NOT_97(G772,G530);
not NOT_98(G773,G548);
not NOT_99(G774,G551);
not NOT_100(G775,G554);
not NOT_101(G776,G557);
nand NAND2_13(G777,G590,G591);
not NOT_102(G780,G366);
not NOT_103(G783,G370);
not NOT_104(G786,G447);
not NOT_105(G789,G451);
not NOT_106(G792,G455);
not NOT_107(G795,G459);
not NOT_108(G798,G463);
not NOT_109(G801,G467);
not NOT_110(G804,G471);
not NOT_111(G807,G475);
not NOT_112(G810,G575);
not NOT_113(G811,G578);
not NOT_114(G812,G479);
not NOT_115(G815,G497);
not NOT_116(G818,G503);
not NOT_117(G821,G507);
not NOT_118(G824,G511);
not NOT_119(G827,G515);
and AND2_8(G830,G147,G593);
and AND2_9(G831,G119,G594);
or OR2_0(G832,G630,G335);
nand NAND2_14(G833,G156,G701);
nand NAND2_15(G834,G539,G703);
nand NAND2_16(G835,G536,G704);
nand NAND2_17(G836,G545,G705);
nand NAND2_18(G837,G542,G706);
nand NAND2_19(G838,G157,G745);
nand NAND2_20(G839,G566,G747);
nand NAND2_21(G840,G563,G748);
nand NAND2_22(G841,G572,G749);
nand NAND2_23(G842,G569,G750);
nand NAND2_24(G843,G530,G771);
nand NAND2_25(G844,G527,G772);
nand NAND2_26(G845,G551,G773);
nand NAND2_27(G846,G548,G774);
nand NAND2_28(G847,G557,G775);
nand NAND2_29(G848,G554,G776);
nand NAND2_30(G849,G578,G810);
nand NAND2_31(G850,G575,G811);
not NOT_120(G851,G830);
not NOT_121(G852,G831);
and AND3_20(G853,G73,G603,G614);
and AND3_21(G854,G41,G301,G614);
and AND3_22(G855,G51,G603,G313);
and AND3_23(G856,G63,G603,G614);
and AND3_24(G857,G31,G301,G614);
and AND3_25(G858,G42,G603,G313);
and AND3_26(G859,G72,G603,G614);
and AND3_27(G860,G40,G301,G614);
and AND3_28(G861,G50,G603,G313);
and AND3_29(G862,G71,G603,G614);
and AND3_30(G863,G39,G301,G614);
and AND3_31(G864,G49,G603,G313);
and AND3_32(G865,G70,G603,G614);
and AND3_33(G866,G38,G301,G614);
and AND3_34(G867,G48,G603,G313);
and AND3_35(G868,G69,G636,G647);
and AND3_36(G869,G37,G342,G647);
and AND3_37(G870,G47,G636,G354);
and AND3_38(G871,G68,G636,G647);
and AND3_39(G872,G36,G342,G647);
and AND3_40(G873,G46,G636,G354);
and AND3_41(G874,G67,G636,G647);
and AND3_42(G875,G35,G342,G647);
and AND2_10(G876,G636,G354);
and AND3_43(G877,G66,G636,G647);
and AND3_44(G878,G34,G342,G647);
and AND3_45(G879,G45,G636,G354);
and AND3_46(G880,G65,G636,G647);
and AND3_47(G881,G33,G342,G647);
and AND3_48(G882,G44,G636,G354);
and AND3_49(G883,G110,G663,G674);
and AND3_50(G884,G80,G374,G674);
and AND3_51(G885,G100,G663,G386);
and AND3_52(G886,G109,G663,G674);
and AND3_53(G887,G79,G374,G674);
and AND3_54(G888,G99,G663,G386);
and AND3_55(G889,G108,G663,G674);
and AND3_56(G890,G78,G374,G674);
and AND3_57(G891,G98,G663,G386);
and AND3_58(G892,G107,G663,G674);
and AND3_59(G893,G77,G374,G674);
and AND3_60(G894,G97,G663,G386);
and AND2_11(G895,G663,G674);
and AND2_12(G896,G374,G674);
and AND2_13(G897,G663,G386);
not NOT_122(G898,G690);
not NOT_123(G901,G694);
nand NAND2_32(G904,G833,G702);
nand NAND2_33(G908,G834,G835);
nand NAND2_34(G912,G836,G837);
not NOT_124(G915,G698);
not NOT_125(G918,G698);
not NOT_126(G921,G780);
not NOT_127(G922,G783);
not NOT_128(G923,G786);
not NOT_129(G924,G789);
not NOT_130(G925,G792);
not NOT_131(G926,G795);
not NOT_132(G927,G798);
not NOT_133(G928,G801);
not NOT_134(G929,G804);
not NOT_135(G930,G807);
and AND3_61(G931,G114,G707,G718);
and AND3_62(G932,G84,G405,G718);
and AND3_63(G933,G104,G707,G417);
and AND3_64(G934,G105,G707,G718);
and AND3_65(G935,G75,G405,G718);
and AND3_66(G936,G95,G707,G417);
and AND3_67(G937,G113,G707,G718);
and AND3_68(G938,G83,G405,G718);
and AND3_69(G939,G103,G707,G417);
and AND3_70(G940,G112,G707,G718);
and AND3_71(G941,G82,G405,G718);
and AND3_72(G942,G102,G707,G417);
and AND3_73(G943,G111,G707,G718);
and AND3_74(G944,G81,G405,G718);
and AND3_75(G945,G101,G707,G417);
and AND2_14(G946,G13,G734);
and AND2_15(G947,G4,G734);
and AND2_16(G948,G14,G734);
and AND2_17(G949,G5,G734);
and AND2_18(G950,G15,G739);
and AND2_19(G951,G16,G739);
and AND2_20(G952,G17,G739);
and AND2_21(G953,G6,G739);
and AND2_22(G954,G18,G739);
nand NAND2_35(G955,G838,G746);
nand NAND2_36(G959,G839,G840);
nand NAND2_37(G963,G841,G842);
and AND2_23(G966,G19,G761);
and AND2_24(G967,G24,G761);
and AND2_25(G968,G20,G761);
and AND2_26(G969,G25,G761);
and AND2_27(G970,G21,G766);
and AND2_28(G971,G26,G766);
and AND2_29(G972,G27,G766);
and AND2_30(G973,G22,G766);
not NOT_136(G974,G812);
not NOT_137(G975,G815);
not NOT_138(G976,G818);
not NOT_139(G977,G821);
not NOT_140(G978,G824);
not NOT_141(G979,G827);
nand NAND2_38(G980,G843,G844);
not NOT_142(G983,G777);
nand NAND2_39(G984,G847,G848);
nand NAND2_40(G987,G845,G846);
nand NAND2_41(G990,G849,G850);
and AND2_31(G993,G851,G852);
or OR4_0(G998,G853,G854,G855,G625);
or OR4_1(G1002,G856,G857,G858,G626);
or OR4_2(G1008,G859,G860,G861,G627);
or OR4_3(G1014,G862,G863,G864,G628);
or OR4_4(G1017,G865,G866,G867,G629);
or OR4_5(G1021,G868,G869,G870,G658);
or OR4_6(G1026,G871,G872,G873,G659);
or OR4_7(G1030,G874,G875,G876,G660);
or OR4_8(G1033,G877,G878,G879,G661);
or OR4_9(G1036,G880,G881,G882,G662);
or OR4_10(G1039,G883,G884,G885,G685);
or OR4_11(G1044,G886,G887,G888,G686);
or OR4_12(G1049,G889,G890,G891,G687);
or OR4_13(G1053,G892,G893,G894,G688);
or OR4_14(G1058,G895,G896,G897,G689);
or OR4_15(G1062,G934,G935,G936,G730);
or OR4_16(G1067,G937,G938,G939,G731);
or OR4_17(G1072,G940,G941,G942,G732);
or OR4_18(G1076,G943,G944,G945,G733);
or OR4_19(G1079,G931,G932,G933,G729);
not NOT_143(G1082,G904);
not NOT_144(G1085,G908);
not NOT_145(G1088,G915);
not NOT_146(G1089,G918);
not NOT_147(G1090,G912);
not NOT_148(G1093,G912);
and AND3_76(G1096,G694,G690,G915);
and AND3_77(G1097,G901,G898,G918);
not NOT_149(G1098,G955);
not NOT_150(G1101,G959);
not NOT_151(G1104,G963);
not NOT_152(G1107,G963);
not NOT_153(G1110,G990);
not NOT_154(G1111,G980);
nand NAND2_42(G1112,G980,G983);
not NOT_155(G1113,G984);
not NOT_156(G1114,G987);
and AND2_32(G1115,G998,G122);
and AND2_33(G1116,G1008,G122);
and AND2_34(G1117,G1002,G122);
and AND4_3(G1118,G288,G116,G28,G993);
and AND4_4(G1119,G288,G116,G993,G286);
not NOT_157(G1120,G998);
not NOT_158(G1123,G1008);
and AND2_35(G1126,G1002,G329);
and AND2_36(G1127,G1008,G329);
and AND2_37(G1128,G1021,G123);
not NOT_159(G1129,G998);
not NOT_160(G1132,G1002);
not NOT_161(G1137,G1008);
not NOT_162(G1144,G1014);
not NOT_163(G1148,G1017);
not NOT_164(G1152,G1021);
not NOT_165(G1159,G1026);
not NOT_166(G1166,G1030);
not NOT_167(G1171,G1033);
not NOT_168(G1176,G1036);
nand NAND2_43(G1181,G519,G1053);
nand NAND2_44(G1184,G522,G1058);
not NOT_169(G1187,G1072);
and AND2_38(G1190,G1039,G284);
not NOT_170(G1193,G1044);
and AND3_78(G1196,G898,G694,G1088);
and AND3_79(G1197,G690,G901,G1089);
and AND2_39(G1198,G1002,G429);
and AND2_40(G1199,G1008,G429);
and AND2_41(G1200,G1014,G429);
and AND2_42(G1201,G1017,G429);
and AND2_43(G1202,G1021,G435);
and AND2_44(G1203,G1026,G435);
and AND2_45(G1204,G1030,G435);
and AND2_46(G1205,G1033,G435);
and AND2_47(G1206,G1036,G435);
not NOT_171(G1207,G1079);
and AND2_48(G1208,G1062,G485);
and AND2_49(G1209,G1067,G485);
and AND2_50(G1210,G1072,G485);
and AND2_51(G1211,G1076,G485);
and AND2_52(G1212,G1039,G491);
and AND2_53(G1213,G1044,G491);
and AND2_54(G1214,G1049,G491);
and AND2_55(G1215,G1053,G491);
not NOT_172(G1216,G1002);
nand NAND2_45(G1219,G777,G1111);
nand NAND2_46(G1220,G987,G1113);
nand NAND2_47(G1221,G984,G1114);
not NOT_173(G1222,G1062);
not NOT_174(G1225,G1072);
not NOT_175(G1228,G1067);
not NOT_176(G1231,G1039);
not NOT_177(G1234,G1076);
not NOT_178(G1237,G1049);
not NOT_179(G1240,G1044);
not NOT_180(G1243,G1058);
not NOT_181(G1246,G1053);
not NOT_182(G1249,G1090);
not NOT_183(G1250,G1093);
nor NOR2_0(G1251,G1196,G1096);
nor NOR2_1(G1252,G1197,G1097);
and AND3_80(G1253,G908,G904,G1090);
and AND3_81(G1254,G1085,G1082,G1093);
or OR2_1(G1255,G973,G1215);
not NOT_184(G1256,G1104);
not NOT_185(G1257,G1107);
and AND3_82(G1258,G959,G955,G1104);
and AND3_83(G1259,G1101,G1098,G1107);
nand NAND2_48(G1260,G1219,G1112);
nand NAND2_49(G1263,G1220,G1221);
or OR2_2(G1266,G946,G1198);
or OR2_3(G1269,G947,G1199);
or OR2_4(G1272,G948,G1200);
or OR2_5(G1275,G949,G1201);
or OR2_6(G1278,G950,G1202);
or OR2_7(G1281,G951,G1203);
or OR2_8(G1284,G952,G1204);
or OR2_9(G1287,G953,G1205);
or OR2_10(G1290,G954,G1206);
or OR2_11(G1293,G966,G1208);
or OR2_12(G1296,G967,G1209);
or OR2_13(G1299,G968,G1210);
or OR2_14(G1302,G969,G1211);
or OR2_15(G1305,G970,G1212);
or OR2_16(G1308,G971,G1213);
or OR2_17(G1311,G972,G1214);
and AND3_84(G1314,G1193,G1190,G30);
not NOT_186(G1320,G1190);
nand NAND2_50(G1321,G283,G1123);
and AND2_56(G1326,G1120,G329);
and AND2_57(G1327,G1148,G123);
and AND2_58(G1328,G1144,G329);
not NOT_187(G1329,G1144);
not NOT_188(G1336,G1148);
not NOT_189(G1342,G1159);
not NOT_190(G1345,G1166);
not NOT_191(G1348,G1171);
not NOT_192(G1351,G1176);
and AND2_59(G1354,G519,G1181);
and AND2_60(G1355,G1181,G1053);
and AND2_61(G1356,G522,G1184);
and AND2_62(G1357,G1184,G1058);
and AND3_85(G1358,G1082,G908,G1249);
and AND3_86(G1359,G904,G1085,G1250);
not NOT_193(G1360,G1222);
nand NAND2_51(G1361,G1222,G1207);
not NOT_194(G1362,G1225);
not NOT_195(G1363,G1228);
not NOT_196(G1364,G1231);
not NOT_197(G1365,G1234);
and AND3_87(G1366,G1098,G959,G1256);
and AND3_88(G1367,G955,G1101,G1257);
not NOT_198(G1368,G1132);
not NOT_199(G1371,G1129);
not NOT_200(G1374,G1137);
not NOT_201(G1377,G1152);
not NOT_202(G1380,G1123);
not NOT_203(G1383,G1216);
not NOT_204(G1384,G1132);
not NOT_205(G1387,G1129);
not NOT_206(G1390,G1137);
not NOT_207(G1393,G1120);
not NOT_208(G1396,G1137);
not NOT_209(G1399,G1137);
nand NAND2_52(G1402,G1252,G1251);
not NOT_210(G1405,G1237);
not NOT_211(G1406,G1240);
not NOT_212(G1407,G1243);
not NOT_213(G1408,G1246);
and AND3_89(G1409,G30,G1193,G1320);
or OR2_18(G1412,G1127,G1327);
or OR2_19(G1415,G1328,G1128);
or OR2_20(G1418,G1354,G1355);
or OR2_21(G1421,G1356,G1357);
nor NOR2_2(G1424,G1358,G1253);
nor NOR2_3(G1425,G1359,G1254);
not NOT_214(G1426,G1260);
not NOT_215(G1427,G1263);
nand NAND2_53(G1428,G1266,G921);
not NOT_216(G1429,G1266);
nand NAND2_54(G1430,G1269,G922);
not NOT_217(G1431,G1269);
nand NAND2_55(G1432,G1272,G923);
not NOT_218(G1433,G1272);
nand NAND2_56(G1434,G1275,G924);
not NOT_219(G1435,G1275);
nand NAND2_57(G1436,G1278,G925);
not NOT_220(G1437,G1278);
nand NAND2_58(G1438,G1281,G926);
not NOT_221(G1439,G1281);
nand NAND2_59(G1440,G1284,G927);
not NOT_222(G1441,G1284);
nand NAND2_60(G1442,G1287,G928);
not NOT_223(G1443,G1287);
nand NAND2_61(G1444,G1290,G929);
not NOT_224(G1445,G1290);
nand NAND2_62(G1446,G1293,G930);
not NOT_225(G1447,G1293);
nand NAND2_63(G1448,G1079,G1360);
nand NAND2_64(G1449,G1228,G1362);
nand NAND2_65(G1450,G1225,G1363);
nand NAND2_66(G1451,G1234,G1364);
nand NAND2_67(G1452,G1231,G1365);
nor NOR2_4(G1453,G1366,G1258);
nor NOR2_5(G1454,G1367,G1259);
nand NAND2_68(G1455,G1296,G974);
not NOT_226(G1456,G1296);
nand NAND2_69(G1457,G1299,G975);
not NOT_227(G1458,G1299);
nand NAND2_70(G1459,G1302,G976);
not NOT_228(G1460,G1302);
nand NAND2_71(G1461,G1305,G977);
not NOT_229(G1462,G1305);
nand NAND2_72(G1463,G1308,G978);
not NOT_230(G1464,G1308);
nand NAND2_73(G1465,G1311,G979);
not NOT_231(G1466,G1311);
nand NAND2_74(G1467,G1240,G1405);
nand NAND2_75(G1468,G1237,G1406);
nand NAND2_76(G1469,G1246,G1407);
nand NAND2_77(G1470,G1243,G1408);
and AND2_63(G1471,G1321,G325);
not NOT_232(G1472,G1314);
not NOT_233(G1475,G1368);
not NOT_234(G1476,G1371);
not NOT_235(G1477,G1374);
not NOT_236(G1478,G1377);
not NOT_237(G1479,G1321);
not NOT_238(G1483,G1384);
not NOT_239(G1484,G1387);
not NOT_240(G1485,G1390);
not NOT_241(G1486,G1393);
not NOT_242(G1487,G1396);
not NOT_243(G1488,G1314);
not NOT_244(G1493,G1314);
and AND2_64(G1497,G1321,G123);
not NOT_245(G1498,G1314);
not NOT_246(G1502,G1314);
nand NAND2_78(G1507,G1402,G1426);
not NOT_247(G1508,G1399);
not NOT_248(G1509,G1402);
nand NAND2_79(G1510,G780,G1429);
nand NAND2_80(G1511,G783,G1431);
nand NAND2_81(G1512,G786,G1433);
nand NAND2_82(G1513,G789,G1435);
nand NAND2_83(G1514,G792,G1437);
nand NAND2_84(G1515,G795,G1439);
nand NAND2_85(G1516,G798,G1441);
nand NAND2_86(G1517,G801,G1443);
nand NAND2_87(G1518,G804,G1445);
nand NAND2_88(G1519,G807,G1447);
nand NAND2_89(G1520,G1448,G1361);
nand NAND2_90(G1524,G1449,G1450);
nand NAND2_91(G1528,G1451,G1452);
nand NAND2_92(G1531,G812,G1456);
nand NAND2_93(G1532,G815,G1458);
nand NAND2_94(G1533,G818,G1460);
nand NAND2_95(G1534,G821,G1462);
nand NAND2_96(G1535,G824,G1464);
nand NAND2_97(G1536,G827,G1466);
not NOT_249(G1537,G1329);
not NOT_250(G1540,G1336);
not NOT_251(G1543,G1345);
not NOT_252(G1546,G1342);
not NOT_253(G1549,G1351);
not NOT_254(G1552,G1348);
not NOT_255(G1555,G1380);
nand NAND2_98(G1556,G1380,G1383);
not NOT_256(G1557,G1329);
not NOT_257(G1560,G1345);
not NOT_258(G1563,G1342);
not NOT_259(G1566,G1351);
not NOT_260(G1569,G1348);
not NOT_261(G1572,G1321);
not NOT_262(G1575,G1329);
not NOT_263(G1578,G1336);
not NOT_264(G1581,G1329);
not NOT_265(G1584,G1336);
nand NAND2_99(G1587,G1425,G1424);
nand NAND2_100(G1590,G1469,G1470);
nand NAND2_101(G1593,G1467,G1468);
nand NAND2_102(G1596,G1454,G1453);
nand NAND2_103(G1599,G1371,G1475);
nand NAND2_104(G1600,G1368,G1476);
nand NAND2_105(G1601,G1387,G1483);
nand NAND2_106(G1602,G1384,G1484);
or OR2_22(G1603,G1126,G1497);
nand NAND2_107(G1606,G1260,G1509);
not NOT_266(G1607,G1418);
not NOT_267(G1610,G1421);
not NOT_268(G1613,G1409);
not NOT_269(G1616,G1409);
nand NAND2_108(G1619,G1428,G1510);
nand NAND2_109(G1620,G1430,G1511);
nand NAND2_110(G1621,G1432,G1512);
nand NAND2_111(G1622,G1434,G1513);
nand NAND2_112(G1623,G1436,G1514);
nand NAND2_113(G1624,G1438,G1515);
nand NAND2_114(G1625,G1440,G1516);
nand NAND2_115(G1626,G1442,G1517);
nand NAND2_116(G1627,G1444,G1518);
nand NAND2_117(G1628,G1446,G1519);
nand NAND2_118(G1629,G1455,G1531);
nand NAND2_119(G1630,G1457,G1532);
nand NAND2_120(G1631,G1459,G1533);
nand NAND2_121(G1632,G1461,G1534);
nand NAND2_122(G1633,G1463,G1535);
nand NAND2_123(G1634,G1465,G1536);
nand NAND2_124(G1635,G1216,G1555);
not NOT_270(G1636,G1472);
and AND2_65(G1640,G1176,G1488);
and AND2_66(G1641,G1062,G1488);
and AND2_67(G1642,G1067,G1488);
and AND2_68(G1643,G1187,G1488);
and AND2_69(G1644,G1152,G1493);
and AND2_70(G1645,G1159,G1493);
nand NAND2_125(G1646,G1599,G1600);
not NOT_271(G1650,G1537);
nand NAND2_126(G1651,G1537,G1477);
nand NAND2_127(G1652,G1540,G1478);
not NOT_272(G1653,G1540);
not NOT_273(G1654,G1479);
nand NAND2_128(G1657,G1601,G1602);
not NOT_274(G1661,G1557);
nand NAND2_129(G1662,G1557,G1485);
not NOT_275(G1663,G1575);
and AND2_71(G1664,G1152,G1498);
and AND2_72(G1665,G1159,G1498);
and AND2_73(G1666,G1176,G1502);
and AND2_74(G1667,G1062,G1502);
and AND2_75(G1668,G1067,G1502);
and AND2_76(G1669,G1187,G1502);
not NOT_276(G1670,G1493);
not NOT_277(G1675,G1578);
not NOT_278(G1676,G1498);
nand NAND2_130(G1681,G1606,G1507);
not NOT_279(G1682,G1581);
not NOT_280(G1683,G1584);
not NOT_281(G1684,G1472);
not NOT_282(G1688,G1587);
nand NAND2_131(G1689,G1587,G1427);
not NOT_283(G1690,G1628);
not NOT_284(G1691,G1627);
not NOT_285(G1692,G1626);
not NOT_286(G1693,G1625);
not NOT_287(G1694,G1624);
not NOT_288(G1695,G1623);
not NOT_289(G1696,G1622);
not NOT_290(G1697,G1621);
not NOT_291(G1698,G1620);
not NOT_292(G1699,G1619);
not NOT_293(G1700,G1634);
not NOT_294(G1701,G1633);
not NOT_295(G1702,G1632);
not NOT_296(G1703,G1631);
not NOT_297(G1704,G1630);
not NOT_298(G1705,G1629);
not NOT_299(G1706,G1520);
not NOT_300(G1709,G1524);
not NOT_301(G1712,G1528);
not NOT_302(G1715,G1528);
not NOT_303(G1718,G1596);
nand NAND2_132(G1719,G1596,G1110);
not NOT_304(G1720,G1543);
not NOT_305(G1721,G1546);
not NOT_306(G1722,G1549);
not NOT_307(G1723,G1552);
not NOT_308(G1724,G1560);
not NOT_309(G1725,G1563);
not NOT_310(G1726,G1566);
not NOT_311(G1727,G1569);
nand NAND2_133(G1728,G1635,G1556);
not NOT_312(G1731,G1572);
not NOT_313(G1732,G1590);
not NOT_314(G1733,G1593);
and AND2_77(G1734,G1421,G1610);
and AND2_78(G1735,G1418,G1607);
nand NAND2_134(G1736,G1374,G1650);
nand NAND2_135(G1737,G1377,G1653);
nand NAND2_136(G1738,G1390,G1661);
not NOT_315(G1739,G1613);
not NOT_316(G1744,G1613);
not NOT_317(G1749,G1681);
nand NAND2_137(G1750,G1263,G1688);
and AND5_0(G1751,G1690,G1691,G1692,G1693,G1694);
and AND5_1(G1752,G1695,G1696,G1697,G1698,G1699);
and AND2_79(G1753,G1255,G1700);
and AND5_2(G1754,G1701,G1702,G1703,G1704,G1705);
nand NAND2_138(G1755,G990,G1718);
not NOT_318(G1756,G1616);
not NOT_319(G1761,G1616);
nand NAND2_139(G1766,G1546,G1720);
nand NAND2_140(G1767,G1543,G1721);
nand NAND2_141(G1768,G1552,G1722);
nand NAND2_142(G1769,G1549,G1723);
nand NAND2_143(G1770,G1563,G1724);
nand NAND2_144(G1771,G1560,G1725);
nand NAND2_145(G1772,G1569,G1726);
nand NAND2_146(G1773,G1566,G1727);
nand NAND2_147(G1774,G1593,G1732);
nand NAND2_148(G1775,G1590,G1733);
or OR2_23(G1776,G1734,G1610);
or OR2_24(G1777,G1735,G1607);
and AND2_80(G1778,G1152,G1670);
and AND2_81(G1779,G1159,G1670);
and AND2_82(G1780,G1166,G1670);
and AND2_83(G1781,G1171,G1670);
not NOT_320(G1782,G1646);
nand NAND2_149(G1785,G1736,G1651);
nand NAND2_150(G1789,G1652,G1737);
not NOT_321(G1792,G1657);
nand NAND2_151(G1795,G1738,G1662);
and AND2_84(G1798,G1152,G1676);
and AND2_85(G1799,G1159,G1676);
and AND2_86(G1800,G1166,G1676);
and AND2_87(G1801,G1171,G1676);
and AND2_88(G1802,G1749,G10);
not NOT_322(G1805,G1636);
nand NAND2_152(G1811,G1750,G1689);
and AND2_89(G1814,G1751,G1752);
and AND2_90(G1815,G1753,G1754);
not NOT_323(G1816,G1684);
not NOT_324(G1822,G1712);
not NOT_325(G1823,G1715);
and AND3_90(G1824,G1524,G1520,G1712);
and AND3_91(G1825,G1709,G1706,G1715);
nand NAND2_153(G1826,G1755,G1719);
not NOT_326(G1829,G1636);
not NOT_327(G1835,G1636);
not NOT_328(G1840,G1684);
not NOT_329(G1846,G1684);
nand NAND2_154(G1851,G1768,G1769);
nand NAND2_155(G1854,G1766,G1767);
not NOT_330(G1857,G1728);
nand NAND2_156(G1858,G1728,G1731);
nand NAND2_157(G1859,G1772,G1773);
nand NAND2_158(G1862,G1770,G1771);
nand NAND2_159(G1865,G1774,G1775);
and AND2_91(G1868,G1640,G1739);
and AND2_92(G1869,G1641,G1739);
and AND2_93(G1870,G1642,G1739);
and AND2_94(G1871,G1643,G1739);
or OR2_25(G1872,G1778,G1644);
or OR2_26(G1873,G1779,G1645);
and AND2_95(G1874,G1780,G598);
and AND2_96(G1875,G1781,G598);
or OR2_27(G1876,G1798,G1664);
or OR2_28(G1877,G1799,G1665);
and AND2_97(G1878,G1800,G631);
and AND2_98(G1879,G1801,G631);
and AND2_99(G1880,G1666,G1744);
and AND2_100(G1881,G1667,G1744);
and AND2_101(G1882,G1668,G1744);
and AND2_102(G1883,G1669,G1744);
and AND3_92(G1884,G1814,G1815,G832);
and AND3_93(G1887,G1706,G1524,G1822);
and AND3_94(G1888,G1520,G1709,G1823);
nand NAND2_160(G1889,G1572,G1857);
not NOT_331(G1890,G1868);
not NOT_332(G1893,G1869);
not NOT_333(G1896,G1870);
not NOT_334(G1899,G1871);
and AND2_103(G1902,G1872,G598);
and AND2_104(G1903,G1873,G598);
not NOT_335(G1904,G1874);
not NOT_336(G1907,G1875);
not NOT_337(G1910,G1785);
not NOT_338(G1913,G1789);
not NOT_339(G1916,G1789);
not NOT_340(G1919,G1795);
not NOT_341(G1922,G1795);
and AND2_105(G1925,G366,G1805);
and AND2_106(G1926,G1876,G631);
and AND2_107(G1927,G1877,G631);
not NOT_342(G1928,G1878);
not NOT_343(G1931,G1879);
not NOT_344(G1934,G1880);
not NOT_345(G1937,G1881);
not NOT_346(G1940,G1882);
not NOT_347(G1943,G1883);
not NOT_348(G1946,G1802);
and AND2_108(G1947,G366,G1816);
not NOT_349(G1948,G1805);
and AND2_109(G1953,G370,G1805);
and AND2_110(G1954,G447,G1805);
and AND2_111(G1955,G451,G1805);
not NOT_350(G1956,G1816);
and AND2_112(G1961,G370,G1816);
and AND2_113(G1962,G447,G1816);
and AND2_114(G1963,G451,G1816);
nor NOR2_6(G1964,G1887,G1824);
nor NOR2_7(G1965,G1888,G1825);
not NOT_351(G1966,G1865);
not NOT_352(G1967,G1829);
and AND2_115(G1970,G455,G1829);
and AND2_116(G1971,G459,G1829);
and AND2_117(G1972,G463,G1829);
and AND2_118(G1973,G467,G1829);
and AND2_119(G1974,G471,G1835);
and AND2_120(G1975,G475,G1835);
and AND2_121(G1976,G479,G1835);
and AND2_122(G1977,G497,G1835);
not NOT_353(G1978,G1840);
and AND2_123(G1981,G455,G1840);
and AND2_124(G1982,G459,G1840);
and AND2_125(G1983,G463,G1840);
and AND2_126(G1984,G467,G1840);
and AND2_127(G1985,G471,G1846);
and AND2_128(G1986,G475,G1846);
and AND2_129(G1987,G479,G1846);
and AND2_130(G1988,G497,G1846);
not NOT_354(G1989,G1851);
not NOT_355(G1990,G1854);
not NOT_356(G1991,G1859);
not NOT_357(G1992,G1862);
nand NAND2_161(G1993,G1858,G1889);
not NOT_358(G1996,G1902);
not NOT_359(G1999,G1903);
not NOT_360(G2002,G1926);
not NOT_361(G2005,G1927);
and AND2_131(G2008,G1972,G751);
and AND2_132(G2011,G1973,G751);
and AND2_133(G2014,G1974,G1756);
and AND2_134(G2017,G1975,G1756);
and AND2_135(G2020,G1976,G1756);
and AND2_136(G2023,G1977,G1756);
and AND2_137(G2026,G1983,G756);
and AND2_138(G2029,G1984,G756);
and AND2_139(G2032,G1985,G1761);
and AND2_140(G2035,G1986,G1761);
and AND2_141(G2038,G1987,G1761);
and AND2_142(G2041,G1988,G1761);
nand NAND2_162(G2044,G1854,G1989);
nand NAND2_163(G2045,G1851,G1990);
nand NAND2_164(G2046,G1862,G1991);
nand NAND2_165(G2047,G1859,G1992);
nand NAND2_166(G2048,G1965,G1964);
not NOT_362(G2051,G1913);
not NOT_363(G2052,G1916);
not NOT_364(G2053,G1919);
not NOT_365(G2054,G1922);
and AND3_95(G2055,G1785,G1646,G1913);
and AND3_96(G2056,G1910,G1782,G1916);
and AND3_97(G2057,G1657,G1479,G1919);
and AND3_98(G2058,G1792,G1654,G1922);
nand NAND2_167(G2059,G1993,G1486);
not NOT_366(G2060,G1993);
and AND2_143(G2061,G479,G1948);
and AND2_144(G2062,G479,G1956);
and AND2_145(G2063,G497,G1948);
and AND2_146(G2064,G503,G1948);
and AND2_147(G2065,G507,G1948);
and AND2_148(G2066,G497,G1956);
and AND2_149(G2067,G503,G1956);
and AND2_150(G2068,G507,G1956);
and AND2_151(G2069,G511,G1967);
and AND2_152(G2070,G515,G1967);
and AND2_153(G2071,G511,G1978);
and AND2_154(G2072,G515,G1978);
nand NAND2_168(G2073,G2044,G2045);
nand NAND2_169(G2076,G2046,G2047);
not NOT_367(G2079,G1899);
not NOT_368(G2082,G1896);
not NOT_369(G2085,G1893);
not NOT_370(G2088,G1890);
not NOT_371(G2091,G1907);
not NOT_372(G2094,G1904);
not NOT_373(G2097,G1943);
not NOT_374(G2100,G1940);
not NOT_375(G2103,G1937);
not NOT_376(G2106,G1934);
not NOT_377(G2109,G1931);
not NOT_378(G2112,G1928);
and AND3_99(G2115,G1782,G1785,G2051);
and AND3_100(G2116,G1646,G1910,G2052);
and AND3_101(G2117,G1654,G1657,G2053);
and AND3_102(G2118,G1479,G1792,G2054);
nand NAND2_170(G2119,G1393,G2060);
or OR2_29(G2120,G2061,G1925);
nand NAND2_171(G2121,G2048,G1966);
and AND2_155(G2122,G2023,G1899);
and AND2_156(G2123,G2020,G1896);
and AND2_157(G2124,G2017,G1893);
and AND2_158(G2125,G1890,G2014);
and AND2_159(G2126,G2011,G1907);
and AND2_160(G2127,G2008,G1904);
or OR2_30(G2128,G2062,G1947);
and AND2_161(G2129,G2041,G1943);
and AND2_162(G2130,G2038,G1940);
and AND2_163(G2131,G2035,G1937);
and AND2_164(G2132,G1934,G2032);
and AND2_165(G2133,G2029,G1931);
and AND2_166(G2134,G2026,G1928);
or OR2_31(G2135,G2063,G1953);
or OR2_32(G2138,G2064,G1954);
or OR2_33(G2141,G2065,G1955);
or OR2_34(G2144,G2066,G1961);
or OR2_35(G2147,G2067,G1962);
or OR2_36(G2150,G2068,G1963);
not NOT_379(G2153,G2048);
or OR2_37(G2154,G2069,G1970);
or OR2_38(G2155,G2070,G1971);
or OR2_39(G2156,G2071,G1981);
or OR2_40(G2157,G2072,G1982);
not NOT_380(G2158,G2023);
not NOT_381(G2161,G2020);
not NOT_382(G2164,G2017);
not NOT_383(G2167,G2014);
not NOT_384(G2170,G2011);
not NOT_385(G2173,G2008);
not NOT_386(G2176,G1999);
not NOT_387(G2179,G1996);
not NOT_388(G2182,G2041);
not NOT_389(G2185,G2038);
not NOT_390(G2188,G2035);
not NOT_391(G2191,G2032);
not NOT_392(G2194,G2029);
not NOT_393(G2197,G2026);
not NOT_394(G2200,G2005);
not NOT_395(G2203,G2002);
nand NAND2_172(G2206,G2059,G2119);
nor NOR2_8(G2207,G2115,G2055);
nor NOR2_9(G2208,G2116,G2056);
nor NOR2_10(G2209,G2117,G2057);
nor NOR2_11(G2210,G2118,G2058);
not NOT_396(G2211,G2073);
not NOT_397(G2212,G2076);
and AND2_167(G2213,G2120,G1132);
nand NAND2_173(G2214,G1865,G2153);
not NOT_398(G2215,G2079);
not NOT_399(G2216,G2082);
not NOT_400(G2217,G2085);
not NOT_401(G2218,G2088);
not NOT_402(G2219,G2091);
not NOT_403(G2220,G2094);
and AND2_168(G2221,G2128,G1132);
not NOT_404(G2222,G2097);
not NOT_405(G2223,G2100);
not NOT_406(G2224,G2103);
not NOT_407(G2225,G2106);
not NOT_408(G2226,G2109);
not NOT_409(G2227,G2112);
and AND2_169(G2228,G2154,G751);
and AND2_170(G2231,G2155,G751);
and AND2_171(G2234,G2156,G756);
and AND2_172(G2237,G2157,G756);
and AND2_173(G2240,G2206,G325);
and AND2_174(G2241,G2138,G1329);
and AND2_175(G2242,G2135,G1137);
nand NAND2_174(G2243,G2214,G2121);
not NOT_410(G2244,G2158);
nand NAND2_175(G2245,G2158,G2215);
not NOT_411(G2246,G2161);
nand NAND2_176(G2247,G2161,G2216);
not NOT_412(G2248,G2164);
nand NAND2_177(G2249,G2164,G2217);
not NOT_413(G2250,G2167);
nand NAND2_178(G2251,G2167,G2218);
not NOT_414(G2252,G2170);
nand NAND2_179(G2253,G2170,G2219);
not NOT_415(G2254,G2173);
nand NAND2_180(G2255,G2173,G2220);
not NOT_416(G2256,G2176);
not NOT_417(G2257,G2179);
and AND2_176(G2258,G2141,G1336);
and AND2_177(G2259,G2147,G1329);
and AND2_178(G2260,G2144,G1137);
not NOT_418(G2261,G2182);
nand NAND2_181(G2262,G2182,G2222);
not NOT_419(G2263,G2185);
nand NAND2_182(G2264,G2185,G2223);
not NOT_420(G2265,G2188);
nand NAND2_183(G2266,G2188,G2224);
not NOT_421(G2267,G2191);
nand NAND2_184(G2268,G2191,G2225);
not NOT_422(G2269,G2194);
nand NAND2_185(G2270,G2194,G2226);
not NOT_423(G2271,G2197);
nand NAND2_186(G2272,G2197,G2227);
not NOT_424(G2273,G2200);
not NOT_425(G2274,G2203);
and AND2_179(G2275,G2150,G1336);
nand NAND2_187(G2276,G2208,G2207);
nand NAND2_188(G2279,G2210,G2209);
not NOT_426(G2282,G2138);
not NOT_427(G2285,G2135);
not NOT_428(G2288,G2141);
not NOT_429(G2291,G2147);
not NOT_430(G2294,G2144);
not NOT_431(G2297,G2150);
not NOT_432(G2300,G2243);
nand NAND2_189(G2301,G2079,G2244);
nand NAND2_190(G2302,G2082,G2246);
nand NAND2_191(G2303,G2085,G2248);
nand NAND2_192(G2304,G2088,G2250);
nand NAND2_193(G2305,G2091,G2252);
nand NAND2_194(G2306,G2094,G2254);
and AND2_180(G2307,G2231,G1999);
and AND2_181(G2308,G2228,G1996);
nand NAND2_195(G2309,G2097,G2261);
nand NAND2_196(G2310,G2100,G2263);
nand NAND2_197(G2311,G2103,G2265);
nand NAND2_198(G2312,G2106,G2267);
nand NAND2_199(G2313,G2109,G2269);
nand NAND2_200(G2314,G2112,G2271);
and AND2_182(G2315,G2237,G2005);
and AND2_183(G2316,G2234,G2002);
not NOT_433(G2317,G2231);
not NOT_434(G2320,G2228);
not NOT_435(G2323,G2237);
not NOT_436(G2326,G2234);
not NOT_437(G2329,G2276);
nand NAND2_201(G2330,G2276,G2211);
not NOT_438(G2331,G2279);
nand NAND2_202(G2332,G2279,G2212);
not NOT_439(G2333,G2282);
nand NAND2_203(G2334,G2282,G1663);
nand NAND2_204(G2335,G2285,G1487);
not NOT_440(G2336,G2285);
and AND2_184(G2337,G2300,G581);
nand NAND2_205(G2340,G2301,G2245);
nand NAND2_206(G2345,G2302,G2247);
nand NAND2_207(G2349,G2303,G2249);
nand NAND2_208(G2352,G2304,G2251);
nand NAND2_209(G2353,G2305,G2253);
nand NAND2_210(G2359,G2306,G2255);
not NOT_441(G2364,G2288);
nand NAND2_211(G2365,G2288,G1675);
not NOT_442(G2366,G2291);
nand NAND2_212(G2367,G2291,G1682);
nand NAND2_213(G2368,G2294,G1508);
not NOT_443(G2369,G2294);
nand NAND2_214(G2370,G2309,G2262);
nand NAND2_215(G2375,G2310,G2264);
nand NAND2_216(G2379,G2311,G2266);
nand NAND2_217(G2382,G2312,G2268);
nand NAND2_218(G2383,G2313,G2270);
nand NAND2_219(G2389,G2314,G2272);
not NOT_444(G2394,G2297);
nand NAND2_220(G2395,G2297,G1683);
nand NAND2_221(G2396,G2073,G2329);
nand NAND2_222(G2397,G2076,G2331);
nand NAND2_223(G2398,G1575,G2333);
nand NAND2_224(G2399,G1396,G2336);
not NOT_445(G2400,G2317);
nand NAND2_225(G2401,G2317,G2256);
not NOT_446(G2402,G2320);
nand NAND2_226(G2403,G2320,G2257);
nand NAND2_227(G2404,G1578,G2364);
nand NAND2_228(G2405,G1581,G2366);
nand NAND2_229(G2406,G1399,G2369);
not NOT_447(G2407,G2323);
nand NAND2_230(G2408,G2323,G2273);
not NOT_448(G2409,G2326);
nand NAND2_231(G2410,G2326,G2274);
nand NAND2_232(G2411,G1584,G2394);
nand NAND2_233(G2412,G2396,G2330);
nand NAND2_234(G2413,G2397,G2332);
nand NAND2_235(G2414,G2398,G2334);
nand NAND2_236(G2417,G2399,G2335);
not NOT_449(G2418,G2337);
nand NAND2_237(G2419,G2176,G2400);
nand NAND2_238(G2420,G2179,G2402);
nand NAND2_239(G2421,G2404,G2365);
and AND4_5(G2422,G2345,G2352,G2349,G2340);
and AND2_185(G2423,G2340,G2123);
and AND3_103(G2424,G2345,G2340,G2124);
and AND4_6(G2425,G2349,G2340,G2125,G2345);
and AND2_186(G2426,G2353,G2127);
and AND3_104(G2427,G2359,G2353,G2307);
nand NAND2_240(G2428,G2405,G2367);
nand NAND2_241(G2431,G2406,G2368);
nand NAND2_242(G2432,G2200,G2407);
nand NAND2_243(G2433,G2203,G2409);
nand NAND2_244(G2434,G2411,G2395);
and AND4_7(G2435,G2375,G2382,G2379,G2370);
and AND2_187(G2436,G2370,G2130);
and AND3_105(G2437,G2375,G2370,G2131);
and AND4_8(G2438,G2379,G2370,G2132,G2375);
and AND2_188(G2439,G2383,G2134);
and AND3_106(G2440,G2389,G2383,G2315);
not NOT_450(G2441,G2412);
and AND2_189(G2442,G2413,G123);
nand NAND2_245(G2443,G2419,G2401);
nand NAND2_246(G2447,G2420,G2403);
not NOT_451(G2450,G2422);
or OR4_20(G2451,G2122,G2423,G2424,G2425);
nand NAND2_247(G2454,G2432,G2408);
nand NAND2_248(G2458,G2433,G2410);
not NOT_452(G2461,G2435);
or OR4_21(G2462,G2129,G2436,G2437,G2438);
and AND2_190(G2465,G2414,G2242);
and AND3_107(G2466,G2417,G2414,G2213);
or OR2_41(G2467,G1326,G2442);
and AND2_191(G2470,G2441,G581);
and AND2_192(G2473,G2428,G2260);
and AND3_108(G2474,G2431,G2428,G2221);
or OR3_0(G2475,G2241,G2465,G2466);
not NOT_453(G2476,G2451);
and AND5_3(G2477,G2359,G2421,G2443,G2353,G2447);
and AND4_9(G2478,G2443,G2353,G2308,G2359);
and AND5_4(G2479,G2447,G2443,G2353,G2258,G2359);
or OR3_1(G2480,G2259,G2473,G2474);
not NOT_454(G2481,G2462);
and AND5_5(G2482,G2389,G2434,G2454,G2383,G2458);
and AND4_10(G2483,G2454,G2383,G2316,G2389);
and AND5_6(G2484,G2458,G2454,G2383,G2275,G2389);
or OR5_0(G2485,G2126,G2426,G2427,G2478,G2479);
and AND2_193(G2486,G2477,G2475);
nand NAND2_249(G2487,G2476,G2450);
not NOT_455(G2488,G2470);
or OR5_1(G2489,G2133,G2439,G2440,G2483,G2484);
and AND2_194(G2490,G2482,G2480);
nand NAND2_250(G2491,G2481,G2461);
or OR2_42(G2492,G2485,G2486);
and AND3_109(G2495,G2418,G2488,G1826);
or OR2_43(G2496,G2489,G2490);
not NOT_456(G2499,G2492);
and AND2_195(G2500,G2487,G2492);
not NOT_457(G2501,G2496);
and AND2_196(G2502,G2491,G2496);
and AND2_197(G2503,G2451,G2499);
and AND2_198(G2504,G2462,G2501);
or OR2_44(G2505,G2503,G2500);
or OR2_45(G2508,G2504,G2502);
nand NAND2_251(G2512,G2508,G2505);
and AND2_199(G2515,G2508,G2512);
and AND2_200(G2516,G2512,G2505);
or OR2_46(G2517,G2515,G2516);
not NOT_458(G2520,G2517);
and AND2_201(G2523,G2517,G2520);
or OR2_47(G2524,G2523,G2520);
and AND3_110(G2527,G1811,G1946,G2524);
and AND3_111(G2528,G2495,G2527,G993);
not NOT_459(G2531,G115);
not NOT_460(G2532,G115);
not NOT_461(G2533,G115);
not NOT_462(G2534,G124);
not NOT_463(G2535,G124);
not NOT_464(G2536,G137);
not NOT_465(G2537,G137);
not NOT_466(G2538,G137);
not NOT_467(G2539,G32);
not NOT_468(G2540,G106);
not NOT_469(G2541,G64);
not NOT_470(G2542,G76);
not NOT_471(G2543,G53);
not NOT_472(G2544,G96);
not NOT_473(G2545,G43);
not NOT_474(G2546,G86);
not NOT_475(G2547,G285);
not NOT_476(G2548,G287);
not NOT_477(G2549,G292);
and AND2_202(G2550,G74,G292);
not NOT_478(G2551,G443);
nand NAND2_252(G2552,G119,G443);
not NOT_479(G2553,G592);
not NOT_480(G2554,G595);
not NOT_481(G2555,G595);
not NOT_482(G2556,G993);
not NOT_483(G2557,G1044);
not NOT_484(G2558,G1049);
not NOT_485(G2559,G1039);
not NOT_486(G2560,G1026);
not NOT_487(G2561,G1021);
not NOT_488(G2562,G1017);
or OR2_48(G2563,G325,G1117);
not NOT_489(G2564,G1118);
not NOT_490(G2565,G1119);
not NOT_491(G2566,G1144);
not NOT_492(G2567,G1148);
not NOT_493(G2568,G1152);
not NOT_494(G2569,G1159);
not NOT_495(G2570,G1166);
not NOT_496(G2571,G1171);
not NOT_497(G2572,G1176);
not NOT_498(G2573,G1412);
not NOT_499(G2574,G1412);
not NOT_500(G2575,G1415);
not NOT_501(G2576,G1415);
or OR2_49(G2577,G1471,G1116);
not NOT_502(G2578,G1603);
not NOT_503(G2579,G1603);
nand NAND2_253(G2580,G1776,G1777);
not NOT_504(G2581,G1802);
not NOT_505(G2582,G1826);
not NOT_506(G2583,G1811);
not NOT_507(G2584,G1884);
not NOT_508(G2585,G1884);
or OR2_50(G2586,G2240,G1115);
not NOT_509(G2587,G2337);
not NOT_510(G2588,G2467);
not NOT_511(G2589,G2467);
not NOT_512(G2590,G2470);
not NOT_513(G2591,G2508);
not NOT_514(G2592,G2524);
not NOT_515(G2593,G2528);
not NOT_516(G2594,G2528);

endmodule