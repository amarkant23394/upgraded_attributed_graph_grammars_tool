module test_I8913(I7139,I6992,I1477,I1470,I8913);
input I7139,I6992,I1477,I1470;
output I8913;
wire I7190,I8896,I6893,I7156,I6872,I5067,I6907,I7269,I7286,I6878;
DFFARX1 I_0(I7156,I1470,I6907,,,I7190,);
nor I_1(I8896,I6893,I6872);
nand I_2(I6893,I7156,I7286);
nand I_3(I8913,I8896,I6878);
DFFARX1 I_4(I7139,I1470,I6907,,,I7156,);
DFFARX1 I_5(I7269,I1470,I6907,,,I6872,);
DFFARX1 I_6(I1470,,,I5067,);
not I_7(I6907,I1477);
DFFARX1 I_8(I5067,I1470,I6907,,,I7269,);
nor I_9(I7286,I7269,I6992);
not I_10(I6878,I7190);
endmodule


