module test_I6303(I2727,I1477,I1470,I4068,I6303);
input I2727,I1477,I1470,I4068;
output I6303;
wire I6781,I6329,I4113,I4308,I4130,I3957,I3983;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
not I_1(I6329,I1477);
DFFARX1 I_2(I1470,I3983,,,I4113,);
DFFARX1 I_3(I2727,I1470,I3983,,,I4308,);
nor I_4(I4130,I4113,I4068);
nand I_5(I3957,I4308,I4130);
DFFARX1 I_6(I6781,I1470,I6329,,,I6303,);
not I_7(I3983,I1477);
endmodule


