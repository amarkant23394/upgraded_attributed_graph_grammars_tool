module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_0,blif_reset_net_5_r_0,N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_0,blif_reset_net_5_r_0;
output N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,n_102_5_r_0,n_452_7_r_0,n_431_5_r_0,n6_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_5_r_0,n6_0,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_37(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_38(n_429_or_0_5_r_0,n38_0,N1507_6_r_3);
DFFARX1 I_39(n_431_5_r_0,blif_clk_net_5_r_0,n6_0,G78_5_r_0,);
nand I_40(n_576_5_r_0,n26_0,N1507_6_r_3);
not I_41(n_102_5_r_0,n27_0);
nand I_42(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_43(n4_7_r_0,blif_clk_net_5_r_0,n6_0,G42_7_r_0,);
nor I_44(n_572_7_r_0,n31_0,N1507_6_r_3);
or I_45(n_573_7_r_0,n29_0,n30_0);
nor I_46(n_549_7_r_0,n29_0,n33_0);
nand I_47(n_569_7_r_0,n28_0,n32_0);
nor I_48(n_452_7_r_0,n30_0,n31_0);
nand I_49(n_431_5_r_0,n_102_5_r_0,n35_0);
not I_50(n6_0,blif_reset_net_5_r_0);
nor I_51(n4_7_r_0,n31_0,n37_0);
nor I_52(n26_0,n27_0,n28_0);
nor I_53(n27_0,n28_0,n44_0);
nand I_54(n28_0,n_573_7_r_3,N1372_1_r_3);
not I_55(n29_0,n32_0);
nor I_56(n30_0,n39_0,N1508_1_r_3);
not I_57(n31_0,n38_0);
nand I_58(n32_0,n41_0,n42_0);
nor I_59(n33_0,n_102_5_r_0,N1507_6_r_3);
nor I_60(n34_0,n27_0,N1507_6_r_3);
nand I_61(n35_0,n29_0,n36_0);
nor I_62(n36_0,n37_0,n38_0);
not I_63(n37_0,n28_0);
nand I_64(n38_0,n40_0,n_569_7_r_3);
nor I_65(n39_0,n_452_7_r_3,N1508_6_r_3);
or I_66(n40_0,n_452_7_r_3,N1508_6_r_3);
nor I_67(n41_0,N1508_6_r_3,N1508_1_r_3);
or I_68(n42_0,n43_0,N1372_1_r_3);
nor I_69(n43_0,N6134_9_r_3,G42_7_r_3);
nor I_70(n44_0,n45_0,G42_7_r_3);
and I_71(n45_0,N1507_6_r_3,n_549_7_r_3);
endmodule


