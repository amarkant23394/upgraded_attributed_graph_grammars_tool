module test_I1767(I1439,I1367,I1477,I1279,I1470,I1699,I1767);
input I1439,I1367,I1477,I1279,I1470,I1699;
output I1767;
wire I1518,I1750,I1733,I1716;
not I_0(I1518,I1477);
or I_1(I1750,I1733,I1279);
and I_2(I1733,I1716,I1439);
nor I_3(I1716,I1699,I1367);
DFFARX1 I_4(I1750,I1470,I1518,,,I1767,);
endmodule


