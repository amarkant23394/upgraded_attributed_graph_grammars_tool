module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_7_r_16,n8_16,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_7_r_16,n8_16,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_16,n35_16,n39_16);
nor I_36(N1508_0_r_16,n39_16,n46_16);
not I_37(N1372_1_r_16,n45_16);
nor I_38(N1508_1_r_16,n53_16,n45_16);
nor I_39(N6147_2_r_16,n37_16,n38_16);
nor I_40(N1507_6_r_16,n44_16,n49_16);
nor I_41(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_42(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_43(n_572_7_r_16,n32_16,n33_16);
nand I_44(n_573_7_r_16,n30_16,n31_16);
nand I_45(n_549_7_r_16,n47_16,G78_5_r_0);
nand I_46(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_47(n_452_7_r_16,n34_16,n35_16);
and I_48(N3_8_l_16,n41_16,G78_5_r_0);
not I_49(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_50(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_51(n29_16,n53_16);
nor I_52(n4_7_r_16,n35_16,n36_16);
nand I_53(n30_16,n_429_or_0_5_r_0,n_547_5_r_0);
not I_54(n31_16,n34_16);
nor I_55(n32_16,n30_16,n_549_7_r_0);
not I_56(n33_16,n_549_7_r_16);
nor I_57(n34_16,n48_16,n_569_7_r_0);
and I_58(n35_16,n50_16,N1371_0_r_0);
not I_59(n36_16,n30_16);
nor I_60(n37_16,n31_16,n40_16);
nand I_61(n38_16,n29_16,n39_16);
not I_62(n39_16,n32_16);
nor I_63(n40_16,G42_7_r_0,n_572_7_r_0);
nand I_64(n41_16,n_576_5_r_0,n_572_7_r_0);
nand I_65(n42_16,n35_16,n43_16);
not I_66(n43_16,n44_16);
nor I_67(n44_16,n32_16,n49_16);
nand I_68(n45_16,n36_16,n40_16);
nor I_69(n46_16,n33_16,n34_16);
nand I_70(n47_16,N1371_0_r_0,n_429_or_0_5_r_0);
or I_71(n48_16,N1508_0_r_0,n_573_7_r_0);
and I_72(n49_16,n35_16,n36_16);
and I_73(n50_16,n51_16,N1508_0_r_0);
nand I_74(n51_16,n47_16,n52_16);
not I_75(n52_16,G78_5_r_0);
endmodule


