module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_17,n6_17,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_17,n6_17,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_17,n6_17,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_17,n6_17,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_17,n6_17,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_17,n6_17,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_17,n6_17,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_17,n6_17,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_17,n6_17,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_34(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_35(n_573_1_r_17,n20_17,n21_17);
nand I_36(n_549_1_r_17,n23_17,n24_17);
nand I_37(n_569_1_r_17,n21_17,n22_17);
not I_38(n_452_1_r_17,n23_17);
DFFARX1 I_39(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_40(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_41(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_42(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_43(n_431_0_l_17,n26_17,G199_4_r_9);
not I_44(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_45(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_46(n20_17,n20_internal_17);
DFFARX1 I_47(n_549_1_r_9,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_48(n_572_1_r_9,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_49(n19_17,n19_internal_17);
nor I_50(n4_1_r_17,n5_17,n25_17);
not I_51(n2_17,n29_17);
DFFARX1 I_52(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_53(n17_17,n17_internal_17);
nor I_54(N1_4_r_17,n29_17,n31_17);
not I_55(n5_17,G214_4_r_9);
and I_56(n21_17,n32_17,G42_1_r_9);
not I_57(n22_17,n25_17);
nand I_58(n23_17,n20_17,n22_17);
nand I_59(n24_17,n19_17,n22_17);
nand I_60(n25_17,n30_17,n_572_1_r_9);
and I_61(n26_17,n27_17,n_569_1_r_9);
nor I_62(n27_17,n28_17,n_573_1_r_9);
not I_63(n28_17,n_42_2_r_9);
nor I_64(n29_17,n28_17,G199_2_r_9);
and I_65(n30_17,n5_17,G199_2_r_9);
nor I_66(n31_17,n21_17,G214_4_r_9);
nor I_67(n32_17,G214_4_r_9,G42_1_r_9);
endmodule


