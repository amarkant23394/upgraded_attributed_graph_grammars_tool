module test_I6315(I1477,I4068,I3963,I2727,I1470,I6315);
input I1477,I4068,I3963,I2727,I1470;
output I6315;
wire I6781,I6442,I6380,I4130,I3983,I6476,I3954,I6346,I6329,I6363,I6459,I3975,I4308,I4113,I3957;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
nor I_1(I6442,I3975,I3954);
DFFARX1 I_2(I6363,I1470,I6329,,,I6380,);
nor I_3(I4130,I4113,I4068);
nand I_4(I6315,I6781,I6476);
not I_5(I3983,I1477);
nor I_6(I6476,I6380,I6459);
not I_7(I3954,I4068);
nand I_8(I6346,I3954);
not I_9(I6329,I1477);
and I_10(I6363,I6346,I3963);
not I_11(I6459,I6442);
nor I_12(I3975,I4308);
DFFARX1 I_13(I2727,I1470,I3983,,,I4308,);
DFFARX1 I_14(I1470,I3983,,,I4113,);
nand I_15(I3957,I4308,I4130);
endmodule


