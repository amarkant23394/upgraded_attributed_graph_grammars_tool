module test_final(IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_102_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13,n4_7_l_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N1371_0_r_13,n59_13,n61_13);
nor I_1(N1508_0_r_13,n59_13,n60_13);
not I_2(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_3(n_431_5_r_13,blif_clk_net_5_r_15,n9_15,G78_5_r_13,);
nand I_4(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_5(n_102_5_r_13,IN_9_7_l_13,IN_10_7_l_13);
nand I_6(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_7(n1_13,blif_clk_net_5_r_15,n9_15,G42_7_r_13,);
nor I_8(n_572_7_r_13,n40_13,n41_13);
nand I_9(n_573_7_r_13,n37_13,n38_13);
nor I_10(n_549_7_r_13,n46_13,n47_13);
nand I_11(n_569_7_r_13,n37_13,n43_13);
nand I_12(n_452_7_r_13,n52_13,n53_13);
nor I_13(n4_7_l_13,G18_7_l_13,IN_1_7_l_13);
DFFARX1 I_14(n4_7_l_13,blif_clk_net_5_r_15,n9_15,n62_13,);
not I_15(n33_13,n62_13);
nand I_16(n_431_5_r_13,n54_13,n55_13);
not I_17(n1_13,n52_13);
nor I_18(n34_13,n35_13,n36_13);
nor I_19(n35_13,G15_7_l_13,n42_13);
nand I_20(n36_13,n50_13,n58_13);
nand I_21(n37_13,n44_13,n45_13);
or I_22(n38_13,IN_3_1_l_13,n39_13);
nand I_23(n39_13,IN_1_1_l_13,IN_2_1_l_13);
not I_24(n40_13,n36_13);
nor I_25(n41_13,IN_10_7_l_13,n35_13);
not I_26(n42_13,IN_4_7_l_13);
or I_27(n43_13,G18_7_l_13,IN_5_7_l_13);
not I_28(n44_13,G15_7_l_13);
not I_29(n45_13,IN_7_7_l_13);
nor I_30(n46_13,n39_13,n40_13);
nor I_31(n47_13,G18_7_l_13,IN_5_7_l_13);
nor I_32(n48_13,n50_13,n51_13);
nor I_33(n49_13,G15_7_l_13,IN_7_7_l_13);
not I_34(n50_13,n59_13);
not I_35(n51_13,n_102_5_r_13);
nand I_36(n52_13,n33_13,n39_13);
nand I_37(n53_13,IN_3_1_l_13,n33_13);
nor I_38(n54_13,IN_5_7_l_13,IN_9_7_l_13);
nand I_39(n55_13,n62_13,n56_13);
nor I_40(n56_13,n39_13,n57_13);
not I_41(n57_13,G18_7_l_13);
or I_42(n58_13,IN_3_10_l_13,IN_4_10_l_13);
nand I_43(n59_13,IN_1_10_l_13,IN_2_10_l_13);
nor I_44(n60_13,IN_5_7_l_13,n51_13);
nor I_45(n61_13,IN_3_1_l_13,n39_13);
and I_46(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_47(N1508_0_r_15,n55_15,N1508_0_r_13);
nor I_48(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_49(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_50(N1372_4_r_15,n39_15);
nor I_51(N1508_4_r_15,n39_15,n43_15);
nand I_52(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_53(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_54(n_576_5_r_15,n31_15,n32_15);
not I_55(n_102_5_r_15,n33_15);
nand I_56(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_57(N1507_6_r_15,n42_15,n46_15);
nand I_58(N1508_6_r_15,n39_15,n40_15);
nand I_59(n_431_5_r_15,n36_15,n37_15);
not I_60(n9_15,blif_reset_net_5_r_15);
nor I_61(n31_15,n33_15,n34_15);
nor I_62(n32_15,n44_15,N1508_0_r_13);
nor I_63(n33_15,n54_15,n55_15);
nand I_64(n34_15,n49_15,n_569_7_r_13);
nand I_65(n35_15,n_547_5_r_13,n_573_7_r_13);
not I_66(n36_15,n32_15);
nand I_67(n37_15,n34_15,n38_15);
not I_68(n38_15,n46_15);
nand I_69(n39_15,n38_15,n41_15);
nand I_70(n40_15,n41_15,n42_15);
and I_71(n41_15,n51_15,n_576_5_r_13);
and I_72(n42_15,n47_15,n_547_5_r_13);
and I_73(n43_15,n34_15,n36_15);
or I_74(n44_15,n_429_or_0_5_r_13,n_452_7_r_13);
not I_75(n45_15,N1372_1_r_15);
nand I_76(n46_15,n53_15,n_547_5_r_13);
nor I_77(n47_15,n34_15,n48_15);
not I_78(n48_15,n_573_7_r_13);
and I_79(n49_15,n50_15,N1371_0_r_13);
nand I_80(n50_15,n51_15,n52_15);
nand I_81(n51_15,N1371_0_r_13,n_429_or_0_5_r_13);
not I_82(n52_15,n_576_5_r_13);
nor I_83(n53_15,n48_15,n_572_7_r_13);
nor I_84(n54_15,G42_7_r_13,n_549_7_r_13);
not I_85(n55_15,G78_5_r_13);
endmodule


