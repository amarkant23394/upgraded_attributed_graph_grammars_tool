module test_final(IN_1_1_l_3,IN_2_1_l_3,IN_3_1_l_3,IN_1_8_l_3,IN_2_8_l_3,IN_3_8_l_3,IN_6_8_l_3,IN_1_10_l_3,IN_2_10_l_3,IN_3_10_l_3,IN_4_10_l_3,blif_clk_net_5_r_4,blif_reset_net_5_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4);
input IN_1_1_l_3,IN_2_1_l_3,IN_3_1_l_3,IN_1_8_l_3,IN_2_8_l_3,IN_3_8_l_3,IN_6_8_l_3,IN_1_10_l_3,IN_2_10_l_3,IN_3_10_l_3,IN_4_10_l_3,blif_clk_net_5_r_4,blif_reset_net_5_r_4;
output N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4;
wire N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1372_10_r_3,N1508_10_r_3,N3_8_l_3,n39_3,n_431_5_r_3,n22_3,n23_3,n24_3,n25_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,N1371_0_r_4,n_102_5_r_4,n_431_5_r_4,n4_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4;
nor I_0(N1371_0_r_3,n39_3,n37_3);
nor I_1(N1508_0_r_3,n25_3,n37_3);
nor I_2(N6147_3_r_3,N1372_10_r_3,n33_3);
nand I_3(n_429_or_0_5_r_3,N1372_10_r_3,n30_3);
DFFARX1 I_4(n_431_5_r_3,blif_clk_net_5_r_4,n4_4,G78_5_r_3,);
nand I_5(n_576_5_r_3,n22_3,n23_3);
not I_6(n_102_5_r_3,n39_3);
nand I_7(n_547_5_r_3,n26_3,n27_3);
not I_8(N1372_10_r_3,n36_3);
nor I_9(N1508_10_r_3,n35_3,n36_3);
and I_10(N3_8_l_3,IN_6_8_l_3,n34_3);
DFFARX1 I_11(N3_8_l_3,blif_clk_net_5_r_4,n4_4,n39_3,);
nand I_12(n_431_5_r_3,n29_3,n30_3);
nor I_13(n22_3,n24_3,n25_3);
nor I_14(n23_3,IN_3_1_l_3,n39_3);
not I_15(n24_3,n27_3);
nand I_16(n25_3,IN_1_1_l_3,IN_2_1_l_3);
nor I_17(n26_3,n39_3,n28_3);
nor I_18(n27_3,IN_1_8_l_3,IN_3_8_l_3);
not I_19(n28_3,n37_3);
nand I_20(n29_3,N1372_10_r_3,n39_3);
nand I_21(n30_3,n31_3,n32_3);
not I_22(n31_3,n25_3);
not I_23(n32_3,IN_3_1_l_3);
nand I_24(n33_3,n24_3,n25_3);
nand I_25(n34_3,IN_2_8_l_3,IN_3_8_l_3);
nor I_26(n35_3,n27_3,n31_3);
nand I_27(n36_3,n28_3,n38_3);
nand I_28(n37_3,IN_1_10_l_3,IN_2_10_l_3);
or I_29(n38_3,IN_3_10_l_3,IN_4_10_l_3);
nor I_30(N1371_0_r_4,n25_4,n29_4);
nor I_31(N1508_0_r_4,n25_4,n32_4);
nor I_32(N6147_2_r_4,n24_4,n31_4);
or I_33(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_34(n_431_5_r_4,blif_clk_net_5_r_4,n4_4,G78_5_r_4,);
nand I_35(n_576_5_r_4,n22_4,n23_4);
nand I_36(n_102_5_r_4,n34_4,n35_4);
nand I_37(n_547_5_r_4,n26_4,n27_4);
nor I_38(N1507_6_r_4,n27_4,n30_4);
nor I_39(N1508_6_r_4,n30_4,n33_4);
nand I_40(n_431_5_r_4,n_102_5_r_4,n28_4);
not I_41(n4_4,blif_reset_net_5_r_4);
nor I_42(n22_4,n24_4,n25_4);
nor I_43(n23_4,n37_4,N1508_0_r_3);
not I_44(n24_4,n_102_5_r_4);
nand I_45(n25_4,G78_5_r_3,n_576_5_r_3);
nor I_46(n26_4,n23_4,n24_4);
not I_47(n27_4,n25_4);
nand I_48(n28_4,n23_4,n29_4);
nor I_49(n29_4,n25_4,N1371_0_r_3);
not I_50(n30_4,n29_4);
nor I_51(n31_4,N1371_0_r_4,n32_4);
nor I_52(n32_4,n23_4,n29_4);
nand I_53(n33_4,n23_4,n24_4);
nor I_54(n34_4,N6147_3_r_3,N1508_0_r_3);
or I_55(n35_4,n36_4,n_102_5_r_3);
nor I_56(n36_4,N1371_0_r_3,n_547_5_r_3);
or I_57(n37_4,n_429_or_0_5_r_3,N1508_10_r_3);
endmodule


