module test_I16661(I1477,I1470,I14588,I16661);
input I1477,I1470,I14588;
output I16661;
wire I16356,I14667,I14856,I13189,I14777,I14808,I14347,I16240,I16644,I14356,I14650,I14421,I14370;
DFFARX1 I_0(I14356,I1470,I16240,,,I16356,);
and I_1(I14667,I14650,I13189);
nor I_2(I14856,I14808,I14421);
DFFARX1 I_3(I1470,,,I13189,);
or I_4(I14777,I14667,I14588);
DFFARX1 I_5(I1470,I14370,,,I14808,);
DFFARX1 I_6(I14777,I1470,I14370,,,I14347,);
nand I_7(I16661,I16644,I16356);
not I_8(I16240,I1477);
DFFARX1 I_9(I14347,I1470,I16240,,,I16644,);
nand I_10(I14356,I14667,I14856);
DFFARX1 I_11(I1470,I14370,,,I14650,);
DFFARX1 I_12(I1470,I14370,,,I14421,);
not I_13(I14370,I1477);
endmodule


