module test_I3217(I1431,I1477,I1470,I3217);
input I1431,I1477,I1470;
output I3217;
wire I2759,I3200;
not I_0(I2759,I1477);
not I_1(I3217,I3200);
DFFARX1 I_2(I1431,I1470,I2759,,,I3200,);
endmodule


