module test_I16568(I14667,I1477,I14350,I14520,I1470,I16568);
input I14667,I1477,I14350,I14520,I1470;
output I16568;
wire I14362,I14344,I16469,I16551,I16435,I14715,I16452,I14901,I14537,I14808,I14335,I14359,I14370,I16534,I16240,I14825;
DFFARX1 I_0(I14825,I1470,I14370,,,I14362,);
nand I_1(I14344,I14537,I14715);
DFFARX1 I_2(I16452,I1470,I16240,,,I16469,);
and I_3(I16551,I16534,I14344);
nand I_4(I16435,I14359,I14350);
not I_5(I14715,I14667);
and I_6(I16452,I16435,I14362);
DFFARX1 I_7(I14808,I1470,I14370,,,I14901,);
DFFARX1 I_8(I14520,I1470,I14370,,,I14537,);
DFFARX1 I_9(I1470,I14370,,,I14808,);
and I_10(I14335,I14808,I14901);
nor I_11(I14359,I14667);
not I_12(I14370,I1477);
nor I_13(I16568,I16551,I16469);
DFFARX1 I_14(I14335,I1470,I16240,,,I16534,);
not I_15(I16240,I1477);
and I_16(I14825,I14808);
endmodule


