module test_I14605(I1477,I13296,I13168,I1470,I13508,I14605);
input I1477,I13296,I13168,I1470,I13508;
output I14605;
wire I13177,I13180,I14503,I14455,I13601,I13186,I14537,I14370,I13197,I13542,I14520,I13159,I14438,I13697,I14472,I13174;
nand I_0(I13177,I13296,I13542);
not I_1(I13180,I13508);
nand I_2(I14503,I13180,I13168);
DFFARX1 I_3(I13177,I1470,I14370,,,I14455,);
and I_4(I14605,I14537,I14472);
DFFARX1 I_5(I1470,I13197,,,I13601,);
nor I_6(I13186,I13601,I13508);
DFFARX1 I_7(I14520,I1470,I14370,,,I14537,);
not I_8(I14370,I1477);
not I_9(I13197,I1477);
nor I_10(I13542,I13508);
and I_11(I14520,I14503,I13174);
DFFARX1 I_12(I13508,I1470,I13197,,,I13159,);
nor I_13(I14438,I13159,I13186);
or I_14(I13697,I13296);
nand I_15(I14472,I14455,I14438);
DFFARX1 I_16(I13697,I1470,I13197,,,I13174,);
endmodule


