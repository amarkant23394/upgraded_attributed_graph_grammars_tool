module test_I13746(I1477,I1470,I13746);
input I1477,I1470;
output I13746;
wire I14083,I11956,I12349,I13775,I14049,I11962,I14066;
DFFARX1 I_0(I14066,I1470,I13775,,,I14083,);
not I_1(I11956,I12349);
DFFARX1 I_2(I1470,,,I12349,);
not I_3(I13746,I14083);
not I_4(I13775,I1477);
DFFARX1 I_5(I11962,I1470,I13775,,,I14049,);
nor I_6(I11962,I12349);
and I_7(I14066,I14049,I11956);
endmodule


