module test_I3538(I1477,I1215,I1423,I2038,I1470,I1207,I1535,I3538);
input I1477,I1215,I1423,I2038,I1470,I1207,I1535;
output I3538;
wire I1518,I1668,I1637,I2072,I1586,I1510,I1603,I1832,I2055,I1492;
not I_0(I1518,I1477);
not I_1(I1668,I1637);
not I_2(I1637,I1215);
and I_3(I2072,I1832,I2055);
nor I_4(I1586,I1535,I1215);
nor I_5(I3538,I1492,I1510);
DFFARX1 I_6(I2072,I1470,I1518,,,I1510,);
nand I_7(I1603,I1586,I1423);
nand I_8(I1832,I1535,I1207);
nand I_9(I2055,I2038,I1603);
nand I_10(I1492,I1603,I1668);
endmodule


