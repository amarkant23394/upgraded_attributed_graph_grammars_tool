module test_I13761(I12380,I11947,I12304,I1477,I1470,I12058,I13761);
input I12380,I11947,I12304,I1477,I1470,I12058;
output I13761;
wire I13826,I13860,I13792,I13891,I13775,I13809,I13843,I12075,I11973,I11959,I11965,I11944;
DFFARX1 I_0(I13809,I1470,I13775,,,I13826,);
nand I_1(I13761,I13891,I13860);
nor I_2(I13860,I13843,I13826);
nand I_3(I13792,I11965);
DFFARX1 I_4(I11944,I1470,I13775,,,I13891,);
not I_5(I13775,I1477);
and I_6(I13809,I13792,I11947);
nor I_7(I13843,I11959,I11965);
DFFARX1 I_8(I12058,I1470,I11973,,,I12075,);
not I_9(I11973,I1477);
nand I_10(I11959,I12058,I12380);
DFFARX1 I_11(I12304,I1470,I11973,,,I11965,);
not I_12(I11944,I12075);
endmodule


