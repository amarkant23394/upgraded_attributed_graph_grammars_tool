module test_I6887(I1477,I5070,I1470,I5642,I6887);
input I1477,I5070,I1470,I5642;
output I6887;
wire I5594,I7427,I7317,I7026,I7057,I5067,I7410,I6907,I7269,I5105,I5082;
DFFARX1 I_0(I1470,I5105,,,I5594,);
not I_1(I7427,I7410);
nor I_2(I7317,I7269,I7057);
not I_3(I7026,I5070);
not I_4(I7057,I7026);
DFFARX1 I_5(I5642,I1470,I5105,,,I5067,);
DFFARX1 I_6(I5082,I1470,I6907,,,I7410,);
not I_7(I6907,I1477);
DFFARX1 I_8(I5067,I1470,I6907,,,I7269,);
nand I_9(I6887,I7427,I7317);
not I_10(I5105,I1477);
not I_11(I5082,I5594);
endmodule


