module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_7_r_3,n10_3,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
not I_36(N1372_1_r_3,n40_3);
nor I_37(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_38(N1507_6_r_3,n31_3,n42_3);
nor I_39(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_40(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_41(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_42(n_573_7_r_3,n30_3,n31_3);
nor I_43(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_44(n_569_7_r_3,n30_3,n32_3);
nor I_45(n_452_7_r_3,n35_3,N1372_1_r_5);
not I_46(N6147_9_r_3,n32_3);
nor I_47(N6134_9_r_3,n36_3,n37_3);
not I_48(I_BUFF_1_9_r_3,n45_3);
nor I_49(n4_7_r_3,I_BUFF_1_9_r_3,N1372_1_r_5);
not I_50(n10_3,blif_reset_net_7_r_3);
not I_51(n30_3,n39_3);
not I_52(n31_3,n35_3);
nand I_53(n32_3,n41_3,N1507_6_r_5);
nor I_54(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_55(n34_3,n46_3,n_573_7_r_5);
nor I_56(n35_3,n43_3,n44_3);
not I_57(n36_3,n34_3);
nor I_58(n37_3,N6147_9_r_3,N1372_1_r_5);
or I_59(n38_3,n_572_7_r_3,n34_3);
nor I_60(n39_3,n44_3,N6147_2_r_5);
nand I_61(n40_3,n39_3,N1372_1_r_5);
nand I_62(n41_3,n_569_7_r_5,N1508_0_r_5);
nor I_63(n42_3,n34_3,n45_3);
not I_64(n43_3,n_572_7_r_5);
nor I_65(n44_3,N1508_0_r_5,G42_7_r_5);
nand I_66(n45_3,n49_3,n50_3);
and I_67(n46_3,n47_3,N1371_0_r_5);
nand I_68(n47_3,n41_3,n48_3);
not I_69(n48_3,N1507_6_r_5);
nor I_70(n49_3,N1508_6_r_5,n_452_7_r_5);
or I_71(n50_3,n51_3,N1372_1_r_5);
nor I_72(n51_3,N1371_0_r_5,N1508_1_r_5);
endmodule


