module test_I1902(I1704,I2138,I1294,I1492,I1301,I1902);
input I1704,I2138,I1294,I1492,I1301;
output I1902;
wire I2172,I1322,I2203,I2234,I1937,I1342,I2155,I1427,I1509,I1304,I1954,I1313;
DFFARX1 I_0(I2155,I1294,I1937,,,I2172,);
nand I_1(I1322,I1427,I1704);
and I_2(I1902,I2234,I2203);
DFFARX1 I_3(I2172,I1294,I1937,,,I2203,);
nand I_4(I2234,I1954,I1304);
not I_5(I1937,I1301);
not I_6(I1342,I1301);
or I_7(I2155,I2138,I1313);
DFFARX1 I_8(I1294,I1342,,,I1427,);
DFFARX1 I_9(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_10(I1509,I1294,I1342,,,I1304,);
not I_11(I1954,I1322);
DFFARX1 I_12(I1427,I1294,I1342,,,I1313,);
endmodule


