module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_5_r_9,n10_9,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_5_r_9,n10_9,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
nor I_40(N6147_2_r_9,n62_9,n46_9);
not I_41(N1372_4_r_9,n59_9);
nor I_42(N1508_4_r_9,n58_9,n59_9);
nand I_43(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_44(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_45(n_576_5_r_9,n39_9,n40_9);
not I_46(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_47(n_547_5_r_9,n43_9,N6147_9_r_8);
and I_48(n_42_8_r_9,n44_9,n_42_8_r_8);
DFFARX1 I_49(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_50(N6147_9_r_9,n41_9,n45_9);
nor I_51(N6134_9_r_9,n45_9,n51_9);
nor I_52(I_BUFF_1_9_r_9,n41_9,N6147_9_r_8);
nor I_53(n4_7_l_9,N1508_1_r_8,n_42_8_r_8);
not I_54(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_55(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_56(N3_8_l_9,n57_9,N1508_6_r_8);
DFFARX1 I_57(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_58(n38_9,n63_9);
nor I_59(n_431_5_r_9,n_42_8_r_8,N6134_9_r_8);
nor I_60(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_61(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_62(n40_9,n41_9);
nand I_63(n41_9,N1371_0_r_8,N1507_6_r_8);
nor I_64(n42_9,N1508_1_r_8,G199_8_r_8);
nor I_65(n43_9,n63_9,n41_9);
nor I_66(n44_9,N1508_1_r_8,N1508_6_r_8);
and I_67(n45_9,n52_9,N1507_6_r_8);
nor I_68(n46_9,n47_9,n48_9);
nor I_69(n47_9,n49_9,n50_9);
not I_70(n48_9,n_429_or_0_5_r_9);
not I_71(n49_9,n42_9);
or I_72(n50_9,n63_9,n51_9);
nor I_73(n51_9,N1371_0_r_8,N1508_10_r_8);
nor I_74(n52_9,n49_9,n_42_8_r_8);
nor I_75(n53_9,n54_9,n55_9);
nor I_76(n54_9,n56_9,n_42_8_r_8);
or I_77(n55_9,n44_9,G199_8_r_8);
not I_78(n56_9,N1507_6_r_8);
nand I_79(n57_9,N1508_10_r_8,G199_8_r_8);
nor I_80(n58_9,n62_9,n60_9);
nand I_81(n59_9,n51_9,n61_9);
nor I_82(n60_9,n38_9,n44_9);
nor I_83(n61_9,N1508_6_r_8,n_42_8_r_8);
endmodule


