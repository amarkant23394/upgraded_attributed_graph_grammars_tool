module test_I5659(I3470,I5187,I1477,I3353,I1470,I5659);
input I3470,I5187,I1477,I3353,I1470;
output I5659;
wire I3368,I5546,I5625,I5204,I5563,I3377,I5529,I5512,I3747,I5105,I5642;
or I_0(I5659,I5642,I5563);
nand I_1(I3368,I3747,I3470);
nor I_2(I5546,I5204,I5529);
DFFARX1 I_3(I3377,I1470,I5105,,,I5625,);
nand I_4(I5204,I5187,I3353);
and I_5(I5563,I5512,I5546);
not I_6(I3377,I3747);
not I_7(I5529,I5512);
DFFARX1 I_8(I3368,I1470,I5105,,,I5512,);
DFFARX1 I_9(I1470,,,I3747,);
not I_10(I5105,I1477);
not I_11(I5642,I5625);
endmodule


