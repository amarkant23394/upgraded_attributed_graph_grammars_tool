module test_I10202(I1477,I7587,I1470,I10202);
input I1477,I7587,I1470;
output I10202;
wire I8107,I6297,I7562,I7652,I7547,I7570,I8090,I7816,I10185,I6380,I7541,I8059,I6318,I7833,I7977,I7669;
not I_0(I8107,I8090);
DFFARX1 I_1(I1470,,,I6297,);
nand I_2(I7562,I8107,I7833);
nor I_3(I7652,I7587,I6297);
not I_4(I7547,I8059);
not I_5(I7570,I1477);
DFFARX1 I_6(I1470,I7570,,,I8090,);
DFFARX1 I_7(I1470,I7570,,,I7816,);
nand I_8(I10185,I7547,I7562);
DFFARX1 I_9(I1470,,,I6380,);
DFFARX1 I_10(I7669,I1470,I7570,,,I7541,);
DFFARX1 I_11(I7977,I1470,I7570,,,I8059,);
not I_12(I6318,I6380);
nor I_13(I7833,I7816,I7669);
and I_14(I10202,I10185,I7541);
DFFARX1 I_15(I1470,I7570,,,I7977,);
nand I_16(I7669,I7652,I6318);
endmodule


