module test_I1959(I1463,I1477,I1215,I1470,I1399,I1383,I1959);
input I1463,I1477,I1215,I1470,I1399,I1383;
output I1959;
wire I1518,I1552,I1880,I1569;
not I_0(I1518,I1477);
nor I_1(I1552,I1215,I1399);
DFFARX1 I_2(I1383,I1470,I1518,,,I1880,);
nand I_3(I1569,I1552,I1463);
nand I_4(I1959,I1880,I1569);
endmodule


