module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_7_r_16,n8_16,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N1371_0_r_16,n35_16,n39_16);
nor I_37(N1508_0_r_16,n39_16,n46_16);
not I_38(N1372_1_r_16,n45_16);
nor I_39(N1508_1_r_16,n53_16,n45_16);
nor I_40(N6147_2_r_16,n37_16,n38_16);
nor I_41(N1507_6_r_16,n44_16,n49_16);
nor I_42(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_43(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_44(n_572_7_r_16,n32_16,n33_16);
nand I_45(n_573_7_r_16,n30_16,n31_16);
nand I_46(n_549_7_r_16,n47_16,N1508_6_r_5);
nand I_47(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_48(n_452_7_r_16,n34_16,n35_16);
and I_49(N3_8_l_16,n41_16,N6147_2_r_5);
not I_50(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_51(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_52(n29_16,n53_16);
nor I_53(n4_7_r_16,n35_16,n36_16);
nand I_54(n30_16,n_452_7_r_5,N1371_0_r_5);
not I_55(n31_16,n34_16);
nor I_56(n32_16,n30_16,G42_7_r_5);
not I_57(n33_16,n_549_7_r_16);
nor I_58(n34_16,n48_16,n_572_7_r_5);
and I_59(n35_16,n50_16,N1371_0_r_5);
not I_60(n36_16,n30_16);
nor I_61(n37_16,n31_16,n40_16);
nand I_62(n38_16,n29_16,n39_16);
not I_63(n39_16,n32_16);
nor I_64(n40_16,N1372_1_r_5,N1508_1_r_5);
nand I_65(n41_16,N1508_1_r_5,N1372_1_r_5);
nand I_66(n42_16,n35_16,n43_16);
not I_67(n43_16,n44_16);
nor I_68(n44_16,n32_16,n49_16);
nand I_69(n45_16,n36_16,n40_16);
nor I_70(n46_16,n33_16,n34_16);
nand I_71(n47_16,N1507_6_r_5,n_569_7_r_5);
or I_72(n48_16,n_573_7_r_5,N1508_0_r_5);
and I_73(n49_16,n35_16,n36_16);
and I_74(n50_16,n51_16,N1508_0_r_5);
nand I_75(n51_16,n47_16,n52_16);
not I_76(n52_16,N1508_6_r_5);
endmodule


