module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_15,n4_15,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_15,n4_15,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_15,n4_15,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_15,n4_15,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_15,n4_15,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_15,n4_15,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_15,n4_15,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_34(n_572_1_r_15,n17_15,n19_15);
nand I_35(n_573_1_r_15,n15_15,n18_15);
nor I_36(n_549_1_r_15,n21_15,n22_15);
nand I_37(n_569_1_r_15,n15_15,n20_15);
nor I_38(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_39(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_40(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_41(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_42(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_43(n4_1_l_15,G42_1_r_13,n_573_1_r_13);
not I_44(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_45(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_46(n15_15,G42_1_l_15);
DFFARX1 I_47(n_573_1_r_13,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_48(n17_15,n17_internal_15);
DFFARX1 I_49(n_266_and_0_3_r_13,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_50(n_572_1_l_15,n_549_1_r_13,n_452_1_r_13);
DFFARX1 I_51(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_52(n14_15,n14_internal_15);
nand I_53(N1_4_r_15,n25_15,n26_15);
or I_54(n_573_1_l_15,G42_1_r_13,P6_5_r_13);
nor I_55(n18_15,ACVQN1_5_r_13,P6_5_r_13);
nand I_56(n19_15,n27_15,n28_15);
nand I_57(n20_15,n30_15,n_572_1_r_13);
not I_58(n21_15,n20_15);
and I_59(n22_15,n17_15,n_572_1_l_15);
nor I_60(n23_15,G42_1_r_13,n_572_1_r_13);
or I_61(n24_15,ACVQN1_5_r_13,P6_5_r_13);
or I_62(n25_15,n_573_1_l_15,n_572_1_r_13);
nand I_63(n26_15,n19_15,n23_15);
not I_64(n27_15,ACVQN1_5_r_13);
nand I_65(n28_15,n29_15,ACVQN2_3_r_13);
not I_66(n29_15,n_452_1_r_13);
endmodule


