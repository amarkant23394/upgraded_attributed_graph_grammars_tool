module test_I6291(I2733,I2742,I1477,I1470,I6291);
input I2733,I2742,I1477,I1470;
output I6291;
wire I4246,I3948,I6688,I6329,I4263,I4068,I4452,I6705,I2724,I3972,I3983;
DFFARX1 I_0(I1470,I3983,,,I4246,);
DFFARX1 I_1(I4452,I1470,I3983,,,I3948,);
DFFARX1 I_2(I3948,I1470,I6329,,,I6688,);
not I_3(I6329,I1477);
and I_4(I4263,I4246,I2733);
nor I_5(I4068,I2742,I2724);
or I_6(I4452,I4263);
and I_7(I6705,I6688,I3972);
DFFARX1 I_8(I6705,I1470,I6329,,,I6291,);
DFFARX1 I_9(I1470,,,I2724,);
or I_10(I3972,I4263,I4068);
not I_11(I3983,I1477);
endmodule


