module test_I14350(I13183,I1477,I13460,I14387,I1470,I13508,I14350);
input I13183,I1477,I13460,I14387,I1470,I13508;
output I14350;
wire I14667,I13177,I14455,I11302,I14421,I11278,I14715,I14650,I14370,I13542,I13296,I13189,I14404,I14732;
and I_0(I14667,I14650,I13189);
nand I_1(I13177,I13296,I13542);
DFFARX1 I_2(I13177,I1470,I14370,,,I14455,);
DFFARX1 I_3(I1470,,,I11302,);
DFFARX1 I_4(I14404,I1470,I14370,,,I14421,);
DFFARX1 I_5(I1470,,,I11278,);
not I_6(I14715,I14667);
nand I_7(I14350,I14455,I14732);
DFFARX1 I_8(I1470,I14370,,,I14650,);
not I_9(I14370,I1477);
nor I_10(I13542,I13508,I13460);
nor I_11(I13296,I11278,I11302);
DFFARX1 I_12(I1470,,,I13189,);
and I_13(I14404,I14387,I13183);
nor I_14(I14732,I14421,I14715);
endmodule


