module test_I8496(I6265,I1477,I8411,I1470,I8496);
input I6265,I1477,I8411,I1470;
output I8496;
wire I5728,I8428,I8216,I8360,I5751,I8445,I5833,I5734,I5719,I8377,I8462;
not I_0(I5728,I5833);
and I_1(I8428,I8411,I5734);
not I_2(I8216,I1477);
not I_3(I8360,I5719);
not I_4(I5751,I1477);
nor I_5(I8496,I8462,I8377);
or I_6(I8445,I8428,I5728);
DFFARX1 I_7(I1470,I5751,,,I5833,);
DFFARX1 I_8(I1470,I5751,,,I5734,);
DFFARX1 I_9(I6265,I1470,I5751,,,I5719,);
not I_10(I8377,I8360);
DFFARX1 I_11(I8445,I1470,I8216,,,I8462,);
endmodule


