module test_I14667(I13231,I1477,I1470,I14667);
input I13231,I1477,I1470;
output I14667;
wire I13313,I13189,I13601,I13197,I11302,I13165,I14650,I13635,I11278,I13296,I13248,I13618,I14370;
DFFARX1 I_0(I1470,I13197,,,I13313,);
and I_1(I14667,I14650,I13189);
DFFARX1 I_2(I13635,I1470,I13197,,,I13189,);
DFFARX1 I_3(I1470,I13197,,,I13601,);
not I_4(I13197,I1477);
DFFARX1 I_5(I1470,,,I11302,);
DFFARX1 I_6(I13248,I1470,I13197,,,I13165,);
DFFARX1 I_7(I13165,I1470,I14370,,,I14650,);
and I_8(I13635,I13296,I13618);
DFFARX1 I_9(I1470,,,I11278,);
nor I_10(I13296,I11278,I11302);
DFFARX1 I_11(I13231,I1470,I13197,,,I13248,);
nand I_12(I13618,I13601,I13313);
not I_13(I14370,I1477);
endmodule


