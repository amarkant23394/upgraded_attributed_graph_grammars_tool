module test_I13189(I1477,I11299,I11293,I1470,I11624,I13189);
input I1477,I11299,I11293,I1470,I11624;
output I13189;
wire I13313,I13601,I13197,I11302,I13635,I11278,I13296,I11310,I13618,I11864;
DFFARX1 I_0(I11293,I1470,I13197,,,I13313,);
DFFARX1 I_1(I13635,I1470,I13197,,,I13189,);
DFFARX1 I_2(I11299,I1470,I13197,,,I13601,);
not I_3(I13197,I1477);
DFFARX1 I_4(I11864,I1470,I11310,,,I11302,);
and I_5(I13635,I13296,I13618);
DFFARX1 I_6(I11624,I1470,I11310,,,I11278,);
nor I_7(I13296,I11278,I11302);
not I_8(I11310,I1477);
nand I_9(I13618,I13601,I13313);
and I_10(I11864,I11624);
endmodule


