module test_I7604(I3963,I3966,I6346,I1477,I6442,I1470,I7604);
input I3963,I3966,I6346,I1477,I6442,I1470;
output I7604;
wire I6781,I6297,I6826,I6329,I6380,I6843,I6493,I6541,I6363,I6294;
DFFARX1 I_0(I1470,I6329,,,I6781,);
DFFARX1 I_1(I6843,I1470,I6329,,,I6297,);
nand I_2(I6826,I6781,I6442);
nor I_3(I7604,I6297,I6294);
not I_4(I6329,I1477);
DFFARX1 I_5(I6363,I1470,I6329,,,I6380,);
and I_6(I6843,I6493,I6826);
DFFARX1 I_7(I3966,I1470,I6329,,,I6493,);
DFFARX1 I_8(I6493,I1470,I6329,,,I6541,);
and I_9(I6363,I6346,I3963);
and I_10(I6294,I6380,I6541);
endmodule


