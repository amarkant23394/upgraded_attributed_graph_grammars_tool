module test_I11105(I1477,I9559,I1470,I11105);
input I1477,I9559,I1470;
output I11105;
wire I10647,I10698,I11009,I11088,I9816,I10766,I9771,I9480,I8178,I9456,I9491,I9477,I9754,I9468,I10681,I9833,I9960,I9864;
not I_0(I10647,I1477);
and I_1(I11105,I10766,I11088);
nand I_2(I10698,I10681,I9456);
DFFARX1 I_3(I9468,I1470,I10647,,,I11009,);
nand I_4(I11088,I11009,I10698);
DFFARX1 I_5(I1470,I9491,,,I9816,);
not I_6(I10766,I9477);
and I_7(I9771,I9754,I8178);
or I_8(I9480,I9771);
DFFARX1 I_9(I1470,,,I8178,);
DFFARX1 I_10(I9960,I1470,I9491,,,I9456,);
not I_11(I9491,I1477);
nor I_12(I9477,I9771,I9833);
DFFARX1 I_13(I1470,I9491,,,I9754,);
DFFARX1 I_14(I9864,I1470,I9491,,,I9468,);
nor I_15(I10681,I9477,I9480);
and I_16(I9833,I9816,I9559);
or I_17(I9960,I9771);
nor I_18(I9864,I9816);
endmodule


