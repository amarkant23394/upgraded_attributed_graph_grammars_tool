module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_8,n8_8,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_8,n8_8,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_8,n8_8,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_8,n8_8,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_8,n8_8,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_8,n8_8,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_8,n8_8,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_8,n8_8,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_33(n_572_1_r_8,n39_8,n23_8);
and I_34(n_549_1_r_8,n38_8,n23_8);
nand I_35(n_569_1_r_8,n38_8,n24_8);
nor I_36(n_452_1_r_8,n25_8,n26_8);
nor I_37(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_38(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_39(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_40(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_41(n_431_0_l_8,n29_8,P6_5_r_16);
not I_42(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_43(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_44(n19_8,G78_0_l_8);
DFFARX1 I_45(n_569_1_r_16,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_46(n22_8,n39_8);
DFFARX1 I_47(G42_1_r_16,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_48(n4_1_r_8,G78_0_l_8,n33_8);
nor I_49(N3_2_r_8,n22_8,n35_8);
nor I_50(N1_4_r_8,n27_8,n37_8);
nand I_51(n23_8,n32_8,n_572_1_r_16);
not I_52(n24_8,n23_8);
nand I_53(n25_8,n36_8,n_452_1_r_16);
nand I_54(n26_8,n27_8,n28_8);
nor I_55(n27_8,n31_8,ACVQN1_5_r_16);
not I_56(n28_8,G199_4_r_16);
and I_57(n29_8,n30_8,n_573_1_r_16);
nor I_58(n30_8,n31_8,G214_4_r_16);
not I_59(n31_8,n_549_1_r_16);
and I_60(n32_8,n28_8,ACVQN1_5_r_16);
nand I_61(n33_8,n28_8,n34_8);
not I_62(n34_8,n25_8);
nor I_63(n35_8,n34_8,G199_4_r_16);
not I_64(n36_8,G42_1_r_16);
nor I_65(n37_8,n19_8,n38_8);
endmodule


