module test_final(IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_102_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13,n4_7_l_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
nor I_0(N1371_0_r_13,n59_13,n61_13);
nor I_1(N1508_0_r_13,n59_13,n60_13);
not I_2(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_3(n_431_5_r_13,blif_clk_net_5_r_7,n6_7,G78_5_r_13,);
nand I_4(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_5(n_102_5_r_13,IN_9_7_l_13,IN_10_7_l_13);
nand I_6(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_7(n1_13,blif_clk_net_5_r_7,n6_7,G42_7_r_13,);
nor I_8(n_572_7_r_13,n40_13,n41_13);
nand I_9(n_573_7_r_13,n37_13,n38_13);
nor I_10(n_549_7_r_13,n46_13,n47_13);
nand I_11(n_569_7_r_13,n37_13,n43_13);
nand I_12(n_452_7_r_13,n52_13,n53_13);
nor I_13(n4_7_l_13,G18_7_l_13,IN_1_7_l_13);
DFFARX1 I_14(n4_7_l_13,blif_clk_net_5_r_7,n6_7,n62_13,);
not I_15(n33_13,n62_13);
nand I_16(n_431_5_r_13,n54_13,n55_13);
not I_17(n1_13,n52_13);
nor I_18(n34_13,n35_13,n36_13);
nor I_19(n35_13,G15_7_l_13,n42_13);
nand I_20(n36_13,n50_13,n58_13);
nand I_21(n37_13,n44_13,n45_13);
or I_22(n38_13,IN_3_1_l_13,n39_13);
nand I_23(n39_13,IN_1_1_l_13,IN_2_1_l_13);
not I_24(n40_13,n36_13);
nor I_25(n41_13,IN_10_7_l_13,n35_13);
not I_26(n42_13,IN_4_7_l_13);
or I_27(n43_13,G18_7_l_13,IN_5_7_l_13);
not I_28(n44_13,G15_7_l_13);
not I_29(n45_13,IN_7_7_l_13);
nor I_30(n46_13,n39_13,n40_13);
nor I_31(n47_13,G18_7_l_13,IN_5_7_l_13);
nor I_32(n48_13,n50_13,n51_13);
nor I_33(n49_13,G15_7_l_13,IN_7_7_l_13);
not I_34(n50_13,n59_13);
not I_35(n51_13,n_102_5_r_13);
nand I_36(n52_13,n33_13,n39_13);
nand I_37(n53_13,IN_3_1_l_13,n33_13);
nor I_38(n54_13,IN_5_7_l_13,IN_9_7_l_13);
nand I_39(n55_13,n62_13,n56_13);
nor I_40(n56_13,n39_13,n57_13);
not I_41(n57_13,G18_7_l_13);
or I_42(n58_13,IN_3_10_l_13,IN_4_10_l_13);
nand I_43(n59_13,IN_1_10_l_13,IN_2_10_l_13);
nor I_44(n60_13,IN_5_7_l_13,n51_13);
nor I_45(n61_13,IN_3_1_l_13,n39_13);
nor I_46(N1371_0_r_7,n53_7,n52_7);
nor I_47(N1508_0_r_7,n51_7,n52_7);
nand I_48(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_49(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_50(n_576_5_r_7,n31_7,n32_7);
nor I_51(n_102_5_r_7,n_549_7_r_13,N1371_0_r_13);
nand I_52(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_53(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_54(n_572_7_r_7,n54_7,n33_7);
nand I_55(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_56(n_549_7_r_7,n53_7,n36_7);
nand I_57(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_58(n_452_7_r_7,n_572_7_r_13,n_569_7_r_13);
nor I_59(n4_7_l_7,n_573_7_r_13,N1508_0_r_13);
not I_60(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_61(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_62(n30_7,n53_7);
and I_63(N3_8_l_7,n50_7,G42_7_r_13);
DFFARX1 I_64(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_65(n_431_5_r_7,n40_7,n41_7);
nor I_66(n4_7_r_7,n54_7,n49_7);
and I_67(n31_7,n_102_5_r_7,n39_7);
not I_68(n32_7,n_573_7_r_13);
nor I_69(n33_7,n34_7,n_576_5_r_13);
and I_70(n34_7,n35_7,N1371_0_r_13);
not I_71(n35_7,G78_5_r_13);
nor I_72(n36_7,n37_7,n_573_7_r_13);
or I_73(n37_7,n54_7,n_549_7_r_13);
or I_74(n38_7,n_429_or_0_5_r_13,n_547_5_r_13);
nor I_75(n39_7,n_452_7_r_7,n_452_7_r_13);
nand I_76(n40_7,n46_7,n47_7);
nand I_77(n41_7,n42_7,n43_7);
nor I_78(n42_7,n44_7,n45_7);
nor I_79(n43_7,n_429_or_0_5_r_13,n_547_5_r_13);
nor I_80(n44_7,N1508_0_r_13,G78_5_r_13);
nor I_81(n45_7,n_576_5_r_13,N1371_0_r_13);
nand I_82(n46_7,n35_7,N1371_0_r_13);
not I_83(n47_7,n_576_5_r_13);
or I_84(n48_7,n_452_7_r_7,n_452_7_r_13);
not I_85(n49_7,n_452_7_r_7);
nand I_86(n50_7,n_429_or_0_5_r_13,G78_5_r_13);
and I_87(n51_7,n_452_7_r_7,n45_7);
not I_88(n52_7,n44_7);
endmodule


