module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_7_r_1,n9_1,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_7_r_1,n9_1,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
and I_40(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_41(N1508_0_r_1,n40_1,n44_1);
nor I_42(N1507_6_r_1,n43_1,n49_1);
nor I_43(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_44(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_45(n_572_7_r_1,n29_1,n30_1);
not I_46(n_573_7_r_1,n_452_7_r_1);
nor I_47(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_48(n_569_7_r_1,n30_1,n31_1);
nor I_49(n_452_7_r_1,n30_1,n32_1);
nor I_50(N6147_9_r_1,n35_1,n36_1);
nand I_51(N6134_9_r_1,n38_1,n39_1);
not I_52(I_BUFF_1_9_r_1,n40_1);
nor I_53(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_54(n9_1,blif_reset_net_7_r_1);
nor I_55(n29_1,n34_1,N1371_0_r_16);
nor I_56(n30_1,n33_1,n34_1);
nor I_57(n31_1,n54_1,N1507_6_r_16);
not I_58(n32_1,n48_1);
nor I_59(n33_1,N1508_1_r_16,n_452_7_r_16);
not I_60(n34_1,N1372_1_r_16);
nor I_61(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_62(n36_1,n29_1);
not I_63(n37_1,n41_1);
nand I_64(n38_1,I_BUFF_1_9_r_1,n_572_7_r_16);
nand I_65(n39_1,n37_1,n40_1);
nand I_66(n40_1,G42_7_r_16,n_569_7_r_16);
nand I_67(n41_1,n52_1,N6147_2_r_16);
or I_68(n42_1,n36_1,n43_1);
nor I_69(n43_1,n32_1,n49_1);
nand I_70(n44_1,n45_1,n46_1);
nand I_71(n45_1,n47_1,n48_1);
not I_72(n46_1,n_572_7_r_16);
not I_73(n47_1,n31_1);
nand I_74(n48_1,n50_1,n_573_7_r_16);
nor I_75(n49_1,n41_1,n47_1);
and I_76(n50_1,n51_1,N1371_0_r_16);
nand I_77(n51_1,n52_1,n53_1);
nand I_78(n52_1,N1508_0_r_16,N1372_1_r_16);
not I_79(n53_1,N6147_2_r_16);
or I_80(n54_1,N1508_6_r_16,N1508_0_r_16);
nor I_81(n55_1,n29_1,n_572_7_r_16);
endmodule


