module test_I5915(I1477,I2328,I2557,I2509,I1470,I2161,I5915);
input I1477,I2328,I2557,I2509,I1470,I2161;
output I5915;
wire I2167,I4629,I2173,I5751,I4595,I4544,I4527,I4561,I4578,I2633;
nand I_0(I2167,I2633,I2328);
nor I_1(I4629,I2167,I2173);
nand I_2(I2173,I2557,I2509);
not I_3(I5751,I1477);
DFFARX1 I_4(I4578,I1470,I4544,,,I4595,);
not I_5(I4544,I1477);
or I_6(I4527,I4629,I4595);
nand I_7(I4561,I2173);
DFFARX1 I_8(I4527,I1470,I5751,,,I5915,);
and I_9(I4578,I4561,I2161);
DFFARX1 I_10(I1470,,,I2633,);
endmodule


