module test_I8184(I1477,I8445,I6127,I1470,I8184);
input I1477,I8445,I6127,I1470;
output I8184;
wire I8527,I8233,I8216,I5751,I5713,I8544,I8561,I5722,I8462;
nand I_0(I8527,I8233,I5713);
not I_1(I8233,I5722);
not I_2(I8216,I1477);
not I_3(I5751,I1477);
DFFARX1 I_4(I6127,I1470,I5751,,,I5713,);
nand I_5(I8544,I8527,I8462);
DFFARX1 I_6(I8561,I1470,I8216,,,I8184,);
and I_7(I8561,I8527,I8544);
DFFARX1 I_8(I1470,I5751,,,I5722,);
DFFARX1 I_9(I8445,I1470,I8216,,,I8462,);
endmodule


