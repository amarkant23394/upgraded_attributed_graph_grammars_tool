module test_I11290(I9320,I1477,I1470,I8848,I11290);
input I9320,I1477,I1470,I8848;
output I11290;
wire I11672,I8854,I11429,I11720,I11813,I8836,I11830,I9179,I9210,I11460,I11310;
DFFARX1 I_0(I8836,I1470,I11310,,,I11672,);
nand I_1(I11290,I11830,I11720);
nor I_2(I8854,I9179,I9320);
not I_3(I11429,I8848);
nor I_4(I11720,I11672,I11460);
DFFARX1 I_5(I8854,I1470,I11310,,,I11813,);
nand I_6(I8836,I9320,I9210);
not I_7(I11830,I11813);
DFFARX1 I_8(I1470,,,I9179,);
nor I_9(I9210,I9179);
not I_10(I11460,I11429);
not I_11(I11310,I1477);
endmodule


