module test_final(G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_14,blif_reset_net_1_r_14,G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14);
input G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_14,blif_reset_net_1_r_14;
output G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14;
wire G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,n_452_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15,n4_1_l_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15,n_452_1_r_14,n4_1_l_14,n3_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14;
DFFARX1 I_0(n_452_1_r_15,blif_clk_net_1_r_14,n3_14,G42_1_r_15,);
and I_1(n_572_1_r_15,n17_15,n19_15);
nand I_2(n_573_1_r_15,n15_15,n18_15);
nor I_3(n_549_1_r_15,n21_15,n22_15);
nand I_4(n_569_1_r_15,n15_15,n20_15);
nor I_5(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_6(G42_1_l_15,blif_clk_net_1_r_14,n3_14,ACVQN2_3_r_15,);
nor I_7(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_8(N1_4_r_15,blif_clk_net_1_r_14,n3_14,G199_4_r_15,);
DFFARX1 I_9(n_573_1_l_15,blif_clk_net_1_r_14,n3_14,G214_4_r_15,);
nor I_10(n4_1_l_15,G18_1_l_15,IN_1_1_l_15);
DFFARX1 I_11(n4_1_l_15,blif_clk_net_1_r_14,n3_14,G42_1_l_15,);
not I_12(n15_15,G42_1_l_15);
DFFARX1 I_13(IN_1_3_l_15,blif_clk_net_1_r_14,n3_14,n17_internal_15,);
not I_14(n17_15,n17_internal_15);
DFFARX1 I_15(IN_2_3_l_15,blif_clk_net_1_r_14,n3_14,n30_15,);
nor I_16(n_572_1_l_15,G15_1_l_15,IN_7_1_l_15);
DFFARX1 I_17(n_572_1_l_15,blif_clk_net_1_r_14,n3_14,n14_internal_15,);
not I_18(n14_15,n14_internal_15);
nand I_19(N1_4_r_15,n25_15,n26_15);
or I_20(n_573_1_l_15,IN_5_1_l_15,IN_9_1_l_15);
nor I_21(n18_15,IN_9_1_l_15,IN_10_1_l_15);
nand I_22(n19_15,n27_15,n28_15);
nand I_23(n20_15,IN_4_3_l_15,n30_15);
not I_24(n21_15,n20_15);
and I_25(n22_15,n17_15,n_572_1_l_15);
nor I_26(n23_15,G18_1_l_15,IN_5_1_l_15);
or I_27(n24_15,IN_9_1_l_15,IN_10_1_l_15);
or I_28(n25_15,G18_1_l_15,n_573_1_l_15);
nand I_29(n26_15,n19_15,n23_15);
not I_30(n27_15,IN_10_1_l_15);
nand I_31(n28_15,IN_4_1_l_15,n29_15);
not I_32(n29_15,G15_1_l_15);
DFFARX1 I_33(n_452_1_r_14,blif_clk_net_1_r_14,n3_14,G42_1_r_14,);
and I_34(n_572_1_r_14,n18_14,n19_14);
nand I_35(n_573_1_r_14,n16_14,n17_14);
nor I_36(n_549_1_r_14,n20_14,n21_14);
or I_37(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_38(n_452_1_r_14,n23_14,G42_1_r_15);
nor I_39(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_40(N3_2_r_14,blif_clk_net_1_r_14,n3_14,G199_2_r_14,);
DFFARX1 I_41(n_572_1_l_14,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_14,);
not I_42(P6_5_r_14,P6_5_r_internal_14);
nor I_43(n4_1_l_14,G42_1_r_15,n_569_1_r_15);
not I_44(n3_14,blif_reset_net_1_r_14);
DFFARX1 I_45(n4_1_l_14,blif_clk_net_1_r_14,n3_14,n15_internal_14,);
not I_46(n15_14,n15_internal_14);
DFFARX1 I_47(n_573_1_r_15,blif_clk_net_1_r_14,n3_14,ACVQN2_3_l_14,);
DFFARX1 I_48(n_266_and_0_3_r_15,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_14,);
and I_49(N3_2_r_14,n26_14,n27_14);
nor I_50(n_572_1_l_14,n_549_1_r_15,ACVQN2_3_r_15);
DFFARX1 I_51(ACVQN2_3_l_14,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_14,);
nor I_52(n16_14,G199_4_r_15,G42_1_r_15);
not I_53(n17_14,n_572_1_l_14);
nor I_54(n18_14,G199_4_r_15,G214_4_r_15);
nand I_55(n19_14,ACVQN1_3_l_14,n_572_1_r_15);
nor I_56(n20_14,n_569_1_r_15,G214_4_r_15);
nor I_57(n21_14,n15_14,n22_14);
nand I_58(n22_14,n24_14,n25_14);
nand I_59(n23_14,n15_14,n24_14);
not I_60(n24_14,G199_4_r_15);
not I_61(n25_14,G214_4_r_15);
nor I_62(n26_14,n20_14,G42_1_r_15);
nand I_63(n27_14,n28_14,n_572_1_r_15);
not I_64(n28_14,ACVQN2_3_r_15);
endmodule


