module test_I1325(I1215,I1294,I1301,I1325);
input I1215,I1294,I1301;
output I1325;
wire I1342,I1780;
not I_0(I1325,I1780);
not I_1(I1342,I1301);
DFFARX1 I_2(I1215,I1294,I1342,,,I1780,);
endmodule


