module Benchmark_testing10000(I1365,I1373,I1381,I1389,I1397,I1405,I1413,I1421,I1429,I1437,I1445,I1453,I1461,I1469,I1477,I1485,I1493,I1501,I1509,I1517,I1525,I1533,I1541,I1549,I1557,I1565,I1573,I1581,I1589,I1597,I1605,I1613,I1621,I1629,I1637,I1645,I1653,I1661,I1669,I1677,I1685,I1693,I1701,I1709,I1717,I1725,I1733,I1741,I1749,I1757,I1765,I1773,I1781,I1789,I1797,I1805,I1813,I1821,I1829,I1837,I1845,I1853,I1861,I1869,I1877,I1885,I1892,I1899,I9941,I9951,I9961,I9971,I9981,I9991,I10001,I10011,I10021,I10031,I18018,I18028,I18038,I18048,I18058,I18068,I18078,I18088,I18098,I26007,I26017,I26027,I26037,I26047,I26057,I26067,I26077,I26087,I34022,I34032,I34042,I34052,I34062,I34072,I34082,I34092,I34102,I42115,I42125,I42135,I42145,I42155,I42165,I42175,I42185,I42195,I50172,I50182,I50192,I50202,I50212,I50222,I50232,I50242,I50252,I50262);
input I1365,I1373,I1381,I1389,I1397,I1405,I1413,I1421,I1429,I1437,I1445,I1453,I1461,I1469,I1477,I1485,I1493,I1501,I1509,I1517,I1525,I1533,I1541,I1549,I1557,I1565,I1573,I1581,I1589,I1597,I1605,I1613,I1621,I1629,I1637,I1645,I1653,I1661,I1669,I1677,I1685,I1693,I1701,I1709,I1717,I1725,I1733,I1741,I1749,I1757,I1765,I1773,I1781,I1789,I1797,I1805,I1813,I1821,I1829,I1837,I1845,I1853,I1861,I1869,I1877,I1885,I1892,I1899;
output I9941,I9951,I9961,I9971,I9981,I9991,I10001,I10011,I10021,I10031,I18018,I18028,I18038,I18048,I18058,I18068,I18078,I18088,I18098,I26007,I26017,I26027,I26037,I26047,I26057,I26067,I26077,I26087,I34022,I34032,I34042,I34052,I34062,I34072,I34082,I34092,I34102,I42115,I42125,I42135,I42145,I42155,I42165,I42175,I42185,I42195,I50172,I50182,I50192,I50202,I50212,I50222,I50232,I50242,I50252,I50262;
wire I1365,I1373,I1381,I1389,I1397,I1405,I1413,I1421,I1429,I1437,I1445,I1453,I1461,I1469,I1477,I1485,I1493,I1501,I1509,I1517,I1525,I1533,I1541,I1549,I1557,I1565,I1573,I1581,I1589,I1597,I1605,I1613,I1621,I1629,I1637,I1645,I1653,I1661,I1669,I1677,I1685,I1693,I1701,I1709,I1717,I1725,I1733,I1741,I1749,I1757,I1765,I1773,I1781,I1789,I1797,I1805,I1813,I1821,I1829,I1837,I1845,I1853,I1861,I1869,I1877,I1885,I1892,I1899,I1909,I1919,I1929,I1939,I1949,I1959,I1969,I1979,I1989,I1999,I2009,I2049,I2052,I2055,I2058,I2061,I2064,I2067,I2070,I2073,I2076,I2092,I2102,I2112,I2122,I2132,I2142,I2152,I2162,I2172,I2182,I2222,I2225,I2228,I2231,I2234,I2237,I2240,I2243,I2246,I2262,I2272,I2282,I2292,I2302,I2312,I2322,I2332,I2342,I2382,I2385,I2388,I2391,I2394,I2397,I2400,I2403,I2406,I2422,I2432,I2442,I2452,I2462,I2472,I2482,I2492,I2502,I2542,I2545,I2548,I2551,I2554,I2557,I2560,I2563,I2566,I2569,I2585,I2595,I2605,I2615,I2625,I2635,I2645,I2655,I2665,I2675,I2715,I2718,I2721,I2724,I2727,I2730,I2733,I2736,I2739,I2755,I2765,I2775,I2785,I2795,I2805,I2815,I2825,I2835,I2875,I2878,I2881,I2884,I2887,I2890,I2893,I2896,I2899,I2902,I2918,I2928,I2938,I2948,I2958,I2968,I2978,I2988,I2998,I3008,I3048,I3051,I3054,I3057,I3060,I3063,I3066,I3069,I3072,I3088,I3098,I3108,I3118,I3128,I3138,I3148,I3158,I3168,I3208,I3211,I3214,I3217,I3220,I3223,I3226,I3229,I3232,I3248,I3258,I3268,I3278,I3288,I3298,I3308,I3318,I3328,I3368,I3371,I3374,I3377,I3380,I3383,I3386,I3389,I3392,I3395,I3411,I3421,I3431,I3441,I3451,I3461,I3471,I3481,I3491,I3501,I3541,I3544,I3547,I3550,I3553,I3556,I3559,I3562,I3565,I3581,I3591,I3601,I3611,I3621,I3631,I3641,I3651,I3661,I3701,I3704,I3707,I3710,I3713,I3716,I3719,I3722,I3725,I3728,I3744,I3754,I3764,I3774,I3784,I3794,I3804,I3814,I3824,I3834,I3874,I3877,I3880,I3883,I3886,I3889,I3892,I3895,I3911,I3921,I3931,I3941,I3951,I3961,I3971,I3981,I4021,I4024,I4027,I4030,I4033,I4036,I4039,I4042,I4045,I4061,I4071,I4081,I4091,I4101,I4111,I4121,I4131,I4141,I4181,I4184,I4187,I4190,I4193,I4196,I4199,I4202,I4205,I4208,I4224,I4234,I4244,I4254,I4264,I4274,I4284,I4294,I4304,I4314,I4354,I4357,I4360,I4363,I4366,I4369,I4372,I4375,I4378,I4381,I4397,I4407,I4417,I4427,I4437,I4447,I4457,I4467,I4477,I4487,I4527,I4530,I4533,I4536,I4539,I4542,I4545,I4548,I4564,I4574,I4584,I4594,I4604,I4614,I4624,I4634,I4674,I4677,I4680,I4683,I4686,I4689,I4692,I4695,I4698,I4714,I4724,I4734,I4744,I4754,I4764,I4774,I4784,I4794,I4834,I4837,I4840,I4843,I4846,I4849,I4852,I4855,I4858,I4874,I4884,I4894,I4904,I4914,I4924,I4934,I4944,I4954,I4994,I4997,I5000,I5003,I5006,I5009,I5012,I5015,I5018,I5034,I5044,I5054,I5064,I5074,I5084,I5094,I5104,I5114,I5154,I5157,I5160,I5163,I5166,I5169,I5172,I5175,I5178,I5194,I5204,I5214,I5224,I5234,I5244,I5254,I5264,I5274,I5314,I5317,I5320,I5323,I5326,I5329,I5332,I5335,I5338,I5354,I5364,I5374,I5384,I5394,I5404,I5414,I5424,I5434,I5474,I5477,I5480,I5483,I5486,I5489,I5492,I5495,I5498,I5514,I5524,I5534,I5544,I5554,I5564,I5574,I5584,I5594,I5634,I5637,I5640,I5643,I5646,I5649,I5652,I5655,I5658,I5661,I5677,I5687,I5697,I5707,I5717,I5727,I5737,I5747,I5757,I5767,I5807,I5810,I5813,I5816,I5819,I5822,I5825,I5828,I5831,I5847,I5857,I5867,I5877,I5887,I5897,I5907,I5917,I5927,I5967,I5970,I5973,I5976,I5979,I5982,I5985,I5988,I5991,I6007,I6017,I6027,I6037,I6047,I6057,I6067,I6077,I6087,I6127,I6130,I6133,I6136,I6139,I6142,I6145,I6148,I6151,I6167,I6177,I6187,I6197,I6207,I6217,I6227,I6237,I6247,I6287,I6290,I6293,I6296,I6299,I6302,I6305,I6308,I6311,I6327,I6337,I6347,I6357,I6367,I6377,I6387,I6397,I6407,I6447,I6450,I6453,I6456,I6459,I6462,I6465,I6468,I6471,I6487,I6497,I6507,I6517,I6527,I6537,I6547,I6557,I6567,I6607,I6610,I6613,I6616,I6619,I6622,I6625,I6628,I6631,I6634,I6650,I6660,I6670,I6680,I6690,I6700,I6710,I6720,I6730,I6740,I6780,I6783,I6786,I6789,I6792,I6795,I6798,I6801,I6804,I6807,I6823,I6833,I6843,I6853,I6863,I6873,I6883,I6893,I6903,I6913,I6953,I6956,I6959,I6962,I6965,I6968,I6971,I6974,I6977,I6993,I7003,I7013,I7023,I7033,I7043,I7053,I7063,I7073,I7113,I7116,I7119,I7122,I7125,I7128,I7131,I7134,I7137,I7140,I7156,I7166,I7176,I7186,I7196,I7206,I7216,I7226,I7236,I7246,I7286,I7289,I7292,I7295,I7298,I7301,I7304,I7307,I7310,I7313,I7329,I7339,I7349,I7359,I7369,I7379,I7389,I7399,I7409,I7419,I7459,I7462,I7465,I7468,I7471,I7474,I7477,I7480,I7483,I7486,I7502,I7512,I7522,I7532,I7542,I7552,I7562,I7572,I7582,I7592,I7632,I7635,I7638,I7641,I7644,I7647,I7650,I7653,I7656,I7672,I7682,I7692,I7702,I7712,I7722,I7732,I7742,I7752,I7792,I7795,I7798,I7801,I7804,I7807,I7810,I7813,I7816,I7832,I7842,I7852,I7862,I7872,I7882,I7892,I7902,I7912,I7952,I7955,I7958,I7961,I7964,I7967,I7970,I7973,I7976,I7992,I8002,I8012,I8022,I8032,I8042,I8052,I8062,I8072,I8112,I8115,I8118,I8121,I8124,I8127,I8130,I8133,I8136,I8152,I8162,I8172,I8182,I8192,I8202,I8212,I8222,I8232,I8272,I8275,I8278,I8281,I8284,I8287,I8290,I8293,I8296,I8299,I8315,I8325,I8335,I8345,I8355,I8365,I8375,I8385,I8395,I8405,I8445,I8448,I8451,I8454,I8457,I8460,I8463,I8466,I8469,I8485,I8495,I8505,I8515,I8525,I8535,I8545,I8555,I8565,I8605,I8608,I8611,I8614,I8617,I8620,I8623,I8626,I8629,I8645,I8655,I8665,I8675,I8685,I8695,I8705,I8715,I8725,I8765,I8768,I8771,I8774,I8777,I8780,I8783,I8786,I8789,I8805,I8815,I8825,I8835,I8845,I8855,I8865,I8875,I8885,I8925,I8928,I8931,I8934,I8937,I8940,I8943,I8946,I8949,I8965,I8975,I8985,I8995,I9005,I9015,I9025,I9035,I9045,I9085,I9088,I9091,I9094,I9097,I9100,I9103,I9106,I9109,I9125,I9135,I9145,I9155,I9165,I9175,I9185,I9195,I9205,I9245,I9248,I9251,I9254,I9257,I9260,I9263,I9266,I9269,I9285,I9295,I9305,I9315,I9325,I9335,I9345,I9355,I9365,I9405,I9408,I9411,I9414,I9417,I9420,I9423,I9426,I9429,I9432,I9448,I9458,I9468,I9478,I9488,I9498,I9508,I9518,I9528,I9538,I9578,I9581,I9584,I9587,I9590,I9593,I9596,I9599,I9602,I9618,I9628,I9638,I9648,I9658,I9668,I9678,I9688,I9698,I9738,I9741,I9744,I9747,I9750,I9753,I9756,I9759,I9762,I9778,I9788,I9798,I9808,I9818,I9828,I9838,I9848,I9858,I9898,I9901,I9904,I9907,I9910,I9913,I9916,I9919,I9922,I9925,I10041,I10051,I10061,I10071,I10081,I10091,I10101,I10111,I10121,I10131,I10141,I10181,I10184,I10187,I10190,I10193,I10196,I10199,I10202,I10205,I10221,I10231,I10241,I10251,I10261,I10271,I10281,I10291,I10301,I10341,I10344,I10347,I10350,I10353,I10356,I10359,I10362,I10365,I10381,I10391,I10401,I10411,I10421,I10431,I10441,I10451,I10461,I10501,I10504,I10507,I10510,I10513,I10516,I10519,I10522,I10525,I10541,I10551,I10561,I10571,I10581,I10591,I10601,I10611,I10621,I10661,I10664,I10667,I10670,I10673,I10676,I10679,I10682,I10698,I10708,I10718,I10728,I10738,I10748,I10758,I10768,I10808,I10811,I10814,I10817,I10820,I10823,I10826,I10829,I10832,I10835,I10851,I10861,I10871,I10881,I10891,I10901,I10911,I10921,I10931,I10941,I10981,I10984,I10987,I10990,I10993,I10996,I10999,I11002,I11005,I11021,I11031,I11041,I11051,I11061,I11071,I11081,I11091,I11101,I11141,I11144,I11147,I11150,I11153,I11156,I11159,I11162,I11165,I11168,I11184,I11194,I11204,I11214,I11224,I11234,I11244,I11254,I11264,I11274,I11314,I11317,I11320,I11323,I11326,I11329,I11332,I11335,I11338,I11354,I11364,I11374,I11384,I11394,I11404,I11414,I11424,I11434,I11474,I11477,I11480,I11483,I11486,I11489,I11492,I11495,I11498,I11501,I11517,I11527,I11537,I11547,I11557,I11567,I11577,I11587,I11597,I11607,I11647,I11650,I11653,I11656,I11659,I11662,I11665,I11668,I11671,I11674,I11690,I11700,I11710,I11720,I11730,I11740,I11750,I11760,I11770,I11780,I11820,I11823,I11826,I11829,I11832,I11835,I11838,I11841,I11844,I11860,I11870,I11880,I11890,I11900,I11910,I11920,I11930,I11940,I11980,I11983,I11986,I11989,I11992,I11995,I11998,I12001,I12004,I12020,I12030,I12040,I12050,I12060,I12070,I12080,I12090,I12100,I12140,I12143,I12146,I12149,I12152,I12155,I12158,I12161,I12177,I12187,I12197,I12207,I12217,I12227,I12237,I12247,I12287,I12290,I12293,I12296,I12299,I12302,I12305,I12308,I12311,I12327,I12337,I12347,I12357,I12367,I12377,I12387,I12397,I12407,I12447,I12450,I12453,I12456,I12459,I12462,I12465,I12468,I12471,I12474,I12490,I12500,I12510,I12520,I12530,I12540,I12550,I12560,I12570,I12580,I12620,I12623,I12626,I12629,I12632,I12635,I12638,I12641,I12644,I12660,I12670,I12680,I12690,I12700,I12710,I12720,I12730,I12740,I12780,I12783,I12786,I12789,I12792,I12795,I12798,I12801,I12804,I12820,I12830,I12840,I12850,I12860,I12870,I12880,I12890,I12900,I12940,I12943,I12946,I12949,I12952,I12955,I12958,I12961,I12977,I12987,I12997,I13007,I13017,I13027,I13037,I13047,I13087,I13090,I13093,I13096,I13099,I13102,I13105,I13108,I13111,I13127,I13137,I13147,I13157,I13167,I13177,I13187,I13197,I13207,I13247,I13250,I13253,I13256,I13259,I13262,I13265,I13268,I13271,I13274,I13290,I13300,I13310,I13320,I13330,I13340,I13350,I13360,I13370,I13380,I13420,I13423,I13426,I13429,I13432,I13435,I13438,I13441,I13444,I13460,I13470,I13480,I13490,I13500,I13510,I13520,I13530,I13540,I13580,I13583,I13586,I13589,I13592,I13595,I13598,I13601,I13604,I13607,I13623,I13633,I13643,I13653,I13663,I13673,I13683,I13693,I13703,I13713,I13753,I13756,I13759,I13762,I13765,I13768,I13771,I13774,I13777,I13793,I13803,I13813,I13823,I13833,I13843,I13853,I13863,I13873,I13913,I13916,I13919,I13922,I13925,I13928,I13931,I13934,I13937,I13940,I13956,I13966,I13976,I13986,I13996,I14006,I14016,I14026,I14036,I14046,I14086,I14089,I14092,I14095,I14098,I14101,I14104,I14107,I14110,I14126,I14136,I14146,I14156,I14166,I14176,I14186,I14196,I14206,I14246,I14249,I14252,I14255,I14258,I14261,I14264,I14267,I14283,I14293,I14303,I14313,I14323,I14333,I14343,I14353,I14393,I14396,I14399,I14402,I14405,I14408,I14411,I14414,I14417,I14433,I14443,I14453,I14463,I14473,I14483,I14493,I14503,I14513,I14553,I14556,I14559,I14562,I14565,I14568,I14571,I14574,I14577,I14593,I14603,I14613,I14623,I14633,I14643,I14653,I14663,I14673,I14713,I14716,I14719,I14722,I14725,I14728,I14731,I14734,I14737,I14753,I14763,I14773,I14783,I14793,I14803,I14813,I14823,I14833,I14873,I14876,I14879,I14882,I14885,I14888,I14891,I14894,I14897,I14913,I14923,I14933,I14943,I14953,I14963,I14973,I14983,I14993,I15033,I15036,I15039,I15042,I15045,I15048,I15051,I15054,I15057,I15060,I15076,I15086,I15096,I15106,I15116,I15126,I15136,I15146,I15156,I15166,I15206,I15209,I15212,I15215,I15218,I15221,I15224,I15227,I15230,I15233,I15249,I15259,I15269,I15279,I15289,I15299,I15309,I15319,I15329,I15339,I15379,I15382,I15385,I15388,I15391,I15394,I15397,I15400,I15403,I15419,I15429,I15439,I15449,I15459,I15469,I15479,I15489,I15499,I15539,I15542,I15545,I15548,I15551,I15554,I15557,I15560,I15563,I15566,I15582,I15592,I15602,I15612,I15622,I15632,I15642,I15652,I15662,I15672,I15712,I15715,I15718,I15721,I15724,I15727,I15730,I15733,I15736,I15752,I15762,I15772,I15782,I15792,I15802,I15812,I15822,I15832,I15872,I15875,I15878,I15881,I15884,I15887,I15890,I15893,I15896,I15912,I15922,I15932,I15942,I15952,I15962,I15972,I15982,I15992,I16032,I16035,I16038,I16041,I16044,I16047,I16050,I16053,I16056,I16072,I16082,I16092,I16102,I16112,I16122,I16132,I16142,I16152,I16192,I16195,I16198,I16201,I16204,I16207,I16210,I16213,I16216,I16232,I16242,I16252,I16262,I16272,I16282,I16292,I16302,I16312,I16352,I16355,I16358,I16361,I16364,I16367,I16370,I16373,I16376,I16392,I16402,I16412,I16422,I16432,I16442,I16452,I16462,I16472,I16512,I16515,I16518,I16521,I16524,I16527,I16530,I16533,I16536,I16539,I16555,I16565,I16575,I16585,I16595,I16605,I16615,I16625,I16635,I16645,I16685,I16688,I16691,I16694,I16697,I16700,I16703,I16706,I16709,I16725,I16735,I16745,I16755,I16765,I16775,I16785,I16795,I16805,I16845,I16848,I16851,I16854,I16857,I16860,I16863,I16866,I16869,I16885,I16895,I16905,I16915,I16925,I16935,I16945,I16955,I16965,I17005,I17008,I17011,I17014,I17017,I17020,I17023,I17026,I17029,I17045,I17055,I17065,I17075,I17085,I17095,I17105,I17115,I17125,I17165,I17168,I17171,I17174,I17177,I17180,I17183,I17186,I17189,I17205,I17215,I17225,I17235,I17245,I17255,I17265,I17275,I17285,I17325,I17328,I17331,I17334,I17337,I17340,I17343,I17346,I17349,I17365,I17375,I17385,I17395,I17405,I17415,I17425,I17435,I17445,I17485,I17488,I17491,I17494,I17497,I17500,I17503,I17506,I17509,I17525,I17535,I17545,I17555,I17565,I17575,I17585,I17595,I17605,I17645,I17648,I17651,I17654,I17657,I17660,I17663,I17666,I17669,I17685,I17695,I17705,I17715,I17725,I17735,I17745,I17755,I17765,I17805,I17808,I17811,I17814,I17817,I17820,I17823,I17826,I17829,I17832,I17848,I17858,I17868,I17878,I17888,I17898,I17908,I17918,I17928,I17938,I17978,I17981,I17984,I17987,I17990,I17993,I17996,I17999,I18002,I18108,I18118,I18128,I18138,I18148,I18158,I18168,I18178,I18188,I18198,I18208,I18248,I18251,I18254,I18257,I18260,I18263,I18266,I18269,I18272,I18288,I18298,I18308,I18318,I18328,I18338,I18348,I18358,I18368,I18408,I18411,I18414,I18417,I18420,I18423,I18426,I18429,I18432,I18448,I18458,I18468,I18478,I18488,I18498,I18508,I18518,I18528,I18568,I18571,I18574,I18577,I18580,I18583,I18586,I18589,I18592,I18608,I18618,I18628,I18638,I18648,I18658,I18668,I18678,I18688,I18728,I18731,I18734,I18737,I18740,I18743,I18746,I18749,I18752,I18768,I18778,I18788,I18798,I18808,I18818,I18828,I18838,I18848,I18888,I18891,I18894,I18897,I18900,I18903,I18906,I18909,I18925,I18935,I18945,I18955,I18965,I18975,I18985,I18995,I19035,I19038,I19041,I19044,I19047,I19050,I19053,I19056,I19059,I19075,I19085,I19095,I19105,I19115,I19125,I19135,I19145,I19155,I19195,I19198,I19201,I19204,I19207,I19210,I19213,I19216,I19219,I19222,I19238,I19248,I19258,I19268,I19278,I19288,I19298,I19308,I19318,I19328,I19368,I19371,I19374,I19377,I19380,I19383,I19386,I19389,I19392,I19408,I19418,I19428,I19438,I19448,I19458,I19468,I19478,I19488,I19528,I19531,I19534,I19537,I19540,I19543,I19546,I19549,I19552,I19568,I19578,I19588,I19598,I19608,I19618,I19628,I19638,I19648,I19688,I19691,I19694,I19697,I19700,I19703,I19706,I19709,I19712,I19728,I19738,I19748,I19758,I19768,I19778,I19788,I19798,I19808,I19848,I19851,I19854,I19857,I19860,I19863,I19866,I19869,I19885,I19895,I19905,I19915,I19925,I19935,I19945,I19955,I19995,I19998,I20001,I20004,I20007,I20010,I20013,I20016,I20019,I20035,I20045,I20055,I20065,I20075,I20085,I20095,I20105,I20115,I20155,I20158,I20161,I20164,I20167,I20170,I20173,I20176,I20192,I20202,I20212,I20222,I20232,I20242,I20252,I20262,I20302,I20305,I20308,I20311,I20314,I20317,I20320,I20323,I20326,I20342,I20352,I20362,I20372,I20382,I20392,I20402,I20412,I20422,I20462,I20465,I20468,I20471,I20474,I20477,I20480,I20483,I20486,I20489,I20505,I20515,I20525,I20535,I20545,I20555,I20565,I20575,I20585,I20595,I20635,I20638,I20641,I20644,I20647,I20650,I20653,I20656,I20659,I20662,I20678,I20688,I20698,I20708,I20718,I20728,I20738,I20748,I20758,I20768,I20808,I20811,I20814,I20817,I20820,I20823,I20826,I20829,I20832,I20835,I20851,I20861,I20871,I20881,I20891,I20901,I20911,I20921,I20931,I20941,I20981,I20984,I20987,I20990,I20993,I20996,I20999,I21002,I21005,I21021,I21031,I21041,I21051,I21061,I21071,I21081,I21091,I21101,I21141,I21144,I21147,I21150,I21153,I21156,I21159,I21162,I21165,I21168,I21184,I21194,I21204,I21214,I21224,I21234,I21244,I21254,I21264,I21274,I21314,I21317,I21320,I21323,I21326,I21329,I21332,I21335,I21338,I21354,I21364,I21374,I21384,I21394,I21404,I21414,I21424,I21434,I21474,I21477,I21480,I21483,I21486,I21489,I21492,I21495,I21511,I21521,I21531,I21541,I21551,I21561,I21571,I21581,I21621,I21624,I21627,I21630,I21633,I21636,I21639,I21642,I21645,I21648,I21664,I21674,I21684,I21694,I21704,I21714,I21724,I21734,I21744,I21754,I21794,I21797,I21800,I21803,I21806,I21809,I21812,I21815,I21818,I21834,I21844,I21854,I21864,I21874,I21884,I21894,I21904,I21914,I21954,I21957,I21960,I21963,I21966,I21969,I21972,I21975,I21978,I21994,I22004,I22014,I22024,I22034,I22044,I22054,I22064,I22074,I22114,I22117,I22120,I22123,I22126,I22129,I22132,I22135,I22138,I22141,I22157,I22167,I22177,I22187,I22197,I22207,I22217,I22227,I22237,I22247,I22287,I22290,I22293,I22296,I22299,I22302,I22305,I22308,I22311,I22327,I22337,I22347,I22357,I22367,I22377,I22387,I22397,I22407,I22447,I22450,I22453,I22456,I22459,I22462,I22465,I22468,I22471,I22487,I22497,I22507,I22517,I22527,I22537,I22547,I22557,I22567,I22607,I22610,I22613,I22616,I22619,I22622,I22625,I22628,I22631,I22647,I22657,I22667,I22677,I22687,I22697,I22707,I22717,I22727,I22767,I22770,I22773,I22776,I22779,I22782,I22785,I22788,I22791,I22807,I22817,I22827,I22837,I22847,I22857,I22867,I22877,I22887,I22927,I22930,I22933,I22936,I22939,I22942,I22945,I22948,I22951,I22967,I22977,I22987,I22997,I23007,I23017,I23027,I23037,I23047,I23087,I23090,I23093,I23096,I23099,I23102,I23105,I23108,I23111,I23114,I23130,I23140,I23150,I23160,I23170,I23180,I23190,I23200,I23210,I23220,I23260,I23263,I23266,I23269,I23272,I23275,I23278,I23281,I23284,I23300,I23310,I23320,I23330,I23340,I23350,I23360,I23370,I23380,I23420,I23423,I23426,I23429,I23432,I23435,I23438,I23441,I23457,I23467,I23477,I23487,I23497,I23507,I23517,I23527,I23567,I23570,I23573,I23576,I23579,I23582,I23585,I23588,I23591,I23607,I23617,I23627,I23637,I23647,I23657,I23667,I23677,I23687,I23727,I23730,I23733,I23736,I23739,I23742,I23745,I23748,I23764,I23774,I23784,I23794,I23804,I23814,I23824,I23834,I23874,I23877,I23880,I23883,I23886,I23889,I23892,I23895,I23898,I23914,I23924,I23934,I23944,I23954,I23964,I23974,I23984,I23994,I24034,I24037,I24040,I24043,I24046,I24049,I24052,I24055,I24058,I24061,I24077,I24087,I24097,I24107,I24117,I24127,I24137,I24147,I24157,I24167,I24207,I24210,I24213,I24216,I24219,I24222,I24225,I24228,I24231,I24247,I24257,I24267,I24277,I24287,I24297,I24307,I24317,I24327,I24367,I24370,I24373,I24376,I24379,I24382,I24385,I24388,I24404,I24414,I24424,I24434,I24444,I24454,I24464,I24474,I24514,I24517,I24520,I24523,I24526,I24529,I24532,I24535,I24538,I24554,I24564,I24574,I24584,I24594,I24604,I24614,I24624,I24634,I24674,I24677,I24680,I24683,I24686,I24689,I24692,I24695,I24698,I24714,I24724,I24734,I24744,I24754,I24764,I24774,I24784,I24794,I24834,I24837,I24840,I24843,I24846,I24849,I24852,I24855,I24858,I24861,I24877,I24887,I24897,I24907,I24917,I24927,I24937,I24947,I24957,I24967,I25007,I25010,I25013,I25016,I25019,I25022,I25025,I25028,I25031,I25047,I25057,I25067,I25077,I25087,I25097,I25107,I25117,I25127,I25167,I25170,I25173,I25176,I25179,I25182,I25185,I25188,I25191,I25194,I25210,I25220,I25230,I25240,I25250,I25260,I25270,I25280,I25290,I25300,I25340,I25343,I25346,I25349,I25352,I25355,I25358,I25361,I25364,I25380,I25390,I25400,I25410,I25420,I25430,I25440,I25450,I25460,I25500,I25503,I25506,I25509,I25512,I25515,I25518,I25521,I25524,I25540,I25550,I25560,I25570,I25580,I25590,I25600,I25610,I25620,I25660,I25663,I25666,I25669,I25672,I25675,I25678,I25681,I25697,I25707,I25717,I25727,I25737,I25747,I25757,I25767,I25807,I25810,I25813,I25816,I25819,I25822,I25825,I25828,I25831,I25847,I25857,I25867,I25877,I25887,I25897,I25907,I25917,I25927,I25967,I25970,I25973,I25976,I25979,I25982,I25985,I25988,I25991,I26097,I26107,I26117,I26127,I26137,I26147,I26157,I26167,I26177,I26187,I26197,I26237,I26240,I26243,I26246,I26249,I26252,I26255,I26258,I26261,I26277,I26287,I26297,I26307,I26317,I26327,I26337,I26347,I26357,I26397,I26400,I26403,I26406,I26409,I26412,I26415,I26418,I26421,I26424,I26440,I26450,I26460,I26470,I26480,I26490,I26500,I26510,I26520,I26530,I26570,I26573,I26576,I26579,I26582,I26585,I26588,I26591,I26594,I26610,I26620,I26630,I26640,I26650,I26660,I26670,I26680,I26690,I26730,I26733,I26736,I26739,I26742,I26745,I26748,I26751,I26767,I26777,I26787,I26797,I26807,I26817,I26827,I26837,I26877,I26880,I26883,I26886,I26889,I26892,I26895,I26898,I26914,I26924,I26934,I26944,I26954,I26964,I26974,I26984,I27024,I27027,I27030,I27033,I27036,I27039,I27042,I27045,I27048,I27064,I27074,I27084,I27094,I27104,I27114,I27124,I27134,I27144,I27184,I27187,I27190,I27193,I27196,I27199,I27202,I27205,I27208,I27211,I27227,I27237,I27247,I27257,I27267,I27277,I27287,I27297,I27307,I27317,I27357,I27360,I27363,I27366,I27369,I27372,I27375,I27378,I27381,I27397,I27407,I27417,I27427,I27437,I27447,I27457,I27467,I27477,I27517,I27520,I27523,I27526,I27529,I27532,I27535,I27538,I27554,I27564,I27574,I27584,I27594,I27604,I27614,I27624,I27664,I27667,I27670,I27673,I27676,I27679,I27682,I27685,I27688,I27704,I27714,I27724,I27734,I27744,I27754,I27764,I27774,I27784,I27824,I27827,I27830,I27833,I27836,I27839,I27842,I27845,I27861,I27871,I27881,I27891,I27901,I27911,I27921,I27931,I27971,I27974,I27977,I27980,I27983,I27986,I27989,I27992,I27995,I28011,I28021,I28031,I28041,I28051,I28061,I28071,I28081,I28091,I28131,I28134,I28137,I28140,I28143,I28146,I28149,I28152,I28155,I28171,I28181,I28191,I28201,I28211,I28221,I28231,I28241,I28251,I28291,I28294,I28297,I28300,I28303,I28306,I28309,I28312,I28315,I28318,I28334,I28344,I28354,I28364,I28374,I28384,I28394,I28404,I28414,I28424,I28464,I28467,I28470,I28473,I28476,I28479,I28482,I28485,I28501,I28511,I28521,I28531,I28541,I28551,I28561,I28571,I28611,I28614,I28617,I28620,I28623,I28626,I28629,I28632,I28635,I28638,I28654,I28664,I28674,I28684,I28694,I28704,I28714,I28724,I28734,I28744,I28784,I28787,I28790,I28793,I28796,I28799,I28802,I28805,I28821,I28831,I28841,I28851,I28861,I28871,I28881,I28891,I28931,I28934,I28937,I28940,I28943,I28946,I28949,I28952,I28955,I28971,I28981,I28991,I29001,I29011,I29021,I29031,I29041,I29051,I29091,I29094,I29097,I29100,I29103,I29106,I29109,I29112,I29115,I29118,I29134,I29144,I29154,I29164,I29174,I29184,I29194,I29204,I29214,I29224,I29264,I29267,I29270,I29273,I29276,I29279,I29282,I29285,I29288,I29304,I29314,I29324,I29334,I29344,I29354,I29364,I29374,I29384,I29424,I29427,I29430,I29433,I29436,I29439,I29442,I29445,I29448,I29451,I29467,I29477,I29487,I29497,I29507,I29517,I29527,I29537,I29547,I29557,I29597,I29600,I29603,I29606,I29609,I29612,I29615,I29618,I29621,I29624,I29640,I29650,I29660,I29670,I29680,I29690,I29700,I29710,I29720,I29730,I29770,I29773,I29776,I29779,I29782,I29785,I29788,I29791,I29794,I29810,I29820,I29830,I29840,I29850,I29860,I29870,I29880,I29890,I29930,I29933,I29936,I29939,I29942,I29945,I29948,I29951,I29954,I29970,I29980,I29990,I30000,I30010,I30020,I30030,I30040,I30050,I30090,I30093,I30096,I30099,I30102,I30105,I30108,I30111,I30114,I30130,I30140,I30150,I30160,I30170,I30180,I30190,I30200,I30210,I30250,I30253,I30256,I30259,I30262,I30265,I30268,I30271,I30274,I30290,I30300,I30310,I30320,I30330,I30340,I30350,I30360,I30370,I30410,I30413,I30416,I30419,I30422,I30425,I30428,I30431,I30447,I30457,I30467,I30477,I30487,I30497,I30507,I30517,I30557,I30560,I30563,I30566,I30569,I30572,I30575,I30578,I30581,I30584,I30600,I30610,I30620,I30630,I30640,I30650,I30660,I30670,I30680,I30690,I30730,I30733,I30736,I30739,I30742,I30745,I30748,I30751,I30767,I30777,I30787,I30797,I30807,I30817,I30827,I30837,I30877,I30880,I30883,I30886,I30889,I30892,I30895,I30898,I30901,I30917,I30927,I30937,I30947,I30957,I30967,I30977,I30987,I30997,I31037,I31040,I31043,I31046,I31049,I31052,I31055,I31058,I31061,I31077,I31087,I31097,I31107,I31117,I31127,I31137,I31147,I31157,I31197,I31200,I31203,I31206,I31209,I31212,I31215,I31218,I31221,I31224,I31240,I31250,I31260,I31270,I31280,I31290,I31300,I31310,I31320,I31330,I31370,I31373,I31376,I31379,I31382,I31385,I31388,I31391,I31394,I31410,I31420,I31430,I31440,I31450,I31460,I31470,I31480,I31490,I31530,I31533,I31536,I31539,I31542,I31545,I31548,I31551,I31554,I31570,I31580,I31590,I31600,I31610,I31620,I31630,I31640,I31650,I31690,I31693,I31696,I31699,I31702,I31705,I31708,I31711,I31714,I31730,I31740,I31750,I31760,I31770,I31780,I31790,I31800,I31810,I31850,I31853,I31856,I31859,I31862,I31865,I31868,I31871,I31874,I31890,I31900,I31910,I31920,I31930,I31940,I31950,I31960,I31970,I32010,I32013,I32016,I32019,I32022,I32025,I32028,I32031,I32047,I32057,I32067,I32077,I32087,I32097,I32107,I32117,I32157,I32160,I32163,I32166,I32169,I32172,I32175,I32178,I32181,I32184,I32200,I32210,I32220,I32230,I32240,I32250,I32260,I32270,I32280,I32290,I32330,I32333,I32336,I32339,I32342,I32345,I32348,I32351,I32354,I32357,I32373,I32383,I32393,I32403,I32413,I32423,I32433,I32443,I32453,I32463,I32503,I32506,I32509,I32512,I32515,I32518,I32521,I32524,I32527,I32543,I32553,I32563,I32573,I32583,I32593,I32603,I32613,I32623,I32663,I32666,I32669,I32672,I32675,I32678,I32681,I32684,I32687,I32703,I32713,I32723,I32733,I32743,I32753,I32763,I32773,I32783,I32823,I32826,I32829,I32832,I32835,I32838,I32841,I32844,I32847,I32863,I32873,I32883,I32893,I32903,I32913,I32923,I32933,I32943,I32983,I32986,I32989,I32992,I32995,I32998,I33001,I33004,I33007,I33010,I33026,I33036,I33046,I33056,I33066,I33076,I33086,I33096,I33106,I33116,I33156,I33159,I33162,I33165,I33168,I33171,I33174,I33177,I33180,I33183,I33199,I33209,I33219,I33229,I33239,I33249,I33259,I33269,I33279,I33289,I33329,I33332,I33335,I33338,I33341,I33344,I33347,I33350,I33353,I33369,I33379,I33389,I33399,I33409,I33419,I33429,I33439,I33449,I33489,I33492,I33495,I33498,I33501,I33504,I33507,I33510,I33513,I33529,I33539,I33549,I33559,I33569,I33579,I33589,I33599,I33609,I33649,I33652,I33655,I33658,I33661,I33664,I33667,I33670,I33673,I33676,I33692,I33702,I33712,I33722,I33732,I33742,I33752,I33762,I33772,I33782,I33822,I33825,I33828,I33831,I33834,I33837,I33840,I33843,I33846,I33862,I33872,I33882,I33892,I33902,I33912,I33922,I33932,I33942,I33982,I33985,I33988,I33991,I33994,I33997,I34000,I34003,I34006,I34112,I34122,I34132,I34142,I34152,I34162,I34172,I34182,I34192,I34202,I34212,I34252,I34255,I34258,I34261,I34264,I34267,I34270,I34273,I34276,I34279,I34295,I34305,I34315,I34325,I34335,I34345,I34355,I34365,I34375,I34385,I34425,I34428,I34431,I34434,I34437,I34440,I34443,I34446,I34449,I34465,I34475,I34485,I34495,I34505,I34515,I34525,I34535,I34545,I34585,I34588,I34591,I34594,I34597,I34600,I34603,I34606,I34609,I34625,I34635,I34645,I34655,I34665,I34675,I34685,I34695,I34705,I34745,I34748,I34751,I34754,I34757,I34760,I34763,I34766,I34769,I34785,I34795,I34805,I34815,I34825,I34835,I34845,I34855,I34865,I34905,I34908,I34911,I34914,I34917,I34920,I34923,I34926,I34929,I34945,I34955,I34965,I34975,I34985,I34995,I35005,I35015,I35025,I35065,I35068,I35071,I35074,I35077,I35080,I35083,I35086,I35089,I35105,I35115,I35125,I35135,I35145,I35155,I35165,I35175,I35185,I35225,I35228,I35231,I35234,I35237,I35240,I35243,I35246,I35249,I35265,I35275,I35285,I35295,I35305,I35315,I35325,I35335,I35345,I35385,I35388,I35391,I35394,I35397,I35400,I35403,I35406,I35422,I35432,I35442,I35452,I35462,I35472,I35482,I35492,I35532,I35535,I35538,I35541,I35544,I35547,I35550,I35553,I35556,I35559,I35575,I35585,I35595,I35605,I35615,I35625,I35635,I35645,I35655,I35665,I35705,I35708,I35711,I35714,I35717,I35720,I35723,I35726,I35729,I35745,I35755,I35765,I35775,I35785,I35795,I35805,I35815,I35825,I35865,I35868,I35871,I35874,I35877,I35880,I35883,I35886,I35889,I35892,I35908,I35918,I35928,I35938,I35948,I35958,I35968,I35978,I35988,I35998,I36038,I36041,I36044,I36047,I36050,I36053,I36056,I36059,I36062,I36078,I36088,I36098,I36108,I36118,I36128,I36138,I36148,I36158,I36198,I36201,I36204,I36207,I36210,I36213,I36216,I36219,I36222,I36238,I36248,I36258,I36268,I36278,I36288,I36298,I36308,I36318,I36358,I36361,I36364,I36367,I36370,I36373,I36376,I36379,I36382,I36385,I36401,I36411,I36421,I36431,I36441,I36451,I36461,I36471,I36481,I36491,I36531,I36534,I36537,I36540,I36543,I36546,I36549,I36552,I36555,I36571,I36581,I36591,I36601,I36611,I36621,I36631,I36641,I36651,I36691,I36694,I36697,I36700,I36703,I36706,I36709,I36712,I36715,I36718,I36734,I36744,I36754,I36764,I36774,I36784,I36794,I36804,I36814,I36824,I36864,I36867,I36870,I36873,I36876,I36879,I36882,I36885,I36888,I36904,I36914,I36924,I36934,I36944,I36954,I36964,I36974,I36984,I37024,I37027,I37030,I37033,I37036,I37039,I37042,I37045,I37061,I37071,I37081,I37091,I37101,I37111,I37121,I37131,I37171,I37174,I37177,I37180,I37183,I37186,I37189,I37192,I37208,I37218,I37228,I37238,I37248,I37258,I37268,I37278,I37318,I37321,I37324,I37327,I37330,I37333,I37336,I37339,I37342,I37345,I37361,I37371,I37381,I37391,I37401,I37411,I37421,I37431,I37441,I37451,I37491,I37494,I37497,I37500,I37503,I37506,I37509,I37512,I37528,I37538,I37548,I37558,I37568,I37578,I37588,I37598,I37638,I37641,I37644,I37647,I37650,I37653,I37656,I37659,I37662,I37678,I37688,I37698,I37708,I37718,I37728,I37738,I37748,I37758,I37798,I37801,I37804,I37807,I37810,I37813,I37816,I37819,I37822,I37825,I37841,I37851,I37861,I37871,I37881,I37891,I37901,I37911,I37921,I37931,I37971,I37974,I37977,I37980,I37983,I37986,I37989,I37992,I37995,I37998,I38014,I38024,I38034,I38044,I38054,I38064,I38074,I38084,I38094,I38104,I38144,I38147,I38150,I38153,I38156,I38159,I38162,I38165,I38168,I38184,I38194,I38204,I38214,I38224,I38234,I38244,I38254,I38264,I38304,I38307,I38310,I38313,I38316,I38319,I38322,I38325,I38328,I38344,I38354,I38364,I38374,I38384,I38394,I38404,I38414,I38424,I38464,I38467,I38470,I38473,I38476,I38479,I38482,I38485,I38488,I38491,I38507,I38517,I38527,I38537,I38547,I38557,I38567,I38577,I38587,I38597,I38637,I38640,I38643,I38646,I38649,I38652,I38655,I38658,I38661,I38677,I38687,I38697,I38707,I38717,I38727,I38737,I38747,I38757,I38797,I38800,I38803,I38806,I38809,I38812,I38815,I38818,I38821,I38837,I38847,I38857,I38867,I38877,I38887,I38897,I38907,I38917,I38957,I38960,I38963,I38966,I38969,I38972,I38975,I38978,I38994,I39004,I39014,I39024,I39034,I39044,I39054,I39064,I39104,I39107,I39110,I39113,I39116,I39119,I39122,I39125,I39128,I39144,I39154,I39164,I39174,I39184,I39194,I39204,I39214,I39224,I39264,I39267,I39270,I39273,I39276,I39279,I39282,I39285,I39288,I39291,I39307,I39317,I39327,I39337,I39347,I39357,I39367,I39377,I39387,I39397,I39437,I39440,I39443,I39446,I39449,I39452,I39455,I39458,I39461,I39477,I39487,I39497,I39507,I39517,I39527,I39537,I39547,I39557,I39597,I39600,I39603,I39606,I39609,I39612,I39615,I39618,I39621,I39624,I39640,I39650,I39660,I39670,I39680,I39690,I39700,I39710,I39720,I39730,I39770,I39773,I39776,I39779,I39782,I39785,I39788,I39791,I39794,I39810,I39820,I39830,I39840,I39850,I39860,I39870,I39880,I39890,I39930,I39933,I39936,I39939,I39942,I39945,I39948,I39951,I39954,I39970,I39980,I39990,I40000,I40010,I40020,I40030,I40040,I40050,I40090,I40093,I40096,I40099,I40102,I40105,I40108,I40111,I40114,I40117,I40133,I40143,I40153,I40163,I40173,I40183,I40193,I40203,I40213,I40223,I40263,I40266,I40269,I40272,I40275,I40278,I40281,I40284,I40287,I40290,I40306,I40316,I40326,I40336,I40346,I40356,I40366,I40376,I40386,I40396,I40436,I40439,I40442,I40445,I40448,I40451,I40454,I40457,I40460,I40476,I40486,I40496,I40506,I40516,I40526,I40536,I40546,I40556,I40596,I40599,I40602,I40605,I40608,I40611,I40614,I40617,I40620,I40636,I40646,I40656,I40666,I40676,I40686,I40696,I40706,I40716,I40756,I40759,I40762,I40765,I40768,I40771,I40774,I40777,I40780,I40796,I40806,I40816,I40826,I40836,I40846,I40856,I40866,I40876,I40916,I40919,I40922,I40925,I40928,I40931,I40934,I40937,I40940,I40943,I40959,I40969,I40979,I40989,I40999,I41009,I41019,I41029,I41039,I41049,I41089,I41092,I41095,I41098,I41101,I41104,I41107,I41110,I41113,I41116,I41132,I41142,I41152,I41162,I41172,I41182,I41192,I41202,I41212,I41222,I41262,I41265,I41268,I41271,I41274,I41277,I41280,I41283,I41286,I41289,I41305,I41315,I41325,I41335,I41345,I41355,I41365,I41375,I41385,I41395,I41435,I41438,I41441,I41444,I41447,I41450,I41453,I41456,I41472,I41482,I41492,I41502,I41512,I41522,I41532,I41542,I41582,I41585,I41588,I41591,I41594,I41597,I41600,I41603,I41606,I41609,I41625,I41635,I41645,I41655,I41665,I41675,I41685,I41695,I41705,I41715,I41755,I41758,I41761,I41764,I41767,I41770,I41773,I41776,I41779,I41795,I41805,I41815,I41825,I41835,I41845,I41855,I41865,I41875,I41915,I41918,I41921,I41924,I41927,I41930,I41933,I41936,I41939,I41955,I41965,I41975,I41985,I41995,I42005,I42015,I42025,I42035,I42075,I42078,I42081,I42084,I42087,I42090,I42093,I42096,I42099,I42205,I42215,I42225,I42235,I42245,I42255,I42265,I42275,I42285,I42295,I42305,I42345,I42348,I42351,I42354,I42357,I42360,I42363,I42366,I42369,I42372,I42388,I42398,I42408,I42418,I42428,I42438,I42448,I42458,I42468,I42478,I42518,I42521,I42524,I42527,I42530,I42533,I42536,I42539,I42542,I42558,I42568,I42578,I42588,I42598,I42608,I42618,I42628,I42638,I42678,I42681,I42684,I42687,I42690,I42693,I42696,I42699,I42702,I42718,I42728,I42738,I42748,I42758,I42768,I42778,I42788,I42798,I42838,I42841,I42844,I42847,I42850,I42853,I42856,I42859,I42862,I42878,I42888,I42898,I42908,I42918,I42928,I42938,I42948,I42958,I42998,I43001,I43004,I43007,I43010,I43013,I43016,I43019,I43022,I43025,I43041,I43051,I43061,I43071,I43081,I43091,I43101,I43111,I43121,I43131,I43171,I43174,I43177,I43180,I43183,I43186,I43189,I43192,I43208,I43218,I43228,I43238,I43248,I43258,I43268,I43278,I43318,I43321,I43324,I43327,I43330,I43333,I43336,I43339,I43342,I43358,I43368,I43378,I43388,I43398,I43408,I43418,I43428,I43438,I43478,I43481,I43484,I43487,I43490,I43493,I43496,I43499,I43502,I43518,I43528,I43538,I43548,I43558,I43568,I43578,I43588,I43598,I43638,I43641,I43644,I43647,I43650,I43653,I43656,I43659,I43662,I43665,I43681,I43691,I43701,I43711,I43721,I43731,I43741,I43751,I43761,I43771,I43811,I43814,I43817,I43820,I43823,I43826,I43829,I43832,I43835,I43851,I43861,I43871,I43881,I43891,I43901,I43911,I43921,I43931,I43971,I43974,I43977,I43980,I43983,I43986,I43989,I43992,I43995,I44011,I44021,I44031,I44041,I44051,I44061,I44071,I44081,I44091,I44131,I44134,I44137,I44140,I44143,I44146,I44149,I44152,I44155,I44158,I44174,I44184,I44194,I44204,I44214,I44224,I44234,I44244,I44254,I44264,I44304,I44307,I44310,I44313,I44316,I44319,I44322,I44325,I44328,I44331,I44347,I44357,I44367,I44377,I44387,I44397,I44407,I44417,I44427,I44437,I44477,I44480,I44483,I44486,I44489,I44492,I44495,I44498,I44501,I44517,I44527,I44537,I44547,I44557,I44567,I44577,I44587,I44597,I44637,I44640,I44643,I44646,I44649,I44652,I44655,I44658,I44661,I44677,I44687,I44697,I44707,I44717,I44727,I44737,I44747,I44757,I44797,I44800,I44803,I44806,I44809,I44812,I44815,I44818,I44821,I44837,I44847,I44857,I44867,I44877,I44887,I44897,I44907,I44917,I44957,I44960,I44963,I44966,I44969,I44972,I44975,I44978,I44981,I44997,I45007,I45017,I45027,I45037,I45047,I45057,I45067,I45077,I45117,I45120,I45123,I45126,I45129,I45132,I45135,I45138,I45141,I45157,I45167,I45177,I45187,I45197,I45207,I45217,I45227,I45237,I45277,I45280,I45283,I45286,I45289,I45292,I45295,I45298,I45301,I45317,I45327,I45337,I45347,I45357,I45367,I45377,I45387,I45397,I45437,I45440,I45443,I45446,I45449,I45452,I45455,I45458,I45461,I45477,I45487,I45497,I45507,I45517,I45527,I45537,I45547,I45557,I45597,I45600,I45603,I45606,I45609,I45612,I45615,I45618,I45621,I45624,I45640,I45650,I45660,I45670,I45680,I45690,I45700,I45710,I45720,I45730,I45770,I45773,I45776,I45779,I45782,I45785,I45788,I45791,I45794,I45810,I45820,I45830,I45840,I45850,I45860,I45870,I45880,I45890,I45930,I45933,I45936,I45939,I45942,I45945,I45948,I45951,I45967,I45977,I45987,I45997,I46007,I46017,I46027,I46037,I46077,I46080,I46083,I46086,I46089,I46092,I46095,I46098,I46101,I46117,I46127,I46137,I46147,I46157,I46167,I46177,I46187,I46197,I46237,I46240,I46243,I46246,I46249,I46252,I46255,I46258,I46261,I46264,I46280,I46290,I46300,I46310,I46320,I46330,I46340,I46350,I46360,I46370,I46410,I46413,I46416,I46419,I46422,I46425,I46428,I46431,I46434,I46450,I46460,I46470,I46480,I46490,I46500,I46510,I46520,I46530,I46570,I46573,I46576,I46579,I46582,I46585,I46588,I46591,I46594,I46597,I46613,I46623,I46633,I46643,I46653,I46663,I46673,I46683,I46693,I46703,I46743,I46746,I46749,I46752,I46755,I46758,I46761,I46764,I46767,I46783,I46793,I46803,I46813,I46823,I46833,I46843,I46853,I46863,I46903,I46906,I46909,I46912,I46915,I46918,I46921,I46924,I46927,I46943,I46953,I46963,I46973,I46983,I46993,I47003,I47013,I47023,I47063,I47066,I47069,I47072,I47075,I47078,I47081,I47084,I47100,I47110,I47120,I47130,I47140,I47150,I47160,I47170,I47210,I47213,I47216,I47219,I47222,I47225,I47228,I47231,I47234,I47250,I47260,I47270,I47280,I47290,I47300,I47310,I47320,I47330,I47370,I47373,I47376,I47379,I47382,I47385,I47388,I47391,I47407,I47417,I47427,I47437,I47447,I47457,I47467,I47477,I47517,I47520,I47523,I47526,I47529,I47532,I47535,I47538,I47541,I47544,I47560,I47570,I47580,I47590,I47600,I47610,I47620,I47630,I47640,I47650,I47690,I47693,I47696,I47699,I47702,I47705,I47708,I47711,I47727,I47737,I47747,I47757,I47767,I47777,I47787,I47797,I47837,I47840,I47843,I47846,I47849,I47852,I47855,I47858,I47861,I47877,I47887,I47897,I47907,I47917,I47927,I47937,I47947,I47957,I47997,I48000,I48003,I48006,I48009,I48012,I48015,I48018,I48021,I48037,I48047,I48057,I48067,I48077,I48087,I48097,I48107,I48117,I48157,I48160,I48163,I48166,I48169,I48172,I48175,I48178,I48181,I48184,I48200,I48210,I48220,I48230,I48240,I48250,I48260,I48270,I48280,I48290,I48330,I48333,I48336,I48339,I48342,I48345,I48348,I48351,I48354,I48357,I48373,I48383,I48393,I48403,I48413,I48423,I48433,I48443,I48453,I48463,I48503,I48506,I48509,I48512,I48515,I48518,I48521,I48524,I48527,I48543,I48553,I48563,I48573,I48583,I48593,I48603,I48613,I48623,I48663,I48666,I48669,I48672,I48675,I48678,I48681,I48684,I48700,I48710,I48720,I48730,I48740,I48750,I48760,I48770,I48810,I48813,I48816,I48819,I48822,I48825,I48828,I48831,I48834,I48837,I48853,I48863,I48873,I48883,I48893,I48903,I48913,I48923,I48933,I48943,I48983,I48986,I48989,I48992,I48995,I48998,I49001,I49004,I49007,I49023,I49033,I49043,I49053,I49063,I49073,I49083,I49093,I49103,I49143,I49146,I49149,I49152,I49155,I49158,I49161,I49164,I49180,I49190,I49200,I49210,I49220,I49230,I49240,I49250,I49290,I49293,I49296,I49299,I49302,I49305,I49308,I49311,I49314,I49317,I49333,I49343,I49353,I49363,I49373,I49383,I49393,I49403,I49413,I49423,I49463,I49466,I49469,I49472,I49475,I49478,I49481,I49484,I49487,I49503,I49513,I49523,I49533,I49543,I49553,I49563,I49573,I49583,I49623,I49626,I49629,I49632,I49635,I49638,I49641,I49644,I49647,I49663,I49673,I49683,I49693,I49703,I49713,I49723,I49733,I49743,I49783,I49786,I49789,I49792,I49795,I49798,I49801,I49804,I49807,I49810,I49826,I49836,I49846,I49856,I49866,I49876,I49886,I49896,I49906,I49916,I49956,I49959,I49962,I49965,I49968,I49971,I49974,I49977,I49980,I49983,I49999,I50009,I50019,I50029,I50039,I50049,I50059,I50069,I50079,I50089,I50129,I50132,I50135,I50138,I50141,I50144,I50147,I50150,I50153,I50156;
IN_INSTANCE I_0 (I1725,I1909);
IN_INSTANCE I_1 (I1437,I1919);
IN_INSTANCE I_2 (I1485,I1929);
IN_INSTANCE I_3 (I1765,I1939);
IN_INSTANCE I_4 (I1509,I1949);
IN_INSTANCE I_5 (I1605,I1959);
IN_INSTANCE I_6 (I1749,I1969);
IN_INSTANCE I_7 (I1653,I1979);
IN_INSTANCE I_8 (I1629,I1989);
IN_INSTANCE I_9 (I1533,I1999);
IN_INSTANCE I_10 (I1445,I2009);
PAT_11 I_11 (I1909,I1919,I1929,I1939,I1949,I1959,I1969,I1979,I1989,I1999,I2009,I2049,I2052,I2055,I2058,I2061,I2064,I2067,I2070,I2073,I2076,I1892,I1899);
OUT_INSTANCE I_12 (I2049,I2092);
OUT_INSTANCE I_13 (I2052,I2102);
OUT_INSTANCE I_14 (I2055,I2112);
OUT_INSTANCE I_15 (I2058,I2122);
OUT_INSTANCE I_16 (I2061,I2132);
OUT_INSTANCE I_17 (I2064,I2142);
OUT_INSTANCE I_18 (I2067,I2152);
OUT_INSTANCE I_19 (I2070,I2162);
OUT_INSTANCE I_20 (I2073,I2172);
OUT_INSTANCE I_21 (I2076,I2182);
PAT_13 I_22 (I2092,I2102,I2132,I2172,I2182,I2142,I2162,I2122,I2152,I2112,I2092,I2222,I2225,I2228,I2231,I2234,I2237,I2240,I2243,I2246,I1892,I1899);
OUT_INSTANCE I_23 (I2222,I2262);
OUT_INSTANCE I_24 (I2225,I2272);
OUT_INSTANCE I_25 (I2228,I2282);
OUT_INSTANCE I_26 (I2231,I2292);
OUT_INSTANCE I_27 (I2234,I2302);
OUT_INSTANCE I_28 (I2237,I2312);
OUT_INSTANCE I_29 (I2240,I2322);
OUT_INSTANCE I_30 (I2243,I2332);
OUT_INSTANCE I_31 (I2246,I2342);
PAT_15 I_32 (I2262,I2302,I2272,I2312,I2262,I2292,I2342,I2332,I2282,I2322,I2272,I2382,I2385,I2388,I2391,I2394,I2397,I2400,I2403,I2406,I1892,I1899);
OUT_INSTANCE I_33 (I2382,I2422);
OUT_INSTANCE I_34 (I2385,I2432);
OUT_INSTANCE I_35 (I2388,I2442);
OUT_INSTANCE I_36 (I2391,I2452);
OUT_INSTANCE I_37 (I2394,I2462);
OUT_INSTANCE I_38 (I2397,I2472);
OUT_INSTANCE I_39 (I2400,I2482);
OUT_INSTANCE I_40 (I2403,I2492);
OUT_INSTANCE I_41 (I2406,I2502);
PAT_6 I_42 (I2432,I2422,I2442,I2492,I2432,I2502,I2452,I2472,I2462,I2482,I2422,I2542,I2545,I2548,I2551,I2554,I2557,I2560,I2563,I2566,I2569,I1892,I1899);
OUT_INSTANCE I_43 (I2542,I2585);
OUT_INSTANCE I_44 (I2545,I2595);
OUT_INSTANCE I_45 (I2548,I2605);
OUT_INSTANCE I_46 (I2551,I2615);
OUT_INSTANCE I_47 (I2554,I2625);
OUT_INSTANCE I_48 (I2557,I2635);
OUT_INSTANCE I_49 (I2560,I2645);
OUT_INSTANCE I_50 (I2563,I2655);
OUT_INSTANCE I_51 (I2566,I2665);
OUT_INSTANCE I_52 (I2569,I2675);
PAT_13 I_53 (I2665,I2605,I2655,I2585,I2595,I2615,I2675,I2625,I2645,I2585,I2635,I2715,I2718,I2721,I2724,I2727,I2730,I2733,I2736,I2739,I1892,I1899);
OUT_INSTANCE I_54 (I2715,I2755);
OUT_INSTANCE I_55 (I2718,I2765);
OUT_INSTANCE I_56 (I2721,I2775);
OUT_INSTANCE I_57 (I2724,I2785);
OUT_INSTANCE I_58 (I2727,I2795);
OUT_INSTANCE I_59 (I2730,I2805);
OUT_INSTANCE I_60 (I2733,I2815);
OUT_INSTANCE I_61 (I2736,I2825);
OUT_INSTANCE I_62 (I2739,I2835);
PAT_17 I_63 (I2835,I2795,I2825,I2815,I2785,I2755,I2765,I2775,I2755,I2805,I2765,I2875,I2878,I2881,I2884,I2887,I2890,I2893,I2896,I2899,I2902,I1892,I1899);
OUT_INSTANCE I_64 (I2875,I2918);
OUT_INSTANCE I_65 (I2878,I2928);
OUT_INSTANCE I_66 (I2881,I2938);
OUT_INSTANCE I_67 (I2884,I2948);
OUT_INSTANCE I_68 (I2887,I2958);
OUT_INSTANCE I_69 (I2890,I2968);
OUT_INSTANCE I_70 (I2893,I2978);
OUT_INSTANCE I_71 (I2896,I2988);
OUT_INSTANCE I_72 (I2899,I2998);
OUT_INSTANCE I_73 (I2902,I3008);
PAT_14 I_74 (I2928,I2978,I2918,I2998,I2948,I2968,I2918,I2988,I2938,I3008,I2958,I3048,I3051,I3054,I3057,I3060,I3063,I3066,I3069,I3072,I1892,I1899);
OUT_INSTANCE I_75 (I3048,I3088);
OUT_INSTANCE I_76 (I3051,I3098);
OUT_INSTANCE I_77 (I3054,I3108);
OUT_INSTANCE I_78 (I3057,I3118);
OUT_INSTANCE I_79 (I3060,I3128);
OUT_INSTANCE I_80 (I3063,I3138);
OUT_INSTANCE I_81 (I3066,I3148);
OUT_INSTANCE I_82 (I3069,I3158);
OUT_INSTANCE I_83 (I3072,I3168);
PAT_13 I_84 (I3118,I3168,I3098,I3128,I3088,I3098,I3148,I3108,I3088,I3158,I3138,I3208,I3211,I3214,I3217,I3220,I3223,I3226,I3229,I3232,I1892,I1899);
OUT_INSTANCE I_85 (I3208,I3248);
OUT_INSTANCE I_86 (I3211,I3258);
OUT_INSTANCE I_87 (I3214,I3268);
OUT_INSTANCE I_88 (I3217,I3278);
OUT_INSTANCE I_89 (I3220,I3288);
OUT_INSTANCE I_90 (I3223,I3298);
OUT_INSTANCE I_91 (I3226,I3308);
OUT_INSTANCE I_92 (I3229,I3318);
OUT_INSTANCE I_93 (I3232,I3328);
PAT_11 I_94 (I3248,I3288,I3298,I3268,I3258,I3328,I3258,I3318,I3278,I3248,I3308,I3368,I3371,I3374,I3377,I3380,I3383,I3386,I3389,I3392,I3395,I1892,I1899);
OUT_INSTANCE I_95 (I3368,I3411);
OUT_INSTANCE I_96 (I3371,I3421);
OUT_INSTANCE I_97 (I3374,I3431);
OUT_INSTANCE I_98 (I3377,I3441);
OUT_INSTANCE I_99 (I3380,I3451);
OUT_INSTANCE I_100 (I3383,I3461);
OUT_INSTANCE I_101 (I3386,I3471);
OUT_INSTANCE I_102 (I3389,I3481);
OUT_INSTANCE I_103 (I3392,I3491);
OUT_INSTANCE I_104 (I3395,I3501);
PAT_9 I_105 (I3431,I3471,I3441,I3481,I3411,I3421,I3451,I3411,I3461,I3491,I3501,I3541,I3544,I3547,I3550,I3553,I3556,I3559,I3562,I3565,I1892,I1899);
OUT_INSTANCE I_106 (I3541,I3581);
OUT_INSTANCE I_107 (I3544,I3591);
OUT_INSTANCE I_108 (I3547,I3601);
OUT_INSTANCE I_109 (I3550,I3611);
OUT_INSTANCE I_110 (I3553,I3621);
OUT_INSTANCE I_111 (I3556,I3631);
OUT_INSTANCE I_112 (I3559,I3641);
OUT_INSTANCE I_113 (I3562,I3651);
OUT_INSTANCE I_114 (I3565,I3661);
PAT_11 I_115 (I3621,I3641,I3661,I3651,I3611,I3591,I3591,I3581,I3631,I3581,I3601,I3701,I3704,I3707,I3710,I3713,I3716,I3719,I3722,I3725,I3728,I1892,I1899);
OUT_INSTANCE I_116 (I3701,I3744);
OUT_INSTANCE I_117 (I3704,I3754);
OUT_INSTANCE I_118 (I3707,I3764);
OUT_INSTANCE I_119 (I3710,I3774);
OUT_INSTANCE I_120 (I3713,I3784);
OUT_INSTANCE I_121 (I3716,I3794);
OUT_INSTANCE I_122 (I3719,I3804);
OUT_INSTANCE I_123 (I3722,I3814);
OUT_INSTANCE I_124 (I3725,I3824);
OUT_INSTANCE I_125 (I3728,I3834);
PAT_10 I_126 (I3794,I3814,I3784,I3764,I3824,I3774,I3834,I3804,I3744,I3754,I3744,I3874,I3877,I3880,I3883,I3886,I3889,I3892,I3895,I1892,I1899);
OUT_INSTANCE I_127 (I3874,I3911);
OUT_INSTANCE I_128 (I3877,I3921);
OUT_INSTANCE I_129 (I3880,I3931);
OUT_INSTANCE I_130 (I3883,I3941);
OUT_INSTANCE I_131 (I3886,I3951);
OUT_INSTANCE I_132 (I3889,I3961);
OUT_INSTANCE I_133 (I3892,I3971);
OUT_INSTANCE I_134 (I3895,I3981);
PAT_14 I_135 (I3911,I3981,I3931,I3961,I3951,I3971,I3941,I3921,I3921,I3931,I3911,I4021,I4024,I4027,I4030,I4033,I4036,I4039,I4042,I4045,I1892,I1899);
OUT_INSTANCE I_136 (I4021,I4061);
OUT_INSTANCE I_137 (I4024,I4071);
OUT_INSTANCE I_138 (I4027,I4081);
OUT_INSTANCE I_139 (I4030,I4091);
OUT_INSTANCE I_140 (I4033,I4101);
OUT_INSTANCE I_141 (I4036,I4111);
OUT_INSTANCE I_142 (I4039,I4121);
OUT_INSTANCE I_143 (I4042,I4131);
OUT_INSTANCE I_144 (I4045,I4141);
PAT_11 I_145 (I4101,I4091,I4081,I4061,I4071,I4071,I4111,I4061,I4131,I4141,I4121,I4181,I4184,I4187,I4190,I4193,I4196,I4199,I4202,I4205,I4208,I1892,I1899);
OUT_INSTANCE I_146 (I4181,I4224);
OUT_INSTANCE I_147 (I4184,I4234);
OUT_INSTANCE I_148 (I4187,I4244);
OUT_INSTANCE I_149 (I4190,I4254);
OUT_INSTANCE I_150 (I4193,I4264);
OUT_INSTANCE I_151 (I4196,I4274);
OUT_INSTANCE I_152 (I4199,I4284);
OUT_INSTANCE I_153 (I4202,I4294);
OUT_INSTANCE I_154 (I4205,I4304);
OUT_INSTANCE I_155 (I4208,I4314);
PAT_6 I_156 (I4224,I4314,I4274,I4304,I4284,I4264,I4234,I4294,I4254,I4244,I4224,I4354,I4357,I4360,I4363,I4366,I4369,I4372,I4375,I4378,I4381,I1892,I1899);
OUT_INSTANCE I_157 (I4354,I4397);
OUT_INSTANCE I_158 (I4357,I4407);
OUT_INSTANCE I_159 (I4360,I4417);
OUT_INSTANCE I_160 (I4363,I4427);
OUT_INSTANCE I_161 (I4366,I4437);
OUT_INSTANCE I_162 (I4369,I4447);
OUT_INSTANCE I_163 (I4372,I4457);
OUT_INSTANCE I_164 (I4375,I4467);
OUT_INSTANCE I_165 (I4378,I4477);
OUT_INSTANCE I_166 (I4381,I4487);
PAT_10 I_167 (I4397,I4447,I4457,I4427,I4397,I4477,I4487,I4407,I4437,I4417,I4467,I4527,I4530,I4533,I4536,I4539,I4542,I4545,I4548,I1892,I1899);
OUT_INSTANCE I_168 (I4527,I4564);
OUT_INSTANCE I_169 (I4530,I4574);
OUT_INSTANCE I_170 (I4533,I4584);
OUT_INSTANCE I_171 (I4536,I4594);
OUT_INSTANCE I_172 (I4539,I4604);
OUT_INSTANCE I_173 (I4542,I4614);
OUT_INSTANCE I_174 (I4545,I4624);
OUT_INSTANCE I_175 (I4548,I4634);
PAT_9 I_176 (I4604,I4564,I4574,I4584,I4564,I4584,I4594,I4574,I4634,I4614,I4624,I4674,I4677,I4680,I4683,I4686,I4689,I4692,I4695,I4698,I1892,I1899);
OUT_INSTANCE I_177 (I4674,I4714);
OUT_INSTANCE I_178 (I4677,I4724);
OUT_INSTANCE I_179 (I4680,I4734);
OUT_INSTANCE I_180 (I4683,I4744);
OUT_INSTANCE I_181 (I4686,I4754);
OUT_INSTANCE I_182 (I4689,I4764);
OUT_INSTANCE I_183 (I4692,I4774);
OUT_INSTANCE I_184 (I4695,I4784);
OUT_INSTANCE I_185 (I4698,I4794);
PAT_2 I_186 (I4764,I4774,I4744,I4794,I4714,I4724,I4734,I4724,I4784,I4754,I4714,I4834,I4837,I4840,I4843,I4846,I4849,I4852,I4855,I4858,I1892,I1899);
OUT_INSTANCE I_187 (I4834,I4874);
OUT_INSTANCE I_188 (I4837,I4884);
OUT_INSTANCE I_189 (I4840,I4894);
OUT_INSTANCE I_190 (I4843,I4904);
OUT_INSTANCE I_191 (I4846,I4914);
OUT_INSTANCE I_192 (I4849,I4924);
OUT_INSTANCE I_193 (I4852,I4934);
OUT_INSTANCE I_194 (I4855,I4944);
OUT_INSTANCE I_195 (I4858,I4954);
PAT_8 I_196 (I4914,I4884,I4904,I4874,I4894,I4944,I4934,I4874,I4924,I4884,I4954,I4994,I4997,I5000,I5003,I5006,I5009,I5012,I5015,I5018,I1892,I1899);
OUT_INSTANCE I_197 (I4994,I5034);
OUT_INSTANCE I_198 (I4997,I5044);
OUT_INSTANCE I_199 (I5000,I5054);
OUT_INSTANCE I_200 (I5003,I5064);
OUT_INSTANCE I_201 (I5006,I5074);
OUT_INSTANCE I_202 (I5009,I5084);
OUT_INSTANCE I_203 (I5012,I5094);
OUT_INSTANCE I_204 (I5015,I5104);
OUT_INSTANCE I_205 (I5018,I5114);
PAT_2 I_206 (I5044,I5094,I5114,I5034,I5074,I5084,I5044,I5104,I5054,I5064,I5034,I5154,I5157,I5160,I5163,I5166,I5169,I5172,I5175,I5178,I1892,I1899);
OUT_INSTANCE I_207 (I5154,I5194);
OUT_INSTANCE I_208 (I5157,I5204);
OUT_INSTANCE I_209 (I5160,I5214);
OUT_INSTANCE I_210 (I5163,I5224);
OUT_INSTANCE I_211 (I5166,I5234);
OUT_INSTANCE I_212 (I5169,I5244);
OUT_INSTANCE I_213 (I5172,I5254);
OUT_INSTANCE I_214 (I5175,I5264);
OUT_INSTANCE I_215 (I5178,I5274);
PAT_13 I_216 (I5224,I5204,I5194,I5264,I5234,I5244,I5204,I5214,I5254,I5274,I5194,I5314,I5317,I5320,I5323,I5326,I5329,I5332,I5335,I5338,I1892,I1899);
OUT_INSTANCE I_217 (I5314,I5354);
OUT_INSTANCE I_218 (I5317,I5364);
OUT_INSTANCE I_219 (I5320,I5374);
OUT_INSTANCE I_220 (I5323,I5384);
OUT_INSTANCE I_221 (I5326,I5394);
OUT_INSTANCE I_222 (I5329,I5404);
OUT_INSTANCE I_223 (I5332,I5414);
OUT_INSTANCE I_224 (I5335,I5424);
OUT_INSTANCE I_225 (I5338,I5434);
PAT_9 I_226 (I5424,I5364,I5364,I5354,I5434,I5374,I5384,I5354,I5394,I5414,I5404,I5474,I5477,I5480,I5483,I5486,I5489,I5492,I5495,I5498,I1892,I1899);
OUT_INSTANCE I_227 (I5474,I5514);
OUT_INSTANCE I_228 (I5477,I5524);
OUT_INSTANCE I_229 (I5480,I5534);
OUT_INSTANCE I_230 (I5483,I5544);
OUT_INSTANCE I_231 (I5486,I5554);
OUT_INSTANCE I_232 (I5489,I5564);
OUT_INSTANCE I_233 (I5492,I5574);
OUT_INSTANCE I_234 (I5495,I5584);
OUT_INSTANCE I_235 (I5498,I5594);
PAT_6 I_236 (I5574,I5514,I5554,I5584,I5514,I5544,I5534,I5594,I5564,I5524,I5524,I5634,I5637,I5640,I5643,I5646,I5649,I5652,I5655,I5658,I5661,I1892,I1899);
OUT_INSTANCE I_237 (I5634,I5677);
OUT_INSTANCE I_238 (I5637,I5687);
OUT_INSTANCE I_239 (I5640,I5697);
OUT_INSTANCE I_240 (I5643,I5707);
OUT_INSTANCE I_241 (I5646,I5717);
OUT_INSTANCE I_242 (I5649,I5727);
OUT_INSTANCE I_243 (I5652,I5737);
OUT_INSTANCE I_244 (I5655,I5747);
OUT_INSTANCE I_245 (I5658,I5757);
OUT_INSTANCE I_246 (I5661,I5767);
PAT_2 I_247 (I5747,I5767,I5707,I5727,I5677,I5697,I5677,I5717,I5687,I5737,I5757,I5807,I5810,I5813,I5816,I5819,I5822,I5825,I5828,I5831,I1892,I1899);
OUT_INSTANCE I_248 (I5807,I5847);
OUT_INSTANCE I_249 (I5810,I5857);
OUT_INSTANCE I_250 (I5813,I5867);
OUT_INSTANCE I_251 (I5816,I5877);
OUT_INSTANCE I_252 (I5819,I5887);
OUT_INSTANCE I_253 (I5822,I5897);
OUT_INSTANCE I_254 (I5825,I5907);
OUT_INSTANCE I_255 (I5828,I5917);
OUT_INSTANCE I_256 (I5831,I5927);
PAT_8 I_257 (I5887,I5857,I5877,I5847,I5867,I5917,I5907,I5847,I5897,I5857,I5927,I5967,I5970,I5973,I5976,I5979,I5982,I5985,I5988,I5991,I1892,I1899);
OUT_INSTANCE I_258 (I5967,I6007);
OUT_INSTANCE I_259 (I5970,I6017);
OUT_INSTANCE I_260 (I5973,I6027);
OUT_INSTANCE I_261 (I5976,I6037);
OUT_INSTANCE I_262 (I5979,I6047);
OUT_INSTANCE I_263 (I5982,I6057);
OUT_INSTANCE I_264 (I5985,I6067);
OUT_INSTANCE I_265 (I5988,I6077);
OUT_INSTANCE I_266 (I5991,I6087);
PAT_2 I_267 (I6017,I6067,I6087,I6007,I6047,I6057,I6017,I6077,I6027,I6037,I6007,I6127,I6130,I6133,I6136,I6139,I6142,I6145,I6148,I6151,I1892,I1899);
OUT_INSTANCE I_268 (I6127,I6167);
OUT_INSTANCE I_269 (I6130,I6177);
OUT_INSTANCE I_270 (I6133,I6187);
OUT_INSTANCE I_271 (I6136,I6197);
OUT_INSTANCE I_272 (I6139,I6207);
OUT_INSTANCE I_273 (I6142,I6217);
OUT_INSTANCE I_274 (I6145,I6227);
OUT_INSTANCE I_275 (I6148,I6237);
OUT_INSTANCE I_276 (I6151,I6247);
PAT_9 I_277 (I6217,I6247,I6167,I6187,I6197,I6227,I6177,I6207,I6237,I6177,I6167,I6287,I6290,I6293,I6296,I6299,I6302,I6305,I6308,I6311,I1892,I1899);
OUT_INSTANCE I_278 (I6287,I6327);
OUT_INSTANCE I_279 (I6290,I6337);
OUT_INSTANCE I_280 (I6293,I6347);
OUT_INSTANCE I_281 (I6296,I6357);
OUT_INSTANCE I_282 (I6299,I6367);
OUT_INSTANCE I_283 (I6302,I6377);
OUT_INSTANCE I_284 (I6305,I6387);
OUT_INSTANCE I_285 (I6308,I6397);
OUT_INSTANCE I_286 (I6311,I6407);
PAT_15 I_287 (I6367,I6397,I6407,I6337,I6387,I6347,I6357,I6327,I6377,I6327,I6337,I6447,I6450,I6453,I6456,I6459,I6462,I6465,I6468,I6471,I1892,I1899);
OUT_INSTANCE I_288 (I6447,I6487);
OUT_INSTANCE I_289 (I6450,I6497);
OUT_INSTANCE I_290 (I6453,I6507);
OUT_INSTANCE I_291 (I6456,I6517);
OUT_INSTANCE I_292 (I6459,I6527);
OUT_INSTANCE I_293 (I6462,I6537);
OUT_INSTANCE I_294 (I6465,I6547);
OUT_INSTANCE I_295 (I6468,I6557);
OUT_INSTANCE I_296 (I6471,I6567);
PAT_16 I_297 (I6497,I6507,I6557,I6497,I6567,I6487,I6537,I6487,I6547,I6517,I6527,I6607,I6610,I6613,I6616,I6619,I6622,I6625,I6628,I6631,I6634,I1892,I1899);
OUT_INSTANCE I_298 (I6607,I6650);
OUT_INSTANCE I_299 (I6610,I6660);
OUT_INSTANCE I_300 (I6613,I6670);
OUT_INSTANCE I_301 (I6616,I6680);
OUT_INSTANCE I_302 (I6619,I6690);
OUT_INSTANCE I_303 (I6622,I6700);
OUT_INSTANCE I_304 (I6625,I6710);
OUT_INSTANCE I_305 (I6628,I6720);
OUT_INSTANCE I_306 (I6631,I6730);
OUT_INSTANCE I_307 (I6634,I6740);
PAT_11 I_308 (I6660,I6650,I6740,I6670,I6720,I6730,I6710,I6650,I6680,I6690,I6700,I6780,I6783,I6786,I6789,I6792,I6795,I6798,I6801,I6804,I6807,I1892,I1899);
OUT_INSTANCE I_309 (I6780,I6823);
OUT_INSTANCE I_310 (I6783,I6833);
OUT_INSTANCE I_311 (I6786,I6843);
OUT_INSTANCE I_312 (I6789,I6853);
OUT_INSTANCE I_313 (I6792,I6863);
OUT_INSTANCE I_314 (I6795,I6873);
OUT_INSTANCE I_315 (I6798,I6883);
OUT_INSTANCE I_316 (I6801,I6893);
OUT_INSTANCE I_317 (I6804,I6903);
OUT_INSTANCE I_318 (I6807,I6913);
PAT_13 I_319 (I6823,I6833,I6863,I6903,I6913,I6873,I6893,I6853,I6883,I6843,I6823,I6953,I6956,I6959,I6962,I6965,I6968,I6971,I6974,I6977,I1892,I1899);
OUT_INSTANCE I_320 (I6953,I6993);
OUT_INSTANCE I_321 (I6956,I7003);
OUT_INSTANCE I_322 (I6959,I7013);
OUT_INSTANCE I_323 (I6962,I7023);
OUT_INSTANCE I_324 (I6965,I7033);
OUT_INSTANCE I_325 (I6968,I7043);
OUT_INSTANCE I_326 (I6971,I7053);
OUT_INSTANCE I_327 (I6974,I7063);
OUT_INSTANCE I_328 (I6977,I7073);
PAT_5 I_329 (I7033,I7003,I7023,I7063,I7003,I7073,I7013,I7043,I6993,I6993,I7053,I7113,I7116,I7119,I7122,I7125,I7128,I7131,I7134,I7137,I7140,I1892,I1899);
OUT_INSTANCE I_330 (I7113,I7156);
OUT_INSTANCE I_331 (I7116,I7166);
OUT_INSTANCE I_332 (I7119,I7176);
OUT_INSTANCE I_333 (I7122,I7186);
OUT_INSTANCE I_334 (I7125,I7196);
OUT_INSTANCE I_335 (I7128,I7206);
OUT_INSTANCE I_336 (I7131,I7216);
OUT_INSTANCE I_337 (I7134,I7226);
OUT_INSTANCE I_338 (I7137,I7236);
OUT_INSTANCE I_339 (I7140,I7246);
PAT_11 I_340 (I7196,I7186,I7166,I7226,I7236,I7156,I7216,I7206,I7246,I7176,I7156,I7286,I7289,I7292,I7295,I7298,I7301,I7304,I7307,I7310,I7313,I1892,I1899);
OUT_INSTANCE I_341 (I7286,I7329);
OUT_INSTANCE I_342 (I7289,I7339);
OUT_INSTANCE I_343 (I7292,I7349);
OUT_INSTANCE I_344 (I7295,I7359);
OUT_INSTANCE I_345 (I7298,I7369);
OUT_INSTANCE I_346 (I7301,I7379);
OUT_INSTANCE I_347 (I7304,I7389);
OUT_INSTANCE I_348 (I7307,I7399);
OUT_INSTANCE I_349 (I7310,I7409);
OUT_INSTANCE I_350 (I7313,I7419);
PAT_17 I_351 (I7369,I7339,I7419,I7329,I7359,I7399,I7389,I7379,I7329,I7409,I7349,I7459,I7462,I7465,I7468,I7471,I7474,I7477,I7480,I7483,I7486,I1892,I1899);
OUT_INSTANCE I_352 (I7459,I7502);
OUT_INSTANCE I_353 (I7462,I7512);
OUT_INSTANCE I_354 (I7465,I7522);
OUT_INSTANCE I_355 (I7468,I7532);
OUT_INSTANCE I_356 (I7471,I7542);
OUT_INSTANCE I_357 (I7474,I7552);
OUT_INSTANCE I_358 (I7477,I7562);
OUT_INSTANCE I_359 (I7480,I7572);
OUT_INSTANCE I_360 (I7483,I7582);
OUT_INSTANCE I_361 (I7486,I7592);
PAT_9 I_362 (I7572,I7512,I7532,I7582,I7522,I7562,I7502,I7542,I7502,I7592,I7552,I7632,I7635,I7638,I7641,I7644,I7647,I7650,I7653,I7656,I1892,I1899);
OUT_INSTANCE I_363 (I7632,I7672);
OUT_INSTANCE I_364 (I7635,I7682);
OUT_INSTANCE I_365 (I7638,I7692);
OUT_INSTANCE I_366 (I7641,I7702);
OUT_INSTANCE I_367 (I7644,I7712);
OUT_INSTANCE I_368 (I7647,I7722);
OUT_INSTANCE I_369 (I7650,I7732);
OUT_INSTANCE I_370 (I7653,I7742);
OUT_INSTANCE I_371 (I7656,I7752);
PAT_13 I_372 (I7672,I7742,I7682,I7732,I7712,I7702,I7752,I7672,I7692,I7722,I7682,I7792,I7795,I7798,I7801,I7804,I7807,I7810,I7813,I7816,I1892,I1899);
OUT_INSTANCE I_373 (I7792,I7832);
OUT_INSTANCE I_374 (I7795,I7842);
OUT_INSTANCE I_375 (I7798,I7852);
OUT_INSTANCE I_376 (I7801,I7862);
OUT_INSTANCE I_377 (I7804,I7872);
OUT_INSTANCE I_378 (I7807,I7882);
OUT_INSTANCE I_379 (I7810,I7892);
OUT_INSTANCE I_380 (I7813,I7902);
OUT_INSTANCE I_381 (I7816,I7912);
PAT_4 I_382 (I7862,I7872,I7912,I7852,I7902,I7892,I7842,I7882,I7842,I7832,I7832,I7952,I7955,I7958,I7961,I7964,I7967,I7970,I7973,I7976,I1892,I1899);
OUT_INSTANCE I_383 (I7952,I7992);
OUT_INSTANCE I_384 (I7955,I8002);
OUT_INSTANCE I_385 (I7958,I8012);
OUT_INSTANCE I_386 (I7961,I8022);
OUT_INSTANCE I_387 (I7964,I8032);
OUT_INSTANCE I_388 (I7967,I8042);
OUT_INSTANCE I_389 (I7970,I8052);
OUT_INSTANCE I_390 (I7973,I8062);
OUT_INSTANCE I_391 (I7976,I8072);
PAT_9 I_392 (I8062,I8002,I8012,I8042,I8052,I7992,I8022,I8002,I8072,I7992,I8032,I8112,I8115,I8118,I8121,I8124,I8127,I8130,I8133,I8136,I1892,I1899);
OUT_INSTANCE I_393 (I8112,I8152);
OUT_INSTANCE I_394 (I8115,I8162);
OUT_INSTANCE I_395 (I8118,I8172);
OUT_INSTANCE I_396 (I8121,I8182);
OUT_INSTANCE I_397 (I8124,I8192);
OUT_INSTANCE I_398 (I8127,I8202);
OUT_INSTANCE I_399 (I8130,I8212);
OUT_INSTANCE I_400 (I8133,I8222);
OUT_INSTANCE I_401 (I8136,I8232);
PAT_5 I_402 (I8222,I8152,I8202,I8152,I8172,I8182,I8162,I8162,I8212,I8192,I8232,I8272,I8275,I8278,I8281,I8284,I8287,I8290,I8293,I8296,I8299,I1892,I1899);
OUT_INSTANCE I_403 (I8272,I8315);
OUT_INSTANCE I_404 (I8275,I8325);
OUT_INSTANCE I_405 (I8278,I8335);
OUT_INSTANCE I_406 (I8281,I8345);
OUT_INSTANCE I_407 (I8284,I8355);
OUT_INSTANCE I_408 (I8287,I8365);
OUT_INSTANCE I_409 (I8290,I8375);
OUT_INSTANCE I_410 (I8293,I8385);
OUT_INSTANCE I_411 (I8296,I8395);
OUT_INSTANCE I_412 (I8299,I8405);
PAT_1 I_413 (I8365,I8325,I8385,I8315,I8335,I8315,I8345,I8395,I8375,I8405,I8355,I8445,I8448,I8451,I8454,I8457,I8460,I8463,I8466,I8469,I1892,I1899);
OUT_INSTANCE I_414 (I8445,I8485);
OUT_INSTANCE I_415 (I8448,I8495);
OUT_INSTANCE I_416 (I8451,I8505);
OUT_INSTANCE I_417 (I8454,I8515);
OUT_INSTANCE I_418 (I8457,I8525);
OUT_INSTANCE I_419 (I8460,I8535);
OUT_INSTANCE I_420 (I8463,I8545);
OUT_INSTANCE I_421 (I8466,I8555);
OUT_INSTANCE I_422 (I8469,I8565);
PAT_13 I_423 (I8515,I8545,I8565,I8485,I8535,I8525,I8555,I8505,I8495,I8485,I8495,I8605,I8608,I8611,I8614,I8617,I8620,I8623,I8626,I8629,I1892,I1899);
OUT_INSTANCE I_424 (I8605,I8645);
OUT_INSTANCE I_425 (I8608,I8655);
OUT_INSTANCE I_426 (I8611,I8665);
OUT_INSTANCE I_427 (I8614,I8675);
OUT_INSTANCE I_428 (I8617,I8685);
OUT_INSTANCE I_429 (I8620,I8695);
OUT_INSTANCE I_430 (I8623,I8705);
OUT_INSTANCE I_431 (I8626,I8715);
OUT_INSTANCE I_432 (I8629,I8725);
PAT_8 I_433 (I8675,I8715,I8685,I8695,I8725,I8655,I8705,I8645,I8655,I8665,I8645,I8765,I8768,I8771,I8774,I8777,I8780,I8783,I8786,I8789,I1892,I1899);
OUT_INSTANCE I_434 (I8765,I8805);
OUT_INSTANCE I_435 (I8768,I8815);
OUT_INSTANCE I_436 (I8771,I8825);
OUT_INSTANCE I_437 (I8774,I8835);
OUT_INSTANCE I_438 (I8777,I8845);
OUT_INSTANCE I_439 (I8780,I8855);
OUT_INSTANCE I_440 (I8783,I8865);
OUT_INSTANCE I_441 (I8786,I8875);
OUT_INSTANCE I_442 (I8789,I8885);
PAT_13 I_443 (I8845,I8875,I8815,I8885,I8825,I8805,I8805,I8835,I8865,I8855,I8815,I8925,I8928,I8931,I8934,I8937,I8940,I8943,I8946,I8949,I1892,I1899);
OUT_INSTANCE I_444 (I8925,I8965);
OUT_INSTANCE I_445 (I8928,I8975);
OUT_INSTANCE I_446 (I8931,I8985);
OUT_INSTANCE I_447 (I8934,I8995);
OUT_INSTANCE I_448 (I8937,I9005);
OUT_INSTANCE I_449 (I8940,I9015);
OUT_INSTANCE I_450 (I8943,I9025);
OUT_INSTANCE I_451 (I8946,I9035);
OUT_INSTANCE I_452 (I8949,I9045);
PAT_7 I_453 (I8995,I9005,I8965,I9015,I9035,I8985,I8975,I9045,I8975,I8965,I9025,I9085,I9088,I9091,I9094,I9097,I9100,I9103,I9106,I9109,I1892,I1899);
OUT_INSTANCE I_454 (I9085,I9125);
OUT_INSTANCE I_455 (I9088,I9135);
OUT_INSTANCE I_456 (I9091,I9145);
OUT_INSTANCE I_457 (I9094,I9155);
OUT_INSTANCE I_458 (I9097,I9165);
OUT_INSTANCE I_459 (I9100,I9175);
OUT_INSTANCE I_460 (I9103,I9185);
OUT_INSTANCE I_461 (I9106,I9195);
OUT_INSTANCE I_462 (I9109,I9205);
PAT_4 I_463 (I9205,I9125,I9125,I9175,I9155,I9135,I9135,I9185,I9195,I9145,I9165,I9245,I9248,I9251,I9254,I9257,I9260,I9263,I9266,I9269,I1892,I1899);
OUT_INSTANCE I_464 (I9245,I9285);
OUT_INSTANCE I_465 (I9248,I9295);
OUT_INSTANCE I_466 (I9251,I9305);
OUT_INSTANCE I_467 (I9254,I9315);
OUT_INSTANCE I_468 (I9257,I9325);
OUT_INSTANCE I_469 (I9260,I9335);
OUT_INSTANCE I_470 (I9263,I9345);
OUT_INSTANCE I_471 (I9266,I9355);
OUT_INSTANCE I_472 (I9269,I9365);
PAT_17 I_473 (I9325,I9315,I9355,I9335,I9285,I9345,I9365,I9295,I9305,I9295,I9285,I9405,I9408,I9411,I9414,I9417,I9420,I9423,I9426,I9429,I9432,I1892,I1899);
OUT_INSTANCE I_474 (I9405,I9448);
OUT_INSTANCE I_475 (I9408,I9458);
OUT_INSTANCE I_476 (I9411,I9468);
OUT_INSTANCE I_477 (I9414,I9478);
OUT_INSTANCE I_478 (I9417,I9488);
OUT_INSTANCE I_479 (I9420,I9498);
OUT_INSTANCE I_480 (I9423,I9508);
OUT_INSTANCE I_481 (I9426,I9518);
OUT_INSTANCE I_482 (I9429,I9528);
OUT_INSTANCE I_483 (I9432,I9538);
PAT_8 I_484 (I9478,I9518,I9538,I9508,I9458,I9488,I9498,I9528,I9468,I9448,I9448,I9578,I9581,I9584,I9587,I9590,I9593,I9596,I9599,I9602,I1892,I1899);
OUT_INSTANCE I_485 (I9578,I9618);
OUT_INSTANCE I_486 (I9581,I9628);
OUT_INSTANCE I_487 (I9584,I9638);
OUT_INSTANCE I_488 (I9587,I9648);
OUT_INSTANCE I_489 (I9590,I9658);
OUT_INSTANCE I_490 (I9593,I9668);
OUT_INSTANCE I_491 (I9596,I9678);
OUT_INSTANCE I_492 (I9599,I9688);
OUT_INSTANCE I_493 (I9602,I9698);
PAT_2 I_494 (I9628,I9678,I9698,I9618,I9658,I9668,I9628,I9688,I9638,I9648,I9618,I9738,I9741,I9744,I9747,I9750,I9753,I9756,I9759,I9762,I1892,I1899);
OUT_INSTANCE I_495 (I9738,I9778);
OUT_INSTANCE I_496 (I9741,I9788);
OUT_INSTANCE I_497 (I9744,I9798);
OUT_INSTANCE I_498 (I9747,I9808);
OUT_INSTANCE I_499 (I9750,I9818);
OUT_INSTANCE I_500 (I9753,I9828);
OUT_INSTANCE I_501 (I9756,I9838);
OUT_INSTANCE I_502 (I9759,I9848);
OUT_INSTANCE I_503 (I9762,I9858);
PAT_5 I_504 (I9848,I9778,I9778,I9818,I9808,I9838,I9798,I9828,I9858,I9788,I9788,I9898,I9901,I9904,I9907,I9910,I9913,I9916,I9919,I9922,I9925,I1892,I1899);
OUT_INSTANCE I_505 (I9898,I9941);
OUT_INSTANCE I_506 (I9901,I9951);
OUT_INSTANCE I_507 (I9904,I9961);
OUT_INSTANCE I_508 (I9907,I9971);
OUT_INSTANCE I_509 (I9910,I9981);
OUT_INSTANCE I_510 (I9913,I9991);
OUT_INSTANCE I_511 (I9916,I10001);
OUT_INSTANCE I_512 (I9919,I10011);
OUT_INSTANCE I_513 (I9922,I10021);
OUT_INSTANCE I_514 (I9925,I10031);
IN_INSTANCE I_515 (I1597,I10041);
IN_INSTANCE I_516 (I1389,I10051);
IN_INSTANCE I_517 (I1885,I10061);
IN_INSTANCE I_518 (I1813,I10071);
IN_INSTANCE I_519 (I1581,I10081);
IN_INSTANCE I_520 (I1557,I10091);
IN_INSTANCE I_521 (I1549,I10101);
IN_INSTANCE I_522 (I1365,I10111);
IN_INSTANCE I_523 (I1421,I10121);
IN_INSTANCE I_524 (I1517,I10131);
IN_INSTANCE I_525 (I1717,I10141);
PAT_9 I_526 (I10041,I10051,I10061,I10071,I10081,I10091,I10101,I10111,I10121,I10131,I10141,I10181,I10184,I10187,I10190,I10193,I10196,I10199,I10202,I10205,I1892,I1899);
OUT_INSTANCE I_527 (I10181,I10221);
OUT_INSTANCE I_528 (I10184,I10231);
OUT_INSTANCE I_529 (I10187,I10241);
OUT_INSTANCE I_530 (I10190,I10251);
OUT_INSTANCE I_531 (I10193,I10261);
OUT_INSTANCE I_532 (I10196,I10271);
OUT_INSTANCE I_533 (I10199,I10281);
OUT_INSTANCE I_534 (I10202,I10291);
OUT_INSTANCE I_535 (I10205,I10301);
PAT_13 I_536 (I10221,I10291,I10231,I10281,I10261,I10251,I10301,I10221,I10241,I10271,I10231,I10341,I10344,I10347,I10350,I10353,I10356,I10359,I10362,I10365,I1892,I1899);
OUT_INSTANCE I_537 (I10341,I10381);
OUT_INSTANCE I_538 (I10344,I10391);
OUT_INSTANCE I_539 (I10347,I10401);
OUT_INSTANCE I_540 (I10350,I10411);
OUT_INSTANCE I_541 (I10353,I10421);
OUT_INSTANCE I_542 (I10356,I10431);
OUT_INSTANCE I_543 (I10359,I10441);
OUT_INSTANCE I_544 (I10362,I10451);
OUT_INSTANCE I_545 (I10365,I10461);
PAT_2 I_546 (I10441,I10421,I10411,I10431,I10381,I10461,I10391,I10451,I10381,I10401,I10391,I10501,I10504,I10507,I10510,I10513,I10516,I10519,I10522,I10525,I1892,I1899);
OUT_INSTANCE I_547 (I10501,I10541);
OUT_INSTANCE I_548 (I10504,I10551);
OUT_INSTANCE I_549 (I10507,I10561);
OUT_INSTANCE I_550 (I10510,I10571);
OUT_INSTANCE I_551 (I10513,I10581);
OUT_INSTANCE I_552 (I10516,I10591);
OUT_INSTANCE I_553 (I10519,I10601);
OUT_INSTANCE I_554 (I10522,I10611);
OUT_INSTANCE I_555 (I10525,I10621);
PAT_12 I_556 (I10571,I10561,I10541,I10551,I10621,I10601,I10611,I10551,I10591,I10541,I10581,I10661,I10664,I10667,I10670,I10673,I10676,I10679,I10682,I1892,I1899);
OUT_INSTANCE I_557 (I10661,I10698);
OUT_INSTANCE I_558 (I10664,I10708);
OUT_INSTANCE I_559 (I10667,I10718);
OUT_INSTANCE I_560 (I10670,I10728);
OUT_INSTANCE I_561 (I10673,I10738);
OUT_INSTANCE I_562 (I10676,I10748);
OUT_INSTANCE I_563 (I10679,I10758);
OUT_INSTANCE I_564 (I10682,I10768);
PAT_17 I_565 (I10748,I10728,I10708,I10698,I10698,I10718,I10718,I10758,I10768,I10708,I10738,I10808,I10811,I10814,I10817,I10820,I10823,I10826,I10829,I10832,I10835,I1892,I1899);
OUT_INSTANCE I_566 (I10808,I10851);
OUT_INSTANCE I_567 (I10811,I10861);
OUT_INSTANCE I_568 (I10814,I10871);
OUT_INSTANCE I_569 (I10817,I10881);
OUT_INSTANCE I_570 (I10820,I10891);
OUT_INSTANCE I_571 (I10823,I10901);
OUT_INSTANCE I_572 (I10826,I10911);
OUT_INSTANCE I_573 (I10829,I10921);
OUT_INSTANCE I_574 (I10832,I10931);
OUT_INSTANCE I_575 (I10835,I10941);
PAT_2 I_576 (I10851,I10911,I10901,I10851,I10881,I10931,I10921,I10871,I10941,I10891,I10861,I10981,I10984,I10987,I10990,I10993,I10996,I10999,I11002,I11005,I1892,I1899);
OUT_INSTANCE I_577 (I10981,I11021);
OUT_INSTANCE I_578 (I10984,I11031);
OUT_INSTANCE I_579 (I10987,I11041);
OUT_INSTANCE I_580 (I10990,I11051);
OUT_INSTANCE I_581 (I10993,I11061);
OUT_INSTANCE I_582 (I10996,I11071);
OUT_INSTANCE I_583 (I10999,I11081);
OUT_INSTANCE I_584 (I11002,I11091);
OUT_INSTANCE I_585 (I11005,I11101);
PAT_6 I_586 (I11101,I11021,I11071,I11061,I11081,I11051,I11031,I11091,I11021,I11041,I11031,I11141,I11144,I11147,I11150,I11153,I11156,I11159,I11162,I11165,I11168,I1892,I1899);
OUT_INSTANCE I_587 (I11141,I11184);
OUT_INSTANCE I_588 (I11144,I11194);
OUT_INSTANCE I_589 (I11147,I11204);
OUT_INSTANCE I_590 (I11150,I11214);
OUT_INSTANCE I_591 (I11153,I11224);
OUT_INSTANCE I_592 (I11156,I11234);
OUT_INSTANCE I_593 (I11159,I11244);
OUT_INSTANCE I_594 (I11162,I11254);
OUT_INSTANCE I_595 (I11165,I11264);
OUT_INSTANCE I_596 (I11168,I11274);
PAT_8 I_597 (I11214,I11234,I11204,I11244,I11184,I11194,I11254,I11184,I11274,I11264,I11224,I11314,I11317,I11320,I11323,I11326,I11329,I11332,I11335,I11338,I1892,I1899);
OUT_INSTANCE I_598 (I11314,I11354);
OUT_INSTANCE I_599 (I11317,I11364);
OUT_INSTANCE I_600 (I11320,I11374);
OUT_INSTANCE I_601 (I11323,I11384);
OUT_INSTANCE I_602 (I11326,I11394);
OUT_INSTANCE I_603 (I11329,I11404);
OUT_INSTANCE I_604 (I11332,I11414);
OUT_INSTANCE I_605 (I11335,I11424);
OUT_INSTANCE I_606 (I11338,I11434);
PAT_17 I_607 (I11434,I11394,I11384,I11364,I11374,I11414,I11354,I11364,I11354,I11404,I11424,I11474,I11477,I11480,I11483,I11486,I11489,I11492,I11495,I11498,I11501,I1892,I1899);
OUT_INSTANCE I_608 (I11474,I11517);
OUT_INSTANCE I_609 (I11477,I11527);
OUT_INSTANCE I_610 (I11480,I11537);
OUT_INSTANCE I_611 (I11483,I11547);
OUT_INSTANCE I_612 (I11486,I11557);
OUT_INSTANCE I_613 (I11489,I11567);
OUT_INSTANCE I_614 (I11492,I11577);
OUT_INSTANCE I_615 (I11495,I11587);
OUT_INSTANCE I_616 (I11498,I11597);
OUT_INSTANCE I_617 (I11501,I11607);
PAT_3 I_618 (I11557,I11567,I11577,I11587,I11517,I11517,I11537,I11597,I11607,I11547,I11527,I11647,I11650,I11653,I11656,I11659,I11662,I11665,I11668,I11671,I11674,I1892,I1899);
OUT_INSTANCE I_619 (I11647,I11690);
OUT_INSTANCE I_620 (I11650,I11700);
OUT_INSTANCE I_621 (I11653,I11710);
OUT_INSTANCE I_622 (I11656,I11720);
OUT_INSTANCE I_623 (I11659,I11730);
OUT_INSTANCE I_624 (I11662,I11740);
OUT_INSTANCE I_625 (I11665,I11750);
OUT_INSTANCE I_626 (I11668,I11760);
OUT_INSTANCE I_627 (I11671,I11770);
OUT_INSTANCE I_628 (I11674,I11780);
PAT_9 I_629 (I11690,I11770,I11710,I11760,I11720,I11700,I11750,I11780,I11690,I11730,I11740,I11820,I11823,I11826,I11829,I11832,I11835,I11838,I11841,I11844,I1892,I1899);
OUT_INSTANCE I_630 (I11820,I11860);
OUT_INSTANCE I_631 (I11823,I11870);
OUT_INSTANCE I_632 (I11826,I11880);
OUT_INSTANCE I_633 (I11829,I11890);
OUT_INSTANCE I_634 (I11832,I11900);
OUT_INSTANCE I_635 (I11835,I11910);
OUT_INSTANCE I_636 (I11838,I11920);
OUT_INSTANCE I_637 (I11841,I11930);
OUT_INSTANCE I_638 (I11844,I11940);
PAT_1 I_639 (I11860,I11920,I11860,I11900,I11870,I11890,I11910,I11930,I11940,I11880,I11870,I11980,I11983,I11986,I11989,I11992,I11995,I11998,I12001,I12004,I1892,I1899);
OUT_INSTANCE I_640 (I11980,I12020);
OUT_INSTANCE I_641 (I11983,I12030);
OUT_INSTANCE I_642 (I11986,I12040);
OUT_INSTANCE I_643 (I11989,I12050);
OUT_INSTANCE I_644 (I11992,I12060);
OUT_INSTANCE I_645 (I11995,I12070);
OUT_INSTANCE I_646 (I11998,I12080);
OUT_INSTANCE I_647 (I12001,I12090);
OUT_INSTANCE I_648 (I12004,I12100);
PAT_10 I_649 (I12070,I12060,I12030,I12020,I12030,I12080,I12040,I12090,I12100,I12050,I12020,I12140,I12143,I12146,I12149,I12152,I12155,I12158,I12161,I1892,I1899);
OUT_INSTANCE I_650 (I12140,I12177);
OUT_INSTANCE I_651 (I12143,I12187);
OUT_INSTANCE I_652 (I12146,I12197);
OUT_INSTANCE I_653 (I12149,I12207);
OUT_INSTANCE I_654 (I12152,I12217);
OUT_INSTANCE I_655 (I12155,I12227);
OUT_INSTANCE I_656 (I12158,I12237);
OUT_INSTANCE I_657 (I12161,I12247);
PAT_13 I_658 (I12197,I12217,I12197,I12187,I12237,I12247,I12177,I12177,I12227,I12187,I12207,I12287,I12290,I12293,I12296,I12299,I12302,I12305,I12308,I12311,I1892,I1899);
OUT_INSTANCE I_659 (I12287,I12327);
OUT_INSTANCE I_660 (I12290,I12337);
OUT_INSTANCE I_661 (I12293,I12347);
OUT_INSTANCE I_662 (I12296,I12357);
OUT_INSTANCE I_663 (I12299,I12367);
OUT_INSTANCE I_664 (I12302,I12377);
OUT_INSTANCE I_665 (I12305,I12387);
OUT_INSTANCE I_666 (I12308,I12397);
OUT_INSTANCE I_667 (I12311,I12407);
PAT_16 I_668 (I12347,I12357,I12387,I12367,I12407,I12327,I12397,I12377,I12337,I12337,I12327,I12447,I12450,I12453,I12456,I12459,I12462,I12465,I12468,I12471,I12474,I1892,I1899);
OUT_INSTANCE I_669 (I12447,I12490);
OUT_INSTANCE I_670 (I12450,I12500);
OUT_INSTANCE I_671 (I12453,I12510);
OUT_INSTANCE I_672 (I12456,I12520);
OUT_INSTANCE I_673 (I12459,I12530);
OUT_INSTANCE I_674 (I12462,I12540);
OUT_INSTANCE I_675 (I12465,I12550);
OUT_INSTANCE I_676 (I12468,I12560);
OUT_INSTANCE I_677 (I12471,I12570);
OUT_INSTANCE I_678 (I12474,I12580);
PAT_13 I_679 (I12530,I12500,I12490,I12510,I12540,I12570,I12560,I12550,I12520,I12490,I12580,I12620,I12623,I12626,I12629,I12632,I12635,I12638,I12641,I12644,I1892,I1899);
OUT_INSTANCE I_680 (I12620,I12660);
OUT_INSTANCE I_681 (I12623,I12670);
OUT_INSTANCE I_682 (I12626,I12680);
OUT_INSTANCE I_683 (I12629,I12690);
OUT_INSTANCE I_684 (I12632,I12700);
OUT_INSTANCE I_685 (I12635,I12710);
OUT_INSTANCE I_686 (I12638,I12720);
OUT_INSTANCE I_687 (I12641,I12730);
OUT_INSTANCE I_688 (I12644,I12740);
PAT_9 I_689 (I12730,I12670,I12670,I12660,I12740,I12680,I12690,I12660,I12700,I12720,I12710,I12780,I12783,I12786,I12789,I12792,I12795,I12798,I12801,I12804,I1892,I1899);
OUT_INSTANCE I_690 (I12780,I12820);
OUT_INSTANCE I_691 (I12783,I12830);
OUT_INSTANCE I_692 (I12786,I12840);
OUT_INSTANCE I_693 (I12789,I12850);
OUT_INSTANCE I_694 (I12792,I12860);
OUT_INSTANCE I_695 (I12795,I12870);
OUT_INSTANCE I_696 (I12798,I12880);
OUT_INSTANCE I_697 (I12801,I12890);
OUT_INSTANCE I_698 (I12804,I12900);
PAT_12 I_699 (I12890,I12880,I12860,I12820,I12850,I12820,I12830,I12840,I12900,I12870,I12830,I12940,I12943,I12946,I12949,I12952,I12955,I12958,I12961,I1892,I1899);
OUT_INSTANCE I_700 (I12940,I12977);
OUT_INSTANCE I_701 (I12943,I12987);
OUT_INSTANCE I_702 (I12946,I12997);
OUT_INSTANCE I_703 (I12949,I13007);
OUT_INSTANCE I_704 (I12952,I13017);
OUT_INSTANCE I_705 (I12955,I13027);
OUT_INSTANCE I_706 (I12958,I13037);
OUT_INSTANCE I_707 (I12961,I13047);
PAT_13 I_708 (I13017,I13027,I12997,I13047,I13037,I12977,I12987,I13007,I12997,I12987,I12977,I13087,I13090,I13093,I13096,I13099,I13102,I13105,I13108,I13111,I1892,I1899);
OUT_INSTANCE I_709 (I13087,I13127);
OUT_INSTANCE I_710 (I13090,I13137);
OUT_INSTANCE I_711 (I13093,I13147);
OUT_INSTANCE I_712 (I13096,I13157);
OUT_INSTANCE I_713 (I13099,I13167);
OUT_INSTANCE I_714 (I13102,I13177);
OUT_INSTANCE I_715 (I13105,I13187);
OUT_INSTANCE I_716 (I13108,I13197);
OUT_INSTANCE I_717 (I13111,I13207);
PAT_6 I_718 (I13127,I13167,I13157,I13197,I13187,I13207,I13127,I13177,I13137,I13137,I13147,I13247,I13250,I13253,I13256,I13259,I13262,I13265,I13268,I13271,I13274,I1892,I1899);
OUT_INSTANCE I_719 (I13247,I13290);
OUT_INSTANCE I_720 (I13250,I13300);
OUT_INSTANCE I_721 (I13253,I13310);
OUT_INSTANCE I_722 (I13256,I13320);
OUT_INSTANCE I_723 (I13259,I13330);
OUT_INSTANCE I_724 (I13262,I13340);
OUT_INSTANCE I_725 (I13265,I13350);
OUT_INSTANCE I_726 (I13268,I13360);
OUT_INSTANCE I_727 (I13271,I13370);
OUT_INSTANCE I_728 (I13274,I13380);
PAT_13 I_729 (I13370,I13310,I13360,I13290,I13300,I13320,I13380,I13330,I13350,I13290,I13340,I13420,I13423,I13426,I13429,I13432,I13435,I13438,I13441,I13444,I1892,I1899);
OUT_INSTANCE I_730 (I13420,I13460);
OUT_INSTANCE I_731 (I13423,I13470);
OUT_INSTANCE I_732 (I13426,I13480);
OUT_INSTANCE I_733 (I13429,I13490);
OUT_INSTANCE I_734 (I13432,I13500);
OUT_INSTANCE I_735 (I13435,I13510);
OUT_INSTANCE I_736 (I13438,I13520);
OUT_INSTANCE I_737 (I13441,I13530);
OUT_INSTANCE I_738 (I13444,I13540);
PAT_6 I_739 (I13460,I13500,I13490,I13530,I13520,I13540,I13460,I13510,I13470,I13470,I13480,I13580,I13583,I13586,I13589,I13592,I13595,I13598,I13601,I13604,I13607,I1892,I1899);
OUT_INSTANCE I_740 (I13580,I13623);
OUT_INSTANCE I_741 (I13583,I13633);
OUT_INSTANCE I_742 (I13586,I13643);
OUT_INSTANCE I_743 (I13589,I13653);
OUT_INSTANCE I_744 (I13592,I13663);
OUT_INSTANCE I_745 (I13595,I13673);
OUT_INSTANCE I_746 (I13598,I13683);
OUT_INSTANCE I_747 (I13601,I13693);
OUT_INSTANCE I_748 (I13604,I13703);
OUT_INSTANCE I_749 (I13607,I13713);
PAT_2 I_750 (I13693,I13713,I13653,I13673,I13623,I13643,I13623,I13663,I13633,I13683,I13703,I13753,I13756,I13759,I13762,I13765,I13768,I13771,I13774,I13777,I1892,I1899);
OUT_INSTANCE I_751 (I13753,I13793);
OUT_INSTANCE I_752 (I13756,I13803);
OUT_INSTANCE I_753 (I13759,I13813);
OUT_INSTANCE I_754 (I13762,I13823);
OUT_INSTANCE I_755 (I13765,I13833);
OUT_INSTANCE I_756 (I13768,I13843);
OUT_INSTANCE I_757 (I13771,I13853);
OUT_INSTANCE I_758 (I13774,I13863);
OUT_INSTANCE I_759 (I13777,I13873);
PAT_11 I_760 (I13803,I13843,I13793,I13833,I13823,I13863,I13853,I13803,I13873,I13813,I13793,I13913,I13916,I13919,I13922,I13925,I13928,I13931,I13934,I13937,I13940,I1892,I1899);
OUT_INSTANCE I_761 (I13913,I13956);
OUT_INSTANCE I_762 (I13916,I13966);
OUT_INSTANCE I_763 (I13919,I13976);
OUT_INSTANCE I_764 (I13922,I13986);
OUT_INSTANCE I_765 (I13925,I13996);
OUT_INSTANCE I_766 (I13928,I14006);
OUT_INSTANCE I_767 (I13931,I14016);
OUT_INSTANCE I_768 (I13934,I14026);
OUT_INSTANCE I_769 (I13937,I14036);
OUT_INSTANCE I_770 (I13940,I14046);
PAT_9 I_771 (I13976,I14016,I13986,I14026,I13956,I13966,I13996,I13956,I14006,I14036,I14046,I14086,I14089,I14092,I14095,I14098,I14101,I14104,I14107,I14110,I1892,I1899);
OUT_INSTANCE I_772 (I14086,I14126);
OUT_INSTANCE I_773 (I14089,I14136);
OUT_INSTANCE I_774 (I14092,I14146);
OUT_INSTANCE I_775 (I14095,I14156);
OUT_INSTANCE I_776 (I14098,I14166);
OUT_INSTANCE I_777 (I14101,I14176);
OUT_INSTANCE I_778 (I14104,I14186);
OUT_INSTANCE I_779 (I14107,I14196);
OUT_INSTANCE I_780 (I14110,I14206);
PAT_10 I_781 (I14196,I14186,I14146,I14136,I14206,I14156,I14176,I14136,I14126,I14126,I14166,I14246,I14249,I14252,I14255,I14258,I14261,I14264,I14267,I1892,I1899);
OUT_INSTANCE I_782 (I14246,I14283);
OUT_INSTANCE I_783 (I14249,I14293);
OUT_INSTANCE I_784 (I14252,I14303);
OUT_INSTANCE I_785 (I14255,I14313);
OUT_INSTANCE I_786 (I14258,I14323);
OUT_INSTANCE I_787 (I14261,I14333);
OUT_INSTANCE I_788 (I14264,I14343);
OUT_INSTANCE I_789 (I14267,I14353);
PAT_13 I_790 (I14303,I14323,I14303,I14293,I14343,I14353,I14283,I14283,I14333,I14293,I14313,I14393,I14396,I14399,I14402,I14405,I14408,I14411,I14414,I14417,I1892,I1899);
OUT_INSTANCE I_791 (I14393,I14433);
OUT_INSTANCE I_792 (I14396,I14443);
OUT_INSTANCE I_793 (I14399,I14453);
OUT_INSTANCE I_794 (I14402,I14463);
OUT_INSTANCE I_795 (I14405,I14473);
OUT_INSTANCE I_796 (I14408,I14483);
OUT_INSTANCE I_797 (I14411,I14493);
OUT_INSTANCE I_798 (I14414,I14503);
OUT_INSTANCE I_799 (I14417,I14513);
PAT_1 I_800 (I14433,I14463,I14443,I14503,I14483,I14453,I14493,I14473,I14443,I14513,I14433,I14553,I14556,I14559,I14562,I14565,I14568,I14571,I14574,I14577,I1892,I1899);
OUT_INSTANCE I_801 (I14553,I14593);
OUT_INSTANCE I_802 (I14556,I14603);
OUT_INSTANCE I_803 (I14559,I14613);
OUT_INSTANCE I_804 (I14562,I14623);
OUT_INSTANCE I_805 (I14565,I14633);
OUT_INSTANCE I_806 (I14568,I14643);
OUT_INSTANCE I_807 (I14571,I14653);
OUT_INSTANCE I_808 (I14574,I14663);
OUT_INSTANCE I_809 (I14577,I14673);
PAT_7 I_810 (I14603,I14623,I14613,I14633,I14653,I14643,I14673,I14663,I14603,I14593,I14593,I14713,I14716,I14719,I14722,I14725,I14728,I14731,I14734,I14737,I1892,I1899);
OUT_INSTANCE I_811 (I14713,I14753);
OUT_INSTANCE I_812 (I14716,I14763);
OUT_INSTANCE I_813 (I14719,I14773);
OUT_INSTANCE I_814 (I14722,I14783);
OUT_INSTANCE I_815 (I14725,I14793);
OUT_INSTANCE I_816 (I14728,I14803);
OUT_INSTANCE I_817 (I14731,I14813);
OUT_INSTANCE I_818 (I14734,I14823);
OUT_INSTANCE I_819 (I14737,I14833);
PAT_14 I_820 (I14803,I14783,I14753,I14763,I14793,I14813,I14773,I14823,I14763,I14753,I14833,I14873,I14876,I14879,I14882,I14885,I14888,I14891,I14894,I14897,I1892,I1899);
OUT_INSTANCE I_821 (I14873,I14913);
OUT_INSTANCE I_822 (I14876,I14923);
OUT_INSTANCE I_823 (I14879,I14933);
OUT_INSTANCE I_824 (I14882,I14943);
OUT_INSTANCE I_825 (I14885,I14953);
OUT_INSTANCE I_826 (I14888,I14963);
OUT_INSTANCE I_827 (I14891,I14973);
OUT_INSTANCE I_828 (I14894,I14983);
OUT_INSTANCE I_829 (I14897,I14993);
PAT_5 I_830 (I14923,I14933,I14923,I14953,I14913,I14983,I14943,I14913,I14993,I14973,I14963,I15033,I15036,I15039,I15042,I15045,I15048,I15051,I15054,I15057,I15060,I1892,I1899);
OUT_INSTANCE I_831 (I15033,I15076);
OUT_INSTANCE I_832 (I15036,I15086);
OUT_INSTANCE I_833 (I15039,I15096);
OUT_INSTANCE I_834 (I15042,I15106);
OUT_INSTANCE I_835 (I15045,I15116);
OUT_INSTANCE I_836 (I15048,I15126);
OUT_INSTANCE I_837 (I15051,I15136);
OUT_INSTANCE I_838 (I15054,I15146);
OUT_INSTANCE I_839 (I15057,I15156);
OUT_INSTANCE I_840 (I15060,I15166);
PAT_6 I_841 (I15136,I15116,I15076,I15096,I15086,I15106,I15126,I15076,I15156,I15146,I15166,I15206,I15209,I15212,I15215,I15218,I15221,I15224,I15227,I15230,I15233,I1892,I1899);
OUT_INSTANCE I_842 (I15206,I15249);
OUT_INSTANCE I_843 (I15209,I15259);
OUT_INSTANCE I_844 (I15212,I15269);
OUT_INSTANCE I_845 (I15215,I15279);
OUT_INSTANCE I_846 (I15218,I15289);
OUT_INSTANCE I_847 (I15221,I15299);
OUT_INSTANCE I_848 (I15224,I15309);
OUT_INSTANCE I_849 (I15227,I15319);
OUT_INSTANCE I_850 (I15230,I15329);
OUT_INSTANCE I_851 (I15233,I15339);
PAT_15 I_852 (I15309,I15279,I15319,I15329,I15299,I15339,I15249,I15269,I15249,I15259,I15289,I15379,I15382,I15385,I15388,I15391,I15394,I15397,I15400,I15403,I1892,I1899);
OUT_INSTANCE I_853 (I15379,I15419);
OUT_INSTANCE I_854 (I15382,I15429);
OUT_INSTANCE I_855 (I15385,I15439);
OUT_INSTANCE I_856 (I15388,I15449);
OUT_INSTANCE I_857 (I15391,I15459);
OUT_INSTANCE I_858 (I15394,I15469);
OUT_INSTANCE I_859 (I15397,I15479);
OUT_INSTANCE I_860 (I15400,I15489);
OUT_INSTANCE I_861 (I15403,I15499);
PAT_5 I_862 (I15429,I15419,I15439,I15499,I15489,I15449,I15479,I15459,I15429,I15469,I15419,I15539,I15542,I15545,I15548,I15551,I15554,I15557,I15560,I15563,I15566,I1892,I1899);
OUT_INSTANCE I_863 (I15539,I15582);
OUT_INSTANCE I_864 (I15542,I15592);
OUT_INSTANCE I_865 (I15545,I15602);
OUT_INSTANCE I_866 (I15548,I15612);
OUT_INSTANCE I_867 (I15551,I15622);
OUT_INSTANCE I_868 (I15554,I15632);
OUT_INSTANCE I_869 (I15557,I15642);
OUT_INSTANCE I_870 (I15560,I15652);
OUT_INSTANCE I_871 (I15563,I15662);
OUT_INSTANCE I_872 (I15566,I15672);
PAT_7 I_873 (I15642,I15652,I15672,I15662,I15612,I15602,I15582,I15622,I15582,I15592,I15632,I15712,I15715,I15718,I15721,I15724,I15727,I15730,I15733,I15736,I1892,I1899);
OUT_INSTANCE I_874 (I15712,I15752);
OUT_INSTANCE I_875 (I15715,I15762);
OUT_INSTANCE I_876 (I15718,I15772);
OUT_INSTANCE I_877 (I15721,I15782);
OUT_INSTANCE I_878 (I15724,I15792);
OUT_INSTANCE I_879 (I15727,I15802);
OUT_INSTANCE I_880 (I15730,I15812);
OUT_INSTANCE I_881 (I15733,I15822);
OUT_INSTANCE I_882 (I15736,I15832);
PAT_4 I_883 (I15832,I15752,I15752,I15802,I15782,I15762,I15762,I15812,I15822,I15772,I15792,I15872,I15875,I15878,I15881,I15884,I15887,I15890,I15893,I15896,I1892,I1899);
OUT_INSTANCE I_884 (I15872,I15912);
OUT_INSTANCE I_885 (I15875,I15922);
OUT_INSTANCE I_886 (I15878,I15932);
OUT_INSTANCE I_887 (I15881,I15942);
OUT_INSTANCE I_888 (I15884,I15952);
OUT_INSTANCE I_889 (I15887,I15962);
OUT_INSTANCE I_890 (I15890,I15972);
OUT_INSTANCE I_891 (I15893,I15982);
OUT_INSTANCE I_892 (I15896,I15992);
PAT_8 I_893 (I15952,I15912,I15982,I15932,I15922,I15992,I15942,I15972,I15922,I15912,I15962,I16032,I16035,I16038,I16041,I16044,I16047,I16050,I16053,I16056,I1892,I1899);
OUT_INSTANCE I_894 (I16032,I16072);
OUT_INSTANCE I_895 (I16035,I16082);
OUT_INSTANCE I_896 (I16038,I16092);
OUT_INSTANCE I_897 (I16041,I16102);
OUT_INSTANCE I_898 (I16044,I16112);
OUT_INSTANCE I_899 (I16047,I16122);
OUT_INSTANCE I_900 (I16050,I16132);
OUT_INSTANCE I_901 (I16053,I16142);
OUT_INSTANCE I_902 (I16056,I16152);
PAT_2 I_903 (I16082,I16132,I16152,I16072,I16112,I16122,I16082,I16142,I16092,I16102,I16072,I16192,I16195,I16198,I16201,I16204,I16207,I16210,I16213,I16216,I1892,I1899);
OUT_INSTANCE I_904 (I16192,I16232);
OUT_INSTANCE I_905 (I16195,I16242);
OUT_INSTANCE I_906 (I16198,I16252);
OUT_INSTANCE I_907 (I16201,I16262);
OUT_INSTANCE I_908 (I16204,I16272);
OUT_INSTANCE I_909 (I16207,I16282);
OUT_INSTANCE I_910 (I16210,I16292);
OUT_INSTANCE I_911 (I16213,I16302);
OUT_INSTANCE I_912 (I16216,I16312);
PAT_4 I_913 (I16232,I16252,I16312,I16292,I16282,I16272,I16242,I16302,I16232,I16242,I16262,I16352,I16355,I16358,I16361,I16364,I16367,I16370,I16373,I16376,I1892,I1899);
OUT_INSTANCE I_914 (I16352,I16392);
OUT_INSTANCE I_915 (I16355,I16402);
OUT_INSTANCE I_916 (I16358,I16412);
OUT_INSTANCE I_917 (I16361,I16422);
OUT_INSTANCE I_918 (I16364,I16432);
OUT_INSTANCE I_919 (I16367,I16442);
OUT_INSTANCE I_920 (I16370,I16452);
OUT_INSTANCE I_921 (I16373,I16462);
OUT_INSTANCE I_922 (I16376,I16472);
PAT_5 I_923 (I16462,I16402,I16402,I16442,I16452,I16432,I16422,I16392,I16412,I16392,I16472,I16512,I16515,I16518,I16521,I16524,I16527,I16530,I16533,I16536,I16539,I1892,I1899);
OUT_INSTANCE I_924 (I16512,I16555);
OUT_INSTANCE I_925 (I16515,I16565);
OUT_INSTANCE I_926 (I16518,I16575);
OUT_INSTANCE I_927 (I16521,I16585);
OUT_INSTANCE I_928 (I16524,I16595);
OUT_INSTANCE I_929 (I16527,I16605);
OUT_INSTANCE I_930 (I16530,I16615);
OUT_INSTANCE I_931 (I16533,I16625);
OUT_INSTANCE I_932 (I16536,I16635);
OUT_INSTANCE I_933 (I16539,I16645);
PAT_9 I_934 (I16605,I16595,I16625,I16615,I16585,I16555,I16575,I16645,I16565,I16635,I16555,I16685,I16688,I16691,I16694,I16697,I16700,I16703,I16706,I16709,I1892,I1899);
OUT_INSTANCE I_935 (I16685,I16725);
OUT_INSTANCE I_936 (I16688,I16735);
OUT_INSTANCE I_937 (I16691,I16745);
OUT_INSTANCE I_938 (I16694,I16755);
OUT_INSTANCE I_939 (I16697,I16765);
OUT_INSTANCE I_940 (I16700,I16775);
OUT_INSTANCE I_941 (I16703,I16785);
OUT_INSTANCE I_942 (I16706,I16795);
OUT_INSTANCE I_943 (I16709,I16805);
PAT_8 I_944 (I16795,I16755,I16785,I16725,I16735,I16775,I16805,I16735,I16745,I16765,I16725,I16845,I16848,I16851,I16854,I16857,I16860,I16863,I16866,I16869,I1892,I1899);
OUT_INSTANCE I_945 (I16845,I16885);
OUT_INSTANCE I_946 (I16848,I16895);
OUT_INSTANCE I_947 (I16851,I16905);
OUT_INSTANCE I_948 (I16854,I16915);
OUT_INSTANCE I_949 (I16857,I16925);
OUT_INSTANCE I_950 (I16860,I16935);
OUT_INSTANCE I_951 (I16863,I16945);
OUT_INSTANCE I_952 (I16866,I16955);
OUT_INSTANCE I_953 (I16869,I16965);
PAT_13 I_954 (I16925,I16955,I16895,I16965,I16905,I16885,I16885,I16915,I16945,I16935,I16895,I17005,I17008,I17011,I17014,I17017,I17020,I17023,I17026,I17029,I1892,I1899);
OUT_INSTANCE I_955 (I17005,I17045);
OUT_INSTANCE I_956 (I17008,I17055);
OUT_INSTANCE I_957 (I17011,I17065);
OUT_INSTANCE I_958 (I17014,I17075);
OUT_INSTANCE I_959 (I17017,I17085);
OUT_INSTANCE I_960 (I17020,I17095);
OUT_INSTANCE I_961 (I17023,I17105);
OUT_INSTANCE I_962 (I17026,I17115);
OUT_INSTANCE I_963 (I17029,I17125);
PAT_4 I_964 (I17075,I17085,I17125,I17065,I17115,I17105,I17055,I17095,I17055,I17045,I17045,I17165,I17168,I17171,I17174,I17177,I17180,I17183,I17186,I17189,I1892,I1899);
OUT_INSTANCE I_965 (I17165,I17205);
OUT_INSTANCE I_966 (I17168,I17215);
OUT_INSTANCE I_967 (I17171,I17225);
OUT_INSTANCE I_968 (I17174,I17235);
OUT_INSTANCE I_969 (I17177,I17245);
OUT_INSTANCE I_970 (I17180,I17255);
OUT_INSTANCE I_971 (I17183,I17265);
OUT_INSTANCE I_972 (I17186,I17275);
OUT_INSTANCE I_973 (I17189,I17285);
PAT_9 I_974 (I17275,I17215,I17225,I17255,I17265,I17205,I17235,I17215,I17285,I17205,I17245,I17325,I17328,I17331,I17334,I17337,I17340,I17343,I17346,I17349,I1892,I1899);
OUT_INSTANCE I_975 (I17325,I17365);
OUT_INSTANCE I_976 (I17328,I17375);
OUT_INSTANCE I_977 (I17331,I17385);
OUT_INSTANCE I_978 (I17334,I17395);
OUT_INSTANCE I_979 (I17337,I17405);
OUT_INSTANCE I_980 (I17340,I17415);
OUT_INSTANCE I_981 (I17343,I17425);
OUT_INSTANCE I_982 (I17346,I17435);
OUT_INSTANCE I_983 (I17349,I17445);
PAT_13 I_984 (I17365,I17435,I17375,I17425,I17405,I17395,I17445,I17365,I17385,I17415,I17375,I17485,I17488,I17491,I17494,I17497,I17500,I17503,I17506,I17509,I1892,I1899);
OUT_INSTANCE I_985 (I17485,I17525);
OUT_INSTANCE I_986 (I17488,I17535);
OUT_INSTANCE I_987 (I17491,I17545);
OUT_INSTANCE I_988 (I17494,I17555);
OUT_INSTANCE I_989 (I17497,I17565);
OUT_INSTANCE I_990 (I17500,I17575);
OUT_INSTANCE I_991 (I17503,I17585);
OUT_INSTANCE I_992 (I17506,I17595);
OUT_INSTANCE I_993 (I17509,I17605);
PAT_4 I_994 (I17555,I17565,I17605,I17545,I17595,I17585,I17535,I17575,I17535,I17525,I17525,I17645,I17648,I17651,I17654,I17657,I17660,I17663,I17666,I17669,I1892,I1899);
OUT_INSTANCE I_995 (I17645,I17685);
OUT_INSTANCE I_996 (I17648,I17695);
OUT_INSTANCE I_997 (I17651,I17705);
OUT_INSTANCE I_998 (I17654,I17715);
OUT_INSTANCE I_999 (I17657,I17725);
OUT_INSTANCE I_1000 (I17660,I17735);
OUT_INSTANCE I_1001 (I17663,I17745);
OUT_INSTANCE I_1002 (I17666,I17755);
OUT_INSTANCE I_1003 (I17669,I17765);
PAT_5 I_1004 (I17755,I17695,I17695,I17735,I17745,I17725,I17715,I17685,I17705,I17685,I17765,I17805,I17808,I17811,I17814,I17817,I17820,I17823,I17826,I17829,I17832,I1892,I1899);
OUT_INSTANCE I_1005 (I17805,I17848);
OUT_INSTANCE I_1006 (I17808,I17858);
OUT_INSTANCE I_1007 (I17811,I17868);
OUT_INSTANCE I_1008 (I17814,I17878);
OUT_INSTANCE I_1009 (I17817,I17888);
OUT_INSTANCE I_1010 (I17820,I17898);
OUT_INSTANCE I_1011 (I17823,I17908);
OUT_INSTANCE I_1012 (I17826,I17918);
OUT_INSTANCE I_1013 (I17829,I17928);
OUT_INSTANCE I_1014 (I17832,I17938);
PAT_2 I_1015 (I17898,I17848,I17888,I17868,I17918,I17858,I17908,I17878,I17928,I17938,I17848,I17978,I17981,I17984,I17987,I17990,I17993,I17996,I17999,I18002,I1892,I1899);
OUT_INSTANCE I_1016 (I17978,I18018);
OUT_INSTANCE I_1017 (I17981,I18028);
OUT_INSTANCE I_1018 (I17984,I18038);
OUT_INSTANCE I_1019 (I17987,I18048);
OUT_INSTANCE I_1020 (I17990,I18058);
OUT_INSTANCE I_1021 (I17993,I18068);
OUT_INSTANCE I_1022 (I17996,I18078);
OUT_INSTANCE I_1023 (I17999,I18088);
OUT_INSTANCE I_1024 (I18002,I18098);
IN_INSTANCE I_1025 (I1589,I18108);
IN_INSTANCE I_1026 (I1621,I18118);
IN_INSTANCE I_1027 (I1821,I18128);
IN_INSTANCE I_1028 (I1781,I18138);
IN_INSTANCE I_1029 (I1645,I18148);
IN_INSTANCE I_1030 (I1845,I18158);
IN_INSTANCE I_1031 (I1477,I18168);
IN_INSTANCE I_1032 (I1637,I18178);
IN_INSTANCE I_1033 (I1861,I18188);
IN_INSTANCE I_1034 (I1413,I18198);
IN_INSTANCE I_1035 (I1789,I18208);
PAT_2 I_1036 (I18108,I18118,I18128,I18138,I18148,I18158,I18168,I18178,I18188,I18198,I18208,I18248,I18251,I18254,I18257,I18260,I18263,I18266,I18269,I18272,I1892,I1899);
OUT_INSTANCE I_1037 (I18248,I18288);
OUT_INSTANCE I_1038 (I18251,I18298);
OUT_INSTANCE I_1039 (I18254,I18308);
OUT_INSTANCE I_1040 (I18257,I18318);
OUT_INSTANCE I_1041 (I18260,I18328);
OUT_INSTANCE I_1042 (I18263,I18338);
OUT_INSTANCE I_1043 (I18266,I18348);
OUT_INSTANCE I_1044 (I18269,I18358);
OUT_INSTANCE I_1045 (I18272,I18368);
PAT_9 I_1046 (I18338,I18368,I18288,I18308,I18318,I18348,I18298,I18328,I18358,I18298,I18288,I18408,I18411,I18414,I18417,I18420,I18423,I18426,I18429,I18432,I1892,I1899);
OUT_INSTANCE I_1047 (I18408,I18448);
OUT_INSTANCE I_1048 (I18411,I18458);
OUT_INSTANCE I_1049 (I18414,I18468);
OUT_INSTANCE I_1050 (I18417,I18478);
OUT_INSTANCE I_1051 (I18420,I18488);
OUT_INSTANCE I_1052 (I18423,I18498);
OUT_INSTANCE I_1053 (I18426,I18508);
OUT_INSTANCE I_1054 (I18429,I18518);
OUT_INSTANCE I_1055 (I18432,I18528);
PAT_2 I_1056 (I18498,I18508,I18478,I18528,I18448,I18458,I18468,I18458,I18518,I18488,I18448,I18568,I18571,I18574,I18577,I18580,I18583,I18586,I18589,I18592,I1892,I1899);
OUT_INSTANCE I_1057 (I18568,I18608);
OUT_INSTANCE I_1058 (I18571,I18618);
OUT_INSTANCE I_1059 (I18574,I18628);
OUT_INSTANCE I_1060 (I18577,I18638);
OUT_INSTANCE I_1061 (I18580,I18648);
OUT_INSTANCE I_1062 (I18583,I18658);
OUT_INSTANCE I_1063 (I18586,I18668);
OUT_INSTANCE I_1064 (I18589,I18678);
OUT_INSTANCE I_1065 (I18592,I18688);
PAT_8 I_1066 (I18648,I18618,I18638,I18608,I18628,I18678,I18668,I18608,I18658,I18618,I18688,I18728,I18731,I18734,I18737,I18740,I18743,I18746,I18749,I18752,I1892,I1899);
OUT_INSTANCE I_1067 (I18728,I18768);
OUT_INSTANCE I_1068 (I18731,I18778);
OUT_INSTANCE I_1069 (I18734,I18788);
OUT_INSTANCE I_1070 (I18737,I18798);
OUT_INSTANCE I_1071 (I18740,I18808);
OUT_INSTANCE I_1072 (I18743,I18818);
OUT_INSTANCE I_1073 (I18746,I18828);
OUT_INSTANCE I_1074 (I18749,I18838);
OUT_INSTANCE I_1075 (I18752,I18848);
PAT_0 I_1076 (I18768,I18828,I18798,I18848,I18808,I18768,I18778,I18788,I18818,I18778,I18838,I18888,I18891,I18894,I18897,I18900,I18903,I18906,I18909,I1892,I1899);
OUT_INSTANCE I_1077 (I18888,I18925);
OUT_INSTANCE I_1078 (I18891,I18935);
OUT_INSTANCE I_1079 (I18894,I18945);
OUT_INSTANCE I_1080 (I18897,I18955);
OUT_INSTANCE I_1081 (I18900,I18965);
OUT_INSTANCE I_1082 (I18903,I18975);
OUT_INSTANCE I_1083 (I18906,I18985);
OUT_INSTANCE I_1084 (I18909,I18995);
PAT_1 I_1085 (I18935,I18925,I18925,I18985,I18935,I18965,I18945,I18975,I18955,I18995,I18945,I19035,I19038,I19041,I19044,I19047,I19050,I19053,I19056,I19059,I1892,I1899);
OUT_INSTANCE I_1086 (I19035,I19075);
OUT_INSTANCE I_1087 (I19038,I19085);
OUT_INSTANCE I_1088 (I19041,I19095);
OUT_INSTANCE I_1089 (I19044,I19105);
OUT_INSTANCE I_1090 (I19047,I19115);
OUT_INSTANCE I_1091 (I19050,I19125);
OUT_INSTANCE I_1092 (I19053,I19135);
OUT_INSTANCE I_1093 (I19056,I19145);
OUT_INSTANCE I_1094 (I19059,I19155);
PAT_11 I_1095 (I19085,I19135,I19125,I19145,I19155,I19085,I19105,I19115,I19075,I19095,I19075,I19195,I19198,I19201,I19204,I19207,I19210,I19213,I19216,I19219,I19222,I1892,I1899);
OUT_INSTANCE I_1096 (I19195,I19238);
OUT_INSTANCE I_1097 (I19198,I19248);
OUT_INSTANCE I_1098 (I19201,I19258);
OUT_INSTANCE I_1099 (I19204,I19268);
OUT_INSTANCE I_1100 (I19207,I19278);
OUT_INSTANCE I_1101 (I19210,I19288);
OUT_INSTANCE I_1102 (I19213,I19298);
OUT_INSTANCE I_1103 (I19216,I19308);
OUT_INSTANCE I_1104 (I19219,I19318);
OUT_INSTANCE I_1105 (I19222,I19328);
PAT_4 I_1106 (I19258,I19328,I19238,I19298,I19268,I19238,I19308,I19248,I19278,I19318,I19288,I19368,I19371,I19374,I19377,I19380,I19383,I19386,I19389,I19392,I1892,I1899);
OUT_INSTANCE I_1107 (I19368,I19408);
OUT_INSTANCE I_1108 (I19371,I19418);
OUT_INSTANCE I_1109 (I19374,I19428);
OUT_INSTANCE I_1110 (I19377,I19438);
OUT_INSTANCE I_1111 (I19380,I19448);
OUT_INSTANCE I_1112 (I19383,I19458);
OUT_INSTANCE I_1113 (I19386,I19468);
OUT_INSTANCE I_1114 (I19389,I19478);
OUT_INSTANCE I_1115 (I19392,I19488);
PAT_13 I_1116 (I19458,I19438,I19478,I19428,I19448,I19408,I19488,I19468,I19418,I19408,I19418,I19528,I19531,I19534,I19537,I19540,I19543,I19546,I19549,I19552,I1892,I1899);
OUT_INSTANCE I_1117 (I19528,I19568);
OUT_INSTANCE I_1118 (I19531,I19578);
OUT_INSTANCE I_1119 (I19534,I19588);
OUT_INSTANCE I_1120 (I19537,I19598);
OUT_INSTANCE I_1121 (I19540,I19608);
OUT_INSTANCE I_1122 (I19543,I19618);
OUT_INSTANCE I_1123 (I19546,I19628);
OUT_INSTANCE I_1124 (I19549,I19638);
OUT_INSTANCE I_1125 (I19552,I19648);
PAT_1 I_1126 (I19568,I19598,I19578,I19638,I19618,I19588,I19628,I19608,I19578,I19648,I19568,I19688,I19691,I19694,I19697,I19700,I19703,I19706,I19709,I19712,I1892,I1899);
OUT_INSTANCE I_1127 (I19688,I19728);
OUT_INSTANCE I_1128 (I19691,I19738);
OUT_INSTANCE I_1129 (I19694,I19748);
OUT_INSTANCE I_1130 (I19697,I19758);
OUT_INSTANCE I_1131 (I19700,I19768);
OUT_INSTANCE I_1132 (I19703,I19778);
OUT_INSTANCE I_1133 (I19706,I19788);
OUT_INSTANCE I_1134 (I19709,I19798);
OUT_INSTANCE I_1135 (I19712,I19808);
PAT_10 I_1136 (I19778,I19768,I19738,I19728,I19738,I19788,I19748,I19798,I19808,I19758,I19728,I19848,I19851,I19854,I19857,I19860,I19863,I19866,I19869,I1892,I1899);
OUT_INSTANCE I_1137 (I19848,I19885);
OUT_INSTANCE I_1138 (I19851,I19895);
OUT_INSTANCE I_1139 (I19854,I19905);
OUT_INSTANCE I_1140 (I19857,I19915);
OUT_INSTANCE I_1141 (I19860,I19925);
OUT_INSTANCE I_1142 (I19863,I19935);
OUT_INSTANCE I_1143 (I19866,I19945);
OUT_INSTANCE I_1144 (I19869,I19955);
PAT_13 I_1145 (I19905,I19925,I19905,I19895,I19945,I19955,I19885,I19885,I19935,I19895,I19915,I19995,I19998,I20001,I20004,I20007,I20010,I20013,I20016,I20019,I1892,I1899);
OUT_INSTANCE I_1146 (I19995,I20035);
OUT_INSTANCE I_1147 (I19998,I20045);
OUT_INSTANCE I_1148 (I20001,I20055);
OUT_INSTANCE I_1149 (I20004,I20065);
OUT_INSTANCE I_1150 (I20007,I20075);
OUT_INSTANCE I_1151 (I20010,I20085);
OUT_INSTANCE I_1152 (I20013,I20095);
OUT_INSTANCE I_1153 (I20016,I20105);
OUT_INSTANCE I_1154 (I20019,I20115);
PAT_12 I_1155 (I20065,I20035,I20035,I20115,I20105,I20045,I20095,I20075,I20045,I20055,I20085,I20155,I20158,I20161,I20164,I20167,I20170,I20173,I20176,I1892,I1899);
OUT_INSTANCE I_1156 (I20155,I20192);
OUT_INSTANCE I_1157 (I20158,I20202);
OUT_INSTANCE I_1158 (I20161,I20212);
OUT_INSTANCE I_1159 (I20164,I20222);
OUT_INSTANCE I_1160 (I20167,I20232);
OUT_INSTANCE I_1161 (I20170,I20242);
OUT_INSTANCE I_1162 (I20173,I20252);
OUT_INSTANCE I_1163 (I20176,I20262);
PAT_14 I_1164 (I20212,I20202,I20202,I20242,I20222,I20262,I20192,I20232,I20192,I20252,I20212,I20302,I20305,I20308,I20311,I20314,I20317,I20320,I20323,I20326,I1892,I1899);
OUT_INSTANCE I_1165 (I20302,I20342);
OUT_INSTANCE I_1166 (I20305,I20352);
OUT_INSTANCE I_1167 (I20308,I20362);
OUT_INSTANCE I_1168 (I20311,I20372);
OUT_INSTANCE I_1169 (I20314,I20382);
OUT_INSTANCE I_1170 (I20317,I20392);
OUT_INSTANCE I_1171 (I20320,I20402);
OUT_INSTANCE I_1172 (I20323,I20412);
OUT_INSTANCE I_1173 (I20326,I20422);
PAT_11 I_1174 (I20382,I20372,I20362,I20342,I20352,I20352,I20392,I20342,I20412,I20422,I20402,I20462,I20465,I20468,I20471,I20474,I20477,I20480,I20483,I20486,I20489,I1892,I1899);
OUT_INSTANCE I_1175 (I20462,I20505);
OUT_INSTANCE I_1176 (I20465,I20515);
OUT_INSTANCE I_1177 (I20468,I20525);
OUT_INSTANCE I_1178 (I20471,I20535);
OUT_INSTANCE I_1179 (I20474,I20545);
OUT_INSTANCE I_1180 (I20477,I20555);
OUT_INSTANCE I_1181 (I20480,I20565);
OUT_INSTANCE I_1182 (I20483,I20575);
OUT_INSTANCE I_1183 (I20486,I20585);
OUT_INSTANCE I_1184 (I20489,I20595);
PAT_5 I_1185 (I20575,I20505,I20595,I20555,I20545,I20585,I20525,I20505,I20565,I20515,I20535,I20635,I20638,I20641,I20644,I20647,I20650,I20653,I20656,I20659,I20662,I1892,I1899);
OUT_INSTANCE I_1186 (I20635,I20678);
OUT_INSTANCE I_1187 (I20638,I20688);
OUT_INSTANCE I_1188 (I20641,I20698);
OUT_INSTANCE I_1189 (I20644,I20708);
OUT_INSTANCE I_1190 (I20647,I20718);
OUT_INSTANCE I_1191 (I20650,I20728);
OUT_INSTANCE I_1192 (I20653,I20738);
OUT_INSTANCE I_1193 (I20656,I20748);
OUT_INSTANCE I_1194 (I20659,I20758);
OUT_INSTANCE I_1195 (I20662,I20768);
PAT_17 I_1196 (I20768,I20688,I20698,I20708,I20678,I20718,I20678,I20758,I20738,I20728,I20748,I20808,I20811,I20814,I20817,I20820,I20823,I20826,I20829,I20832,I20835,I1892,I1899);
OUT_INSTANCE I_1197 (I20808,I20851);
OUT_INSTANCE I_1198 (I20811,I20861);
OUT_INSTANCE I_1199 (I20814,I20871);
OUT_INSTANCE I_1200 (I20817,I20881);
OUT_INSTANCE I_1201 (I20820,I20891);
OUT_INSTANCE I_1202 (I20823,I20901);
OUT_INSTANCE I_1203 (I20826,I20911);
OUT_INSTANCE I_1204 (I20829,I20921);
OUT_INSTANCE I_1205 (I20832,I20931);
OUT_INSTANCE I_1206 (I20835,I20941);
PAT_9 I_1207 (I20921,I20861,I20881,I20931,I20871,I20911,I20851,I20891,I20851,I20941,I20901,I20981,I20984,I20987,I20990,I20993,I20996,I20999,I21002,I21005,I1892,I1899);
OUT_INSTANCE I_1208 (I20981,I21021);
OUT_INSTANCE I_1209 (I20984,I21031);
OUT_INSTANCE I_1210 (I20987,I21041);
OUT_INSTANCE I_1211 (I20990,I21051);
OUT_INSTANCE I_1212 (I20993,I21061);
OUT_INSTANCE I_1213 (I20996,I21071);
OUT_INSTANCE I_1214 (I20999,I21081);
OUT_INSTANCE I_1215 (I21002,I21091);
OUT_INSTANCE I_1216 (I21005,I21101);
PAT_17 I_1217 (I21031,I21051,I21101,I21071,I21081,I21041,I21021,I21061,I21021,I21031,I21091,I21141,I21144,I21147,I21150,I21153,I21156,I21159,I21162,I21165,I21168,I1892,I1899);
OUT_INSTANCE I_1218 (I21141,I21184);
OUT_INSTANCE I_1219 (I21144,I21194);
OUT_INSTANCE I_1220 (I21147,I21204);
OUT_INSTANCE I_1221 (I21150,I21214);
OUT_INSTANCE I_1222 (I21153,I21224);
OUT_INSTANCE I_1223 (I21156,I21234);
OUT_INSTANCE I_1224 (I21159,I21244);
OUT_INSTANCE I_1225 (I21162,I21254);
OUT_INSTANCE I_1226 (I21165,I21264);
OUT_INSTANCE I_1227 (I21168,I21274);
PAT_4 I_1228 (I21214,I21184,I21244,I21234,I21274,I21264,I21194,I21184,I21204,I21224,I21254,I21314,I21317,I21320,I21323,I21326,I21329,I21332,I21335,I21338,I1892,I1899);
OUT_INSTANCE I_1229 (I21314,I21354);
OUT_INSTANCE I_1230 (I21317,I21364);
OUT_INSTANCE I_1231 (I21320,I21374);
OUT_INSTANCE I_1232 (I21323,I21384);
OUT_INSTANCE I_1233 (I21326,I21394);
OUT_INSTANCE I_1234 (I21329,I21404);
OUT_INSTANCE I_1235 (I21332,I21414);
OUT_INSTANCE I_1236 (I21335,I21424);
OUT_INSTANCE I_1237 (I21338,I21434);
PAT_12 I_1238 (I21354,I21364,I21424,I21434,I21404,I21374,I21394,I21384,I21354,I21414,I21364,I21474,I21477,I21480,I21483,I21486,I21489,I21492,I21495,I1892,I1899);
OUT_INSTANCE I_1239 (I21474,I21511);
OUT_INSTANCE I_1240 (I21477,I21521);
OUT_INSTANCE I_1241 (I21480,I21531);
OUT_INSTANCE I_1242 (I21483,I21541);
OUT_INSTANCE I_1243 (I21486,I21551);
OUT_INSTANCE I_1244 (I21489,I21561);
OUT_INSTANCE I_1245 (I21492,I21571);
OUT_INSTANCE I_1246 (I21495,I21581);
PAT_5 I_1247 (I21541,I21561,I21581,I21531,I21531,I21511,I21571,I21511,I21521,I21521,I21551,I21621,I21624,I21627,I21630,I21633,I21636,I21639,I21642,I21645,I21648,I1892,I1899);
OUT_INSTANCE I_1248 (I21621,I21664);
OUT_INSTANCE I_1249 (I21624,I21674);
OUT_INSTANCE I_1250 (I21627,I21684);
OUT_INSTANCE I_1251 (I21630,I21694);
OUT_INSTANCE I_1252 (I21633,I21704);
OUT_INSTANCE I_1253 (I21636,I21714);
OUT_INSTANCE I_1254 (I21639,I21724);
OUT_INSTANCE I_1255 (I21642,I21734);
OUT_INSTANCE I_1256 (I21645,I21744);
OUT_INSTANCE I_1257 (I21648,I21754);
PAT_9 I_1258 (I21714,I21704,I21734,I21724,I21694,I21664,I21684,I21754,I21674,I21744,I21664,I21794,I21797,I21800,I21803,I21806,I21809,I21812,I21815,I21818,I1892,I1899);
OUT_INSTANCE I_1259 (I21794,I21834);
OUT_INSTANCE I_1260 (I21797,I21844);
OUT_INSTANCE I_1261 (I21800,I21854);
OUT_INSTANCE I_1262 (I21803,I21864);
OUT_INSTANCE I_1263 (I21806,I21874);
OUT_INSTANCE I_1264 (I21809,I21884);
OUT_INSTANCE I_1265 (I21812,I21894);
OUT_INSTANCE I_1266 (I21815,I21904);
OUT_INSTANCE I_1267 (I21818,I21914);
PAT_13 I_1268 (I21834,I21904,I21844,I21894,I21874,I21864,I21914,I21834,I21854,I21884,I21844,I21954,I21957,I21960,I21963,I21966,I21969,I21972,I21975,I21978,I1892,I1899);
OUT_INSTANCE I_1269 (I21954,I21994);
OUT_INSTANCE I_1270 (I21957,I22004);
OUT_INSTANCE I_1271 (I21960,I22014);
OUT_INSTANCE I_1272 (I21963,I22024);
OUT_INSTANCE I_1273 (I21966,I22034);
OUT_INSTANCE I_1274 (I21969,I22044);
OUT_INSTANCE I_1275 (I21972,I22054);
OUT_INSTANCE I_1276 (I21975,I22064);
OUT_INSTANCE I_1277 (I21978,I22074);
PAT_6 I_1278 (I21994,I22034,I22024,I22064,I22054,I22074,I21994,I22044,I22004,I22004,I22014,I22114,I22117,I22120,I22123,I22126,I22129,I22132,I22135,I22138,I22141,I1892,I1899);
OUT_INSTANCE I_1279 (I22114,I22157);
OUT_INSTANCE I_1280 (I22117,I22167);
OUT_INSTANCE I_1281 (I22120,I22177);
OUT_INSTANCE I_1282 (I22123,I22187);
OUT_INSTANCE I_1283 (I22126,I22197);
OUT_INSTANCE I_1284 (I22129,I22207);
OUT_INSTANCE I_1285 (I22132,I22217);
OUT_INSTANCE I_1286 (I22135,I22227);
OUT_INSTANCE I_1287 (I22138,I22237);
OUT_INSTANCE I_1288 (I22141,I22247);
PAT_8 I_1289 (I22187,I22207,I22177,I22217,I22157,I22167,I22227,I22157,I22247,I22237,I22197,I22287,I22290,I22293,I22296,I22299,I22302,I22305,I22308,I22311,I1892,I1899);
OUT_INSTANCE I_1290 (I22287,I22327);
OUT_INSTANCE I_1291 (I22290,I22337);
OUT_INSTANCE I_1292 (I22293,I22347);
OUT_INSTANCE I_1293 (I22296,I22357);
OUT_INSTANCE I_1294 (I22299,I22367);
OUT_INSTANCE I_1295 (I22302,I22377);
OUT_INSTANCE I_1296 (I22305,I22387);
OUT_INSTANCE I_1297 (I22308,I22397);
OUT_INSTANCE I_1298 (I22311,I22407);
PAT_9 I_1299 (I22337,I22367,I22337,I22327,I22377,I22347,I22397,I22357,I22387,I22327,I22407,I22447,I22450,I22453,I22456,I22459,I22462,I22465,I22468,I22471,I1892,I1899);
OUT_INSTANCE I_1300 (I22447,I22487);
OUT_INSTANCE I_1301 (I22450,I22497);
OUT_INSTANCE I_1302 (I22453,I22507);
OUT_INSTANCE I_1303 (I22456,I22517);
OUT_INSTANCE I_1304 (I22459,I22527);
OUT_INSTANCE I_1305 (I22462,I22537);
OUT_INSTANCE I_1306 (I22465,I22547);
OUT_INSTANCE I_1307 (I22468,I22557);
OUT_INSTANCE I_1308 (I22471,I22567);
PAT_7 I_1309 (I22507,I22537,I22487,I22557,I22527,I22487,I22497,I22567,I22547,I22497,I22517,I22607,I22610,I22613,I22616,I22619,I22622,I22625,I22628,I22631,I1892,I1899);
OUT_INSTANCE I_1310 (I22607,I22647);
OUT_INSTANCE I_1311 (I22610,I22657);
OUT_INSTANCE I_1312 (I22613,I22667);
OUT_INSTANCE I_1313 (I22616,I22677);
OUT_INSTANCE I_1314 (I22619,I22687);
OUT_INSTANCE I_1315 (I22622,I22697);
OUT_INSTANCE I_1316 (I22625,I22707);
OUT_INSTANCE I_1317 (I22628,I22717);
OUT_INSTANCE I_1318 (I22631,I22727);
PAT_15 I_1319 (I22707,I22657,I22657,I22697,I22647,I22727,I22667,I22687,I22717,I22647,I22677,I22767,I22770,I22773,I22776,I22779,I22782,I22785,I22788,I22791,I1892,I1899);
OUT_INSTANCE I_1320 (I22767,I22807);
OUT_INSTANCE I_1321 (I22770,I22817);
OUT_INSTANCE I_1322 (I22773,I22827);
OUT_INSTANCE I_1323 (I22776,I22837);
OUT_INSTANCE I_1324 (I22779,I22847);
OUT_INSTANCE I_1325 (I22782,I22857);
OUT_INSTANCE I_1326 (I22785,I22867);
OUT_INSTANCE I_1327 (I22788,I22877);
OUT_INSTANCE I_1328 (I22791,I22887);
PAT_9 I_1329 (I22807,I22877,I22837,I22817,I22857,I22817,I22867,I22887,I22827,I22807,I22847,I22927,I22930,I22933,I22936,I22939,I22942,I22945,I22948,I22951,I1892,I1899);
OUT_INSTANCE I_1330 (I22927,I22967);
OUT_INSTANCE I_1331 (I22930,I22977);
OUT_INSTANCE I_1332 (I22933,I22987);
OUT_INSTANCE I_1333 (I22936,I22997);
OUT_INSTANCE I_1334 (I22939,I23007);
OUT_INSTANCE I_1335 (I22942,I23017);
OUT_INSTANCE I_1336 (I22945,I23027);
OUT_INSTANCE I_1337 (I22948,I23037);
OUT_INSTANCE I_1338 (I22951,I23047);
PAT_5 I_1339 (I23037,I22967,I23017,I22967,I22987,I22997,I22977,I22977,I23027,I23007,I23047,I23087,I23090,I23093,I23096,I23099,I23102,I23105,I23108,I23111,I23114,I1892,I1899);
OUT_INSTANCE I_1340 (I23087,I23130);
OUT_INSTANCE I_1341 (I23090,I23140);
OUT_INSTANCE I_1342 (I23093,I23150);
OUT_INSTANCE I_1343 (I23096,I23160);
OUT_INSTANCE I_1344 (I23099,I23170);
OUT_INSTANCE I_1345 (I23102,I23180);
OUT_INSTANCE I_1346 (I23105,I23190);
OUT_INSTANCE I_1347 (I23108,I23200);
OUT_INSTANCE I_1348 (I23111,I23210);
OUT_INSTANCE I_1349 (I23114,I23220);
PAT_13 I_1350 (I23150,I23180,I23130,I23140,I23210,I23160,I23200,I23130,I23190,I23220,I23170,I23260,I23263,I23266,I23269,I23272,I23275,I23278,I23281,I23284,I1892,I1899);
OUT_INSTANCE I_1351 (I23260,I23300);
OUT_INSTANCE I_1352 (I23263,I23310);
OUT_INSTANCE I_1353 (I23266,I23320);
OUT_INSTANCE I_1354 (I23269,I23330);
OUT_INSTANCE I_1355 (I23272,I23340);
OUT_INSTANCE I_1356 (I23275,I23350);
OUT_INSTANCE I_1357 (I23278,I23360);
OUT_INSTANCE I_1358 (I23281,I23370);
OUT_INSTANCE I_1359 (I23284,I23380);
PAT_12 I_1360 (I23330,I23300,I23300,I23380,I23370,I23310,I23360,I23340,I23310,I23320,I23350,I23420,I23423,I23426,I23429,I23432,I23435,I23438,I23441,I1892,I1899);
OUT_INSTANCE I_1361 (I23420,I23457);
OUT_INSTANCE I_1362 (I23423,I23467);
OUT_INSTANCE I_1363 (I23426,I23477);
OUT_INSTANCE I_1364 (I23429,I23487);
OUT_INSTANCE I_1365 (I23432,I23497);
OUT_INSTANCE I_1366 (I23435,I23507);
OUT_INSTANCE I_1367 (I23438,I23517);
OUT_INSTANCE I_1368 (I23441,I23527);
PAT_13 I_1369 (I23497,I23507,I23477,I23527,I23517,I23457,I23467,I23487,I23477,I23467,I23457,I23567,I23570,I23573,I23576,I23579,I23582,I23585,I23588,I23591,I1892,I1899);
OUT_INSTANCE I_1370 (I23567,I23607);
OUT_INSTANCE I_1371 (I23570,I23617);
OUT_INSTANCE I_1372 (I23573,I23627);
OUT_INSTANCE I_1373 (I23576,I23637);
OUT_INSTANCE I_1374 (I23579,I23647);
OUT_INSTANCE I_1375 (I23582,I23657);
OUT_INSTANCE I_1376 (I23585,I23667);
OUT_INSTANCE I_1377 (I23588,I23677);
OUT_INSTANCE I_1378 (I23591,I23687);
PAT_0 I_1379 (I23627,I23637,I23607,I23607,I23647,I23677,I23687,I23657,I23667,I23617,I23617,I23727,I23730,I23733,I23736,I23739,I23742,I23745,I23748,I1892,I1899);
OUT_INSTANCE I_1380 (I23727,I23764);
OUT_INSTANCE I_1381 (I23730,I23774);
OUT_INSTANCE I_1382 (I23733,I23784);
OUT_INSTANCE I_1383 (I23736,I23794);
OUT_INSTANCE I_1384 (I23739,I23804);
OUT_INSTANCE I_1385 (I23742,I23814);
OUT_INSTANCE I_1386 (I23745,I23824);
OUT_INSTANCE I_1387 (I23748,I23834);
PAT_13 I_1388 (I23794,I23824,I23764,I23774,I23774,I23784,I23804,I23784,I23764,I23814,I23834,I23874,I23877,I23880,I23883,I23886,I23889,I23892,I23895,I23898,I1892,I1899);
OUT_INSTANCE I_1389 (I23874,I23914);
OUT_INSTANCE I_1390 (I23877,I23924);
OUT_INSTANCE I_1391 (I23880,I23934);
OUT_INSTANCE I_1392 (I23883,I23944);
OUT_INSTANCE I_1393 (I23886,I23954);
OUT_INSTANCE I_1394 (I23889,I23964);
OUT_INSTANCE I_1395 (I23892,I23974);
OUT_INSTANCE I_1396 (I23895,I23984);
OUT_INSTANCE I_1397 (I23898,I23994);
PAT_6 I_1398 (I23914,I23954,I23944,I23984,I23974,I23994,I23914,I23964,I23924,I23924,I23934,I24034,I24037,I24040,I24043,I24046,I24049,I24052,I24055,I24058,I24061,I1892,I1899);
OUT_INSTANCE I_1399 (I24034,I24077);
OUT_INSTANCE I_1400 (I24037,I24087);
OUT_INSTANCE I_1401 (I24040,I24097);
OUT_INSTANCE I_1402 (I24043,I24107);
OUT_INSTANCE I_1403 (I24046,I24117);
OUT_INSTANCE I_1404 (I24049,I24127);
OUT_INSTANCE I_1405 (I24052,I24137);
OUT_INSTANCE I_1406 (I24055,I24147);
OUT_INSTANCE I_1407 (I24058,I24157);
OUT_INSTANCE I_1408 (I24061,I24167);
PAT_2 I_1409 (I24147,I24167,I24107,I24127,I24077,I24097,I24077,I24117,I24087,I24137,I24157,I24207,I24210,I24213,I24216,I24219,I24222,I24225,I24228,I24231,I1892,I1899);
OUT_INSTANCE I_1410 (I24207,I24247);
OUT_INSTANCE I_1411 (I24210,I24257);
OUT_INSTANCE I_1412 (I24213,I24267);
OUT_INSTANCE I_1413 (I24216,I24277);
OUT_INSTANCE I_1414 (I24219,I24287);
OUT_INSTANCE I_1415 (I24222,I24297);
OUT_INSTANCE I_1416 (I24225,I24307);
OUT_INSTANCE I_1417 (I24228,I24317);
OUT_INSTANCE I_1418 (I24231,I24327);
PAT_12 I_1419 (I24277,I24267,I24247,I24257,I24327,I24307,I24317,I24257,I24297,I24247,I24287,I24367,I24370,I24373,I24376,I24379,I24382,I24385,I24388,I1892,I1899);
OUT_INSTANCE I_1420 (I24367,I24404);
OUT_INSTANCE I_1421 (I24370,I24414);
OUT_INSTANCE I_1422 (I24373,I24424);
OUT_INSTANCE I_1423 (I24376,I24434);
OUT_INSTANCE I_1424 (I24379,I24444);
OUT_INSTANCE I_1425 (I24382,I24454);
OUT_INSTANCE I_1426 (I24385,I24464);
OUT_INSTANCE I_1427 (I24388,I24474);
PAT_13 I_1428 (I24444,I24454,I24424,I24474,I24464,I24404,I24414,I24434,I24424,I24414,I24404,I24514,I24517,I24520,I24523,I24526,I24529,I24532,I24535,I24538,I1892,I1899);
OUT_INSTANCE I_1429 (I24514,I24554);
OUT_INSTANCE I_1430 (I24517,I24564);
OUT_INSTANCE I_1431 (I24520,I24574);
OUT_INSTANCE I_1432 (I24523,I24584);
OUT_INSTANCE I_1433 (I24526,I24594);
OUT_INSTANCE I_1434 (I24529,I24604);
OUT_INSTANCE I_1435 (I24532,I24614);
OUT_INSTANCE I_1436 (I24535,I24624);
OUT_INSTANCE I_1437 (I24538,I24634);
PAT_4 I_1438 (I24584,I24594,I24634,I24574,I24624,I24614,I24564,I24604,I24564,I24554,I24554,I24674,I24677,I24680,I24683,I24686,I24689,I24692,I24695,I24698,I1892,I1899);
OUT_INSTANCE I_1439 (I24674,I24714);
OUT_INSTANCE I_1440 (I24677,I24724);
OUT_INSTANCE I_1441 (I24680,I24734);
OUT_INSTANCE I_1442 (I24683,I24744);
OUT_INSTANCE I_1443 (I24686,I24754);
OUT_INSTANCE I_1444 (I24689,I24764);
OUT_INSTANCE I_1445 (I24692,I24774);
OUT_INSTANCE I_1446 (I24695,I24784);
OUT_INSTANCE I_1447 (I24698,I24794);
PAT_5 I_1448 (I24784,I24724,I24724,I24764,I24774,I24754,I24744,I24714,I24734,I24714,I24794,I24834,I24837,I24840,I24843,I24846,I24849,I24852,I24855,I24858,I24861,I1892,I1899);
OUT_INSTANCE I_1449 (I24834,I24877);
OUT_INSTANCE I_1450 (I24837,I24887);
OUT_INSTANCE I_1451 (I24840,I24897);
OUT_INSTANCE I_1452 (I24843,I24907);
OUT_INSTANCE I_1453 (I24846,I24917);
OUT_INSTANCE I_1454 (I24849,I24927);
OUT_INSTANCE I_1455 (I24852,I24937);
OUT_INSTANCE I_1456 (I24855,I24947);
OUT_INSTANCE I_1457 (I24858,I24957);
OUT_INSTANCE I_1458 (I24861,I24967);
PAT_15 I_1459 (I24937,I24887,I24877,I24877,I24927,I24917,I24957,I24907,I24947,I24897,I24967,I25007,I25010,I25013,I25016,I25019,I25022,I25025,I25028,I25031,I1892,I1899);
OUT_INSTANCE I_1460 (I25007,I25047);
OUT_INSTANCE I_1461 (I25010,I25057);
OUT_INSTANCE I_1462 (I25013,I25067);
OUT_INSTANCE I_1463 (I25016,I25077);
OUT_INSTANCE I_1464 (I25019,I25087);
OUT_INSTANCE I_1465 (I25022,I25097);
OUT_INSTANCE I_1466 (I25025,I25107);
OUT_INSTANCE I_1467 (I25028,I25117);
OUT_INSTANCE I_1468 (I25031,I25127);
PAT_11 I_1469 (I25117,I25057,I25047,I25097,I25067,I25047,I25107,I25127,I25087,I25057,I25077,I25167,I25170,I25173,I25176,I25179,I25182,I25185,I25188,I25191,I25194,I1892,I1899);
OUT_INSTANCE I_1470 (I25167,I25210);
OUT_INSTANCE I_1471 (I25170,I25220);
OUT_INSTANCE I_1472 (I25173,I25230);
OUT_INSTANCE I_1473 (I25176,I25240);
OUT_INSTANCE I_1474 (I25179,I25250);
OUT_INSTANCE I_1475 (I25182,I25260);
OUT_INSTANCE I_1476 (I25185,I25270);
OUT_INSTANCE I_1477 (I25188,I25280);
OUT_INSTANCE I_1478 (I25191,I25290);
OUT_INSTANCE I_1479 (I25194,I25300);
PAT_4 I_1480 (I25230,I25300,I25210,I25270,I25240,I25210,I25280,I25220,I25250,I25290,I25260,I25340,I25343,I25346,I25349,I25352,I25355,I25358,I25361,I25364,I1892,I1899);
OUT_INSTANCE I_1481 (I25340,I25380);
OUT_INSTANCE I_1482 (I25343,I25390);
OUT_INSTANCE I_1483 (I25346,I25400);
OUT_INSTANCE I_1484 (I25349,I25410);
OUT_INSTANCE I_1485 (I25352,I25420);
OUT_INSTANCE I_1486 (I25355,I25430);
OUT_INSTANCE I_1487 (I25358,I25440);
OUT_INSTANCE I_1488 (I25361,I25450);
OUT_INSTANCE I_1489 (I25364,I25460);
PAT_7 I_1490 (I25430,I25410,I25400,I25380,I25420,I25440,I25390,I25390,I25450,I25460,I25380,I25500,I25503,I25506,I25509,I25512,I25515,I25518,I25521,I25524,I1892,I1899);
OUT_INSTANCE I_1491 (I25500,I25540);
OUT_INSTANCE I_1492 (I25503,I25550);
OUT_INSTANCE I_1493 (I25506,I25560);
OUT_INSTANCE I_1494 (I25509,I25570);
OUT_INSTANCE I_1495 (I25512,I25580);
OUT_INSTANCE I_1496 (I25515,I25590);
OUT_INSTANCE I_1497 (I25518,I25600);
OUT_INSTANCE I_1498 (I25521,I25610);
OUT_INSTANCE I_1499 (I25524,I25620);
PAT_10 I_1500 (I25540,I25550,I25540,I25610,I25570,I25580,I25550,I25620,I25590,I25560,I25600,I25660,I25663,I25666,I25669,I25672,I25675,I25678,I25681,I1892,I1899);
OUT_INSTANCE I_1501 (I25660,I25697);
OUT_INSTANCE I_1502 (I25663,I25707);
OUT_INSTANCE I_1503 (I25666,I25717);
OUT_INSTANCE I_1504 (I25669,I25727);
OUT_INSTANCE I_1505 (I25672,I25737);
OUT_INSTANCE I_1506 (I25675,I25747);
OUT_INSTANCE I_1507 (I25678,I25757);
OUT_INSTANCE I_1508 (I25681,I25767);
PAT_4 I_1509 (I25747,I25737,I25707,I25767,I25697,I25707,I25727,I25717,I25757,I25697,I25717,I25807,I25810,I25813,I25816,I25819,I25822,I25825,I25828,I25831,I1892,I1899);
OUT_INSTANCE I_1510 (I25807,I25847);
OUT_INSTANCE I_1511 (I25810,I25857);
OUT_INSTANCE I_1512 (I25813,I25867);
OUT_INSTANCE I_1513 (I25816,I25877);
OUT_INSTANCE I_1514 (I25819,I25887);
OUT_INSTANCE I_1515 (I25822,I25897);
OUT_INSTANCE I_1516 (I25825,I25907);
OUT_INSTANCE I_1517 (I25828,I25917);
OUT_INSTANCE I_1518 (I25831,I25927);
PAT_9 I_1519 (I25917,I25857,I25867,I25897,I25907,I25847,I25877,I25857,I25927,I25847,I25887,I25967,I25970,I25973,I25976,I25979,I25982,I25985,I25988,I25991,I1892,I1899);
OUT_INSTANCE I_1520 (I25967,I26007);
OUT_INSTANCE I_1521 (I25970,I26017);
OUT_INSTANCE I_1522 (I25973,I26027);
OUT_INSTANCE I_1523 (I25976,I26037);
OUT_INSTANCE I_1524 (I25979,I26047);
OUT_INSTANCE I_1525 (I25982,I26057);
OUT_INSTANCE I_1526 (I25985,I26067);
OUT_INSTANCE I_1527 (I25988,I26077);
OUT_INSTANCE I_1528 (I25991,I26087);
IN_INSTANCE I_1529 (I1397,I26097);
IN_INSTANCE I_1530 (I1869,I26107);
IN_INSTANCE I_1531 (I1661,I26117);
IN_INSTANCE I_1532 (I1453,I26127);
IN_INSTANCE I_1533 (I1525,I26137);
IN_INSTANCE I_1534 (I1805,I26147);
IN_INSTANCE I_1535 (I1677,I26157);
IN_INSTANCE I_1536 (I1757,I26167);
IN_INSTANCE I_1537 (I1541,I26177);
IN_INSTANCE I_1538 (I1877,I26187);
IN_INSTANCE I_1539 (I1613,I26197);
PAT_2 I_1540 (I26097,I26107,I26117,I26127,I26137,I26147,I26157,I26167,I26177,I26187,I26197,I26237,I26240,I26243,I26246,I26249,I26252,I26255,I26258,I26261,I1892,I1899);
OUT_INSTANCE I_1541 (I26237,I26277);
OUT_INSTANCE I_1542 (I26240,I26287);
OUT_INSTANCE I_1543 (I26243,I26297);
OUT_INSTANCE I_1544 (I26246,I26307);
OUT_INSTANCE I_1545 (I26249,I26317);
OUT_INSTANCE I_1546 (I26252,I26327);
OUT_INSTANCE I_1547 (I26255,I26337);
OUT_INSTANCE I_1548 (I26258,I26347);
OUT_INSTANCE I_1549 (I26261,I26357);
PAT_5 I_1550 (I26347,I26277,I26277,I26317,I26307,I26337,I26297,I26327,I26357,I26287,I26287,I26397,I26400,I26403,I26406,I26409,I26412,I26415,I26418,I26421,I26424,I1892,I1899);
OUT_INSTANCE I_1551 (I26397,I26440);
OUT_INSTANCE I_1552 (I26400,I26450);
OUT_INSTANCE I_1553 (I26403,I26460);
OUT_INSTANCE I_1554 (I26406,I26470);
OUT_INSTANCE I_1555 (I26409,I26480);
OUT_INSTANCE I_1556 (I26412,I26490);
OUT_INSTANCE I_1557 (I26415,I26500);
OUT_INSTANCE I_1558 (I26418,I26510);
OUT_INSTANCE I_1559 (I26421,I26520);
OUT_INSTANCE I_1560 (I26424,I26530);
PAT_1 I_1561 (I26490,I26450,I26510,I26440,I26460,I26440,I26470,I26520,I26500,I26530,I26480,I26570,I26573,I26576,I26579,I26582,I26585,I26588,I26591,I26594,I1892,I1899);
OUT_INSTANCE I_1562 (I26570,I26610);
OUT_INSTANCE I_1563 (I26573,I26620);
OUT_INSTANCE I_1564 (I26576,I26630);
OUT_INSTANCE I_1565 (I26579,I26640);
OUT_INSTANCE I_1566 (I26582,I26650);
OUT_INSTANCE I_1567 (I26585,I26660);
OUT_INSTANCE I_1568 (I26588,I26670);
OUT_INSTANCE I_1569 (I26591,I26680);
OUT_INSTANCE I_1570 (I26594,I26690);
PAT_12 I_1571 (I26650,I26630,I26690,I26610,I26640,I26610,I26620,I26680,I26660,I26620,I26670,I26730,I26733,I26736,I26739,I26742,I26745,I26748,I26751,I1892,I1899);
OUT_INSTANCE I_1572 (I26730,I26767);
OUT_INSTANCE I_1573 (I26733,I26777);
OUT_INSTANCE I_1574 (I26736,I26787);
OUT_INSTANCE I_1575 (I26739,I26797);
OUT_INSTANCE I_1576 (I26742,I26807);
OUT_INSTANCE I_1577 (I26745,I26817);
OUT_INSTANCE I_1578 (I26748,I26827);
OUT_INSTANCE I_1579 (I26751,I26837);
PAT_10 I_1580 (I26767,I26837,I26807,I26817,I26787,I26777,I26767,I26827,I26787,I26797,I26777,I26877,I26880,I26883,I26886,I26889,I26892,I26895,I26898,I1892,I1899);
OUT_INSTANCE I_1581 (I26877,I26914);
OUT_INSTANCE I_1582 (I26880,I26924);
OUT_INSTANCE I_1583 (I26883,I26934);
OUT_INSTANCE I_1584 (I26886,I26944);
OUT_INSTANCE I_1585 (I26889,I26954);
OUT_INSTANCE I_1586 (I26892,I26964);
OUT_INSTANCE I_1587 (I26895,I26974);
OUT_INSTANCE I_1588 (I26898,I26984);
PAT_9 I_1589 (I26954,I26914,I26924,I26934,I26914,I26934,I26944,I26924,I26984,I26964,I26974,I27024,I27027,I27030,I27033,I27036,I27039,I27042,I27045,I27048,I1892,I1899);
OUT_INSTANCE I_1590 (I27024,I27064);
OUT_INSTANCE I_1591 (I27027,I27074);
OUT_INSTANCE I_1592 (I27030,I27084);
OUT_INSTANCE I_1593 (I27033,I27094);
OUT_INSTANCE I_1594 (I27036,I27104);
OUT_INSTANCE I_1595 (I27039,I27114);
OUT_INSTANCE I_1596 (I27042,I27124);
OUT_INSTANCE I_1597 (I27045,I27134);
OUT_INSTANCE I_1598 (I27048,I27144);
PAT_6 I_1599 (I27124,I27064,I27104,I27134,I27064,I27094,I27084,I27144,I27114,I27074,I27074,I27184,I27187,I27190,I27193,I27196,I27199,I27202,I27205,I27208,I27211,I1892,I1899);
OUT_INSTANCE I_1600 (I27184,I27227);
OUT_INSTANCE I_1601 (I27187,I27237);
OUT_INSTANCE I_1602 (I27190,I27247);
OUT_INSTANCE I_1603 (I27193,I27257);
OUT_INSTANCE I_1604 (I27196,I27267);
OUT_INSTANCE I_1605 (I27199,I27277);
OUT_INSTANCE I_1606 (I27202,I27287);
OUT_INSTANCE I_1607 (I27205,I27297);
OUT_INSTANCE I_1608 (I27208,I27307);
OUT_INSTANCE I_1609 (I27211,I27317);
PAT_9 I_1610 (I27227,I27317,I27307,I27247,I27267,I27237,I27277,I27227,I27287,I27257,I27297,I27357,I27360,I27363,I27366,I27369,I27372,I27375,I27378,I27381,I1892,I1899);
OUT_INSTANCE I_1611 (I27357,I27397);
OUT_INSTANCE I_1612 (I27360,I27407);
OUT_INSTANCE I_1613 (I27363,I27417);
OUT_INSTANCE I_1614 (I27366,I27427);
OUT_INSTANCE I_1615 (I27369,I27437);
OUT_INSTANCE I_1616 (I27372,I27447);
OUT_INSTANCE I_1617 (I27375,I27457);
OUT_INSTANCE I_1618 (I27378,I27467);
OUT_INSTANCE I_1619 (I27381,I27477);
PAT_0 I_1620 (I27427,I27467,I27397,I27407,I27417,I27397,I27447,I27457,I27437,I27477,I27407,I27517,I27520,I27523,I27526,I27529,I27532,I27535,I27538,I1892,I1899);
OUT_INSTANCE I_1621 (I27517,I27554);
OUT_INSTANCE I_1622 (I27520,I27564);
OUT_INSTANCE I_1623 (I27523,I27574);
OUT_INSTANCE I_1624 (I27526,I27584);
OUT_INSTANCE I_1625 (I27529,I27594);
OUT_INSTANCE I_1626 (I27532,I27604);
OUT_INSTANCE I_1627 (I27535,I27614);
OUT_INSTANCE I_1628 (I27538,I27624);
PAT_9 I_1629 (I27574,I27614,I27564,I27594,I27604,I27564,I27554,I27584,I27624,I27574,I27554,I27664,I27667,I27670,I27673,I27676,I27679,I27682,I27685,I27688,I1892,I1899);
OUT_INSTANCE I_1630 (I27664,I27704);
OUT_INSTANCE I_1631 (I27667,I27714);
OUT_INSTANCE I_1632 (I27670,I27724);
OUT_INSTANCE I_1633 (I27673,I27734);
OUT_INSTANCE I_1634 (I27676,I27744);
OUT_INSTANCE I_1635 (I27679,I27754);
OUT_INSTANCE I_1636 (I27682,I27764);
OUT_INSTANCE I_1637 (I27685,I27774);
OUT_INSTANCE I_1638 (I27688,I27784);
PAT_10 I_1639 (I27774,I27764,I27724,I27714,I27784,I27734,I27754,I27714,I27704,I27704,I27744,I27824,I27827,I27830,I27833,I27836,I27839,I27842,I27845,I1892,I1899);
OUT_INSTANCE I_1640 (I27824,I27861);
OUT_INSTANCE I_1641 (I27827,I27871);
OUT_INSTANCE I_1642 (I27830,I27881);
OUT_INSTANCE I_1643 (I27833,I27891);
OUT_INSTANCE I_1644 (I27836,I27901);
OUT_INSTANCE I_1645 (I27839,I27911);
OUT_INSTANCE I_1646 (I27842,I27921);
OUT_INSTANCE I_1647 (I27845,I27931);
PAT_15 I_1648 (I27911,I27921,I27881,I27901,I27861,I27861,I27881,I27931,I27891,I27871,I27871,I27971,I27974,I27977,I27980,I27983,I27986,I27989,I27992,I27995,I1892,I1899);
OUT_INSTANCE I_1649 (I27971,I28011);
OUT_INSTANCE I_1650 (I27974,I28021);
OUT_INSTANCE I_1651 (I27977,I28031);
OUT_INSTANCE I_1652 (I27980,I28041);
OUT_INSTANCE I_1653 (I27983,I28051);
OUT_INSTANCE I_1654 (I27986,I28061);
OUT_INSTANCE I_1655 (I27989,I28071);
OUT_INSTANCE I_1656 (I27992,I28081);
OUT_INSTANCE I_1657 (I27995,I28091);
PAT_2 I_1658 (I28021,I28021,I28031,I28051,I28011,I28011,I28041,I28091,I28071,I28081,I28061,I28131,I28134,I28137,I28140,I28143,I28146,I28149,I28152,I28155,I1892,I1899);
OUT_INSTANCE I_1659 (I28131,I28171);
OUT_INSTANCE I_1660 (I28134,I28181);
OUT_INSTANCE I_1661 (I28137,I28191);
OUT_INSTANCE I_1662 (I28140,I28201);
OUT_INSTANCE I_1663 (I28143,I28211);
OUT_INSTANCE I_1664 (I28146,I28221);
OUT_INSTANCE I_1665 (I28149,I28231);
OUT_INSTANCE I_1666 (I28152,I28241);
OUT_INSTANCE I_1667 (I28155,I28251);
PAT_5 I_1668 (I28241,I28171,I28171,I28211,I28201,I28231,I28191,I28221,I28251,I28181,I28181,I28291,I28294,I28297,I28300,I28303,I28306,I28309,I28312,I28315,I28318,I1892,I1899);
OUT_INSTANCE I_1669 (I28291,I28334);
OUT_INSTANCE I_1670 (I28294,I28344);
OUT_INSTANCE I_1671 (I28297,I28354);
OUT_INSTANCE I_1672 (I28300,I28364);
OUT_INSTANCE I_1673 (I28303,I28374);
OUT_INSTANCE I_1674 (I28306,I28384);
OUT_INSTANCE I_1675 (I28309,I28394);
OUT_INSTANCE I_1676 (I28312,I28404);
OUT_INSTANCE I_1677 (I28315,I28414);
OUT_INSTANCE I_1678 (I28318,I28424);
PAT_0 I_1679 (I28404,I28334,I28424,I28414,I28334,I28394,I28374,I28344,I28364,I28384,I28354,I28464,I28467,I28470,I28473,I28476,I28479,I28482,I28485,I1892,I1899);
OUT_INSTANCE I_1680 (I28464,I28501);
OUT_INSTANCE I_1681 (I28467,I28511);
OUT_INSTANCE I_1682 (I28470,I28521);
OUT_INSTANCE I_1683 (I28473,I28531);
OUT_INSTANCE I_1684 (I28476,I28541);
OUT_INSTANCE I_1685 (I28479,I28551);
OUT_INSTANCE I_1686 (I28482,I28561);
OUT_INSTANCE I_1687 (I28485,I28571);
PAT_5 I_1688 (I28571,I28511,I28561,I28501,I28511,I28521,I28541,I28521,I28531,I28551,I28501,I28611,I28614,I28617,I28620,I28623,I28626,I28629,I28632,I28635,I28638,I1892,I1899);
OUT_INSTANCE I_1689 (I28611,I28654);
OUT_INSTANCE I_1690 (I28614,I28664);
OUT_INSTANCE I_1691 (I28617,I28674);
OUT_INSTANCE I_1692 (I28620,I28684);
OUT_INSTANCE I_1693 (I28623,I28694);
OUT_INSTANCE I_1694 (I28626,I28704);
OUT_INSTANCE I_1695 (I28629,I28714);
OUT_INSTANCE I_1696 (I28632,I28724);
OUT_INSTANCE I_1697 (I28635,I28734);
OUT_INSTANCE I_1698 (I28638,I28744);
PAT_10 I_1699 (I28734,I28744,I28674,I28694,I28704,I28724,I28664,I28654,I28654,I28684,I28714,I28784,I28787,I28790,I28793,I28796,I28799,I28802,I28805,I1892,I1899);
OUT_INSTANCE I_1700 (I28784,I28821);
OUT_INSTANCE I_1701 (I28787,I28831);
OUT_INSTANCE I_1702 (I28790,I28841);
OUT_INSTANCE I_1703 (I28793,I28851);
OUT_INSTANCE I_1704 (I28796,I28861);
OUT_INSTANCE I_1705 (I28799,I28871);
OUT_INSTANCE I_1706 (I28802,I28881);
OUT_INSTANCE I_1707 (I28805,I28891);
PAT_15 I_1708 (I28871,I28881,I28841,I28861,I28821,I28821,I28841,I28891,I28851,I28831,I28831,I28931,I28934,I28937,I28940,I28943,I28946,I28949,I28952,I28955,I1892,I1899);
OUT_INSTANCE I_1709 (I28931,I28971);
OUT_INSTANCE I_1710 (I28934,I28981);
OUT_INSTANCE I_1711 (I28937,I28991);
OUT_INSTANCE I_1712 (I28940,I29001);
OUT_INSTANCE I_1713 (I28943,I29011);
OUT_INSTANCE I_1714 (I28946,I29021);
OUT_INSTANCE I_1715 (I28949,I29031);
OUT_INSTANCE I_1716 (I28952,I29041);
OUT_INSTANCE I_1717 (I28955,I29051);
PAT_5 I_1718 (I28981,I28971,I28991,I29051,I29041,I29001,I29031,I29011,I28981,I29021,I28971,I29091,I29094,I29097,I29100,I29103,I29106,I29109,I29112,I29115,I29118,I1892,I1899);
OUT_INSTANCE I_1719 (I29091,I29134);
OUT_INSTANCE I_1720 (I29094,I29144);
OUT_INSTANCE I_1721 (I29097,I29154);
OUT_INSTANCE I_1722 (I29100,I29164);
OUT_INSTANCE I_1723 (I29103,I29174);
OUT_INSTANCE I_1724 (I29106,I29184);
OUT_INSTANCE I_1725 (I29109,I29194);
OUT_INSTANCE I_1726 (I29112,I29204);
OUT_INSTANCE I_1727 (I29115,I29214);
OUT_INSTANCE I_1728 (I29118,I29224);
PAT_2 I_1729 (I29184,I29134,I29174,I29154,I29204,I29144,I29194,I29164,I29214,I29224,I29134,I29264,I29267,I29270,I29273,I29276,I29279,I29282,I29285,I29288,I1892,I1899);
OUT_INSTANCE I_1730 (I29264,I29304);
OUT_INSTANCE I_1731 (I29267,I29314);
OUT_INSTANCE I_1732 (I29270,I29324);
OUT_INSTANCE I_1733 (I29273,I29334);
OUT_INSTANCE I_1734 (I29276,I29344);
OUT_INSTANCE I_1735 (I29279,I29354);
OUT_INSTANCE I_1736 (I29282,I29364);
OUT_INSTANCE I_1737 (I29285,I29374);
OUT_INSTANCE I_1738 (I29288,I29384);
PAT_5 I_1739 (I29374,I29304,I29304,I29344,I29334,I29364,I29324,I29354,I29384,I29314,I29314,I29424,I29427,I29430,I29433,I29436,I29439,I29442,I29445,I29448,I29451,I1892,I1899);
OUT_INSTANCE I_1740 (I29424,I29467);
OUT_INSTANCE I_1741 (I29427,I29477);
OUT_INSTANCE I_1742 (I29430,I29487);
OUT_INSTANCE I_1743 (I29433,I29497);
OUT_INSTANCE I_1744 (I29436,I29507);
OUT_INSTANCE I_1745 (I29439,I29517);
OUT_INSTANCE I_1746 (I29442,I29527);
OUT_INSTANCE I_1747 (I29445,I29537);
OUT_INSTANCE I_1748 (I29448,I29547);
OUT_INSTANCE I_1749 (I29451,I29557);
PAT_6 I_1750 (I29527,I29507,I29467,I29487,I29477,I29497,I29517,I29467,I29547,I29537,I29557,I29597,I29600,I29603,I29606,I29609,I29612,I29615,I29618,I29621,I29624,I1892,I1899);
OUT_INSTANCE I_1751 (I29597,I29640);
OUT_INSTANCE I_1752 (I29600,I29650);
OUT_INSTANCE I_1753 (I29603,I29660);
OUT_INSTANCE I_1754 (I29606,I29670);
OUT_INSTANCE I_1755 (I29609,I29680);
OUT_INSTANCE I_1756 (I29612,I29690);
OUT_INSTANCE I_1757 (I29615,I29700);
OUT_INSTANCE I_1758 (I29618,I29710);
OUT_INSTANCE I_1759 (I29621,I29720);
OUT_INSTANCE I_1760 (I29624,I29730);
PAT_9 I_1761 (I29640,I29730,I29720,I29660,I29680,I29650,I29690,I29640,I29700,I29670,I29710,I29770,I29773,I29776,I29779,I29782,I29785,I29788,I29791,I29794,I1892,I1899);
OUT_INSTANCE I_1762 (I29770,I29810);
OUT_INSTANCE I_1763 (I29773,I29820);
OUT_INSTANCE I_1764 (I29776,I29830);
OUT_INSTANCE I_1765 (I29779,I29840);
OUT_INSTANCE I_1766 (I29782,I29850);
OUT_INSTANCE I_1767 (I29785,I29860);
OUT_INSTANCE I_1768 (I29788,I29870);
OUT_INSTANCE I_1769 (I29791,I29880);
OUT_INSTANCE I_1770 (I29794,I29890);
PAT_14 I_1771 (I29840,I29810,I29890,I29830,I29820,I29810,I29860,I29880,I29850,I29820,I29870,I29930,I29933,I29936,I29939,I29942,I29945,I29948,I29951,I29954,I1892,I1899);
OUT_INSTANCE I_1772 (I29930,I29970);
OUT_INSTANCE I_1773 (I29933,I29980);
OUT_INSTANCE I_1774 (I29936,I29990);
OUT_INSTANCE I_1775 (I29939,I30000);
OUT_INSTANCE I_1776 (I29942,I30010);
OUT_INSTANCE I_1777 (I29945,I30020);
OUT_INSTANCE I_1778 (I29948,I30030);
OUT_INSTANCE I_1779 (I29951,I30040);
OUT_INSTANCE I_1780 (I29954,I30050);
PAT_2 I_1781 (I30030,I30050,I30000,I29970,I29980,I29980,I30020,I29970,I30040,I29990,I30010,I30090,I30093,I30096,I30099,I30102,I30105,I30108,I30111,I30114,I1892,I1899);
OUT_INSTANCE I_1782 (I30090,I30130);
OUT_INSTANCE I_1783 (I30093,I30140);
OUT_INSTANCE I_1784 (I30096,I30150);
OUT_INSTANCE I_1785 (I30099,I30160);
OUT_INSTANCE I_1786 (I30102,I30170);
OUT_INSTANCE I_1787 (I30105,I30180);
OUT_INSTANCE I_1788 (I30108,I30190);
OUT_INSTANCE I_1789 (I30111,I30200);
OUT_INSTANCE I_1790 (I30114,I30210);
PAT_15 I_1791 (I30140,I30180,I30200,I30210,I30150,I30190,I30130,I30160,I30130,I30170,I30140,I30250,I30253,I30256,I30259,I30262,I30265,I30268,I30271,I30274,I1892,I1899);
OUT_INSTANCE I_1792 (I30250,I30290);
OUT_INSTANCE I_1793 (I30253,I30300);
OUT_INSTANCE I_1794 (I30256,I30310);
OUT_INSTANCE I_1795 (I30259,I30320);
OUT_INSTANCE I_1796 (I30262,I30330);
OUT_INSTANCE I_1797 (I30265,I30340);
OUT_INSTANCE I_1798 (I30268,I30350);
OUT_INSTANCE I_1799 (I30271,I30360);
OUT_INSTANCE I_1800 (I30274,I30370);
PAT_12 I_1801 (I30350,I30360,I30370,I30330,I30320,I30300,I30290,I30340,I30310,I30290,I30300,I30410,I30413,I30416,I30419,I30422,I30425,I30428,I30431,I1892,I1899);
OUT_INSTANCE I_1802 (I30410,I30447);
OUT_INSTANCE I_1803 (I30413,I30457);
OUT_INSTANCE I_1804 (I30416,I30467);
OUT_INSTANCE I_1805 (I30419,I30477);
OUT_INSTANCE I_1806 (I30422,I30487);
OUT_INSTANCE I_1807 (I30425,I30497);
OUT_INSTANCE I_1808 (I30428,I30507);
OUT_INSTANCE I_1809 (I30431,I30517);
PAT_17 I_1810 (I30497,I30477,I30457,I30447,I30447,I30467,I30467,I30507,I30517,I30457,I30487,I30557,I30560,I30563,I30566,I30569,I30572,I30575,I30578,I30581,I30584,I1892,I1899);
OUT_INSTANCE I_1811 (I30557,I30600);
OUT_INSTANCE I_1812 (I30560,I30610);
OUT_INSTANCE I_1813 (I30563,I30620);
OUT_INSTANCE I_1814 (I30566,I30630);
OUT_INSTANCE I_1815 (I30569,I30640);
OUT_INSTANCE I_1816 (I30572,I30650);
OUT_INSTANCE I_1817 (I30575,I30660);
OUT_INSTANCE I_1818 (I30578,I30670);
OUT_INSTANCE I_1819 (I30581,I30680);
OUT_INSTANCE I_1820 (I30584,I30690);
PAT_12 I_1821 (I30680,I30620,I30600,I30660,I30640,I30670,I30610,I30690,I30600,I30630,I30650,I30730,I30733,I30736,I30739,I30742,I30745,I30748,I30751,I1892,I1899);
OUT_INSTANCE I_1822 (I30730,I30767);
OUT_INSTANCE I_1823 (I30733,I30777);
OUT_INSTANCE I_1824 (I30736,I30787);
OUT_INSTANCE I_1825 (I30739,I30797);
OUT_INSTANCE I_1826 (I30742,I30807);
OUT_INSTANCE I_1827 (I30745,I30817);
OUT_INSTANCE I_1828 (I30748,I30827);
OUT_INSTANCE I_1829 (I30751,I30837);
PAT_7 I_1830 (I30787,I30797,I30767,I30807,I30827,I30787,I30837,I30817,I30777,I30777,I30767,I30877,I30880,I30883,I30886,I30889,I30892,I30895,I30898,I30901,I1892,I1899);
OUT_INSTANCE I_1831 (I30877,I30917);
OUT_INSTANCE I_1832 (I30880,I30927);
OUT_INSTANCE I_1833 (I30883,I30937);
OUT_INSTANCE I_1834 (I30886,I30947);
OUT_INSTANCE I_1835 (I30889,I30957);
OUT_INSTANCE I_1836 (I30892,I30967);
OUT_INSTANCE I_1837 (I30895,I30977);
OUT_INSTANCE I_1838 (I30898,I30987);
OUT_INSTANCE I_1839 (I30901,I30997);
PAT_4 I_1840 (I30997,I30917,I30917,I30967,I30947,I30927,I30927,I30977,I30987,I30937,I30957,I31037,I31040,I31043,I31046,I31049,I31052,I31055,I31058,I31061,I1892,I1899);
OUT_INSTANCE I_1841 (I31037,I31077);
OUT_INSTANCE I_1842 (I31040,I31087);
OUT_INSTANCE I_1843 (I31043,I31097);
OUT_INSTANCE I_1844 (I31046,I31107);
OUT_INSTANCE I_1845 (I31049,I31117);
OUT_INSTANCE I_1846 (I31052,I31127);
OUT_INSTANCE I_1847 (I31055,I31137);
OUT_INSTANCE I_1848 (I31058,I31147);
OUT_INSTANCE I_1849 (I31061,I31157);
PAT_6 I_1850 (I31077,I31097,I31087,I31127,I31137,I31117,I31157,I31147,I31077,I31107,I31087,I31197,I31200,I31203,I31206,I31209,I31212,I31215,I31218,I31221,I31224,I1892,I1899);
OUT_INSTANCE I_1851 (I31197,I31240);
OUT_INSTANCE I_1852 (I31200,I31250);
OUT_INSTANCE I_1853 (I31203,I31260);
OUT_INSTANCE I_1854 (I31206,I31270);
OUT_INSTANCE I_1855 (I31209,I31280);
OUT_INSTANCE I_1856 (I31212,I31290);
OUT_INSTANCE I_1857 (I31215,I31300);
OUT_INSTANCE I_1858 (I31218,I31310);
OUT_INSTANCE I_1859 (I31221,I31320);
OUT_INSTANCE I_1860 (I31224,I31330);
PAT_1 I_1861 (I31330,I31300,I31260,I31270,I31310,I31280,I31290,I31240,I31250,I31240,I31320,I31370,I31373,I31376,I31379,I31382,I31385,I31388,I31391,I31394,I1892,I1899);
OUT_INSTANCE I_1862 (I31370,I31410);
OUT_INSTANCE I_1863 (I31373,I31420);
OUT_INSTANCE I_1864 (I31376,I31430);
OUT_INSTANCE I_1865 (I31379,I31440);
OUT_INSTANCE I_1866 (I31382,I31450);
OUT_INSTANCE I_1867 (I31385,I31460);
OUT_INSTANCE I_1868 (I31388,I31470);
OUT_INSTANCE I_1869 (I31391,I31480);
OUT_INSTANCE I_1870 (I31394,I31490);
PAT_2 I_1871 (I31410,I31430,I31410,I31460,I31420,I31420,I31440,I31450,I31470,I31490,I31480,I31530,I31533,I31536,I31539,I31542,I31545,I31548,I31551,I31554,I1892,I1899);
OUT_INSTANCE I_1872 (I31530,I31570);
OUT_INSTANCE I_1873 (I31533,I31580);
OUT_INSTANCE I_1874 (I31536,I31590);
OUT_INSTANCE I_1875 (I31539,I31600);
OUT_INSTANCE I_1876 (I31542,I31610);
OUT_INSTANCE I_1877 (I31545,I31620);
OUT_INSTANCE I_1878 (I31548,I31630);
OUT_INSTANCE I_1879 (I31551,I31640);
OUT_INSTANCE I_1880 (I31554,I31650);
PAT_9 I_1881 (I31620,I31650,I31570,I31590,I31600,I31630,I31580,I31610,I31640,I31580,I31570,I31690,I31693,I31696,I31699,I31702,I31705,I31708,I31711,I31714,I1892,I1899);
OUT_INSTANCE I_1882 (I31690,I31730);
OUT_INSTANCE I_1883 (I31693,I31740);
OUT_INSTANCE I_1884 (I31696,I31750);
OUT_INSTANCE I_1885 (I31699,I31760);
OUT_INSTANCE I_1886 (I31702,I31770);
OUT_INSTANCE I_1887 (I31705,I31780);
OUT_INSTANCE I_1888 (I31708,I31790);
OUT_INSTANCE I_1889 (I31711,I31800);
OUT_INSTANCE I_1890 (I31714,I31810);
PAT_4 I_1891 (I31730,I31810,I31790,I31750,I31740,I31800,I31740,I31730,I31780,I31760,I31770,I31850,I31853,I31856,I31859,I31862,I31865,I31868,I31871,I31874,I1892,I1899);
OUT_INSTANCE I_1892 (I31850,I31890);
OUT_INSTANCE I_1893 (I31853,I31900);
OUT_INSTANCE I_1894 (I31856,I31910);
OUT_INSTANCE I_1895 (I31859,I31920);
OUT_INSTANCE I_1896 (I31862,I31930);
OUT_INSTANCE I_1897 (I31865,I31940);
OUT_INSTANCE I_1898 (I31868,I31950);
OUT_INSTANCE I_1899 (I31871,I31960);
OUT_INSTANCE I_1900 (I31874,I31970);
PAT_12 I_1901 (I31890,I31900,I31960,I31970,I31940,I31910,I31930,I31920,I31890,I31950,I31900,I32010,I32013,I32016,I32019,I32022,I32025,I32028,I32031,I1892,I1899);
OUT_INSTANCE I_1902 (I32010,I32047);
OUT_INSTANCE I_1903 (I32013,I32057);
OUT_INSTANCE I_1904 (I32016,I32067);
OUT_INSTANCE I_1905 (I32019,I32077);
OUT_INSTANCE I_1906 (I32022,I32087);
OUT_INSTANCE I_1907 (I32025,I32097);
OUT_INSTANCE I_1908 (I32028,I32107);
OUT_INSTANCE I_1909 (I32031,I32117);
PAT_5 I_1910 (I32077,I32097,I32117,I32067,I32067,I32047,I32107,I32047,I32057,I32057,I32087,I32157,I32160,I32163,I32166,I32169,I32172,I32175,I32178,I32181,I32184,I1892,I1899);
OUT_INSTANCE I_1911 (I32157,I32200);
OUT_INSTANCE I_1912 (I32160,I32210);
OUT_INSTANCE I_1913 (I32163,I32220);
OUT_INSTANCE I_1914 (I32166,I32230);
OUT_INSTANCE I_1915 (I32169,I32240);
OUT_INSTANCE I_1916 (I32172,I32250);
OUT_INSTANCE I_1917 (I32175,I32260);
OUT_INSTANCE I_1918 (I32178,I32270);
OUT_INSTANCE I_1919 (I32181,I32280);
OUT_INSTANCE I_1920 (I32184,I32290);
PAT_17 I_1921 (I32290,I32210,I32220,I32230,I32200,I32240,I32200,I32280,I32260,I32250,I32270,I32330,I32333,I32336,I32339,I32342,I32345,I32348,I32351,I32354,I32357,I1892,I1899);
OUT_INSTANCE I_1922 (I32330,I32373);
OUT_INSTANCE I_1923 (I32333,I32383);
OUT_INSTANCE I_1924 (I32336,I32393);
OUT_INSTANCE I_1925 (I32339,I32403);
OUT_INSTANCE I_1926 (I32342,I32413);
OUT_INSTANCE I_1927 (I32345,I32423);
OUT_INSTANCE I_1928 (I32348,I32433);
OUT_INSTANCE I_1929 (I32351,I32443);
OUT_INSTANCE I_1930 (I32354,I32453);
OUT_INSTANCE I_1931 (I32357,I32463);
PAT_7 I_1932 (I32433,I32403,I32423,I32383,I32413,I32443,I32463,I32373,I32453,I32393,I32373,I32503,I32506,I32509,I32512,I32515,I32518,I32521,I32524,I32527,I1892,I1899);
OUT_INSTANCE I_1933 (I32503,I32543);
OUT_INSTANCE I_1934 (I32506,I32553);
OUT_INSTANCE I_1935 (I32509,I32563);
OUT_INSTANCE I_1936 (I32512,I32573);
OUT_INSTANCE I_1937 (I32515,I32583);
OUT_INSTANCE I_1938 (I32518,I32593);
OUT_INSTANCE I_1939 (I32521,I32603);
OUT_INSTANCE I_1940 (I32524,I32613);
OUT_INSTANCE I_1941 (I32527,I32623);
PAT_4 I_1942 (I32623,I32543,I32543,I32593,I32573,I32553,I32553,I32603,I32613,I32563,I32583,I32663,I32666,I32669,I32672,I32675,I32678,I32681,I32684,I32687,I1892,I1899);
OUT_INSTANCE I_1943 (I32663,I32703);
OUT_INSTANCE I_1944 (I32666,I32713);
OUT_INSTANCE I_1945 (I32669,I32723);
OUT_INSTANCE I_1946 (I32672,I32733);
OUT_INSTANCE I_1947 (I32675,I32743);
OUT_INSTANCE I_1948 (I32678,I32753);
OUT_INSTANCE I_1949 (I32681,I32763);
OUT_INSTANCE I_1950 (I32684,I32773);
OUT_INSTANCE I_1951 (I32687,I32783);
PAT_8 I_1952 (I32743,I32703,I32773,I32723,I32713,I32783,I32733,I32763,I32713,I32703,I32753,I32823,I32826,I32829,I32832,I32835,I32838,I32841,I32844,I32847,I1892,I1899);
OUT_INSTANCE I_1953 (I32823,I32863);
OUT_INSTANCE I_1954 (I32826,I32873);
OUT_INSTANCE I_1955 (I32829,I32883);
OUT_INSTANCE I_1956 (I32832,I32893);
OUT_INSTANCE I_1957 (I32835,I32903);
OUT_INSTANCE I_1958 (I32838,I32913);
OUT_INSTANCE I_1959 (I32841,I32923);
OUT_INSTANCE I_1960 (I32844,I32933);
OUT_INSTANCE I_1961 (I32847,I32943);
PAT_5 I_1962 (I32883,I32943,I32863,I32933,I32893,I32903,I32873,I32863,I32873,I32913,I32923,I32983,I32986,I32989,I32992,I32995,I32998,I33001,I33004,I33007,I33010,I1892,I1899);
OUT_INSTANCE I_1963 (I32983,I33026);
OUT_INSTANCE I_1964 (I32986,I33036);
OUT_INSTANCE I_1965 (I32989,I33046);
OUT_INSTANCE I_1966 (I32992,I33056);
OUT_INSTANCE I_1967 (I32995,I33066);
OUT_INSTANCE I_1968 (I32998,I33076);
OUT_INSTANCE I_1969 (I33001,I33086);
OUT_INSTANCE I_1970 (I33004,I33096);
OUT_INSTANCE I_1971 (I33007,I33106);
OUT_INSTANCE I_1972 (I33010,I33116);
PAT_6 I_1973 (I33086,I33066,I33026,I33046,I33036,I33056,I33076,I33026,I33106,I33096,I33116,I33156,I33159,I33162,I33165,I33168,I33171,I33174,I33177,I33180,I33183,I1892,I1899);
OUT_INSTANCE I_1974 (I33156,I33199);
OUT_INSTANCE I_1975 (I33159,I33209);
OUT_INSTANCE I_1976 (I33162,I33219);
OUT_INSTANCE I_1977 (I33165,I33229);
OUT_INSTANCE I_1978 (I33168,I33239);
OUT_INSTANCE I_1979 (I33171,I33249);
OUT_INSTANCE I_1980 (I33174,I33259);
OUT_INSTANCE I_1981 (I33177,I33269);
OUT_INSTANCE I_1982 (I33180,I33279);
OUT_INSTANCE I_1983 (I33183,I33289);
PAT_8 I_1984 (I33229,I33249,I33219,I33259,I33199,I33209,I33269,I33199,I33289,I33279,I33239,I33329,I33332,I33335,I33338,I33341,I33344,I33347,I33350,I33353,I1892,I1899);
OUT_INSTANCE I_1985 (I33329,I33369);
OUT_INSTANCE I_1986 (I33332,I33379);
OUT_INSTANCE I_1987 (I33335,I33389);
OUT_INSTANCE I_1988 (I33338,I33399);
OUT_INSTANCE I_1989 (I33341,I33409);
OUT_INSTANCE I_1990 (I33344,I33419);
OUT_INSTANCE I_1991 (I33347,I33429);
OUT_INSTANCE I_1992 (I33350,I33439);
OUT_INSTANCE I_1993 (I33353,I33449);
PAT_13 I_1994 (I33409,I33439,I33379,I33449,I33389,I33369,I33369,I33399,I33429,I33419,I33379,I33489,I33492,I33495,I33498,I33501,I33504,I33507,I33510,I33513,I1892,I1899);
OUT_INSTANCE I_1995 (I33489,I33529);
OUT_INSTANCE I_1996 (I33492,I33539);
OUT_INSTANCE I_1997 (I33495,I33549);
OUT_INSTANCE I_1998 (I33498,I33559);
OUT_INSTANCE I_1999 (I33501,I33569);
OUT_INSTANCE I_2000 (I33504,I33579);
OUT_INSTANCE I_2001 (I33507,I33589);
OUT_INSTANCE I_2002 (I33510,I33599);
OUT_INSTANCE I_2003 (I33513,I33609);
PAT_17 I_2004 (I33609,I33569,I33599,I33589,I33559,I33529,I33539,I33549,I33529,I33579,I33539,I33649,I33652,I33655,I33658,I33661,I33664,I33667,I33670,I33673,I33676,I1892,I1899);
OUT_INSTANCE I_2005 (I33649,I33692);
OUT_INSTANCE I_2006 (I33652,I33702);
OUT_INSTANCE I_2007 (I33655,I33712);
OUT_INSTANCE I_2008 (I33658,I33722);
OUT_INSTANCE I_2009 (I33661,I33732);
OUT_INSTANCE I_2010 (I33664,I33742);
OUT_INSTANCE I_2011 (I33667,I33752);
OUT_INSTANCE I_2012 (I33670,I33762);
OUT_INSTANCE I_2013 (I33673,I33772);
OUT_INSTANCE I_2014 (I33676,I33782);
PAT_9 I_2015 (I33762,I33702,I33722,I33772,I33712,I33752,I33692,I33732,I33692,I33782,I33742,I33822,I33825,I33828,I33831,I33834,I33837,I33840,I33843,I33846,I1892,I1899);
OUT_INSTANCE I_2016 (I33822,I33862);
OUT_INSTANCE I_2017 (I33825,I33872);
OUT_INSTANCE I_2018 (I33828,I33882);
OUT_INSTANCE I_2019 (I33831,I33892);
OUT_INSTANCE I_2020 (I33834,I33902);
OUT_INSTANCE I_2021 (I33837,I33912);
OUT_INSTANCE I_2022 (I33840,I33922);
OUT_INSTANCE I_2023 (I33843,I33932);
OUT_INSTANCE I_2024 (I33846,I33942);
PAT_2 I_2025 (I33912,I33922,I33892,I33942,I33862,I33872,I33882,I33872,I33932,I33902,I33862,I33982,I33985,I33988,I33991,I33994,I33997,I34000,I34003,I34006,I1892,I1899);
OUT_INSTANCE I_2026 (I33982,I34022);
OUT_INSTANCE I_2027 (I33985,I34032);
OUT_INSTANCE I_2028 (I33988,I34042);
OUT_INSTANCE I_2029 (I33991,I34052);
OUT_INSTANCE I_2030 (I33994,I34062);
OUT_INSTANCE I_2031 (I33997,I34072);
OUT_INSTANCE I_2032 (I34000,I34082);
OUT_INSTANCE I_2033 (I34003,I34092);
OUT_INSTANCE I_2034 (I34006,I34102);
IN_INSTANCE I_2035 (I1429,I34112);
IN_INSTANCE I_2036 (I1685,I34122);
IN_INSTANCE I_2037 (I1733,I34132);
IN_INSTANCE I_2038 (I1837,I34142);
IN_INSTANCE I_2039 (I1701,I34152);
IN_INSTANCE I_2040 (I1829,I34162);
IN_INSTANCE I_2041 (I1501,I34172);
IN_INSTANCE I_2042 (I1709,I34182);
IN_INSTANCE I_2043 (I1741,I34192);
IN_INSTANCE I_2044 (I1405,I34202);
IN_INSTANCE I_2045 (I1693,I34212);
PAT_5 I_2046 (I34112,I34122,I34132,I34142,I34152,I34162,I34172,I34182,I34192,I34202,I34212,I34252,I34255,I34258,I34261,I34264,I34267,I34270,I34273,I34276,I34279,I1892,I1899);
OUT_INSTANCE I_2047 (I34252,I34295);
OUT_INSTANCE I_2048 (I34255,I34305);
OUT_INSTANCE I_2049 (I34258,I34315);
OUT_INSTANCE I_2050 (I34261,I34325);
OUT_INSTANCE I_2051 (I34264,I34335);
OUT_INSTANCE I_2052 (I34267,I34345);
OUT_INSTANCE I_2053 (I34270,I34355);
OUT_INSTANCE I_2054 (I34273,I34365);
OUT_INSTANCE I_2055 (I34276,I34375);
OUT_INSTANCE I_2056 (I34279,I34385);
PAT_4 I_2057 (I34355,I34375,I34385,I34315,I34325,I34365,I34305,I34295,I34335,I34345,I34295,I34425,I34428,I34431,I34434,I34437,I34440,I34443,I34446,I34449,I1892,I1899);
OUT_INSTANCE I_2058 (I34425,I34465);
OUT_INSTANCE I_2059 (I34428,I34475);
OUT_INSTANCE I_2060 (I34431,I34485);
OUT_INSTANCE I_2061 (I34434,I34495);
OUT_INSTANCE I_2062 (I34437,I34505);
OUT_INSTANCE I_2063 (I34440,I34515);
OUT_INSTANCE I_2064 (I34443,I34525);
OUT_INSTANCE I_2065 (I34446,I34535);
OUT_INSTANCE I_2066 (I34449,I34545);
PAT_9 I_2067 (I34535,I34475,I34485,I34515,I34525,I34465,I34495,I34475,I34545,I34465,I34505,I34585,I34588,I34591,I34594,I34597,I34600,I34603,I34606,I34609,I1892,I1899);
OUT_INSTANCE I_2068 (I34585,I34625);
OUT_INSTANCE I_2069 (I34588,I34635);
OUT_INSTANCE I_2070 (I34591,I34645);
OUT_INSTANCE I_2071 (I34594,I34655);
OUT_INSTANCE I_2072 (I34597,I34665);
OUT_INSTANCE I_2073 (I34600,I34675);
OUT_INSTANCE I_2074 (I34603,I34685);
OUT_INSTANCE I_2075 (I34606,I34695);
OUT_INSTANCE I_2076 (I34609,I34705);
PAT_2 I_2077 (I34675,I34685,I34655,I34705,I34625,I34635,I34645,I34635,I34695,I34665,I34625,I34745,I34748,I34751,I34754,I34757,I34760,I34763,I34766,I34769,I1892,I1899);
OUT_INSTANCE I_2078 (I34745,I34785);
OUT_INSTANCE I_2079 (I34748,I34795);
OUT_INSTANCE I_2080 (I34751,I34805);
OUT_INSTANCE I_2081 (I34754,I34815);
OUT_INSTANCE I_2082 (I34757,I34825);
OUT_INSTANCE I_2083 (I34760,I34835);
OUT_INSTANCE I_2084 (I34763,I34845);
OUT_INSTANCE I_2085 (I34766,I34855);
OUT_INSTANCE I_2086 (I34769,I34865);
PAT_9 I_2087 (I34835,I34865,I34785,I34805,I34815,I34845,I34795,I34825,I34855,I34795,I34785,I34905,I34908,I34911,I34914,I34917,I34920,I34923,I34926,I34929,I1892,I1899);
OUT_INSTANCE I_2088 (I34905,I34945);
OUT_INSTANCE I_2089 (I34908,I34955);
OUT_INSTANCE I_2090 (I34911,I34965);
OUT_INSTANCE I_2091 (I34914,I34975);
OUT_INSTANCE I_2092 (I34917,I34985);
OUT_INSTANCE I_2093 (I34920,I34995);
OUT_INSTANCE I_2094 (I34923,I35005);
OUT_INSTANCE I_2095 (I34926,I35015);
OUT_INSTANCE I_2096 (I34929,I35025);
PAT_8 I_2097 (I35015,I34975,I35005,I34945,I34955,I34995,I35025,I34955,I34965,I34985,I34945,I35065,I35068,I35071,I35074,I35077,I35080,I35083,I35086,I35089,I1892,I1899);
OUT_INSTANCE I_2098 (I35065,I35105);
OUT_INSTANCE I_2099 (I35068,I35115);
OUT_INSTANCE I_2100 (I35071,I35125);
OUT_INSTANCE I_2101 (I35074,I35135);
OUT_INSTANCE I_2102 (I35077,I35145);
OUT_INSTANCE I_2103 (I35080,I35155);
OUT_INSTANCE I_2104 (I35083,I35165);
OUT_INSTANCE I_2105 (I35086,I35175);
OUT_INSTANCE I_2106 (I35089,I35185);
PAT_9 I_2107 (I35115,I35145,I35115,I35105,I35155,I35125,I35175,I35135,I35165,I35105,I35185,I35225,I35228,I35231,I35234,I35237,I35240,I35243,I35246,I35249,I1892,I1899);
OUT_INSTANCE I_2108 (I35225,I35265);
OUT_INSTANCE I_2109 (I35228,I35275);
OUT_INSTANCE I_2110 (I35231,I35285);
OUT_INSTANCE I_2111 (I35234,I35295);
OUT_INSTANCE I_2112 (I35237,I35305);
OUT_INSTANCE I_2113 (I35240,I35315);
OUT_INSTANCE I_2114 (I35243,I35325);
OUT_INSTANCE I_2115 (I35246,I35335);
OUT_INSTANCE I_2116 (I35249,I35345);
PAT_0 I_2117 (I35295,I35335,I35265,I35275,I35285,I35265,I35315,I35325,I35305,I35345,I35275,I35385,I35388,I35391,I35394,I35397,I35400,I35403,I35406,I1892,I1899);
OUT_INSTANCE I_2118 (I35385,I35422);
OUT_INSTANCE I_2119 (I35388,I35432);
OUT_INSTANCE I_2120 (I35391,I35442);
OUT_INSTANCE I_2121 (I35394,I35452);
OUT_INSTANCE I_2122 (I35397,I35462);
OUT_INSTANCE I_2123 (I35400,I35472);
OUT_INSTANCE I_2124 (I35403,I35482);
OUT_INSTANCE I_2125 (I35406,I35492);
PAT_5 I_2126 (I35492,I35432,I35482,I35422,I35432,I35442,I35462,I35442,I35452,I35472,I35422,I35532,I35535,I35538,I35541,I35544,I35547,I35550,I35553,I35556,I35559,I1892,I1899);
OUT_INSTANCE I_2127 (I35532,I35575);
OUT_INSTANCE I_2128 (I35535,I35585);
OUT_INSTANCE I_2129 (I35538,I35595);
OUT_INSTANCE I_2130 (I35541,I35605);
OUT_INSTANCE I_2131 (I35544,I35615);
OUT_INSTANCE I_2132 (I35547,I35625);
OUT_INSTANCE I_2133 (I35550,I35635);
OUT_INSTANCE I_2134 (I35553,I35645);
OUT_INSTANCE I_2135 (I35556,I35655);
OUT_INSTANCE I_2136 (I35559,I35665);
PAT_9 I_2137 (I35625,I35615,I35645,I35635,I35605,I35575,I35595,I35665,I35585,I35655,I35575,I35705,I35708,I35711,I35714,I35717,I35720,I35723,I35726,I35729,I1892,I1899);
OUT_INSTANCE I_2138 (I35705,I35745);
OUT_INSTANCE I_2139 (I35708,I35755);
OUT_INSTANCE I_2140 (I35711,I35765);
OUT_INSTANCE I_2141 (I35714,I35775);
OUT_INSTANCE I_2142 (I35717,I35785);
OUT_INSTANCE I_2143 (I35720,I35795);
OUT_INSTANCE I_2144 (I35723,I35805);
OUT_INSTANCE I_2145 (I35726,I35815);
OUT_INSTANCE I_2146 (I35729,I35825);
PAT_5 I_2147 (I35815,I35745,I35795,I35745,I35765,I35775,I35755,I35755,I35805,I35785,I35825,I35865,I35868,I35871,I35874,I35877,I35880,I35883,I35886,I35889,I35892,I1892,I1899);
OUT_INSTANCE I_2148 (I35865,I35908);
OUT_INSTANCE I_2149 (I35868,I35918);
OUT_INSTANCE I_2150 (I35871,I35928);
OUT_INSTANCE I_2151 (I35874,I35938);
OUT_INSTANCE I_2152 (I35877,I35948);
OUT_INSTANCE I_2153 (I35880,I35958);
OUT_INSTANCE I_2154 (I35883,I35968);
OUT_INSTANCE I_2155 (I35886,I35978);
OUT_INSTANCE I_2156 (I35889,I35988);
OUT_INSTANCE I_2157 (I35892,I35998);
PAT_4 I_2158 (I35968,I35988,I35998,I35928,I35938,I35978,I35918,I35908,I35948,I35958,I35908,I36038,I36041,I36044,I36047,I36050,I36053,I36056,I36059,I36062,I1892,I1899);
OUT_INSTANCE I_2159 (I36038,I36078);
OUT_INSTANCE I_2160 (I36041,I36088);
OUT_INSTANCE I_2161 (I36044,I36098);
OUT_INSTANCE I_2162 (I36047,I36108);
OUT_INSTANCE I_2163 (I36050,I36118);
OUT_INSTANCE I_2164 (I36053,I36128);
OUT_INSTANCE I_2165 (I36056,I36138);
OUT_INSTANCE I_2166 (I36059,I36148);
OUT_INSTANCE I_2167 (I36062,I36158);
PAT_2 I_2168 (I36108,I36088,I36088,I36158,I36078,I36138,I36128,I36098,I36078,I36118,I36148,I36198,I36201,I36204,I36207,I36210,I36213,I36216,I36219,I36222,I1892,I1899);
OUT_INSTANCE I_2169 (I36198,I36238);
OUT_INSTANCE I_2170 (I36201,I36248);
OUT_INSTANCE I_2171 (I36204,I36258);
OUT_INSTANCE I_2172 (I36207,I36268);
OUT_INSTANCE I_2173 (I36210,I36278);
OUT_INSTANCE I_2174 (I36213,I36288);
OUT_INSTANCE I_2175 (I36216,I36298);
OUT_INSTANCE I_2176 (I36219,I36308);
OUT_INSTANCE I_2177 (I36222,I36318);
PAT_6 I_2178 (I36318,I36238,I36288,I36278,I36298,I36268,I36248,I36308,I36238,I36258,I36248,I36358,I36361,I36364,I36367,I36370,I36373,I36376,I36379,I36382,I36385,I1892,I1899);
OUT_INSTANCE I_2179 (I36358,I36401);
OUT_INSTANCE I_2180 (I36361,I36411);
OUT_INSTANCE I_2181 (I36364,I36421);
OUT_INSTANCE I_2182 (I36367,I36431);
OUT_INSTANCE I_2183 (I36370,I36441);
OUT_INSTANCE I_2184 (I36373,I36451);
OUT_INSTANCE I_2185 (I36376,I36461);
OUT_INSTANCE I_2186 (I36379,I36471);
OUT_INSTANCE I_2187 (I36382,I36481);
OUT_INSTANCE I_2188 (I36385,I36491);
PAT_15 I_2189 (I36461,I36431,I36471,I36481,I36451,I36491,I36401,I36421,I36401,I36411,I36441,I36531,I36534,I36537,I36540,I36543,I36546,I36549,I36552,I36555,I1892,I1899);
OUT_INSTANCE I_2190 (I36531,I36571);
OUT_INSTANCE I_2191 (I36534,I36581);
OUT_INSTANCE I_2192 (I36537,I36591);
OUT_INSTANCE I_2193 (I36540,I36601);
OUT_INSTANCE I_2194 (I36543,I36611);
OUT_INSTANCE I_2195 (I36546,I36621);
OUT_INSTANCE I_2196 (I36549,I36631);
OUT_INSTANCE I_2197 (I36552,I36641);
OUT_INSTANCE I_2198 (I36555,I36651);
PAT_11 I_2199 (I36641,I36581,I36571,I36621,I36591,I36571,I36631,I36651,I36611,I36581,I36601,I36691,I36694,I36697,I36700,I36703,I36706,I36709,I36712,I36715,I36718,I1892,I1899);
OUT_INSTANCE I_2200 (I36691,I36734);
OUT_INSTANCE I_2201 (I36694,I36744);
OUT_INSTANCE I_2202 (I36697,I36754);
OUT_INSTANCE I_2203 (I36700,I36764);
OUT_INSTANCE I_2204 (I36703,I36774);
OUT_INSTANCE I_2205 (I36706,I36784);
OUT_INSTANCE I_2206 (I36709,I36794);
OUT_INSTANCE I_2207 (I36712,I36804);
OUT_INSTANCE I_2208 (I36715,I36814);
OUT_INSTANCE I_2209 (I36718,I36824);
PAT_8 I_2210 (I36764,I36784,I36794,I36814,I36804,I36774,I36734,I36734,I36824,I36744,I36754,I36864,I36867,I36870,I36873,I36876,I36879,I36882,I36885,I36888,I1892,I1899);
OUT_INSTANCE I_2211 (I36864,I36904);
OUT_INSTANCE I_2212 (I36867,I36914);
OUT_INSTANCE I_2213 (I36870,I36924);
OUT_INSTANCE I_2214 (I36873,I36934);
OUT_INSTANCE I_2215 (I36876,I36944);
OUT_INSTANCE I_2216 (I36879,I36954);
OUT_INSTANCE I_2217 (I36882,I36964);
OUT_INSTANCE I_2218 (I36885,I36974);
OUT_INSTANCE I_2219 (I36888,I36984);
PAT_12 I_2220 (I36904,I36914,I36914,I36984,I36934,I36964,I36974,I36944,I36924,I36954,I36904,I37024,I37027,I37030,I37033,I37036,I37039,I37042,I37045,I1892,I1899);
OUT_INSTANCE I_2221 (I37024,I37061);
OUT_INSTANCE I_2222 (I37027,I37071);
OUT_INSTANCE I_2223 (I37030,I37081);
OUT_INSTANCE I_2224 (I37033,I37091);
OUT_INSTANCE I_2225 (I37036,I37101);
OUT_INSTANCE I_2226 (I37039,I37111);
OUT_INSTANCE I_2227 (I37042,I37121);
OUT_INSTANCE I_2228 (I37045,I37131);
PAT_10 I_2229 (I37061,I37131,I37101,I37111,I37081,I37071,I37061,I37121,I37081,I37091,I37071,I37171,I37174,I37177,I37180,I37183,I37186,I37189,I37192,I1892,I1899);
OUT_INSTANCE I_2230 (I37171,I37208);
OUT_INSTANCE I_2231 (I37174,I37218);
OUT_INSTANCE I_2232 (I37177,I37228);
OUT_INSTANCE I_2233 (I37180,I37238);
OUT_INSTANCE I_2234 (I37183,I37248);
OUT_INSTANCE I_2235 (I37186,I37258);
OUT_INSTANCE I_2236 (I37189,I37268);
OUT_INSTANCE I_2237 (I37192,I37278);
PAT_6 I_2238 (I37278,I37258,I37238,I37218,I37208,I37228,I37208,I37228,I37218,I37248,I37268,I37318,I37321,I37324,I37327,I37330,I37333,I37336,I37339,I37342,I37345,I1892,I1899);
OUT_INSTANCE I_2239 (I37318,I37361);
OUT_INSTANCE I_2240 (I37321,I37371);
OUT_INSTANCE I_2241 (I37324,I37381);
OUT_INSTANCE I_2242 (I37327,I37391);
OUT_INSTANCE I_2243 (I37330,I37401);
OUT_INSTANCE I_2244 (I37333,I37411);
OUT_INSTANCE I_2245 (I37336,I37421);
OUT_INSTANCE I_2246 (I37339,I37431);
OUT_INSTANCE I_2247 (I37342,I37441);
OUT_INSTANCE I_2248 (I37345,I37451);
PAT_10 I_2249 (I37361,I37411,I37421,I37391,I37361,I37441,I37451,I37371,I37401,I37381,I37431,I37491,I37494,I37497,I37500,I37503,I37506,I37509,I37512,I1892,I1899);
OUT_INSTANCE I_2250 (I37491,I37528);
OUT_INSTANCE I_2251 (I37494,I37538);
OUT_INSTANCE I_2252 (I37497,I37548);
OUT_INSTANCE I_2253 (I37500,I37558);
OUT_INSTANCE I_2254 (I37503,I37568);
OUT_INSTANCE I_2255 (I37506,I37578);
OUT_INSTANCE I_2256 (I37509,I37588);
OUT_INSTANCE I_2257 (I37512,I37598);
PAT_9 I_2258 (I37568,I37528,I37538,I37548,I37528,I37548,I37558,I37538,I37598,I37578,I37588,I37638,I37641,I37644,I37647,I37650,I37653,I37656,I37659,I37662,I1892,I1899);
OUT_INSTANCE I_2259 (I37638,I37678);
OUT_INSTANCE I_2260 (I37641,I37688);
OUT_INSTANCE I_2261 (I37644,I37698);
OUT_INSTANCE I_2262 (I37647,I37708);
OUT_INSTANCE I_2263 (I37650,I37718);
OUT_INSTANCE I_2264 (I37653,I37728);
OUT_INSTANCE I_2265 (I37656,I37738);
OUT_INSTANCE I_2266 (I37659,I37748);
OUT_INSTANCE I_2267 (I37662,I37758);
PAT_6 I_2268 (I37738,I37678,I37718,I37748,I37678,I37708,I37698,I37758,I37728,I37688,I37688,I37798,I37801,I37804,I37807,I37810,I37813,I37816,I37819,I37822,I37825,I1892,I1899);
OUT_INSTANCE I_2269 (I37798,I37841);
OUT_INSTANCE I_2270 (I37801,I37851);
OUT_INSTANCE I_2271 (I37804,I37861);
OUT_INSTANCE I_2272 (I37807,I37871);
OUT_INSTANCE I_2273 (I37810,I37881);
OUT_INSTANCE I_2274 (I37813,I37891);
OUT_INSTANCE I_2275 (I37816,I37901);
OUT_INSTANCE I_2276 (I37819,I37911);
OUT_INSTANCE I_2277 (I37822,I37921);
OUT_INSTANCE I_2278 (I37825,I37931);
PAT_17 I_2279 (I37881,I37891,I37911,I37871,I37851,I37921,I37901,I37841,I37931,I37861,I37841,I37971,I37974,I37977,I37980,I37983,I37986,I37989,I37992,I37995,I37998,I1892,I1899);
OUT_INSTANCE I_2280 (I37971,I38014);
OUT_INSTANCE I_2281 (I37974,I38024);
OUT_INSTANCE I_2282 (I37977,I38034);
OUT_INSTANCE I_2283 (I37980,I38044);
OUT_INSTANCE I_2284 (I37983,I38054);
OUT_INSTANCE I_2285 (I37986,I38064);
OUT_INSTANCE I_2286 (I37989,I38074);
OUT_INSTANCE I_2287 (I37992,I38084);
OUT_INSTANCE I_2288 (I37995,I38094);
OUT_INSTANCE I_2289 (I37998,I38104);
PAT_13 I_2290 (I38074,I38084,I38034,I38014,I38054,I38094,I38024,I38064,I38014,I38104,I38044,I38144,I38147,I38150,I38153,I38156,I38159,I38162,I38165,I38168,I1892,I1899);
OUT_INSTANCE I_2291 (I38144,I38184);
OUT_INSTANCE I_2292 (I38147,I38194);
OUT_INSTANCE I_2293 (I38150,I38204);
OUT_INSTANCE I_2294 (I38153,I38214);
OUT_INSTANCE I_2295 (I38156,I38224);
OUT_INSTANCE I_2296 (I38159,I38234);
OUT_INSTANCE I_2297 (I38162,I38244);
OUT_INSTANCE I_2298 (I38165,I38254);
OUT_INSTANCE I_2299 (I38168,I38264);
PAT_2 I_2300 (I38244,I38224,I38214,I38234,I38184,I38264,I38194,I38254,I38184,I38204,I38194,I38304,I38307,I38310,I38313,I38316,I38319,I38322,I38325,I38328,I1892,I1899);
OUT_INSTANCE I_2301 (I38304,I38344);
OUT_INSTANCE I_2302 (I38307,I38354);
OUT_INSTANCE I_2303 (I38310,I38364);
OUT_INSTANCE I_2304 (I38313,I38374);
OUT_INSTANCE I_2305 (I38316,I38384);
OUT_INSTANCE I_2306 (I38319,I38394);
OUT_INSTANCE I_2307 (I38322,I38404);
OUT_INSTANCE I_2308 (I38325,I38414);
OUT_INSTANCE I_2309 (I38328,I38424);
PAT_16 I_2310 (I38404,I38344,I38414,I38374,I38344,I38384,I38364,I38354,I38354,I38424,I38394,I38464,I38467,I38470,I38473,I38476,I38479,I38482,I38485,I38488,I38491,I1892,I1899);
OUT_INSTANCE I_2311 (I38464,I38507);
OUT_INSTANCE I_2312 (I38467,I38517);
OUT_INSTANCE I_2313 (I38470,I38527);
OUT_INSTANCE I_2314 (I38473,I38537);
OUT_INSTANCE I_2315 (I38476,I38547);
OUT_INSTANCE I_2316 (I38479,I38557);
OUT_INSTANCE I_2317 (I38482,I38567);
OUT_INSTANCE I_2318 (I38485,I38577);
OUT_INSTANCE I_2319 (I38488,I38587);
OUT_INSTANCE I_2320 (I38491,I38597);
PAT_13 I_2321 (I38547,I38517,I38507,I38527,I38557,I38587,I38577,I38567,I38537,I38507,I38597,I38637,I38640,I38643,I38646,I38649,I38652,I38655,I38658,I38661,I1892,I1899);
OUT_INSTANCE I_2322 (I38637,I38677);
OUT_INSTANCE I_2323 (I38640,I38687);
OUT_INSTANCE I_2324 (I38643,I38697);
OUT_INSTANCE I_2325 (I38646,I38707);
OUT_INSTANCE I_2326 (I38649,I38717);
OUT_INSTANCE I_2327 (I38652,I38727);
OUT_INSTANCE I_2328 (I38655,I38737);
OUT_INSTANCE I_2329 (I38658,I38747);
OUT_INSTANCE I_2330 (I38661,I38757);
PAT_1 I_2331 (I38677,I38707,I38687,I38747,I38727,I38697,I38737,I38717,I38687,I38757,I38677,I38797,I38800,I38803,I38806,I38809,I38812,I38815,I38818,I38821,I1892,I1899);
OUT_INSTANCE I_2332 (I38797,I38837);
OUT_INSTANCE I_2333 (I38800,I38847);
OUT_INSTANCE I_2334 (I38803,I38857);
OUT_INSTANCE I_2335 (I38806,I38867);
OUT_INSTANCE I_2336 (I38809,I38877);
OUT_INSTANCE I_2337 (I38812,I38887);
OUT_INSTANCE I_2338 (I38815,I38897);
OUT_INSTANCE I_2339 (I38818,I38907);
OUT_INSTANCE I_2340 (I38821,I38917);
PAT_12 I_2341 (I38877,I38857,I38917,I38837,I38867,I38837,I38847,I38907,I38887,I38847,I38897,I38957,I38960,I38963,I38966,I38969,I38972,I38975,I38978,I1892,I1899);
OUT_INSTANCE I_2342 (I38957,I38994);
OUT_INSTANCE I_2343 (I38960,I39004);
OUT_INSTANCE I_2344 (I38963,I39014);
OUT_INSTANCE I_2345 (I38966,I39024);
OUT_INSTANCE I_2346 (I38969,I39034);
OUT_INSTANCE I_2347 (I38972,I39044);
OUT_INSTANCE I_2348 (I38975,I39054);
OUT_INSTANCE I_2349 (I38978,I39064);
PAT_1 I_2350 (I39044,I39004,I39054,I39024,I38994,I39004,I39034,I38994,I39064,I39014,I39014,I39104,I39107,I39110,I39113,I39116,I39119,I39122,I39125,I39128,I1892,I1899);
OUT_INSTANCE I_2351 (I39104,I39144);
OUT_INSTANCE I_2352 (I39107,I39154);
OUT_INSTANCE I_2353 (I39110,I39164);
OUT_INSTANCE I_2354 (I39113,I39174);
OUT_INSTANCE I_2355 (I39116,I39184);
OUT_INSTANCE I_2356 (I39119,I39194);
OUT_INSTANCE I_2357 (I39122,I39204);
OUT_INSTANCE I_2358 (I39125,I39214);
OUT_INSTANCE I_2359 (I39128,I39224);
PAT_6 I_2360 (I39174,I39144,I39154,I39164,I39214,I39224,I39204,I39144,I39194,I39184,I39154,I39264,I39267,I39270,I39273,I39276,I39279,I39282,I39285,I39288,I39291,I1892,I1899);
OUT_INSTANCE I_2361 (I39264,I39307);
OUT_INSTANCE I_2362 (I39267,I39317);
OUT_INSTANCE I_2363 (I39270,I39327);
OUT_INSTANCE I_2364 (I39273,I39337);
OUT_INSTANCE I_2365 (I39276,I39347);
OUT_INSTANCE I_2366 (I39279,I39357);
OUT_INSTANCE I_2367 (I39282,I39367);
OUT_INSTANCE I_2368 (I39285,I39377);
OUT_INSTANCE I_2369 (I39288,I39387);
OUT_INSTANCE I_2370 (I39291,I39397);
PAT_2 I_2371 (I39377,I39397,I39337,I39357,I39307,I39327,I39307,I39347,I39317,I39367,I39387,I39437,I39440,I39443,I39446,I39449,I39452,I39455,I39458,I39461,I1892,I1899);
OUT_INSTANCE I_2372 (I39437,I39477);
OUT_INSTANCE I_2373 (I39440,I39487);
OUT_INSTANCE I_2374 (I39443,I39497);
OUT_INSTANCE I_2375 (I39446,I39507);
OUT_INSTANCE I_2376 (I39449,I39517);
OUT_INSTANCE I_2377 (I39452,I39527);
OUT_INSTANCE I_2378 (I39455,I39537);
OUT_INSTANCE I_2379 (I39458,I39547);
OUT_INSTANCE I_2380 (I39461,I39557);
PAT_11 I_2381 (I39487,I39527,I39477,I39517,I39507,I39547,I39537,I39487,I39557,I39497,I39477,I39597,I39600,I39603,I39606,I39609,I39612,I39615,I39618,I39621,I39624,I1892,I1899);
OUT_INSTANCE I_2382 (I39597,I39640);
OUT_INSTANCE I_2383 (I39600,I39650);
OUT_INSTANCE I_2384 (I39603,I39660);
OUT_INSTANCE I_2385 (I39606,I39670);
OUT_INSTANCE I_2386 (I39609,I39680);
OUT_INSTANCE I_2387 (I39612,I39690);
OUT_INSTANCE I_2388 (I39615,I39700);
OUT_INSTANCE I_2389 (I39618,I39710);
OUT_INSTANCE I_2390 (I39621,I39720);
OUT_INSTANCE I_2391 (I39624,I39730);
PAT_9 I_2392 (I39660,I39700,I39670,I39710,I39640,I39650,I39680,I39640,I39690,I39720,I39730,I39770,I39773,I39776,I39779,I39782,I39785,I39788,I39791,I39794,I1892,I1899);
OUT_INSTANCE I_2393 (I39770,I39810);
OUT_INSTANCE I_2394 (I39773,I39820);
OUT_INSTANCE I_2395 (I39776,I39830);
OUT_INSTANCE I_2396 (I39779,I39840);
OUT_INSTANCE I_2397 (I39782,I39850);
OUT_INSTANCE I_2398 (I39785,I39860);
OUT_INSTANCE I_2399 (I39788,I39870);
OUT_INSTANCE I_2400 (I39791,I39880);
OUT_INSTANCE I_2401 (I39794,I39890);
PAT_2 I_2402 (I39860,I39870,I39840,I39890,I39810,I39820,I39830,I39820,I39880,I39850,I39810,I39930,I39933,I39936,I39939,I39942,I39945,I39948,I39951,I39954,I1892,I1899);
OUT_INSTANCE I_2403 (I39930,I39970);
OUT_INSTANCE I_2404 (I39933,I39980);
OUT_INSTANCE I_2405 (I39936,I39990);
OUT_INSTANCE I_2406 (I39939,I40000);
OUT_INSTANCE I_2407 (I39942,I40010);
OUT_INSTANCE I_2408 (I39945,I40020);
OUT_INSTANCE I_2409 (I39948,I40030);
OUT_INSTANCE I_2410 (I39951,I40040);
OUT_INSTANCE I_2411 (I39954,I40050);
PAT_17 I_2412 (I39970,I39970,I40010,I39980,I39990,I40030,I40020,I40050,I39980,I40000,I40040,I40090,I40093,I40096,I40099,I40102,I40105,I40108,I40111,I40114,I40117,I1892,I1899);
OUT_INSTANCE I_2413 (I40090,I40133);
OUT_INSTANCE I_2414 (I40093,I40143);
OUT_INSTANCE I_2415 (I40096,I40153);
OUT_INSTANCE I_2416 (I40099,I40163);
OUT_INSTANCE I_2417 (I40102,I40173);
OUT_INSTANCE I_2418 (I40105,I40183);
OUT_INSTANCE I_2419 (I40108,I40193);
OUT_INSTANCE I_2420 (I40111,I40203);
OUT_INSTANCE I_2421 (I40114,I40213);
OUT_INSTANCE I_2422 (I40117,I40223);
PAT_16 I_2423 (I40133,I40213,I40133,I40203,I40193,I40153,I40173,I40143,I40223,I40183,I40163,I40263,I40266,I40269,I40272,I40275,I40278,I40281,I40284,I40287,I40290,I1892,I1899);
OUT_INSTANCE I_2424 (I40263,I40306);
OUT_INSTANCE I_2425 (I40266,I40316);
OUT_INSTANCE I_2426 (I40269,I40326);
OUT_INSTANCE I_2427 (I40272,I40336);
OUT_INSTANCE I_2428 (I40275,I40346);
OUT_INSTANCE I_2429 (I40278,I40356);
OUT_INSTANCE I_2430 (I40281,I40366);
OUT_INSTANCE I_2431 (I40284,I40376);
OUT_INSTANCE I_2432 (I40287,I40386);
OUT_INSTANCE I_2433 (I40290,I40396);
PAT_4 I_2434 (I40346,I40366,I40316,I40356,I40306,I40326,I40336,I40376,I40386,I40306,I40396,I40436,I40439,I40442,I40445,I40448,I40451,I40454,I40457,I40460,I1892,I1899);
OUT_INSTANCE I_2435 (I40436,I40476);
OUT_INSTANCE I_2436 (I40439,I40486);
OUT_INSTANCE I_2437 (I40442,I40496);
OUT_INSTANCE I_2438 (I40445,I40506);
OUT_INSTANCE I_2439 (I40448,I40516);
OUT_INSTANCE I_2440 (I40451,I40526);
OUT_INSTANCE I_2441 (I40454,I40536);
OUT_INSTANCE I_2442 (I40457,I40546);
OUT_INSTANCE I_2443 (I40460,I40556);
PAT_1 I_2444 (I40476,I40546,I40536,I40486,I40526,I40476,I40486,I40556,I40506,I40496,I40516,I40596,I40599,I40602,I40605,I40608,I40611,I40614,I40617,I40620,I1892,I1899);
OUT_INSTANCE I_2445 (I40596,I40636);
OUT_INSTANCE I_2446 (I40599,I40646);
OUT_INSTANCE I_2447 (I40602,I40656);
OUT_INSTANCE I_2448 (I40605,I40666);
OUT_INSTANCE I_2449 (I40608,I40676);
OUT_INSTANCE I_2450 (I40611,I40686);
OUT_INSTANCE I_2451 (I40614,I40696);
OUT_INSTANCE I_2452 (I40617,I40706);
OUT_INSTANCE I_2453 (I40620,I40716);
PAT_7 I_2454 (I40646,I40666,I40656,I40676,I40696,I40686,I40716,I40706,I40646,I40636,I40636,I40756,I40759,I40762,I40765,I40768,I40771,I40774,I40777,I40780,I1892,I1899);
OUT_INSTANCE I_2455 (I40756,I40796);
OUT_INSTANCE I_2456 (I40759,I40806);
OUT_INSTANCE I_2457 (I40762,I40816);
OUT_INSTANCE I_2458 (I40765,I40826);
OUT_INSTANCE I_2459 (I40768,I40836);
OUT_INSTANCE I_2460 (I40771,I40846);
OUT_INSTANCE I_2461 (I40774,I40856);
OUT_INSTANCE I_2462 (I40777,I40866);
OUT_INSTANCE I_2463 (I40780,I40876);
PAT_6 I_2464 (I40796,I40856,I40796,I40826,I40846,I40806,I40866,I40816,I40876,I40806,I40836,I40916,I40919,I40922,I40925,I40928,I40931,I40934,I40937,I40940,I40943,I1892,I1899);
OUT_INSTANCE I_2465 (I40916,I40959);
OUT_INSTANCE I_2466 (I40919,I40969);
OUT_INSTANCE I_2467 (I40922,I40979);
OUT_INSTANCE I_2468 (I40925,I40989);
OUT_INSTANCE I_2469 (I40928,I40999);
OUT_INSTANCE I_2470 (I40931,I41009);
OUT_INSTANCE I_2471 (I40934,I41019);
OUT_INSTANCE I_2472 (I40937,I41029);
OUT_INSTANCE I_2473 (I40940,I41039);
OUT_INSTANCE I_2474 (I40943,I41049);
PAT_5 I_2475 (I41029,I40959,I40979,I40989,I41009,I41019,I40959,I41039,I40969,I40999,I41049,I41089,I41092,I41095,I41098,I41101,I41104,I41107,I41110,I41113,I41116,I1892,I1899);
OUT_INSTANCE I_2476 (I41089,I41132);
OUT_INSTANCE I_2477 (I41092,I41142);
OUT_INSTANCE I_2478 (I41095,I41152);
OUT_INSTANCE I_2479 (I41098,I41162);
OUT_INSTANCE I_2480 (I41101,I41172);
OUT_INSTANCE I_2481 (I41104,I41182);
OUT_INSTANCE I_2482 (I41107,I41192);
OUT_INSTANCE I_2483 (I41110,I41202);
OUT_INSTANCE I_2484 (I41113,I41212);
OUT_INSTANCE I_2485 (I41116,I41222);
PAT_6 I_2486 (I41192,I41172,I41132,I41152,I41142,I41162,I41182,I41132,I41212,I41202,I41222,I41262,I41265,I41268,I41271,I41274,I41277,I41280,I41283,I41286,I41289,I1892,I1899);
OUT_INSTANCE I_2487 (I41262,I41305);
OUT_INSTANCE I_2488 (I41265,I41315);
OUT_INSTANCE I_2489 (I41268,I41325);
OUT_INSTANCE I_2490 (I41271,I41335);
OUT_INSTANCE I_2491 (I41274,I41345);
OUT_INSTANCE I_2492 (I41277,I41355);
OUT_INSTANCE I_2493 (I41280,I41365);
OUT_INSTANCE I_2494 (I41283,I41375);
OUT_INSTANCE I_2495 (I41286,I41385);
OUT_INSTANCE I_2496 (I41289,I41395);
PAT_10 I_2497 (I41305,I41355,I41365,I41335,I41305,I41385,I41395,I41315,I41345,I41325,I41375,I41435,I41438,I41441,I41444,I41447,I41450,I41453,I41456,I1892,I1899);
OUT_INSTANCE I_2498 (I41435,I41472);
OUT_INSTANCE I_2499 (I41438,I41482);
OUT_INSTANCE I_2500 (I41441,I41492);
OUT_INSTANCE I_2501 (I41444,I41502);
OUT_INSTANCE I_2502 (I41447,I41512);
OUT_INSTANCE I_2503 (I41450,I41522);
OUT_INSTANCE I_2504 (I41453,I41532);
OUT_INSTANCE I_2505 (I41456,I41542);
PAT_11 I_2506 (I41502,I41512,I41542,I41522,I41532,I41472,I41472,I41492,I41482,I41482,I41492,I41582,I41585,I41588,I41591,I41594,I41597,I41600,I41603,I41606,I41609,I1892,I1899);
OUT_INSTANCE I_2507 (I41582,I41625);
OUT_INSTANCE I_2508 (I41585,I41635);
OUT_INSTANCE I_2509 (I41588,I41645);
OUT_INSTANCE I_2510 (I41591,I41655);
OUT_INSTANCE I_2511 (I41594,I41665);
OUT_INSTANCE I_2512 (I41597,I41675);
OUT_INSTANCE I_2513 (I41600,I41685);
OUT_INSTANCE I_2514 (I41603,I41695);
OUT_INSTANCE I_2515 (I41606,I41705);
OUT_INSTANCE I_2516 (I41609,I41715);
PAT_2 I_2517 (I41625,I41705,I41665,I41645,I41675,I41685,I41635,I41715,I41695,I41655,I41625,I41755,I41758,I41761,I41764,I41767,I41770,I41773,I41776,I41779,I1892,I1899);
OUT_INSTANCE I_2518 (I41755,I41795);
OUT_INSTANCE I_2519 (I41758,I41805);
OUT_INSTANCE I_2520 (I41761,I41815);
OUT_INSTANCE I_2521 (I41764,I41825);
OUT_INSTANCE I_2522 (I41767,I41835);
OUT_INSTANCE I_2523 (I41770,I41845);
OUT_INSTANCE I_2524 (I41773,I41855);
OUT_INSTANCE I_2525 (I41776,I41865);
OUT_INSTANCE I_2526 (I41779,I41875);
PAT_4 I_2527 (I41795,I41815,I41875,I41855,I41845,I41835,I41805,I41865,I41795,I41805,I41825,I41915,I41918,I41921,I41924,I41927,I41930,I41933,I41936,I41939,I1892,I1899);
OUT_INSTANCE I_2528 (I41915,I41955);
OUT_INSTANCE I_2529 (I41918,I41965);
OUT_INSTANCE I_2530 (I41921,I41975);
OUT_INSTANCE I_2531 (I41924,I41985);
OUT_INSTANCE I_2532 (I41927,I41995);
OUT_INSTANCE I_2533 (I41930,I42005);
OUT_INSTANCE I_2534 (I41933,I42015);
OUT_INSTANCE I_2535 (I41936,I42025);
OUT_INSTANCE I_2536 (I41939,I42035);
PAT_9 I_2537 (I42025,I41965,I41975,I42005,I42015,I41955,I41985,I41965,I42035,I41955,I41995,I42075,I42078,I42081,I42084,I42087,I42090,I42093,I42096,I42099,I1892,I1899);
OUT_INSTANCE I_2538 (I42075,I42115);
OUT_INSTANCE I_2539 (I42078,I42125);
OUT_INSTANCE I_2540 (I42081,I42135);
OUT_INSTANCE I_2541 (I42084,I42145);
OUT_INSTANCE I_2542 (I42087,I42155);
OUT_INSTANCE I_2543 (I42090,I42165);
OUT_INSTANCE I_2544 (I42093,I42175);
OUT_INSTANCE I_2545 (I42096,I42185);
OUT_INSTANCE I_2546 (I42099,I42195);
IN_INSTANCE I_2547 (I1573,I42205);
IN_INSTANCE I_2548 (I1565,I42215);
IN_INSTANCE I_2549 (I1669,I42225);
IN_INSTANCE I_2550 (I1773,I42235);
IN_INSTANCE I_2551 (I1853,I42245);
IN_INSTANCE I_2552 (I1469,I42255);
IN_INSTANCE I_2553 (I1373,I42265);
IN_INSTANCE I_2554 (I1493,I42275);
IN_INSTANCE I_2555 (I1797,I42285);
IN_INSTANCE I_2556 (I1461,I42295);
IN_INSTANCE I_2557 (I1381,I42305);
PAT_11 I_2558 (I42205,I42215,I42225,I42235,I42245,I42255,I42265,I42275,I42285,I42295,I42305,I42345,I42348,I42351,I42354,I42357,I42360,I42363,I42366,I42369,I42372,I1892,I1899);
OUT_INSTANCE I_2559 (I42345,I42388);
OUT_INSTANCE I_2560 (I42348,I42398);
OUT_INSTANCE I_2561 (I42351,I42408);
OUT_INSTANCE I_2562 (I42354,I42418);
OUT_INSTANCE I_2563 (I42357,I42428);
OUT_INSTANCE I_2564 (I42360,I42438);
OUT_INSTANCE I_2565 (I42363,I42448);
OUT_INSTANCE I_2566 (I42366,I42458);
OUT_INSTANCE I_2567 (I42369,I42468);
OUT_INSTANCE I_2568 (I42372,I42478);
PAT_4 I_2569 (I42408,I42478,I42388,I42448,I42418,I42388,I42458,I42398,I42428,I42468,I42438,I42518,I42521,I42524,I42527,I42530,I42533,I42536,I42539,I42542,I1892,I1899);
OUT_INSTANCE I_2570 (I42518,I42558);
OUT_INSTANCE I_2571 (I42521,I42568);
OUT_INSTANCE I_2572 (I42524,I42578);
OUT_INSTANCE I_2573 (I42527,I42588);
OUT_INSTANCE I_2574 (I42530,I42598);
OUT_INSTANCE I_2575 (I42533,I42608);
OUT_INSTANCE I_2576 (I42536,I42618);
OUT_INSTANCE I_2577 (I42539,I42628);
OUT_INSTANCE I_2578 (I42542,I42638);
PAT_9 I_2579 (I42628,I42568,I42578,I42608,I42618,I42558,I42588,I42568,I42638,I42558,I42598,I42678,I42681,I42684,I42687,I42690,I42693,I42696,I42699,I42702,I1892,I1899);
OUT_INSTANCE I_2580 (I42678,I42718);
OUT_INSTANCE I_2581 (I42681,I42728);
OUT_INSTANCE I_2582 (I42684,I42738);
OUT_INSTANCE I_2583 (I42687,I42748);
OUT_INSTANCE I_2584 (I42690,I42758);
OUT_INSTANCE I_2585 (I42693,I42768);
OUT_INSTANCE I_2586 (I42696,I42778);
OUT_INSTANCE I_2587 (I42699,I42788);
OUT_INSTANCE I_2588 (I42702,I42798);
PAT_1 I_2589 (I42718,I42778,I42718,I42758,I42728,I42748,I42768,I42788,I42798,I42738,I42728,I42838,I42841,I42844,I42847,I42850,I42853,I42856,I42859,I42862,I1892,I1899);
OUT_INSTANCE I_2590 (I42838,I42878);
OUT_INSTANCE I_2591 (I42841,I42888);
OUT_INSTANCE I_2592 (I42844,I42898);
OUT_INSTANCE I_2593 (I42847,I42908);
OUT_INSTANCE I_2594 (I42850,I42918);
OUT_INSTANCE I_2595 (I42853,I42928);
OUT_INSTANCE I_2596 (I42856,I42938);
OUT_INSTANCE I_2597 (I42859,I42948);
OUT_INSTANCE I_2598 (I42862,I42958);
PAT_5 I_2599 (I42938,I42948,I42888,I42918,I42908,I42898,I42928,I42958,I42888,I42878,I42878,I42998,I43001,I43004,I43007,I43010,I43013,I43016,I43019,I43022,I43025,I1892,I1899);
OUT_INSTANCE I_2600 (I42998,I43041);
OUT_INSTANCE I_2601 (I43001,I43051);
OUT_INSTANCE I_2602 (I43004,I43061);
OUT_INSTANCE I_2603 (I43007,I43071);
OUT_INSTANCE I_2604 (I43010,I43081);
OUT_INSTANCE I_2605 (I43013,I43091);
OUT_INSTANCE I_2606 (I43016,I43101);
OUT_INSTANCE I_2607 (I43019,I43111);
OUT_INSTANCE I_2608 (I43022,I43121);
OUT_INSTANCE I_2609 (I43025,I43131);
PAT_10 I_2610 (I43121,I43131,I43061,I43081,I43091,I43111,I43051,I43041,I43041,I43071,I43101,I43171,I43174,I43177,I43180,I43183,I43186,I43189,I43192,I1892,I1899);
OUT_INSTANCE I_2611 (I43171,I43208);
OUT_INSTANCE I_2612 (I43174,I43218);
OUT_INSTANCE I_2613 (I43177,I43228);
OUT_INSTANCE I_2614 (I43180,I43238);
OUT_INSTANCE I_2615 (I43183,I43248);
OUT_INSTANCE I_2616 (I43186,I43258);
OUT_INSTANCE I_2617 (I43189,I43268);
OUT_INSTANCE I_2618 (I43192,I43278);
PAT_9 I_2619 (I43248,I43208,I43218,I43228,I43208,I43228,I43238,I43218,I43278,I43258,I43268,I43318,I43321,I43324,I43327,I43330,I43333,I43336,I43339,I43342,I1892,I1899);
OUT_INSTANCE I_2620 (I43318,I43358);
OUT_INSTANCE I_2621 (I43321,I43368);
OUT_INSTANCE I_2622 (I43324,I43378);
OUT_INSTANCE I_2623 (I43327,I43388);
OUT_INSTANCE I_2624 (I43330,I43398);
OUT_INSTANCE I_2625 (I43333,I43408);
OUT_INSTANCE I_2626 (I43336,I43418);
OUT_INSTANCE I_2627 (I43339,I43428);
OUT_INSTANCE I_2628 (I43342,I43438);
PAT_2 I_2629 (I43408,I43418,I43388,I43438,I43358,I43368,I43378,I43368,I43428,I43398,I43358,I43478,I43481,I43484,I43487,I43490,I43493,I43496,I43499,I43502,I1892,I1899);
OUT_INSTANCE I_2630 (I43478,I43518);
OUT_INSTANCE I_2631 (I43481,I43528);
OUT_INSTANCE I_2632 (I43484,I43538);
OUT_INSTANCE I_2633 (I43487,I43548);
OUT_INSTANCE I_2634 (I43490,I43558);
OUT_INSTANCE I_2635 (I43493,I43568);
OUT_INSTANCE I_2636 (I43496,I43578);
OUT_INSTANCE I_2637 (I43499,I43588);
OUT_INSTANCE I_2638 (I43502,I43598);
PAT_17 I_2639 (I43518,I43518,I43558,I43528,I43538,I43578,I43568,I43598,I43528,I43548,I43588,I43638,I43641,I43644,I43647,I43650,I43653,I43656,I43659,I43662,I43665,I1892,I1899);
OUT_INSTANCE I_2640 (I43638,I43681);
OUT_INSTANCE I_2641 (I43641,I43691);
OUT_INSTANCE I_2642 (I43644,I43701);
OUT_INSTANCE I_2643 (I43647,I43711);
OUT_INSTANCE I_2644 (I43650,I43721);
OUT_INSTANCE I_2645 (I43653,I43731);
OUT_INSTANCE I_2646 (I43656,I43741);
OUT_INSTANCE I_2647 (I43659,I43751);
OUT_INSTANCE I_2648 (I43662,I43761);
OUT_INSTANCE I_2649 (I43665,I43771);
PAT_14 I_2650 (I43691,I43741,I43681,I43761,I43711,I43731,I43681,I43751,I43701,I43771,I43721,I43811,I43814,I43817,I43820,I43823,I43826,I43829,I43832,I43835,I1892,I1899);
OUT_INSTANCE I_2651 (I43811,I43851);
OUT_INSTANCE I_2652 (I43814,I43861);
OUT_INSTANCE I_2653 (I43817,I43871);
OUT_INSTANCE I_2654 (I43820,I43881);
OUT_INSTANCE I_2655 (I43823,I43891);
OUT_INSTANCE I_2656 (I43826,I43901);
OUT_INSTANCE I_2657 (I43829,I43911);
OUT_INSTANCE I_2658 (I43832,I43921);
OUT_INSTANCE I_2659 (I43835,I43931);
PAT_9 I_2660 (I43881,I43921,I43851,I43911,I43861,I43871,I43931,I43861,I43891,I43851,I43901,I43971,I43974,I43977,I43980,I43983,I43986,I43989,I43992,I43995,I1892,I1899);
OUT_INSTANCE I_2661 (I43971,I44011);
OUT_INSTANCE I_2662 (I43974,I44021);
OUT_INSTANCE I_2663 (I43977,I44031);
OUT_INSTANCE I_2664 (I43980,I44041);
OUT_INSTANCE I_2665 (I43983,I44051);
OUT_INSTANCE I_2666 (I43986,I44061);
OUT_INSTANCE I_2667 (I43989,I44071);
OUT_INSTANCE I_2668 (I43992,I44081);
OUT_INSTANCE I_2669 (I43995,I44091);
PAT_6 I_2670 (I44071,I44011,I44051,I44081,I44011,I44041,I44031,I44091,I44061,I44021,I44021,I44131,I44134,I44137,I44140,I44143,I44146,I44149,I44152,I44155,I44158,I1892,I1899);
OUT_INSTANCE I_2671 (I44131,I44174);
OUT_INSTANCE I_2672 (I44134,I44184);
OUT_INSTANCE I_2673 (I44137,I44194);
OUT_INSTANCE I_2674 (I44140,I44204);
OUT_INSTANCE I_2675 (I44143,I44214);
OUT_INSTANCE I_2676 (I44146,I44224);
OUT_INSTANCE I_2677 (I44149,I44234);
OUT_INSTANCE I_2678 (I44152,I44244);
OUT_INSTANCE I_2679 (I44155,I44254);
OUT_INSTANCE I_2680 (I44158,I44264);
PAT_5 I_2681 (I44244,I44174,I44194,I44204,I44224,I44234,I44174,I44254,I44184,I44214,I44264,I44304,I44307,I44310,I44313,I44316,I44319,I44322,I44325,I44328,I44331,I1892,I1899);
OUT_INSTANCE I_2682 (I44304,I44347);
OUT_INSTANCE I_2683 (I44307,I44357);
OUT_INSTANCE I_2684 (I44310,I44367);
OUT_INSTANCE I_2685 (I44313,I44377);
OUT_INSTANCE I_2686 (I44316,I44387);
OUT_INSTANCE I_2687 (I44319,I44397);
OUT_INSTANCE I_2688 (I44322,I44407);
OUT_INSTANCE I_2689 (I44325,I44417);
OUT_INSTANCE I_2690 (I44328,I44427);
OUT_INSTANCE I_2691 (I44331,I44437);
PAT_13 I_2692 (I44367,I44397,I44347,I44357,I44427,I44377,I44417,I44347,I44407,I44437,I44387,I44477,I44480,I44483,I44486,I44489,I44492,I44495,I44498,I44501,I1892,I1899);
OUT_INSTANCE I_2693 (I44477,I44517);
OUT_INSTANCE I_2694 (I44480,I44527);
OUT_INSTANCE I_2695 (I44483,I44537);
OUT_INSTANCE I_2696 (I44486,I44547);
OUT_INSTANCE I_2697 (I44489,I44557);
OUT_INSTANCE I_2698 (I44492,I44567);
OUT_INSTANCE I_2699 (I44495,I44577);
OUT_INSTANCE I_2700 (I44498,I44587);
OUT_INSTANCE I_2701 (I44501,I44597);
PAT_2 I_2702 (I44577,I44557,I44547,I44567,I44517,I44597,I44527,I44587,I44517,I44537,I44527,I44637,I44640,I44643,I44646,I44649,I44652,I44655,I44658,I44661,I1892,I1899);
OUT_INSTANCE I_2703 (I44637,I44677);
OUT_INSTANCE I_2704 (I44640,I44687);
OUT_INSTANCE I_2705 (I44643,I44697);
OUT_INSTANCE I_2706 (I44646,I44707);
OUT_INSTANCE I_2707 (I44649,I44717);
OUT_INSTANCE I_2708 (I44652,I44727);
OUT_INSTANCE I_2709 (I44655,I44737);
OUT_INSTANCE I_2710 (I44658,I44747);
OUT_INSTANCE I_2711 (I44661,I44757);
PAT_8 I_2712 (I44717,I44687,I44707,I44677,I44697,I44747,I44737,I44677,I44727,I44687,I44757,I44797,I44800,I44803,I44806,I44809,I44812,I44815,I44818,I44821,I1892,I1899);
OUT_INSTANCE I_2713 (I44797,I44837);
OUT_INSTANCE I_2714 (I44800,I44847);
OUT_INSTANCE I_2715 (I44803,I44857);
OUT_INSTANCE I_2716 (I44806,I44867);
OUT_INSTANCE I_2717 (I44809,I44877);
OUT_INSTANCE I_2718 (I44812,I44887);
OUT_INSTANCE I_2719 (I44815,I44897);
OUT_INSTANCE I_2720 (I44818,I44907);
OUT_INSTANCE I_2721 (I44821,I44917);
PAT_14 I_2722 (I44857,I44897,I44847,I44837,I44847,I44917,I44837,I44877,I44887,I44907,I44867,I44957,I44960,I44963,I44966,I44969,I44972,I44975,I44978,I44981,I1892,I1899);
OUT_INSTANCE I_2723 (I44957,I44997);
OUT_INSTANCE I_2724 (I44960,I45007);
OUT_INSTANCE I_2725 (I44963,I45017);
OUT_INSTANCE I_2726 (I44966,I45027);
OUT_INSTANCE I_2727 (I44969,I45037);
OUT_INSTANCE I_2728 (I44972,I45047);
OUT_INSTANCE I_2729 (I44975,I45057);
OUT_INSTANCE I_2730 (I44978,I45067);
OUT_INSTANCE I_2731 (I44981,I45077);
PAT_4 I_2732 (I45027,I45047,I45017,I44997,I45077,I45037,I44997,I45007,I45067,I45007,I45057,I45117,I45120,I45123,I45126,I45129,I45132,I45135,I45138,I45141,I1892,I1899);
OUT_INSTANCE I_2733 (I45117,I45157);
OUT_INSTANCE I_2734 (I45120,I45167);
OUT_INSTANCE I_2735 (I45123,I45177);
OUT_INSTANCE I_2736 (I45126,I45187);
OUT_INSTANCE I_2737 (I45129,I45197);
OUT_INSTANCE I_2738 (I45132,I45207);
OUT_INSTANCE I_2739 (I45135,I45217);
OUT_INSTANCE I_2740 (I45138,I45227);
OUT_INSTANCE I_2741 (I45141,I45237);
PAT_2 I_2742 (I45187,I45167,I45167,I45237,I45157,I45217,I45207,I45177,I45157,I45197,I45227,I45277,I45280,I45283,I45286,I45289,I45292,I45295,I45298,I45301,I1892,I1899);
OUT_INSTANCE I_2743 (I45277,I45317);
OUT_INSTANCE I_2744 (I45280,I45327);
OUT_INSTANCE I_2745 (I45283,I45337);
OUT_INSTANCE I_2746 (I45286,I45347);
OUT_INSTANCE I_2747 (I45289,I45357);
OUT_INSTANCE I_2748 (I45292,I45367);
OUT_INSTANCE I_2749 (I45295,I45377);
OUT_INSTANCE I_2750 (I45298,I45387);
OUT_INSTANCE I_2751 (I45301,I45397);
PAT_4 I_2752 (I45317,I45337,I45397,I45377,I45367,I45357,I45327,I45387,I45317,I45327,I45347,I45437,I45440,I45443,I45446,I45449,I45452,I45455,I45458,I45461,I1892,I1899);
OUT_INSTANCE I_2753 (I45437,I45477);
OUT_INSTANCE I_2754 (I45440,I45487);
OUT_INSTANCE I_2755 (I45443,I45497);
OUT_INSTANCE I_2756 (I45446,I45507);
OUT_INSTANCE I_2757 (I45449,I45517);
OUT_INSTANCE I_2758 (I45452,I45527);
OUT_INSTANCE I_2759 (I45455,I45537);
OUT_INSTANCE I_2760 (I45458,I45547);
OUT_INSTANCE I_2761 (I45461,I45557);
PAT_6 I_2762 (I45477,I45497,I45487,I45527,I45537,I45517,I45557,I45547,I45477,I45507,I45487,I45597,I45600,I45603,I45606,I45609,I45612,I45615,I45618,I45621,I45624,I1892,I1899);
OUT_INSTANCE I_2763 (I45597,I45640);
OUT_INSTANCE I_2764 (I45600,I45650);
OUT_INSTANCE I_2765 (I45603,I45660);
OUT_INSTANCE I_2766 (I45606,I45670);
OUT_INSTANCE I_2767 (I45609,I45680);
OUT_INSTANCE I_2768 (I45612,I45690);
OUT_INSTANCE I_2769 (I45615,I45700);
OUT_INSTANCE I_2770 (I45618,I45710);
OUT_INSTANCE I_2771 (I45621,I45720);
OUT_INSTANCE I_2772 (I45624,I45730);
PAT_4 I_2773 (I45640,I45690,I45650,I45660,I45670,I45640,I45730,I45700,I45710,I45680,I45720,I45770,I45773,I45776,I45779,I45782,I45785,I45788,I45791,I45794,I1892,I1899);
OUT_INSTANCE I_2774 (I45770,I45810);
OUT_INSTANCE I_2775 (I45773,I45820);
OUT_INSTANCE I_2776 (I45776,I45830);
OUT_INSTANCE I_2777 (I45779,I45840);
OUT_INSTANCE I_2778 (I45782,I45850);
OUT_INSTANCE I_2779 (I45785,I45860);
OUT_INSTANCE I_2780 (I45788,I45870);
OUT_INSTANCE I_2781 (I45791,I45880);
OUT_INSTANCE I_2782 (I45794,I45890);
PAT_10 I_2783 (I45810,I45810,I45890,I45820,I45840,I45870,I45860,I45820,I45880,I45830,I45850,I45930,I45933,I45936,I45939,I45942,I45945,I45948,I45951,I1892,I1899);
OUT_INSTANCE I_2784 (I45930,I45967);
OUT_INSTANCE I_2785 (I45933,I45977);
OUT_INSTANCE I_2786 (I45936,I45987);
OUT_INSTANCE I_2787 (I45939,I45997);
OUT_INSTANCE I_2788 (I45942,I46007);
OUT_INSTANCE I_2789 (I45945,I46017);
OUT_INSTANCE I_2790 (I45948,I46027);
OUT_INSTANCE I_2791 (I45951,I46037);
PAT_13 I_2792 (I45987,I46007,I45987,I45977,I46027,I46037,I45967,I45967,I46017,I45977,I45997,I46077,I46080,I46083,I46086,I46089,I46092,I46095,I46098,I46101,I1892,I1899);
OUT_INSTANCE I_2793 (I46077,I46117);
OUT_INSTANCE I_2794 (I46080,I46127);
OUT_INSTANCE I_2795 (I46083,I46137);
OUT_INSTANCE I_2796 (I46086,I46147);
OUT_INSTANCE I_2797 (I46089,I46157);
OUT_INSTANCE I_2798 (I46092,I46167);
OUT_INSTANCE I_2799 (I46095,I46177);
OUT_INSTANCE I_2800 (I46098,I46187);
OUT_INSTANCE I_2801 (I46101,I46197);
PAT_11 I_2802 (I46117,I46157,I46167,I46137,I46127,I46197,I46127,I46187,I46147,I46117,I46177,I46237,I46240,I46243,I46246,I46249,I46252,I46255,I46258,I46261,I46264,I1892,I1899);
OUT_INSTANCE I_2803 (I46237,I46280);
OUT_INSTANCE I_2804 (I46240,I46290);
OUT_INSTANCE I_2805 (I46243,I46300);
OUT_INSTANCE I_2806 (I46246,I46310);
OUT_INSTANCE I_2807 (I46249,I46320);
OUT_INSTANCE I_2808 (I46252,I46330);
OUT_INSTANCE I_2809 (I46255,I46340);
OUT_INSTANCE I_2810 (I46258,I46350);
OUT_INSTANCE I_2811 (I46261,I46360);
OUT_INSTANCE I_2812 (I46264,I46370);
PAT_15 I_2813 (I46360,I46290,I46310,I46340,I46330,I46280,I46320,I46350,I46280,I46300,I46370,I46410,I46413,I46416,I46419,I46422,I46425,I46428,I46431,I46434,I1892,I1899);
OUT_INSTANCE I_2814 (I46410,I46450);
OUT_INSTANCE I_2815 (I46413,I46460);
OUT_INSTANCE I_2816 (I46416,I46470);
OUT_INSTANCE I_2817 (I46419,I46480);
OUT_INSTANCE I_2818 (I46422,I46490);
OUT_INSTANCE I_2819 (I46425,I46500);
OUT_INSTANCE I_2820 (I46428,I46510);
OUT_INSTANCE I_2821 (I46431,I46520);
OUT_INSTANCE I_2822 (I46434,I46530);
PAT_6 I_2823 (I46460,I46450,I46470,I46520,I46460,I46530,I46480,I46500,I46490,I46510,I46450,I46570,I46573,I46576,I46579,I46582,I46585,I46588,I46591,I46594,I46597,I1892,I1899);
OUT_INSTANCE I_2824 (I46570,I46613);
OUT_INSTANCE I_2825 (I46573,I46623);
OUT_INSTANCE I_2826 (I46576,I46633);
OUT_INSTANCE I_2827 (I46579,I46643);
OUT_INSTANCE I_2828 (I46582,I46653);
OUT_INSTANCE I_2829 (I46585,I46663);
OUT_INSTANCE I_2830 (I46588,I46673);
OUT_INSTANCE I_2831 (I46591,I46683);
OUT_INSTANCE I_2832 (I46594,I46693);
OUT_INSTANCE I_2833 (I46597,I46703);
PAT_15 I_2834 (I46673,I46643,I46683,I46693,I46663,I46703,I46613,I46633,I46613,I46623,I46653,I46743,I46746,I46749,I46752,I46755,I46758,I46761,I46764,I46767,I1892,I1899);
OUT_INSTANCE I_2835 (I46743,I46783);
OUT_INSTANCE I_2836 (I46746,I46793);
OUT_INSTANCE I_2837 (I46749,I46803);
OUT_INSTANCE I_2838 (I46752,I46813);
OUT_INSTANCE I_2839 (I46755,I46823);
OUT_INSTANCE I_2840 (I46758,I46833);
OUT_INSTANCE I_2841 (I46761,I46843);
OUT_INSTANCE I_2842 (I46764,I46853);
OUT_INSTANCE I_2843 (I46767,I46863);
PAT_8 I_2844 (I46853,I46783,I46783,I46813,I46803,I46793,I46843,I46833,I46793,I46863,I46823,I46903,I46906,I46909,I46912,I46915,I46918,I46921,I46924,I46927,I1892,I1899);
OUT_INSTANCE I_2845 (I46903,I46943);
OUT_INSTANCE I_2846 (I46906,I46953);
OUT_INSTANCE I_2847 (I46909,I46963);
OUT_INSTANCE I_2848 (I46912,I46973);
OUT_INSTANCE I_2849 (I46915,I46983);
OUT_INSTANCE I_2850 (I46918,I46993);
OUT_INSTANCE I_2851 (I46921,I47003);
OUT_INSTANCE I_2852 (I46924,I47013);
OUT_INSTANCE I_2853 (I46927,I47023);
PAT_10 I_2854 (I46963,I46943,I46953,I47023,I47003,I46953,I46983,I46943,I47013,I46993,I46973,I47063,I47066,I47069,I47072,I47075,I47078,I47081,I47084,I1892,I1899);
OUT_INSTANCE I_2855 (I47063,I47100);
OUT_INSTANCE I_2856 (I47066,I47110);
OUT_INSTANCE I_2857 (I47069,I47120);
OUT_INSTANCE I_2858 (I47072,I47130);
OUT_INSTANCE I_2859 (I47075,I47140);
OUT_INSTANCE I_2860 (I47078,I47150);
OUT_INSTANCE I_2861 (I47081,I47160);
OUT_INSTANCE I_2862 (I47084,I47170);
PAT_15 I_2863 (I47150,I47160,I47120,I47140,I47100,I47100,I47120,I47170,I47130,I47110,I47110,I47210,I47213,I47216,I47219,I47222,I47225,I47228,I47231,I47234,I1892,I1899);
OUT_INSTANCE I_2864 (I47210,I47250);
OUT_INSTANCE I_2865 (I47213,I47260);
OUT_INSTANCE I_2866 (I47216,I47270);
OUT_INSTANCE I_2867 (I47219,I47280);
OUT_INSTANCE I_2868 (I47222,I47290);
OUT_INSTANCE I_2869 (I47225,I47300);
OUT_INSTANCE I_2870 (I47228,I47310);
OUT_INSTANCE I_2871 (I47231,I47320);
OUT_INSTANCE I_2872 (I47234,I47330);
PAT_10 I_2873 (I47260,I47290,I47270,I47250,I47320,I47330,I47280,I47250,I47260,I47310,I47300,I47370,I47373,I47376,I47379,I47382,I47385,I47388,I47391,I1892,I1899);
OUT_INSTANCE I_2874 (I47370,I47407);
OUT_INSTANCE I_2875 (I47373,I47417);
OUT_INSTANCE I_2876 (I47376,I47427);
OUT_INSTANCE I_2877 (I47379,I47437);
OUT_INSTANCE I_2878 (I47382,I47447);
OUT_INSTANCE I_2879 (I47385,I47457);
OUT_INSTANCE I_2880 (I47388,I47467);
OUT_INSTANCE I_2881 (I47391,I47477);
PAT_6 I_2882 (I47477,I47457,I47437,I47417,I47407,I47427,I47407,I47427,I47417,I47447,I47467,I47517,I47520,I47523,I47526,I47529,I47532,I47535,I47538,I47541,I47544,I1892,I1899);
OUT_INSTANCE I_2883 (I47517,I47560);
OUT_INSTANCE I_2884 (I47520,I47570);
OUT_INSTANCE I_2885 (I47523,I47580);
OUT_INSTANCE I_2886 (I47526,I47590);
OUT_INSTANCE I_2887 (I47529,I47600);
OUT_INSTANCE I_2888 (I47532,I47610);
OUT_INSTANCE I_2889 (I47535,I47620);
OUT_INSTANCE I_2890 (I47538,I47630);
OUT_INSTANCE I_2891 (I47541,I47640);
OUT_INSTANCE I_2892 (I47544,I47650);
PAT_10 I_2893 (I47560,I47610,I47620,I47590,I47560,I47640,I47650,I47570,I47600,I47580,I47630,I47690,I47693,I47696,I47699,I47702,I47705,I47708,I47711,I1892,I1899);
OUT_INSTANCE I_2894 (I47690,I47727);
OUT_INSTANCE I_2895 (I47693,I47737);
OUT_INSTANCE I_2896 (I47696,I47747);
OUT_INSTANCE I_2897 (I47699,I47757);
OUT_INSTANCE I_2898 (I47702,I47767);
OUT_INSTANCE I_2899 (I47705,I47777);
OUT_INSTANCE I_2900 (I47708,I47787);
OUT_INSTANCE I_2901 (I47711,I47797);
PAT_1 I_2902 (I47747,I47747,I47777,I47727,I47767,I47737,I47787,I47727,I47797,I47757,I47737,I47837,I47840,I47843,I47846,I47849,I47852,I47855,I47858,I47861,I1892,I1899);
OUT_INSTANCE I_2903 (I47837,I47877);
OUT_INSTANCE I_2904 (I47840,I47887);
OUT_INSTANCE I_2905 (I47843,I47897);
OUT_INSTANCE I_2906 (I47846,I47907);
OUT_INSTANCE I_2907 (I47849,I47917);
OUT_INSTANCE I_2908 (I47852,I47927);
OUT_INSTANCE I_2909 (I47855,I47937);
OUT_INSTANCE I_2910 (I47858,I47947);
OUT_INSTANCE I_2911 (I47861,I47957);
PAT_7 I_2912 (I47887,I47907,I47897,I47917,I47937,I47927,I47957,I47947,I47887,I47877,I47877,I47997,I48000,I48003,I48006,I48009,I48012,I48015,I48018,I48021,I1892,I1899);
OUT_INSTANCE I_2913 (I47997,I48037);
OUT_INSTANCE I_2914 (I48000,I48047);
OUT_INSTANCE I_2915 (I48003,I48057);
OUT_INSTANCE I_2916 (I48006,I48067);
OUT_INSTANCE I_2917 (I48009,I48077);
OUT_INSTANCE I_2918 (I48012,I48087);
OUT_INSTANCE I_2919 (I48015,I48097);
OUT_INSTANCE I_2920 (I48018,I48107);
OUT_INSTANCE I_2921 (I48021,I48117);
PAT_6 I_2922 (I48037,I48097,I48037,I48067,I48087,I48047,I48107,I48057,I48117,I48047,I48077,I48157,I48160,I48163,I48166,I48169,I48172,I48175,I48178,I48181,I48184,I1892,I1899);
OUT_INSTANCE I_2923 (I48157,I48200);
OUT_INSTANCE I_2924 (I48160,I48210);
OUT_INSTANCE I_2925 (I48163,I48220);
OUT_INSTANCE I_2926 (I48166,I48230);
OUT_INSTANCE I_2927 (I48169,I48240);
OUT_INSTANCE I_2928 (I48172,I48250);
OUT_INSTANCE I_2929 (I48175,I48260);
OUT_INSTANCE I_2930 (I48178,I48270);
OUT_INSTANCE I_2931 (I48181,I48280);
OUT_INSTANCE I_2932 (I48184,I48290);
PAT_5 I_2933 (I48270,I48200,I48220,I48230,I48250,I48260,I48200,I48280,I48210,I48240,I48290,I48330,I48333,I48336,I48339,I48342,I48345,I48348,I48351,I48354,I48357,I1892,I1899);
OUT_INSTANCE I_2934 (I48330,I48373);
OUT_INSTANCE I_2935 (I48333,I48383);
OUT_INSTANCE I_2936 (I48336,I48393);
OUT_INSTANCE I_2937 (I48339,I48403);
OUT_INSTANCE I_2938 (I48342,I48413);
OUT_INSTANCE I_2939 (I48345,I48423);
OUT_INSTANCE I_2940 (I48348,I48433);
OUT_INSTANCE I_2941 (I48351,I48443);
OUT_INSTANCE I_2942 (I48354,I48453);
OUT_INSTANCE I_2943 (I48357,I48463);
PAT_13 I_2944 (I48393,I48423,I48373,I48383,I48453,I48403,I48443,I48373,I48433,I48463,I48413,I48503,I48506,I48509,I48512,I48515,I48518,I48521,I48524,I48527,I1892,I1899);
OUT_INSTANCE I_2945 (I48503,I48543);
OUT_INSTANCE I_2946 (I48506,I48553);
OUT_INSTANCE I_2947 (I48509,I48563);
OUT_INSTANCE I_2948 (I48512,I48573);
OUT_INSTANCE I_2949 (I48515,I48583);
OUT_INSTANCE I_2950 (I48518,I48593);
OUT_INSTANCE I_2951 (I48521,I48603);
OUT_INSTANCE I_2952 (I48524,I48613);
OUT_INSTANCE I_2953 (I48527,I48623);
PAT_10 I_2954 (I48613,I48593,I48573,I48553,I48623,I48553,I48583,I48543,I48543,I48603,I48563,I48663,I48666,I48669,I48672,I48675,I48678,I48681,I48684,I1892,I1899);
OUT_INSTANCE I_2955 (I48663,I48700);
OUT_INSTANCE I_2956 (I48666,I48710);
OUT_INSTANCE I_2957 (I48669,I48720);
OUT_INSTANCE I_2958 (I48672,I48730);
OUT_INSTANCE I_2959 (I48675,I48740);
OUT_INSTANCE I_2960 (I48678,I48750);
OUT_INSTANCE I_2961 (I48681,I48760);
OUT_INSTANCE I_2962 (I48684,I48770);
PAT_6 I_2963 (I48770,I48750,I48730,I48710,I48700,I48720,I48700,I48720,I48710,I48740,I48760,I48810,I48813,I48816,I48819,I48822,I48825,I48828,I48831,I48834,I48837,I1892,I1899);
OUT_INSTANCE I_2964 (I48810,I48853);
OUT_INSTANCE I_2965 (I48813,I48863);
OUT_INSTANCE I_2966 (I48816,I48873);
OUT_INSTANCE I_2967 (I48819,I48883);
OUT_INSTANCE I_2968 (I48822,I48893);
OUT_INSTANCE I_2969 (I48825,I48903);
OUT_INSTANCE I_2970 (I48828,I48913);
OUT_INSTANCE I_2971 (I48831,I48923);
OUT_INSTANCE I_2972 (I48834,I48933);
OUT_INSTANCE I_2973 (I48837,I48943);
PAT_4 I_2974 (I48853,I48903,I48863,I48873,I48883,I48853,I48943,I48913,I48923,I48893,I48933,I48983,I48986,I48989,I48992,I48995,I48998,I49001,I49004,I49007,I1892,I1899);
OUT_INSTANCE I_2975 (I48983,I49023);
OUT_INSTANCE I_2976 (I48986,I49033);
OUT_INSTANCE I_2977 (I48989,I49043);
OUT_INSTANCE I_2978 (I48992,I49053);
OUT_INSTANCE I_2979 (I48995,I49063);
OUT_INSTANCE I_2980 (I48998,I49073);
OUT_INSTANCE I_2981 (I49001,I49083);
OUT_INSTANCE I_2982 (I49004,I49093);
OUT_INSTANCE I_2983 (I49007,I49103);
PAT_10 I_2984 (I49023,I49023,I49103,I49033,I49053,I49083,I49073,I49033,I49093,I49043,I49063,I49143,I49146,I49149,I49152,I49155,I49158,I49161,I49164,I1892,I1899);
OUT_INSTANCE I_2985 (I49143,I49180);
OUT_INSTANCE I_2986 (I49146,I49190);
OUT_INSTANCE I_2987 (I49149,I49200);
OUT_INSTANCE I_2988 (I49152,I49210);
OUT_INSTANCE I_2989 (I49155,I49220);
OUT_INSTANCE I_2990 (I49158,I49230);
OUT_INSTANCE I_2991 (I49161,I49240);
OUT_INSTANCE I_2992 (I49164,I49250);
PAT_6 I_2993 (I49250,I49230,I49210,I49190,I49180,I49200,I49180,I49200,I49190,I49220,I49240,I49290,I49293,I49296,I49299,I49302,I49305,I49308,I49311,I49314,I49317,I1892,I1899);
OUT_INSTANCE I_2994 (I49290,I49333);
OUT_INSTANCE I_2995 (I49293,I49343);
OUT_INSTANCE I_2996 (I49296,I49353);
OUT_INSTANCE I_2997 (I49299,I49363);
OUT_INSTANCE I_2998 (I49302,I49373);
OUT_INSTANCE I_2999 (I49305,I49383);
OUT_INSTANCE I_3000 (I49308,I49393);
OUT_INSTANCE I_3001 (I49311,I49403);
OUT_INSTANCE I_3002 (I49314,I49413);
OUT_INSTANCE I_3003 (I49317,I49423);
PAT_15 I_3004 (I49393,I49363,I49403,I49413,I49383,I49423,I49333,I49353,I49333,I49343,I49373,I49463,I49466,I49469,I49472,I49475,I49478,I49481,I49484,I49487,I1892,I1899);
OUT_INSTANCE I_3005 (I49463,I49503);
OUT_INSTANCE I_3006 (I49466,I49513);
OUT_INSTANCE I_3007 (I49469,I49523);
OUT_INSTANCE I_3008 (I49472,I49533);
OUT_INSTANCE I_3009 (I49475,I49543);
OUT_INSTANCE I_3010 (I49478,I49553);
OUT_INSTANCE I_3011 (I49481,I49563);
OUT_INSTANCE I_3012 (I49484,I49573);
OUT_INSTANCE I_3013 (I49487,I49583);
PAT_4 I_3014 (I49543,I49563,I49503,I49513,I49523,I49503,I49583,I49573,I49533,I49553,I49513,I49623,I49626,I49629,I49632,I49635,I49638,I49641,I49644,I49647,I1892,I1899);
OUT_INSTANCE I_3015 (I49623,I49663);
OUT_INSTANCE I_3016 (I49626,I49673);
OUT_INSTANCE I_3017 (I49629,I49683);
OUT_INSTANCE I_3018 (I49632,I49693);
OUT_INSTANCE I_3019 (I49635,I49703);
OUT_INSTANCE I_3020 (I49638,I49713);
OUT_INSTANCE I_3021 (I49641,I49723);
OUT_INSTANCE I_3022 (I49644,I49733);
OUT_INSTANCE I_3023 (I49647,I49743);
PAT_6 I_3024 (I49663,I49683,I49673,I49713,I49723,I49703,I49743,I49733,I49663,I49693,I49673,I49783,I49786,I49789,I49792,I49795,I49798,I49801,I49804,I49807,I49810,I1892,I1899);
OUT_INSTANCE I_3025 (I49783,I49826);
OUT_INSTANCE I_3026 (I49786,I49836);
OUT_INSTANCE I_3027 (I49789,I49846);
OUT_INSTANCE I_3028 (I49792,I49856);
OUT_INSTANCE I_3029 (I49795,I49866);
OUT_INSTANCE I_3030 (I49798,I49876);
OUT_INSTANCE I_3031 (I49801,I49886);
OUT_INSTANCE I_3032 (I49804,I49896);
OUT_INSTANCE I_3033 (I49807,I49906);
OUT_INSTANCE I_3034 (I49810,I49916);
PAT_17 I_3035 (I49866,I49876,I49896,I49856,I49836,I49906,I49886,I49826,I49916,I49846,I49826,I49956,I49959,I49962,I49965,I49968,I49971,I49974,I49977,I49980,I49983,I1892,I1899);
OUT_INSTANCE I_3036 (I49956,I49999);
OUT_INSTANCE I_3037 (I49959,I50009);
OUT_INSTANCE I_3038 (I49962,I50019);
OUT_INSTANCE I_3039 (I49965,I50029);
OUT_INSTANCE I_3040 (I49968,I50039);
OUT_INSTANCE I_3041 (I49971,I50049);
OUT_INSTANCE I_3042 (I49974,I50059);
OUT_INSTANCE I_3043 (I49977,I50069);
OUT_INSTANCE I_3044 (I49980,I50079);
OUT_INSTANCE I_3045 (I49983,I50089);
PAT_5 I_3046 (I50039,I50019,I50009,I50079,I50029,I50049,I50059,I49999,I49999,I50069,I50089,I50129,I50132,I50135,I50138,I50141,I50144,I50147,I50150,I50153,I50156,I1892,I1899);
OUT_INSTANCE I_3047 (I50129,I50172);
OUT_INSTANCE I_3048 (I50132,I50182);
OUT_INSTANCE I_3049 (I50135,I50192);
OUT_INSTANCE I_3050 (I50138,I50202);
OUT_INSTANCE I_3051 (I50141,I50212);
OUT_INSTANCE I_3052 (I50144,I50222);
OUT_INSTANCE I_3053 (I50147,I50232);
OUT_INSTANCE I_3054 (I50150,I50242);
OUT_INSTANCE I_3055 (I50153,I50252);
OUT_INSTANCE I_3056 (I50156,I50262);
endmodule


