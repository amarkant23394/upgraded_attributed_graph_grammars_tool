module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_5_r_7,n6_7,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_5_r_7,n6_7,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N1371_0_r_7,n53_7,n52_7);
nor I_41(N1508_0_r_7,n51_7,n52_7);
nand I_42(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_43(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_44(n_576_5_r_7,n31_7,n32_7);
nor I_45(n_102_5_r_7,N1371_0_r_16,n_572_7_r_16);
nand I_46(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_47(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_48(n_572_7_r_7,n54_7,n33_7);
nand I_49(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_50(n_549_7_r_7,n53_7,n36_7);
nand I_51(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_52(n_452_7_r_7,N1372_1_r_16,n_569_7_r_16);
nor I_53(n4_7_l_7,N1508_1_r_16,N6147_2_r_16);
not I_54(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_55(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_56(n30_7,n53_7);
and I_57(N3_8_l_7,n50_7,N1507_6_r_16);
DFFARX1 I_58(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_59(n_431_5_r_7,n40_7,n41_7);
nor I_60(n4_7_r_7,n54_7,n49_7);
and I_61(n31_7,n_102_5_r_7,n39_7);
not I_62(n32_7,N1508_1_r_16);
nor I_63(n33_7,n34_7,n_452_7_r_16);
and I_64(n34_7,n35_7,N1508_0_r_16);
not I_65(n35_7,N1371_0_r_16);
nor I_66(n36_7,n37_7,N1508_1_r_16);
or I_67(n37_7,n54_7,N1371_0_r_16);
or I_68(n38_7,N1508_6_r_16,G42_7_r_16);
nor I_69(n39_7,n_452_7_r_7,N1508_0_r_16);
nand I_70(n40_7,n46_7,n47_7);
nand I_71(n41_7,n42_7,n43_7);
nor I_72(n42_7,n44_7,n45_7);
nor I_73(n43_7,N1508_6_r_16,G42_7_r_16);
nor I_74(n44_7,n_573_7_r_16,N1371_0_r_16);
nor I_75(n45_7,n_572_7_r_16,n_452_7_r_16);
nand I_76(n46_7,n35_7,N1508_0_r_16);
not I_77(n47_7,n_452_7_r_16);
or I_78(n48_7,n_452_7_r_7,N1508_0_r_16);
not I_79(n49_7,n_452_7_r_7);
nand I_80(n50_7,N1508_6_r_16,N1372_1_r_16);
and I_81(n51_7,n_452_7_r_7,n45_7);
not I_82(n52_7,n44_7);
endmodule


