module test_I2914(I2005,I1316,I2798,I1294,I2488,I2070,I1301,I1917,I1988,I2914);
input I2005,I1316,I2798,I1294,I2488,I2070,I1301,I1917,I1988;
output I2914;
wire I2668,I1911,I1914,I2583,I2313,I2022,I2897,I2600,I2849,I2832,I2344,I2651,I2685,I2815,I1923;
nand I_0(I2668,I2651,I1914);
nand I_1(I1911,I2070,I2488);
DFFARX1 I_2(I1294,,,I1914,);
not I_3(I2583,I1301);
DFFARX1 I_4(I1294,,,I2313,);
nand I_5(I2022,I2005,I1316);
nand I_6(I2897,I2600,I1923);
not I_7(I2600,I1911);
nor I_8(I2849,I2832,I2685);
DFFARX1 I_9(I2815,I1294,I2583,,,I2832,);
nor I_10(I2344,I2313,I1988);
nor I_11(I2651,I2600);
not I_12(I2685,I2668);
and I_13(I2914,I2897,I2849);
or I_14(I2815,I2798,I1917);
nand I_15(I1923,I2022,I2344);
endmodule


