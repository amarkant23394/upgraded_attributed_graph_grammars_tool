module test_I13860(I1477,I12024,I12041,I10026,I11953,I12106,I12524,I1470,I13860);
input I1477,I12024,I12041,I10026,I11953,I12106,I12524,I1470;
output I13860;
wire I13792,I12058,I12380,I13775,I13843,I11965,I11947,I12287,I12349,I13809,I13826,I12304,I11973,I11959;
nor I_0(I13860,I13843,I13826);
nand I_1(I13792,I11953,I11965);
nand I_2(I12058,I12041,I10026);
nor I_3(I12380,I12349,I12024);
not I_4(I13775,I1477);
nor I_5(I13843,I11959,I11965);
DFFARX1 I_6(I12304,I1470,I11973,,,I11965,);
nand I_7(I11947,I12106,I12524);
nand I_8(I12287,I12024);
DFFARX1 I_9(I1470,I11973,,,I12349,);
and I_10(I13809,I13792,I11947);
DFFARX1 I_11(I13809,I1470,I13775,,,I13826,);
and I_12(I12304,I12106,I12287);
not I_13(I11973,I1477);
nand I_14(I11959,I12058,I12380);
endmodule


