module test_I10609(I9833,I1477,I9771,I1470,I10609);
input I9833,I1477,I9771,I1470;
output I10609;
wire I9477,I10647,I11105,I10698,I10766,I9468,I10681,I11009,I9456,I11088;
nor I_0(I9477,I9771,I9833);
not I_1(I10647,I1477);
and I_2(I11105,I10766,I11088);
nand I_3(I10698,I10681,I9456);
not I_4(I10766,I9477);
DFFARX1 I_5(I1470,,,I9468,);
nor I_6(I10681,I9477);
DFFARX1 I_7(I9468,I1470,I10647,,,I11009,);
DFFARX1 I_8(I1470,,,I9456,);
nand I_9(I11088,I11009,I10698);
DFFARX1 I_10(I11105,I1470,I10647,,,I10609,);
endmodule


