module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_7,n8_7,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_7,n8_7,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_7,n8_7,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_7,n8_7,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_7,n8_7,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_7,n8_7,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_34(n_572_1_r_7,n30_7,n31_7);
nand I_35(n_573_1_r_7,n28_7,n_573_1_r_13);
nor I_36(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_37(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_38(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_39(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_40(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_41(P6_5_r_7,P6_5_r_internal_7);
or I_42(n_431_0_l_7,n36_7,n_572_1_r_13);
not I_43(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_44(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_45(n27_7,n43_7);
DFFARX1 I_46(n_266_and_0_3_r_13,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_47(G42_1_r_13,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_48(n4_1_r_7,n30_7,n38_7);
nor I_49(N1_4_r_7,n27_7,n40_7);
nand I_50(n26_7,n39_7,n_572_1_r_13);
not I_51(n5_7,n_452_1_r_13);
DFFARX1 I_52(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_53(n28_7,n26_7,n29_7);
not I_54(n29_7,ACVQN1_5_r_13);
not I_55(n30_7,n_549_1_r_13);
nand I_56(n31_7,n27_7,n29_7);
nor I_57(n32_7,ACVQN1_5_l_7,n34_7);
nor I_58(n33_7,n29_7,n_452_1_r_13);
not I_59(n34_7,n_573_1_r_13);
nor I_60(n35_7,n43_7,n44_7);
and I_61(n36_7,n37_7,G42_1_r_13);
nor I_62(n37_7,n30_7,ACVQN2_3_r_13);
nand I_63(n38_7,n29_7,n_452_1_r_13);
nor I_64(n39_7,n_452_1_r_13,P6_5_r_13);
nor I_65(n40_7,n44_7,n41_7);
nor I_66(n41_7,n34_7,n42_7);
nand I_67(n42_7,n5_7,ACVQN1_5_r_13);
endmodule


