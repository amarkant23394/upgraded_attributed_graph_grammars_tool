module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_5_r_9,n10_9,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N6147_2_r_9,n62_9,n46_9);
not I_37(N1372_4_r_9,n59_9);
nor I_38(N1508_4_r_9,n58_9,n59_9);
nand I_39(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_40(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_41(n_576_5_r_9,n39_9,n40_9);
not I_42(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_43(n_547_5_r_9,n43_9,N1372_1_r_5);
and I_44(n_42_8_r_9,n44_9,N1371_0_r_5);
DFFARX1 I_45(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_46(N6147_9_r_9,n41_9,n45_9);
nor I_47(N6134_9_r_9,n45_9,n51_9);
nor I_48(I_BUFF_1_9_r_9,n41_9,N1372_1_r_5);
nor I_49(n4_7_l_9,N1371_0_r_5,N1508_1_r_5);
not I_50(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_51(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_52(N3_8_l_9,n57_9,N1507_6_r_5);
DFFARX1 I_53(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_54(n38_9,n63_9);
nor I_55(n_431_5_r_9,N1508_0_r_5,N1372_1_r_5);
nor I_56(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_57(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_58(n40_9,n41_9);
nand I_59(n41_9,G42_7_r_5,n_573_7_r_5);
nor I_60(n42_9,N1508_1_r_5,N6147_2_r_5);
nor I_61(n43_9,n63_9,n41_9);
nor I_62(n44_9,N6147_2_r_5,N1508_6_r_5);
and I_63(n45_9,n52_9,n_572_7_r_5);
nor I_64(n46_9,n47_9,n48_9);
nor I_65(n47_9,n49_9,n50_9);
not I_66(n48_9,n_429_or_0_5_r_9);
not I_67(n49_9,n42_9);
or I_68(n50_9,n63_9,n51_9);
nor I_69(n51_9,N1371_0_r_5,n_452_7_r_5);
nor I_70(n52_9,n49_9,N1372_1_r_5);
nor I_71(n53_9,n54_9,n55_9);
nor I_72(n54_9,n56_9,N1372_1_r_5);
or I_73(n55_9,n44_9,N1508_1_r_5);
not I_74(n56_9,n_572_7_r_5);
nand I_75(n57_9,n_569_7_r_5,n_452_7_r_5);
nor I_76(n58_9,n62_9,n60_9);
nand I_77(n59_9,n51_9,n61_9);
nor I_78(n60_9,n38_9,n44_9);
nor I_79(n61_9,N1508_6_r_5,N1371_0_r_5);
endmodule


