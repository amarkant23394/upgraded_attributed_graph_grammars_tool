module test_I2815(I1328,I1923,I2155,I1294,I1331,I1301,I2815);
input I1328,I1923,I2155,I1294,I1331,I1301;
output I2815;
wire I2172,I2764,I2798,I1917,I2781,I1905,I1899,I2313,I1937,I2505,I2389,I2406,I2488;
DFFARX1 I_0(I2155,I1294,I1937,,,I2172,);
or I_1(I2815,I2798,I1917);
not I_2(I2764,I1923);
and I_3(I2798,I2781,I1899);
nand I_4(I1917,I2406,I2505);
nor I_5(I2781,I2764,I1905);
DFFARX1 I_6(I2172,I1294,I1937,,,I1905,);
DFFARX1 I_7(I2172,I1294,I1937,,,I1899,);
DFFARX1 I_8(I1331,I1294,I1937,,,I2313,);
not I_9(I1937,I1301);
nor I_10(I2505,I2313,I2488);
DFFARX1 I_11(I1328,I1294,I1937,,,I2389,);
not I_12(I2406,I2389);
not I_13(I2488,I2406);
endmodule


