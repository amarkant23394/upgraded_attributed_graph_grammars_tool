module Benchmark_testing35000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2859,I2866,I7840,I7831,I7828,I7834,I7822,I7816,I7837,I7825,I7819,I53138,I53150,I53159,I53162,I53147,I53156,I53144,I53153,I53141,I72712,I72688,I72700,I72694,I72709,I72703,I72697,I72691,I72706,I82232,I82208,I82220,I82214,I82229,I82223,I82217,I82211,I82226,I84612,I84588,I84600,I84594,I84609,I84603,I84597,I84591,I84606,I224437,I224434,I224419,I224431,I224425,I224413,I224422,I224428,I224416,I240768,I240765,I240756,I240759,I240753,I240762,I240750,I240774,I240771,I263888,I263885,I263876,I263879,I263873,I263882,I263870,I263894,I263891,I287005,I287008,I286990,I286999,I287011,I287002,I286993,I286996,I287014,I315327,I315330,I315312,I315321,I315333,I315324,I315315,I315318,I315336,I345318,I345321,I345312,I345303,I345306,I345315,I345300,I345309,I412590,I412593,I412569,I412581,I412596,I412584,I412578,I412572,I412575,I412587,I430950,I430932,I430935,I430944,I430947,I430941,I430929,I430938,I487061,I487049,I487070,I487046,I487067,I487058,I487064,I487055,I487052,I503730,I503709,I503712,I503727,I503724,I503721,I503718,I503706,I503715,I504274,I504253,I504256,I504271,I504268,I504265,I504262,I504250,I504259,I550238,I550253,I550235,I550247,I550262,I550259,I550256,I550250,I550244,I550241);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2859,I2866;
output I7840,I7831,I7828,I7834,I7822,I7816,I7837,I7825,I7819,I53138,I53150,I53159,I53162,I53147,I53156,I53144,I53153,I53141,I72712,I72688,I72700,I72694,I72709,I72703,I72697,I72691,I72706,I82232,I82208,I82220,I82214,I82229,I82223,I82217,I82211,I82226,I84612,I84588,I84600,I84594,I84609,I84603,I84597,I84591,I84606,I224437,I224434,I224419,I224431,I224425,I224413,I224422,I224428,I224416,I240768,I240765,I240756,I240759,I240753,I240762,I240750,I240774,I240771,I263888,I263885,I263876,I263879,I263873,I263882,I263870,I263894,I263891,I287005,I287008,I286990,I286999,I287011,I287002,I286993,I286996,I287014,I315327,I315330,I315312,I315321,I315333,I315324,I315315,I315318,I315336,I345318,I345321,I345312,I345303,I345306,I345315,I345300,I345309,I412590,I412593,I412569,I412581,I412596,I412584,I412578,I412572,I412575,I412587,I430950,I430932,I430935,I430944,I430947,I430941,I430929,I430938,I487061,I487049,I487070,I487046,I487067,I487058,I487064,I487055,I487052,I503730,I503709,I503712,I503727,I503724,I503721,I503718,I503706,I503715,I504274,I504253,I504256,I504271,I504268,I504265,I504262,I504250,I504259,I550238,I550253,I550235,I550247,I550262,I550259,I550256,I550250,I550244,I550241;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2859,I2866,I2898,I43137,I2924,I2932,I43128,I2949,I2890,I43149,I2989,I2997,I3014,I43125,I3031,I3048,I3065,I2869,I3096,I3113,I3130,I43134,I2872,I3161,I3178,I43146,I3195,I43143,I3212,I3229,I3246,I2881,I3277,I43140,I3294,I3311,I2887,I3342,I2884,I3373,I43131,I3399,I3407,I3424,I2878,I2875,I3493,I309556,I3519,I3527,I309535,I3544,I3485,I309544,I3584,I3592,I3609,I309550,I3626,I309547,I3643,I3660,I3464,I3691,I3708,I3725,I309538,I309532,I3467,I3756,I3773,I309553,I3790,I3807,I3824,I3841,I3476,I3872,I309541,I3889,I3906,I3482,I3937,I3479,I3968,I3994,I4002,I4019,I3473,I3470,I4088,I163534,I4114,I4122,I163525,I4139,I4080,I163528,I4179,I4187,I4204,I163522,I4221,I163531,I4238,I4255,I4059,I4286,I4303,I4320,I163519,I163537,I4062,I4351,I4368,I4385,I163543,I4402,I4419,I4436,I4071,I4467,I163540,I4484,I4501,I4077,I4532,I4074,I4563,I163546,I4589,I4597,I4614,I4068,I4065,I4686,I120332,I4712,I4729,I4737,I4754,I120329,I120323,I4771,I120317,I4797,I4678,I4669,I120305,I4842,I4850,I120314,I4867,I4666,I120311,I4907,I4915,I4672,I4660,I4960,I120308,I120326,I4977,I5003,I5011,I4654,I5042,I5059,I120320,I5076,I5093,I5110,I4675,I5141,I4663,I4657,I5213,I474932,I5239,I5256,I5264,I5281,I474920,I474911,I5298,I474908,I5324,I5205,I5196,I474914,I5369,I5377,I474926,I5394,I5193,I474923,I5434,I5442,I5199,I5187,I5487,I474917,I5504,I474929,I5530,I5538,I5181,I5569,I5586,I5603,I5620,I5637,I5202,I5668,I5190,I5184,I5740,I176507,I5766,I5783,I5791,I5808,I176510,I5825,I176531,I5851,I5732,I5723,I176519,I5896,I5904,I176522,I5921,I5720,I176528,I5961,I5969,I5726,I5714,I6014,I176525,I176513,I6031,I176516,I6057,I6065,I5708,I6096,I6113,I176534,I6130,I6147,I6164,I5729,I6195,I5717,I5711,I6267,I150898,I6293,I6310,I6318,I6335,I150895,I150889,I6352,I150883,I6378,I6259,I6250,I150871,I6423,I6431,I150880,I6448,I6247,I150877,I6488,I6496,I6253,I6241,I6541,I150874,I150892,I6558,I6584,I6592,I6235,I6623,I6640,I150886,I6657,I6674,I6691,I6256,I6722,I6244,I6238,I6794,I520570,I6820,I6837,I6845,I6862,I520588,I520582,I6879,I520591,I6905,I6786,I6777,I520576,I6950,I6958,I520585,I6975,I6774,I520573,I7015,I7023,I6780,I6768,I7068,I520594,I520579,I7085,I7111,I7119,I6762,I7150,I7167,I7184,I7201,I7218,I6783,I7249,I6771,I6765,I7321,I172699,I7347,I7364,I7372,I7389,I172702,I7406,I172723,I7432,I7313,I7304,I172711,I7477,I7485,I172714,I7502,I7301,I172720,I7542,I7550,I7307,I7295,I7595,I172717,I172705,I7612,I172708,I7638,I7646,I7289,I7677,I7694,I172726,I7711,I7728,I7745,I7310,I7776,I7298,I7292,I7848,I295666,I7874,I7891,I7899,I7916,I295681,I295684,I7933,I295663,I7959,I295669,I8004,I8012,I295675,I8029,I8069,I8077,I8122,I295678,I295660,I8139,I295672,I8165,I8173,I8204,I8221,I8238,I8255,I8272,I8303,I8375,I77454,I8401,I8418,I8426,I8443,I77472,I77457,I8460,I77460,I8486,I8367,I8358,I77448,I8531,I8539,I77451,I8556,I8355,I77463,I8596,I8604,I8361,I8349,I8649,I77469,I77466,I8666,I8692,I8700,I8343,I8731,I8748,I8765,I8782,I8799,I8364,I8830,I8352,I8346,I8902,I568680,I8928,I8945,I8953,I8970,I568683,I568689,I8987,I568698,I9013,I8894,I8885,I568701,I9058,I9066,I568692,I9083,I8882,I9123,I9131,I8888,I8876,I9176,I568707,I568686,I9193,I568695,I9219,I9227,I8870,I9258,I9275,I568704,I9292,I9309,I9326,I8891,I9357,I8879,I8873,I9429,I510234,I9455,I9472,I9480,I9497,I510252,I510246,I9514,I510255,I9540,I9421,I9412,I510240,I9585,I9593,I510249,I9610,I9409,I510237,I9650,I9658,I9415,I9403,I9703,I510258,I510243,I9720,I9746,I9754,I9397,I9785,I9802,I9819,I9836,I9853,I9418,I9884,I9406,I9400,I9956,I567490,I9982,I9999,I10007,I10024,I567493,I567499,I10041,I567508,I10067,I9948,I9939,I567511,I10112,I10120,I567502,I10137,I9936,I10177,I10185,I9942,I9930,I10230,I567517,I567496,I10247,I567505,I10273,I10281,I9924,I10312,I10329,I567514,I10346,I10363,I10380,I9945,I10411,I9933,I9927,I10483,I485914,I10509,I10526,I10534,I10551,I485902,I485893,I10568,I485890,I10594,I10475,I10466,I485896,I10639,I10647,I485908,I10664,I10463,I485905,I10704,I10712,I10469,I10457,I10757,I485899,I10774,I485911,I10800,I10808,I10451,I10839,I10856,I10873,I10890,I10907,I10472,I10938,I10460,I10454,I11010,I155114,I11036,I11053,I11061,I11078,I155111,I155105,I11095,I155099,I11121,I11002,I10993,I155087,I11166,I11174,I155096,I11191,I10990,I155093,I11231,I11239,I10996,I10984,I11284,I155090,I155108,I11301,I11327,I11335,I10978,I11366,I11383,I155102,I11400,I11417,I11434,I10999,I11465,I10987,I10981,I11537,I233829,I11563,I11580,I11588,I11605,I233814,I233832,I11622,I233826,I11648,I11529,I11520,I233823,I11693,I11701,I11718,I11517,I233817,I11758,I11766,I11523,I11511,I11811,I233838,I233820,I11828,I233835,I11854,I11862,I11505,I11893,I11910,I11927,I11944,I11961,I11526,I11992,I11514,I11508,I12064,I190651,I12090,I12107,I12115,I12132,I190654,I12149,I190675,I12175,I12056,I12047,I190663,I12220,I12228,I190666,I12245,I12044,I190672,I12285,I12293,I12050,I12038,I12338,I190669,I190657,I12355,I190660,I12381,I12389,I12032,I12420,I12437,I190678,I12454,I12471,I12488,I12053,I12519,I12041,I12035,I12591,I12617,I12634,I12642,I12659,I12676,I12702,I12583,I12574,I12747,I12755,I12772,I12571,I12812,I12820,I12577,I12565,I12865,I12882,I12908,I12916,I12559,I12947,I12964,I12981,I12998,I13015,I12580,I13046,I12568,I12562,I13118,I97684,I13144,I13161,I13169,I13186,I97702,I97687,I13203,I97690,I13229,I13110,I13101,I97678,I13274,I13282,I97681,I13299,I13098,I97693,I13339,I13347,I13104,I13092,I13392,I97699,I97696,I13409,I13435,I13443,I13086,I13474,I13491,I13508,I13525,I13542,I13107,I13573,I13095,I13089,I13645,I400965,I13671,I13688,I13696,I13713,I400941,I400968,I13730,I400953,I13756,I13637,I13628,I400959,I13801,I13809,I400944,I13826,I13625,I400962,I13866,I13874,I13631,I13619,I13919,I400947,I400950,I13936,I13962,I13970,I13613,I14001,I14018,I400956,I14035,I14052,I14069,I13634,I14100,I13622,I13616,I14172,I164600,I14198,I14215,I14223,I14240,I164597,I164591,I14257,I164585,I14283,I14164,I14155,I164573,I14328,I14336,I164582,I14353,I14152,I164579,I14393,I14401,I14158,I14146,I14446,I164576,I164594,I14463,I14489,I14497,I14140,I14528,I14545,I164588,I14562,I14579,I14596,I14161,I14627,I14149,I14143,I14699,I138777,I14725,I14742,I14750,I14767,I138774,I138768,I14784,I138762,I14810,I14691,I14682,I138750,I14855,I14863,I138759,I14880,I14679,I138756,I14920,I14928,I14685,I14673,I14973,I138753,I138771,I14990,I15016,I15024,I14667,I15055,I15072,I138765,I15089,I15106,I15123,I14688,I15154,I14676,I14670,I15226,I555590,I15252,I15269,I15277,I15294,I555593,I555599,I15311,I555608,I15337,I15218,I15209,I555611,I15382,I15390,I555602,I15407,I15206,I15447,I15455,I15212,I15200,I15500,I555617,I555596,I15517,I555605,I15543,I15551,I15194,I15582,I15599,I555614,I15616,I15633,I15650,I15215,I15681,I15203,I15197,I15753,I363754,I15779,I15796,I15804,I15821,I363745,I363766,I15838,I363748,I15864,I15745,I15736,I15909,I15917,I363763,I15934,I15733,I363757,I15974,I15982,I15739,I15727,I16027,I363751,I363760,I16044,I16070,I16078,I15721,I16109,I16126,I16143,I16160,I16177,I15742,I16208,I15730,I15724,I16280,I167803,I16306,I16323,I16331,I16348,I167806,I16365,I167827,I16391,I16272,I16263,I167815,I16436,I16444,I167818,I16461,I16260,I167824,I16501,I16509,I16266,I16254,I16554,I167821,I167809,I16571,I167812,I16597,I16605,I16248,I16636,I16653,I167830,I16670,I16687,I16704,I16269,I16735,I16257,I16251,I16807,I212522,I16833,I16850,I16858,I16875,I212528,I212516,I16892,I212513,I16918,I16799,I16790,I212525,I16963,I16971,I212519,I16988,I16787,I212537,I17028,I17036,I16793,I16781,I17081,I212531,I212534,I17098,I17124,I17132,I16775,I17163,I17180,I17197,I17214,I17231,I16796,I17262,I16784,I16778,I17334,I433740,I17360,I17377,I17385,I17402,I433734,I433755,I17419,I17445,I17326,I17317,I433737,I17490,I17498,I433746,I17515,I17314,I17555,I17563,I17320,I17308,I17608,I433752,I17625,I433743,I17651,I17659,I17302,I17690,I17707,I433749,I17724,I17741,I17758,I17323,I17789,I17311,I17305,I17861,I146682,I17887,I17904,I17912,I17929,I146679,I146673,I17946,I146667,I17972,I17853,I17844,I146655,I18017,I18025,I146664,I18042,I17841,I146661,I18082,I18090,I17847,I17835,I18135,I146658,I146676,I18152,I18178,I18186,I17829,I18217,I18234,I146670,I18251,I18268,I18285,I17850,I18316,I17838,I17832,I18388,I319364,I18414,I18431,I18439,I18456,I319379,I319382,I18473,I319361,I18499,I18380,I18371,I319367,I18544,I18552,I319373,I18569,I18368,I18609,I18617,I18374,I18362,I18662,I319376,I319358,I18679,I319370,I18705,I18713,I18356,I18744,I18761,I18778,I18795,I18812,I18377,I18843,I18365,I18359,I18915,I433179,I18941,I18958,I18966,I18983,I433173,I433194,I19000,I19026,I18907,I18898,I433176,I19071,I19079,I433185,I19096,I18895,I19136,I19144,I18901,I18889,I19189,I433191,I19206,I433182,I19232,I19240,I18883,I19271,I19288,I433188,I19305,I19322,I19339,I18904,I19370,I18892,I18886,I19442,I279482,I19468,I19485,I19493,I19510,I279497,I279500,I19527,I279479,I19553,I19434,I19425,I279485,I19598,I19606,I279491,I19623,I19422,I19663,I19671,I19428,I19416,I19716,I279494,I279476,I19733,I279488,I19759,I19767,I19410,I19798,I19815,I19832,I19849,I19866,I19431,I19897,I19419,I19413,I19969,I202619,I19995,I20012,I20020,I20037,I202622,I20054,I202643,I20080,I19961,I19952,I202631,I20125,I20133,I202634,I20150,I19949,I202640,I20190,I20198,I19955,I19943,I20243,I202637,I202625,I20260,I202628,I20286,I20294,I19937,I20325,I20342,I202646,I20359,I20376,I20393,I19958,I20424,I19946,I19940,I20496,I502074,I20522,I20539,I20547,I20564,I502092,I502086,I20581,I502095,I20607,I20488,I20479,I502080,I20652,I20660,I502089,I20677,I20476,I502077,I20717,I20725,I20482,I20470,I20770,I502098,I502083,I20787,I20813,I20821,I20464,I20852,I20869,I20886,I20903,I20920,I20485,I20951,I20473,I20467,I21023,I62585,I21049,I21057,I21074,I62579,I62573,I21091,I62594,I21117,I62591,I21134,I21142,I62588,I21159,I20991,I21190,I21207,I21003,I21247,I21012,I21269,I62576,I21286,I62597,I21312,I21329,I21015,I21351,I21000,I21382,I62582,I21399,I21416,I21433,I21009,I21464,I20997,I21006,I20994,I21550,I459886,I21576,I21584,I21601,I459901,I459880,I21618,I459883,I21644,I459904,I21661,I21669,I21686,I21518,I21717,I21734,I21530,I21774,I21539,I21796,I459892,I459889,I21813,I459895,I21839,I21856,I21542,I21878,I21527,I21909,I459898,I21926,I21943,I21960,I21536,I21991,I21524,I21533,I21521,I22077,I91740,I22103,I22111,I22128,I91734,I91728,I22145,I91749,I22171,I91746,I22188,I22196,I91743,I22213,I22045,I22244,I22261,I22057,I22301,I22066,I22323,I91731,I22340,I91752,I22366,I22383,I22069,I22405,I22054,I22436,I91737,I22453,I22470,I22487,I22063,I22518,I22051,I22060,I22048,I22604,I70915,I22630,I22638,I22655,I70909,I70903,I22672,I70924,I22698,I70921,I22715,I22723,I70918,I22740,I22572,I22771,I22788,I22584,I22828,I22593,I22850,I70906,I22867,I70927,I22893,I22910,I22596,I22932,I22581,I22963,I70912,I22980,I22997,I23014,I22590,I23045,I22578,I22587,I22575,I23131,I265038,I23157,I23165,I23182,I265029,I265047,I23199,I265026,I23225,I23242,I23250,I265032,I23267,I23099,I23298,I23315,I23111,I23355,I23120,I23377,I265044,I265035,I23394,I265050,I23420,I23437,I23123,I23459,I23108,I23490,I265041,I23507,I23524,I23541,I23117,I23572,I23105,I23114,I23102,I23658,I222036,I23684,I23692,I23709,I222057,I222051,I23726,I222033,I23752,I23769,I23777,I222045,I23794,I23626,I23825,I23842,I23638,I222042,I23882,I23647,I23904,I222048,I222039,I23921,I23947,I23964,I23650,I23986,I23635,I24017,I222054,I24034,I24051,I24068,I23644,I24099,I23632,I23641,I23629,I24185,I514048,I24211,I24219,I24236,I514042,I514063,I24253,I514054,I24279,I514045,I24296,I24304,I514057,I24321,I24153,I24352,I24369,I24165,I24409,I24174,I24431,I514066,I514051,I24448,I24474,I24491,I24177,I24513,I24162,I24544,I514060,I24561,I24578,I24595,I24171,I24626,I24159,I24168,I24156,I24712,I102450,I24738,I24746,I24763,I102444,I102438,I24780,I102459,I24806,I102456,I24823,I24831,I102453,I24848,I24680,I24879,I24896,I24692,I24936,I24701,I24958,I102441,I24975,I102462,I25001,I25018,I24704,I25040,I24689,I25071,I102447,I25088,I25105,I25122,I24698,I25153,I24686,I24695,I24683,I25239,I25265,I25273,I25290,I25307,I25333,I25350,I25358,I25375,I25207,I25406,I25423,I25219,I25463,I25228,I25485,I25502,I25528,I25545,I25231,I25567,I25216,I25598,I25615,I25632,I25649,I25225,I25680,I25213,I25222,I25210,I25766,I366916,I25792,I25800,I25817,I366913,I366928,I25834,I366910,I25860,I366907,I25877,I25885,I25902,I25734,I25933,I25950,I25746,I25990,I25755,I26012,I366922,I26029,I366925,I26055,I26072,I25758,I26094,I25743,I26125,I366919,I26142,I26159,I26176,I25752,I26207,I25740,I25749,I25737,I26293,I373767,I26319,I26327,I26344,I373764,I373779,I26361,I373761,I26387,I373758,I26404,I26412,I26429,I26261,I26460,I26477,I26273,I26517,I26282,I26539,I373773,I26556,I373776,I26582,I26599,I26285,I26621,I26270,I26652,I373770,I26669,I26686,I26703,I26279,I26734,I26267,I26276,I26264,I26820,I535564,I26846,I26854,I26871,I535570,I535588,I26888,I535585,I26914,I535582,I26931,I26939,I535576,I26956,I26788,I26987,I27004,I26800,I27044,I26809,I27066,I535579,I535567,I27083,I535591,I27109,I27126,I26812,I27148,I26797,I27179,I535573,I27196,I27213,I27230,I26806,I27261,I26794,I26803,I26791,I27347,I83410,I27373,I27381,I27398,I83404,I83398,I27415,I83419,I27441,I83416,I27458,I27466,I83413,I27483,I27315,I27514,I27531,I27327,I27571,I27336,I27593,I83401,I27610,I83422,I27636,I27653,I27339,I27675,I27324,I27706,I83407,I27723,I27740,I27757,I27333,I27788,I27321,I27330,I27318,I27874,I544297,I27900,I27908,I27925,I544291,I544312,I27942,I544288,I27968,I544309,I27985,I27993,I544306,I28010,I27842,I28041,I28058,I27854,I544294,I28098,I27863,I28120,I544303,I544300,I28137,I544285,I28163,I28180,I27866,I28202,I27851,I28233,I28250,I28267,I28284,I27860,I28315,I27848,I27857,I27845,I28401,I115589,I28427,I28435,I28452,I115571,I115586,I28469,I115562,I28495,I115565,I28512,I28520,I115580,I28537,I28369,I28568,I28585,I28381,I115583,I28625,I28390,I28647,I115574,I28664,I115568,I28690,I28707,I28393,I28729,I28378,I28760,I115577,I28777,I28794,I28811,I28387,I28842,I28375,I28384,I28372,I28928,I306654,I28954,I28962,I28979,I306645,I306663,I28996,I306642,I29022,I29039,I29047,I306648,I29064,I28896,I29095,I29112,I28908,I29152,I28917,I29174,I306660,I306651,I29191,I306666,I29217,I29234,I28920,I29256,I28905,I29287,I306657,I29304,I29321,I29338,I28914,I29369,I28902,I28911,I28899,I29455,I121386,I29481,I29489,I29506,I121368,I121383,I29523,I121359,I29549,I121362,I29566,I29574,I121377,I29591,I29423,I29622,I29639,I29435,I121380,I29679,I29444,I29701,I121371,I29718,I121365,I29744,I29761,I29447,I29783,I29432,I29814,I121374,I29831,I29848,I29865,I29441,I29896,I29429,I29438,I29426,I29982,I127710,I30008,I30016,I30033,I127692,I127707,I30050,I127683,I30076,I127686,I30093,I30101,I127701,I30118,I29950,I30149,I30166,I29962,I127704,I30206,I29971,I30228,I127695,I30245,I127689,I30271,I30288,I29974,I30310,I29959,I30341,I127698,I30358,I30375,I30392,I29968,I30423,I29956,I29965,I29953,I30509,I314168,I30535,I30543,I30560,I314159,I314177,I30577,I314156,I30603,I30620,I30628,I314162,I30645,I30477,I30676,I30693,I30489,I30733,I30498,I30755,I314174,I314165,I30772,I314180,I30798,I30815,I30501,I30837,I30486,I30868,I314171,I30885,I30902,I30919,I30495,I30950,I30483,I30492,I30480,I31036,I468556,I31062,I31070,I31087,I468571,I468550,I31104,I468553,I31130,I468574,I31147,I31155,I31172,I31004,I31203,I31220,I31016,I31260,I31025,I31282,I468562,I468559,I31299,I468565,I31325,I31342,I31028,I31364,I31013,I31395,I468568,I31412,I31429,I31446,I31022,I31477,I31010,I31019,I31007,I31563,I192845,I31589,I31597,I31614,I192839,I192830,I31631,I192851,I31657,I192833,I31674,I31682,I192827,I31699,I31531,I31730,I31747,I31543,I31787,I31552,I31809,I192854,I192836,I31826,I192842,I31852,I31869,I31555,I31891,I31540,I31922,I192848,I31939,I31956,I31973,I31549,I32004,I31537,I31546,I31534,I32090,I78650,I32116,I32124,I32141,I78644,I78638,I32158,I78659,I32184,I78656,I32201,I32209,I78653,I32226,I32058,I32257,I32274,I32070,I32314,I32079,I32336,I78641,I32353,I78662,I32379,I32396,I32082,I32418,I32067,I32449,I78647,I32466,I32483,I32500,I32076,I32531,I32064,I32073,I32061,I32617,I335296,I32643,I32651,I32668,I335293,I335308,I32685,I335290,I32711,I335287,I32728,I32736,I32753,I32585,I32784,I32801,I32597,I32841,I32606,I32863,I335302,I32880,I335305,I32906,I32923,I32609,I32945,I32594,I32976,I335299,I32993,I33010,I33027,I32603,I33058,I32591,I32600,I32588,I33144,I281800,I33170,I33178,I33195,I281791,I281809,I33212,I281788,I33238,I33255,I33263,I281794,I33280,I33112,I33311,I33328,I33124,I33368,I33133,I33390,I281806,I281797,I33407,I281812,I33433,I33450,I33136,I33472,I33121,I33503,I281803,I33520,I33537,I33554,I33130,I33585,I33118,I33127,I33115,I33671,I100070,I33697,I33705,I33722,I100064,I100058,I33739,I100079,I33765,I100076,I33782,I33790,I100073,I33807,I33639,I33838,I33855,I33651,I33895,I33660,I33917,I100061,I33934,I100082,I33960,I33977,I33663,I33999,I33648,I34030,I100067,I34047,I34064,I34081,I33657,I34112,I33645,I33654,I33642,I34198,I469134,I34224,I34232,I34249,I469149,I469128,I34266,I469131,I34292,I469152,I34309,I34317,I34334,I34166,I34365,I34382,I34178,I34422,I34187,I34444,I469140,I469137,I34461,I469143,I34487,I34504,I34190,I34526,I34175,I34557,I469146,I34574,I34591,I34608,I34184,I34639,I34172,I34181,I34169,I34725,I402242,I34751,I34759,I34776,I402260,I402254,I34793,I402233,I34819,I402251,I34836,I34844,I402236,I34861,I34693,I34892,I34909,I34705,I402248,I34949,I34714,I34971,I402257,I402245,I34988,I402239,I35014,I35031,I34717,I35053,I34702,I35084,I35101,I35118,I35135,I34711,I35166,I34699,I34708,I34696,I35252,I213706,I35278,I35286,I35303,I213727,I213721,I35320,I213703,I35346,I35363,I35371,I213715,I35388,I35220,I35419,I35436,I35232,I213712,I35476,I35241,I35498,I213718,I213709,I35515,I35541,I35558,I35244,I35580,I35229,I35611,I213724,I35628,I35645,I35662,I35238,I35693,I35226,I35235,I35223,I35779,I503168,I35805,I35813,I35830,I503162,I503183,I35847,I503174,I35873,I503165,I35890,I35898,I503177,I35915,I35747,I35946,I35963,I35759,I36003,I35768,I36025,I503186,I503171,I36042,I36068,I36085,I35771,I36107,I35756,I36138,I503180,I36155,I36172,I36189,I35765,I36220,I35753,I35762,I35750,I36306,I367443,I36332,I36340,I36357,I367440,I367455,I36374,I367437,I36400,I367434,I36417,I36425,I36442,I36274,I36473,I36490,I36286,I36530,I36295,I36552,I367449,I36569,I367452,I36595,I36612,I36298,I36634,I36283,I36665,I367446,I36682,I36699,I36716,I36292,I36747,I36280,I36289,I36277,I36833,I340566,I36859,I36867,I36884,I340563,I340578,I36901,I340560,I36927,I340557,I36944,I36952,I36969,I36801,I37000,I37017,I36813,I37057,I36822,I37079,I340572,I37096,I340575,I37122,I37139,I36825,I37161,I36810,I37192,I340569,I37209,I37226,I37243,I36819,I37274,I36807,I36816,I36804,I37360,I418392,I37386,I37394,I37411,I418410,I418404,I37428,I418383,I37454,I418401,I37471,I37479,I418386,I37496,I37328,I37527,I37544,I37340,I418398,I37584,I37349,I37606,I418407,I418395,I37623,I418389,I37649,I37666,I37352,I37688,I37337,I37719,I37736,I37753,I37770,I37346,I37801,I37334,I37343,I37331,I37887,I243649,I37913,I37921,I37938,I243661,I243646,I37955,I243640,I37981,I243655,I37998,I38006,I243643,I38023,I37855,I38054,I38071,I37867,I243652,I38111,I37876,I38133,I243658,I243664,I38150,I38176,I38193,I37879,I38215,I37864,I38246,I38263,I38280,I38297,I37873,I38328,I37861,I37870,I37858,I38414,I439347,I38440,I38448,I38465,I439344,I439350,I38482,I38508,I38525,I38533,I38550,I38382,I38581,I38598,I38394,I439353,I38638,I38403,I38660,I439356,I439365,I38677,I439359,I38703,I38720,I38406,I38742,I38391,I38773,I439362,I38790,I38807,I38824,I38400,I38855,I38388,I38397,I38385,I38941,I557982,I38967,I38975,I38992,I557976,I557997,I39009,I557973,I39035,I557994,I39052,I39060,I557991,I39077,I38909,I39108,I39125,I38921,I557979,I39165,I38930,I39187,I557988,I557985,I39204,I557970,I39230,I39247,I38933,I39269,I38918,I39300,I39317,I39334,I39351,I38927,I39382,I38915,I38924,I38912,I39468,I403534,I39494,I39502,I39519,I403552,I403546,I39536,I403525,I39562,I403543,I39579,I39587,I403528,I39604,I39436,I39635,I39652,I39448,I403540,I39692,I39457,I39714,I403549,I403537,I39731,I403531,I39757,I39774,I39460,I39796,I39445,I39827,I39844,I39861,I39878,I39454,I39909,I39442,I39451,I39439,I39995,I40021,I40029,I40046,I40063,I40089,I40106,I40114,I40131,I39963,I40162,I40179,I39975,I40219,I39984,I40241,I40258,I40284,I40301,I39987,I40323,I39972,I40354,I40371,I40388,I40405,I39981,I40436,I39969,I39978,I39966,I40522,I271974,I40548,I40556,I40573,I271965,I271983,I40590,I271962,I40616,I40633,I40641,I271968,I40658,I40490,I40689,I40706,I40502,I40746,I40511,I40768,I271980,I271971,I40785,I271986,I40811,I40828,I40514,I40850,I40499,I40881,I271977,I40898,I40915,I40932,I40508,I40963,I40496,I40505,I40493,I41049,I497456,I41075,I41083,I41100,I497471,I497450,I41117,I497453,I41143,I497474,I41160,I41168,I41185,I41017,I41216,I41233,I41029,I41273,I41038,I41295,I497462,I497459,I41312,I497465,I41338,I41355,I41041,I41377,I41026,I41408,I497468,I41425,I41442,I41459,I41035,I41490,I41023,I41032,I41020,I41576,I557387,I41602,I41610,I41627,I557381,I557402,I41644,I557378,I41670,I557399,I41687,I41695,I557396,I41712,I41544,I41743,I41760,I41556,I557384,I41800,I41565,I41822,I557393,I557390,I41839,I557375,I41865,I41882,I41568,I41904,I41553,I41935,I41952,I41969,I41986,I41562,I42017,I41550,I41559,I41547,I42103,I261567,I42129,I42137,I42154,I261579,I261564,I42171,I261558,I42197,I261573,I42214,I42222,I261561,I42239,I42071,I42270,I42287,I42083,I261570,I42327,I42092,I42349,I261576,I261582,I42366,I42392,I42409,I42095,I42431,I42080,I42462,I42479,I42496,I42513,I42089,I42544,I42077,I42086,I42074,I42630,I369551,I42656,I42664,I42681,I369548,I369563,I42698,I369545,I42724,I369542,I42741,I42749,I42766,I42598,I42797,I42814,I42610,I42854,I42619,I42876,I369557,I42893,I369560,I42919,I42936,I42622,I42958,I42607,I42989,I369554,I43006,I43023,I43040,I42616,I43071,I42604,I42613,I42601,I43157,I43183,I43191,I43208,I43225,I43251,I43268,I43276,I43293,I43324,I43341,I43381,I43403,I43420,I43446,I43463,I43485,I43516,I43533,I43550,I43567,I43598,I43684,I151952,I43710,I43718,I43735,I151934,I151949,I43752,I151925,I43778,I151928,I43795,I43803,I151943,I43820,I43652,I43851,I43868,I43664,I151946,I43908,I43673,I43930,I151937,I43947,I151931,I43973,I43990,I43676,I44012,I43661,I44043,I151940,I44060,I44077,I44094,I43670,I44125,I43658,I43667,I43655,I44211,I406118,I44237,I44245,I44262,I406136,I406130,I44279,I406109,I44305,I406127,I44322,I44330,I406112,I44347,I44179,I44378,I44395,I44191,I406124,I44435,I44200,I44457,I406133,I406121,I44474,I406115,I44500,I44517,I44203,I44539,I44188,I44570,I44587,I44604,I44621,I44197,I44652,I44185,I44194,I44182,I44738,I164073,I44764,I44772,I44789,I164055,I164070,I44806,I164046,I44832,I164049,I44849,I44857,I164064,I44874,I44706,I44905,I44922,I44718,I164067,I44962,I44727,I44984,I164058,I45001,I164052,I45027,I45044,I44730,I45066,I44715,I45097,I164061,I45114,I45131,I45148,I44724,I45179,I44712,I44721,I44709,I45265,I441030,I45291,I45299,I45316,I441027,I441033,I45333,I45359,I45376,I45384,I45401,I45233,I45432,I45449,I45245,I441036,I45489,I45254,I45511,I441039,I441048,I45528,I441042,I45554,I45571,I45257,I45593,I45242,I45624,I441045,I45641,I45658,I45675,I45251,I45706,I45239,I45248,I45236,I45792,I481850,I45818,I45826,I45843,I481865,I481844,I45860,I481847,I45886,I481868,I45903,I45911,I45928,I45760,I45959,I45976,I45772,I46016,I45781,I46038,I481856,I481853,I46055,I481859,I46081,I46098,I45784,I46120,I45769,I46151,I481862,I46168,I46185,I46202,I45778,I46233,I45766,I45775,I45763,I46319,I569882,I46345,I46353,I46370,I569876,I569897,I46387,I569873,I46413,I569894,I46430,I46438,I569891,I46455,I46287,I46486,I46503,I46299,I569879,I46543,I46308,I46565,I569888,I569885,I46582,I569870,I46608,I46625,I46311,I46647,I46296,I46678,I46695,I46712,I46729,I46305,I46760,I46293,I46302,I46290,I46846,I566907,I46872,I46880,I46897,I566901,I566922,I46914,I566898,I46940,I566919,I46957,I46965,I566916,I46982,I46814,I47013,I47030,I46826,I566904,I47070,I46835,I47092,I566913,I566910,I47109,I566895,I47135,I47152,I46838,I47174,I46823,I47205,I47222,I47239,I47256,I46832,I47287,I46820,I46829,I46817,I47373,I357957,I47399,I47407,I47424,I357954,I357969,I47441,I357951,I47467,I357948,I47484,I47492,I47509,I47341,I47540,I47557,I47353,I47597,I47362,I47619,I357963,I47636,I357966,I47662,I47679,I47365,I47701,I47350,I47732,I357960,I47749,I47766,I47783,I47359,I47814,I47347,I47356,I47344,I47900,I397074,I47926,I47934,I47951,I397092,I397086,I47968,I397065,I47994,I397083,I48011,I48019,I397068,I48036,I47868,I48067,I48084,I47880,I397080,I48124,I47889,I48146,I397089,I397077,I48163,I397071,I48189,I48206,I47892,I48228,I47877,I48259,I48276,I48293,I48310,I47886,I48341,I47874,I47883,I47871,I48427,I258099,I48453,I48461,I48478,I258111,I258096,I48495,I258090,I48521,I258105,I48538,I48546,I258093,I48563,I48395,I48594,I48611,I48407,I258102,I48651,I48416,I48673,I258108,I258114,I48690,I48716,I48733,I48419,I48755,I48404,I48786,I48803,I48820,I48837,I48413,I48868,I48401,I48410,I48398,I48954,I488208,I48980,I48988,I49005,I488223,I488202,I49022,I488205,I49048,I488226,I49065,I49073,I49090,I48922,I49121,I49138,I48934,I49178,I48943,I49200,I488214,I488211,I49217,I488217,I49243,I49260,I48946,I49282,I48931,I49313,I488220,I49330,I49347,I49364,I48940,I49395,I48928,I48937,I48925,I49481,I106020,I49507,I49515,I49532,I106014,I106008,I49549,I106029,I49575,I106026,I49592,I49600,I106023,I49617,I49449,I49648,I49665,I49461,I49705,I49470,I49727,I106011,I49744,I106032,I49770,I49787,I49473,I49809,I49458,I49840,I106017,I49857,I49874,I49891,I49467,I49922,I49455,I49464,I49452,I50008,I199917,I50034,I50042,I50059,I199911,I199902,I50076,I199923,I50102,I199905,I50119,I50127,I199899,I50144,I49976,I50175,I50192,I49988,I50232,I49997,I50254,I199926,I199908,I50271,I199914,I50297,I50314,I50000,I50336,I49985,I50367,I199920,I50384,I50401,I50418,I49994,I50449,I49982,I49991,I49979,I50535,I565122,I50561,I50569,I50586,I565116,I565137,I50603,I565113,I50629,I565134,I50646,I50654,I565131,I50671,I50503,I50702,I50719,I50515,I565119,I50759,I50524,I50781,I565128,I565125,I50798,I565110,I50824,I50841,I50527,I50863,I50512,I50894,I50911,I50928,I50945,I50521,I50976,I50509,I50518,I50506,I51062,I399012,I51088,I51096,I51113,I399030,I399024,I51130,I399003,I51156,I399021,I51173,I51181,I399006,I51198,I51030,I51229,I51246,I51042,I399018,I51286,I51051,I51308,I399027,I399015,I51325,I399009,I51351,I51368,I51054,I51390,I51039,I51421,I51438,I51455,I51472,I51048,I51503,I51036,I51045,I51033,I51589,I489364,I51615,I51623,I51640,I489379,I489358,I51657,I489361,I51683,I489382,I51700,I51708,I51725,I51557,I51756,I51773,I51569,I51813,I51578,I51835,I489370,I489367,I51852,I489373,I51878,I51895,I51581,I51917,I51566,I51948,I489376,I51965,I51982,I51999,I51575,I52030,I51563,I51572,I51560,I52116,I287580,I52142,I52150,I52167,I287571,I287589,I52184,I287568,I52210,I52227,I52235,I287574,I52252,I52084,I52283,I52300,I52096,I52340,I52105,I52362,I287586,I287577,I52379,I287592,I52405,I52422,I52108,I52444,I52093,I52475,I287583,I52492,I52509,I52526,I52102,I52557,I52090,I52099,I52087,I52643,I297984,I52669,I52677,I52694,I297975,I297993,I52711,I297972,I52737,I52754,I52762,I297978,I52779,I52611,I52810,I52827,I52623,I52867,I52632,I52889,I297990,I297981,I52906,I297996,I52932,I52949,I52635,I52971,I52620,I53002,I297987,I53019,I53036,I53053,I52629,I53084,I52617,I52626,I52614,I53170,I506976,I53196,I53204,I53221,I506970,I506991,I53238,I506982,I53264,I506973,I53281,I53289,I506985,I53306,I53337,I53354,I53394,I53416,I506994,I506979,I53433,I53459,I53476,I53498,I53529,I506988,I53546,I53563,I53580,I53611,I53697,I323994,I53723,I53731,I53748,I323985,I324003,I53765,I323982,I53791,I53808,I53816,I323988,I53833,I53665,I53864,I53881,I53677,I53921,I53686,I53943,I324000,I323991,I53960,I324006,I53986,I54003,I53689,I54025,I53674,I54056,I323997,I54073,I54090,I54107,I53683,I54138,I53671,I53680,I53668,I54224,I54250,I54258,I54275,I54292,I54318,I54335,I54343,I54360,I54192,I54391,I54408,I54204,I54448,I54213,I54470,I54487,I54513,I54530,I54216,I54552,I54201,I54583,I54600,I54617,I54634,I54210,I54665,I54198,I54207,I54195,I54751,I162492,I54777,I54785,I54802,I162474,I162489,I54819,I162465,I54845,I162468,I54862,I54870,I162483,I54887,I54719,I54918,I54935,I54731,I162486,I54975,I54740,I54997,I162477,I55014,I162471,I55040,I55057,I54743,I55079,I54728,I55110,I162480,I55127,I55144,I55161,I54737,I55192,I54725,I54734,I54722,I55278,I454106,I55304,I55312,I55329,I454121,I454100,I55346,I454103,I55372,I454124,I55389,I55397,I55414,I55246,I55445,I55462,I55258,I55502,I55267,I55524,I454112,I454109,I55541,I454115,I55567,I55584,I55270,I55606,I55255,I55637,I454118,I55654,I55671,I55688,I55264,I55719,I55252,I55261,I55249,I55805,I374294,I55831,I55839,I55856,I374291,I374306,I55873,I374288,I55899,I374285,I55916,I55924,I55941,I55773,I55972,I55989,I55785,I56029,I55794,I56051,I374300,I56068,I374303,I56094,I56111,I55797,I56133,I55782,I56164,I374297,I56181,I56198,I56215,I55791,I56246,I55779,I55788,I55776,I56332,I561552,I56358,I56366,I56383,I561546,I561567,I56400,I561543,I56426,I561564,I56443,I56451,I561561,I56468,I56300,I56499,I56516,I56312,I561549,I56556,I56321,I56578,I561558,I561555,I56595,I561540,I56621,I56638,I56324,I56660,I56309,I56691,I56708,I56725,I56742,I56318,I56773,I56306,I56315,I56303,I56859,I56885,I56893,I56910,I56927,I56953,I56970,I56978,I56995,I56827,I57026,I57043,I56839,I57083,I56848,I57105,I57122,I57148,I57165,I56851,I57187,I56836,I57218,I57235,I57252,I57269,I56845,I57300,I56833,I56842,I56830,I57386,I365335,I57412,I57420,I57437,I365332,I365347,I57454,I365329,I57480,I365326,I57497,I57505,I57522,I57354,I57553,I57570,I57366,I57610,I57375,I57632,I365341,I57649,I365344,I57675,I57692,I57378,I57714,I57363,I57745,I365338,I57762,I57779,I57796,I57372,I57827,I57360,I57369,I57357,I57913,I236713,I57939,I57947,I57964,I236725,I236710,I57981,I236704,I58007,I236719,I58024,I58032,I236707,I58049,I57881,I58080,I58097,I57893,I236716,I58137,I57902,I58159,I236722,I236728,I58176,I58202,I58219,I57905,I58241,I57890,I58272,I58289,I58306,I58323,I57899,I58354,I57887,I57896,I57884,I58443,I144556,I58469,I58477,I144553,I58503,I58511,I144550,I58528,I144562,I58545,I58420,I58576,I144571,I58414,I58607,I144568,I58624,I58641,I144547,I58658,I58675,I58692,I58429,I58426,I58432,I58751,I58768,I58785,I144559,I144574,I58811,I58411,I58842,I58850,I144565,I58435,I58881,I58898,I58915,I58417,I58946,I58963,I58408,I58423,I59038,I371129,I59064,I59072,I59098,I59106,I371126,I59123,I371138,I59140,I59015,I59171,I371132,I59009,I59202,I371144,I59219,I59236,I371135,I371123,I59253,I59270,I59287,I59024,I59021,I59027,I59346,I59363,I59380,I59406,I59006,I59437,I59445,I371141,I59030,I59476,I59493,I59510,I59012,I59541,I59558,I59003,I59018,I59633,I251169,I59659,I59667,I251154,I59693,I59701,I251178,I59718,I251157,I59735,I59610,I59766,I251160,I59604,I59797,I251163,I59814,I59831,I251166,I251172,I59848,I59865,I59882,I59619,I59616,I59622,I59941,I59958,I59975,I251175,I60001,I59601,I60032,I60040,I59625,I60071,I60088,I60105,I59607,I60136,I60153,I59598,I59613,I60228,I284100,I60254,I60262,I284121,I60288,I60296,I60313,I284112,I60330,I60205,I60361,I284109,I60199,I60392,I284118,I60409,I60426,I284103,I60443,I60460,I60477,I60214,I60211,I60217,I60536,I60553,I60570,I284124,I284106,I60596,I60196,I60627,I60635,I284115,I60220,I60666,I60683,I60700,I60202,I60731,I60748,I60193,I60208,I60823,I521117,I60849,I60857,I521114,I60883,I60891,I521132,I60908,I521126,I60925,I60800,I60956,I521120,I60794,I60987,I61004,I61021,I521123,I521129,I61038,I61055,I61072,I60809,I60806,I60812,I61131,I61148,I61165,I521135,I61191,I60791,I61222,I61230,I521138,I60815,I61261,I61278,I61295,I60797,I61326,I61343,I60788,I60803,I61418,I149299,I61444,I61452,I149296,I61478,I61486,I149293,I61503,I149305,I61520,I61395,I61551,I149314,I61389,I61582,I149311,I61599,I61616,I149290,I61633,I61650,I61667,I61404,I61401,I61407,I61726,I61743,I61760,I149302,I149317,I61786,I61386,I61817,I61825,I149308,I61410,I61856,I61873,I61890,I61392,I61921,I61938,I61383,I61398,I62013,I62039,I62047,I62073,I62081,I62098,I62115,I61990,I62146,I61984,I62177,I62194,I62211,I62228,I62245,I62262,I61999,I61996,I62002,I62321,I62338,I62355,I62381,I61981,I62412,I62420,I62005,I62451,I62468,I62485,I61987,I62516,I62533,I61978,I61993,I62605,I148763,I62631,I62648,I62670,I148778,I62696,I62704,I62721,I148775,I62738,I62755,I62772,I148772,I62789,I148787,I62806,I148784,I62823,I62854,I62871,I62888,I62905,I62950,I148781,I62995,I63012,I148769,I63029,I148790,I63046,I148766,I63072,I63080,I63134,I63142,I63200,I63226,I63243,I63192,I63265,I63291,I63299,I63316,I63333,I63350,I63367,I63384,I63401,I63418,I63168,I63449,I63466,I63483,I63500,I63180,I63174,I63545,I63189,I63183,I63590,I63607,I63624,I63641,I63667,I63675,I63177,I63171,I63729,I63737,I63186,I63795,I156141,I63821,I63838,I63787,I63860,I156156,I63886,I63894,I63911,I156153,I63928,I63945,I63962,I156150,I63979,I156165,I63996,I156162,I64013,I63763,I64044,I64061,I64078,I64095,I63775,I63769,I64140,I156159,I63784,I63778,I64185,I64202,I156147,I64219,I156168,I64236,I156144,I64262,I64270,I63772,I63766,I64324,I64332,I63781,I64390,I495138,I64416,I64433,I64382,I64455,I64481,I64489,I64506,I495141,I64523,I495153,I64540,I64557,I495159,I64574,I495150,I64591,I495156,I64608,I64358,I64639,I64656,I64673,I64690,I64370,I64364,I64735,I495147,I64379,I64373,I64780,I64797,I495144,I64814,I495162,I64831,I64857,I64865,I64367,I64361,I64919,I64927,I64376,I64985,I549661,I65011,I65028,I64977,I65050,I549652,I65076,I65084,I65101,I549646,I65118,I549640,I65135,I65152,I549667,I65169,I65186,I549664,I65203,I64953,I65234,I65251,I65268,I65285,I64965,I64959,I65330,I549649,I64974,I64968,I65375,I65392,I549655,I65409,I549658,I65426,I549643,I65452,I65460,I64962,I64956,I65514,I65522,I64971,I65580,I191219,I65606,I65623,I65572,I65645,I191207,I65671,I65679,I65696,I191216,I65713,I191213,I65730,I65747,I191204,I65764,I191210,I65781,I191195,I65798,I65548,I65829,I65846,I65863,I65880,I65560,I65554,I65925,I65569,I65563,I65970,I65987,I191201,I66004,I191198,I66021,I191222,I66047,I66055,I65557,I65551,I66109,I66117,I65566,I66175,I112400,I66201,I66218,I66167,I66240,I112415,I66266,I66274,I66291,I112412,I66308,I66325,I66342,I112409,I66359,I112424,I66376,I112421,I66393,I66143,I66424,I66441,I66458,I66475,I66155,I66149,I66520,I112418,I66164,I66158,I66565,I66582,I112406,I66599,I112427,I66616,I112403,I66642,I66650,I66152,I66146,I66704,I66712,I66161,I66770,I245389,I66796,I66813,I66762,I66835,I245380,I66861,I66869,I66886,I245398,I66903,I245395,I66920,I66937,I245374,I66954,I245377,I66971,I245386,I66988,I66738,I67019,I67036,I67053,I67070,I66750,I66744,I67115,I245392,I66759,I66753,I67160,I67177,I67194,I245383,I67211,I67237,I67245,I66747,I66741,I67299,I67307,I66756,I67365,I67391,I67408,I67357,I67430,I67456,I67464,I67481,I67498,I67515,I67532,I67549,I67566,I67583,I67333,I67614,I67631,I67648,I67665,I67345,I67339,I67710,I67354,I67348,I67755,I67772,I67789,I67806,I67832,I67840,I67342,I67336,I67894,I67902,I67351,I67960,I334239,I67986,I68003,I67952,I68025,I334233,I68051,I68059,I68076,I334251,I68093,I68110,I68127,I68144,I334245,I68161,I334236,I68178,I67928,I68209,I68226,I68243,I68260,I67940,I67934,I68305,I334248,I67949,I67943,I68350,I68367,I334254,I68384,I68401,I334242,I68427,I68435,I67937,I67931,I68489,I68497,I67946,I68555,I360062,I68581,I68598,I68547,I68620,I360056,I68646,I68654,I68671,I360074,I68688,I68705,I68722,I68739,I360068,I68756,I360059,I68773,I68523,I68804,I68821,I68838,I68855,I68535,I68529,I68900,I360071,I68544,I68538,I68945,I68962,I360077,I68979,I68996,I360065,I69022,I69030,I68532,I68526,I69084,I69092,I68541,I69150,I295094,I69176,I69193,I69142,I69215,I295091,I69241,I69249,I69266,I295097,I69283,I295082,I69300,I69317,I295085,I69334,I295106,I69351,I295103,I69368,I69118,I69399,I69416,I69433,I69450,I69130,I69124,I69495,I69139,I69133,I69540,I69557,I295088,I69574,I295100,I69591,I69617,I69625,I69127,I69121,I69679,I69687,I69136,I69745,I318214,I69771,I69788,I69737,I69810,I318211,I69836,I69844,I69861,I318217,I69878,I318202,I69895,I69912,I318205,I69929,I318226,I69946,I318223,I69963,I69713,I69994,I70011,I70028,I70045,I69725,I69719,I70090,I69734,I69728,I70135,I70152,I318208,I70169,I318220,I70186,I70212,I70220,I69722,I69716,I70274,I70282,I69731,I70340,I393204,I70366,I70383,I70332,I70405,I393213,I70431,I70439,I70456,I393201,I70473,I393192,I70490,I70507,I393198,I70524,I393216,I70541,I393189,I70558,I70308,I70589,I70606,I70623,I70640,I70320,I70314,I70685,I393195,I70329,I70323,I70730,I70747,I393207,I70764,I70781,I393210,I70807,I70815,I70317,I70311,I70869,I70877,I70326,I70935,I165100,I70961,I70978,I71000,I165115,I71026,I71034,I71051,I165112,I71068,I71085,I71102,I165109,I71119,I165124,I71136,I165121,I71153,I71184,I71201,I71218,I71235,I71280,I165118,I71325,I71342,I165106,I71359,I165127,I71376,I165103,I71402,I71410,I71464,I71472,I71530,I424200,I71556,I71573,I71522,I71595,I424209,I71621,I71629,I71646,I424203,I71663,I424197,I71680,I71697,I424212,I71714,I71731,I424206,I71748,I71498,I71779,I71796,I71813,I71830,I71510,I71504,I71875,I71519,I71513,I71920,I71937,I424218,I71954,I424215,I71971,I71997,I72005,I71507,I71501,I72059,I72067,I71516,I72125,I345833,I72151,I72168,I72117,I72190,I345827,I72216,I72224,I72241,I345845,I72258,I72275,I72292,I72309,I345839,I72326,I345830,I72343,I72093,I72374,I72391,I72408,I72425,I72105,I72099,I72470,I345842,I72114,I72108,I72515,I72532,I345848,I72549,I72566,I345836,I72592,I72600,I72102,I72096,I72654,I72662,I72111,I72720,I359008,I72746,I72763,I72785,I359002,I72811,I72819,I72836,I359020,I72853,I72870,I72887,I72904,I359014,I72921,I359005,I72938,I72969,I72986,I73003,I73020,I73065,I359017,I73110,I73127,I359023,I73144,I73161,I359011,I73187,I73195,I73249,I73257,I73315,I225615,I73341,I73358,I73307,I73380,I225609,I73406,I73414,I73431,I225624,I73448,I225621,I73465,I73482,I225612,I73499,I225603,I73516,I225606,I73533,I73283,I73564,I73581,I73598,I73615,I73295,I73289,I73660,I225627,I73304,I73298,I73705,I73722,I225618,I73739,I73756,I73782,I73790,I73292,I73286,I73844,I73852,I73301,I73910,I73936,I73953,I73902,I73975,I74001,I74009,I74026,I74043,I74060,I74077,I74094,I74111,I74128,I73878,I74159,I74176,I74193,I74210,I73890,I73884,I74255,I73899,I73893,I74300,I74317,I74334,I74351,I74377,I74385,I73887,I73881,I74439,I74447,I73896,I74505,I240187,I74531,I74548,I74497,I74570,I240178,I74596,I74604,I74621,I240196,I74638,I240193,I74655,I74672,I240172,I74689,I240175,I74706,I240184,I74723,I74473,I74754,I74771,I74788,I74805,I74485,I74479,I74850,I240190,I74494,I74488,I74895,I74912,I74929,I240181,I74946,I74972,I74980,I74482,I74476,I75034,I75042,I74491,I75100,I430371,I75126,I75143,I75092,I75165,I430380,I75191,I75199,I75216,I430374,I75233,I430368,I75250,I75267,I430383,I75284,I75301,I430377,I75318,I75068,I75349,I75366,I75383,I75400,I75080,I75074,I75445,I75089,I75083,I75490,I75507,I430389,I75524,I430386,I75541,I75567,I75575,I75077,I75071,I75629,I75637,I75086,I75695,I145601,I75721,I75738,I75687,I75760,I145616,I75786,I75794,I75811,I145613,I75828,I75845,I75862,I145610,I75879,I145625,I75896,I145622,I75913,I75663,I75944,I75961,I75978,I75995,I75675,I75669,I76040,I145619,I75684,I75678,I76085,I76102,I145607,I76119,I145628,I76136,I145604,I76162,I76170,I75672,I75666,I76224,I76232,I75681,I76290,I190131,I76316,I76333,I76282,I76355,I190119,I76381,I76389,I76406,I190128,I76423,I190125,I76440,I76457,I190116,I76474,I190122,I76491,I190107,I76508,I76258,I76539,I76556,I76573,I76590,I76270,I76264,I76635,I76279,I76273,I76680,I76697,I190113,I76714,I190110,I76731,I190134,I76757,I76765,I76267,I76261,I76819,I76827,I76276,I76885,I76911,I76928,I76877,I76950,I76976,I76984,I77001,I77018,I77035,I77052,I77069,I77086,I77103,I76853,I77134,I77151,I77168,I77185,I76865,I76859,I77230,I76874,I76868,I77275,I77292,I77309,I77326,I77352,I77360,I76862,I76856,I77414,I77422,I76871,I77480,I302608,I77506,I77523,I77545,I302605,I77571,I77579,I77596,I302611,I77613,I302596,I77630,I77647,I302599,I77664,I302620,I77681,I302617,I77698,I77729,I77746,I77763,I77780,I77825,I77870,I77887,I302602,I77904,I302614,I77921,I77947,I77955,I78009,I78017,I78075,I146128,I78101,I78118,I78067,I78140,I146143,I78166,I78174,I78191,I146140,I78208,I78225,I78242,I146137,I78259,I146152,I78276,I146149,I78293,I78043,I78324,I78341,I78358,I78375,I78055,I78049,I78420,I146146,I78064,I78058,I78465,I78482,I146134,I78499,I146155,I78516,I146131,I78542,I78550,I78052,I78046,I78604,I78612,I78061,I78670,I505900,I78696,I78713,I78735,I505885,I78761,I78769,I78786,I505903,I78803,I78820,I78837,I505906,I78854,I505897,I78871,I505894,I78888,I78919,I78936,I78953,I78970,I79015,I505891,I79060,I79077,I505882,I79094,I505888,I79111,I79137,I79145,I79199,I79207,I79265,I500340,I79291,I79308,I79257,I79330,I79356,I79364,I79381,I500343,I79398,I500355,I79415,I79432,I500361,I79449,I500352,I79466,I500358,I79483,I79233,I79514,I79531,I79548,I79565,I79245,I79239,I79610,I500349,I79254,I79248,I79655,I79672,I500346,I79689,I500364,I79706,I79732,I79740,I79242,I79236,I79794,I79802,I79251,I79860,I562751,I79886,I79903,I79852,I79925,I562742,I79951,I79959,I79976,I562736,I79993,I562730,I80010,I80027,I562757,I80044,I80061,I562754,I80078,I79828,I80109,I80126,I80143,I80160,I79840,I79834,I80205,I562739,I79849,I79843,I80250,I80267,I562745,I80284,I562748,I80301,I562733,I80327,I80335,I79837,I79831,I80389,I80397,I79846,I80455,I434859,I80481,I80498,I80447,I80520,I434868,I80546,I80554,I80571,I434862,I80588,I434856,I80605,I80622,I434871,I80639,I80656,I434865,I80673,I80423,I80704,I80721,I80738,I80755,I80435,I80429,I80800,I80444,I80438,I80845,I80862,I434877,I80879,I434874,I80896,I80922,I80930,I80432,I80426,I80984,I80992,I80441,I81050,I157195,I81076,I81093,I81042,I81115,I157210,I81141,I81149,I81166,I157207,I81183,I81200,I81217,I157204,I81234,I157219,I81251,I157216,I81268,I81018,I81299,I81316,I81333,I81350,I81030,I81024,I81395,I157213,I81039,I81033,I81440,I81457,I157201,I81474,I157222,I81491,I157198,I81517,I81525,I81027,I81021,I81579,I81587,I81036,I81645,I352157,I81671,I81688,I81637,I81710,I352151,I81736,I81744,I81761,I352169,I81778,I81795,I81812,I81829,I352163,I81846,I352154,I81863,I81613,I81894,I81911,I81928,I81945,I81625,I81619,I81990,I352166,I81634,I81628,I82035,I82052,I352172,I82069,I82086,I352160,I82112,I82120,I81622,I81616,I82174,I82182,I81631,I82240,I161411,I82266,I82283,I82305,I161426,I82331,I82339,I82356,I161423,I82373,I82390,I82407,I161420,I82424,I161435,I82441,I161432,I82458,I82489,I82506,I82523,I82540,I82585,I161429,I82630,I82647,I161417,I82664,I161438,I82681,I161414,I82707,I82715,I82769,I82777,I82835,I440469,I82861,I82878,I82827,I82900,I440478,I82926,I82934,I82951,I440472,I82968,I440466,I82985,I83002,I440481,I83019,I83036,I440475,I83053,I82803,I83084,I83101,I83118,I83135,I82815,I82809,I83180,I82824,I82818,I83225,I83242,I440487,I83259,I440484,I83276,I83302,I83310,I82812,I82806,I83364,I83372,I82821,I83430,I299140,I83456,I83473,I83495,I299137,I83521,I83529,I83546,I299143,I83563,I299128,I83580,I83597,I299131,I83614,I299152,I83631,I299149,I83648,I83679,I83696,I83713,I83730,I83775,I83820,I83837,I299134,I83854,I299146,I83871,I83897,I83905,I83959,I83967,I84025,I214905,I84051,I84068,I84017,I84090,I214899,I84116,I84124,I84141,I214914,I84158,I214911,I84175,I84192,I214902,I84209,I214893,I84226,I214896,I84243,I83993,I84274,I84291,I84308,I84325,I84005,I83999,I84370,I214917,I84014,I84008,I84415,I84432,I214908,I84449,I84466,I84492,I84500,I84002,I83996,I84554,I84562,I84011,I84620,I118197,I84646,I84663,I84685,I118212,I84711,I84719,I84736,I118209,I84753,I84770,I84787,I118206,I84804,I118221,I84821,I118218,I84838,I84869,I84886,I84903,I84920,I84965,I118215,I85010,I85027,I118203,I85044,I118224,I85061,I118200,I85087,I85095,I85149,I85157,I85215,I512428,I85241,I85258,I85207,I85280,I512413,I85306,I85314,I85331,I512431,I85348,I85365,I85382,I512434,I85399,I512425,I85416,I512422,I85433,I85183,I85464,I85481,I85498,I85515,I85195,I85189,I85560,I512419,I85204,I85198,I85605,I85622,I512410,I85639,I512416,I85656,I85682,I85690,I85192,I85186,I85744,I85752,I85201,I85810,I191763,I85836,I85853,I85802,I85875,I191751,I85901,I85909,I85926,I191760,I85943,I191757,I85960,I85977,I191748,I85994,I191754,I86011,I191739,I86028,I85778,I86059,I86076,I86093,I86110,I85790,I85784,I86155,I85799,I85793,I86200,I86217,I191745,I86234,I191742,I86251,I191766,I86277,I86285,I85787,I85781,I86339,I86347,I85796,I86405,I392558,I86431,I86448,I86397,I86470,I392567,I86496,I86504,I86521,I392555,I86538,I392546,I86555,I86572,I392552,I86589,I392570,I86606,I392543,I86623,I86373,I86654,I86671,I86688,I86705,I86385,I86379,I86750,I392549,I86394,I86388,I86795,I86812,I392561,I86829,I86846,I392564,I86872,I86880,I86382,I86376,I86934,I86942,I86391,I87000,I429249,I87026,I87043,I86992,I87065,I429258,I87091,I87099,I87116,I429252,I87133,I429246,I87150,I87167,I429261,I87184,I87201,I429255,I87218,I86968,I87249,I87266,I87283,I87300,I86980,I86974,I87345,I86989,I86983,I87390,I87407,I429267,I87424,I429264,I87441,I87467,I87475,I86977,I86971,I87529,I87537,I86986,I87595,I109765,I87621,I87638,I87587,I87660,I109780,I87686,I87694,I87711,I109777,I87728,I87745,I87762,I109774,I87779,I109789,I87796,I109786,I87813,I87563,I87844,I87861,I87878,I87895,I87575,I87569,I87940,I109783,I87584,I87578,I87985,I88002,I109771,I88019,I109792,I88036,I109768,I88062,I88070,I87572,I87566,I88124,I88132,I87581,I88190,I364805,I88216,I88233,I88182,I88255,I364799,I88281,I88289,I88306,I364817,I88323,I88340,I88357,I88374,I364811,I88391,I364802,I88408,I88158,I88439,I88456,I88473,I88490,I88170,I88164,I88535,I364814,I88179,I88173,I88580,I88597,I364820,I88614,I88631,I364808,I88657,I88665,I88167,I88161,I88719,I88727,I88176,I88785,I88811,I88828,I88777,I88850,I88876,I88884,I88901,I88918,I88935,I88952,I88969,I88986,I89003,I88753,I89034,I89051,I89068,I89085,I88765,I88759,I89130,I88774,I88768,I89175,I89192,I89209,I89226,I89252,I89260,I88762,I88756,I89314,I89322,I88771,I89380,I454678,I89406,I89423,I89372,I89445,I89471,I89479,I89496,I454681,I89513,I454693,I89530,I89547,I454699,I89564,I454690,I89581,I454696,I89598,I89348,I89629,I89646,I89663,I89680,I89360,I89354,I89725,I454687,I89369,I89363,I89770,I89787,I454684,I89804,I454702,I89821,I89847,I89855,I89357,I89351,I89909,I89917,I89366,I89975,I504812,I90001,I90018,I89967,I90040,I504797,I90066,I90074,I90091,I504815,I90108,I90125,I90142,I504818,I90159,I504809,I90176,I504806,I90193,I89943,I90224,I90241,I90258,I90275,I89955,I89949,I90320,I504803,I89964,I89958,I90365,I90382,I504794,I90399,I504800,I90416,I90442,I90450,I89952,I89946,I90504,I90512,I89961,I90570,I184691,I90596,I90613,I90562,I90635,I184679,I90661,I90669,I90686,I184688,I90703,I184685,I90720,I90737,I184676,I90754,I184682,I90771,I184667,I90788,I90538,I90819,I90836,I90853,I90870,I90550,I90544,I90915,I90559,I90553,I90960,I90977,I184673,I90994,I184670,I91011,I184694,I91037,I91045,I90547,I90541,I91099,I91107,I90556,I91165,I323416,I91191,I91208,I91157,I91230,I323413,I91256,I91264,I91281,I323419,I91298,I323404,I91315,I91332,I323407,I91349,I323428,I91366,I323425,I91383,I91133,I91414,I91431,I91448,I91465,I91145,I91139,I91510,I91154,I91148,I91555,I91572,I323410,I91589,I323422,I91606,I91632,I91640,I91142,I91136,I91694,I91702,I91151,I91760,I91786,I91803,I91825,I91851,I91859,I91876,I91893,I91910,I91927,I91944,I91961,I91978,I92009,I92026,I92043,I92060,I92105,I92150,I92167,I92184,I92201,I92227,I92235,I92289,I92297,I92355,I488780,I92381,I92398,I92347,I92420,I92446,I92454,I92471,I488783,I92488,I488795,I92505,I92522,I488801,I92539,I488792,I92556,I488798,I92573,I92323,I92604,I92621,I92638,I92655,I92335,I92329,I92700,I488789,I92344,I92338,I92745,I92762,I488786,I92779,I488804,I92796,I92822,I92830,I92332,I92326,I92884,I92892,I92341,I92950,I250591,I92976,I92993,I92942,I93015,I250582,I93041,I93049,I93066,I250600,I93083,I250597,I93100,I93117,I250576,I93134,I250579,I93151,I250588,I93168,I92918,I93199,I93216,I93233,I93250,I92930,I92924,I93295,I250594,I92939,I92933,I93340,I93357,I93374,I250585,I93391,I93417,I93425,I92927,I92921,I93479,I93487,I92936,I93545,I277754,I93571,I93588,I93537,I93610,I277751,I93636,I93644,I93661,I277757,I93678,I277742,I93695,I93712,I277745,I93729,I277766,I93746,I277763,I93763,I93513,I93794,I93811,I93828,I93845,I93525,I93519,I93890,I93534,I93528,I93935,I93952,I277748,I93969,I277760,I93986,I94012,I94020,I93522,I93516,I94074,I94082,I93531,I94140,I135061,I94166,I94183,I94132,I94205,I135076,I94231,I94239,I94256,I135073,I94273,I94290,I94307,I135070,I94324,I135085,I94341,I135082,I94358,I94108,I94389,I94406,I94423,I94440,I94120,I94114,I94485,I135079,I94129,I94123,I94530,I94547,I135067,I94564,I135088,I94581,I135064,I94607,I94615,I94117,I94111,I94669,I94677,I94126,I94735,I244811,I94761,I94778,I94727,I94800,I244802,I94826,I94834,I94851,I244820,I94868,I244817,I94885,I94902,I244796,I94919,I244799,I94936,I244808,I94953,I94703,I94984,I95001,I95018,I95035,I94715,I94709,I95080,I244814,I94724,I94718,I95125,I95142,I95159,I244805,I95176,I95202,I95210,I94712,I94706,I95264,I95272,I94721,I95330,I117670,I95356,I95373,I95322,I95395,I117685,I95421,I95429,I95446,I117682,I95463,I95480,I95497,I117679,I95514,I117694,I95531,I117691,I95548,I95298,I95579,I95596,I95613,I95630,I95310,I95304,I95675,I117688,I95319,I95313,I95720,I95737,I117676,I95754,I117697,I95771,I117673,I95797,I95805,I95307,I95301,I95859,I95867,I95316,I95925,I122940,I95951,I95968,I95917,I95990,I122955,I96016,I96024,I96041,I122952,I96058,I96075,I96092,I122949,I96109,I122964,I96126,I122961,I96143,I95893,I96174,I96191,I96208,I96225,I95905,I95899,I96270,I122958,I95914,I95908,I96315,I96332,I122946,I96349,I122967,I96366,I122943,I96392,I96400,I95902,I95896,I96454,I96462,I95911,I96520,I475486,I96546,I96563,I96512,I96585,I96611,I96619,I96636,I475489,I96653,I475501,I96670,I96687,I475507,I96704,I475498,I96721,I475504,I96738,I96488,I96769,I96786,I96803,I96820,I96500,I96494,I96865,I475495,I96509,I96503,I96910,I96927,I475492,I96944,I475510,I96961,I96987,I96995,I96497,I96491,I97049,I97057,I96506,I97115,I180883,I97141,I97158,I97107,I97180,I180871,I97206,I97214,I97231,I180880,I97248,I180877,I97265,I97282,I180868,I97299,I180874,I97316,I180859,I97333,I97083,I97364,I97381,I97398,I97415,I97095,I97089,I97460,I97104,I97098,I97505,I97522,I180865,I97539,I180862,I97556,I180886,I97582,I97590,I97092,I97086,I97644,I97652,I97101,I97710,I302030,I97736,I97753,I97775,I302027,I97801,I97809,I97826,I302033,I97843,I302018,I97860,I97877,I302021,I97894,I302042,I97911,I302039,I97928,I97959,I97976,I97993,I98010,I98055,I98100,I98117,I302024,I98134,I302036,I98151,I98177,I98185,I98239,I98247,I98305,I361643,I98331,I98348,I98297,I98370,I361637,I98396,I98404,I98421,I361655,I98438,I98455,I98472,I98489,I361649,I98506,I361640,I98523,I98273,I98554,I98571,I98588,I98605,I98285,I98279,I98650,I361652,I98294,I98288,I98695,I98712,I361658,I98729,I98746,I361646,I98772,I98780,I98282,I98276,I98834,I98842,I98291,I98900,I462192,I98926,I98943,I98892,I98965,I98991,I98999,I99016,I462195,I99033,I462207,I99050,I99067,I462213,I99084,I462204,I99101,I462210,I99118,I98868,I99149,I99166,I99183,I99200,I98880,I98874,I99245,I462201,I98889,I98883,I99290,I99307,I462198,I99324,I462216,I99341,I99367,I99375,I98877,I98871,I99429,I99437,I98886,I99495,I370075,I99521,I99538,I99487,I99560,I370069,I99586,I99594,I99611,I370087,I99628,I99645,I99662,I99679,I370081,I99696,I370072,I99713,I99463,I99744,I99761,I99778,I99795,I99475,I99469,I99840,I370084,I99484,I99478,I99885,I99902,I370090,I99919,I99936,I370078,I99962,I99970,I99472,I99466,I100024,I100032,I99481,I100090,I230939,I100116,I100133,I100155,I230930,I100181,I100189,I100206,I230948,I100223,I230945,I100240,I100257,I230924,I100274,I230927,I100291,I230936,I100308,I100339,I100356,I100373,I100390,I100435,I230942,I100480,I100497,I100514,I230933,I100531,I100557,I100565,I100619,I100627,I100685,I516780,I100711,I100728,I100677,I100750,I516765,I100776,I100784,I100801,I516783,I100818,I100835,I100852,I516786,I100869,I516777,I100886,I516774,I100903,I100653,I100934,I100951,I100968,I100985,I100665,I100659,I101030,I516771,I100674,I100668,I101075,I101092,I516762,I101109,I516768,I101126,I101152,I101160,I100662,I100656,I101214,I101222,I100671,I101280,I415814,I101306,I101323,I101272,I101345,I415823,I101371,I101379,I101396,I415811,I101413,I415802,I101430,I101447,I415808,I101464,I415826,I101481,I415799,I101498,I101248,I101529,I101546,I101563,I101580,I101260,I101254,I101625,I415805,I101269,I101263,I101670,I101687,I415817,I101704,I101721,I415820,I101747,I101755,I101257,I101251,I101809,I101817,I101266,I101875,I158776,I101901,I101918,I101867,I101940,I158791,I101966,I101974,I101991,I158788,I102008,I102025,I102042,I158785,I102059,I158800,I102076,I158797,I102093,I101843,I102124,I102141,I102158,I102175,I101855,I101849,I102220,I158794,I101864,I101858,I102265,I102282,I158782,I102299,I158803,I102316,I158779,I102342,I102350,I101852,I101846,I102404,I102412,I101861,I102470,I265616,I102496,I102513,I102535,I265613,I102561,I102569,I102586,I265619,I102603,I265604,I102620,I102637,I265607,I102654,I265628,I102671,I265625,I102688,I102719,I102736,I102753,I102770,I102815,I102860,I102877,I265610,I102894,I265622,I102911,I102937,I102945,I102999,I103007,I103065,I434298,I103091,I103108,I103057,I103130,I434307,I103156,I103164,I103181,I434301,I103198,I434295,I103215,I103232,I434310,I103249,I103266,I434304,I103283,I103033,I103314,I103331,I103348,I103365,I103045,I103039,I103410,I103054,I103048,I103455,I103472,I434316,I103489,I434313,I103506,I103532,I103540,I103042,I103036,I103594,I103602,I103051,I103660,I528631,I103686,I103703,I103652,I103725,I528643,I103751,I103759,I103776,I528637,I103793,I528649,I103810,I103827,I528634,I103844,I528646,I103861,I528628,I103878,I103628,I103909,I103926,I103943,I103960,I103640,I103634,I104005,I528640,I103649,I103643,I104050,I104067,I104084,I104101,I528652,I104127,I104135,I103637,I103631,I104189,I104197,I103646,I104255,I134007,I104281,I104298,I104247,I104320,I134022,I104346,I104354,I104371,I134019,I104388,I104405,I104422,I134016,I104439,I134031,I104456,I134028,I104473,I104223,I104504,I104521,I104538,I104555,I104235,I104229,I104600,I134025,I104244,I104238,I104645,I104662,I134013,I104679,I134034,I104696,I134010,I104722,I104730,I104232,I104226,I104784,I104792,I104241,I104850,I219070,I104876,I104893,I104842,I104915,I219064,I104941,I104949,I104966,I219079,I104983,I219076,I105000,I105017,I219067,I105034,I219058,I105051,I219061,I105068,I104818,I105099,I105116,I105133,I105150,I104830,I104824,I105195,I219082,I104839,I104833,I105240,I105257,I219073,I105274,I105291,I105317,I105325,I104827,I104821,I105379,I105387,I104836,I105445,I339509,I105471,I105488,I105437,I105510,I339503,I105536,I105544,I105561,I339521,I105578,I105595,I105612,I105629,I339515,I105646,I339506,I105663,I105413,I105694,I105711,I105728,I105745,I105425,I105419,I105790,I339518,I105434,I105428,I105835,I105852,I339524,I105869,I105886,I339512,I105912,I105920,I105422,I105416,I105974,I105982,I105431,I106040,I150344,I106066,I106083,I106105,I150359,I106131,I106139,I106156,I150356,I106173,I106190,I106207,I150353,I106224,I150368,I106241,I150365,I106258,I106289,I106306,I106323,I106340,I106385,I150362,I106430,I106447,I150350,I106464,I150371,I106481,I150347,I106507,I106515,I106569,I106577,I106638,I106664,I106672,I106689,I106715,I106606,I106737,I106763,I106771,I106788,I106814,I106630,I106836,I106612,I106876,I106893,I106901,I106918,I106615,I106949,I106966,I106992,I107000,I106603,I106621,I107045,I107062,I106624,I106609,I106618,I106627,I107165,I107191,I107199,I107216,I107242,I107133,I107264,I107290,I107298,I107315,I107341,I107157,I107363,I107139,I107403,I107420,I107428,I107445,I107142,I107476,I107493,I107519,I107527,I107130,I107148,I107572,I107589,I107151,I107136,I107145,I107154,I107692,I107718,I107726,I107743,I107769,I107660,I107791,I107817,I107825,I107842,I107868,I107684,I107890,I107666,I107930,I107947,I107955,I107972,I107669,I108003,I108020,I108046,I108054,I107657,I107675,I108099,I108116,I107678,I107663,I107672,I107681,I108219,I341087,I108245,I108253,I341090,I341084,I108270,I341096,I108296,I108187,I108318,I341099,I108344,I108352,I108369,I108395,I108211,I108417,I108193,I341102,I108457,I108474,I108482,I108499,I108196,I108530,I341093,I108547,I108573,I108581,I108184,I108202,I108626,I341105,I108643,I108205,I108190,I108199,I108208,I108746,I283534,I108772,I108780,I283525,I283540,I108797,I283546,I108823,I108714,I108845,I283531,I108871,I108879,I108896,I108922,I108738,I108944,I108720,I283528,I108984,I109001,I109009,I109026,I108723,I109057,I283522,I283537,I109074,I109100,I109108,I108711,I108729,I109153,I283543,I109170,I108732,I108717,I108726,I108735,I109273,I249435,I109299,I109307,I249420,I249423,I109324,I249438,I109350,I109241,I109372,I249432,I109398,I109406,I109423,I109449,I109265,I109471,I109247,I249429,I109511,I109528,I109536,I109553,I109250,I109584,I249444,I109601,I249441,I109627,I109635,I109238,I109256,I109680,I249426,I109697,I109259,I109244,I109253,I109262,I109800,I109826,I109834,I109851,I109877,I109899,I109925,I109933,I109950,I109976,I109998,I110038,I110055,I110063,I110080,I110111,I110128,I110154,I110162,I110207,I110224,I110327,I205895,I110353,I110361,I205907,I205886,I110378,I205910,I110404,I110295,I110426,I205901,I110452,I110460,I205883,I110477,I110503,I110319,I110525,I110301,I205898,I110565,I110582,I110590,I110607,I110304,I110638,I205889,I110655,I205892,I110681,I110689,I110292,I110310,I110734,I205904,I110751,I110313,I110298,I110307,I110316,I110854,I110880,I110888,I110905,I110931,I110822,I110953,I110979,I110987,I111004,I111030,I110846,I111052,I110828,I111092,I111109,I111117,I111134,I110831,I111165,I111182,I111208,I111216,I110819,I110837,I111261,I111278,I110840,I110825,I110834,I110843,I111381,I448898,I111407,I111415,I448913,I111432,I448916,I111458,I111349,I111480,I448922,I111506,I111514,I448904,I111531,I111557,I111373,I111579,I111355,I448901,I111619,I111636,I111644,I111661,I111358,I111692,I448907,I111709,I448919,I111735,I111743,I111346,I111364,I111788,I448910,I111805,I111367,I111352,I111361,I111370,I111908,I458146,I111934,I111942,I458161,I111959,I458164,I111985,I111876,I112007,I458170,I112033,I112041,I458152,I112058,I112084,I111900,I112106,I111882,I458149,I112146,I112163,I112171,I112188,I111885,I112219,I458155,I112236,I458167,I112262,I112270,I111873,I111891,I112315,I458158,I112332,I111894,I111879,I111888,I111897,I112435,I349519,I112461,I112469,I349522,I349516,I112486,I349528,I112512,I112534,I349531,I112560,I112568,I112585,I112611,I112633,I349534,I112673,I112690,I112698,I112715,I112746,I349525,I112763,I112789,I112797,I112842,I349537,I112859,I112962,I230361,I112988,I112996,I230346,I230349,I113013,I230364,I113039,I112930,I113061,I230358,I113087,I113095,I113112,I113138,I112954,I113160,I112936,I230355,I113200,I113217,I113225,I113242,I112939,I113273,I230370,I113290,I230367,I113316,I113324,I112927,I112945,I113369,I230352,I113386,I112948,I112933,I112942,I112951,I113489,I113515,I113523,I113540,I113566,I113457,I113588,I113614,I113622,I113639,I113665,I113481,I113687,I113463,I113727,I113744,I113752,I113769,I113466,I113800,I113817,I113843,I113851,I113454,I113472,I113896,I113913,I113475,I113460,I113469,I113478,I114016,I114042,I114050,I114067,I114093,I113984,I114115,I114141,I114149,I114166,I114192,I114008,I114214,I113990,I114254,I114271,I114279,I114296,I113993,I114327,I114344,I114370,I114378,I113981,I113999,I114423,I114440,I114002,I113987,I113996,I114005,I114543,I522863,I114569,I114577,I522860,I522851,I114594,I522848,I114620,I114511,I114642,I522857,I114668,I114676,I522866,I114693,I114719,I114535,I114741,I114517,I522869,I114781,I114798,I114806,I114823,I114520,I114854,I522854,I114871,I522872,I114897,I114905,I114508,I114526,I114950,I114967,I114529,I114514,I114523,I114532,I115070,I356370,I115096,I115104,I356373,I356367,I115121,I356379,I115147,I115038,I115169,I356382,I115195,I115203,I115220,I115246,I115062,I115268,I115044,I356385,I115308,I115325,I115333,I115350,I115047,I115381,I356376,I115398,I115424,I115432,I115035,I115053,I115477,I356388,I115494,I115056,I115041,I115050,I115059,I115597,I115623,I115631,I115648,I115674,I115696,I115722,I115730,I115747,I115773,I115795,I115835,I115852,I115860,I115877,I115908,I115925,I115951,I115959,I116004,I116021,I116124,I483000,I116150,I116158,I483015,I116175,I483018,I116201,I116092,I116223,I483024,I116249,I116257,I483006,I116274,I116300,I116116,I116322,I116098,I483003,I116362,I116379,I116387,I116404,I116101,I116435,I483009,I116452,I483021,I116478,I116486,I116089,I116107,I116531,I483012,I116548,I116110,I116095,I116104,I116113,I116651,I314746,I116677,I116685,I314737,I314752,I116702,I314758,I116728,I116619,I116750,I314743,I116776,I116784,I116801,I116827,I116643,I116849,I116625,I314740,I116889,I116906,I116914,I116931,I116628,I116962,I314734,I314749,I116979,I117005,I117013,I116616,I116634,I117058,I314755,I117075,I116637,I116622,I116631,I116640,I117178,I117204,I117212,I117229,I117255,I117146,I117277,I117303,I117311,I117328,I117354,I117170,I117376,I117152,I117416,I117433,I117441,I117458,I117155,I117489,I117506,I117532,I117540,I117143,I117161,I117585,I117602,I117164,I117149,I117158,I117167,I117705,I474330,I117731,I117739,I474345,I117756,I474348,I117782,I117804,I474354,I117830,I117838,I474336,I117855,I117881,I117903,I474333,I117943,I117960,I117968,I117985,I118016,I474339,I118033,I474351,I118059,I118067,I118112,I474342,I118129,I118232,I360586,I118258,I118266,I360589,I360583,I118283,I360595,I118309,I118331,I360598,I118357,I118365,I118382,I118408,I118430,I360601,I118470,I118487,I118495,I118512,I118543,I360592,I118560,I118586,I118594,I118639,I360604,I118656,I118759,I533845,I118785,I118793,I533842,I533833,I118810,I533830,I118836,I118727,I118858,I533839,I118884,I118892,I533848,I118909,I118935,I118751,I118957,I118733,I533851,I118997,I119014,I119022,I119039,I118736,I119070,I533836,I119087,I533854,I119113,I119121,I118724,I118742,I119166,I119183,I118745,I118730,I118739,I118748,I119286,I119312,I119320,I119337,I119363,I119254,I119385,I119411,I119419,I119436,I119462,I119278,I119484,I119260,I119524,I119541,I119549,I119566,I119263,I119597,I119614,I119640,I119648,I119251,I119269,I119693,I119710,I119272,I119257,I119266,I119275,I119813,I493982,I119839,I119847,I493997,I119864,I494000,I119890,I119781,I119912,I494006,I119938,I119946,I493988,I119963,I119989,I119805,I120011,I119787,I493985,I120051,I120068,I120076,I120093,I119790,I120124,I493991,I120141,I494003,I120167,I120175,I119778,I119796,I120220,I493994,I120237,I119799,I119784,I119793,I119802,I120340,I229783,I120366,I120374,I229768,I229771,I120391,I229786,I120417,I120439,I229780,I120465,I120473,I120490,I120516,I120538,I229777,I120578,I120595,I120603,I120620,I120651,I229792,I120668,I229789,I120694,I120702,I120747,I229774,I120764,I120867,I350046,I120893,I120901,I350049,I350043,I120918,I350055,I120944,I120835,I120966,I350058,I120992,I121000,I121017,I121043,I120859,I121065,I120841,I350061,I121105,I121122,I121130,I121147,I120844,I121178,I350052,I121195,I121221,I121229,I120832,I120850,I121274,I350064,I121291,I120853,I120838,I120847,I120856,I121394,I562156,I121420,I121428,I562135,I121445,I562162,I121471,I121493,I562150,I121519,I121527,I562153,I121544,I121570,I121592,I562144,I121632,I121649,I121657,I121674,I121705,I562141,I562138,I121722,I562159,I121748,I121756,I121801,I562147,I121818,I121921,I121947,I121955,I121972,I121998,I121889,I122020,I122046,I122054,I122071,I122097,I121913,I122119,I121895,I122159,I122176,I122184,I122201,I121898,I122232,I122249,I122275,I122283,I121886,I121904,I122328,I122345,I121907,I121892,I121901,I121910,I122448,I338979,I122474,I122482,I338982,I338976,I122499,I338988,I122525,I122416,I122547,I338991,I122573,I122581,I122598,I122624,I122440,I122646,I122422,I338994,I122686,I122703,I122711,I122728,I122425,I122759,I338985,I122776,I122802,I122810,I122413,I122431,I122855,I338997,I122872,I122434,I122419,I122428,I122437,I122975,I247701,I123001,I123009,I247686,I247689,I123026,I247704,I123052,I123074,I247698,I123100,I123108,I123125,I123151,I123173,I247695,I123213,I123230,I123238,I123255,I123286,I247710,I123303,I247707,I123329,I123337,I123382,I247692,I123399,I123502,I543711,I123528,I123536,I543690,I123553,I543717,I123579,I123470,I123601,I543705,I123627,I123635,I543708,I123652,I123678,I123494,I123700,I123476,I543699,I123740,I123757,I123765,I123782,I123479,I123813,I543696,I543693,I123830,I543714,I123856,I123864,I123467,I123485,I123909,I543702,I123926,I123488,I123473,I123482,I123491,I124029,I535001,I124055,I124063,I534998,I534989,I124080,I534986,I124106,I123997,I124128,I534995,I124154,I124162,I535004,I124179,I124205,I124021,I124227,I124003,I535007,I124267,I124284,I124292,I124309,I124006,I124340,I534992,I124357,I535010,I124383,I124391,I123994,I124012,I124436,I124453,I124015,I124000,I124009,I124018,I124556,I338452,I124582,I124590,I338455,I338449,I124607,I338461,I124633,I124524,I124655,I338464,I124681,I124689,I124706,I124732,I124548,I124754,I124530,I338467,I124794,I124811,I124819,I124836,I124533,I124867,I338458,I124884,I124910,I124918,I124521,I124539,I124963,I338470,I124980,I124542,I124527,I124536,I124545,I125083,I444396,I125109,I125117,I444393,I125134,I444405,I125160,I125051,I125182,I125208,I125216,I444411,I125233,I125259,I125075,I125281,I125057,I444399,I125321,I125338,I125346,I125363,I125060,I125394,I444408,I444414,I125411,I125437,I125445,I125048,I125066,I125490,I444402,I125507,I125069,I125054,I125063,I125072,I125610,I510796,I125636,I125644,I510778,I510802,I125661,I510793,I125687,I125578,I125709,I510799,I125735,I125743,I510787,I125760,I125786,I125602,I125808,I125584,I125848,I125865,I125873,I125890,I125587,I125921,I510784,I510781,I125938,I510790,I125964,I125972,I125575,I125593,I126017,I126034,I125596,I125581,I125590,I125599,I126137,I168903,I126163,I126171,I168915,I168894,I126188,I168918,I126214,I126105,I126236,I168909,I126262,I126270,I168891,I126287,I126313,I126129,I126335,I126111,I168906,I126375,I126392,I126400,I126417,I126114,I126448,I168897,I126465,I168900,I126491,I126499,I126102,I126120,I126544,I168912,I126561,I126123,I126108,I126117,I126126,I126664,I537247,I126690,I126698,I537274,I537250,I126715,I537259,I126741,I126632,I126763,I126789,I126797,I537271,I126814,I126840,I126656,I126862,I126638,I537253,I126902,I126919,I126927,I126944,I126641,I126975,I537268,I537256,I126992,I537262,I127018,I127026,I126629,I126647,I127071,I537265,I127088,I126650,I126635,I126644,I126653,I127191,I274864,I127217,I127225,I274855,I274870,I127242,I274876,I127268,I127159,I127290,I274861,I127316,I127324,I127341,I127367,I127183,I127389,I127165,I274858,I127429,I127446,I127454,I127471,I127168,I127502,I274852,I274867,I127519,I127545,I127553,I127156,I127174,I127598,I274873,I127615,I127177,I127162,I127171,I127180,I127718,I388024,I127744,I127752,I388021,I388039,I127769,I388030,I127795,I127817,I388045,I127843,I127851,I388027,I127868,I127894,I127916,I388033,I127956,I127973,I127981,I127998,I128029,I388048,I128046,I388036,I128072,I128080,I128125,I388042,I128142,I128245,I175431,I128271,I128279,I175443,I175422,I128296,I175446,I128322,I128213,I128344,I175437,I128370,I128378,I175419,I128395,I128421,I128237,I128443,I128219,I175434,I128483,I128500,I128508,I128525,I128222,I128556,I175425,I128573,I175428,I128599,I128607,I128210,I128228,I128652,I175440,I128669,I128231,I128216,I128225,I128234,I128772,I128798,I128806,I128823,I128849,I128740,I128871,I128897,I128905,I128922,I128948,I128764,I128970,I128746,I129010,I129027,I129035,I129052,I128749,I129083,I129100,I129126,I129134,I128737,I128755,I129179,I129196,I128758,I128743,I128752,I128761,I129299,I329774,I129325,I129333,I329765,I329780,I129350,I329786,I129376,I129267,I129398,I329771,I129424,I129432,I129449,I129475,I129291,I129497,I129273,I329768,I129537,I129554,I129562,I129579,I129276,I129610,I329762,I329777,I129627,I129653,I129661,I129264,I129282,I129706,I329783,I129723,I129285,I129270,I129279,I129288,I129826,I505356,I129852,I129860,I505338,I505362,I129877,I505353,I129903,I129794,I129925,I505359,I129951,I129959,I505347,I129976,I130002,I129818,I130024,I129800,I130064,I130081,I130089,I130106,I129803,I130137,I505344,I505341,I130154,I505350,I130180,I130188,I129791,I129809,I130233,I130250,I129812,I129797,I129806,I129815,I130353,I130379,I130387,I130404,I130430,I130321,I130452,I130478,I130486,I130503,I130529,I130345,I130551,I130327,I130591,I130608,I130616,I130633,I130330,I130664,I130681,I130707,I130715,I130318,I130336,I130760,I130777,I130339,I130324,I130333,I130342,I130880,I486468,I130906,I130914,I486483,I130931,I486486,I130957,I130848,I130979,I486492,I131005,I131013,I486474,I131030,I131056,I130872,I131078,I130854,I486471,I131118,I131135,I131143,I131160,I130857,I131191,I486477,I131208,I486489,I131234,I131242,I130845,I130863,I131287,I486480,I131304,I130866,I130851,I130860,I130869,I131407,I288158,I131433,I131441,I288149,I288164,I131458,I288170,I131484,I131375,I131506,I288155,I131532,I131540,I131557,I131583,I131399,I131605,I131381,I288152,I131645,I131662,I131670,I131687,I131384,I131718,I288146,I288161,I131735,I131761,I131769,I131372,I131390,I131814,I288167,I131831,I131393,I131378,I131387,I131396,I131934,I229176,I131960,I131968,I229188,I131985,I229173,I132011,I131902,I132033,I229197,I132059,I132067,I229194,I132084,I132110,I131926,I132132,I131908,I229185,I132172,I132189,I132197,I132214,I131911,I132245,I229182,I132262,I229191,I132288,I132296,I131899,I131917,I132341,I229179,I132358,I131920,I131905,I131914,I131923,I132461,I400298,I132487,I132495,I400295,I400313,I132512,I400304,I132538,I132429,I132560,I400319,I132586,I132594,I400301,I132611,I132637,I132453,I132659,I132435,I400307,I132699,I132716,I132724,I132741,I132438,I132772,I400322,I132789,I400310,I132815,I132823,I132426,I132444,I132868,I400316,I132885,I132447,I132432,I132441,I132450,I132988,I280644,I133014,I133022,I280635,I280650,I133039,I280656,I133065,I132956,I133087,I280641,I133113,I133121,I133138,I133164,I132980,I133186,I132962,I280638,I133226,I133243,I133251,I133268,I132965,I133299,I280632,I280647,I133316,I133342,I133350,I132953,I132971,I133395,I280653,I133412,I132974,I132959,I132968,I132977,I133515,I133541,I133549,I133566,I133592,I133483,I133614,I133640,I133648,I133665,I133691,I133507,I133713,I133489,I133753,I133770,I133778,I133795,I133492,I133826,I133843,I133869,I133877,I133480,I133498,I133922,I133939,I133501,I133486,I133495,I133504,I134042,I134068,I134076,I134093,I134119,I134141,I134167,I134175,I134192,I134218,I134240,I134280,I134297,I134305,I134322,I134353,I134370,I134396,I134404,I134449,I134466,I134569,I300874,I134595,I134603,I300865,I300880,I134620,I300886,I134646,I134537,I134668,I300871,I134694,I134702,I134719,I134745,I134561,I134767,I134543,I300868,I134807,I134824,I134832,I134849,I134546,I134880,I300862,I300877,I134897,I134923,I134931,I134534,I134552,I134976,I300883,I134993,I134555,I134540,I134549,I134558,I135096,I328040,I135122,I135130,I328031,I328046,I135147,I328052,I135173,I135195,I328037,I135221,I135229,I135246,I135272,I135294,I328034,I135334,I135351,I135359,I135376,I135407,I328028,I328043,I135424,I135450,I135458,I135503,I328049,I135520,I135623,I384794,I135649,I135657,I384791,I384809,I135674,I384800,I135700,I135591,I135722,I384815,I135748,I135756,I384797,I135773,I135799,I135615,I135821,I135597,I384803,I135861,I135878,I135886,I135903,I135600,I135934,I384818,I135951,I384806,I135977,I135985,I135588,I135606,I136030,I384812,I136047,I135609,I135594,I135603,I135612,I136150,I278332,I136176,I136184,I278323,I278338,I136201,I278344,I136227,I136118,I136249,I278329,I136275,I136283,I136300,I136326,I136142,I136348,I136124,I278326,I136388,I136405,I136413,I136430,I136127,I136461,I278320,I278335,I136478,I136504,I136512,I136115,I136133,I136557,I278341,I136574,I136136,I136121,I136130,I136139,I136677,I443835,I136703,I136711,I443832,I136728,I443844,I136754,I136645,I136776,I136802,I136810,I443850,I136827,I136853,I136669,I136875,I136651,I443838,I136915,I136932,I136940,I136957,I136654,I136988,I443847,I443853,I137005,I137031,I137039,I136642,I136660,I137084,I443841,I137101,I136663,I136648,I136657,I136666,I137204,I137230,I137238,I137255,I137281,I137172,I137303,I137329,I137337,I137354,I137380,I137196,I137402,I137178,I137442,I137459,I137467,I137484,I137181,I137515,I137532,I137558,I137566,I137169,I137187,I137611,I137628,I137190,I137175,I137184,I137193,I137731,I341614,I137757,I137765,I341617,I341611,I137782,I341623,I137808,I137699,I137830,I341626,I137856,I137864,I137881,I137907,I137723,I137929,I137705,I341629,I137969,I137986,I137994,I138011,I137708,I138042,I341620,I138059,I138085,I138093,I137696,I137714,I138138,I341632,I138155,I137717,I137702,I137711,I137720,I138258,I138284,I138292,I138309,I138335,I138226,I138357,I138383,I138391,I138408,I138434,I138250,I138456,I138232,I138496,I138513,I138521,I138538,I138235,I138569,I138586,I138612,I138620,I138223,I138241,I138665,I138682,I138244,I138229,I138238,I138247,I138785,I336344,I138811,I138819,I336347,I336341,I138836,I336353,I138862,I138884,I336356,I138910,I138918,I138935,I138961,I138983,I336359,I139023,I139040,I139048,I139065,I139096,I336350,I139113,I139139,I139147,I139192,I336362,I139209,I139312,I139338,I139346,I139363,I139389,I139280,I139411,I139437,I139445,I139462,I139488,I139304,I139510,I139286,I139550,I139567,I139575,I139592,I139289,I139623,I139640,I139666,I139674,I139277,I139295,I139719,I139736,I139298,I139283,I139292,I139301,I139839,I558586,I139865,I139873,I558565,I139890,I558592,I139916,I139807,I139938,I558580,I139964,I139972,I558583,I139989,I140015,I139831,I140037,I139813,I558574,I140077,I140094,I140102,I140119,I139816,I140150,I558571,I558568,I140167,I558589,I140193,I140201,I139804,I139822,I140246,I558577,I140263,I139825,I139810,I139819,I139828,I140366,I140392,I140400,I140417,I140443,I140334,I140465,I140491,I140499,I140516,I140542,I140358,I140564,I140340,I140604,I140621,I140629,I140646,I140343,I140677,I140694,I140720,I140728,I140331,I140349,I140773,I140790,I140352,I140337,I140346,I140355,I140893,I252903,I140919,I140927,I252888,I252891,I140944,I252906,I140970,I140861,I140992,I252900,I141018,I141026,I141043,I141069,I140885,I141091,I140867,I252897,I141131,I141148,I141156,I141173,I140870,I141204,I252912,I141221,I252909,I141247,I141255,I140858,I140876,I141300,I252894,I141317,I140879,I140864,I140873,I140882,I141420,I141446,I141454,I141471,I141497,I141388,I141519,I141545,I141553,I141570,I141596,I141412,I141618,I141394,I141658,I141675,I141683,I141700,I141397,I141731,I141748,I141774,I141782,I141385,I141403,I141827,I141844,I141406,I141391,I141400,I141409,I141947,I141973,I141981,I141998,I142024,I141915,I142046,I142072,I142080,I142097,I142123,I141939,I142145,I141921,I142185,I142202,I142210,I142227,I141924,I142258,I142275,I142301,I142309,I141912,I141930,I142354,I142371,I141933,I141918,I141927,I141936,I142474,I142500,I142508,I142525,I142551,I142442,I142573,I142599,I142607,I142624,I142650,I142466,I142672,I142448,I142712,I142729,I142737,I142754,I142451,I142785,I142802,I142828,I142836,I142439,I142457,I142881,I142898,I142460,I142445,I142454,I142463,I143001,I185223,I143027,I143035,I185235,I185214,I143052,I185238,I143078,I142969,I143100,I185229,I143126,I143134,I185211,I143151,I143177,I142993,I143199,I142975,I185226,I143239,I143256,I143264,I143281,I142978,I143312,I185217,I143329,I185220,I143355,I143363,I142966,I142984,I143408,I185232,I143425,I142987,I142972,I142981,I142990,I143528,I172167,I143554,I143562,I172179,I172158,I143579,I172182,I143605,I143496,I143627,I172173,I143653,I143661,I172155,I143678,I143704,I143520,I143726,I143502,I172170,I143766,I143783,I143791,I143808,I143505,I143839,I172161,I143856,I172164,I143882,I143890,I143493,I143511,I143935,I172176,I143952,I143514,I143499,I143508,I143517,I144055,I432615,I144081,I144089,I432612,I144106,I432624,I144132,I144023,I144154,I144180,I144188,I432630,I144205,I144231,I144047,I144253,I144029,I432618,I144293,I144310,I144318,I144335,I144032,I144366,I432627,I432633,I144383,I144409,I144417,I144020,I144038,I144462,I432621,I144479,I144041,I144026,I144035,I144044,I144582,I563941,I144608,I144616,I563920,I144633,I563947,I144659,I144681,I563935,I144707,I144715,I563938,I144732,I144758,I144780,I563929,I144820,I144837,I144845,I144862,I144893,I563926,I563923,I144910,I563944,I144936,I144944,I144989,I563932,I145006,I145109,I299718,I145135,I145143,I299709,I299724,I145160,I299730,I145186,I145077,I145208,I299715,I145234,I145242,I145259,I145285,I145101,I145307,I145083,I299712,I145347,I145364,I145372,I145389,I145086,I145420,I299706,I299721,I145437,I145463,I145471,I145074,I145092,I145516,I299727,I145533,I145095,I145080,I145089,I145098,I145636,I145662,I145670,I145687,I145713,I145735,I145761,I145769,I145786,I145812,I145834,I145874,I145891,I145899,I145916,I145947,I145964,I145990,I145998,I146043,I146060,I146163,I146189,I146197,I146214,I146240,I146262,I146288,I146296,I146313,I146339,I146361,I146401,I146418,I146426,I146443,I146474,I146491,I146517,I146525,I146570,I146587,I146690,I405466,I146716,I146724,I405463,I405481,I146741,I405472,I146767,I146789,I405487,I146815,I146823,I405469,I146840,I146866,I146888,I405475,I146928,I146945,I146953,I146970,I147001,I405490,I147018,I405478,I147044,I147052,I147097,I405484,I147114,I147217,I552041,I147243,I147251,I552020,I147268,I552047,I147294,I147185,I147316,I552035,I147342,I147350,I552038,I147367,I147393,I147209,I147415,I147191,I552029,I147455,I147472,I147480,I147497,I147194,I147528,I552026,I552023,I147545,I552044,I147571,I147579,I147182,I147200,I147624,I552032,I147641,I147203,I147188,I147197,I147206,I147744,I200999,I147770,I147778,I201011,I200990,I147795,I201014,I147821,I147712,I147843,I201005,I147869,I147877,I200987,I147894,I147920,I147736,I147942,I147718,I201002,I147982,I147999,I148007,I148024,I147721,I148055,I200993,I148072,I200996,I148098,I148106,I147709,I147727,I148151,I201008,I148168,I147730,I147715,I147724,I147733,I148271,I206983,I148297,I148305,I206995,I206974,I148322,I206998,I148348,I148239,I148370,I206989,I148396,I148404,I206971,I148421,I148447,I148263,I148469,I148245,I206986,I148509,I148526,I148534,I148551,I148248,I148582,I206977,I148599,I206980,I148625,I148633,I148236,I148254,I148678,I206992,I148695,I148257,I148242,I148251,I148260,I148798,I487624,I148824,I148832,I487639,I148849,I487642,I148875,I148897,I487648,I148923,I148931,I487630,I148948,I148974,I148996,I487627,I149036,I149053,I149061,I149078,I149109,I487633,I149126,I487645,I149152,I149160,I149205,I487636,I149222,I149325,I149351,I149359,I149376,I149402,I149424,I149450,I149458,I149475,I149501,I149523,I149563,I149580,I149588,I149605,I149636,I149653,I149679,I149687,I149732,I149749,I149852,I149878,I149886,I149903,I149929,I149820,I149951,I149977,I149985,I150002,I150028,I149844,I150050,I149826,I150090,I150107,I150115,I150132,I149829,I150163,I150180,I150206,I150214,I149817,I149835,I150259,I150276,I149838,I149823,I149832,I149841,I150379,I410634,I150405,I150413,I410631,I410649,I150430,I410640,I150456,I150478,I410655,I150504,I150512,I410637,I150529,I150555,I150577,I410643,I150617,I150634,I150642,I150659,I150690,I410658,I150707,I410646,I150733,I150741,I150786,I410652,I150803,I150906,I490514,I150932,I150940,I490529,I150957,I490532,I150983,I151005,I490538,I151031,I151039,I490520,I151056,I151082,I151104,I490517,I151144,I151161,I151169,I151186,I151217,I490523,I151234,I490535,I151260,I151268,I151313,I490526,I151330,I151433,I239031,I151459,I151467,I239016,I239019,I151484,I239034,I151510,I151401,I151532,I239028,I151558,I151566,I151583,I151609,I151425,I151631,I151407,I239025,I151671,I151688,I151696,I151713,I151410,I151744,I239040,I151761,I239037,I151787,I151795,I151398,I151416,I151840,I239022,I151857,I151419,I151404,I151413,I151422,I151960,I269084,I151986,I151994,I269075,I269090,I152011,I269096,I152037,I152059,I269081,I152085,I152093,I152110,I152136,I152158,I269078,I152198,I152215,I152223,I152240,I152271,I269072,I269087,I152288,I152314,I152322,I152367,I269093,I152384,I152487,I563346,I152513,I152521,I563325,I152538,I563352,I152564,I152455,I152586,I563340,I152612,I152620,I563343,I152637,I152663,I152479,I152685,I152461,I563334,I152725,I152742,I152750,I152767,I152464,I152798,I563331,I563328,I152815,I563349,I152841,I152849,I152452,I152470,I152894,I563337,I152911,I152473,I152458,I152467,I152476,I153014,I480110,I153040,I153048,I480125,I153065,I480128,I153091,I152982,I153113,I480134,I153139,I153147,I480116,I153164,I153190,I153006,I153212,I152988,I480113,I153252,I153269,I153277,I153294,I152991,I153325,I480119,I153342,I480131,I153368,I153376,I152979,I152997,I153421,I480122,I153438,I153000,I152985,I152994,I153003,I153541,I165639,I153567,I153575,I165651,I165630,I153592,I165654,I153618,I153509,I153640,I165645,I153666,I153674,I165627,I153691,I153717,I153533,I153739,I153515,I165642,I153779,I153796,I153804,I153821,I153518,I153852,I165633,I153869,I165636,I153895,I153903,I153506,I153524,I153948,I165648,I153965,I153527,I153512,I153521,I153530,I154068,I184135,I154094,I154102,I184147,I184126,I154119,I184150,I154145,I154036,I154167,I184141,I154193,I154201,I184123,I154218,I154244,I154060,I154266,I154042,I184138,I154306,I154323,I154331,I154348,I154045,I154379,I184129,I154396,I184132,I154422,I154430,I154033,I154051,I154475,I184144,I154492,I154054,I154039,I154048,I154057,I154595,I242499,I154621,I154629,I242484,I242487,I154646,I242502,I154672,I154563,I154694,I242496,I154720,I154728,I154745,I154771,I154587,I154793,I154569,I242493,I154833,I154850,I154858,I154875,I154572,I154906,I242508,I154923,I242505,I154949,I154957,I154560,I154578,I155002,I242490,I155019,I154581,I154566,I154575,I154584,I155122,I370599,I155148,I155156,I370602,I370596,I155173,I370608,I155199,I155221,I370611,I155247,I155255,I155272,I155298,I155320,I370614,I155360,I155377,I155385,I155402,I155433,I370605,I155450,I155476,I155484,I155529,I370617,I155546,I155649,I269662,I155675,I155683,I269653,I269668,I155700,I269674,I155726,I155617,I155748,I269659,I155774,I155782,I155799,I155825,I155641,I155847,I155623,I269656,I155887,I155904,I155912,I155929,I155626,I155960,I269650,I269665,I155977,I156003,I156011,I155614,I155632,I156056,I269671,I156073,I155635,I155620,I155629,I155638,I156176,I461036,I156202,I156210,I461051,I156227,I461054,I156253,I156275,I461060,I156301,I156309,I461042,I156326,I156352,I156374,I461039,I156414,I156431,I156439,I156456,I156487,I461045,I156504,I461057,I156530,I156538,I156583,I461048,I156600,I156703,I498606,I156729,I156737,I498621,I156754,I498624,I156780,I156671,I156802,I498630,I156828,I156836,I498612,I156853,I156879,I156695,I156901,I156677,I498609,I156941,I156958,I156966,I156983,I156680,I157014,I498615,I157031,I498627,I157057,I157065,I156668,I156686,I157110,I498618,I157127,I156689,I156674,I156683,I156692,I157230,I515148,I157256,I157264,I515130,I515154,I157281,I515145,I157307,I157329,I515151,I157355,I157363,I515139,I157380,I157406,I157428,I157468,I157485,I157493,I157510,I157541,I515136,I515133,I157558,I515142,I157584,I157592,I157637,I157654,I157757,I157783,I157791,I157808,I157834,I157725,I157856,I157882,I157890,I157907,I157933,I157749,I157955,I157731,I157995,I158012,I158020,I158037,I157734,I158068,I158085,I158111,I158119,I157722,I157740,I158164,I158181,I157743,I157728,I157737,I157746,I158284,I425883,I158310,I158318,I425880,I158335,I425892,I158361,I158252,I158383,I158409,I158417,I425898,I158434,I158460,I158276,I158482,I158258,I425886,I158522,I158539,I158547,I158564,I158261,I158595,I425895,I425901,I158612,I158638,I158646,I158249,I158267,I158691,I425889,I158708,I158270,I158255,I158264,I158273,I158811,I422262,I158837,I158845,I422259,I422277,I158862,I422268,I158888,I158910,I422283,I158936,I158944,I422265,I158961,I158987,I159009,I422271,I159049,I159066,I159074,I159091,I159122,I422286,I159139,I422274,I159165,I159173,I159218,I422280,I159235,I159338,I477798,I159364,I159372,I477813,I159389,I477816,I159415,I159306,I159437,I477822,I159463,I159471,I477804,I159488,I159514,I159330,I159536,I159312,I477801,I159576,I159593,I159601,I159618,I159315,I159649,I477807,I159666,I477819,I159692,I159700,I159303,I159321,I159745,I477810,I159762,I159324,I159309,I159318,I159327,I159865,I404820,I159891,I159899,I404817,I404835,I159916,I404826,I159942,I159833,I159964,I404841,I159990,I159998,I404823,I160015,I160041,I159857,I160063,I159839,I404829,I160103,I160120,I160128,I160145,I159842,I160176,I404844,I160193,I404832,I160219,I160227,I159830,I159848,I160272,I404838,I160289,I159851,I159836,I159845,I159854,I160392,I372180,I160418,I160426,I372183,I372177,I160443,I372189,I160469,I160360,I160491,I372192,I160517,I160525,I160542,I160568,I160384,I160590,I160366,I372195,I160630,I160647,I160655,I160672,I160369,I160703,I372186,I160720,I160746,I160754,I160357,I160375,I160799,I372198,I160816,I160378,I160363,I160372,I160381,I160919,I296828,I160945,I160953,I296819,I296834,I160970,I296840,I160996,I160887,I161018,I296825,I161044,I161052,I161069,I161095,I160911,I161117,I160893,I296822,I161157,I161174,I161182,I161199,I160896,I161230,I296816,I296831,I161247,I161273,I161281,I160884,I160902,I161326,I296837,I161343,I160905,I160890,I160899,I160908,I161446,I492826,I161472,I161480,I492841,I161497,I492844,I161523,I161545,I492850,I161571,I161579,I492832,I161596,I161622,I161644,I492829,I161684,I161701,I161709,I161726,I161757,I492835,I161774,I492847,I161800,I161808,I161853,I492838,I161870,I161973,I452944,I161999,I162007,I452959,I162024,I452962,I162050,I161941,I162072,I452968,I162098,I162106,I452950,I162123,I162149,I161965,I162171,I161947,I452947,I162211,I162228,I162236,I162253,I161950,I162284,I452953,I162301,I452965,I162327,I162335,I161938,I161956,I162380,I452956,I162397,I161959,I161944,I161953,I161962,I162500,I198279,I162526,I162534,I198291,I198270,I162551,I198294,I162577,I162599,I198285,I162625,I162633,I198267,I162650,I162676,I162698,I198282,I162738,I162755,I162763,I162780,I162811,I198273,I162828,I198276,I162854,I162862,I162907,I198288,I162924,I163027,I163053,I163061,I163078,I163104,I162995,I163126,I163152,I163160,I163177,I163203,I163019,I163225,I163001,I163265,I163282,I163290,I163307,I163004,I163338,I163355,I163381,I163389,I162992,I163010,I163434,I163451,I163013,I162998,I163007,I163016,I163554,I313012,I163580,I163588,I313003,I313018,I163605,I313024,I163631,I163653,I313009,I163679,I163687,I163704,I163730,I163752,I313006,I163792,I163809,I163817,I163834,I163865,I313000,I313015,I163882,I163908,I163916,I163961,I313021,I163978,I164081,I291048,I164107,I164115,I291039,I291054,I164132,I291060,I164158,I164180,I291045,I164206,I164214,I164231,I164257,I164279,I291042,I164319,I164336,I164344,I164361,I164392,I291036,I291051,I164409,I164435,I164443,I164488,I291057,I164505,I164608,I384148,I164634,I164642,I384145,I384163,I164659,I384154,I164685,I164707,I384169,I164733,I164741,I384151,I164758,I164784,I164806,I384157,I164846,I164863,I164871,I164888,I164919,I384172,I164936,I384160,I164962,I164970,I165015,I384166,I165032,I165135,I404174,I165161,I165169,I404171,I404189,I165186,I404180,I165212,I165234,I404195,I165260,I165268,I404177,I165285,I165311,I165333,I404183,I165373,I165390,I165398,I165415,I165446,I404198,I165463,I404186,I165489,I165497,I165542,I404192,I165559,I165662,I260405,I165688,I165705,I165727,I165744,I260402,I260423,I165761,I260426,I165787,I165795,I260411,I165821,I165829,I260414,I165846,I260417,I165886,I165894,I165939,I260408,I165956,I260420,I165982,I166004,I166021,I166038,I166069,I166086,I166117,I166206,I215491,I166232,I166249,I166198,I166271,I166288,I215494,I215512,I166305,I215500,I166331,I166339,I166365,I166373,I215509,I166390,I166177,I215503,I166430,I166438,I166171,I166186,I166483,I215506,I215488,I166500,I215497,I166526,I166174,I166548,I166565,I166582,I166189,I166613,I166630,I166180,I166661,I166183,I166195,I166192,I166750,I166776,I166793,I166742,I166815,I166832,I166849,I166875,I166883,I166909,I166917,I166934,I166721,I166974,I166982,I166715,I166730,I167027,I167044,I167070,I166718,I167092,I167109,I167126,I166733,I167157,I167174,I166724,I167205,I166727,I166739,I166736,I167294,I445515,I167320,I167337,I167286,I167359,I167376,I445533,I167393,I445527,I167419,I167427,I445521,I167453,I167461,I445530,I167478,I167265,I445518,I167518,I167526,I167259,I167274,I167571,I445536,I167588,I167614,I167262,I167636,I167653,I167670,I167277,I167701,I167718,I445524,I167268,I167749,I167271,I167283,I167280,I167838,I484737,I167864,I167881,I167903,I167920,I484749,I167937,I484740,I167963,I167971,I484758,I167997,I168005,I484734,I168022,I484752,I168062,I168070,I168115,I484746,I484743,I168132,I484755,I168158,I168180,I168197,I168214,I168245,I168262,I168293,I168382,I237285,I168408,I168425,I168374,I168447,I168464,I237282,I237303,I168481,I237306,I168507,I168515,I237291,I168541,I168549,I237294,I168566,I168353,I237297,I168606,I168614,I168347,I168362,I168659,I237288,I168676,I237300,I168702,I168350,I168724,I168741,I168758,I168365,I168789,I168806,I168356,I168837,I168359,I168371,I168368,I168926,I168952,I168969,I168991,I169008,I169025,I169051,I169059,I169085,I169093,I169110,I169150,I169158,I169203,I169220,I169246,I169268,I169285,I169302,I169333,I169350,I169381,I169470,I256937,I169496,I169513,I169462,I169535,I169552,I256934,I256955,I169569,I256958,I169595,I169603,I256943,I169629,I169637,I256946,I169654,I169441,I256949,I169694,I169702,I169435,I169450,I169747,I256940,I169764,I256952,I169790,I169438,I169812,I169829,I169846,I169453,I169877,I169894,I169444,I169925,I169447,I169459,I169456,I170014,I306067,I170040,I170057,I170006,I170079,I170096,I306088,I306079,I170113,I170139,I170147,I306073,I170173,I170181,I306070,I170198,I169985,I306064,I170238,I170246,I169979,I169994,I170291,I306076,I170308,I306085,I170334,I169982,I170356,I170373,I170390,I169997,I170421,I170438,I306082,I169988,I170469,I169991,I170003,I170000,I170558,I281213,I170584,I170601,I170550,I170623,I170640,I281234,I281225,I170657,I170683,I170691,I281219,I170717,I170725,I281216,I170742,I170529,I281210,I170782,I170790,I170523,I170538,I170835,I281222,I170852,I281231,I170878,I170526,I170900,I170917,I170934,I170541,I170965,I170982,I281228,I170532,I171013,I170535,I170547,I170544,I171102,I171128,I171145,I171094,I171167,I171184,I171201,I171227,I171235,I171261,I171269,I171286,I171073,I171326,I171334,I171067,I171082,I171379,I171396,I171422,I171070,I171444,I171461,I171478,I171085,I171509,I171526,I171076,I171557,I171079,I171091,I171088,I171646,I171672,I171689,I171638,I171711,I171728,I171745,I171771,I171779,I171805,I171813,I171830,I171617,I171870,I171878,I171611,I171626,I171923,I171940,I171966,I171614,I171988,I172005,I172022,I171629,I172053,I172070,I171620,I172101,I171623,I171635,I171632,I172190,I509149,I172216,I172233,I172255,I172272,I509161,I509164,I172289,I509167,I172315,I172323,I509152,I172349,I172357,I509158,I172374,I509146,I172414,I172422,I172467,I509170,I172484,I509155,I172510,I172532,I172549,I172566,I172597,I172614,I172645,I172734,I491095,I172760,I172777,I172799,I172816,I491107,I172833,I491098,I172859,I172867,I491116,I172893,I172901,I491092,I172918,I491110,I172958,I172966,I173011,I491104,I491101,I173028,I491113,I173054,I173076,I173093,I173110,I173141,I173158,I173189,I173278,I173304,I173321,I173270,I173343,I173360,I173377,I173403,I173411,I173437,I173445,I173462,I173249,I173502,I173510,I173243,I173258,I173555,I173572,I173598,I173246,I173620,I173637,I173654,I173261,I173685,I173702,I173252,I173733,I173255,I173267,I173264,I173822,I173848,I173865,I173814,I173887,I173904,I173921,I173947,I173955,I173981,I173989,I174006,I173793,I174046,I174054,I173787,I173802,I174099,I174116,I174142,I173790,I174164,I174181,I174198,I173805,I174229,I174246,I173796,I174277,I173799,I173811,I173808,I174366,I408699,I174392,I174409,I174358,I174431,I174448,I408714,I408702,I174465,I408693,I174491,I174499,I408705,I174525,I174533,I408696,I174550,I174337,I408711,I174590,I174598,I174331,I174346,I174643,I408720,I408708,I174660,I408717,I174686,I174334,I174708,I174725,I174742,I174349,I174773,I174790,I174340,I174821,I174343,I174355,I174352,I174910,I174936,I174953,I174902,I174975,I174992,I175009,I175035,I175043,I175069,I175077,I175094,I174881,I175134,I175142,I174875,I174890,I175187,I175204,I175230,I174878,I175252,I175269,I175286,I174893,I175317,I175334,I174884,I175365,I174887,I174899,I174896,I175454,I175480,I175497,I175519,I175536,I175553,I175579,I175587,I175613,I175621,I175638,I175678,I175686,I175731,I175748,I175774,I175796,I175813,I175830,I175861,I175878,I175909,I175998,I517309,I176024,I176041,I175990,I176063,I176080,I517321,I517324,I176097,I517327,I176123,I176131,I517312,I176157,I176165,I517318,I176182,I175969,I517306,I176222,I176230,I175963,I175978,I176275,I517330,I176292,I517315,I176318,I175966,I176340,I176357,I176374,I175981,I176405,I176422,I175972,I176453,I175975,I175987,I175984,I176542,I450635,I176568,I176585,I176607,I176624,I450647,I176641,I450638,I176667,I176675,I450656,I176701,I176709,I450632,I176726,I450650,I176766,I176774,I176819,I450644,I450641,I176836,I450653,I176862,I176884,I176901,I176918,I176949,I176966,I176997,I177086,I496297,I177112,I177129,I177078,I177151,I177168,I496309,I177185,I496300,I177211,I177219,I496318,I177245,I177253,I496294,I177270,I177057,I496312,I177310,I177318,I177051,I177066,I177363,I496306,I496303,I177380,I496315,I177406,I177054,I177428,I177445,I177462,I177069,I177493,I177510,I177060,I177541,I177063,I177075,I177072,I177630,I525178,I177656,I177673,I177622,I177695,I177712,I525175,I525172,I177729,I525160,I177755,I177763,I525184,I177789,I177797,I525169,I177814,I177601,I525163,I177854,I177862,I177595,I177610,I177907,I525166,I177924,I525181,I177950,I177598,I177972,I177989,I178006,I177613,I178037,I178054,I177604,I178085,I177607,I177619,I177616,I178174,I178200,I178217,I178166,I178239,I178256,I178273,I178299,I178307,I178333,I178341,I178358,I178145,I178398,I178406,I178139,I178154,I178451,I178468,I178494,I178142,I178516,I178533,I178550,I178157,I178581,I178598,I178148,I178629,I178151,I178163,I178160,I178718,I322251,I178744,I178761,I178710,I178783,I178800,I322272,I322263,I178817,I178843,I178851,I322257,I178877,I178885,I322254,I178902,I178689,I322248,I178942,I178950,I178683,I178698,I178995,I322260,I179012,I322269,I179038,I178686,I179060,I179077,I179094,I178701,I179125,I179142,I322266,I178692,I179173,I178695,I178707,I178704,I179262,I179288,I179305,I179254,I179327,I179344,I179361,I179387,I179395,I179421,I179429,I179446,I179233,I179486,I179494,I179227,I179242,I179539,I179556,I179582,I179230,I179604,I179621,I179638,I179245,I179669,I179686,I179236,I179717,I179239,I179251,I179248,I179806,I289883,I179832,I179849,I179798,I179871,I179888,I289904,I289895,I179905,I179931,I179939,I289889,I179965,I179973,I289886,I179990,I179777,I289880,I180030,I180038,I179771,I179786,I180083,I289892,I180100,I289901,I180126,I179774,I180148,I180165,I180182,I179789,I180213,I180230,I289898,I179780,I180261,I179783,I179795,I179792,I180350,I411283,I180376,I180393,I180342,I180415,I180432,I411298,I411286,I180449,I411277,I180475,I180483,I411289,I180509,I180517,I411280,I180534,I180321,I411295,I180574,I180582,I180315,I180330,I180627,I411304,I411292,I180644,I411301,I180670,I180318,I180692,I180709,I180726,I180333,I180757,I180774,I180324,I180805,I180327,I180339,I180336,I180894,I391903,I180920,I180937,I180959,I180976,I391918,I391906,I180993,I391897,I181019,I181027,I391909,I181053,I181061,I391900,I181078,I391915,I181118,I181126,I181171,I391924,I391912,I181188,I391921,I181214,I181236,I181253,I181270,I181301,I181318,I181349,I181438,I450057,I181464,I181481,I181430,I181503,I181520,I450069,I181537,I450060,I181563,I181571,I450078,I181597,I181605,I450054,I181622,I181409,I450072,I181662,I181670,I181403,I181418,I181715,I450066,I450063,I181732,I450075,I181758,I181406,I181780,I181797,I181814,I181421,I181845,I181862,I181412,I181893,I181415,I181427,I181424,I181982,I489939,I182008,I182025,I181974,I182047,I182064,I489951,I182081,I489942,I182107,I182115,I489960,I182141,I182149,I489936,I182166,I181953,I489954,I182206,I182214,I181947,I181962,I182259,I489948,I489945,I182276,I489957,I182302,I181950,I182324,I182341,I182358,I181965,I182389,I182406,I181956,I182437,I181959,I181971,I181968,I182526,I182552,I182569,I182518,I182591,I182608,I182625,I182651,I182659,I182685,I182693,I182710,I182497,I182750,I182758,I182491,I182506,I182803,I182820,I182846,I182494,I182868,I182885,I182902,I182509,I182933,I182950,I182500,I182981,I182503,I182515,I182512,I183070,I301443,I183096,I183113,I183062,I183135,I183152,I301464,I301455,I183169,I183195,I183203,I301449,I183229,I183237,I301446,I183254,I183041,I301440,I183294,I183302,I183035,I183050,I183347,I301452,I183364,I301461,I183390,I183038,I183412,I183429,I183446,I183053,I183477,I183494,I301458,I183044,I183525,I183047,I183059,I183056,I183614,I226201,I183640,I183657,I183606,I183679,I183696,I226204,I226222,I183713,I226210,I183739,I183747,I183773,I183781,I226219,I183798,I183585,I226213,I183838,I183846,I183579,I183594,I183891,I226216,I226198,I183908,I226207,I183934,I183582,I183956,I183973,I183990,I183597,I184021,I184038,I183588,I184069,I183591,I183603,I183600,I184158,I214301,I184184,I184201,I184223,I184240,I214304,I214322,I184257,I214310,I184283,I184291,I184317,I184325,I214319,I184342,I214313,I184382,I184390,I184435,I214316,I214298,I184452,I214307,I184478,I184500,I184517,I184534,I184565,I184582,I184613,I184702,I184728,I184745,I184767,I184784,I184801,I184827,I184835,I184861,I184869,I184886,I184926,I184934,I184979,I184996,I185022,I185044,I185061,I185078,I185109,I185126,I185157,I185246,I185272,I185289,I185311,I185328,I185345,I185371,I185379,I185405,I185413,I185430,I185470,I185478,I185523,I185540,I185566,I185588,I185605,I185622,I185653,I185670,I185701,I185790,I395133,I185816,I185833,I185782,I185855,I185872,I395148,I395136,I185889,I395127,I185915,I185923,I395139,I185949,I185957,I395130,I185974,I185761,I395145,I186014,I186022,I185755,I185770,I186067,I395154,I395142,I186084,I395151,I186110,I185758,I186132,I186149,I186166,I185773,I186197,I186214,I185764,I186245,I185767,I185779,I185776,I186334,I378983,I186360,I186377,I186326,I186399,I186416,I378998,I378986,I186433,I378977,I186459,I186467,I378989,I186493,I186501,I378980,I186518,I186305,I378995,I186558,I186566,I186299,I186314,I186611,I379004,I378992,I186628,I379001,I186654,I186302,I186676,I186693,I186710,I186317,I186741,I186758,I186308,I186789,I186311,I186323,I186320,I186878,I186904,I186921,I186870,I186943,I186960,I186977,I187003,I187011,I187037,I187045,I187062,I186849,I187102,I187110,I186843,I186858,I187155,I187172,I187198,I186846,I187220,I187237,I187254,I186861,I187285,I187302,I186852,I187333,I186855,I186867,I186864,I187422,I187448,I187465,I187414,I187487,I187504,I187521,I187547,I187555,I187581,I187589,I187606,I187393,I187646,I187654,I187387,I187402,I187699,I187716,I187742,I187390,I187764,I187781,I187798,I187405,I187829,I187846,I187396,I187877,I187399,I187411,I187408,I187966,I187992,I188009,I187958,I188031,I188048,I188065,I188091,I188099,I188125,I188133,I188150,I187937,I188190,I188198,I187931,I187946,I188243,I188260,I188286,I187934,I188308,I188325,I188342,I187949,I188373,I188390,I187940,I188421,I187943,I187955,I187952,I188510,I188536,I188553,I188502,I188575,I188592,I188609,I188635,I188643,I188669,I188677,I188694,I188481,I188734,I188742,I188475,I188490,I188787,I188804,I188830,I188478,I188852,I188869,I188886,I188493,I188917,I188934,I188484,I188965,I188487,I188499,I188496,I189054,I189080,I189097,I189046,I189119,I189136,I189153,I189179,I189187,I189213,I189221,I189238,I189025,I189278,I189286,I189019,I189034,I189331,I189348,I189374,I189022,I189396,I189413,I189430,I189037,I189461,I189478,I189028,I189509,I189031,I189043,I189040,I189598,I402885,I189624,I189641,I189590,I189663,I189680,I402900,I402888,I189697,I402879,I189723,I189731,I402891,I189757,I189765,I402882,I189782,I189569,I402897,I189822,I189830,I189563,I189578,I189875,I402906,I402894,I189892,I402903,I189918,I189566,I189940,I189957,I189974,I189581,I190005,I190022,I189572,I190053,I189575,I189587,I189584,I190142,I220251,I190168,I190185,I190207,I190224,I220254,I220272,I190241,I220260,I190267,I190275,I190301,I190309,I220269,I190326,I220263,I190366,I190374,I190419,I220266,I220248,I190436,I220257,I190462,I190484,I190501,I190518,I190549,I190566,I190597,I190686,I541337,I190712,I190729,I190751,I190768,I541313,I541334,I190785,I541331,I190811,I190819,I541310,I190845,I190853,I541322,I190870,I541325,I190910,I190918,I190963,I541328,I541316,I190980,I541319,I191006,I191028,I191045,I191062,I191093,I191110,I191141,I191230,I523444,I191256,I191273,I191295,I191312,I523441,I523438,I191329,I523426,I191355,I191363,I523450,I191389,I191397,I523435,I191414,I523429,I191454,I191462,I191507,I523432,I191524,I523447,I191550,I191572,I191589,I191606,I191637,I191654,I191685,I191774,I409991,I191800,I191817,I191839,I191856,I410006,I409994,I191873,I409985,I191899,I191907,I409997,I191933,I191941,I409988,I191958,I410003,I191998,I192006,I192051,I410012,I410000,I192068,I410009,I192094,I192116,I192133,I192150,I192181,I192198,I192229,I192318,I192344,I192361,I192310,I192383,I192400,I192417,I192443,I192451,I192477,I192485,I192502,I192289,I192542,I192550,I192283,I192298,I192595,I192612,I192638,I192286,I192660,I192677,I192694,I192301,I192725,I192742,I192292,I192773,I192295,I192307,I192304,I192862,I192888,I192905,I192927,I192944,I192961,I192987,I192995,I193021,I193029,I193046,I193086,I193094,I193139,I193156,I193182,I193204,I193221,I193238,I193269,I193286,I193317,I193406,I252313,I193432,I193449,I193398,I193471,I193488,I252310,I252331,I193505,I252334,I193531,I193539,I252319,I193565,I193573,I252322,I193590,I193377,I252325,I193630,I193638,I193371,I193386,I193683,I252316,I193700,I252328,I193726,I193374,I193748,I193765,I193782,I193389,I193813,I193830,I193380,I193861,I193383,I193395,I193392,I193950,I395779,I193976,I193993,I193942,I194015,I194032,I395794,I395782,I194049,I395773,I194075,I194083,I395785,I194109,I194117,I395776,I194134,I193921,I395791,I194174,I194182,I193915,I193930,I194227,I395800,I395788,I194244,I395797,I194270,I193918,I194292,I194309,I194326,I193933,I194357,I194374,I193924,I194405,I193927,I193939,I193936,I194494,I241909,I194520,I194537,I194486,I194559,I194576,I241906,I241927,I194593,I241930,I194619,I194627,I241915,I194653,I194661,I241918,I194678,I194465,I241921,I194718,I194726,I194459,I194474,I194771,I241912,I194788,I241924,I194814,I194462,I194836,I194853,I194870,I194477,I194901,I194918,I194468,I194949,I194471,I194483,I194480,I195038,I346893,I195064,I195081,I195030,I195103,I195120,I346887,I346884,I195137,I346899,I195163,I195171,I195197,I195205,I346881,I195222,I195009,I195262,I195270,I195003,I195018,I195315,I346896,I346890,I195332,I195358,I195006,I195380,I195397,I195414,I195021,I195445,I195462,I346902,I195012,I195493,I195015,I195027,I195024,I195582,I294507,I195608,I195625,I195574,I195647,I195664,I294528,I294519,I195681,I195707,I195715,I294513,I195741,I195749,I294510,I195766,I195553,I294504,I195806,I195814,I195547,I195562,I195859,I294516,I195876,I294525,I195902,I195550,I195924,I195941,I195958,I195565,I195989,I196006,I294522,I195556,I196037,I195559,I195571,I195568,I196126,I467975,I196152,I196169,I196118,I196191,I196208,I467987,I196225,I467978,I196251,I196259,I467996,I196285,I196293,I467972,I196310,I196097,I467990,I196350,I196358,I196091,I196106,I196403,I467984,I467981,I196420,I467993,I196446,I196094,I196468,I196485,I196502,I196109,I196533,I196550,I196100,I196581,I196103,I196115,I196112,I196670,I196696,I196713,I196662,I196735,I196752,I196769,I196795,I196803,I196829,I196837,I196854,I196641,I196894,I196902,I196635,I196650,I196947,I196964,I196990,I196638,I197012,I197029,I197046,I196653,I197077,I197094,I196644,I197125,I196647,I196659,I196656,I197214,I531536,I197240,I197257,I197206,I197279,I197296,I531533,I531530,I197313,I531518,I197339,I197347,I531542,I197373,I197381,I531527,I197398,I197185,I531521,I197438,I197446,I197179,I197194,I197491,I531524,I197508,I531539,I197534,I197182,I197556,I197573,I197590,I197197,I197621,I197638,I197188,I197669,I197191,I197203,I197200,I197758,I350582,I197784,I197801,I197750,I197823,I197840,I350576,I350573,I197857,I350588,I197883,I197891,I197917,I197925,I350570,I197942,I197729,I197982,I197990,I197723,I197738,I198035,I350585,I350579,I198052,I198078,I197726,I198100,I198117,I198134,I197741,I198165,I198182,I350591,I197732,I198213,I197735,I197747,I197744,I198302,I322829,I198328,I198345,I198367,I198384,I322850,I322841,I198401,I198427,I198435,I322835,I198461,I198469,I322832,I198486,I322826,I198526,I198534,I198579,I322838,I198596,I322847,I198622,I198644,I198661,I198678,I198709,I198726,I322844,I198757,I198846,I198872,I198889,I198838,I198911,I198928,I198945,I198971,I198979,I199005,I199013,I199030,I198817,I199070,I199078,I198811,I198826,I199123,I199140,I199166,I198814,I199188,I199205,I199222,I198829,I199253,I199270,I198820,I199301,I198823,I198835,I198832,I199390,I199416,I199433,I199382,I199455,I199472,I199489,I199515,I199523,I199549,I199557,I199574,I199361,I199614,I199622,I199355,I199370,I199667,I199684,I199710,I199358,I199732,I199749,I199766,I199373,I199797,I199814,I199364,I199845,I199367,I199379,I199376,I199934,I199960,I199977,I199999,I200016,I200033,I200059,I200067,I200093,I200101,I200118,I200158,I200166,I200211,I200228,I200254,I200276,I200293,I200310,I200341,I200358,I200389,I200478,I443271,I200504,I200521,I200470,I200543,I200560,I443289,I200577,I443283,I200603,I200611,I443277,I200637,I200645,I443286,I200662,I200449,I443274,I200702,I200710,I200443,I200458,I200755,I443292,I200772,I200798,I200446,I200820,I200837,I200854,I200461,I200885,I200902,I443280,I200452,I200933,I200455,I200467,I200464,I201022,I415159,I201048,I201065,I201087,I201104,I415174,I415162,I201121,I415153,I201147,I201155,I415165,I201181,I201189,I415156,I201206,I415171,I201246,I201254,I201299,I415180,I415168,I201316,I415177,I201342,I201364,I201381,I201398,I201429,I201446,I201477,I201566,I263295,I201592,I201609,I201558,I201631,I201648,I263292,I263313,I201665,I263316,I201691,I201699,I263301,I201725,I201733,I263304,I201750,I201537,I263307,I201790,I201798,I201531,I201546,I201843,I263298,I201860,I263310,I201886,I201534,I201908,I201925,I201942,I201549,I201973,I201990,I201540,I202021,I201543,I201555,I201552,I202110,I202136,I202153,I202102,I202175,I202192,I202209,I202235,I202243,I202269,I202277,I202294,I202081,I202334,I202342,I202075,I202090,I202387,I202404,I202430,I202078,I202452,I202469,I202486,I202093,I202517,I202534,I202084,I202565,I202087,I202099,I202096,I202654,I202680,I202697,I202719,I202736,I202753,I202779,I202787,I202813,I202821,I202838,I202878,I202886,I202931,I202948,I202974,I202996,I203013,I203030,I203061,I203078,I203109,I203198,I260983,I203224,I203241,I203190,I203263,I203280,I260980,I261001,I203297,I261004,I203323,I203331,I260989,I203357,I203365,I260992,I203382,I203169,I260995,I203422,I203430,I203163,I203178,I203475,I260986,I203492,I260998,I203518,I203166,I203540,I203557,I203574,I203181,I203605,I203622,I203172,I203653,I203175,I203187,I203184,I203742,I464507,I203768,I203785,I203734,I203807,I203824,I464519,I203841,I464510,I203867,I203875,I464528,I203901,I203909,I464504,I203926,I203713,I464522,I203966,I203974,I203707,I203722,I204019,I464516,I464513,I204036,I464525,I204062,I203710,I204084,I204101,I204118,I203725,I204149,I204166,I203716,I204197,I203719,I203731,I203728,I204286,I204312,I204329,I204278,I204351,I204368,I204385,I204411,I204419,I204445,I204453,I204470,I204257,I204510,I204518,I204251,I204266,I204563,I204580,I204606,I204254,I204628,I204645,I204662,I204269,I204693,I204710,I204260,I204741,I204263,I204275,I204272,I204830,I495719,I204856,I204873,I204822,I204895,I204912,I495731,I204929,I495722,I204955,I204963,I495740,I204989,I204997,I495716,I205014,I204801,I495734,I205054,I205062,I204795,I204810,I205107,I495728,I495725,I205124,I495737,I205150,I204798,I205172,I205189,I205206,I204813,I205237,I205254,I204804,I205285,I204807,I204819,I204816,I205374,I444954,I205400,I205417,I205366,I205439,I205456,I444972,I205473,I444966,I205499,I205507,I444960,I205533,I205541,I444969,I205558,I205345,I444957,I205598,I205606,I205339,I205354,I205651,I444975,I205668,I205694,I205342,I205716,I205733,I205750,I205357,I205781,I205798,I444963,I205348,I205829,I205351,I205363,I205360,I205918,I432051,I205944,I205961,I205983,I206000,I432069,I206017,I432063,I206043,I206051,I432057,I206077,I206085,I432066,I206102,I432054,I206142,I206150,I206195,I432072,I206212,I206238,I206260,I206277,I206294,I206325,I206342,I432060,I206373,I206462,I216681,I206488,I206505,I206454,I206527,I206544,I216684,I216702,I206561,I216690,I206587,I206595,I206621,I206629,I216699,I206646,I206433,I216693,I206686,I206694,I206427,I206442,I206739,I216696,I216678,I206756,I216687,I206782,I206430,I206804,I206821,I206838,I206445,I206869,I206886,I206436,I206917,I206439,I206451,I206448,I207006,I207032,I207049,I207071,I207088,I207105,I207131,I207139,I207165,I207173,I207190,I207230,I207238,I207283,I207300,I207326,I207348,I207365,I207382,I207413,I207430,I207461,I207550,I207576,I207593,I207542,I207615,I207632,I207649,I207675,I207683,I207709,I207717,I207734,I207521,I207774,I207782,I207515,I207530,I207827,I207844,I207870,I207518,I207892,I207909,I207926,I207533,I207957,I207974,I207524,I208005,I207527,I207539,I207536,I208094,I262717,I208120,I208137,I208086,I208159,I208176,I262714,I262735,I208193,I262738,I208219,I208227,I262723,I208253,I208261,I262726,I208278,I208065,I262729,I208318,I208326,I208059,I208074,I208371,I262720,I208388,I262732,I208414,I208062,I208436,I208453,I208470,I208077,I208501,I208518,I208068,I208549,I208071,I208083,I208080,I208638,I248845,I208664,I208681,I208630,I208703,I208720,I248842,I248863,I208737,I248866,I208763,I208771,I248851,I208797,I208805,I248854,I208822,I208609,I248857,I208862,I208870,I208603,I208618,I208915,I248848,I208932,I248860,I208958,I208606,I208980,I208997,I209014,I208621,I209045,I209062,I208612,I209093,I208615,I208627,I208624,I209182,I511325,I209208,I209225,I209174,I209247,I209264,I511337,I511340,I209281,I511343,I209307,I209315,I511328,I209341,I209349,I511334,I209366,I209153,I511322,I209406,I209414,I209147,I209162,I209459,I511346,I209476,I511331,I209502,I209150,I209524,I209541,I209558,I209165,I209589,I209606,I209156,I209637,I209159,I209171,I209168,I209726,I354798,I209752,I209769,I209718,I209791,I209808,I354792,I354789,I209825,I354804,I209851,I209859,I209885,I209893,I354786,I209910,I209697,I209950,I209958,I209691,I209706,I210003,I354801,I354795,I210020,I210046,I209694,I210068,I210085,I210102,I209709,I210133,I210150,I354807,I209700,I210181,I209703,I209715,I209712,I210270,I387381,I210296,I210313,I210262,I210335,I210352,I387396,I387384,I210369,I387375,I210395,I210403,I387387,I210429,I210437,I387378,I210454,I210241,I387393,I210494,I210502,I210235,I210250,I210547,I387402,I387390,I210564,I387399,I210590,I210238,I210612,I210629,I210646,I210253,I210677,I210694,I210244,I210725,I210247,I210259,I210256,I210814,I210840,I210857,I210806,I210879,I210896,I210913,I210939,I210947,I210973,I210981,I210998,I210785,I211038,I211046,I210779,I210794,I211091,I211108,I211134,I210782,I211156,I211173,I211190,I210797,I211221,I211238,I210788,I211269,I210791,I210803,I210800,I211355,I317055,I211381,I211398,I211347,I317049,I211429,I211437,I317046,I211454,I211471,I317058,I211488,I317061,I211505,I211522,I211539,I211344,I211570,I317070,I211587,I317064,I211604,I211329,I211341,I211649,I211666,I211335,I211697,I317052,I211714,I211323,I211745,I317067,I211762,I211779,I211805,I211813,I211332,I211844,I211861,I211338,I211892,I211326,I211950,I211976,I211993,I211942,I212024,I212032,I212049,I212066,I212083,I212100,I212117,I212134,I211939,I212165,I212182,I212199,I211924,I211936,I212244,I212261,I211930,I212292,I212309,I211918,I212340,I212357,I212374,I212400,I212408,I211927,I212439,I212456,I211933,I212487,I211921,I212545,I247111,I212571,I212588,I247123,I212619,I212627,I247108,I212644,I212661,I247126,I212678,I247117,I212695,I212712,I212729,I212760,I247129,I212777,I247132,I212794,I212839,I212856,I212887,I212904,I212935,I247120,I212952,I247114,I212969,I212995,I213003,I213034,I213051,I213082,I213140,I213166,I213183,I213132,I213214,I213222,I213239,I213256,I213273,I213290,I213307,I213324,I213129,I213355,I213372,I213389,I213114,I213126,I213434,I213451,I213120,I213482,I213499,I213108,I213530,I213547,I213564,I213590,I213598,I213117,I213629,I213646,I213123,I213677,I213111,I213735,I376408,I213761,I213778,I376396,I213809,I213817,I376393,I213834,I213851,I376405,I213868,I376402,I213885,I213902,I213919,I213950,I376411,I213967,I376414,I213984,I214029,I214046,I214077,I376417,I214094,I214125,I376420,I214142,I376399,I214159,I214185,I214193,I214224,I214241,I214272,I214330,I214356,I214373,I214404,I214412,I214429,I214446,I214463,I214480,I214497,I214514,I214545,I214562,I214579,I214624,I214641,I214672,I214689,I214720,I214737,I214754,I214780,I214788,I214819,I214836,I214867,I214925,I393850,I214951,I214968,I393838,I214999,I215007,I393835,I215024,I215041,I393847,I215058,I393844,I215075,I215092,I215109,I215140,I393853,I215157,I393856,I215174,I215219,I215236,I215267,I393859,I215284,I215315,I393862,I215332,I393841,I215349,I215375,I215383,I215414,I215431,I215462,I215520,I215546,I215563,I215594,I215602,I215619,I215636,I215653,I215670,I215687,I215704,I215735,I215752,I215769,I215814,I215831,I215862,I215879,I215910,I215927,I215944,I215970,I215978,I216009,I216026,I216057,I216115,I216141,I216158,I216107,I216189,I216197,I216214,I216231,I216248,I216265,I216282,I216299,I216104,I216330,I216347,I216364,I216089,I216101,I216409,I216426,I216095,I216457,I216474,I216083,I216505,I216522,I216539,I216565,I216573,I216092,I216604,I216621,I216098,I216652,I216086,I216710,I526325,I216736,I216753,I526331,I216784,I216792,I526319,I216809,I216826,I526322,I216843,I526328,I216860,I216877,I216894,I216925,I216942,I526337,I216959,I217004,I217021,I217052,I526316,I217069,I217100,I526340,I217117,I217134,I526334,I217160,I217168,I217199,I217216,I217247,I217305,I291623,I217331,I217348,I217297,I291617,I217379,I217387,I291614,I217404,I217421,I291626,I217438,I291629,I217455,I217472,I217489,I217294,I217520,I291638,I217537,I291632,I217554,I217279,I217291,I217599,I217616,I217285,I217647,I291620,I217664,I217273,I217695,I291635,I217712,I217729,I217755,I217763,I217282,I217794,I217811,I217288,I217842,I217276,I217900,I236129,I217926,I217943,I217892,I236141,I217974,I217982,I236126,I217999,I218016,I236144,I218033,I236135,I218050,I218067,I218084,I217889,I218115,I236147,I218132,I236150,I218149,I217874,I217886,I218194,I218211,I217880,I218242,I218259,I217868,I218290,I236138,I218307,I236132,I218324,I218350,I218358,I217877,I218389,I218406,I217883,I218437,I217871,I218495,I218521,I218538,I218487,I218569,I218577,I218594,I218611,I218628,I218645,I218662,I218679,I218484,I218710,I218727,I218744,I218469,I218481,I218789,I218806,I218475,I218837,I218854,I218463,I218885,I218902,I218919,I218945,I218953,I218472,I218984,I219001,I218478,I219032,I218466,I219090,I501514,I219116,I219133,I501496,I219164,I219172,I501502,I219189,I219206,I501517,I219223,I501508,I219240,I219257,I219274,I219305,I501520,I219322,I501499,I219339,I219384,I219401,I219432,I501505,I219449,I219480,I501511,I219497,I219514,I219540,I219548,I219579,I219596,I219627,I219685,I219711,I219728,I219677,I219759,I219767,I219784,I219801,I219818,I219835,I219852,I219869,I219674,I219900,I219917,I219934,I219659,I219671,I219979,I219996,I219665,I220027,I220044,I219653,I220075,I220092,I220109,I220135,I220143,I219662,I220174,I220191,I219668,I220222,I219656,I220280,I304917,I220306,I220323,I304911,I220354,I220362,I304908,I220379,I220396,I304920,I220413,I304923,I220430,I220447,I220464,I220495,I304932,I220512,I304926,I220529,I220574,I220591,I220622,I304914,I220639,I220670,I304929,I220687,I220704,I220730,I220738,I220769,I220786,I220817,I220875,I347417,I220901,I220918,I220867,I347414,I220949,I220957,I220974,I220991,I347411,I221008,I347426,I221025,I221042,I221059,I220864,I221090,I347420,I221107,I347408,I221124,I220849,I220861,I221169,I221186,I220855,I221217,I347429,I221234,I220843,I221265,I221282,I347423,I221299,I221325,I221333,I220852,I221364,I221381,I220858,I221412,I220846,I221470,I221496,I221513,I221462,I221544,I221552,I221569,I221586,I221603,I221620,I221637,I221654,I221459,I221685,I221702,I221719,I221444,I221456,I221764,I221781,I221450,I221812,I221829,I221438,I221860,I221877,I221894,I221920,I221928,I221447,I221959,I221976,I221453,I222007,I221441,I222065,I235551,I222091,I222108,I235563,I222139,I222147,I235548,I222164,I222181,I235566,I222198,I235557,I222215,I222232,I222249,I222280,I235569,I222297,I235572,I222314,I222359,I222376,I222407,I222424,I222455,I235560,I222472,I235554,I222489,I222515,I222523,I222554,I222571,I222602,I222660,I222686,I222703,I222652,I222734,I222742,I222759,I222776,I222793,I222810,I222827,I222844,I222649,I222875,I222892,I222909,I222634,I222646,I222954,I222971,I222640,I223002,I223019,I222628,I223050,I223067,I223084,I223110,I223118,I222637,I223149,I223166,I222643,I223197,I222631,I223255,I255781,I223281,I223298,I223247,I255793,I223329,I223337,I255778,I223354,I223371,I255796,I223388,I255787,I223405,I223422,I223439,I223244,I223470,I255799,I223487,I255802,I223504,I223229,I223241,I223549,I223566,I223235,I223597,I223614,I223223,I223645,I255790,I223662,I255784,I223679,I223705,I223713,I223232,I223744,I223761,I223238,I223792,I223226,I223850,I446076,I223876,I223893,I223842,I446079,I223924,I223932,I446082,I223949,I223966,I446094,I223983,I446085,I224000,I224017,I224034,I223839,I224065,I446091,I224082,I224099,I223824,I223836,I224144,I224161,I223830,I224192,I224209,I223818,I224240,I446088,I224257,I224274,I446097,I224300,I224308,I223827,I224339,I224356,I223833,I224387,I223821,I224445,I367970,I224471,I224488,I367967,I224519,I224527,I224544,I224561,I367964,I224578,I367979,I224595,I224612,I224629,I224660,I367973,I224677,I367961,I224694,I224739,I224756,I224787,I367982,I224804,I224835,I224852,I367976,I224869,I224895,I224903,I224934,I224951,I224982,I225040,I292779,I225066,I225083,I225032,I292773,I225114,I225122,I292770,I225139,I225156,I292782,I225173,I292785,I225190,I225207,I225224,I225029,I225255,I292794,I225272,I292788,I225289,I225014,I225026,I225334,I225351,I225020,I225382,I292776,I225399,I225008,I225430,I292791,I225447,I225464,I225490,I225498,I225017,I225529,I225546,I225023,I225577,I225011,I225635,I437661,I225661,I225678,I437664,I225709,I225717,I437667,I225734,I225751,I437679,I225768,I437670,I225785,I225802,I225819,I225850,I437676,I225867,I225884,I225929,I225946,I225977,I225994,I226025,I437673,I226042,I226059,I437682,I226085,I226093,I226124,I226141,I226172,I226230,I375348,I226256,I226273,I375345,I226304,I226312,I226329,I226346,I375342,I226363,I375357,I226380,I226397,I226414,I226445,I375351,I226462,I375339,I226479,I226524,I226541,I226572,I375360,I226589,I226620,I226637,I375354,I226654,I226680,I226688,I226719,I226736,I226767,I226825,I538384,I226851,I226868,I226817,I538390,I226899,I226907,I538393,I226924,I226941,I538396,I226958,I538381,I226975,I226992,I227009,I226814,I227040,I538387,I227057,I538369,I227074,I226799,I226811,I227119,I227136,I226805,I227167,I227184,I226793,I227215,I538378,I227232,I538375,I227249,I538372,I227275,I227283,I226802,I227314,I227331,I226808,I227362,I226796,I227420,I227446,I227463,I227412,I227494,I227502,I227519,I227536,I227553,I227570,I227587,I227604,I227409,I227635,I227652,I227669,I227394,I227406,I227714,I227731,I227400,I227762,I227779,I227388,I227810,I227827,I227844,I227870,I227878,I227397,I227909,I227926,I227403,I227957,I227391,I228015,I228041,I228058,I228007,I228089,I228097,I228114,I228131,I228148,I228165,I228182,I228199,I228004,I228230,I228247,I228264,I227989,I228001,I228309,I228326,I227995,I228357,I228374,I227983,I228405,I228422,I228439,I228465,I228473,I227992,I228504,I228521,I227998,I228552,I227986,I228610,I228636,I228653,I228602,I228684,I228692,I228709,I228726,I228743,I228760,I228777,I228794,I228599,I228825,I228842,I228859,I228584,I228596,I228904,I228921,I228590,I228952,I228969,I228578,I229000,I229017,I229034,I229060,I229068,I228587,I229099,I229116,I228593,I229147,I228581,I229205,I458742,I229231,I229248,I458724,I229279,I229287,I458730,I229304,I229321,I458745,I229338,I458736,I229355,I229372,I229389,I229420,I458748,I229437,I458727,I229454,I229499,I229516,I229547,I458733,I229564,I229595,I458739,I229612,I229629,I229655,I229663,I229694,I229711,I229742,I229800,I463348,I229826,I229834,I463354,I229860,I229868,I229885,I463351,I229902,I229919,I463369,I229936,I229967,I229984,I230001,I463372,I230018,I230063,I230108,I463357,I230125,I230142,I230173,I463363,I230190,I463360,I230207,I463366,I230233,I230241,I230286,I230303,I230320,I230378,I230404,I230412,I230438,I230446,I230463,I230480,I230497,I230514,I230545,I230562,I230579,I230596,I230641,I230686,I230703,I230720,I230751,I230768,I230785,I230811,I230819,I230864,I230881,I230898,I230956,I423557,I230982,I230990,I423554,I231016,I231024,I423551,I231041,I423578,I231058,I231075,I423566,I231092,I231123,I231140,I231157,I423572,I231174,I423563,I231219,I231264,I423560,I231281,I231298,I231329,I423575,I231346,I423569,I231363,I231389,I231397,I231442,I231459,I231476,I231534,I231560,I231568,I231594,I231602,I231619,I231636,I231653,I231670,I231520,I231701,I231718,I231735,I231752,I231517,I231508,I231797,I231511,I231505,I231842,I231859,I231876,I231514,I231907,I231924,I231941,I231967,I231975,I231502,I231526,I232020,I232037,I232054,I231523,I232112,I232138,I232146,I232172,I232180,I232197,I232214,I232231,I232248,I232098,I232279,I232296,I232313,I232330,I232095,I232086,I232375,I232089,I232083,I232420,I232437,I232454,I232092,I232485,I232502,I232519,I232545,I232553,I232080,I232104,I232598,I232615,I232632,I232101,I232690,I232716,I232724,I232750,I232758,I232775,I232792,I232809,I232826,I232676,I232857,I232874,I232891,I232908,I232673,I232664,I232953,I232667,I232661,I232998,I233015,I233032,I232670,I233063,I233080,I233097,I233123,I233131,I232658,I232682,I233176,I233193,I233210,I232679,I233268,I391257,I233294,I233302,I391254,I233328,I233336,I391251,I233353,I391278,I233370,I233387,I391266,I233404,I233254,I233435,I233452,I233469,I391272,I233486,I391263,I233251,I233242,I233531,I233245,I233239,I233576,I391260,I233593,I233610,I233248,I233641,I391275,I233658,I391269,I233675,I233701,I233709,I233236,I233260,I233754,I233771,I233788,I233257,I233846,I436560,I233872,I233880,I436551,I233906,I233914,I436545,I233931,I436557,I233948,I233965,I436548,I233982,I234013,I234030,I234047,I436554,I234064,I436539,I234109,I234154,I234171,I234188,I234219,I436542,I234236,I234253,I234279,I234287,I234332,I234349,I234366,I234424,I442170,I234450,I234458,I442161,I234484,I234492,I442155,I234509,I442167,I234526,I234543,I442158,I234560,I234410,I234591,I234608,I234625,I442164,I234642,I442149,I234407,I234398,I234687,I234401,I234395,I234732,I234749,I234766,I234404,I234797,I442152,I234814,I234831,I234857,I234865,I234392,I234416,I234910,I234927,I234944,I234413,I235002,I235028,I235036,I235062,I235070,I235087,I235104,I235121,I235138,I234988,I235169,I235186,I235203,I235220,I234985,I234976,I235265,I234979,I234973,I235310,I235327,I235344,I234982,I235375,I235392,I235409,I235435,I235443,I234970,I234994,I235488,I235505,I235522,I234991,I235580,I235606,I235614,I235640,I235648,I235665,I235682,I235699,I235716,I235747,I235764,I235781,I235798,I235843,I235888,I235905,I235922,I235953,I235970,I235987,I236013,I236021,I236066,I236083,I236100,I236158,I236184,I236192,I236218,I236226,I236243,I236260,I236277,I236294,I236325,I236342,I236359,I236376,I236421,I236466,I236483,I236500,I236531,I236548,I236565,I236591,I236599,I236644,I236661,I236678,I236736,I236762,I236770,I236796,I236804,I236821,I236838,I236855,I236872,I236903,I236920,I236937,I236954,I236999,I237044,I237061,I237078,I237109,I237126,I237143,I237169,I237177,I237222,I237239,I237256,I237314,I237340,I237348,I237374,I237382,I237399,I237416,I237433,I237450,I237481,I237498,I237515,I237532,I237577,I237622,I237639,I237656,I237687,I237704,I237721,I237747,I237755,I237800,I237817,I237834,I237892,I435438,I237918,I237926,I435429,I237952,I237960,I435423,I237977,I435435,I237994,I238011,I435426,I238028,I237878,I238059,I238076,I238093,I435432,I238110,I435417,I237875,I237866,I238155,I237869,I237863,I238200,I238217,I238234,I237872,I238265,I435420,I238282,I238299,I238325,I238333,I237860,I237884,I238378,I238395,I238412,I237881,I238470,I238496,I238504,I238530,I238538,I238555,I238572,I238589,I238606,I238456,I238637,I238654,I238671,I238688,I238453,I238444,I238733,I238447,I238441,I238778,I238795,I238812,I238450,I238843,I238860,I238877,I238903,I238911,I238438,I238462,I238956,I238973,I238990,I238459,I239048,I239074,I239082,I239108,I239116,I239133,I239150,I239167,I239184,I239215,I239232,I239249,I239266,I239311,I239356,I239373,I239390,I239421,I239438,I239455,I239481,I239489,I239534,I239551,I239568,I239626,I271384,I239652,I239660,I271396,I239686,I239694,I271387,I239711,I271390,I239728,I239745,I271393,I239762,I239612,I239793,I239810,I239827,I239844,I271399,I239609,I239600,I239889,I239603,I239597,I239934,I271405,I239951,I239968,I239606,I239999,I240016,I271402,I240033,I271408,I240059,I240067,I239594,I239618,I240112,I240129,I240146,I239615,I240204,I478954,I240230,I240238,I478960,I240264,I240272,I240289,I478957,I240306,I240323,I478975,I240340,I240371,I240388,I240405,I478978,I240422,I240467,I240512,I478963,I240529,I240546,I240577,I478969,I240594,I478966,I240611,I478972,I240637,I240645,I240690,I240707,I240724,I240782,I240808,I240816,I240842,I240850,I240867,I240884,I240901,I240918,I240949,I240966,I240983,I241000,I241045,I241090,I241107,I241124,I241155,I241172,I241189,I241215,I241223,I241268,I241285,I241302,I241360,I506444,I241386,I241394,I506438,I241420,I241428,I506447,I241445,I506426,I241462,I241479,I506435,I241496,I241346,I241527,I241544,I241561,I506450,I241578,I506429,I241343,I241334,I241623,I241337,I241331,I241668,I506432,I241685,I241702,I241340,I241733,I506441,I241750,I241767,I241793,I241801,I241328,I241352,I241846,I241863,I241880,I241349,I241938,I241964,I241972,I241998,I242006,I242023,I242040,I242057,I242074,I242105,I242122,I242139,I242156,I242201,I242246,I242263,I242280,I242311,I242328,I242345,I242371,I242379,I242424,I242441,I242458,I242516,I242542,I242550,I242576,I242584,I242601,I242618,I242635,I242652,I242683,I242700,I242717,I242734,I242779,I242824,I242841,I242858,I242889,I242906,I242923,I242949,I242957,I243002,I243019,I243036,I243094,I243120,I243128,I243154,I243162,I243179,I243196,I243213,I243230,I243080,I243261,I243278,I243295,I243312,I243077,I243068,I243357,I243071,I243065,I243402,I243419,I243436,I243074,I243467,I243484,I243501,I243527,I243535,I243062,I243086,I243580,I243597,I243614,I243083,I243672,I378337,I243698,I243706,I378334,I243732,I243740,I378331,I243757,I378358,I243774,I243791,I378346,I243808,I243839,I243856,I243873,I378352,I243890,I378343,I243935,I243980,I378340,I243997,I244014,I244045,I378355,I244062,I378349,I244079,I244105,I244113,I244158,I244175,I244192,I244250,I359535,I244276,I244284,I244310,I244318,I359532,I244335,I359547,I244352,I244369,I359541,I244386,I244236,I244417,I244434,I244451,I359538,I244468,I359529,I244233,I244224,I244513,I244227,I244221,I244558,I359550,I244575,I244592,I244230,I244623,I244640,I244657,I359544,I244683,I244691,I244218,I244242,I244736,I244753,I244770,I244239,I244828,I435999,I244854,I244862,I435990,I244888,I244896,I435984,I244913,I435996,I244930,I244947,I435987,I244964,I244995,I245012,I245029,I435993,I245046,I435978,I245091,I245136,I245153,I245170,I245201,I435981,I245218,I245235,I245261,I245269,I245314,I245331,I245348,I245406,I530374,I245432,I245440,I530386,I245466,I245474,I530377,I245491,I530365,I245508,I245525,I530362,I245542,I245573,I245590,I245607,I530368,I245624,I245669,I245714,I530383,I245731,I245748,I245779,I530371,I245796,I245813,I530380,I245839,I245847,I245892,I245909,I245926,I245984,I548450,I246010,I246018,I246044,I246052,I548474,I246069,I548456,I246086,I246103,I548471,I246120,I245970,I246151,I246168,I246185,I548453,I246202,I548462,I245967,I245958,I246247,I245961,I245955,I246292,I548459,I246309,I246326,I245964,I246357,I548468,I246374,I548477,I246391,I548465,I246417,I246425,I245952,I245976,I246470,I246487,I246504,I245973,I246562,I332658,I246588,I246596,I246622,I246630,I332655,I246647,I332670,I246664,I246681,I332664,I246698,I246548,I246729,I246746,I246763,I332661,I246780,I332652,I246545,I246536,I246825,I246539,I246533,I246870,I332673,I246887,I246904,I246542,I246935,I246952,I246969,I332667,I246995,I247003,I246530,I246554,I247048,I247065,I247082,I246551,I247140,I310688,I247166,I247174,I310700,I247200,I247208,I310691,I247225,I310694,I247242,I247259,I310697,I247276,I247307,I247324,I247341,I247358,I310703,I247403,I247448,I310709,I247465,I247482,I247513,I247530,I310706,I247547,I310712,I247573,I247581,I247626,I247643,I247660,I247718,I285834,I247744,I247752,I285846,I247778,I247786,I285837,I247803,I285840,I247820,I247837,I285843,I247854,I247885,I247902,I247919,I247936,I285849,I247981,I248026,I285855,I248043,I248060,I248091,I248108,I285852,I248125,I285858,I248151,I248159,I248204,I248221,I248238,I248296,I564515,I248322,I248330,I248356,I248364,I564539,I248381,I564521,I248398,I248415,I564536,I248432,I248282,I248463,I248480,I248497,I564518,I248514,I564527,I248279,I248270,I248559,I248273,I248267,I248604,I564524,I248621,I248638,I248276,I248669,I564533,I248686,I564542,I248703,I564530,I248729,I248737,I248264,I248288,I248782,I248799,I248816,I248285,I248874,I419035,I248900,I248908,I419032,I248934,I248942,I419029,I248959,I419056,I248976,I248993,I419044,I249010,I249041,I249058,I249075,I419050,I249092,I419041,I249137,I249182,I419038,I249199,I249216,I249247,I419053,I249264,I419047,I249281,I249307,I249315,I249360,I249377,I249394,I249452,I342144,I249478,I249486,I249512,I249520,I342141,I249537,I342156,I249554,I249571,I342150,I249588,I249619,I249636,I249653,I342147,I249670,I342138,I249715,I249760,I342159,I249777,I249794,I249825,I249842,I249859,I342153,I249885,I249893,I249938,I249955,I249972,I250030,I250056,I250064,I250090,I250098,I250115,I250132,I250149,I250166,I250016,I250197,I250214,I250231,I250248,I250013,I250004,I250293,I250007,I250001,I250338,I250355,I250372,I250010,I250403,I250420,I250437,I250463,I250471,I249998,I250022,I250516,I250533,I250550,I250019,I250608,I250634,I250642,I250668,I250676,I250693,I250710,I250727,I250744,I250775,I250792,I250809,I250826,I250871,I250916,I250933,I250950,I250981,I250998,I251015,I251041,I251049,I251094,I251111,I251128,I251186,I355319,I251212,I251220,I251246,I251254,I355316,I251271,I355331,I251288,I251305,I355325,I251322,I251353,I251370,I251387,I355322,I251404,I355313,I251449,I251494,I355334,I251511,I251528,I251559,I251576,I251593,I355328,I251619,I251627,I251672,I251689,I251706,I251764,I251790,I251798,I251824,I251832,I251849,I251866,I251883,I251900,I251750,I251931,I251948,I251965,I251982,I251747,I251738,I252027,I251741,I251735,I252072,I252089,I252106,I251744,I252137,I252154,I252171,I252197,I252205,I251732,I251756,I252250,I252267,I252284,I251753,I252342,I252368,I252376,I252402,I252410,I252427,I252444,I252461,I252478,I252509,I252526,I252543,I252560,I252605,I252650,I252667,I252684,I252715,I252732,I252749,I252775,I252783,I252828,I252845,I252862,I252920,I252946,I252954,I252980,I252988,I253005,I253022,I253039,I253056,I253087,I253104,I253121,I253138,I253183,I253228,I253245,I253262,I253293,I253310,I253327,I253353,I253361,I253406,I253423,I253440,I253498,I293348,I253524,I253532,I293360,I253558,I253566,I293351,I253583,I293354,I253600,I253617,I293357,I253634,I253484,I253665,I253682,I253699,I253716,I293363,I253481,I253472,I253761,I253475,I253469,I253806,I293369,I253823,I253840,I253478,I253871,I253888,I293366,I253905,I293372,I253931,I253939,I253466,I253490,I253984,I254001,I254018,I253487,I254076,I420327,I254102,I254110,I420324,I254136,I254144,I420321,I254161,I420348,I254178,I254195,I420336,I254212,I254062,I254243,I254260,I254277,I420342,I254294,I420333,I254059,I254050,I254339,I254053,I254047,I254384,I420330,I254401,I254418,I254056,I254449,I420345,I254466,I420339,I254483,I254509,I254517,I254044,I254068,I254562,I254579,I254596,I254065,I254654,I455834,I254680,I254688,I455840,I254714,I254722,I254739,I455837,I254756,I254773,I455855,I254790,I254640,I254821,I254838,I254855,I455858,I254872,I254637,I254628,I254917,I254631,I254625,I254962,I455843,I254979,I254996,I254634,I255027,I455849,I255044,I455846,I255061,I455852,I255087,I255095,I254622,I254646,I255140,I255157,I255174,I254643,I255232,I255258,I255266,I255292,I255300,I255317,I255334,I255351,I255368,I255218,I255399,I255416,I255433,I255450,I255215,I255206,I255495,I255209,I255203,I255540,I255557,I255574,I255212,I255605,I255622,I255639,I255665,I255673,I255200,I255224,I255718,I255735,I255752,I255221,I255810,I255836,I255844,I255870,I255878,I255895,I255912,I255929,I255946,I255977,I255994,I256011,I256028,I256073,I256118,I256135,I256152,I256183,I256200,I256217,I256243,I256251,I256296,I256313,I256330,I256388,I354265,I256414,I256422,I256448,I256456,I354262,I256473,I354277,I256490,I256507,I354271,I256524,I256374,I256555,I256572,I256589,I354268,I256606,I354259,I256371,I256362,I256651,I256365,I256359,I256696,I354280,I256713,I256730,I256368,I256761,I256778,I256795,I354274,I256821,I256829,I256356,I256380,I256874,I256891,I256908,I256377,I256966,I256992,I257000,I257026,I257034,I257051,I257068,I257085,I257102,I257133,I257150,I257167,I257184,I257229,I257274,I257291,I257308,I257339,I257356,I257373,I257399,I257407,I257452,I257469,I257486,I257544,I325138,I257570,I257578,I325150,I257604,I257612,I325141,I257629,I325144,I257646,I257663,I325147,I257680,I257530,I257711,I257728,I257745,I257762,I325153,I257527,I257518,I257807,I257521,I257515,I257852,I325159,I257869,I257886,I257524,I257917,I257934,I325156,I257951,I325162,I257977,I257985,I257512,I257536,I258030,I258047,I258064,I257533,I258122,I258148,I258156,I258182,I258190,I258207,I258224,I258241,I258258,I258289,I258306,I258323,I258340,I258385,I258430,I258447,I258464,I258495,I258512,I258529,I258555,I258563,I258608,I258625,I258642,I258700,I307798,I258726,I258734,I307810,I258760,I258768,I307801,I258785,I307804,I258802,I258819,I307807,I258836,I258686,I258867,I258884,I258901,I258918,I307813,I258683,I258674,I258963,I258677,I258671,I259008,I307819,I259025,I259042,I258680,I259073,I259090,I307816,I259107,I307822,I259133,I259141,I258668,I258692,I259186,I259203,I259220,I258689,I259278,I374818,I259304,I259312,I259338,I259346,I374815,I259363,I374830,I259380,I259397,I374824,I259414,I259264,I259445,I259462,I259479,I374821,I259496,I374812,I259261,I259252,I259541,I259255,I259249,I259586,I374833,I259603,I259620,I259258,I259651,I259668,I259685,I374827,I259711,I259719,I259246,I259270,I259764,I259781,I259798,I259267,I259856,I259882,I259890,I259916,I259924,I259941,I259958,I259975,I259992,I259842,I260023,I260040,I260057,I260074,I259839,I259830,I260119,I259833,I259827,I260164,I260181,I260198,I259836,I260229,I260246,I260263,I260289,I260297,I259824,I259848,I260342,I260359,I260376,I259845,I260434,I260460,I260468,I260494,I260502,I260519,I260536,I260553,I260570,I260601,I260618,I260635,I260652,I260697,I260742,I260759,I260776,I260807,I260824,I260841,I260867,I260875,I260920,I260937,I260954,I261012,I543095,I261038,I261046,I261072,I261080,I543119,I261097,I543101,I261114,I261131,I543116,I261148,I261179,I261196,I261213,I543098,I261230,I543107,I261275,I261320,I543104,I261337,I261354,I261385,I543113,I261402,I543122,I261419,I543110,I261445,I261453,I261498,I261515,I261532,I261590,I261616,I261624,I261650,I261658,I261675,I261692,I261709,I261726,I261757,I261774,I261791,I261808,I261853,I261898,I261915,I261932,I261963,I261980,I261997,I262023,I262031,I262076,I262093,I262110,I262168,I556185,I262194,I262202,I262228,I262236,I556209,I262253,I556191,I262270,I262287,I556206,I262304,I262154,I262335,I262352,I262369,I556188,I262386,I556197,I262151,I262142,I262431,I262145,I262139,I262476,I556194,I262493,I262510,I262148,I262541,I556203,I262558,I556212,I262575,I556200,I262601,I262609,I262136,I262160,I262654,I262671,I262688,I262157,I262746,I262772,I262780,I262806,I262814,I262831,I262848,I262865,I262882,I262913,I262930,I262947,I262964,I263009,I263054,I263071,I263088,I263119,I263136,I263153,I263179,I263187,I263232,I263249,I263266,I263324,I499762,I263350,I263358,I499768,I263384,I263392,I263409,I499765,I263426,I263443,I499783,I263460,I263491,I263508,I263525,I499786,I263542,I263587,I263632,I499771,I263649,I263666,I263697,I499777,I263714,I499774,I263731,I499780,I263757,I263765,I263810,I263827,I263844,I263902,I315890,I263928,I263936,I315902,I263962,I263970,I315893,I263987,I315896,I264004,I264021,I315899,I264038,I264069,I264086,I264103,I264120,I315905,I264165,I264210,I315911,I264227,I264244,I264275,I264292,I315908,I264309,I315914,I264335,I264343,I264388,I264405,I264422,I264480,I353738,I264506,I264514,I264540,I264548,I353735,I264565,I353750,I264582,I264599,I353744,I264616,I264466,I264647,I264664,I264681,I353741,I264698,I353732,I264463,I264454,I264743,I264457,I264451,I264788,I353753,I264805,I264822,I264460,I264853,I264870,I264887,I353747,I264913,I264921,I264448,I264472,I264966,I264983,I265000,I264469,I265058,I265084,I265092,I265109,I265126,I265152,I265160,I265186,I265194,I265211,I265228,I265245,I265285,I265293,I265310,I265327,I265344,I265375,I265392,I265418,I265426,I265457,I265488,I265505,I265536,I265636,I459320,I265662,I265670,I265687,I459302,I459314,I265704,I459317,I265730,I265738,I459311,I459308,I265764,I265772,I265789,I265806,I265823,I459326,I265863,I265871,I265888,I265905,I265922,I265953,I459305,I265970,I265996,I266004,I266035,I266066,I266083,I266114,I459323,I266214,I266240,I266248,I266265,I266282,I266308,I266316,I266342,I266350,I266367,I266384,I266401,I266197,I266441,I266449,I266466,I266483,I266500,I266200,I266531,I266548,I266574,I266582,I266182,I266613,I266191,I266644,I266661,I266203,I266692,I266194,I266185,I266188,I266206,I266792,I266818,I266826,I266843,I266860,I266886,I266894,I266920,I266928,I266945,I266962,I266979,I266775,I267019,I267027,I267044,I267061,I267078,I266778,I267109,I267126,I267152,I267160,I266760,I267191,I266769,I267222,I267239,I266781,I267270,I266772,I266763,I266766,I266784,I267370,I267396,I267404,I267421,I267438,I267464,I267472,I267498,I267506,I267523,I267540,I267557,I267353,I267597,I267605,I267622,I267639,I267656,I267356,I267687,I267704,I267730,I267738,I267338,I267769,I267347,I267800,I267817,I267359,I267848,I267350,I267341,I267344,I267362,I267948,I544907,I267974,I267982,I267999,I544892,I544880,I268016,I544895,I268042,I268050,I544898,I268076,I268084,I268101,I268118,I268135,I267931,I544886,I268175,I268183,I268200,I268217,I268234,I267934,I268265,I544883,I544889,I268282,I544904,I268308,I268316,I267916,I268347,I267925,I268378,I268395,I267937,I268426,I544901,I267928,I267919,I267922,I267940,I268526,I268552,I268560,I268577,I268594,I268620,I268628,I268654,I268662,I268679,I268696,I268713,I268509,I268753,I268761,I268778,I268795,I268812,I268512,I268843,I268860,I268886,I268894,I268494,I268925,I268503,I268956,I268973,I268515,I269004,I268506,I268497,I268500,I268518,I269104,I269130,I269138,I269155,I269172,I269198,I269206,I269232,I269240,I269257,I269274,I269291,I269331,I269339,I269356,I269373,I269390,I269421,I269438,I269464,I269472,I269503,I269534,I269551,I269582,I269682,I269708,I269716,I269733,I269750,I269776,I269784,I269810,I269818,I269835,I269852,I269869,I269909,I269917,I269934,I269951,I269968,I269999,I270016,I270042,I270050,I270081,I270112,I270129,I270160,I270260,I529206,I270286,I270294,I270311,I529230,I529212,I270328,I529218,I270354,I270362,I529224,I529209,I270388,I270396,I270413,I270430,I270447,I270243,I529221,I270487,I270495,I270512,I270529,I270546,I270246,I270577,I529227,I529215,I270594,I270620,I270628,I270228,I270659,I270237,I270690,I270707,I270249,I270738,I270240,I270231,I270234,I270252,I270838,I511866,I270864,I270872,I270889,I511869,I511878,I270906,I511881,I270932,I270940,I511890,I511872,I270966,I270974,I270991,I271008,I271025,I270821,I271065,I271073,I271090,I271107,I271124,I270824,I271155,I511887,I271172,I511884,I271198,I271206,I270806,I271237,I270815,I271268,I271285,I270827,I271316,I511875,I270818,I270809,I270812,I270830,I271416,I470302,I271442,I271450,I271467,I470284,I470296,I271484,I470299,I271510,I271518,I470293,I470290,I271544,I271552,I271569,I271586,I271603,I470308,I271643,I271651,I271668,I271685,I271702,I271733,I470287,I271750,I271776,I271784,I271815,I271846,I271863,I271894,I470305,I271994,I272020,I272028,I272045,I272062,I272088,I272096,I272122,I272130,I272147,I272164,I272181,I272221,I272229,I272246,I272263,I272280,I272311,I272328,I272354,I272362,I272393,I272424,I272441,I272472,I272572,I272598,I272606,I272623,I272640,I272666,I272674,I272700,I272708,I272725,I272742,I272759,I272555,I272799,I272807,I272824,I272841,I272858,I272558,I272889,I272906,I272932,I272940,I272540,I272971,I272549,I273002,I273019,I272561,I273050,I272552,I272543,I272546,I272564,I273150,I481284,I273176,I273184,I273201,I481266,I481278,I273218,I481281,I273244,I273252,I481275,I481272,I273278,I273286,I273303,I273320,I273337,I273133,I481290,I273377,I273385,I273402,I273419,I273436,I273136,I273467,I481269,I273484,I273510,I273518,I273118,I273549,I273127,I273580,I273597,I273139,I273628,I481287,I273130,I273121,I273124,I273142,I273728,I273754,I273762,I273779,I273796,I273822,I273830,I273856,I273864,I273881,I273898,I273915,I273711,I273955,I273963,I273980,I273997,I274014,I273714,I274045,I274062,I274088,I274096,I273696,I274127,I273705,I274158,I274175,I273717,I274206,I273708,I273699,I273702,I273720,I274306,I427008,I274332,I274340,I274357,I427005,I427023,I274374,I427020,I274400,I274408,I427002,I274434,I274442,I274459,I274476,I274493,I274289,I427014,I274533,I274541,I274558,I274575,I274592,I274292,I274623,I427017,I274640,I274666,I274674,I274274,I274705,I274283,I274736,I274753,I274295,I274784,I427011,I274286,I274277,I274280,I274298,I274884,I274910,I274918,I274935,I274952,I274978,I274986,I275012,I275020,I275037,I275054,I275071,I275111,I275119,I275136,I275153,I275170,I275201,I275218,I275244,I275252,I275283,I275314,I275331,I275362,I275462,I275488,I275496,I275513,I275530,I275556,I275564,I275590,I275598,I275615,I275632,I275649,I275445,I275689,I275697,I275714,I275731,I275748,I275448,I275779,I275796,I275822,I275830,I275430,I275861,I275439,I275892,I275909,I275451,I275940,I275442,I275433,I275436,I275454,I276040,I276066,I276074,I276091,I276108,I276134,I276142,I276168,I276176,I276193,I276210,I276227,I276023,I276267,I276275,I276292,I276309,I276326,I276026,I276357,I276374,I276400,I276408,I276008,I276439,I276017,I276470,I276487,I276029,I276518,I276020,I276011,I276014,I276032,I276618,I276644,I276652,I276669,I276686,I276712,I276720,I276746,I276754,I276771,I276788,I276805,I276601,I276845,I276853,I276870,I276887,I276904,I276604,I276935,I276952,I276978,I276986,I276586,I277017,I276595,I277048,I277065,I276607,I277096,I276598,I276589,I276592,I276610,I277196,I522270,I277222,I277230,I277247,I522294,I522276,I277264,I522282,I277290,I277298,I522288,I522273,I277324,I277332,I277349,I277366,I277383,I277179,I522285,I277423,I277431,I277448,I277465,I277482,I277182,I277513,I522291,I522279,I277530,I277556,I277564,I277164,I277595,I277173,I277626,I277643,I277185,I277674,I277176,I277167,I277170,I277188,I277774,I386107,I277800,I277808,I277825,I386083,I386098,I277842,I386110,I277868,I277876,I386095,I386086,I277902,I277910,I277927,I277944,I277961,I278001,I278009,I278026,I278043,I278060,I278091,I386101,I386092,I278108,I386104,I278134,I278142,I278173,I278204,I278221,I278252,I386089,I278352,I278378,I278386,I278403,I278420,I278446,I278454,I278480,I278488,I278505,I278522,I278539,I278579,I278587,I278604,I278621,I278638,I278669,I278686,I278712,I278720,I278751,I278782,I278799,I278830,I278930,I278956,I278964,I278981,I278998,I279024,I279032,I279058,I279066,I279083,I279100,I279117,I278913,I279157,I279165,I279182,I279199,I279216,I278916,I279247,I279264,I279290,I279298,I278898,I279329,I278907,I279360,I279377,I278919,I279408,I278910,I278901,I278904,I278922,I279508,I279534,I279542,I279559,I279576,I279602,I279610,I279636,I279644,I279661,I279678,I279695,I279735,I279743,I279760,I279777,I279794,I279825,I279842,I279868,I279876,I279907,I279938,I279955,I279986,I280086,I280112,I280120,I280137,I280154,I280180,I280188,I280214,I280222,I280239,I280256,I280273,I280069,I280313,I280321,I280338,I280355,I280372,I280072,I280403,I280420,I280446,I280454,I280054,I280485,I280063,I280516,I280533,I280075,I280564,I280066,I280057,I280060,I280078,I280664,I437106,I280690,I280698,I280715,I437103,I437121,I280732,I437118,I280758,I280766,I437100,I280792,I280800,I280817,I280834,I280851,I437112,I280891,I280899,I280916,I280933,I280950,I280981,I437115,I280998,I281024,I281032,I281063,I281094,I281111,I281142,I437109,I281242,I281268,I281276,I281293,I281310,I281336,I281344,I281370,I281378,I281395,I281412,I281429,I281469,I281477,I281494,I281511,I281528,I281559,I281576,I281602,I281610,I281641,I281672,I281689,I281720,I281820,I281846,I281854,I281871,I281888,I281914,I281922,I281948,I281956,I281973,I281990,I282007,I282047,I282055,I282072,I282089,I282106,I282137,I282154,I282180,I282188,I282219,I282250,I282267,I282298,I282398,I362706,I282424,I282432,I282449,I362694,I362712,I282466,I362709,I282492,I282500,I362700,I362697,I282526,I282534,I282551,I282568,I282585,I282381,I362691,I282625,I282633,I282650,I282667,I282684,I282384,I282715,I282732,I282758,I282766,I282366,I282797,I282375,I282828,I282845,I282387,I282876,I362703,I282378,I282369,I282372,I282390,I282976,I414531,I283002,I283010,I283027,I414507,I414522,I283044,I414534,I283070,I283078,I414519,I414510,I283104,I283112,I283129,I283146,I283163,I282959,I283203,I283211,I283228,I283245,I283262,I282962,I283293,I414525,I414516,I283310,I414528,I283336,I283344,I282944,I283375,I282953,I283406,I283423,I282965,I283454,I414513,I282956,I282947,I282950,I282968,I283554,I283580,I283588,I283605,I283622,I283648,I283656,I283682,I283690,I283707,I283724,I283741,I283781,I283789,I283806,I283823,I283840,I283871,I283888,I283914,I283922,I283953,I283984,I284001,I284032,I284132,I284158,I284166,I284183,I284200,I284226,I284234,I284260,I284268,I284285,I284302,I284319,I284359,I284367,I284384,I284401,I284418,I284449,I284466,I284492,I284500,I284531,I284562,I284579,I284610,I284710,I407425,I284736,I284744,I284761,I407401,I407416,I284778,I407428,I284804,I284812,I407413,I407404,I284838,I284846,I284863,I284880,I284897,I284693,I284937,I284945,I284962,I284979,I284996,I284696,I285027,I407419,I407410,I285044,I407422,I285070,I285078,I284678,I285109,I284687,I285140,I285157,I284699,I285188,I407407,I284690,I284681,I284684,I284702,I285288,I285314,I285322,I285339,I285356,I285382,I285390,I285416,I285424,I285441,I285458,I285475,I285271,I285515,I285523,I285540,I285557,I285574,I285274,I285605,I285622,I285648,I285656,I285256,I285687,I285265,I285718,I285735,I285277,I285766,I285268,I285259,I285262,I285280,I285866,I285892,I285900,I285917,I285934,I285960,I285968,I285994,I286002,I286019,I286036,I286053,I286093,I286101,I286118,I286135,I286152,I286183,I286200,I286226,I286234,I286265,I286296,I286313,I286344,I286444,I286470,I286478,I286495,I286512,I286538,I286546,I286572,I286580,I286597,I286614,I286631,I286427,I286671,I286679,I286696,I286713,I286730,I286430,I286761,I286778,I286804,I286812,I286412,I286843,I286421,I286874,I286891,I286433,I286922,I286424,I286415,I286418,I286436,I287022,I287048,I287056,I287073,I287090,I287116,I287124,I287150,I287158,I287175,I287192,I287209,I287249,I287257,I287274,I287291,I287308,I287339,I287356,I287382,I287390,I287421,I287452,I287469,I287500,I287600,I287626,I287634,I287651,I287668,I287694,I287702,I287728,I287736,I287753,I287770,I287787,I287827,I287835,I287852,I287869,I287886,I287917,I287934,I287960,I287968,I287999,I288030,I288047,I288078,I288178,I288204,I288212,I288229,I288246,I288272,I288280,I288306,I288314,I288331,I288348,I288365,I288405,I288413,I288430,I288447,I288464,I288495,I288512,I288538,I288546,I288577,I288608,I288625,I288656,I288756,I288782,I288790,I288807,I288824,I288850,I288858,I288884,I288892,I288909,I288926,I288943,I288739,I288983,I288991,I289008,I289025,I289042,I288742,I289073,I289090,I289116,I289124,I288724,I289155,I288733,I289186,I289203,I288745,I289234,I288736,I288727,I288730,I288748,I289334,I289360,I289368,I289385,I289402,I289428,I289436,I289462,I289470,I289487,I289504,I289521,I289317,I289561,I289569,I289586,I289603,I289620,I289320,I289651,I289668,I289694,I289702,I289302,I289733,I289311,I289764,I289781,I289323,I289812,I289314,I289305,I289308,I289326,I289912,I289938,I289946,I289963,I289980,I290006,I290014,I290040,I290048,I290065,I290082,I290099,I290139,I290147,I290164,I290181,I290198,I290229,I290246,I290272,I290280,I290311,I290342,I290359,I290390,I290490,I290516,I290524,I290541,I290558,I290584,I290592,I290618,I290626,I290643,I290660,I290677,I290473,I290717,I290725,I290742,I290759,I290776,I290476,I290807,I290824,I290850,I290858,I290458,I290889,I290467,I290920,I290937,I290479,I290968,I290470,I290461,I290464,I290482,I291068,I291094,I291102,I291119,I291136,I291162,I291170,I291196,I291204,I291221,I291238,I291255,I291295,I291303,I291320,I291337,I291354,I291385,I291402,I291428,I291436,I291467,I291498,I291515,I291546,I291646,I539552,I291672,I291680,I291697,I539537,I539525,I291714,I539540,I291740,I291748,I539543,I291774,I291782,I291799,I291816,I291833,I539531,I291873,I291881,I291898,I291915,I291932,I291963,I539528,I539534,I291980,I539549,I292006,I292014,I292045,I292076,I292093,I292124,I539546,I292224,I292250,I292258,I292275,I292292,I292318,I292326,I292352,I292360,I292377,I292394,I292411,I292207,I292451,I292459,I292476,I292493,I292510,I292210,I292541,I292558,I292584,I292592,I292192,I292623,I292201,I292654,I292671,I292213,I292702,I292204,I292195,I292198,I292216,I292802,I372719,I292828,I292836,I292853,I372707,I372725,I292870,I372722,I292896,I292904,I372713,I372710,I292930,I292938,I292955,I292972,I292989,I372704,I293029,I293037,I293054,I293071,I293088,I293119,I293136,I293162,I293170,I293201,I293232,I293249,I293280,I372716,I293380,I293406,I293414,I293431,I293448,I293474,I293482,I293508,I293516,I293533,I293550,I293567,I293607,I293615,I293632,I293649,I293666,I293697,I293714,I293740,I293748,I293779,I293810,I293827,I293858,I293958,I293984,I293992,I294009,I294026,I294052,I294060,I294086,I294094,I294111,I294128,I294145,I293941,I294185,I294193,I294210,I294227,I294244,I293944,I294275,I294292,I294318,I294326,I293926,I294357,I293935,I294388,I294405,I293947,I294436,I293938,I293929,I293932,I293950,I294536,I294562,I294570,I294587,I294604,I294630,I294638,I294664,I294672,I294689,I294706,I294723,I294763,I294771,I294788,I294805,I294822,I294853,I294870,I294896,I294904,I294935,I294966,I294983,I295014,I295114,I340045,I295140,I295148,I295165,I340033,I340051,I295182,I340048,I295208,I295216,I340039,I340036,I295242,I295250,I295267,I295284,I295301,I340030,I295341,I295349,I295366,I295383,I295400,I295431,I295448,I295474,I295482,I295513,I295544,I295561,I295592,I340042,I295692,I518394,I295718,I295726,I295743,I518397,I518406,I295760,I518409,I295786,I295794,I518418,I518400,I295820,I295828,I295845,I295862,I295879,I295919,I295927,I295944,I295961,I295978,I296009,I518415,I296026,I518412,I296052,I296060,I296091,I296122,I296139,I296170,I518403,I296270,I547882,I296296,I296304,I296321,I547867,I547855,I296338,I547870,I296364,I296372,I547873,I296398,I296406,I296423,I296440,I296457,I296253,I547861,I296497,I296505,I296522,I296539,I296556,I296256,I296587,I547858,I547864,I296604,I547879,I296630,I296638,I296238,I296669,I296247,I296700,I296717,I296259,I296748,I547876,I296250,I296241,I296244,I296262,I296848,I296874,I296882,I296899,I296916,I296942,I296950,I296976,I296984,I297001,I297018,I297035,I297075,I297083,I297100,I297117,I297134,I297165,I297182,I297208,I297216,I297247,I297278,I297295,I297326,I297426,I366395,I297452,I297460,I297477,I366383,I366401,I297494,I366398,I297520,I297528,I366389,I366386,I297554,I297562,I297579,I297596,I297613,I297409,I366380,I297653,I297661,I297678,I297695,I297712,I297412,I297743,I297760,I297786,I297794,I297394,I297825,I297403,I297856,I297873,I297415,I297904,I366392,I297406,I297397,I297400,I297418,I298004,I516218,I298030,I298038,I298055,I516221,I516230,I298072,I516233,I298098,I298106,I516242,I516224,I298132,I298140,I298157,I298174,I298191,I298231,I298239,I298256,I298273,I298290,I298321,I516239,I298338,I516236,I298364,I298372,I298403,I298434,I298451,I298482,I516227,I298582,I298608,I298616,I298633,I298650,I298676,I298684,I298710,I298718,I298735,I298752,I298769,I298565,I298809,I298817,I298834,I298851,I298868,I298568,I298899,I298916,I298942,I298950,I298550,I298981,I298559,I299012,I299029,I298571,I299060,I298562,I298553,I298556,I298574,I299160,I553832,I299186,I299194,I299211,I553817,I553805,I299228,I553820,I299254,I299262,I553823,I299288,I299296,I299313,I299330,I299347,I553811,I299387,I299395,I299412,I299429,I299446,I299477,I553808,I553814,I299494,I553829,I299520,I299528,I299559,I299590,I299607,I299638,I553826,I299738,I299764,I299772,I299789,I299806,I299832,I299840,I299866,I299874,I299891,I299908,I299925,I299965,I299973,I299990,I300007,I300024,I300055,I300072,I300098,I300106,I300137,I300168,I300185,I300216,I300316,I524004,I300342,I300350,I300367,I524028,I524010,I300384,I524016,I300410,I300418,I524022,I524007,I300444,I300452,I300469,I300486,I300503,I300299,I524019,I300543,I300551,I300568,I300585,I300602,I300302,I300633,I524025,I524013,I300650,I300676,I300684,I300284,I300715,I300293,I300746,I300763,I300305,I300794,I300296,I300287,I300290,I300308,I300894,I482440,I300920,I300928,I300945,I482422,I482434,I300962,I482437,I300988,I300996,I482431,I482428,I301022,I301030,I301047,I301064,I301081,I482446,I301121,I301129,I301146,I301163,I301180,I301211,I482425,I301228,I301254,I301262,I301293,I301324,I301341,I301372,I482443,I301472,I447204,I301498,I301506,I301523,I447201,I447219,I301540,I447216,I301566,I301574,I447198,I301600,I301608,I301625,I301642,I301659,I447210,I301699,I301707,I301724,I301741,I301758,I301789,I447213,I301806,I301832,I301840,I301871,I301902,I301919,I301950,I447207,I302050,I530940,I302076,I302084,I302101,I530964,I530946,I302118,I530952,I302144,I302152,I530958,I530943,I302178,I302186,I302203,I302220,I302237,I530955,I302277,I302285,I302302,I302319,I302336,I302367,I530961,I530949,I302384,I302410,I302418,I302449,I302480,I302497,I302528,I302628,I365868,I302654,I302662,I302679,I365856,I365874,I302696,I365871,I302722,I302730,I365862,I365859,I302756,I302764,I302781,I302798,I302815,I365853,I302855,I302863,I302880,I302897,I302914,I302945,I302962,I302988,I302996,I303027,I303058,I303075,I303106,I365865,I303206,I485330,I303232,I303240,I303257,I485312,I485324,I303274,I485327,I303300,I303308,I485321,I485318,I303334,I303342,I303359,I303376,I303393,I303189,I485336,I303433,I303441,I303458,I303475,I303492,I303192,I303523,I485315,I303540,I303566,I303574,I303174,I303605,I303183,I303636,I303653,I303195,I303684,I485333,I303186,I303177,I303180,I303198,I303784,I357436,I303810,I303818,I303835,I357424,I357442,I303852,I357439,I303878,I303886,I357430,I357427,I303912,I303920,I303937,I303954,I303971,I303767,I357421,I304011,I304019,I304036,I304053,I304070,I303770,I304101,I304118,I304144,I304152,I303752,I304183,I303761,I304214,I304231,I303773,I304262,I357433,I303764,I303755,I303758,I303776,I304362,I333721,I304388,I304396,I304413,I333709,I333727,I304430,I333724,I304456,I304464,I333715,I333712,I304490,I304498,I304515,I304532,I304549,I304345,I333706,I304589,I304597,I304614,I304631,I304648,I304348,I304679,I304696,I304722,I304730,I304330,I304761,I304339,I304792,I304809,I304351,I304840,I333718,I304342,I304333,I304336,I304354,I304940,I304966,I304974,I304991,I305008,I305034,I305042,I305068,I305076,I305093,I305110,I305127,I305167,I305175,I305192,I305209,I305226,I305257,I305274,I305300,I305308,I305339,I305370,I305387,I305418,I305518,I380293,I305544,I305552,I305569,I380269,I380284,I305586,I380296,I305612,I305620,I380281,I380272,I305646,I305654,I305671,I305688,I305705,I305501,I305745,I305753,I305770,I305787,I305804,I305504,I305835,I380287,I380278,I305852,I380290,I305878,I305886,I305486,I305917,I305495,I305948,I305965,I305507,I305996,I380275,I305498,I305489,I305492,I305510,I306096,I306122,I306130,I306147,I306164,I306190,I306198,I306224,I306232,I306249,I306266,I306283,I306323,I306331,I306348,I306365,I306382,I306413,I306430,I306456,I306464,I306495,I306526,I306543,I306574,I306674,I306700,I306708,I306725,I306742,I306768,I306776,I306802,I306810,I306827,I306844,I306861,I306901,I306909,I306926,I306943,I306960,I306991,I307008,I307034,I307042,I307073,I307104,I307121,I307152,I307252,I465100,I307278,I307286,I307303,I465082,I465094,I307320,I465097,I307346,I307354,I465091,I465088,I307380,I307388,I307405,I307422,I307439,I307235,I465106,I307479,I307487,I307504,I307521,I307538,I307238,I307569,I465085,I307586,I307612,I307620,I307220,I307651,I307229,I307682,I307699,I307241,I307730,I465103,I307232,I307223,I307226,I307244,I307830,I307856,I307864,I307881,I307898,I307924,I307932,I307958,I307966,I307983,I308000,I308017,I308057,I308065,I308082,I308099,I308116,I308147,I308164,I308190,I308198,I308229,I308260,I308277,I308308,I308408,I351639,I308434,I308442,I308459,I351627,I351645,I308476,I351642,I308502,I308510,I351633,I351630,I308536,I308544,I308561,I308578,I308595,I308391,I351624,I308635,I308643,I308660,I308677,I308694,I308394,I308725,I308742,I308768,I308776,I308376,I308807,I308385,I308838,I308855,I308397,I308886,I351636,I308388,I308379,I308382,I308400,I308986,I534408,I309012,I309020,I309037,I534432,I534414,I309054,I534420,I309080,I309088,I534426,I534411,I309114,I309122,I309139,I309156,I309173,I308969,I534423,I309213,I309221,I309238,I309255,I309272,I308972,I309303,I534429,I534417,I309320,I309346,I309354,I308954,I309385,I308963,I309416,I309433,I308975,I309464,I308966,I308957,I308960,I308978,I309564,I309590,I309598,I309615,I309632,I309658,I309666,I309692,I309700,I309717,I309734,I309751,I309791,I309799,I309816,I309833,I309850,I309881,I309898,I309924,I309932,I309963,I309994,I310011,I310042,I310142,I310168,I310176,I310193,I310210,I310236,I310244,I310270,I310278,I310295,I310312,I310329,I310125,I310369,I310377,I310394,I310411,I310428,I310128,I310459,I310476,I310502,I310510,I310110,I310541,I310119,I310572,I310589,I310131,I310620,I310122,I310113,I310116,I310134,I310720,I310746,I310754,I310771,I310788,I310814,I310822,I310848,I310856,I310873,I310890,I310907,I310947,I310955,I310972,I310989,I311006,I311037,I311054,I311080,I311088,I311119,I311150,I311167,I311198,I311298,I455274,I311324,I311332,I311349,I455256,I455268,I311366,I455271,I311392,I311400,I455265,I455262,I311426,I311434,I311451,I311468,I311485,I311281,I455280,I311525,I311533,I311550,I311567,I311584,I311284,I311615,I455259,I311632,I311658,I311666,I311266,I311697,I311275,I311728,I311745,I311287,I311776,I455277,I311278,I311269,I311272,I311290,I311876,I311902,I311910,I311927,I311944,I311970,I311978,I312004,I312012,I312029,I312046,I312063,I311859,I312103,I312111,I312128,I312145,I312162,I311862,I312193,I312210,I312236,I312244,I311844,I312275,I311853,I312306,I312323,I311865,I312354,I311856,I311847,I311850,I311868,I312454,I499202,I312480,I312488,I312505,I499184,I499196,I312522,I499199,I312548,I312556,I499193,I499190,I312582,I312590,I312607,I312624,I312641,I312437,I499208,I312681,I312689,I312706,I312723,I312740,I312440,I312771,I499187,I312788,I312814,I312822,I312422,I312853,I312431,I312884,I312901,I312443,I312932,I499205,I312434,I312425,I312428,I312446,I313032,I536140,I313058,I313066,I313083,I536128,I536146,I313100,I536137,I313126,I313134,I536152,I536149,I313160,I313168,I313185,I313202,I313219,I536131,I313259,I313267,I313284,I313301,I313318,I313349,I536125,I313366,I536134,I313392,I313400,I313431,I313462,I313479,I313510,I536143,I313610,I313636,I313644,I313661,I313678,I313704,I313712,I313738,I313746,I313763,I313780,I313797,I313593,I313837,I313845,I313862,I313879,I313896,I313596,I313927,I313944,I313970,I313978,I313578,I314009,I313587,I314040,I314057,I313599,I314088,I313590,I313581,I313584,I313602,I314188,I314214,I314222,I314239,I314256,I314282,I314290,I314316,I314324,I314341,I314358,I314375,I314415,I314423,I314440,I314457,I314474,I314505,I314522,I314548,I314556,I314587,I314618,I314635,I314666,I314766,I420991,I314792,I314800,I314817,I420967,I420982,I314834,I420994,I314860,I314868,I420979,I420970,I314894,I314902,I314919,I314936,I314953,I314993,I315001,I315018,I315035,I315052,I315083,I420985,I420976,I315100,I420988,I315126,I315134,I315165,I315196,I315213,I315244,I420973,I315344,I315370,I315378,I315395,I315412,I315438,I315446,I315472,I315480,I315497,I315514,I315531,I315571,I315579,I315596,I315613,I315630,I315661,I315678,I315704,I315712,I315743,I315774,I315791,I315822,I315922,I315948,I315956,I315973,I315990,I316016,I316024,I316050,I316058,I316075,I316092,I316109,I316149,I316157,I316174,I316191,I316208,I316239,I316256,I316282,I316290,I316321,I316352,I316369,I316400,I316500,I316526,I316534,I316551,I316568,I316594,I316602,I316628,I316636,I316653,I316670,I316687,I316483,I316727,I316735,I316752,I316769,I316786,I316486,I316817,I316834,I316860,I316868,I316468,I316899,I316477,I316930,I316947,I316489,I316978,I316480,I316471,I316474,I316492,I317078,I317104,I317112,I317129,I317146,I317172,I317180,I317206,I317214,I317231,I317248,I317265,I317305,I317313,I317330,I317347,I317364,I317395,I317412,I317438,I317446,I317477,I317508,I317525,I317556,I317656,I508058,I317682,I317690,I317707,I508061,I508070,I317724,I508073,I317750,I317758,I508082,I508064,I317784,I317792,I317809,I317826,I317843,I317639,I317883,I317891,I317908,I317925,I317942,I317642,I317973,I508079,I317990,I508076,I318016,I318024,I317624,I318055,I317633,I318086,I318103,I317645,I318134,I508067,I317636,I317627,I317630,I317648,I318234,I568112,I318260,I318268,I318285,I568097,I568085,I318302,I568100,I318328,I318336,I568103,I318362,I318370,I318387,I318404,I318421,I568091,I318461,I318469,I318486,I318503,I318520,I318551,I568088,I568094,I318568,I568109,I318594,I318602,I318633,I318664,I318681,I318712,I568106,I318812,I318838,I318846,I318863,I318880,I318906,I318914,I318940,I318948,I318965,I318982,I318999,I318795,I319039,I319047,I319064,I319081,I319098,I318798,I319129,I319146,I319172,I319180,I318780,I319211,I318789,I319242,I319259,I318801,I319290,I318792,I318783,I318786,I318804,I319390,I319416,I319424,I319441,I319458,I319484,I319492,I319518,I319526,I319543,I319560,I319577,I319617,I319625,I319642,I319659,I319676,I319707,I319724,I319750,I319758,I319789,I319820,I319837,I319868,I319968,I532096,I319994,I320002,I320019,I532120,I532102,I320036,I532108,I320062,I320070,I532114,I532099,I320096,I320104,I320121,I320138,I320155,I319951,I532111,I320195,I320203,I320220,I320237,I320254,I319954,I320285,I532117,I532105,I320302,I320328,I320336,I319936,I320367,I319945,I320398,I320415,I319957,I320446,I319948,I319939,I319942,I319960,I320546,I320572,I320580,I320597,I320614,I320640,I320648,I320674,I320682,I320699,I320716,I320733,I320529,I320773,I320781,I320798,I320815,I320832,I320532,I320863,I320880,I320906,I320914,I320514,I320945,I320523,I320976,I320993,I320535,I321024,I320526,I320517,I320520,I320538,I321124,I467412,I321150,I321158,I321175,I467394,I467406,I321192,I467409,I321218,I321226,I467403,I467400,I321252,I321260,I321277,I321294,I321311,I321107,I467418,I321351,I321359,I321376,I321393,I321410,I321110,I321441,I467397,I321458,I321484,I321492,I321092,I321523,I321101,I321554,I321571,I321113,I321602,I467415,I321104,I321095,I321098,I321116,I321702,I466834,I321728,I321736,I321753,I466816,I466828,I321770,I466831,I321796,I321804,I466825,I466822,I321830,I321838,I321855,I321872,I321889,I321685,I466840,I321929,I321937,I321954,I321971,I321988,I321688,I322019,I466819,I322036,I322062,I322070,I321670,I322101,I321679,I322132,I322149,I321691,I322180,I466837,I321682,I321673,I321676,I321694,I322280,I322306,I322314,I322331,I322348,I322374,I322382,I322408,I322416,I322433,I322450,I322467,I322507,I322515,I322532,I322549,I322566,I322597,I322614,I322640,I322648,I322679,I322710,I322727,I322758,I322858,I322884,I322892,I322909,I322926,I322952,I322960,I322986,I322994,I323011,I323028,I323045,I323085,I323093,I323110,I323127,I323144,I323175,I323192,I323218,I323226,I323257,I323288,I323305,I323336,I323436,I323462,I323470,I323487,I323504,I323530,I323538,I323564,I323572,I323589,I323606,I323623,I323663,I323671,I323688,I323705,I323722,I323753,I323770,I323796,I323804,I323835,I323866,I323883,I323914,I324014,I324040,I324048,I324065,I324082,I324108,I324116,I324142,I324150,I324167,I324184,I324201,I324241,I324249,I324266,I324283,I324300,I324331,I324348,I324374,I324382,I324413,I324444,I324461,I324492,I324592,I457008,I324618,I324626,I324643,I456990,I457002,I324660,I457005,I324686,I324694,I456999,I456996,I324720,I324728,I324745,I324762,I324779,I324575,I457014,I324819,I324827,I324844,I324861,I324878,I324578,I324909,I456993,I324926,I324952,I324960,I324560,I324991,I324569,I325022,I325039,I324581,I325070,I457011,I324572,I324563,I324566,I324584,I325170,I428691,I325196,I325204,I325221,I428688,I428706,I325238,I428703,I325264,I325272,I428685,I325298,I325306,I325323,I325340,I325357,I428697,I325397,I325405,I325422,I325439,I325456,I325487,I428700,I325504,I325530,I325538,I325569,I325600,I325617,I325648,I428694,I325748,I325774,I325782,I325799,I325816,I325842,I325850,I325876,I325884,I325901,I325918,I325935,I325731,I325975,I325983,I326000,I326017,I326034,I325734,I326065,I326082,I326108,I326116,I325716,I326147,I325725,I326178,I326195,I325737,I326226,I325728,I325719,I325722,I325740,I326326,I383523,I326352,I326360,I326377,I383499,I383514,I326394,I383526,I326420,I326428,I383511,I383502,I326454,I326462,I326479,I326496,I326513,I326309,I326553,I326561,I326578,I326595,I326612,I326312,I326643,I383517,I383508,I326660,I383520,I326686,I326694,I326294,I326725,I326303,I326756,I326773,I326315,I326804,I383505,I326306,I326297,I326300,I326318,I326904,I326930,I326938,I326955,I326972,I326998,I327006,I327032,I327040,I327057,I327074,I327091,I326887,I327131,I327139,I327156,I327173,I327190,I326890,I327221,I327238,I327264,I327272,I326872,I327303,I326881,I327334,I327351,I326893,I327382,I326884,I326875,I326878,I326896,I327482,I327508,I327516,I327533,I327550,I327576,I327584,I327610,I327618,I327635,I327652,I327669,I327465,I327709,I327717,I327734,I327751,I327768,I327468,I327799,I327816,I327842,I327850,I327450,I327881,I327459,I327912,I327929,I327471,I327960,I327462,I327453,I327456,I327474,I328060,I328086,I328094,I328111,I328128,I328154,I328162,I328188,I328196,I328213,I328230,I328247,I328287,I328295,I328312,I328329,I328346,I328377,I328394,I328420,I328428,I328459,I328490,I328507,I328538,I328638,I328664,I328672,I328689,I328706,I328732,I328740,I328766,I328774,I328791,I328808,I328825,I328621,I328865,I328873,I328890,I328907,I328924,I328624,I328955,I328972,I328998,I329006,I328606,I329037,I328615,I329068,I329085,I328627,I329116,I328618,I328609,I328612,I328630,I329216,I394505,I329242,I329250,I329267,I394481,I394496,I329284,I394508,I329310,I329318,I394493,I394484,I329344,I329352,I329369,I329386,I329403,I329199,I329443,I329451,I329468,I329485,I329502,I329202,I329533,I394499,I394490,I329550,I394502,I329576,I329584,I329184,I329615,I329193,I329646,I329663,I329205,I329694,I394487,I329196,I329187,I329190,I329208,I329794,I329820,I329828,I329845,I329862,I329888,I329896,I329922,I329930,I329947,I329964,I329981,I330021,I330029,I330046,I330063,I330080,I330111,I330128,I330154,I330162,I330193,I330224,I330241,I330272,I330372,I362179,I330398,I330406,I330423,I362167,I362185,I330440,I362182,I330466,I330474,I362173,I362170,I330500,I330508,I330525,I330542,I330559,I330355,I362164,I330599,I330607,I330624,I330641,I330658,I330358,I330689,I330706,I330732,I330740,I330340,I330771,I330349,I330802,I330819,I330361,I330850,I362176,I330352,I330343,I330346,I330364,I330950,I381585,I330976,I330984,I331001,I381561,I381576,I331018,I381588,I331044,I331052,I381573,I381564,I331078,I331086,I331103,I331120,I331137,I330933,I331177,I331185,I331202,I331219,I331236,I330936,I331267,I381579,I381570,I331284,I381582,I331310,I331318,I330918,I331349,I330927,I331380,I331397,I330939,I331428,I381567,I330930,I330921,I330924,I330942,I331528,I355855,I331554,I331562,I331579,I355843,I355861,I331596,I355858,I331622,I331630,I355849,I355846,I331656,I331664,I331681,I331698,I331715,I331511,I355840,I331755,I331763,I331780,I331797,I331814,I331514,I331845,I331862,I331888,I331896,I331496,I331927,I331505,I331958,I331975,I331517,I332006,I355852,I331508,I331499,I331502,I331520,I332106,I408071,I332132,I332140,I332157,I408047,I408062,I332174,I408074,I332200,I332208,I408059,I408050,I332234,I332242,I332259,I332276,I332293,I332089,I332333,I332341,I332358,I332375,I332392,I332092,I332423,I408065,I408056,I332440,I408068,I332466,I332474,I332074,I332505,I332083,I332536,I332553,I332095,I332584,I408053,I332086,I332077,I332080,I332098,I332681,I461632,I332707,I332715,I332732,I461614,I332749,I461620,I332775,I461617,I332806,I332814,I461626,I332831,I332857,I332865,I461638,I332905,I332941,I461629,I461623,I332958,I332984,I332992,I333009,I333040,I461635,I333057,I333074,I333105,I333136,I333153,I333208,I460476,I333234,I333242,I333259,I460458,I333276,I460464,I333302,I333197,I460461,I333333,I333341,I460470,I333358,I333384,I333392,I333200,I460482,I333432,I333191,I333182,I333468,I460473,I460467,I333485,I333511,I333519,I333536,I333185,I333567,I460479,I333584,I333601,I333194,I333632,I333179,I333663,I333680,I333188,I333735,I333761,I333769,I333786,I333803,I333829,I333860,I333868,I333885,I333911,I333919,I333959,I333995,I334012,I334038,I334046,I334063,I334094,I334111,I334128,I334159,I334190,I334207,I334262,I334288,I334296,I334313,I334330,I334356,I334387,I334395,I334412,I334438,I334446,I334486,I334522,I334539,I334565,I334573,I334590,I334621,I334638,I334655,I334686,I334717,I334734,I334789,I334815,I334823,I334840,I334857,I334883,I334778,I334914,I334922,I334939,I334965,I334973,I334781,I335013,I334772,I334763,I335049,I335066,I335092,I335100,I335117,I334766,I335148,I335165,I335182,I334775,I335213,I334760,I335244,I335261,I334769,I335316,I335342,I335350,I335367,I335384,I335410,I335441,I335449,I335466,I335492,I335500,I335540,I335576,I335593,I335619,I335627,I335644,I335675,I335692,I335709,I335740,I335771,I335788,I335843,I335869,I335877,I335894,I335911,I335937,I335832,I335968,I335976,I335993,I336019,I336027,I335835,I336067,I335826,I335817,I336103,I336120,I336146,I336154,I336171,I335820,I336202,I336219,I336236,I335829,I336267,I335814,I336298,I336315,I335823,I336370,I336396,I336404,I336421,I336438,I336464,I336495,I336503,I336520,I336546,I336554,I336594,I336630,I336647,I336673,I336681,I336698,I336729,I336746,I336763,I336794,I336825,I336842,I336897,I336923,I336931,I336948,I336965,I336991,I336886,I337022,I337030,I337047,I337073,I337081,I336889,I337121,I336880,I336871,I337157,I337174,I337200,I337208,I337225,I336874,I337256,I337273,I337290,I336883,I337321,I336868,I337352,I337369,I336877,I337424,I337450,I337458,I337475,I337492,I337518,I337413,I337549,I337557,I337574,I337600,I337608,I337416,I337648,I337407,I337398,I337684,I337701,I337727,I337735,I337752,I337401,I337783,I337800,I337817,I337410,I337848,I337395,I337879,I337896,I337404,I337951,I337977,I337985,I338002,I338019,I338045,I337940,I338076,I338084,I338101,I338127,I338135,I337943,I338175,I337934,I337925,I338211,I338228,I338254,I338262,I338279,I337928,I338310,I338327,I338344,I337937,I338375,I337922,I338406,I338423,I337931,I338478,I338504,I338512,I338529,I338546,I338572,I338603,I338611,I338628,I338654,I338662,I338702,I338738,I338755,I338781,I338789,I338806,I338837,I338854,I338871,I338902,I338933,I338950,I339005,I417094,I339031,I339039,I339056,I417109,I417091,I339073,I339099,I417100,I339130,I339138,I417118,I339155,I339181,I339189,I417115,I339229,I339265,I417112,I417103,I339282,I417097,I339308,I339316,I339333,I339364,I417106,I339381,I339398,I339429,I339460,I339477,I339532,I339558,I339566,I339583,I339600,I339626,I339657,I339665,I339682,I339708,I339716,I339756,I339792,I339809,I339835,I339843,I339860,I339891,I339908,I339925,I339956,I339987,I340004,I340059,I340085,I340093,I340110,I340127,I340153,I340184,I340192,I340209,I340235,I340243,I340283,I340319,I340336,I340362,I340370,I340387,I340418,I340435,I340452,I340483,I340514,I340531,I340586,I340612,I340620,I340637,I340654,I340680,I340711,I340719,I340736,I340762,I340770,I340810,I340846,I340863,I340889,I340897,I340914,I340945,I340962,I340979,I341010,I341041,I341058,I341113,I491688,I341139,I341147,I341164,I491670,I341181,I491676,I341207,I491673,I341238,I341246,I491682,I341263,I341289,I341297,I491694,I341337,I341373,I491685,I491679,I341390,I341416,I341424,I341441,I341472,I491691,I341489,I341506,I341537,I341568,I341585,I341640,I513510,I341666,I341674,I341691,I513516,I513498,I341708,I513507,I341734,I513513,I341765,I341773,I513501,I341790,I341816,I341824,I513519,I341864,I341900,I513504,I341917,I513522,I341943,I341951,I341968,I341999,I342016,I342033,I342064,I342095,I342112,I342167,I342193,I342201,I342218,I342235,I342261,I342292,I342300,I342317,I342343,I342351,I342391,I342427,I342444,I342470,I342478,I342495,I342526,I342543,I342560,I342591,I342622,I342639,I342694,I536692,I342720,I342728,I342745,I536686,I536704,I342762,I536689,I342788,I342683,I536710,I342819,I342827,I536695,I342844,I342870,I342878,I342686,I536707,I342918,I342677,I342668,I342954,I536698,I536713,I342971,I536701,I342997,I343005,I343022,I342671,I343053,I343070,I343087,I342680,I343118,I342665,I343149,I343166,I342674,I343221,I484174,I343247,I343255,I343272,I484156,I343289,I484162,I343315,I343210,I484159,I343346,I343354,I484168,I343371,I343397,I343405,I343213,I484180,I343445,I343204,I343195,I343481,I484171,I484165,I343498,I343524,I343532,I343549,I343198,I343580,I484177,I343597,I343614,I343207,I343645,I343192,I343676,I343693,I343201,I343748,I469724,I343774,I343782,I343799,I469706,I343816,I469712,I343842,I343737,I469709,I343873,I343881,I469718,I343898,I343924,I343932,I343740,I469730,I343972,I343731,I343722,I344008,I469721,I469715,I344025,I344051,I344059,I344076,I343725,I344107,I469727,I344124,I344141,I343734,I344172,I343719,I344203,I344220,I343728,I344275,I344301,I344309,I344326,I344343,I344369,I344264,I344400,I344408,I344425,I344451,I344459,I344267,I344499,I344258,I344249,I344535,I344552,I344578,I344586,I344603,I344252,I344634,I344651,I344668,I344261,I344699,I344246,I344730,I344747,I344255,I344802,I344828,I344836,I344853,I344870,I344896,I344791,I344927,I344935,I344952,I344978,I344986,I344794,I345026,I344785,I344776,I345062,I345079,I345105,I345113,I345130,I344779,I345161,I345178,I345195,I344788,I345226,I344773,I345257,I345274,I344782,I345329,I345355,I345363,I345380,I345397,I345423,I345454,I345462,I345479,I345505,I345513,I345553,I345589,I345606,I345632,I345640,I345657,I345688,I345705,I345722,I345753,I345784,I345801,I345856,I452384,I345882,I345890,I345907,I452366,I345924,I452372,I345950,I452369,I345981,I345989,I452378,I346006,I346032,I346040,I452390,I346080,I346116,I452381,I452375,I346133,I346159,I346167,I346184,I346215,I452387,I346232,I346249,I346280,I346311,I346328,I346383,I346409,I346417,I346434,I346451,I346477,I346372,I346508,I346516,I346533,I346559,I346567,I346375,I346607,I346366,I346357,I346643,I346660,I346686,I346694,I346711,I346360,I346742,I346759,I346776,I346369,I346807,I346354,I346838,I346855,I346363,I346910,I398360,I346936,I346944,I346961,I398375,I398357,I346978,I347004,I398366,I347035,I347043,I398384,I347060,I347086,I347094,I398381,I347134,I347170,I398378,I398369,I347187,I398363,I347213,I347221,I347238,I347269,I398372,I347286,I347303,I347334,I347365,I347382,I347437,I347463,I347471,I347488,I347505,I347531,I347562,I347570,I347587,I347613,I347621,I347661,I347697,I347714,I347740,I347748,I347765,I347796,I347813,I347830,I347861,I347892,I347909,I347964,I347990,I347998,I348015,I348032,I348058,I347953,I348089,I348097,I348114,I348140,I348148,I347956,I348188,I347947,I347938,I348224,I348241,I348267,I348275,I348292,I347941,I348323,I348340,I348357,I347950,I348388,I347935,I348419,I348436,I347944,I348491,I348517,I348525,I348542,I348559,I348585,I348480,I348616,I348624,I348641,I348667,I348675,I348483,I348715,I348474,I348465,I348751,I348768,I348794,I348802,I348819,I348468,I348850,I348867,I348884,I348477,I348915,I348462,I348946,I348963,I348471,I349018,I439914,I349044,I349052,I349069,I439923,I439911,I349086,I439908,I349112,I349007,I349143,I349151,I439905,I349168,I349194,I349202,I349010,I349242,I349001,I348992,I349278,I439926,I439917,I349295,I439920,I349321,I349329,I349346,I348995,I349377,I349394,I349411,I349004,I349442,I348989,I349473,I349490,I348998,I349545,I441597,I349571,I349579,I349596,I441606,I441594,I349613,I441591,I349639,I349670,I349678,I441588,I349695,I349721,I349729,I349769,I349805,I441609,I441600,I349822,I441603,I349848,I349856,I349873,I349904,I349921,I349938,I349969,I350000,I350017,I350072,I350098,I350106,I350123,I350140,I350166,I350197,I350205,I350222,I350248,I350256,I350296,I350332,I350349,I350375,I350383,I350400,I350431,I350448,I350465,I350496,I350527,I350544,I350599,I350625,I350633,I350650,I350667,I350693,I350724,I350732,I350749,I350775,I350783,I350823,I350859,I350876,I350902,I350910,I350927,I350958,I350975,I350992,I351023,I351054,I351071,I351126,I569290,I351152,I351160,I351177,I569287,I569296,I351194,I569275,I351220,I351115,I569278,I351251,I351259,I569293,I351276,I351302,I351310,I351118,I569299,I351350,I351109,I351100,I351386,I569281,I569302,I351403,I569284,I351429,I351437,I351454,I351103,I351485,I351502,I351519,I351112,I351550,I351097,I351581,I351598,I351106,I351653,I351679,I351687,I351704,I351721,I351747,I351778,I351786,I351803,I351829,I351837,I351877,I351913,I351930,I351956,I351964,I351981,I352012,I352029,I352046,I352077,I352108,I352125,I352180,I401590,I352206,I352214,I352231,I401605,I401587,I352248,I352274,I401596,I352305,I352313,I401614,I352330,I352356,I352364,I401611,I352404,I352440,I401608,I401599,I352457,I401593,I352483,I352491,I352508,I352539,I401602,I352556,I352573,I352604,I352635,I352652,I352707,I546680,I352733,I352741,I352758,I546677,I546686,I352775,I546665,I352801,I352696,I546668,I352832,I352840,I546683,I352857,I352883,I352891,I352699,I546689,I352931,I352690,I352681,I352967,I546671,I546692,I352984,I546674,I353010,I353018,I353035,I352684,I353066,I353083,I353100,I352693,I353131,I352678,I353162,I353179,I352687,I353234,I353260,I353268,I353285,I353302,I353328,I353223,I353359,I353367,I353384,I353410,I353418,I353226,I353458,I353217,I353208,I353494,I353511,I353537,I353545,I353562,I353211,I353593,I353610,I353627,I353220,I353658,I353205,I353689,I353706,I353214,I353761,I353787,I353795,I353812,I353829,I353855,I353886,I353894,I353911,I353937,I353945,I353985,I354021,I354038,I354064,I354072,I354089,I354120,I354137,I354154,I354185,I354216,I354233,I354288,I354314,I354322,I354339,I354356,I354382,I354413,I354421,I354438,I354464,I354472,I354512,I354548,I354565,I354591,I354599,I354616,I354647,I354664,I354681,I354712,I354743,I354760,I354815,I354841,I354849,I354866,I354883,I354909,I354940,I354948,I354965,I354991,I354999,I355039,I355075,I355092,I355118,I355126,I355143,I355174,I355191,I355208,I355239,I355270,I355287,I355342,I355368,I355376,I355393,I355410,I355436,I355467,I355475,I355492,I355518,I355526,I355566,I355602,I355619,I355645,I355653,I355670,I355701,I355718,I355735,I355766,I355797,I355814,I355869,I355895,I355903,I355920,I355937,I355963,I355994,I356002,I356019,I356045,I356053,I356093,I356129,I356146,I356172,I356180,I356197,I356228,I356245,I356262,I356293,I356324,I356341,I356396,I356422,I356430,I356447,I356464,I356490,I356521,I356529,I356546,I356572,I356580,I356620,I356656,I356673,I356699,I356707,I356724,I356755,I356772,I356789,I356820,I356851,I356868,I356923,I356949,I356957,I356974,I356991,I357017,I356912,I357048,I357056,I357073,I357099,I357107,I356915,I357147,I356906,I356897,I357183,I357200,I357226,I357234,I357251,I356900,I357282,I357299,I357316,I356909,I357347,I356894,I357378,I357395,I356903,I357450,I502630,I357476,I357484,I357501,I502636,I502618,I357518,I502627,I357544,I502633,I357575,I357583,I502621,I357600,I357626,I357634,I502639,I357674,I357710,I502624,I357727,I502642,I357753,I357761,I357778,I357809,I357826,I357843,I357874,I357905,I357922,I357977,I358003,I358011,I358028,I358045,I358071,I358102,I358110,I358127,I358153,I358161,I358201,I358237,I358254,I358280,I358288,I358305,I358336,I358353,I358370,I358401,I358432,I358449,I358504,I358530,I358538,I358555,I358572,I358598,I358493,I358629,I358637,I358654,I358680,I358688,I358496,I358728,I358487,I358478,I358764,I358781,I358807,I358815,I358832,I358481,I358863,I358880,I358897,I358490,I358928,I358475,I358959,I358976,I358484,I359031,I382210,I359057,I359065,I359082,I382225,I382207,I359099,I359125,I382216,I359156,I359164,I382234,I359181,I359207,I359215,I382231,I359255,I359291,I382228,I382219,I359308,I382213,I359334,I359342,I359359,I359390,I382222,I359407,I359424,I359455,I359486,I359503,I359558,I532692,I359584,I359592,I359609,I532674,I532677,I359626,I532689,I359652,I532698,I359683,I359691,I532683,I359708,I359734,I359742,I532695,I359782,I359818,I532686,I532680,I359835,I359861,I359869,I359886,I359917,I359934,I359951,I359982,I360013,I360030,I360085,I360111,I360119,I360136,I360153,I360179,I360210,I360218,I360235,I360261,I360269,I360309,I360345,I360362,I360388,I360396,I360413,I360444,I360461,I360478,I360509,I360540,I360557,I360612,I421616,I360638,I360646,I360663,I421631,I421613,I360680,I360706,I421622,I360737,I360745,I421640,I360762,I360788,I360796,I421637,I360836,I360872,I421634,I421625,I360889,I421619,I360915,I360923,I360940,I360971,I421628,I360988,I361005,I361036,I361067,I361084,I361139,I361165,I361173,I361190,I361207,I361233,I361128,I361264,I361272,I361289,I361315,I361323,I361131,I361363,I361122,I361113,I361399,I361416,I361442,I361450,I361467,I361116,I361498,I361515,I361532,I361125,I361563,I361110,I361594,I361611,I361119,I361666,I361692,I361700,I361717,I361734,I361760,I361791,I361799,I361816,I361842,I361850,I361890,I361926,I361943,I361969,I361977,I361994,I362025,I362042,I362059,I362090,I362121,I362138,I362193,I453540,I362219,I362227,I362244,I453522,I362261,I453528,I362287,I453525,I362318,I362326,I453534,I362343,I362369,I362377,I453546,I362417,I362453,I453537,I453531,I362470,I362496,I362504,I362521,I362552,I453543,I362569,I362586,I362617,I362648,I362665,I362720,I362746,I362754,I362771,I362788,I362814,I362845,I362853,I362870,I362896,I362904,I362944,I362980,I362997,I363023,I363031,I363048,I363079,I363096,I363113,I363144,I363175,I363192,I363247,I363273,I363281,I363298,I363315,I363341,I363236,I363372,I363380,I363397,I363423,I363431,I363239,I363471,I363230,I363221,I363507,I363524,I363550,I363558,I363575,I363224,I363606,I363623,I363640,I363233,I363671,I363218,I363702,I363719,I363227,I363774,I363800,I363808,I363825,I363842,I363868,I363899,I363907,I363924,I363950,I363958,I363998,I364034,I364051,I364077,I364085,I364102,I364133,I364150,I364167,I364198,I364229,I364246,I364301,I364327,I364335,I364352,I364369,I364395,I364290,I364426,I364434,I364451,I364477,I364485,I364293,I364525,I364284,I364275,I364561,I364578,I364604,I364612,I364629,I364278,I364660,I364677,I364694,I364287,I364725,I364272,I364756,I364773,I364281,I364828,I528068,I364854,I364862,I364879,I528050,I528053,I364896,I528065,I364922,I528074,I364953,I364961,I528059,I364978,I365004,I365012,I528071,I365052,I365088,I528062,I528056,I365105,I365131,I365139,I365156,I365187,I365204,I365221,I365252,I365283,I365300,I365355,I365381,I365389,I365406,I365423,I365449,I365480,I365488,I365505,I365531,I365539,I365579,I365615,I365632,I365658,I365666,I365683,I365714,I365731,I365748,I365779,I365810,I365827,I365882,I413218,I365908,I365916,I365933,I413233,I413215,I365950,I365976,I413224,I366007,I366015,I413242,I366032,I366058,I366066,I413239,I366106,I366142,I413236,I413227,I366159,I413221,I366185,I366193,I366210,I366241,I413230,I366258,I366275,I366306,I366337,I366354,I366409,I366435,I366443,I366460,I366477,I366503,I366534,I366542,I366559,I366585,I366593,I366633,I366669,I366686,I366712,I366720,I366737,I366768,I366785,I366802,I366833,I366864,I366881,I366936,I555010,I366962,I366970,I366987,I555007,I555016,I367004,I554995,I367030,I554998,I367061,I367069,I555013,I367086,I367112,I367120,I555019,I367160,I367196,I555001,I555022,I367213,I555004,I367239,I367247,I367264,I367295,I367312,I367329,I367360,I367391,I367408,I367463,I367489,I367497,I367514,I367531,I367557,I367588,I367596,I367613,I367639,I367647,I367687,I367723,I367740,I367766,I367774,I367791,I367822,I367839,I367856,I367887,I367918,I367935,I367990,I538945,I368016,I368024,I368041,I538942,I538951,I368058,I538930,I368084,I538933,I368115,I368123,I538948,I368140,I368166,I368174,I538954,I368214,I368250,I538936,I538957,I368267,I538939,I368293,I368301,I368318,I368349,I368366,I368383,I368414,I368445,I368462,I368517,I368543,I368551,I368568,I368585,I368611,I368506,I368642,I368650,I368667,I368693,I368701,I368509,I368741,I368500,I368491,I368777,I368794,I368820,I368828,I368845,I368494,I368876,I368893,I368910,I368503,I368941,I368488,I368972,I368989,I368497,I369044,I473770,I369070,I369078,I369095,I473752,I369112,I473758,I369138,I369033,I473755,I369169,I369177,I473764,I369194,I369220,I369228,I369036,I473776,I369268,I369027,I369018,I369304,I473767,I473761,I369321,I369347,I369355,I369372,I369021,I369403,I473773,I369420,I369437,I369030,I369468,I369015,I369499,I369516,I369024,I369571,I369597,I369605,I369622,I369639,I369665,I369696,I369704,I369721,I369747,I369755,I369795,I369831,I369848,I369874,I369882,I369899,I369930,I369947,I369964,I369995,I370026,I370043,I370098,I370124,I370132,I370149,I370166,I370192,I370223,I370231,I370248,I370274,I370282,I370322,I370358,I370375,I370401,I370409,I370426,I370457,I370474,I370491,I370522,I370553,I370570,I370625,I370651,I370659,I370676,I370693,I370719,I370750,I370758,I370775,I370801,I370809,I370849,I370885,I370902,I370928,I370936,I370953,I370984,I371001,I371018,I371049,I371080,I371097,I371152,I527490,I371178,I371186,I371203,I527472,I527475,I371220,I527487,I371246,I527496,I371277,I371285,I527481,I371302,I371328,I371336,I527493,I371376,I371412,I527484,I527478,I371429,I371455,I371463,I371480,I371511,I371528,I371545,I371576,I371607,I371624,I371679,I371705,I371713,I371730,I371747,I371773,I371668,I371804,I371812,I371829,I371855,I371863,I371671,I371903,I371662,I371653,I371939,I371956,I371982,I371990,I372007,I371656,I372038,I372055,I372072,I371665,I372103,I371650,I372134,I372151,I371659,I372206,I372232,I372240,I372257,I372274,I372300,I372331,I372339,I372356,I372382,I372390,I372430,I372466,I372483,I372509,I372517,I372534,I372565,I372582,I372599,I372630,I372661,I372678,I372733,I372759,I372767,I372784,I372801,I372827,I372858,I372866,I372883,I372909,I372917,I372957,I372993,I373010,I373036,I373044,I373061,I373092,I373109,I373126,I373157,I373188,I373205,I373260,I397714,I373286,I373294,I373311,I397729,I397711,I373328,I373354,I373249,I397720,I373385,I373393,I397738,I373410,I373436,I373444,I373252,I397735,I373484,I373243,I373234,I373520,I397732,I397723,I373537,I397717,I373563,I373571,I373588,I373237,I373619,I397726,I373636,I373653,I373246,I373684,I373231,I373715,I373732,I373240,I373787,I373813,I373821,I373838,I373855,I373881,I373912,I373920,I373937,I373963,I373971,I374011,I374047,I374064,I374090,I374098,I374115,I374146,I374163,I374180,I374211,I374242,I374259,I374314,I374340,I374348,I374365,I374382,I374408,I374439,I374447,I374464,I374490,I374498,I374538,I374574,I374591,I374617,I374625,I374642,I374673,I374690,I374707,I374738,I374769,I374786,I374841,I374867,I374875,I374892,I374909,I374935,I374966,I374974,I374991,I375017,I375025,I375065,I375101,I375118,I375144,I375152,I375169,I375200,I375217,I375234,I375265,I375296,I375313,I375368,I375394,I375402,I375419,I375436,I375462,I375493,I375501,I375518,I375544,I375552,I375592,I375628,I375645,I375671,I375679,I375696,I375727,I375744,I375761,I375792,I375823,I375840,I375895,I375921,I375929,I375946,I375963,I375989,I375884,I376020,I376028,I376045,I376071,I376079,I375887,I376119,I375878,I375869,I376155,I376172,I376198,I376206,I376223,I375872,I376254,I376271,I376288,I375881,I376319,I375866,I376350,I376367,I375875,I376428,I376454,I376471,I376479,I376496,I376513,I376530,I376547,I376564,I376595,I376612,I376643,I376660,I376677,I376708,I376748,I376756,I376773,I376790,I376807,I376838,I376855,I376872,I376898,I376920,I376937,I376968,I377013,I377074,I377100,I377117,I377125,I377142,I377159,I377176,I377193,I377210,I377060,I377241,I377258,I377063,I377289,I377306,I377323,I377039,I377354,I377051,I377394,I377402,I377419,I377436,I377453,I377066,I377484,I377501,I377518,I377544,I377054,I377566,I377583,I377048,I377614,I377042,I377045,I377659,I377057,I377720,I377746,I377763,I377771,I377788,I377805,I377822,I377839,I377856,I377706,I377887,I377904,I377709,I377935,I377952,I377969,I377685,I378000,I377697,I378040,I378048,I378065,I378082,I378099,I377712,I378130,I378147,I378164,I378190,I377700,I378212,I378229,I377694,I378260,I377688,I377691,I378305,I377703,I378366,I378392,I378409,I378417,I378434,I378451,I378468,I378485,I378502,I378533,I378550,I378581,I378598,I378615,I378646,I378686,I378694,I378711,I378728,I378745,I378776,I378793,I378810,I378836,I378858,I378875,I378906,I378951,I379012,I379038,I379055,I379063,I379080,I379097,I379114,I379131,I379148,I379179,I379196,I379227,I379244,I379261,I379292,I379332,I379340,I379357,I379374,I379391,I379422,I379439,I379456,I379482,I379504,I379521,I379552,I379597,I379658,I466256,I379684,I466238,I379701,I379709,I379726,I466247,I379743,I466259,I379760,I466241,I379777,I466250,I379794,I379644,I379825,I379842,I379647,I379873,I379890,I466262,I379907,I379623,I379938,I379635,I379978,I379986,I380003,I380020,I380037,I379650,I380068,I466244,I380085,I466253,I380102,I380128,I379638,I380150,I380167,I379632,I380198,I379626,I379629,I380243,I379641,I380304,I380330,I380347,I380355,I380372,I380389,I380406,I380423,I380440,I380471,I380488,I380519,I380536,I380553,I380584,I380624,I380632,I380649,I380666,I380683,I380714,I380731,I380748,I380774,I380796,I380813,I380844,I380889,I380950,I380976,I380993,I381001,I381018,I381035,I381052,I381069,I381086,I380936,I381117,I381134,I380939,I381165,I381182,I381199,I380915,I381230,I380927,I381270,I381278,I381295,I381312,I381329,I380942,I381360,I381377,I381394,I381420,I380930,I381442,I381459,I380924,I381490,I380918,I380921,I381535,I380933,I381596,I381622,I381639,I381647,I381664,I381681,I381698,I381715,I381732,I381763,I381780,I381811,I381828,I381845,I381876,I381916,I381924,I381941,I381958,I381975,I382006,I382023,I382040,I382066,I382088,I382105,I382136,I382181,I382242,I382268,I382285,I382293,I382310,I382327,I382344,I382361,I382378,I382409,I382426,I382457,I382474,I382491,I382522,I382562,I382570,I382587,I382604,I382621,I382652,I382669,I382686,I382712,I382734,I382751,I382782,I382827,I382888,I382914,I382931,I382939,I382956,I382973,I382990,I383007,I383024,I382874,I383055,I383072,I382877,I383103,I383120,I383137,I382853,I383168,I382865,I383208,I383216,I383233,I383250,I383267,I382880,I383298,I383315,I383332,I383358,I382868,I383380,I383397,I382862,I383428,I382856,I382859,I383473,I382871,I383534,I383560,I383577,I383585,I383602,I383619,I383636,I383653,I383670,I383701,I383718,I383749,I383766,I383783,I383814,I383854,I383862,I383879,I383896,I383913,I383944,I383961,I383978,I384004,I384026,I384043,I384074,I384119,I384180,I384206,I384223,I384231,I384248,I384265,I384282,I384299,I384316,I384347,I384364,I384395,I384412,I384429,I384460,I384500,I384508,I384525,I384542,I384559,I384590,I384607,I384624,I384650,I384672,I384689,I384720,I384765,I384826,I384852,I384869,I384877,I384894,I384911,I384928,I384945,I384962,I384993,I385010,I385041,I385058,I385075,I385106,I385146,I385154,I385171,I385188,I385205,I385236,I385253,I385270,I385296,I385318,I385335,I385366,I385411,I385472,I385498,I385515,I385523,I385540,I385557,I385574,I385591,I385608,I385458,I385639,I385656,I385461,I385687,I385704,I385721,I385437,I385752,I385449,I385792,I385800,I385817,I385834,I385851,I385464,I385882,I385899,I385916,I385942,I385452,I385964,I385981,I385446,I386012,I385440,I385443,I386057,I385455,I386118,I451228,I386144,I451210,I386161,I386169,I386186,I451219,I386203,I451231,I386220,I451213,I386237,I451222,I386254,I386285,I386302,I386333,I386350,I451234,I386367,I386398,I386438,I386446,I386463,I386480,I386497,I386528,I451216,I386545,I451225,I386562,I386588,I386610,I386627,I386658,I386703,I386764,I386790,I386807,I386815,I386832,I386849,I386866,I386883,I386900,I386750,I386931,I386948,I386753,I386979,I386996,I387013,I386729,I387044,I386741,I387084,I387092,I387109,I387126,I387143,I386756,I387174,I387191,I387208,I387234,I386744,I387256,I387273,I386738,I387304,I386732,I386735,I387349,I386747,I387410,I387436,I387453,I387461,I387478,I387495,I387512,I387529,I387546,I387577,I387594,I387625,I387642,I387659,I387690,I387730,I387738,I387755,I387772,I387789,I387820,I387837,I387854,I387880,I387902,I387919,I387950,I387995,I388056,I388082,I388099,I388107,I388124,I388141,I388158,I388175,I388192,I388223,I388240,I388271,I388288,I388305,I388336,I388376,I388384,I388401,I388418,I388435,I388466,I388483,I388500,I388526,I388548,I388565,I388596,I388641,I388702,I388728,I388745,I388753,I388770,I388787,I388804,I388821,I388838,I388688,I388869,I388886,I388691,I388917,I388934,I388951,I388667,I388982,I388679,I389022,I389030,I389047,I389064,I389081,I388694,I389112,I389129,I389146,I389172,I388682,I389194,I389211,I388676,I389242,I388670,I388673,I389287,I388685,I389348,I389374,I389391,I389399,I389416,I389433,I389450,I389467,I389484,I389334,I389515,I389532,I389337,I389563,I389580,I389597,I389313,I389628,I389325,I389668,I389676,I389693,I389710,I389727,I389340,I389758,I389775,I389792,I389818,I389328,I389840,I389857,I389322,I389888,I389316,I389319,I389933,I389331,I389994,I390020,I390037,I390045,I390062,I390079,I390096,I390113,I390130,I389980,I390161,I390178,I389983,I390209,I390226,I390243,I389959,I390274,I389971,I390314,I390322,I390339,I390356,I390373,I389986,I390404,I390421,I390438,I390464,I389974,I390486,I390503,I389968,I390534,I389962,I389965,I390579,I389977,I390640,I476082,I390666,I476064,I390683,I390691,I390708,I476073,I390725,I476085,I390742,I476067,I390759,I476076,I390776,I390626,I390807,I390824,I390629,I390855,I390872,I476088,I390889,I390605,I390920,I390617,I390960,I390968,I390985,I391002,I391019,I390632,I391050,I476070,I391067,I476079,I391084,I391110,I390620,I391132,I391149,I390614,I391180,I390608,I390611,I391225,I390623,I391286,I391312,I391329,I391337,I391354,I391371,I391388,I391405,I391422,I391453,I391470,I391501,I391518,I391535,I391566,I391606,I391614,I391631,I391648,I391665,I391696,I391713,I391730,I391756,I391778,I391795,I391826,I391871,I391932,I391958,I391975,I391983,I392000,I392017,I392034,I392051,I392068,I392099,I392116,I392147,I392164,I392181,I392212,I392252,I392260,I392277,I392294,I392311,I392342,I392359,I392376,I392402,I392424,I392441,I392472,I392517,I392578,I392604,I392621,I392629,I392646,I392663,I392680,I392697,I392714,I392745,I392762,I392793,I392810,I392827,I392858,I392898,I392906,I392923,I392940,I392957,I392988,I393005,I393022,I393048,I393070,I393087,I393118,I393163,I393224,I393250,I393267,I393275,I393292,I393309,I393326,I393343,I393360,I393391,I393408,I393439,I393456,I393473,I393504,I393544,I393552,I393569,I393586,I393603,I393634,I393651,I393668,I393694,I393716,I393733,I393764,I393809,I393870,I393896,I393913,I393921,I393938,I393955,I393972,I393989,I394006,I394037,I394054,I394085,I394102,I394119,I394150,I394190,I394198,I394215,I394232,I394249,I394280,I394297,I394314,I394340,I394362,I394379,I394410,I394455,I394516,I483596,I394542,I483578,I394559,I394567,I394584,I483587,I394601,I483599,I394618,I483581,I394635,I483590,I394652,I394683,I394700,I394731,I394748,I483602,I394765,I394796,I394836,I394844,I394861,I394878,I394895,I394926,I483584,I394943,I483593,I394960,I394986,I395008,I395025,I395056,I395101,I395162,I395188,I395205,I395213,I395230,I395247,I395264,I395281,I395298,I395329,I395346,I395377,I395394,I395411,I395442,I395482,I395490,I395507,I395524,I395541,I395572,I395589,I395606,I395632,I395654,I395671,I395702,I395747,I395808,I395834,I395851,I395859,I395876,I395893,I395910,I395927,I395944,I395975,I395992,I396023,I396040,I396057,I396088,I396128,I396136,I396153,I396170,I396187,I396218,I396235,I396252,I396278,I396300,I396317,I396348,I396393,I396454,I396480,I396497,I396505,I396522,I396539,I396556,I396573,I396590,I396440,I396621,I396638,I396443,I396669,I396686,I396703,I396419,I396734,I396431,I396774,I396782,I396799,I396816,I396833,I396446,I396864,I396881,I396898,I396924,I396434,I396946,I396963,I396428,I396994,I396422,I396425,I397039,I396437,I397100,I397126,I397143,I397151,I397168,I397185,I397202,I397219,I397236,I397267,I397284,I397315,I397332,I397349,I397380,I397420,I397428,I397445,I397462,I397479,I397510,I397527,I397544,I397570,I397592,I397609,I397640,I397685,I397746,I500936,I397772,I500918,I397789,I397797,I397814,I500927,I397831,I500939,I397848,I500921,I397865,I500930,I397882,I397913,I397930,I397961,I397978,I500942,I397995,I398026,I398066,I398074,I398091,I398108,I398125,I398156,I500924,I398173,I500933,I398190,I398216,I398238,I398255,I398286,I398331,I398392,I451806,I398418,I451788,I398435,I398443,I398460,I451797,I398477,I451809,I398494,I451791,I398511,I451800,I398528,I398559,I398576,I398607,I398624,I451812,I398641,I398672,I398712,I398720,I398737,I398754,I398771,I398802,I451794,I398819,I451803,I398836,I398862,I398884,I398901,I398932,I398977,I399038,I399064,I399081,I399089,I399106,I399123,I399140,I399157,I399174,I399205,I399222,I399253,I399270,I399287,I399318,I399358,I399366,I399383,I399400,I399417,I399448,I399465,I399482,I399508,I399530,I399547,I399578,I399623,I399684,I399710,I399727,I399735,I399752,I399769,I399786,I399803,I399820,I399670,I399851,I399868,I399673,I399899,I399916,I399933,I399649,I399964,I399661,I400004,I400012,I400029,I400046,I400063,I399676,I400094,I400111,I400128,I400154,I399664,I400176,I400193,I399658,I400224,I399652,I399655,I400269,I399667,I400330,I400356,I400373,I400381,I400398,I400415,I400432,I400449,I400466,I400497,I400514,I400545,I400562,I400579,I400610,I400650,I400658,I400675,I400692,I400709,I400740,I400757,I400774,I400800,I400822,I400839,I400870,I400915,I400976,I401002,I401019,I401027,I401044,I401061,I401078,I401095,I401112,I401143,I401160,I401191,I401208,I401225,I401256,I401296,I401304,I401321,I401338,I401355,I401386,I401403,I401420,I401446,I401468,I401485,I401516,I401561,I401622,I401648,I401665,I401673,I401690,I401707,I401724,I401741,I401758,I401789,I401806,I401837,I401854,I401871,I401902,I401942,I401950,I401967,I401984,I402001,I402032,I402049,I402066,I402092,I402114,I402131,I402162,I402207,I402268,I547260,I402294,I547284,I402311,I402319,I402336,I547266,I402353,I547275,I402370,I402387,I547281,I402404,I402435,I402452,I402483,I402500,I547278,I402517,I402548,I402588,I402596,I402613,I402630,I547272,I402647,I402678,I547263,I402695,I547287,I402712,I547269,I402738,I402760,I402777,I402808,I402853,I402914,I438783,I402940,I438786,I402957,I402965,I402982,I402999,I438795,I403016,I438804,I403033,I438792,I403050,I403081,I403098,I403129,I403146,I438798,I403163,I403194,I403234,I403242,I403259,I403276,I438789,I403293,I403324,I438801,I403341,I403358,I403384,I403406,I403423,I403454,I403499,I403560,I517868,I403586,I517874,I403603,I403611,I403628,I517871,I403645,I517850,I403662,I517853,I403679,I517859,I403696,I403727,I403744,I403775,I403792,I403809,I403840,I403880,I403888,I403905,I403922,I517862,I403939,I403970,I403987,I517856,I404004,I517865,I404030,I404052,I404069,I404100,I404145,I404206,I404232,I404249,I404257,I404274,I404291,I404308,I404325,I404342,I404373,I404390,I404421,I404438,I404455,I404486,I404526,I404534,I404551,I404568,I404585,I404616,I404633,I404650,I404676,I404698,I404715,I404746,I404791,I404852,I404878,I404895,I404903,I404920,I404937,I404954,I404971,I404988,I405019,I405036,I405067,I405084,I405101,I405132,I405172,I405180,I405197,I405214,I405231,I405262,I405279,I405296,I405322,I405344,I405361,I405392,I405437,I405498,I405524,I405541,I405549,I405566,I405583,I405600,I405617,I405634,I405665,I405682,I405713,I405730,I405747,I405778,I405818,I405826,I405843,I405860,I405877,I405908,I405925,I405942,I405968,I405990,I406007,I406038,I406083,I406144,I406170,I406187,I406195,I406212,I406229,I406246,I406263,I406280,I406311,I406328,I406359,I406376,I406393,I406424,I406464,I406472,I406489,I406506,I406523,I406554,I406571,I406588,I406614,I406636,I406653,I406684,I406729,I406790,I406816,I406833,I406841,I406858,I406875,I406892,I406909,I406926,I406776,I406957,I406974,I406779,I407005,I407022,I407039,I406755,I407070,I406767,I407110,I407118,I407135,I407152,I407169,I406782,I407200,I407217,I407234,I407260,I406770,I407282,I407299,I406764,I407330,I406758,I406761,I407375,I406773,I407436,I407462,I407479,I407487,I407504,I407521,I407538,I407555,I407572,I407603,I407620,I407651,I407668,I407685,I407716,I407756,I407764,I407781,I407798,I407815,I407846,I407863,I407880,I407906,I407928,I407945,I407976,I408021,I408082,I447759,I408108,I447762,I408125,I408133,I408150,I408167,I447771,I408184,I447780,I408201,I447768,I408218,I408249,I408266,I408297,I408314,I447774,I408331,I408362,I408402,I408410,I408427,I408444,I447765,I408461,I408492,I447777,I408509,I408526,I408552,I408574,I408591,I408622,I408667,I408728,I540715,I408754,I540739,I408771,I408779,I408796,I540721,I408813,I540730,I408830,I408847,I540736,I408864,I408895,I408912,I408943,I408960,I540733,I408977,I409008,I409048,I409056,I409073,I409090,I540727,I409107,I409138,I540718,I409155,I540742,I409172,I540724,I409198,I409220,I409237,I409268,I409313,I409374,I409400,I409417,I409425,I409442,I409459,I409476,I409493,I409510,I409360,I409541,I409558,I409363,I409589,I409606,I409623,I409339,I409654,I409351,I409694,I409702,I409719,I409736,I409753,I409366,I409784,I409801,I409818,I409844,I409354,I409866,I409883,I409348,I409914,I409342,I409345,I409959,I409357,I410020,I456430,I410046,I456412,I410063,I410071,I410088,I456421,I410105,I456433,I410122,I456415,I410139,I456424,I410156,I410187,I410204,I410235,I410252,I456436,I410269,I410300,I410340,I410348,I410365,I410382,I410399,I410430,I456418,I410447,I456427,I410464,I410490,I410512,I410529,I410560,I410605,I410666,I410692,I410709,I410717,I410734,I410751,I410768,I410785,I410802,I410833,I410850,I410881,I410898,I410915,I410946,I410986,I410994,I411011,I411028,I411045,I411076,I411093,I411110,I411136,I411158,I411175,I411206,I411251,I411312,I411338,I411355,I411363,I411380,I411397,I411414,I411431,I411448,I411479,I411496,I411527,I411544,I411561,I411592,I411632,I411640,I411657,I411674,I411691,I411722,I411739,I411756,I411782,I411804,I411821,I411852,I411897,I411958,I411984,I412001,I412009,I412026,I412043,I412060,I412077,I412094,I411944,I412125,I412142,I411947,I412173,I412190,I412207,I411923,I412238,I411935,I412278,I412286,I412303,I412320,I412337,I411950,I412368,I412385,I412402,I412428,I411938,I412450,I412467,I411932,I412498,I411926,I411929,I412543,I411941,I412604,I412630,I412647,I412655,I412672,I412689,I412706,I412723,I412740,I412771,I412788,I412819,I412836,I412853,I412884,I412924,I412932,I412949,I412966,I412983,I413014,I413031,I413048,I413074,I413096,I413113,I413144,I413189,I413250,I566300,I413276,I566324,I413293,I413301,I413318,I566306,I413335,I566315,I413352,I413369,I566321,I413386,I413417,I413434,I413465,I413482,I566318,I413499,I413530,I413570,I413578,I413595,I413612,I566312,I413629,I413660,I566303,I413677,I566327,I413694,I566309,I413720,I413742,I413759,I413790,I413835,I413896,I413922,I413939,I413947,I413964,I413981,I413998,I414015,I414032,I413882,I414063,I414080,I413885,I414111,I414128,I414145,I413861,I414176,I413873,I414216,I414224,I414241,I414258,I414275,I413888,I414306,I414323,I414340,I414366,I413876,I414388,I414405,I413870,I414436,I413864,I413867,I414481,I413879,I414542,I414568,I414585,I414593,I414610,I414627,I414644,I414661,I414678,I414709,I414726,I414757,I414774,I414791,I414822,I414862,I414870,I414887,I414904,I414921,I414952,I414969,I414986,I415012,I415034,I415051,I415082,I415127,I415188,I415214,I415231,I415239,I415256,I415273,I415290,I415307,I415324,I415355,I415372,I415403,I415420,I415437,I415468,I415508,I415516,I415533,I415550,I415567,I415598,I415615,I415632,I415658,I415680,I415697,I415728,I415773,I415834,I415860,I415877,I415885,I415902,I415919,I415936,I415953,I415970,I416001,I416018,I416049,I416066,I416083,I416114,I416154,I416162,I416179,I416196,I416213,I416244,I416261,I416278,I416304,I416326,I416343,I416374,I416419,I416480,I565705,I416506,I565729,I416523,I416531,I416548,I565711,I416565,I565720,I416582,I416599,I565726,I416616,I416466,I416647,I416664,I416469,I416695,I416712,I565723,I416729,I416445,I416760,I416457,I416800,I416808,I416825,I416842,I565717,I416859,I416472,I416890,I565708,I416907,I565732,I416924,I565714,I416950,I416460,I416972,I416989,I416454,I417020,I416448,I416451,I417065,I416463,I417126,I477238,I417152,I477220,I417169,I417177,I417194,I477229,I417211,I477241,I417228,I477223,I417245,I477232,I417262,I417293,I417310,I417341,I417358,I477244,I417375,I417406,I417446,I417454,I417471,I417488,I417505,I417536,I477226,I417553,I477235,I417570,I417596,I417618,I417635,I417666,I417711,I417772,I492266,I417798,I492248,I417815,I417823,I417840,I492257,I417857,I492269,I417874,I492251,I417891,I492260,I417908,I417758,I417939,I417956,I417761,I417987,I418004,I492272,I418021,I417737,I418052,I417749,I418092,I418100,I418117,I418134,I418151,I417764,I418182,I492254,I418199,I492263,I418216,I418242,I417752,I418264,I418281,I417746,I418312,I417740,I417743,I418357,I417755,I418418,I418444,I418461,I418469,I418486,I418503,I418520,I418537,I418554,I418585,I418602,I418633,I418650,I418667,I418698,I418738,I418746,I418763,I418780,I418797,I418828,I418845,I418862,I418888,I418910,I418927,I418958,I419003,I419064,I419090,I419107,I419115,I419132,I419149,I419166,I419183,I419200,I419231,I419248,I419279,I419296,I419313,I419344,I419384,I419392,I419409,I419426,I419443,I419474,I419491,I419508,I419534,I419556,I419573,I419604,I419649,I419710,I419736,I419753,I419761,I419778,I419795,I419812,I419829,I419846,I419696,I419877,I419894,I419699,I419925,I419942,I419959,I419675,I419990,I419687,I420030,I420038,I420055,I420072,I420089,I419702,I420120,I420137,I420154,I420180,I419690,I420202,I420219,I419684,I420250,I419678,I419681,I420295,I419693,I420356,I420382,I420399,I420407,I420424,I420441,I420458,I420475,I420492,I420523,I420540,I420571,I420588,I420605,I420636,I420676,I420684,I420701,I420718,I420735,I420766,I420783,I420800,I420826,I420848,I420865,I420896,I420941,I421002,I421028,I421045,I421053,I421070,I421087,I421104,I421121,I421138,I421169,I421186,I421217,I421234,I421251,I421282,I421322,I421330,I421347,I421364,I421381,I421412,I421429,I421446,I421472,I421494,I421511,I421542,I421587,I421648,I421674,I421691,I421699,I421716,I421733,I421750,I421767,I421784,I421815,I421832,I421863,I421880,I421897,I421928,I421968,I421976,I421993,I422010,I422027,I422058,I422075,I422092,I422118,I422140,I422157,I422188,I422233,I422294,I425319,I422320,I425322,I422337,I422345,I422362,I422379,I425331,I422396,I425340,I422413,I425328,I422430,I422461,I422478,I422509,I422526,I425334,I422543,I422574,I422614,I422622,I422639,I422656,I425325,I422673,I422704,I425337,I422721,I422738,I422764,I422786,I422803,I422834,I422879,I422940,I479550,I422966,I479532,I422983,I422991,I423008,I479541,I423025,I479553,I423042,I479535,I423059,I479544,I423076,I422926,I423107,I423124,I422929,I423155,I423172,I479556,I423189,I422905,I423220,I422917,I423260,I423268,I423285,I423302,I423319,I422932,I423350,I479538,I423367,I479547,I423384,I423410,I422920,I423432,I423449,I422914,I423480,I422908,I422911,I423525,I422923,I423586,I423612,I423629,I423637,I423654,I423671,I423688,I423705,I423722,I423753,I423770,I423801,I423818,I423835,I423866,I423906,I423914,I423931,I423948,I423965,I423996,I424013,I424030,I424056,I424078,I424095,I424126,I424171,I424226,I424252,I424269,I424291,I424317,I424325,I424342,I424359,I424376,I424393,I424410,I424427,I424458,I424489,I424506,I424523,I424540,I424571,I424616,I424633,I424650,I424676,I424684,I424715,I424732,I424787,I529787,I424813,I424830,I424779,I424852,I529784,I424878,I424886,I529790,I424903,I424920,I529799,I424937,I529793,I424954,I424971,I529805,I424988,I424761,I425019,I424764,I425050,I529802,I425067,I425084,I425101,I424773,I425132,I424776,I424770,I425177,I529796,I425194,I529808,I425211,I425237,I425245,I424758,I425276,I425293,I424767,I425348,I559770,I425374,I425391,I425413,I559764,I425439,I425447,I559755,I425464,I425481,I559782,I425498,I559767,I559776,I425515,I425532,I559761,I425549,I425580,I425611,I559779,I425628,I425645,I425662,I425693,I425738,I559773,I425755,I425772,I559758,I425798,I425806,I425837,I425854,I425909,I425935,I425952,I425974,I426000,I426008,I426025,I426042,I426059,I426076,I426093,I426110,I426141,I426172,I426189,I426206,I426223,I426254,I426299,I426316,I426333,I426359,I426367,I426398,I426415,I426470,I426496,I426513,I426462,I426535,I426561,I426569,I426586,I426603,I426620,I426637,I426654,I426671,I426444,I426702,I426447,I426733,I426750,I426767,I426784,I426456,I426815,I426459,I426453,I426860,I426877,I426894,I426920,I426928,I426441,I426959,I426976,I426450,I427031,I427057,I427074,I427096,I427122,I427130,I427147,I427164,I427181,I427198,I427215,I427232,I427263,I427294,I427311,I427328,I427345,I427376,I427421,I427438,I427455,I427481,I427489,I427520,I427537,I427592,I427618,I427635,I427584,I427657,I427683,I427691,I427708,I427725,I427742,I427759,I427776,I427793,I427566,I427824,I427569,I427855,I427872,I427889,I427906,I427578,I427937,I427581,I427575,I427982,I427999,I428016,I428042,I428050,I427563,I428081,I428098,I427572,I428153,I428179,I428196,I428145,I428218,I428244,I428252,I428269,I428286,I428303,I428320,I428337,I428354,I428127,I428385,I428130,I428416,I428433,I428450,I428467,I428139,I428498,I428142,I428136,I428543,I428560,I428577,I428603,I428611,I428124,I428642,I428659,I428133,I428714,I428740,I428757,I428779,I428805,I428813,I428830,I428847,I428864,I428881,I428898,I428915,I428946,I428977,I428994,I429011,I429028,I429059,I429104,I429121,I429138,I429164,I429172,I429203,I429220,I429275,I559175,I429301,I429318,I429340,I559169,I429366,I429374,I559160,I429391,I429408,I559187,I429425,I559172,I559181,I429442,I429459,I559166,I429476,I429507,I429538,I559184,I429555,I429572,I429589,I429620,I429665,I559178,I429682,I429699,I559163,I429725,I429733,I429764,I429781,I429836,I429862,I429879,I429828,I429901,I429927,I429935,I429952,I429969,I429986,I430003,I430020,I430037,I429810,I430068,I429813,I430099,I430116,I430133,I430150,I429822,I430181,I429825,I429819,I430226,I430243,I430260,I430286,I430294,I429807,I430325,I430342,I429816,I430397,I430423,I430440,I430462,I430488,I430496,I430513,I430530,I430547,I430564,I430581,I430598,I430629,I430660,I430677,I430694,I430711,I430742,I430787,I430804,I430821,I430847,I430855,I430886,I430903,I430958,I560960,I430984,I431001,I431023,I560954,I431049,I431057,I560945,I431074,I431091,I560972,I431108,I560957,I560966,I431125,I431142,I560951,I431159,I431190,I431221,I560969,I431238,I431255,I431272,I431303,I431348,I560963,I431365,I431382,I560948,I431408,I431416,I431447,I431464,I431519,I431545,I431562,I431511,I431584,I431610,I431618,I431635,I431652,I431669,I431686,I431703,I431720,I431493,I431751,I431496,I431782,I431799,I431816,I431833,I431505,I431864,I431508,I431502,I431909,I431926,I431943,I431969,I431977,I431490,I432008,I432025,I431499,I432080,I432106,I432123,I432145,I432171,I432179,I432196,I432213,I432230,I432247,I432264,I432281,I432312,I432343,I432360,I432377,I432394,I432425,I432470,I432487,I432504,I432530,I432538,I432569,I432586,I432641,I432667,I432684,I432706,I432732,I432740,I432757,I432774,I432791,I432808,I432825,I432842,I432873,I432904,I432921,I432938,I432955,I432986,I433031,I433048,I433065,I433091,I433099,I433130,I433147,I433202,I512960,I433228,I433245,I433267,I512966,I433293,I433301,I512975,I433318,I433335,I512954,I433352,I512957,I433369,I433386,I512969,I433403,I433434,I433465,I512963,I433482,I433499,I433516,I433547,I433592,I512978,I433609,I433626,I512972,I433652,I433660,I433691,I433708,I433763,I463941,I433789,I433806,I433828,I463932,I433854,I433862,I463929,I433879,I433896,I463938,I433913,I463947,I433930,I433947,I463926,I433964,I433995,I434026,I463935,I434043,I434060,I434077,I434108,I434153,I463950,I434170,I434187,I463944,I434213,I434221,I434252,I434269,I434324,I496887,I434350,I434367,I434389,I496878,I434415,I434423,I496875,I434440,I434457,I496884,I434474,I496893,I434491,I434508,I496872,I434525,I434556,I434587,I496881,I434604,I434621,I434638,I434669,I434714,I496896,I434731,I434748,I496890,I434774,I434782,I434813,I434830,I434885,I525741,I434911,I434928,I434950,I525738,I434976,I434984,I525744,I435001,I435018,I525753,I435035,I525747,I435052,I435069,I525759,I435086,I435117,I435148,I525756,I435165,I435182,I435199,I435230,I435275,I525750,I435292,I525762,I435309,I435335,I435343,I435374,I435391,I435446,I473189,I435472,I435489,I435511,I473180,I435537,I435545,I473177,I435562,I435579,I473186,I435596,I473195,I435613,I435630,I473174,I435647,I435678,I435709,I473183,I435726,I435743,I435760,I435791,I435836,I473198,I435853,I435870,I473192,I435896,I435904,I435935,I435952,I436007,I436033,I436050,I436072,I436098,I436106,I436123,I436140,I436157,I436174,I436191,I436208,I436239,I436270,I436287,I436304,I436321,I436352,I436397,I436414,I436431,I436457,I436465,I436496,I436513,I436568,I436594,I436611,I436633,I436659,I436667,I436684,I436701,I436718,I436735,I436752,I436769,I436800,I436831,I436848,I436865,I436882,I436913,I436958,I436975,I436992,I437018,I437026,I437057,I437074,I437129,I493419,I437155,I437172,I437194,I493410,I437220,I437228,I493407,I437245,I437262,I493416,I437279,I493425,I437296,I437313,I493404,I437330,I437361,I437392,I493413,I437409,I437426,I437443,I437474,I437519,I493428,I437536,I437553,I493422,I437579,I437587,I437618,I437635,I437690,I437716,I437733,I437755,I437781,I437789,I437806,I437823,I437840,I437857,I437874,I437891,I437922,I437953,I437970,I437987,I438004,I438035,I438080,I438097,I438114,I438140,I438148,I438179,I438196,I438251,I462785,I438277,I438294,I438243,I438316,I462776,I438342,I438350,I462773,I438367,I438384,I462782,I438401,I462791,I438418,I438435,I462770,I438452,I438225,I438483,I438228,I438514,I462779,I438531,I438548,I438565,I438237,I438596,I438240,I438234,I438641,I462794,I438658,I438675,I462788,I438701,I438709,I438222,I438740,I438757,I438231,I438812,I438838,I438855,I438877,I438903,I438911,I438928,I438945,I438962,I438979,I438996,I439013,I439044,I439075,I439092,I439109,I439126,I439157,I439202,I439219,I439236,I439262,I439270,I439301,I439318,I439373,I439399,I439416,I439438,I439464,I439472,I439489,I439506,I439523,I439540,I439557,I439574,I439605,I439636,I439653,I439670,I439687,I439718,I439763,I439780,I439797,I439823,I439831,I439862,I439879,I439934,I439960,I439977,I439999,I440025,I440033,I440050,I440067,I440084,I440101,I440118,I440135,I440166,I440197,I440214,I440231,I440248,I440279,I440324,I440341,I440358,I440384,I440392,I440423,I440440,I440495,I440521,I440538,I440560,I440586,I440594,I440611,I440628,I440645,I440662,I440679,I440696,I440727,I440758,I440775,I440792,I440809,I440840,I440885,I440902,I440919,I440945,I440953,I440984,I441001,I441056,I441082,I441099,I441121,I441147,I441155,I441172,I441189,I441206,I441223,I441240,I441257,I441288,I441319,I441336,I441353,I441370,I441401,I441446,I441463,I441480,I441506,I441514,I441545,I441562,I441617,I441643,I441660,I441682,I441708,I441716,I441733,I441750,I441767,I441784,I441801,I441818,I441849,I441880,I441897,I441914,I441931,I441962,I442007,I442024,I442041,I442067,I442075,I442106,I442123,I442178,I524585,I442204,I442221,I442243,I524582,I442269,I442277,I524588,I442294,I442311,I524597,I442328,I524591,I442345,I442362,I524603,I442379,I442410,I442441,I524600,I442458,I442475,I442492,I442523,I442568,I524594,I442585,I524606,I442602,I442628,I442636,I442667,I442684,I442739,I442765,I442782,I442731,I442804,I442830,I442838,I442855,I442872,I442889,I442906,I442923,I442940,I442713,I442971,I442716,I443002,I443019,I443036,I443053,I442725,I443084,I442728,I442722,I443129,I443146,I443163,I443189,I443197,I442710,I443228,I443245,I442719,I443300,I443326,I443343,I443365,I443391,I443399,I443416,I443433,I443450,I443467,I443484,I443501,I443532,I443563,I443580,I443597,I443614,I443645,I443690,I443707,I443724,I443750,I443758,I443789,I443806,I443861,I443887,I443904,I443926,I443952,I443960,I443977,I443994,I444011,I444028,I444045,I444062,I444093,I444124,I444141,I444158,I444175,I444206,I444251,I444268,I444285,I444311,I444319,I444350,I444367,I444422,I444448,I444465,I444487,I444513,I444521,I444538,I444555,I444572,I444589,I444606,I444623,I444654,I444685,I444702,I444719,I444736,I444767,I444812,I444829,I444846,I444872,I444880,I444911,I444928,I444983,I553225,I445009,I445026,I445048,I553219,I445074,I445082,I553210,I445099,I445116,I553237,I445133,I553222,I553231,I445150,I445167,I553216,I445184,I445215,I445246,I553234,I445263,I445280,I445297,I445328,I445373,I553228,I445390,I445407,I553213,I445433,I445441,I445472,I445489,I445544,I445570,I445587,I445609,I445635,I445643,I445660,I445677,I445694,I445711,I445728,I445745,I445776,I445807,I445824,I445841,I445858,I445889,I445934,I445951,I445968,I445994,I446002,I446033,I446050,I446105,I541920,I446131,I446148,I446170,I541914,I446196,I446204,I541905,I446221,I446238,I541932,I446255,I541917,I541926,I446272,I446289,I541911,I446306,I446337,I446368,I541929,I446385,I446402,I446419,I446450,I446495,I541923,I446512,I446529,I541908,I446555,I446563,I446594,I446611,I446666,I446692,I446709,I446658,I446731,I446757,I446765,I446782,I446799,I446816,I446833,I446850,I446867,I446640,I446898,I446643,I446929,I446946,I446963,I446980,I446652,I447011,I446655,I446649,I447056,I447073,I447090,I447116,I447124,I446637,I447155,I447172,I446646,I447227,I546085,I447253,I447270,I447292,I546079,I447318,I447326,I546070,I447343,I447360,I546097,I447377,I546082,I546091,I447394,I447411,I546076,I447428,I447459,I447490,I546094,I447507,I447524,I447541,I447572,I447617,I546088,I447634,I447651,I546073,I447677,I447685,I447716,I447733,I447788,I447814,I447831,I447853,I447879,I447887,I447904,I447921,I447938,I447955,I447972,I447989,I448020,I448051,I448068,I448085,I448102,I448133,I448178,I448195,I448212,I448238,I448246,I448277,I448294,I448352,I448378,I448386,I448335,I448426,I448434,I448451,I448468,I448323,I448508,I448344,I448530,I448547,I448573,I448581,I448598,I448615,I448632,I448649,I448320,I448341,I448694,I448332,I448725,I448742,I448768,I448776,I448338,I448807,I448824,I448841,I448858,I448329,I448326,I448930,I448956,I448964,I449004,I449012,I449029,I449046,I449086,I449108,I449125,I449151,I449159,I449176,I449193,I449210,I449227,I449272,I449303,I449320,I449346,I449354,I449385,I449402,I449419,I449436,I449508,I449534,I449542,I449491,I449582,I449590,I449607,I449624,I449479,I449664,I449500,I449686,I449703,I449729,I449737,I449754,I449771,I449788,I449805,I449476,I449497,I449850,I449488,I449881,I449898,I449924,I449932,I449494,I449963,I449980,I449997,I450014,I449485,I449482,I450086,I450112,I450120,I450160,I450168,I450185,I450202,I450242,I450264,I450281,I450307,I450315,I450332,I450349,I450366,I450383,I450428,I450459,I450476,I450502,I450510,I450541,I450558,I450575,I450592,I450664,I450690,I450698,I450738,I450746,I450763,I450780,I450820,I450842,I450859,I450885,I450893,I450910,I450927,I450944,I450961,I451006,I451037,I451054,I451080,I451088,I451119,I451136,I451153,I451170,I451242,I451268,I451276,I451316,I451324,I451341,I451358,I451398,I451420,I451437,I451463,I451471,I451488,I451505,I451522,I451539,I451584,I451615,I451632,I451658,I451666,I451697,I451714,I451731,I451748,I451820,I451846,I451854,I451894,I451902,I451919,I451936,I451976,I451998,I452015,I452041,I452049,I452066,I452083,I452100,I452117,I452162,I452193,I452210,I452236,I452244,I452275,I452292,I452309,I452326,I452398,I452424,I452432,I452472,I452480,I452497,I452514,I452554,I452576,I452593,I452619,I452627,I452644,I452661,I452678,I452695,I452740,I452771,I452788,I452814,I452822,I452853,I452870,I452887,I452904,I452976,I453002,I453010,I453050,I453058,I453075,I453092,I453132,I453154,I453171,I453197,I453205,I453222,I453239,I453256,I453273,I453318,I453349,I453366,I453392,I453400,I453431,I453448,I453465,I453482,I453554,I453580,I453588,I453628,I453636,I453653,I453670,I453710,I453732,I453749,I453775,I453783,I453800,I453817,I453834,I453851,I453896,I453927,I453944,I453970,I453978,I454009,I454026,I454043,I454060,I454132,I454158,I454166,I454206,I454214,I454231,I454248,I454288,I454310,I454327,I454353,I454361,I454378,I454395,I454412,I454429,I454474,I454505,I454522,I454548,I454556,I454587,I454604,I454621,I454638,I454710,I552642,I454736,I454744,I552624,I552615,I454784,I454792,I552630,I454809,I552618,I454826,I454866,I454888,I552627,I454905,I454931,I454939,I454956,I552636,I454973,I454990,I455007,I455052,I552639,I455083,I455100,I552633,I552621,I455126,I455134,I455165,I455182,I455199,I455216,I455288,I455314,I455322,I455362,I455370,I455387,I455404,I455444,I455466,I455483,I455509,I455517,I455534,I455551,I455568,I455585,I455630,I455661,I455678,I455704,I455712,I455743,I455760,I455777,I455794,I455866,I455892,I455900,I455940,I455948,I455965,I455982,I456022,I456044,I456061,I456087,I456095,I456112,I456129,I456146,I456163,I456208,I456239,I456256,I456282,I456290,I456321,I456338,I456355,I456372,I456444,I456470,I456478,I456518,I456526,I456543,I456560,I456600,I456622,I456639,I456665,I456673,I456690,I456707,I456724,I456741,I456786,I456817,I456834,I456860,I456868,I456899,I456916,I456933,I456950,I457022,I457048,I457056,I457096,I457104,I457121,I457138,I457178,I457200,I457217,I457243,I457251,I457268,I457285,I457302,I457319,I457364,I457395,I457412,I457438,I457446,I457477,I457494,I457511,I457528,I457600,I457626,I457634,I457583,I457674,I457682,I457699,I457716,I457571,I457756,I457592,I457778,I457795,I457821,I457829,I457846,I457863,I457880,I457897,I457568,I457589,I457942,I457580,I457973,I457990,I458016,I458024,I457586,I458055,I458072,I458089,I458106,I457577,I457574,I458178,I556807,I458204,I458212,I556789,I556780,I458252,I458260,I556795,I458277,I556783,I458294,I458334,I458356,I556792,I458373,I458399,I458407,I458424,I556801,I458441,I458458,I458475,I458520,I556804,I458551,I458568,I556798,I556786,I458594,I458602,I458633,I458650,I458667,I458684,I458756,I458782,I458790,I458830,I458838,I458855,I458872,I458912,I458934,I458951,I458977,I458985,I459002,I459019,I459036,I459053,I459098,I459129,I459146,I459172,I459180,I459211,I459228,I459245,I459262,I459334,I459360,I459368,I459408,I459416,I459433,I459450,I459490,I459512,I459529,I459555,I459563,I459580,I459597,I459614,I459631,I459676,I459707,I459724,I459750,I459758,I459789,I459806,I459823,I459840,I459912,I459938,I459946,I459986,I459994,I460011,I460028,I460068,I460090,I460107,I460133,I460141,I460158,I460175,I460192,I460209,I460254,I460285,I460302,I460328,I460336,I460367,I460384,I460401,I460418,I460490,I460516,I460524,I460564,I460572,I460589,I460606,I460646,I460668,I460685,I460711,I460719,I460736,I460753,I460770,I460787,I460832,I460863,I460880,I460906,I460914,I460945,I460962,I460979,I460996,I461068,I461094,I461102,I461142,I461150,I461167,I461184,I461224,I461246,I461263,I461289,I461297,I461314,I461331,I461348,I461365,I461410,I461441,I461458,I461484,I461492,I461523,I461540,I461557,I461574,I461646,I461672,I461680,I461720,I461728,I461745,I461762,I461802,I461824,I461841,I461867,I461875,I461892,I461909,I461926,I461943,I461988,I462019,I462036,I462062,I462070,I462101,I462118,I462135,I462152,I462224,I462250,I462258,I462298,I462306,I462323,I462340,I462380,I462402,I462419,I462445,I462453,I462470,I462487,I462504,I462521,I462566,I462597,I462614,I462640,I462648,I462679,I462696,I462713,I462730,I462802,I519503,I462828,I462836,I519497,I519482,I462876,I462884,I519488,I462901,I519500,I462918,I462958,I462980,I462997,I463023,I463031,I463048,I519506,I463065,I519494,I463082,I463099,I463144,I519485,I463175,I463192,I519491,I463218,I463226,I463257,I463274,I463291,I463308,I463380,I463406,I463414,I463454,I463462,I463479,I463496,I463536,I463558,I463575,I463601,I463609,I463626,I463643,I463660,I463677,I463722,I463753,I463770,I463796,I463804,I463835,I463852,I463869,I463886,I463958,I463984,I463992,I464032,I464040,I464057,I464074,I464114,I464136,I464153,I464179,I464187,I464204,I464221,I464238,I464255,I464300,I464331,I464348,I464374,I464382,I464413,I464430,I464447,I464464,I464536,I464562,I464570,I464610,I464618,I464635,I464652,I464692,I464714,I464731,I464757,I464765,I464782,I464799,I464816,I464833,I464878,I464909,I464926,I464952,I464960,I464991,I465008,I465025,I465042,I465114,I465140,I465148,I465188,I465196,I465213,I465230,I465270,I465292,I465309,I465335,I465343,I465360,I465377,I465394,I465411,I465456,I465487,I465504,I465530,I465538,I465569,I465586,I465603,I465620,I465692,I465718,I465726,I465675,I465766,I465774,I465791,I465808,I465663,I465848,I465684,I465870,I465887,I465913,I465921,I465938,I465955,I465972,I465989,I465660,I465681,I466034,I465672,I466065,I466082,I466108,I466116,I465678,I466147,I466164,I466181,I466198,I465669,I465666,I466270,I549072,I466296,I466304,I549054,I549045,I466344,I466352,I549060,I466369,I549048,I466386,I466426,I466448,I549057,I466465,I466491,I466499,I466516,I549066,I466533,I466550,I466567,I466612,I549069,I466643,I466660,I549063,I549051,I466686,I466694,I466725,I466742,I466759,I466776,I466848,I466874,I466882,I466922,I466930,I466947,I466964,I467004,I467026,I467043,I467069,I467077,I467094,I467111,I467128,I467145,I467190,I467221,I467238,I467264,I467272,I467303,I467320,I467337,I467354,I467426,I518959,I467452,I467460,I518953,I518938,I467500,I467508,I518944,I467525,I518956,I467542,I467582,I467604,I467621,I467647,I467655,I467672,I518962,I467689,I518950,I467706,I467723,I467768,I518941,I467799,I467816,I518947,I467842,I467850,I467881,I467898,I467915,I467932,I468004,I468030,I468038,I468078,I468086,I468103,I468120,I468160,I468182,I468199,I468225,I468233,I468250,I468267,I468284,I468301,I468346,I468377,I468394,I468420,I468428,I468459,I468476,I468493,I468510,I468582,I468608,I468616,I468656,I468664,I468681,I468698,I468738,I468760,I468777,I468803,I468811,I468828,I468845,I468862,I468879,I468924,I468955,I468972,I468998,I469006,I469037,I469054,I469071,I469088,I469160,I469186,I469194,I469234,I469242,I469259,I469276,I469316,I469338,I469355,I469381,I469389,I469406,I469423,I469440,I469457,I469502,I469533,I469550,I469576,I469584,I469615,I469632,I469649,I469666,I469738,I469764,I469772,I469812,I469820,I469837,I469854,I469894,I469916,I469933,I469959,I469967,I469984,I470001,I470018,I470035,I470080,I470111,I470128,I470154,I470162,I470193,I470210,I470227,I470244,I470316,I470342,I470350,I470390,I470398,I470415,I470432,I470472,I470494,I470511,I470537,I470545,I470562,I470579,I470596,I470613,I470658,I470689,I470706,I470732,I470740,I470771,I470788,I470805,I470822,I470894,I545502,I470920,I470928,I545484,I470877,I545475,I470968,I470976,I545490,I470993,I545478,I471010,I470865,I471050,I470886,I471072,I545487,I471089,I471115,I471123,I471140,I545496,I471157,I471174,I471191,I470862,I470883,I471236,I545499,I470874,I471267,I471284,I545493,I545481,I471310,I471318,I470880,I471349,I471366,I471383,I471400,I470871,I470868,I471472,I471498,I471506,I471455,I471546,I471554,I471571,I471588,I471443,I471628,I471464,I471650,I471667,I471693,I471701,I471718,I471735,I471752,I471769,I471440,I471461,I471814,I471452,I471845,I471862,I471888,I471896,I471458,I471927,I471944,I471961,I471978,I471449,I471446,I472050,I472076,I472084,I472033,I472124,I472132,I472149,I472166,I472021,I472206,I472042,I472228,I472245,I472271,I472279,I472296,I472313,I472330,I472347,I472018,I472039,I472392,I472030,I472423,I472440,I472466,I472474,I472036,I472505,I472522,I472539,I472556,I472027,I472024,I472628,I472654,I472662,I472611,I472702,I472710,I472727,I472744,I472599,I472784,I472620,I472806,I472823,I472849,I472857,I472874,I472891,I472908,I472925,I472596,I472617,I472970,I472608,I473001,I473018,I473044,I473052,I472614,I473083,I473100,I473117,I473134,I472605,I472602,I473206,I473232,I473240,I473280,I473288,I473305,I473322,I473362,I473384,I473401,I473427,I473435,I473452,I473469,I473486,I473503,I473548,I473579,I473596,I473622,I473630,I473661,I473678,I473695,I473712,I473784,I473810,I473818,I473858,I473866,I473883,I473900,I473940,I473962,I473979,I474005,I474013,I474030,I474047,I474064,I474081,I474126,I474157,I474174,I474200,I474208,I474239,I474256,I474273,I474290,I474362,I474388,I474396,I474436,I474444,I474461,I474478,I474518,I474540,I474557,I474583,I474591,I474608,I474625,I474642,I474659,I474704,I474735,I474752,I474778,I474786,I474817,I474834,I474851,I474868,I474940,I474966,I474974,I475014,I475022,I475039,I475056,I475096,I475118,I475135,I475161,I475169,I475186,I475203,I475220,I475237,I475282,I475313,I475330,I475356,I475364,I475395,I475412,I475429,I475446,I475518,I475544,I475552,I475592,I475600,I475617,I475634,I475674,I475696,I475713,I475739,I475747,I475764,I475781,I475798,I475815,I475860,I475891,I475908,I475934,I475942,I475973,I475990,I476007,I476024,I476096,I476122,I476130,I476170,I476178,I476195,I476212,I476252,I476274,I476291,I476317,I476325,I476342,I476359,I476376,I476393,I476438,I476469,I476486,I476512,I476520,I476551,I476568,I476585,I476602,I476674,I476700,I476708,I476657,I476748,I476756,I476773,I476790,I476645,I476830,I476666,I476852,I476869,I476895,I476903,I476920,I476937,I476954,I476971,I476642,I476663,I477016,I476654,I477047,I477064,I477090,I477098,I476660,I477129,I477146,I477163,I477180,I476651,I476648,I477252,I477278,I477286,I477326,I477334,I477351,I477368,I477408,I477430,I477447,I477473,I477481,I477498,I477515,I477532,I477549,I477594,I477625,I477642,I477668,I477676,I477707,I477724,I477741,I477758,I477830,I477856,I477864,I477904,I477912,I477929,I477946,I477986,I478008,I478025,I478051,I478059,I478076,I478093,I478110,I478127,I478172,I478203,I478220,I478246,I478254,I478285,I478302,I478319,I478336,I478408,I478434,I478442,I478391,I478482,I478490,I478507,I478524,I478379,I478564,I478400,I478586,I478603,I478629,I478637,I478654,I478671,I478688,I478705,I478376,I478397,I478750,I478388,I478781,I478798,I478824,I478832,I478394,I478863,I478880,I478897,I478914,I478385,I478382,I478986,I479012,I479020,I479060,I479068,I479085,I479102,I479142,I479164,I479181,I479207,I479215,I479232,I479249,I479266,I479283,I479328,I479359,I479376,I479402,I479410,I479441,I479458,I479475,I479492,I479564,I479590,I479598,I479638,I479646,I479663,I479680,I479720,I479742,I479759,I479785,I479793,I479810,I479827,I479844,I479861,I479906,I479937,I479954,I479980,I479988,I480019,I480036,I480053,I480070,I480142,I480168,I480176,I480216,I480224,I480241,I480258,I480298,I480320,I480337,I480363,I480371,I480388,I480405,I480422,I480439,I480484,I480515,I480532,I480558,I480566,I480597,I480614,I480631,I480648,I480720,I480746,I480754,I480703,I480794,I480802,I480819,I480836,I480691,I480876,I480712,I480898,I480915,I480941,I480949,I480966,I480983,I481000,I481017,I480688,I480709,I481062,I480700,I481093,I481110,I481136,I481144,I480706,I481175,I481192,I481209,I481226,I480697,I480694,I481298,I481324,I481332,I481372,I481380,I481397,I481414,I481454,I481476,I481493,I481519,I481527,I481544,I481561,I481578,I481595,I481640,I481671,I481688,I481714,I481722,I481753,I481770,I481787,I481804,I481876,I481902,I481910,I481950,I481958,I481975,I481992,I482032,I482054,I482071,I482097,I482105,I482122,I482139,I482156,I482173,I482218,I482249,I482266,I482292,I482300,I482331,I482348,I482365,I482382,I482454,I482480,I482488,I482528,I482536,I482553,I482570,I482610,I482632,I482649,I482675,I482683,I482700,I482717,I482734,I482751,I482796,I482827,I482844,I482870,I482878,I482909,I482926,I482943,I482960,I483032,I540147,I483058,I483066,I540129,I540120,I483106,I483114,I540135,I483131,I540123,I483148,I483188,I483210,I540132,I483227,I483253,I483261,I483278,I540141,I483295,I483312,I483329,I483374,I540144,I483405,I483422,I540138,I540126,I483448,I483456,I483487,I483504,I483521,I483538,I483610,I483636,I483644,I483684,I483692,I483709,I483726,I483766,I483788,I483805,I483831,I483839,I483856,I483873,I483890,I483907,I483952,I483983,I484000,I484026,I484034,I484065,I484082,I484099,I484116,I484188,I484214,I484222,I484262,I484270,I484287,I484304,I484344,I484366,I484383,I484409,I484417,I484434,I484451,I484468,I484485,I484530,I484561,I484578,I484604,I484612,I484643,I484660,I484677,I484694,I484766,I484792,I484800,I484840,I484848,I484865,I484882,I484922,I484944,I484961,I484987,I484995,I485012,I485029,I485046,I485063,I485108,I485139,I485156,I485182,I485190,I485221,I485238,I485255,I485272,I485344,I485370,I485378,I485418,I485426,I485443,I485460,I485500,I485522,I485539,I485565,I485573,I485590,I485607,I485624,I485641,I485686,I485717,I485734,I485760,I485768,I485799,I485816,I485833,I485850,I485922,I485948,I485956,I485996,I486004,I486021,I486038,I486078,I486100,I486117,I486143,I486151,I486168,I486185,I486202,I486219,I486264,I486295,I486312,I486338,I486346,I486377,I486394,I486411,I486428,I486500,I486526,I486534,I486574,I486582,I486599,I486616,I486656,I486678,I486695,I486721,I486729,I486746,I486763,I486780,I486797,I486842,I486873,I486890,I486916,I486924,I486955,I486972,I486989,I487006,I487078,I487104,I487112,I487152,I487160,I487177,I487194,I487234,I487256,I487273,I487299,I487307,I487324,I487341,I487358,I487375,I487420,I487451,I487468,I487494,I487502,I487533,I487550,I487567,I487584,I487656,I487682,I487690,I487730,I487738,I487755,I487772,I487812,I487834,I487851,I487877,I487885,I487902,I487919,I487936,I487953,I487998,I488029,I488046,I488072,I488080,I488111,I488128,I488145,I488162,I488234,I488260,I488268,I488308,I488316,I488333,I488350,I488390,I488412,I488429,I488455,I488463,I488480,I488497,I488514,I488531,I488576,I488607,I488624,I488650,I488658,I488689,I488706,I488723,I488740,I488812,I488838,I488846,I488886,I488894,I488911,I488928,I488968,I488990,I489007,I489033,I489041,I489058,I489075,I489092,I489109,I489154,I489185,I489202,I489228,I489236,I489267,I489284,I489301,I489318,I489390,I489416,I489424,I489464,I489472,I489489,I489506,I489546,I489568,I489585,I489611,I489619,I489636,I489653,I489670,I489687,I489732,I489763,I489780,I489806,I489814,I489845,I489862,I489879,I489896,I489968,I489994,I490002,I490042,I490050,I490067,I490084,I490124,I490146,I490163,I490189,I490197,I490214,I490231,I490248,I490265,I490310,I490341,I490358,I490384,I490392,I490423,I490440,I490457,I490474,I490546,I490572,I490580,I490620,I490628,I490645,I490662,I490702,I490724,I490741,I490767,I490775,I490792,I490809,I490826,I490843,I490888,I490919,I490936,I490962,I490970,I491001,I491018,I491035,I491052,I491124,I526918,I491150,I491158,I526900,I526909,I491198,I491206,I526894,I491223,I526906,I491240,I491280,I491302,I526897,I491319,I491345,I491353,I491370,I491387,I491404,I491421,I491466,I526915,I491497,I491514,I526903,I526912,I491540,I491548,I491579,I491596,I491613,I491630,I491702,I491728,I491736,I491776,I491784,I491801,I491818,I491858,I491880,I491897,I491923,I491931,I491948,I491965,I491982,I491999,I492044,I492075,I492092,I492118,I492126,I492157,I492174,I492191,I492208,I492280,I492306,I492314,I492354,I492362,I492379,I492396,I492436,I492458,I492475,I492501,I492509,I492526,I492543,I492560,I492577,I492622,I492653,I492670,I492696,I492704,I492735,I492752,I492769,I492786,I492858,I492884,I492892,I492932,I492940,I492957,I492974,I493014,I493036,I493053,I493079,I493087,I493104,I493121,I493138,I493155,I493200,I493231,I493248,I493274,I493282,I493313,I493330,I493347,I493364,I493436,I493462,I493470,I493510,I493518,I493535,I493552,I493592,I493614,I493631,I493657,I493665,I493682,I493699,I493716,I493733,I493778,I493809,I493826,I493852,I493860,I493891,I493908,I493925,I493942,I494014,I494040,I494048,I494088,I494096,I494113,I494130,I494170,I494192,I494209,I494235,I494243,I494260,I494277,I494294,I494311,I494356,I494387,I494404,I494430,I494438,I494469,I494486,I494503,I494520,I494592,I494618,I494626,I494575,I494666,I494674,I494691,I494708,I494563,I494748,I494584,I494770,I494787,I494813,I494821,I494838,I494855,I494872,I494889,I494560,I494581,I494934,I494572,I494965,I494982,I495008,I495016,I494578,I495047,I495064,I495081,I495098,I494569,I494566,I495170,I495196,I495204,I495244,I495252,I495269,I495286,I495326,I495348,I495365,I495391,I495399,I495416,I495433,I495450,I495467,I495512,I495543,I495560,I495586,I495594,I495625,I495642,I495659,I495676,I495748,I495774,I495782,I495822,I495830,I495847,I495864,I495904,I495926,I495943,I495969,I495977,I495994,I496011,I496028,I496045,I496090,I496121,I496138,I496164,I496172,I496203,I496220,I496237,I496254,I496326,I496352,I496360,I496400,I496408,I496425,I496442,I496482,I496504,I496521,I496547,I496555,I496572,I496589,I496606,I496623,I496668,I496699,I496716,I496742,I496750,I496781,I496798,I496815,I496832,I496904,I496930,I496938,I496978,I496986,I497003,I497020,I497060,I497082,I497099,I497125,I497133,I497150,I497167,I497184,I497201,I497246,I497277,I497294,I497320,I497328,I497359,I497376,I497393,I497410,I497482,I497508,I497516,I497556,I497564,I497581,I497598,I497638,I497660,I497677,I497703,I497711,I497728,I497745,I497762,I497779,I497824,I497855,I497872,I497898,I497906,I497937,I497954,I497971,I497988,I498060,I498086,I498094,I498043,I498134,I498142,I498159,I498176,I498031,I498216,I498052,I498238,I498255,I498281,I498289,I498306,I498323,I498340,I498357,I498028,I498049,I498402,I498040,I498433,I498450,I498476,I498484,I498046,I498515,I498532,I498549,I498566,I498037,I498034,I498638,I498664,I498672,I498712,I498720,I498737,I498754,I498794,I498816,I498833,I498859,I498867,I498884,I498901,I498918,I498935,I498980,I499011,I499028,I499054,I499062,I499093,I499110,I499127,I499144,I499216,I499242,I499250,I499290,I499298,I499315,I499332,I499372,I499394,I499411,I499437,I499445,I499462,I499479,I499496,I499513,I499558,I499589,I499606,I499632,I499640,I499671,I499688,I499705,I499722,I499794,I499820,I499828,I499868,I499876,I499893,I499910,I499950,I499972,I499989,I500015,I500023,I500040,I500057,I500074,I500091,I500136,I500167,I500184,I500210,I500218,I500249,I500266,I500283,I500300,I500372,I500398,I500406,I500446,I500454,I500471,I500488,I500528,I500550,I500567,I500593,I500601,I500618,I500635,I500652,I500669,I500714,I500745,I500762,I500788,I500796,I500827,I500844,I500861,I500878,I500950,I500976,I500984,I501024,I501032,I501049,I501066,I501106,I501128,I501145,I501171,I501179,I501196,I501213,I501230,I501247,I501292,I501323,I501340,I501366,I501374,I501405,I501422,I501439,I501456,I501528,I501554,I501562,I501602,I501610,I501627,I501644,I501684,I501706,I501723,I501749,I501757,I501774,I501791,I501808,I501825,I501870,I501901,I501918,I501944,I501952,I501983,I502000,I502017,I502034,I502106,I502132,I502140,I502166,I502183,I502205,I502222,I502239,I502256,I502273,I502304,I502321,I502338,I502355,I502400,I502417,I502434,I502493,I502519,I502527,I502544,I502561,I502592,I502650,I502676,I502684,I502710,I502727,I502749,I502766,I502783,I502800,I502817,I502848,I502865,I502882,I502899,I502944,I502961,I502978,I503037,I503063,I503071,I503088,I503105,I503136,I503194,I503220,I503228,I503254,I503271,I503293,I503310,I503327,I503344,I503361,I503392,I503409,I503426,I503443,I503488,I503505,I503522,I503581,I503607,I503615,I503632,I503649,I503680,I503738,I503764,I503772,I503798,I503815,I503837,I503854,I503871,I503888,I503905,I503936,I503953,I503970,I503987,I504032,I504049,I504066,I504125,I504151,I504159,I504176,I504193,I504224,I504282,I504308,I504316,I504342,I504359,I504381,I504398,I504415,I504432,I504449,I504480,I504497,I504514,I504531,I504576,I504593,I504610,I504669,I504695,I504703,I504720,I504737,I504768,I504826,I504852,I504860,I504886,I504903,I504925,I504942,I504959,I504976,I504993,I505024,I505041,I505058,I505075,I505120,I505137,I505154,I505213,I505239,I505247,I505264,I505281,I505312,I505370,I505396,I505404,I505430,I505447,I505469,I505486,I505503,I505520,I505537,I505568,I505585,I505602,I505619,I505664,I505681,I505698,I505757,I505783,I505791,I505808,I505825,I505856,I505914,I505940,I505948,I505974,I505991,I506013,I506030,I506047,I506064,I506081,I506112,I506129,I506146,I506163,I506208,I506225,I506242,I506301,I506327,I506335,I506352,I506369,I506400,I506458,I506484,I506492,I506518,I506535,I506557,I506574,I506591,I506608,I506625,I506656,I506673,I506690,I506707,I506752,I506769,I506786,I506845,I506871,I506879,I506896,I506913,I506944,I507002,I507028,I507036,I507062,I507079,I507101,I507118,I507135,I507152,I507169,I507200,I507217,I507234,I507251,I507296,I507313,I507330,I507389,I507415,I507423,I507440,I507457,I507488,I507546,I507572,I507580,I507606,I507623,I507538,I507645,I507662,I507679,I507696,I507713,I507517,I507744,I507761,I507778,I507795,I507520,I507535,I507840,I507857,I507874,I507532,I507529,I507526,I507933,I507959,I507967,I507984,I508001,I507514,I508032,I507523,I508090,I542527,I508116,I508124,I542512,I542506,I508150,I508167,I508189,I542500,I508206,I542521,I508223,I542509,I508240,I508257,I508288,I542518,I508305,I542524,I508322,I542515,I508339,I508384,I542503,I508401,I508418,I508477,I508503,I508511,I508528,I508545,I508576,I508634,I508660,I508668,I508694,I508711,I508626,I508733,I508750,I508767,I508784,I508801,I508605,I508832,I508849,I508866,I508883,I508608,I508623,I508928,I508945,I508962,I508620,I508617,I508614,I509021,I509047,I509055,I509072,I509089,I508602,I509120,I508611,I509178,I509204,I509212,I509238,I509255,I509277,I509294,I509311,I509328,I509345,I509376,I509393,I509410,I509427,I509472,I509489,I509506,I509565,I509591,I509599,I509616,I509633,I509664,I509722,I560377,I509748,I509756,I560362,I560356,I509782,I509799,I509714,I509821,I560350,I509838,I560371,I509855,I560359,I509872,I509889,I509693,I509920,I560368,I509937,I560374,I509954,I560365,I509971,I509696,I509711,I510016,I560353,I510033,I510050,I509708,I509705,I509702,I510109,I510135,I510143,I510160,I510177,I509690,I510208,I509699,I510266,I510292,I510300,I510326,I510343,I510365,I510382,I510399,I510416,I510433,I510464,I510481,I510498,I510515,I510560,I510577,I510594,I510653,I510679,I510687,I510704,I510721,I510752,I510810,I510836,I510844,I510870,I510887,I510909,I510926,I510943,I510960,I510977,I511008,I511025,I511042,I511059,I511104,I511121,I511138,I511197,I511223,I511231,I511248,I511265,I511296,I511354,I511380,I511388,I511414,I511431,I511453,I511470,I511487,I511504,I511521,I511552,I511569,I511586,I511603,I511648,I511665,I511682,I511741,I511767,I511775,I511792,I511809,I511840,I511898,I511924,I511932,I511958,I511975,I511997,I512014,I512031,I512048,I512065,I512096,I512113,I512130,I512147,I512192,I512209,I512226,I512285,I512311,I512319,I512336,I512353,I512384,I512442,I512468,I512476,I512502,I512519,I512541,I512558,I512575,I512592,I512609,I512640,I512657,I512674,I512691,I512736,I512753,I512770,I512829,I512855,I512863,I512880,I512897,I512928,I512986,I513012,I513020,I513046,I513063,I513085,I513102,I513119,I513136,I513153,I513184,I513201,I513218,I513235,I513280,I513297,I513314,I513373,I513399,I513407,I513424,I513441,I513472,I513530,I521701,I513556,I513564,I521710,I521713,I513590,I513607,I513629,I521707,I513646,I521704,I513663,I521698,I513680,I513697,I513728,I521695,I513745,I521692,I513762,I513779,I513824,I513841,I513858,I513917,I521716,I513943,I513951,I513968,I513985,I514016,I514074,I514100,I514108,I514134,I514151,I514173,I514190,I514207,I514224,I514241,I514272,I514289,I514306,I514323,I514368,I514385,I514402,I514461,I514487,I514495,I514512,I514529,I514560,I514618,I514644,I514652,I514678,I514695,I514610,I514717,I514734,I514751,I514768,I514785,I514589,I514816,I514833,I514850,I514867,I514592,I514607,I514912,I514929,I514946,I514604,I514601,I514598,I515005,I515031,I515039,I515056,I515073,I514586,I515104,I514595,I515162,I515188,I515196,I515222,I515239,I515261,I515278,I515295,I515312,I515329,I515360,I515377,I515394,I515411,I515456,I515473,I515490,I515549,I515575,I515583,I515600,I515617,I515648,I515706,I515732,I515740,I515766,I515783,I515698,I515805,I515822,I515839,I515856,I515873,I515677,I515904,I515921,I515938,I515955,I515680,I515695,I516000,I516017,I516034,I515692,I515689,I515686,I516093,I516119,I516127,I516144,I516161,I515674,I516192,I515683,I516250,I516276,I516284,I516310,I516327,I516349,I516366,I516383,I516400,I516417,I516448,I516465,I516482,I516499,I516544,I516561,I516578,I516637,I516663,I516671,I516688,I516705,I516736,I516794,I516820,I516828,I516854,I516871,I516893,I516910,I516927,I516944,I516961,I516992,I517009,I517026,I517043,I517088,I517105,I517122,I517181,I517207,I517215,I517232,I517249,I517280,I517338,I517364,I517372,I517398,I517415,I517437,I517454,I517471,I517488,I517505,I517536,I517553,I517570,I517587,I517632,I517649,I517666,I517725,I517751,I517759,I517776,I517793,I517824,I517882,I517908,I517916,I517942,I517959,I517981,I517998,I518015,I518032,I518049,I518080,I518097,I518114,I518131,I518176,I518193,I518210,I518269,I518295,I518303,I518320,I518337,I518368,I518426,I518452,I518460,I518486,I518503,I518525,I518542,I518559,I518576,I518593,I518624,I518641,I518658,I518675,I518720,I518737,I518754,I518813,I518839,I518847,I518864,I518881,I518912,I518970,I554427,I518996,I519004,I554412,I554406,I519030,I519047,I519069,I554400,I519086,I554421,I519103,I554409,I519120,I519137,I519168,I554418,I519185,I554424,I519202,I554415,I519219,I519264,I554403,I519281,I519298,I519357,I519383,I519391,I519408,I519425,I519456,I519514,I519540,I519548,I519574,I519591,I519613,I519630,I519647,I519664,I519681,I519712,I519729,I519746,I519763,I519808,I519825,I519842,I519901,I519927,I519935,I519952,I519969,I520000,I520058,I520084,I520092,I520118,I520135,I520050,I520157,I520174,I520191,I520208,I520225,I520029,I520256,I520273,I520290,I520307,I520032,I520047,I520352,I520369,I520386,I520044,I520041,I520038,I520445,I520471,I520479,I520496,I520513,I520026,I520544,I520035,I520602,I520628,I520636,I520662,I520679,I520701,I520718,I520735,I520752,I520769,I520800,I520817,I520834,I520851,I520896,I520913,I520930,I520989,I521015,I521023,I521040,I521057,I521088,I521146,I550854,I521172,I521180,I550845,I521197,I550830,I521223,I521231,I521248,I550833,I521265,I550842,I521282,I521299,I550839,I521330,I550851,I521347,I521364,I521395,I550836,I521412,I521452,I521460,I521491,I550857,I521508,I521525,I521542,I521573,I521604,I550848,I521630,I521652,I521724,I521750,I521758,I521775,I521801,I521809,I521826,I521843,I521860,I521877,I521908,I521925,I521942,I521973,I521990,I522030,I522038,I522069,I522086,I522103,I522120,I522151,I522182,I522208,I522230,I522302,I522328,I522336,I522353,I522379,I522387,I522404,I522421,I522438,I522455,I522486,I522503,I522520,I522551,I522568,I522608,I522616,I522647,I522664,I522681,I522698,I522729,I522760,I522786,I522808,I522880,I522906,I522914,I522931,I522957,I522965,I522982,I522999,I523016,I523033,I523064,I523081,I523098,I523129,I523146,I523186,I523194,I523225,I523242,I523259,I523276,I523307,I523338,I523364,I523386,I523458,I523484,I523492,I523509,I523535,I523543,I523560,I523577,I523594,I523611,I523642,I523659,I523676,I523707,I523724,I523764,I523772,I523803,I523820,I523837,I523854,I523885,I523916,I523942,I523964,I524036,I524062,I524070,I524087,I524113,I524121,I524138,I524155,I524172,I524189,I524220,I524237,I524254,I524285,I524302,I524342,I524350,I524381,I524398,I524415,I524432,I524463,I524494,I524520,I524542,I524614,I524640,I524648,I524665,I524691,I524699,I524716,I524733,I524750,I524767,I524798,I524815,I524832,I524863,I524880,I524920,I524928,I524959,I524976,I524993,I525010,I525041,I525072,I525098,I525120,I525192,I525218,I525226,I525243,I525269,I525277,I525294,I525311,I525328,I525345,I525376,I525393,I525410,I525441,I525458,I525498,I525506,I525537,I525554,I525571,I525588,I525619,I525650,I525676,I525698,I525770,I525796,I525804,I525821,I525847,I525855,I525872,I525889,I525906,I525923,I525954,I525971,I525988,I526019,I526036,I526076,I526084,I526115,I526132,I526149,I526166,I526197,I526228,I526254,I526276,I526348,I551449,I526374,I526382,I551440,I526399,I551425,I526425,I526433,I526450,I551428,I526467,I551437,I526484,I526501,I551434,I526532,I551446,I526549,I526566,I526597,I551431,I526614,I526654,I526662,I526693,I551452,I526710,I526727,I526744,I526775,I526806,I551443,I526832,I526854,I526926,I526952,I526960,I526977,I527003,I527011,I527028,I527045,I527062,I527079,I527110,I527127,I527144,I527175,I527192,I527232,I527240,I527271,I527288,I527305,I527322,I527353,I527384,I527410,I527432,I527504,I527530,I527538,I527555,I527581,I527589,I527606,I527623,I527640,I527657,I527688,I527705,I527722,I527753,I527770,I527810,I527818,I527849,I527866,I527883,I527900,I527931,I527962,I527988,I528010,I528082,I528108,I528116,I528133,I528159,I528167,I528184,I528201,I528218,I528235,I528266,I528283,I528300,I528331,I528348,I528388,I528396,I528427,I528444,I528461,I528478,I528509,I528540,I528566,I528588,I528660,I528686,I528694,I528711,I528737,I528745,I528762,I528779,I528796,I528813,I528844,I528861,I528878,I528909,I528926,I528966,I528974,I529005,I529022,I529039,I529056,I529087,I529118,I529144,I529166,I529238,I529264,I529272,I529289,I529315,I529323,I529340,I529357,I529374,I529391,I529422,I529439,I529456,I529487,I529504,I529544,I529552,I529583,I529600,I529617,I529634,I529665,I529696,I529722,I529744,I529816,I529842,I529850,I529867,I529893,I529901,I529918,I529935,I529952,I529969,I530000,I530017,I530034,I530065,I530082,I530122,I530130,I530161,I530178,I530195,I530212,I530243,I530274,I530300,I530322,I530394,I530420,I530428,I530445,I530471,I530479,I530496,I530513,I530530,I530547,I530578,I530595,I530612,I530643,I530660,I530700,I530708,I530739,I530756,I530773,I530790,I530821,I530852,I530878,I530900,I530972,I530998,I531006,I531023,I531049,I531057,I531074,I531091,I531108,I531125,I531156,I531173,I531190,I531221,I531238,I531278,I531286,I531317,I531334,I531351,I531368,I531399,I531430,I531456,I531478,I531550,I531576,I531584,I531601,I531627,I531635,I531652,I531669,I531686,I531703,I531734,I531751,I531768,I531799,I531816,I531856,I531864,I531895,I531912,I531929,I531946,I531977,I532008,I532034,I532056,I532128,I537826,I532154,I532162,I537820,I532179,I537835,I532205,I532213,I532230,I537811,I532247,I537808,I532264,I532281,I537814,I532312,I532329,I537823,I532346,I532377,I537817,I532394,I532434,I532442,I532473,I537832,I532490,I532507,I532524,I532555,I532586,I537829,I532612,I532634,I532706,I532732,I532740,I532757,I532783,I532791,I532808,I532825,I532842,I532859,I532890,I532907,I532924,I532955,I532972,I533012,I533020,I533051,I533068,I533085,I533102,I533133,I533164,I533190,I533212,I533284,I533310,I533318,I533335,I533361,I533369,I533386,I533403,I533420,I533437,I533276,I533468,I533485,I533502,I533255,I533533,I533550,I533261,I533590,I533598,I533270,I533629,I533646,I533663,I533680,I533273,I533711,I533252,I533742,I533768,I533267,I533790,I533264,I533258,I533862,I533888,I533896,I533913,I533939,I533947,I533964,I533981,I533998,I534015,I534046,I534063,I534080,I534111,I534128,I534168,I534176,I534207,I534224,I534241,I534258,I534289,I534320,I534346,I534368,I534440,I534466,I534474,I534491,I534517,I534525,I534542,I534559,I534576,I534593,I534624,I534641,I534658,I534689,I534706,I534746,I534754,I534785,I534802,I534819,I534836,I534867,I534898,I534924,I534946,I535018,I535044,I535052,I535069,I535095,I535103,I535120,I535137,I535154,I535171,I535202,I535219,I535236,I535267,I535284,I535324,I535332,I535363,I535380,I535397,I535414,I535445,I535476,I535502,I535524,I535599,I535625,I535633,I535650,I535676,I535684,I535701,I535718,I535749,I535780,I535797,I535814,I535831,I535848,I535879,I535938,I535955,I535981,I536003,I536029,I536037,I536054,I536085,I536160,I536186,I536194,I536211,I536237,I536245,I536262,I536279,I536310,I536341,I536358,I536375,I536392,I536409,I536440,I536499,I536516,I536542,I536564,I536590,I536598,I536615,I536646,I536721,I536747,I536755,I536772,I536798,I536806,I536823,I536840,I536871,I536902,I536919,I536936,I536953,I536970,I537001,I537060,I537077,I537103,I537125,I537151,I537159,I537176,I537207,I537282,I537308,I537316,I537333,I537359,I537367,I537384,I537401,I537432,I537463,I537480,I537497,I537514,I537531,I537562,I537621,I537638,I537664,I537686,I537712,I537720,I537737,I537768,I537843,I537869,I537877,I537894,I537920,I537928,I537945,I537962,I537993,I538024,I538041,I538058,I538075,I538092,I538123,I538182,I538199,I538225,I538247,I538273,I538281,I538298,I538329,I538404,I538430,I538438,I538455,I538481,I538489,I538506,I538523,I538554,I538585,I538602,I538619,I538636,I538653,I538684,I538743,I538760,I538786,I538808,I538834,I538842,I538859,I538890,I538965,I538991,I539008,I539016,I539061,I539078,I539095,I539112,I539129,I539146,I539163,I539194,I539211,I539256,I539273,I539290,I539321,I539347,I539355,I539386,I539403,I539420,I539446,I539454,I539471,I539560,I539586,I539603,I539611,I539656,I539673,I539690,I539707,I539724,I539741,I539758,I539789,I539806,I539851,I539868,I539885,I539916,I539942,I539950,I539981,I539998,I540015,I540041,I540049,I540066,I540155,I540181,I540198,I540206,I540251,I540268,I540285,I540302,I540319,I540336,I540353,I540384,I540401,I540446,I540463,I540480,I540511,I540537,I540545,I540576,I540593,I540610,I540636,I540644,I540661,I540750,I540776,I540793,I540801,I540846,I540863,I540880,I540897,I540914,I540931,I540948,I540979,I540996,I541041,I541058,I541075,I541106,I541132,I541140,I541171,I541188,I541205,I541231,I541239,I541256,I541345,I541371,I541388,I541396,I541441,I541458,I541475,I541492,I541509,I541526,I541543,I541574,I541591,I541636,I541653,I541670,I541701,I541727,I541735,I541766,I541783,I541800,I541826,I541834,I541851,I541940,I541966,I541983,I541991,I542036,I542053,I542070,I542087,I542104,I542121,I542138,I542169,I542186,I542231,I542248,I542265,I542296,I542322,I542330,I542361,I542378,I542395,I542421,I542429,I542446,I542535,I542561,I542578,I542586,I542631,I542648,I542665,I542682,I542699,I542716,I542733,I542764,I542781,I542826,I542843,I542860,I542891,I542917,I542925,I542956,I542973,I542990,I543016,I543024,I543041,I543130,I543156,I543173,I543181,I543226,I543243,I543260,I543277,I543294,I543311,I543328,I543359,I543376,I543421,I543438,I543455,I543486,I543512,I543520,I543551,I543568,I543585,I543611,I543619,I543636,I543725,I543751,I543768,I543776,I543821,I543838,I543855,I543872,I543889,I543906,I543923,I543954,I543971,I544016,I544033,I544050,I544081,I544107,I544115,I544146,I544163,I544180,I544206,I544214,I544231,I544320,I544346,I544363,I544371,I544416,I544433,I544450,I544467,I544484,I544501,I544518,I544549,I544566,I544611,I544628,I544645,I544676,I544702,I544710,I544741,I544758,I544775,I544801,I544809,I544826,I544915,I544941,I544958,I544966,I545011,I545028,I545045,I545062,I545079,I545096,I545113,I545144,I545161,I545206,I545223,I545240,I545271,I545297,I545305,I545336,I545353,I545370,I545396,I545404,I545421,I545510,I545536,I545553,I545561,I545606,I545623,I545640,I545657,I545674,I545691,I545708,I545739,I545756,I545801,I545818,I545835,I545866,I545892,I545900,I545931,I545948,I545965,I545991,I545999,I546016,I546105,I546131,I546148,I546156,I546201,I546218,I546235,I546252,I546269,I546286,I546303,I546334,I546351,I546396,I546413,I546430,I546461,I546487,I546495,I546526,I546543,I546560,I546586,I546594,I546611,I546700,I546726,I546743,I546751,I546796,I546813,I546830,I546847,I546864,I546881,I546898,I546929,I546946,I546991,I547008,I547025,I547056,I547082,I547090,I547121,I547138,I547155,I547181,I547189,I547206,I547295,I547321,I547338,I547346,I547391,I547408,I547425,I547442,I547459,I547476,I547493,I547524,I547541,I547586,I547603,I547620,I547651,I547677,I547685,I547716,I547733,I547750,I547776,I547784,I547801,I547890,I547916,I547933,I547941,I547986,I548003,I548020,I548037,I548054,I548071,I548088,I548119,I548136,I548181,I548198,I548215,I548246,I548272,I548280,I548311,I548328,I548345,I548371,I548379,I548396,I548485,I548511,I548528,I548536,I548581,I548598,I548615,I548632,I548649,I548666,I548683,I548714,I548731,I548776,I548793,I548810,I548841,I548867,I548875,I548906,I548923,I548940,I548966,I548974,I548991,I549080,I549106,I549123,I549131,I549176,I549193,I549210,I549227,I549244,I549261,I549278,I549309,I549326,I549371,I549388,I549405,I549436,I549462,I549470,I549501,I549518,I549535,I549561,I549569,I549586,I549675,I549701,I549718,I549726,I549771,I549788,I549805,I549822,I549839,I549856,I549873,I549904,I549921,I549966,I549983,I550000,I550031,I550057,I550065,I550096,I550113,I550130,I550156,I550164,I550181,I550270,I550296,I550313,I550321,I550366,I550383,I550400,I550417,I550434,I550451,I550468,I550499,I550516,I550561,I550578,I550595,I550626,I550652,I550660,I550691,I550708,I550725,I550751,I550759,I550776,I550865,I550891,I550908,I550916,I550961,I550978,I550995,I551012,I551029,I551046,I551063,I551094,I551111,I551156,I551173,I551190,I551221,I551247,I551255,I551286,I551303,I551320,I551346,I551354,I551371,I551460,I551486,I551503,I551511,I551556,I551573,I551590,I551607,I551624,I551641,I551658,I551689,I551706,I551751,I551768,I551785,I551816,I551842,I551850,I551881,I551898,I551915,I551941,I551949,I551966,I552055,I552081,I552098,I552106,I552151,I552168,I552185,I552202,I552219,I552236,I552253,I552284,I552301,I552346,I552363,I552380,I552411,I552437,I552445,I552476,I552493,I552510,I552536,I552544,I552561,I552650,I552676,I552693,I552701,I552746,I552763,I552780,I552797,I552814,I552831,I552848,I552879,I552896,I552941,I552958,I552975,I553006,I553032,I553040,I553071,I553088,I553105,I553131,I553139,I553156,I553245,I553271,I553288,I553296,I553341,I553358,I553375,I553392,I553409,I553426,I553443,I553474,I553491,I553536,I553553,I553570,I553601,I553627,I553635,I553666,I553683,I553700,I553726,I553734,I553751,I553840,I553866,I553883,I553891,I553936,I553953,I553970,I553987,I554004,I554021,I554038,I554069,I554086,I554131,I554148,I554165,I554196,I554222,I554230,I554261,I554278,I554295,I554321,I554329,I554346,I554435,I554461,I554478,I554486,I554531,I554548,I554565,I554582,I554599,I554616,I554633,I554664,I554681,I554726,I554743,I554760,I554791,I554817,I554825,I554856,I554873,I554890,I554916,I554924,I554941,I555030,I555056,I555073,I555081,I555126,I555143,I555160,I555177,I555194,I555211,I555228,I555259,I555276,I555321,I555338,I555355,I555386,I555412,I555420,I555451,I555468,I555485,I555511,I555519,I555536,I555625,I555651,I555668,I555676,I555721,I555738,I555755,I555772,I555789,I555806,I555823,I555854,I555871,I555916,I555933,I555950,I555981,I556007,I556015,I556046,I556063,I556080,I556106,I556114,I556131,I556220,I556246,I556263,I556271,I556316,I556333,I556350,I556367,I556384,I556401,I556418,I556449,I556466,I556511,I556528,I556545,I556576,I556602,I556610,I556641,I556658,I556675,I556701,I556709,I556726,I556815,I556841,I556858,I556866,I556911,I556928,I556945,I556962,I556979,I556996,I557013,I557044,I557061,I557106,I557123,I557140,I557171,I557197,I557205,I557236,I557253,I557270,I557296,I557304,I557321,I557410,I557436,I557453,I557461,I557506,I557523,I557540,I557557,I557574,I557591,I557608,I557639,I557656,I557701,I557718,I557735,I557766,I557792,I557800,I557831,I557848,I557865,I557891,I557899,I557916,I558005,I558031,I558048,I558056,I558101,I558118,I558135,I558152,I558169,I558186,I558203,I558234,I558251,I558296,I558313,I558330,I558361,I558387,I558395,I558426,I558443,I558460,I558486,I558494,I558511,I558600,I558626,I558643,I558651,I558696,I558713,I558730,I558747,I558764,I558781,I558798,I558829,I558846,I558891,I558908,I558925,I558956,I558982,I558990,I559021,I559038,I559055,I559081,I559089,I559106,I559195,I559221,I559238,I559246,I559291,I559308,I559325,I559342,I559359,I559376,I559393,I559424,I559441,I559486,I559503,I559520,I559551,I559577,I559585,I559616,I559633,I559650,I559676,I559684,I559701,I559790,I559816,I559833,I559841,I559886,I559903,I559920,I559937,I559954,I559971,I559988,I560019,I560036,I560081,I560098,I560115,I560146,I560172,I560180,I560211,I560228,I560245,I560271,I560279,I560296,I560385,I560411,I560428,I560436,I560481,I560498,I560515,I560532,I560549,I560566,I560583,I560614,I560631,I560676,I560693,I560710,I560741,I560767,I560775,I560806,I560823,I560840,I560866,I560874,I560891,I560980,I561006,I561023,I561031,I561076,I561093,I561110,I561127,I561144,I561161,I561178,I561209,I561226,I561271,I561288,I561305,I561336,I561362,I561370,I561401,I561418,I561435,I561461,I561469,I561486,I561575,I561601,I561618,I561626,I561671,I561688,I561705,I561722,I561739,I561756,I561773,I561804,I561821,I561866,I561883,I561900,I561931,I561957,I561965,I561996,I562013,I562030,I562056,I562064,I562081,I562170,I562196,I562213,I562221,I562266,I562283,I562300,I562317,I562334,I562351,I562368,I562399,I562416,I562461,I562478,I562495,I562526,I562552,I562560,I562591,I562608,I562625,I562651,I562659,I562676,I562765,I562791,I562808,I562816,I562861,I562878,I562895,I562912,I562929,I562946,I562963,I562994,I563011,I563056,I563073,I563090,I563121,I563147,I563155,I563186,I563203,I563220,I563246,I563254,I563271,I563360,I563386,I563403,I563411,I563456,I563473,I563490,I563507,I563524,I563541,I563558,I563589,I563606,I563651,I563668,I563685,I563716,I563742,I563750,I563781,I563798,I563815,I563841,I563849,I563866,I563955,I563981,I563998,I564006,I564051,I564068,I564085,I564102,I564119,I564136,I564153,I564184,I564201,I564246,I564263,I564280,I564311,I564337,I564345,I564376,I564393,I564410,I564436,I564444,I564461,I564550,I564576,I564593,I564601,I564646,I564663,I564680,I564697,I564714,I564731,I564748,I564779,I564796,I564841,I564858,I564875,I564906,I564932,I564940,I564971,I564988,I565005,I565031,I565039,I565056,I565145,I565171,I565188,I565196,I565241,I565258,I565275,I565292,I565309,I565326,I565343,I565374,I565391,I565436,I565453,I565470,I565501,I565527,I565535,I565566,I565583,I565600,I565626,I565634,I565651,I565740,I565766,I565783,I565791,I565836,I565853,I565870,I565887,I565904,I565921,I565938,I565969,I565986,I566031,I566048,I566065,I566096,I566122,I566130,I566161,I566178,I566195,I566221,I566229,I566246,I566335,I566361,I566378,I566386,I566431,I566448,I566465,I566482,I566499,I566516,I566533,I566564,I566581,I566626,I566643,I566660,I566691,I566717,I566725,I566756,I566773,I566790,I566816,I566824,I566841,I566930,I566956,I566973,I566981,I567026,I567043,I567060,I567077,I567094,I567111,I567128,I567159,I567176,I567221,I567238,I567255,I567286,I567312,I567320,I567351,I567368,I567385,I567411,I567419,I567436,I567525,I567551,I567568,I567576,I567621,I567638,I567655,I567672,I567689,I567706,I567723,I567754,I567771,I567816,I567833,I567850,I567881,I567907,I567915,I567946,I567963,I567980,I568006,I568014,I568031,I568120,I568146,I568163,I568171,I568216,I568233,I568250,I568267,I568284,I568301,I568318,I568349,I568366,I568411,I568428,I568445,I568476,I568502,I568510,I568541,I568558,I568575,I568601,I568609,I568626,I568715,I568741,I568758,I568766,I568811,I568828,I568845,I568862,I568879,I568896,I568913,I568944,I568961,I569006,I569023,I569040,I569071,I569097,I569105,I569136,I569153,I569170,I569196,I569204,I569221,I569310,I569336,I569353,I569361,I569406,I569423,I569440,I569457,I569474,I569491,I569508,I569539,I569556,I569601,I569618,I569635,I569666,I569692,I569700,I569731,I569748,I569765,I569791,I569799,I569816,I569905,I569931,I569948,I569956,I570001,I570018,I570035,I570052,I570069,I570086,I570103,I570134,I570151,I570196,I570213,I570230,I570261,I570287,I570295,I570326,I570343,I570360,I570386,I570394,I570411;
not I_0 (I2898,I2866);
DFFARX1 I_1 (I43137,I2859,I2898,I2924,);
nand I_2 (I2932,I2924,I43128);
not I_3 (I2949,I2932);
DFFARX1 I_4 (I2949,I2859,I2898,I2890,);
DFFARX1 I_5 (I43149,I2859,I2898,I2989,);
not I_6 (I2997,I2989);
not I_7 (I3014,I43125);
not I_8 (I3031,I43125);
nand I_9 (I3048,I2997,I3031);
nor I_10 (I3065,I3048,I43125);
DFFARX1 I_11 (I3065,I2859,I2898,I2869,);
nor I_12 (I3096,I43125,I43125);
nand I_13 (I3113,I2989,I3096);
nor I_14 (I3130,I43134,I43128);
nor I_15 (I2872,I3048,I43134);
not I_16 (I3161,I43134);
not I_17 (I3178,I43146);
nand I_18 (I3195,I3178,I43143);
nand I_19 (I3212,I3014,I3195);
not I_20 (I3229,I3212);
nor I_21 (I3246,I43146,I43128);
nor I_22 (I2881,I3229,I3246);
nor I_23 (I3277,I43140,I43146);
and I_24 (I3294,I3277,I3130);
nor I_25 (I3311,I3212,I3294);
DFFARX1 I_26 (I3311,I2859,I2898,I2887,);
nor I_27 (I3342,I2932,I3294);
DFFARX1 I_28 (I3342,I2859,I2898,I2884,);
nor I_29 (I3373,I43140,I43131);
DFFARX1 I_30 (I3373,I2859,I2898,I3399,);
nor I_31 (I3407,I3399,I43125);
nand I_32 (I3424,I3407,I3014);
nand I_33 (I2878,I3424,I3113);
nand I_34 (I2875,I3407,I3161);
not I_35 (I3493,I2866);
DFFARX1 I_36 (I309556,I2859,I3493,I3519,);
nand I_37 (I3527,I3519,I309535);
not I_38 (I3544,I3527);
DFFARX1 I_39 (I3544,I2859,I3493,I3485,);
DFFARX1 I_40 (I309544,I2859,I3493,I3584,);
not I_41 (I3592,I3584);
not I_42 (I3609,I309550);
not I_43 (I3626,I309547);
nand I_44 (I3643,I3592,I3626);
nor I_45 (I3660,I3643,I309550);
DFFARX1 I_46 (I3660,I2859,I3493,I3464,);
nor I_47 (I3691,I309547,I309550);
nand I_48 (I3708,I3584,I3691);
nor I_49 (I3725,I309538,I309532);
nor I_50 (I3467,I3643,I309538);
not I_51 (I3756,I309538);
not I_52 (I3773,I309553);
nand I_53 (I3790,I3773,I309535);
nand I_54 (I3807,I3609,I3790);
not I_55 (I3824,I3807);
nor I_56 (I3841,I309553,I309532);
nor I_57 (I3476,I3824,I3841);
nor I_58 (I3872,I309541,I309553);
and I_59 (I3889,I3872,I3725);
nor I_60 (I3906,I3807,I3889);
DFFARX1 I_61 (I3906,I2859,I3493,I3482,);
nor I_62 (I3937,I3527,I3889);
DFFARX1 I_63 (I3937,I2859,I3493,I3479,);
nor I_64 (I3968,I309541,I309532);
DFFARX1 I_65 (I3968,I2859,I3493,I3994,);
nor I_66 (I4002,I3994,I309547);
nand I_67 (I4019,I4002,I3609);
nand I_68 (I3473,I4019,I3708);
nand I_69 (I3470,I4002,I3756);
not I_70 (I4088,I2866);
DFFARX1 I_71 (I163534,I2859,I4088,I4114,);
nand I_72 (I4122,I4114,I163525);
not I_73 (I4139,I4122);
DFFARX1 I_74 (I4139,I2859,I4088,I4080,);
DFFARX1 I_75 (I163528,I2859,I4088,I4179,);
not I_76 (I4187,I4179);
not I_77 (I4204,I163522);
not I_78 (I4221,I163531);
nand I_79 (I4238,I4187,I4221);
nor I_80 (I4255,I4238,I163522);
DFFARX1 I_81 (I4255,I2859,I4088,I4059,);
nor I_82 (I4286,I163531,I163522);
nand I_83 (I4303,I4179,I4286);
nor I_84 (I4320,I163519,I163537);
nor I_85 (I4062,I4238,I163519);
not I_86 (I4351,I163519);
not I_87 (I4368,I163519);
nand I_88 (I4385,I4368,I163543);
nand I_89 (I4402,I4204,I4385);
not I_90 (I4419,I4402);
nor I_91 (I4436,I163519,I163537);
nor I_92 (I4071,I4419,I4436);
nor I_93 (I4467,I163540,I163519);
and I_94 (I4484,I4467,I4320);
nor I_95 (I4501,I4402,I4484);
DFFARX1 I_96 (I4501,I2859,I4088,I4077,);
nor I_97 (I4532,I4122,I4484);
DFFARX1 I_98 (I4532,I2859,I4088,I4074,);
nor I_99 (I4563,I163540,I163546);
DFFARX1 I_100 (I4563,I2859,I4088,I4589,);
nor I_101 (I4597,I4589,I163531);
nand I_102 (I4614,I4597,I4204);
nand I_103 (I4068,I4614,I4303);
nand I_104 (I4065,I4597,I4351);
not I_105 (I4686,I2866);
DFFARX1 I_106 (I120332,I2859,I4686,I4712,);
DFFARX1 I_107 (I4712,I2859,I4686,I4729,);
not I_108 (I4737,I4729);
nand I_109 (I4754,I120329,I120323);
and I_110 (I4771,I4754,I120317);
DFFARX1 I_111 (I4771,I2859,I4686,I4797,);
DFFARX1 I_112 (I4797,I2859,I4686,I4678,);
DFFARX1 I_113 (I4797,I2859,I4686,I4669,);
DFFARX1 I_114 (I120305,I2859,I4686,I4842,);
nand I_115 (I4850,I4842,I120314);
not I_116 (I4867,I4850);
nor I_117 (I4666,I4712,I4867);
DFFARX1 I_118 (I120311,I2859,I4686,I4907,);
not I_119 (I4915,I4907);
nor I_120 (I4672,I4915,I4737);
nand I_121 (I4660,I4915,I4850);
nand I_122 (I4960,I120308,I120326);
and I_123 (I4977,I4960,I120305);
DFFARX1 I_124 (I4977,I2859,I4686,I5003,);
nor I_125 (I5011,I5003,I4712);
DFFARX1 I_126 (I5011,I2859,I4686,I4654,);
not I_127 (I5042,I5003);
nor I_128 (I5059,I120320,I120326);
not I_129 (I5076,I5059);
nor I_130 (I5093,I4850,I5076);
nor I_131 (I5110,I5042,I5093);
DFFARX1 I_132 (I5110,I2859,I4686,I4675,);
nor I_133 (I5141,I5003,I5076);
nor I_134 (I4663,I4867,I5141);
nor I_135 (I4657,I5003,I5059);
not I_136 (I5213,I2866);
DFFARX1 I_137 (I474932,I2859,I5213,I5239,);
DFFARX1 I_138 (I5239,I2859,I5213,I5256,);
not I_139 (I5264,I5256);
nand I_140 (I5281,I474920,I474911);
and I_141 (I5298,I5281,I474908);
DFFARX1 I_142 (I5298,I2859,I5213,I5324,);
DFFARX1 I_143 (I5324,I2859,I5213,I5205,);
DFFARX1 I_144 (I5324,I2859,I5213,I5196,);
DFFARX1 I_145 (I474914,I2859,I5213,I5369,);
nand I_146 (I5377,I5369,I474926);
not I_147 (I5394,I5377);
nor I_148 (I5193,I5239,I5394);
DFFARX1 I_149 (I474923,I2859,I5213,I5434,);
not I_150 (I5442,I5434);
nor I_151 (I5199,I5442,I5264);
nand I_152 (I5187,I5442,I5377);
nand I_153 (I5487,I474917,I474911);
and I_154 (I5504,I5487,I474929);
DFFARX1 I_155 (I5504,I2859,I5213,I5530,);
nor I_156 (I5538,I5530,I5239);
DFFARX1 I_157 (I5538,I2859,I5213,I5181,);
not I_158 (I5569,I5530);
nor I_159 (I5586,I474908,I474911);
not I_160 (I5603,I5586);
nor I_161 (I5620,I5377,I5603);
nor I_162 (I5637,I5569,I5620);
DFFARX1 I_163 (I5637,I2859,I5213,I5202,);
nor I_164 (I5668,I5530,I5603);
nor I_165 (I5190,I5394,I5668);
nor I_166 (I5184,I5530,I5586);
not I_167 (I5740,I2866);
DFFARX1 I_168 (I176507,I2859,I5740,I5766,);
DFFARX1 I_169 (I5766,I2859,I5740,I5783,);
not I_170 (I5791,I5783);
nand I_171 (I5808,I176507,I176510);
and I_172 (I5825,I5808,I176531);
DFFARX1 I_173 (I5825,I2859,I5740,I5851,);
DFFARX1 I_174 (I5851,I2859,I5740,I5732,);
DFFARX1 I_175 (I5851,I2859,I5740,I5723,);
DFFARX1 I_176 (I176519,I2859,I5740,I5896,);
nand I_177 (I5904,I5896,I176522);
not I_178 (I5921,I5904);
nor I_179 (I5720,I5766,I5921);
DFFARX1 I_180 (I176528,I2859,I5740,I5961,);
not I_181 (I5969,I5961);
nor I_182 (I5726,I5969,I5791);
nand I_183 (I5714,I5969,I5904);
nand I_184 (I6014,I176525,I176513);
and I_185 (I6031,I6014,I176516);
DFFARX1 I_186 (I6031,I2859,I5740,I6057,);
nor I_187 (I6065,I6057,I5766);
DFFARX1 I_188 (I6065,I2859,I5740,I5708,);
not I_189 (I6096,I6057);
nor I_190 (I6113,I176534,I176513);
not I_191 (I6130,I6113);
nor I_192 (I6147,I5904,I6130);
nor I_193 (I6164,I6096,I6147);
DFFARX1 I_194 (I6164,I2859,I5740,I5729,);
nor I_195 (I6195,I6057,I6130);
nor I_196 (I5717,I5921,I6195);
nor I_197 (I5711,I6057,I6113);
not I_198 (I6267,I2866);
DFFARX1 I_199 (I150898,I2859,I6267,I6293,);
DFFARX1 I_200 (I6293,I2859,I6267,I6310,);
not I_201 (I6318,I6310);
nand I_202 (I6335,I150895,I150889);
and I_203 (I6352,I6335,I150883);
DFFARX1 I_204 (I6352,I2859,I6267,I6378,);
DFFARX1 I_205 (I6378,I2859,I6267,I6259,);
DFFARX1 I_206 (I6378,I2859,I6267,I6250,);
DFFARX1 I_207 (I150871,I2859,I6267,I6423,);
nand I_208 (I6431,I6423,I150880);
not I_209 (I6448,I6431);
nor I_210 (I6247,I6293,I6448);
DFFARX1 I_211 (I150877,I2859,I6267,I6488,);
not I_212 (I6496,I6488);
nor I_213 (I6253,I6496,I6318);
nand I_214 (I6241,I6496,I6431);
nand I_215 (I6541,I150874,I150892);
and I_216 (I6558,I6541,I150871);
DFFARX1 I_217 (I6558,I2859,I6267,I6584,);
nor I_218 (I6592,I6584,I6293);
DFFARX1 I_219 (I6592,I2859,I6267,I6235,);
not I_220 (I6623,I6584);
nor I_221 (I6640,I150886,I150892);
not I_222 (I6657,I6640);
nor I_223 (I6674,I6431,I6657);
nor I_224 (I6691,I6623,I6674);
DFFARX1 I_225 (I6691,I2859,I6267,I6256,);
nor I_226 (I6722,I6584,I6657);
nor I_227 (I6244,I6448,I6722);
nor I_228 (I6238,I6584,I6640);
not I_229 (I6794,I2866);
DFFARX1 I_230 (I520570,I2859,I6794,I6820,);
DFFARX1 I_231 (I6820,I2859,I6794,I6837,);
not I_232 (I6845,I6837);
nand I_233 (I6862,I520588,I520582);
and I_234 (I6879,I6862,I520591);
DFFARX1 I_235 (I6879,I2859,I6794,I6905,);
DFFARX1 I_236 (I6905,I2859,I6794,I6786,);
DFFARX1 I_237 (I6905,I2859,I6794,I6777,);
DFFARX1 I_238 (I520576,I2859,I6794,I6950,);
nand I_239 (I6958,I6950,I520585);
not I_240 (I6975,I6958);
nor I_241 (I6774,I6820,I6975);
DFFARX1 I_242 (I520573,I2859,I6794,I7015,);
not I_243 (I7023,I7015);
nor I_244 (I6780,I7023,I6845);
nand I_245 (I6768,I7023,I6958);
nand I_246 (I7068,I520594,I520579);
and I_247 (I7085,I7068,I520573);
DFFARX1 I_248 (I7085,I2859,I6794,I7111,);
nor I_249 (I7119,I7111,I6820);
DFFARX1 I_250 (I7119,I2859,I6794,I6762,);
not I_251 (I7150,I7111);
nor I_252 (I7167,I520570,I520579);
not I_253 (I7184,I7167);
nor I_254 (I7201,I6958,I7184);
nor I_255 (I7218,I7150,I7201);
DFFARX1 I_256 (I7218,I2859,I6794,I6783,);
nor I_257 (I7249,I7111,I7184);
nor I_258 (I6771,I6975,I7249);
nor I_259 (I6765,I7111,I7167);
not I_260 (I7321,I2866);
DFFARX1 I_261 (I172699,I2859,I7321,I7347,);
DFFARX1 I_262 (I7347,I2859,I7321,I7364,);
not I_263 (I7372,I7364);
nand I_264 (I7389,I172699,I172702);
and I_265 (I7406,I7389,I172723);
DFFARX1 I_266 (I7406,I2859,I7321,I7432,);
DFFARX1 I_267 (I7432,I2859,I7321,I7313,);
DFFARX1 I_268 (I7432,I2859,I7321,I7304,);
DFFARX1 I_269 (I172711,I2859,I7321,I7477,);
nand I_270 (I7485,I7477,I172714);
not I_271 (I7502,I7485);
nor I_272 (I7301,I7347,I7502);
DFFARX1 I_273 (I172720,I2859,I7321,I7542,);
not I_274 (I7550,I7542);
nor I_275 (I7307,I7550,I7372);
nand I_276 (I7295,I7550,I7485);
nand I_277 (I7595,I172717,I172705);
and I_278 (I7612,I7595,I172708);
DFFARX1 I_279 (I7612,I2859,I7321,I7638,);
nor I_280 (I7646,I7638,I7347);
DFFARX1 I_281 (I7646,I2859,I7321,I7289,);
not I_282 (I7677,I7638);
nor I_283 (I7694,I172726,I172705);
not I_284 (I7711,I7694);
nor I_285 (I7728,I7485,I7711);
nor I_286 (I7745,I7677,I7728);
DFFARX1 I_287 (I7745,I2859,I7321,I7310,);
nor I_288 (I7776,I7638,I7711);
nor I_289 (I7298,I7502,I7776);
nor I_290 (I7292,I7638,I7694);
not I_291 (I7848,I2866);
DFFARX1 I_292 (I295666,I2859,I7848,I7874,);
DFFARX1 I_293 (I7874,I2859,I7848,I7891,);
not I_294 (I7899,I7891);
nand I_295 (I7916,I295681,I295684);
and I_296 (I7933,I7916,I295663);
DFFARX1 I_297 (I7933,I2859,I7848,I7959,);
DFFARX1 I_298 (I7959,I2859,I7848,I7840,);
DFFARX1 I_299 (I7959,I2859,I7848,I7831,);
DFFARX1 I_300 (I295669,I2859,I7848,I8004,);
nand I_301 (I8012,I8004,I295675);
not I_302 (I8029,I8012);
nor I_303 (I7828,I7874,I8029);
DFFARX1 I_304 (I295663,I2859,I7848,I8069,);
not I_305 (I8077,I8069);
nor I_306 (I7834,I8077,I7899);
nand I_307 (I7822,I8077,I8012);
nand I_308 (I8122,I295678,I295660);
and I_309 (I8139,I8122,I295672);
DFFARX1 I_310 (I8139,I2859,I7848,I8165,);
nor I_311 (I8173,I8165,I7874);
DFFARX1 I_312 (I8173,I2859,I7848,I7816,);
not I_313 (I8204,I8165);
nor I_314 (I8221,I295660,I295660);
not I_315 (I8238,I8221);
nor I_316 (I8255,I8012,I8238);
nor I_317 (I8272,I8204,I8255);
DFFARX1 I_318 (I8272,I2859,I7848,I7837,);
nor I_319 (I8303,I8165,I8238);
nor I_320 (I7825,I8029,I8303);
nor I_321 (I7819,I8165,I8221);
not I_322 (I8375,I2866);
DFFARX1 I_323 (I77454,I2859,I8375,I8401,);
DFFARX1 I_324 (I8401,I2859,I8375,I8418,);
not I_325 (I8426,I8418);
nand I_326 (I8443,I77472,I77457);
and I_327 (I8460,I8443,I77460);
DFFARX1 I_328 (I8460,I2859,I8375,I8486,);
DFFARX1 I_329 (I8486,I2859,I8375,I8367,);
DFFARX1 I_330 (I8486,I2859,I8375,I8358,);
DFFARX1 I_331 (I77448,I2859,I8375,I8531,);
nand I_332 (I8539,I8531,I77451);
not I_333 (I8556,I8539);
nor I_334 (I8355,I8401,I8556);
DFFARX1 I_335 (I77463,I2859,I8375,I8596,);
not I_336 (I8604,I8596);
nor I_337 (I8361,I8604,I8426);
nand I_338 (I8349,I8604,I8539);
nand I_339 (I8649,I77469,I77466);
and I_340 (I8666,I8649,I77451);
DFFARX1 I_341 (I8666,I2859,I8375,I8692,);
nor I_342 (I8700,I8692,I8401);
DFFARX1 I_343 (I8700,I2859,I8375,I8343,);
not I_344 (I8731,I8692);
nor I_345 (I8748,I77448,I77466);
not I_346 (I8765,I8748);
nor I_347 (I8782,I8539,I8765);
nor I_348 (I8799,I8731,I8782);
DFFARX1 I_349 (I8799,I2859,I8375,I8364,);
nor I_350 (I8830,I8692,I8765);
nor I_351 (I8352,I8556,I8830);
nor I_352 (I8346,I8692,I8748);
not I_353 (I8902,I2866);
DFFARX1 I_354 (I568680,I2859,I8902,I8928,);
DFFARX1 I_355 (I8928,I2859,I8902,I8945,);
not I_356 (I8953,I8945);
nand I_357 (I8970,I568683,I568689);
and I_358 (I8987,I8970,I568698);
DFFARX1 I_359 (I8987,I2859,I8902,I9013,);
DFFARX1 I_360 (I9013,I2859,I8902,I8894,);
DFFARX1 I_361 (I9013,I2859,I8902,I8885,);
DFFARX1 I_362 (I568701,I2859,I8902,I9058,);
nand I_363 (I9066,I9058,I568692);
not I_364 (I9083,I9066);
nor I_365 (I8882,I8928,I9083);
DFFARX1 I_366 (I568680,I2859,I8902,I9123,);
not I_367 (I9131,I9123);
nor I_368 (I8888,I9131,I8953);
nand I_369 (I8876,I9131,I9066);
nand I_370 (I9176,I568707,I568686);
and I_371 (I9193,I9176,I568695);
DFFARX1 I_372 (I9193,I2859,I8902,I9219,);
nor I_373 (I9227,I9219,I8928);
DFFARX1 I_374 (I9227,I2859,I8902,I8870,);
not I_375 (I9258,I9219);
nor I_376 (I9275,I568704,I568686);
not I_377 (I9292,I9275);
nor I_378 (I9309,I9066,I9292);
nor I_379 (I9326,I9258,I9309);
DFFARX1 I_380 (I9326,I2859,I8902,I8891,);
nor I_381 (I9357,I9219,I9292);
nor I_382 (I8879,I9083,I9357);
nor I_383 (I8873,I9219,I9275);
not I_384 (I9429,I2866);
DFFARX1 I_385 (I510234,I2859,I9429,I9455,);
DFFARX1 I_386 (I9455,I2859,I9429,I9472,);
not I_387 (I9480,I9472);
nand I_388 (I9497,I510252,I510246);
and I_389 (I9514,I9497,I510255);
DFFARX1 I_390 (I9514,I2859,I9429,I9540,);
DFFARX1 I_391 (I9540,I2859,I9429,I9421,);
DFFARX1 I_392 (I9540,I2859,I9429,I9412,);
DFFARX1 I_393 (I510240,I2859,I9429,I9585,);
nand I_394 (I9593,I9585,I510249);
not I_395 (I9610,I9593);
nor I_396 (I9409,I9455,I9610);
DFFARX1 I_397 (I510237,I2859,I9429,I9650,);
not I_398 (I9658,I9650);
nor I_399 (I9415,I9658,I9480);
nand I_400 (I9403,I9658,I9593);
nand I_401 (I9703,I510258,I510243);
and I_402 (I9720,I9703,I510237);
DFFARX1 I_403 (I9720,I2859,I9429,I9746,);
nor I_404 (I9754,I9746,I9455);
DFFARX1 I_405 (I9754,I2859,I9429,I9397,);
not I_406 (I9785,I9746);
nor I_407 (I9802,I510234,I510243);
not I_408 (I9819,I9802);
nor I_409 (I9836,I9593,I9819);
nor I_410 (I9853,I9785,I9836);
DFFARX1 I_411 (I9853,I2859,I9429,I9418,);
nor I_412 (I9884,I9746,I9819);
nor I_413 (I9406,I9610,I9884);
nor I_414 (I9400,I9746,I9802);
not I_415 (I9956,I2866);
DFFARX1 I_416 (I567490,I2859,I9956,I9982,);
DFFARX1 I_417 (I9982,I2859,I9956,I9999,);
not I_418 (I10007,I9999);
nand I_419 (I10024,I567493,I567499);
and I_420 (I10041,I10024,I567508);
DFFARX1 I_421 (I10041,I2859,I9956,I10067,);
DFFARX1 I_422 (I10067,I2859,I9956,I9948,);
DFFARX1 I_423 (I10067,I2859,I9956,I9939,);
DFFARX1 I_424 (I567511,I2859,I9956,I10112,);
nand I_425 (I10120,I10112,I567502);
not I_426 (I10137,I10120);
nor I_427 (I9936,I9982,I10137);
DFFARX1 I_428 (I567490,I2859,I9956,I10177,);
not I_429 (I10185,I10177);
nor I_430 (I9942,I10185,I10007);
nand I_431 (I9930,I10185,I10120);
nand I_432 (I10230,I567517,I567496);
and I_433 (I10247,I10230,I567505);
DFFARX1 I_434 (I10247,I2859,I9956,I10273,);
nor I_435 (I10281,I10273,I9982);
DFFARX1 I_436 (I10281,I2859,I9956,I9924,);
not I_437 (I10312,I10273);
nor I_438 (I10329,I567514,I567496);
not I_439 (I10346,I10329);
nor I_440 (I10363,I10120,I10346);
nor I_441 (I10380,I10312,I10363);
DFFARX1 I_442 (I10380,I2859,I9956,I9945,);
nor I_443 (I10411,I10273,I10346);
nor I_444 (I9933,I10137,I10411);
nor I_445 (I9927,I10273,I10329);
not I_446 (I10483,I2866);
DFFARX1 I_447 (I485914,I2859,I10483,I10509,);
DFFARX1 I_448 (I10509,I2859,I10483,I10526,);
not I_449 (I10534,I10526);
nand I_450 (I10551,I485902,I485893);
and I_451 (I10568,I10551,I485890);
DFFARX1 I_452 (I10568,I2859,I10483,I10594,);
DFFARX1 I_453 (I10594,I2859,I10483,I10475,);
DFFARX1 I_454 (I10594,I2859,I10483,I10466,);
DFFARX1 I_455 (I485896,I2859,I10483,I10639,);
nand I_456 (I10647,I10639,I485908);
not I_457 (I10664,I10647);
nor I_458 (I10463,I10509,I10664);
DFFARX1 I_459 (I485905,I2859,I10483,I10704,);
not I_460 (I10712,I10704);
nor I_461 (I10469,I10712,I10534);
nand I_462 (I10457,I10712,I10647);
nand I_463 (I10757,I485899,I485893);
and I_464 (I10774,I10757,I485911);
DFFARX1 I_465 (I10774,I2859,I10483,I10800,);
nor I_466 (I10808,I10800,I10509);
DFFARX1 I_467 (I10808,I2859,I10483,I10451,);
not I_468 (I10839,I10800);
nor I_469 (I10856,I485890,I485893);
not I_470 (I10873,I10856);
nor I_471 (I10890,I10647,I10873);
nor I_472 (I10907,I10839,I10890);
DFFARX1 I_473 (I10907,I2859,I10483,I10472,);
nor I_474 (I10938,I10800,I10873);
nor I_475 (I10460,I10664,I10938);
nor I_476 (I10454,I10800,I10856);
not I_477 (I11010,I2866);
DFFARX1 I_478 (I155114,I2859,I11010,I11036,);
DFFARX1 I_479 (I11036,I2859,I11010,I11053,);
not I_480 (I11061,I11053);
nand I_481 (I11078,I155111,I155105);
and I_482 (I11095,I11078,I155099);
DFFARX1 I_483 (I11095,I2859,I11010,I11121,);
DFFARX1 I_484 (I11121,I2859,I11010,I11002,);
DFFARX1 I_485 (I11121,I2859,I11010,I10993,);
DFFARX1 I_486 (I155087,I2859,I11010,I11166,);
nand I_487 (I11174,I11166,I155096);
not I_488 (I11191,I11174);
nor I_489 (I10990,I11036,I11191);
DFFARX1 I_490 (I155093,I2859,I11010,I11231,);
not I_491 (I11239,I11231);
nor I_492 (I10996,I11239,I11061);
nand I_493 (I10984,I11239,I11174);
nand I_494 (I11284,I155090,I155108);
and I_495 (I11301,I11284,I155087);
DFFARX1 I_496 (I11301,I2859,I11010,I11327,);
nor I_497 (I11335,I11327,I11036);
DFFARX1 I_498 (I11335,I2859,I11010,I10978,);
not I_499 (I11366,I11327);
nor I_500 (I11383,I155102,I155108);
not I_501 (I11400,I11383);
nor I_502 (I11417,I11174,I11400);
nor I_503 (I11434,I11366,I11417);
DFFARX1 I_504 (I11434,I2859,I11010,I10999,);
nor I_505 (I11465,I11327,I11400);
nor I_506 (I10987,I11191,I11465);
nor I_507 (I10981,I11327,I11383);
not I_508 (I11537,I2866);
DFFARX1 I_509 (I233829,I2859,I11537,I11563,);
DFFARX1 I_510 (I11563,I2859,I11537,I11580,);
not I_511 (I11588,I11580);
nand I_512 (I11605,I233814,I233832);
and I_513 (I11622,I11605,I233826);
DFFARX1 I_514 (I11622,I2859,I11537,I11648,);
DFFARX1 I_515 (I11648,I2859,I11537,I11529,);
DFFARX1 I_516 (I11648,I2859,I11537,I11520,);
DFFARX1 I_517 (I233823,I2859,I11537,I11693,);
nand I_518 (I11701,I11693,I233814);
not I_519 (I11718,I11701);
nor I_520 (I11517,I11563,I11718);
DFFARX1 I_521 (I233817,I2859,I11537,I11758,);
not I_522 (I11766,I11758);
nor I_523 (I11523,I11766,I11588);
nand I_524 (I11511,I11766,I11701);
nand I_525 (I11811,I233838,I233820);
and I_526 (I11828,I11811,I233835);
DFFARX1 I_527 (I11828,I2859,I11537,I11854,);
nor I_528 (I11862,I11854,I11563);
DFFARX1 I_529 (I11862,I2859,I11537,I11505,);
not I_530 (I11893,I11854);
nor I_531 (I11910,I233817,I233820);
not I_532 (I11927,I11910);
nor I_533 (I11944,I11701,I11927);
nor I_534 (I11961,I11893,I11944);
DFFARX1 I_535 (I11961,I2859,I11537,I11526,);
nor I_536 (I11992,I11854,I11927);
nor I_537 (I11514,I11718,I11992);
nor I_538 (I11508,I11854,I11910);
not I_539 (I12064,I2866);
DFFARX1 I_540 (I190651,I2859,I12064,I12090,);
DFFARX1 I_541 (I12090,I2859,I12064,I12107,);
not I_542 (I12115,I12107);
nand I_543 (I12132,I190651,I190654);
and I_544 (I12149,I12132,I190675);
DFFARX1 I_545 (I12149,I2859,I12064,I12175,);
DFFARX1 I_546 (I12175,I2859,I12064,I12056,);
DFFARX1 I_547 (I12175,I2859,I12064,I12047,);
DFFARX1 I_548 (I190663,I2859,I12064,I12220,);
nand I_549 (I12228,I12220,I190666);
not I_550 (I12245,I12228);
nor I_551 (I12044,I12090,I12245);
DFFARX1 I_552 (I190672,I2859,I12064,I12285,);
not I_553 (I12293,I12285);
nor I_554 (I12050,I12293,I12115);
nand I_555 (I12038,I12293,I12228);
nand I_556 (I12338,I190669,I190657);
and I_557 (I12355,I12338,I190660);
DFFARX1 I_558 (I12355,I2859,I12064,I12381,);
nor I_559 (I12389,I12381,I12090);
DFFARX1 I_560 (I12389,I2859,I12064,I12032,);
not I_561 (I12420,I12381);
nor I_562 (I12437,I190678,I190657);
not I_563 (I12454,I12437);
nor I_564 (I12471,I12228,I12454);
nor I_565 (I12488,I12420,I12471);
DFFARX1 I_566 (I12488,I2859,I12064,I12053,);
nor I_567 (I12519,I12381,I12454);
nor I_568 (I12041,I12245,I12519);
nor I_569 (I12035,I12381,I12437);
not I_570 (I12591,I2866);
DFFARX1 I_571 (I1508,I2859,I12591,I12617,);
DFFARX1 I_572 (I12617,I2859,I12591,I12634,);
not I_573 (I12642,I12634);
nand I_574 (I12659,I1444,I1940);
and I_575 (I12676,I12659,I1908);
DFFARX1 I_576 (I12676,I2859,I12591,I12702,);
DFFARX1 I_577 (I12702,I2859,I12591,I12583,);
DFFARX1 I_578 (I12702,I2859,I12591,I12574,);
DFFARX1 I_579 (I2732,I2859,I12591,I12747,);
nand I_580 (I12755,I12747,I2468);
not I_581 (I12772,I12755);
nor I_582 (I12571,I12617,I12772);
DFFARX1 I_583 (I2044,I2859,I12591,I12812,);
not I_584 (I12820,I12812);
nor I_585 (I12577,I12820,I12642);
nand I_586 (I12565,I12820,I12755);
nand I_587 (I12865,I2716,I2164);
and I_588 (I12882,I12865,I1436);
DFFARX1 I_589 (I12882,I2859,I12591,I12908,);
nor I_590 (I12916,I12908,I12617);
DFFARX1 I_591 (I12916,I2859,I12591,I12559,);
not I_592 (I12947,I12908);
nor I_593 (I12964,I1812,I2164);
not I_594 (I12981,I12964);
nor I_595 (I12998,I12755,I12981);
nor I_596 (I13015,I12947,I12998);
DFFARX1 I_597 (I13015,I2859,I12591,I12580,);
nor I_598 (I13046,I12908,I12981);
nor I_599 (I12568,I12772,I13046);
nor I_600 (I12562,I12908,I12964);
not I_601 (I13118,I2866);
DFFARX1 I_602 (I97684,I2859,I13118,I13144,);
DFFARX1 I_603 (I13144,I2859,I13118,I13161,);
not I_604 (I13169,I13161);
nand I_605 (I13186,I97702,I97687);
and I_606 (I13203,I13186,I97690);
DFFARX1 I_607 (I13203,I2859,I13118,I13229,);
DFFARX1 I_608 (I13229,I2859,I13118,I13110,);
DFFARX1 I_609 (I13229,I2859,I13118,I13101,);
DFFARX1 I_610 (I97678,I2859,I13118,I13274,);
nand I_611 (I13282,I13274,I97681);
not I_612 (I13299,I13282);
nor I_613 (I13098,I13144,I13299);
DFFARX1 I_614 (I97693,I2859,I13118,I13339,);
not I_615 (I13347,I13339);
nor I_616 (I13104,I13347,I13169);
nand I_617 (I13092,I13347,I13282);
nand I_618 (I13392,I97699,I97696);
and I_619 (I13409,I13392,I97681);
DFFARX1 I_620 (I13409,I2859,I13118,I13435,);
nor I_621 (I13443,I13435,I13144);
DFFARX1 I_622 (I13443,I2859,I13118,I13086,);
not I_623 (I13474,I13435);
nor I_624 (I13491,I97678,I97696);
not I_625 (I13508,I13491);
nor I_626 (I13525,I13282,I13508);
nor I_627 (I13542,I13474,I13525);
DFFARX1 I_628 (I13542,I2859,I13118,I13107,);
nor I_629 (I13573,I13435,I13508);
nor I_630 (I13095,I13299,I13573);
nor I_631 (I13089,I13435,I13491);
not I_632 (I13645,I2866);
DFFARX1 I_633 (I400965,I2859,I13645,I13671,);
DFFARX1 I_634 (I13671,I2859,I13645,I13688,);
not I_635 (I13696,I13688);
nand I_636 (I13713,I400941,I400968);
and I_637 (I13730,I13713,I400953);
DFFARX1 I_638 (I13730,I2859,I13645,I13756,);
DFFARX1 I_639 (I13756,I2859,I13645,I13637,);
DFFARX1 I_640 (I13756,I2859,I13645,I13628,);
DFFARX1 I_641 (I400959,I2859,I13645,I13801,);
nand I_642 (I13809,I13801,I400944);
not I_643 (I13826,I13809);
nor I_644 (I13625,I13671,I13826);
DFFARX1 I_645 (I400962,I2859,I13645,I13866,);
not I_646 (I13874,I13866);
nor I_647 (I13631,I13874,I13696);
nand I_648 (I13619,I13874,I13809);
nand I_649 (I13919,I400947,I400950);
and I_650 (I13936,I13919,I400941);
DFFARX1 I_651 (I13936,I2859,I13645,I13962,);
nor I_652 (I13970,I13962,I13671);
DFFARX1 I_653 (I13970,I2859,I13645,I13613,);
not I_654 (I14001,I13962);
nor I_655 (I14018,I400956,I400950);
not I_656 (I14035,I14018);
nor I_657 (I14052,I13809,I14035);
nor I_658 (I14069,I14001,I14052);
DFFARX1 I_659 (I14069,I2859,I13645,I13634,);
nor I_660 (I14100,I13962,I14035);
nor I_661 (I13622,I13826,I14100);
nor I_662 (I13616,I13962,I14018);
not I_663 (I14172,I2866);
DFFARX1 I_664 (I164600,I2859,I14172,I14198,);
DFFARX1 I_665 (I14198,I2859,I14172,I14215,);
not I_666 (I14223,I14215);
nand I_667 (I14240,I164597,I164591);
and I_668 (I14257,I14240,I164585);
DFFARX1 I_669 (I14257,I2859,I14172,I14283,);
DFFARX1 I_670 (I14283,I2859,I14172,I14164,);
DFFARX1 I_671 (I14283,I2859,I14172,I14155,);
DFFARX1 I_672 (I164573,I2859,I14172,I14328,);
nand I_673 (I14336,I14328,I164582);
not I_674 (I14353,I14336);
nor I_675 (I14152,I14198,I14353);
DFFARX1 I_676 (I164579,I2859,I14172,I14393,);
not I_677 (I14401,I14393);
nor I_678 (I14158,I14401,I14223);
nand I_679 (I14146,I14401,I14336);
nand I_680 (I14446,I164576,I164594);
and I_681 (I14463,I14446,I164573);
DFFARX1 I_682 (I14463,I2859,I14172,I14489,);
nor I_683 (I14497,I14489,I14198);
DFFARX1 I_684 (I14497,I2859,I14172,I14140,);
not I_685 (I14528,I14489);
nor I_686 (I14545,I164588,I164594);
not I_687 (I14562,I14545);
nor I_688 (I14579,I14336,I14562);
nor I_689 (I14596,I14528,I14579);
DFFARX1 I_690 (I14596,I2859,I14172,I14161,);
nor I_691 (I14627,I14489,I14562);
nor I_692 (I14149,I14353,I14627);
nor I_693 (I14143,I14489,I14545);
not I_694 (I14699,I2866);
DFFARX1 I_695 (I138777,I2859,I14699,I14725,);
DFFARX1 I_696 (I14725,I2859,I14699,I14742,);
not I_697 (I14750,I14742);
nand I_698 (I14767,I138774,I138768);
and I_699 (I14784,I14767,I138762);
DFFARX1 I_700 (I14784,I2859,I14699,I14810,);
DFFARX1 I_701 (I14810,I2859,I14699,I14691,);
DFFARX1 I_702 (I14810,I2859,I14699,I14682,);
DFFARX1 I_703 (I138750,I2859,I14699,I14855,);
nand I_704 (I14863,I14855,I138759);
not I_705 (I14880,I14863);
nor I_706 (I14679,I14725,I14880);
DFFARX1 I_707 (I138756,I2859,I14699,I14920,);
not I_708 (I14928,I14920);
nor I_709 (I14685,I14928,I14750);
nand I_710 (I14673,I14928,I14863);
nand I_711 (I14973,I138753,I138771);
and I_712 (I14990,I14973,I138750);
DFFARX1 I_713 (I14990,I2859,I14699,I15016,);
nor I_714 (I15024,I15016,I14725);
DFFARX1 I_715 (I15024,I2859,I14699,I14667,);
not I_716 (I15055,I15016);
nor I_717 (I15072,I138765,I138771);
not I_718 (I15089,I15072);
nor I_719 (I15106,I14863,I15089);
nor I_720 (I15123,I15055,I15106);
DFFARX1 I_721 (I15123,I2859,I14699,I14688,);
nor I_722 (I15154,I15016,I15089);
nor I_723 (I14676,I14880,I15154);
nor I_724 (I14670,I15016,I15072);
not I_725 (I15226,I2866);
DFFARX1 I_726 (I555590,I2859,I15226,I15252,);
DFFARX1 I_727 (I15252,I2859,I15226,I15269,);
not I_728 (I15277,I15269);
nand I_729 (I15294,I555593,I555599);
and I_730 (I15311,I15294,I555608);
DFFARX1 I_731 (I15311,I2859,I15226,I15337,);
DFFARX1 I_732 (I15337,I2859,I15226,I15218,);
DFFARX1 I_733 (I15337,I2859,I15226,I15209,);
DFFARX1 I_734 (I555611,I2859,I15226,I15382,);
nand I_735 (I15390,I15382,I555602);
not I_736 (I15407,I15390);
nor I_737 (I15206,I15252,I15407);
DFFARX1 I_738 (I555590,I2859,I15226,I15447,);
not I_739 (I15455,I15447);
nor I_740 (I15212,I15455,I15277);
nand I_741 (I15200,I15455,I15390);
nand I_742 (I15500,I555617,I555596);
and I_743 (I15517,I15500,I555605);
DFFARX1 I_744 (I15517,I2859,I15226,I15543,);
nor I_745 (I15551,I15543,I15252);
DFFARX1 I_746 (I15551,I2859,I15226,I15194,);
not I_747 (I15582,I15543);
nor I_748 (I15599,I555614,I555596);
not I_749 (I15616,I15599);
nor I_750 (I15633,I15390,I15616);
nor I_751 (I15650,I15582,I15633);
DFFARX1 I_752 (I15650,I2859,I15226,I15215,);
nor I_753 (I15681,I15543,I15616);
nor I_754 (I15203,I15407,I15681);
nor I_755 (I15197,I15543,I15599);
not I_756 (I15753,I2866);
DFFARX1 I_757 (I363754,I2859,I15753,I15779,);
DFFARX1 I_758 (I15779,I2859,I15753,I15796,);
not I_759 (I15804,I15796);
nand I_760 (I15821,I363745,I363766);
and I_761 (I15838,I15821,I363748);
DFFARX1 I_762 (I15838,I2859,I15753,I15864,);
DFFARX1 I_763 (I15864,I2859,I15753,I15745,);
DFFARX1 I_764 (I15864,I2859,I15753,I15736,);
DFFARX1 I_765 (I363748,I2859,I15753,I15909,);
nand I_766 (I15917,I15909,I363763);
not I_767 (I15934,I15917);
nor I_768 (I15733,I15779,I15934);
DFFARX1 I_769 (I363757,I2859,I15753,I15974,);
not I_770 (I15982,I15974);
nor I_771 (I15739,I15982,I15804);
nand I_772 (I15727,I15982,I15917);
nand I_773 (I16027,I363751,I363760);
and I_774 (I16044,I16027,I363745);
DFFARX1 I_775 (I16044,I2859,I15753,I16070,);
nor I_776 (I16078,I16070,I15779);
DFFARX1 I_777 (I16078,I2859,I15753,I15721,);
not I_778 (I16109,I16070);
nor I_779 (I16126,I363751,I363760);
not I_780 (I16143,I16126);
nor I_781 (I16160,I15917,I16143);
nor I_782 (I16177,I16109,I16160);
DFFARX1 I_783 (I16177,I2859,I15753,I15742,);
nor I_784 (I16208,I16070,I16143);
nor I_785 (I15730,I15934,I16208);
nor I_786 (I15724,I16070,I16126);
not I_787 (I16280,I2866);
DFFARX1 I_788 (I167803,I2859,I16280,I16306,);
DFFARX1 I_789 (I16306,I2859,I16280,I16323,);
not I_790 (I16331,I16323);
nand I_791 (I16348,I167803,I167806);
and I_792 (I16365,I16348,I167827);
DFFARX1 I_793 (I16365,I2859,I16280,I16391,);
DFFARX1 I_794 (I16391,I2859,I16280,I16272,);
DFFARX1 I_795 (I16391,I2859,I16280,I16263,);
DFFARX1 I_796 (I167815,I2859,I16280,I16436,);
nand I_797 (I16444,I16436,I167818);
not I_798 (I16461,I16444);
nor I_799 (I16260,I16306,I16461);
DFFARX1 I_800 (I167824,I2859,I16280,I16501,);
not I_801 (I16509,I16501);
nor I_802 (I16266,I16509,I16331);
nand I_803 (I16254,I16509,I16444);
nand I_804 (I16554,I167821,I167809);
and I_805 (I16571,I16554,I167812);
DFFARX1 I_806 (I16571,I2859,I16280,I16597,);
nor I_807 (I16605,I16597,I16306);
DFFARX1 I_808 (I16605,I2859,I16280,I16248,);
not I_809 (I16636,I16597);
nor I_810 (I16653,I167830,I167809);
not I_811 (I16670,I16653);
nor I_812 (I16687,I16444,I16670);
nor I_813 (I16704,I16636,I16687);
DFFARX1 I_814 (I16704,I2859,I16280,I16269,);
nor I_815 (I16735,I16597,I16670);
nor I_816 (I16257,I16461,I16735);
nor I_817 (I16251,I16597,I16653);
not I_818 (I16807,I2866);
DFFARX1 I_819 (I212522,I2859,I16807,I16833,);
DFFARX1 I_820 (I16833,I2859,I16807,I16850,);
not I_821 (I16858,I16850);
nand I_822 (I16875,I212528,I212516);
and I_823 (I16892,I16875,I212513);
DFFARX1 I_824 (I16892,I2859,I16807,I16918,);
DFFARX1 I_825 (I16918,I2859,I16807,I16799,);
DFFARX1 I_826 (I16918,I2859,I16807,I16790,);
DFFARX1 I_827 (I212525,I2859,I16807,I16963,);
nand I_828 (I16971,I16963,I212519);
not I_829 (I16988,I16971);
nor I_830 (I16787,I16833,I16988);
DFFARX1 I_831 (I212537,I2859,I16807,I17028,);
not I_832 (I17036,I17028);
nor I_833 (I16793,I17036,I16858);
nand I_834 (I16781,I17036,I16971);
nand I_835 (I17081,I212531,I212534);
and I_836 (I17098,I17081,I212516);
DFFARX1 I_837 (I17098,I2859,I16807,I17124,);
nor I_838 (I17132,I17124,I16833);
DFFARX1 I_839 (I17132,I2859,I16807,I16775,);
not I_840 (I17163,I17124);
nor I_841 (I17180,I212513,I212534);
not I_842 (I17197,I17180);
nor I_843 (I17214,I16971,I17197);
nor I_844 (I17231,I17163,I17214);
DFFARX1 I_845 (I17231,I2859,I16807,I16796,);
nor I_846 (I17262,I17124,I17197);
nor I_847 (I16784,I16988,I17262);
nor I_848 (I16778,I17124,I17180);
not I_849 (I17334,I2866);
DFFARX1 I_850 (I433740,I2859,I17334,I17360,);
DFFARX1 I_851 (I17360,I2859,I17334,I17377,);
not I_852 (I17385,I17377);
nand I_853 (I17402,I433734,I433755);
and I_854 (I17419,I17402,I433740);
DFFARX1 I_855 (I17419,I2859,I17334,I17445,);
DFFARX1 I_856 (I17445,I2859,I17334,I17326,);
DFFARX1 I_857 (I17445,I2859,I17334,I17317,);
DFFARX1 I_858 (I433737,I2859,I17334,I17490,);
nand I_859 (I17498,I17490,I433746);
not I_860 (I17515,I17498);
nor I_861 (I17314,I17360,I17515);
DFFARX1 I_862 (I433734,I2859,I17334,I17555,);
not I_863 (I17563,I17555);
nor I_864 (I17320,I17563,I17385);
nand I_865 (I17308,I17563,I17498);
nand I_866 (I17608,I433737,I433752);
and I_867 (I17625,I17608,I433743);
DFFARX1 I_868 (I17625,I2859,I17334,I17651,);
nor I_869 (I17659,I17651,I17360);
DFFARX1 I_870 (I17659,I2859,I17334,I17302,);
not I_871 (I17690,I17651);
nor I_872 (I17707,I433749,I433752);
not I_873 (I17724,I17707);
nor I_874 (I17741,I17498,I17724);
nor I_875 (I17758,I17690,I17741);
DFFARX1 I_876 (I17758,I2859,I17334,I17323,);
nor I_877 (I17789,I17651,I17724);
nor I_878 (I17311,I17515,I17789);
nor I_879 (I17305,I17651,I17707);
not I_880 (I17861,I2866);
DFFARX1 I_881 (I146682,I2859,I17861,I17887,);
DFFARX1 I_882 (I17887,I2859,I17861,I17904,);
not I_883 (I17912,I17904);
nand I_884 (I17929,I146679,I146673);
and I_885 (I17946,I17929,I146667);
DFFARX1 I_886 (I17946,I2859,I17861,I17972,);
DFFARX1 I_887 (I17972,I2859,I17861,I17853,);
DFFARX1 I_888 (I17972,I2859,I17861,I17844,);
DFFARX1 I_889 (I146655,I2859,I17861,I18017,);
nand I_890 (I18025,I18017,I146664);
not I_891 (I18042,I18025);
nor I_892 (I17841,I17887,I18042);
DFFARX1 I_893 (I146661,I2859,I17861,I18082,);
not I_894 (I18090,I18082);
nor I_895 (I17847,I18090,I17912);
nand I_896 (I17835,I18090,I18025);
nand I_897 (I18135,I146658,I146676);
and I_898 (I18152,I18135,I146655);
DFFARX1 I_899 (I18152,I2859,I17861,I18178,);
nor I_900 (I18186,I18178,I17887);
DFFARX1 I_901 (I18186,I2859,I17861,I17829,);
not I_902 (I18217,I18178);
nor I_903 (I18234,I146670,I146676);
not I_904 (I18251,I18234);
nor I_905 (I18268,I18025,I18251);
nor I_906 (I18285,I18217,I18268);
DFFARX1 I_907 (I18285,I2859,I17861,I17850,);
nor I_908 (I18316,I18178,I18251);
nor I_909 (I17838,I18042,I18316);
nor I_910 (I17832,I18178,I18234);
not I_911 (I18388,I2866);
DFFARX1 I_912 (I319364,I2859,I18388,I18414,);
DFFARX1 I_913 (I18414,I2859,I18388,I18431,);
not I_914 (I18439,I18431);
nand I_915 (I18456,I319379,I319382);
and I_916 (I18473,I18456,I319361);
DFFARX1 I_917 (I18473,I2859,I18388,I18499,);
DFFARX1 I_918 (I18499,I2859,I18388,I18380,);
DFFARX1 I_919 (I18499,I2859,I18388,I18371,);
DFFARX1 I_920 (I319367,I2859,I18388,I18544,);
nand I_921 (I18552,I18544,I319373);
not I_922 (I18569,I18552);
nor I_923 (I18368,I18414,I18569);
DFFARX1 I_924 (I319361,I2859,I18388,I18609,);
not I_925 (I18617,I18609);
nor I_926 (I18374,I18617,I18439);
nand I_927 (I18362,I18617,I18552);
nand I_928 (I18662,I319376,I319358);
and I_929 (I18679,I18662,I319370);
DFFARX1 I_930 (I18679,I2859,I18388,I18705,);
nor I_931 (I18713,I18705,I18414);
DFFARX1 I_932 (I18713,I2859,I18388,I18356,);
not I_933 (I18744,I18705);
nor I_934 (I18761,I319358,I319358);
not I_935 (I18778,I18761);
nor I_936 (I18795,I18552,I18778);
nor I_937 (I18812,I18744,I18795);
DFFARX1 I_938 (I18812,I2859,I18388,I18377,);
nor I_939 (I18843,I18705,I18778);
nor I_940 (I18365,I18569,I18843);
nor I_941 (I18359,I18705,I18761);
not I_942 (I18915,I2866);
DFFARX1 I_943 (I433179,I2859,I18915,I18941,);
DFFARX1 I_944 (I18941,I2859,I18915,I18958,);
not I_945 (I18966,I18958);
nand I_946 (I18983,I433173,I433194);
and I_947 (I19000,I18983,I433179);
DFFARX1 I_948 (I19000,I2859,I18915,I19026,);
DFFARX1 I_949 (I19026,I2859,I18915,I18907,);
DFFARX1 I_950 (I19026,I2859,I18915,I18898,);
DFFARX1 I_951 (I433176,I2859,I18915,I19071,);
nand I_952 (I19079,I19071,I433185);
not I_953 (I19096,I19079);
nor I_954 (I18895,I18941,I19096);
DFFARX1 I_955 (I433173,I2859,I18915,I19136,);
not I_956 (I19144,I19136);
nor I_957 (I18901,I19144,I18966);
nand I_958 (I18889,I19144,I19079);
nand I_959 (I19189,I433176,I433191);
and I_960 (I19206,I19189,I433182);
DFFARX1 I_961 (I19206,I2859,I18915,I19232,);
nor I_962 (I19240,I19232,I18941);
DFFARX1 I_963 (I19240,I2859,I18915,I18883,);
not I_964 (I19271,I19232);
nor I_965 (I19288,I433188,I433191);
not I_966 (I19305,I19288);
nor I_967 (I19322,I19079,I19305);
nor I_968 (I19339,I19271,I19322);
DFFARX1 I_969 (I19339,I2859,I18915,I18904,);
nor I_970 (I19370,I19232,I19305);
nor I_971 (I18892,I19096,I19370);
nor I_972 (I18886,I19232,I19288);
not I_973 (I19442,I2866);
DFFARX1 I_974 (I279482,I2859,I19442,I19468,);
DFFARX1 I_975 (I19468,I2859,I19442,I19485,);
not I_976 (I19493,I19485);
nand I_977 (I19510,I279497,I279500);
and I_978 (I19527,I19510,I279479);
DFFARX1 I_979 (I19527,I2859,I19442,I19553,);
DFFARX1 I_980 (I19553,I2859,I19442,I19434,);
DFFARX1 I_981 (I19553,I2859,I19442,I19425,);
DFFARX1 I_982 (I279485,I2859,I19442,I19598,);
nand I_983 (I19606,I19598,I279491);
not I_984 (I19623,I19606);
nor I_985 (I19422,I19468,I19623);
DFFARX1 I_986 (I279479,I2859,I19442,I19663,);
not I_987 (I19671,I19663);
nor I_988 (I19428,I19671,I19493);
nand I_989 (I19416,I19671,I19606);
nand I_990 (I19716,I279494,I279476);
and I_991 (I19733,I19716,I279488);
DFFARX1 I_992 (I19733,I2859,I19442,I19759,);
nor I_993 (I19767,I19759,I19468);
DFFARX1 I_994 (I19767,I2859,I19442,I19410,);
not I_995 (I19798,I19759);
nor I_996 (I19815,I279476,I279476);
not I_997 (I19832,I19815);
nor I_998 (I19849,I19606,I19832);
nor I_999 (I19866,I19798,I19849);
DFFARX1 I_1000 (I19866,I2859,I19442,I19431,);
nor I_1001 (I19897,I19759,I19832);
nor I_1002 (I19419,I19623,I19897);
nor I_1003 (I19413,I19759,I19815);
not I_1004 (I19969,I2866);
DFFARX1 I_1005 (I202619,I2859,I19969,I19995,);
DFFARX1 I_1006 (I19995,I2859,I19969,I20012,);
not I_1007 (I20020,I20012);
nand I_1008 (I20037,I202619,I202622);
and I_1009 (I20054,I20037,I202643);
DFFARX1 I_1010 (I20054,I2859,I19969,I20080,);
DFFARX1 I_1011 (I20080,I2859,I19969,I19961,);
DFFARX1 I_1012 (I20080,I2859,I19969,I19952,);
DFFARX1 I_1013 (I202631,I2859,I19969,I20125,);
nand I_1014 (I20133,I20125,I202634);
not I_1015 (I20150,I20133);
nor I_1016 (I19949,I19995,I20150);
DFFARX1 I_1017 (I202640,I2859,I19969,I20190,);
not I_1018 (I20198,I20190);
nor I_1019 (I19955,I20198,I20020);
nand I_1020 (I19943,I20198,I20133);
nand I_1021 (I20243,I202637,I202625);
and I_1022 (I20260,I20243,I202628);
DFFARX1 I_1023 (I20260,I2859,I19969,I20286,);
nor I_1024 (I20294,I20286,I19995);
DFFARX1 I_1025 (I20294,I2859,I19969,I19937,);
not I_1026 (I20325,I20286);
nor I_1027 (I20342,I202646,I202625);
not I_1028 (I20359,I20342);
nor I_1029 (I20376,I20133,I20359);
nor I_1030 (I20393,I20325,I20376);
DFFARX1 I_1031 (I20393,I2859,I19969,I19958,);
nor I_1032 (I20424,I20286,I20359);
nor I_1033 (I19946,I20150,I20424);
nor I_1034 (I19940,I20286,I20342);
not I_1035 (I20496,I2866);
DFFARX1 I_1036 (I502074,I2859,I20496,I20522,);
DFFARX1 I_1037 (I20522,I2859,I20496,I20539,);
not I_1038 (I20547,I20539);
nand I_1039 (I20564,I502092,I502086);
and I_1040 (I20581,I20564,I502095);
DFFARX1 I_1041 (I20581,I2859,I20496,I20607,);
DFFARX1 I_1042 (I20607,I2859,I20496,I20488,);
DFFARX1 I_1043 (I20607,I2859,I20496,I20479,);
DFFARX1 I_1044 (I502080,I2859,I20496,I20652,);
nand I_1045 (I20660,I20652,I502089);
not I_1046 (I20677,I20660);
nor I_1047 (I20476,I20522,I20677);
DFFARX1 I_1048 (I502077,I2859,I20496,I20717,);
not I_1049 (I20725,I20717);
nor I_1050 (I20482,I20725,I20547);
nand I_1051 (I20470,I20725,I20660);
nand I_1052 (I20770,I502098,I502083);
and I_1053 (I20787,I20770,I502077);
DFFARX1 I_1054 (I20787,I2859,I20496,I20813,);
nor I_1055 (I20821,I20813,I20522);
DFFARX1 I_1056 (I20821,I2859,I20496,I20464,);
not I_1057 (I20852,I20813);
nor I_1058 (I20869,I502074,I502083);
not I_1059 (I20886,I20869);
nor I_1060 (I20903,I20660,I20886);
nor I_1061 (I20920,I20852,I20903);
DFFARX1 I_1062 (I20920,I2859,I20496,I20485,);
nor I_1063 (I20951,I20813,I20886);
nor I_1064 (I20473,I20677,I20951);
nor I_1065 (I20467,I20813,I20869);
not I_1066 (I21023,I2866);
DFFARX1 I_1067 (I62585,I2859,I21023,I21049,);
not I_1068 (I21057,I21049);
nand I_1069 (I21074,I62579,I62573);
and I_1070 (I21091,I21074,I62594);
DFFARX1 I_1071 (I21091,I2859,I21023,I21117,);
DFFARX1 I_1072 (I62591,I2859,I21023,I21134,);
and I_1073 (I21142,I21134,I62588);
nor I_1074 (I21159,I21117,I21142);
DFFARX1 I_1075 (I21159,I2859,I21023,I20991,);
nand I_1076 (I21190,I21134,I62588);
nand I_1077 (I21207,I21057,I21190);
not I_1078 (I21003,I21207);
DFFARX1 I_1079 (I62573,I2859,I21023,I21247,);
DFFARX1 I_1080 (I21247,I2859,I21023,I21012,);
nand I_1081 (I21269,I62576,I62576);
and I_1082 (I21286,I21269,I62597);
DFFARX1 I_1083 (I21286,I2859,I21023,I21312,);
DFFARX1 I_1084 (I21312,I2859,I21023,I21329,);
not I_1085 (I21015,I21329);
not I_1086 (I21351,I21312);
nand I_1087 (I21000,I21351,I21190);
nor I_1088 (I21382,I62582,I62576);
not I_1089 (I21399,I21382);
nor I_1090 (I21416,I21351,I21399);
nor I_1091 (I21433,I21057,I21416);
DFFARX1 I_1092 (I21433,I2859,I21023,I21009,);
nor I_1093 (I21464,I21117,I21399);
nor I_1094 (I20997,I21312,I21464);
nor I_1095 (I21006,I21247,I21382);
nor I_1096 (I20994,I21117,I21382);
not I_1097 (I21550,I2866);
DFFARX1 I_1098 (I459886,I2859,I21550,I21576,);
not I_1099 (I21584,I21576);
nand I_1100 (I21601,I459901,I459880);
and I_1101 (I21618,I21601,I459883);
DFFARX1 I_1102 (I21618,I2859,I21550,I21644,);
DFFARX1 I_1103 (I459904,I2859,I21550,I21661,);
and I_1104 (I21669,I21661,I459883);
nor I_1105 (I21686,I21644,I21669);
DFFARX1 I_1106 (I21686,I2859,I21550,I21518,);
nand I_1107 (I21717,I21661,I459883);
nand I_1108 (I21734,I21584,I21717);
not I_1109 (I21530,I21734);
DFFARX1 I_1110 (I459880,I2859,I21550,I21774,);
DFFARX1 I_1111 (I21774,I2859,I21550,I21539,);
nand I_1112 (I21796,I459892,I459889);
and I_1113 (I21813,I21796,I459895);
DFFARX1 I_1114 (I21813,I2859,I21550,I21839,);
DFFARX1 I_1115 (I21839,I2859,I21550,I21856,);
not I_1116 (I21542,I21856);
not I_1117 (I21878,I21839);
nand I_1118 (I21527,I21878,I21717);
nor I_1119 (I21909,I459898,I459889);
not I_1120 (I21926,I21909);
nor I_1121 (I21943,I21878,I21926);
nor I_1122 (I21960,I21584,I21943);
DFFARX1 I_1123 (I21960,I2859,I21550,I21536,);
nor I_1124 (I21991,I21644,I21926);
nor I_1125 (I21524,I21839,I21991);
nor I_1126 (I21533,I21774,I21909);
nor I_1127 (I21521,I21644,I21909);
not I_1128 (I22077,I2866);
DFFARX1 I_1129 (I91740,I2859,I22077,I22103,);
not I_1130 (I22111,I22103);
nand I_1131 (I22128,I91734,I91728);
and I_1132 (I22145,I22128,I91749);
DFFARX1 I_1133 (I22145,I2859,I22077,I22171,);
DFFARX1 I_1134 (I91746,I2859,I22077,I22188,);
and I_1135 (I22196,I22188,I91743);
nor I_1136 (I22213,I22171,I22196);
DFFARX1 I_1137 (I22213,I2859,I22077,I22045,);
nand I_1138 (I22244,I22188,I91743);
nand I_1139 (I22261,I22111,I22244);
not I_1140 (I22057,I22261);
DFFARX1 I_1141 (I91728,I2859,I22077,I22301,);
DFFARX1 I_1142 (I22301,I2859,I22077,I22066,);
nand I_1143 (I22323,I91731,I91731);
and I_1144 (I22340,I22323,I91752);
DFFARX1 I_1145 (I22340,I2859,I22077,I22366,);
DFFARX1 I_1146 (I22366,I2859,I22077,I22383,);
not I_1147 (I22069,I22383);
not I_1148 (I22405,I22366);
nand I_1149 (I22054,I22405,I22244);
nor I_1150 (I22436,I91737,I91731);
not I_1151 (I22453,I22436);
nor I_1152 (I22470,I22405,I22453);
nor I_1153 (I22487,I22111,I22470);
DFFARX1 I_1154 (I22487,I2859,I22077,I22063,);
nor I_1155 (I22518,I22171,I22453);
nor I_1156 (I22051,I22366,I22518);
nor I_1157 (I22060,I22301,I22436);
nor I_1158 (I22048,I22171,I22436);
not I_1159 (I22604,I2866);
DFFARX1 I_1160 (I70915,I2859,I22604,I22630,);
not I_1161 (I22638,I22630);
nand I_1162 (I22655,I70909,I70903);
and I_1163 (I22672,I22655,I70924);
DFFARX1 I_1164 (I22672,I2859,I22604,I22698,);
DFFARX1 I_1165 (I70921,I2859,I22604,I22715,);
and I_1166 (I22723,I22715,I70918);
nor I_1167 (I22740,I22698,I22723);
DFFARX1 I_1168 (I22740,I2859,I22604,I22572,);
nand I_1169 (I22771,I22715,I70918);
nand I_1170 (I22788,I22638,I22771);
not I_1171 (I22584,I22788);
DFFARX1 I_1172 (I70903,I2859,I22604,I22828,);
DFFARX1 I_1173 (I22828,I2859,I22604,I22593,);
nand I_1174 (I22850,I70906,I70906);
and I_1175 (I22867,I22850,I70927);
DFFARX1 I_1176 (I22867,I2859,I22604,I22893,);
DFFARX1 I_1177 (I22893,I2859,I22604,I22910,);
not I_1178 (I22596,I22910);
not I_1179 (I22932,I22893);
nand I_1180 (I22581,I22932,I22771);
nor I_1181 (I22963,I70912,I70906);
not I_1182 (I22980,I22963);
nor I_1183 (I22997,I22932,I22980);
nor I_1184 (I23014,I22638,I22997);
DFFARX1 I_1185 (I23014,I2859,I22604,I22590,);
nor I_1186 (I23045,I22698,I22980);
nor I_1187 (I22578,I22893,I23045);
nor I_1188 (I22587,I22828,I22963);
nor I_1189 (I22575,I22698,I22963);
not I_1190 (I23131,I2866);
DFFARX1 I_1191 (I265038,I2859,I23131,I23157,);
not I_1192 (I23165,I23157);
nand I_1193 (I23182,I265029,I265047);
and I_1194 (I23199,I23182,I265026);
DFFARX1 I_1195 (I23199,I2859,I23131,I23225,);
DFFARX1 I_1196 (I265029,I2859,I23131,I23242,);
and I_1197 (I23250,I23242,I265032);
nor I_1198 (I23267,I23225,I23250);
DFFARX1 I_1199 (I23267,I2859,I23131,I23099,);
nand I_1200 (I23298,I23242,I265032);
nand I_1201 (I23315,I23165,I23298);
not I_1202 (I23111,I23315);
DFFARX1 I_1203 (I265026,I2859,I23131,I23355,);
DFFARX1 I_1204 (I23355,I2859,I23131,I23120,);
nand I_1205 (I23377,I265044,I265035);
and I_1206 (I23394,I23377,I265050);
DFFARX1 I_1207 (I23394,I2859,I23131,I23420,);
DFFARX1 I_1208 (I23420,I2859,I23131,I23437,);
not I_1209 (I23123,I23437);
not I_1210 (I23459,I23420);
nand I_1211 (I23108,I23459,I23298);
nor I_1212 (I23490,I265041,I265035);
not I_1213 (I23507,I23490);
nor I_1214 (I23524,I23459,I23507);
nor I_1215 (I23541,I23165,I23524);
DFFARX1 I_1216 (I23541,I2859,I23131,I23117,);
nor I_1217 (I23572,I23225,I23507);
nor I_1218 (I23105,I23420,I23572);
nor I_1219 (I23114,I23355,I23490);
nor I_1220 (I23102,I23225,I23490);
not I_1221 (I23658,I2866);
DFFARX1 I_1222 (I222036,I2859,I23658,I23684,);
not I_1223 (I23692,I23684);
nand I_1224 (I23709,I222057,I222051);
and I_1225 (I23726,I23709,I222033);
DFFARX1 I_1226 (I23726,I2859,I23658,I23752,);
DFFARX1 I_1227 (I222036,I2859,I23658,I23769,);
and I_1228 (I23777,I23769,I222045);
nor I_1229 (I23794,I23752,I23777);
DFFARX1 I_1230 (I23794,I2859,I23658,I23626,);
nand I_1231 (I23825,I23769,I222045);
nand I_1232 (I23842,I23692,I23825);
not I_1233 (I23638,I23842);
DFFARX1 I_1234 (I222042,I2859,I23658,I23882,);
DFFARX1 I_1235 (I23882,I2859,I23658,I23647,);
nand I_1236 (I23904,I222048,I222039);
and I_1237 (I23921,I23904,I222033);
DFFARX1 I_1238 (I23921,I2859,I23658,I23947,);
DFFARX1 I_1239 (I23947,I2859,I23658,I23964,);
not I_1240 (I23650,I23964);
not I_1241 (I23986,I23947);
nand I_1242 (I23635,I23986,I23825);
nor I_1243 (I24017,I222054,I222039);
not I_1244 (I24034,I24017);
nor I_1245 (I24051,I23986,I24034);
nor I_1246 (I24068,I23692,I24051);
DFFARX1 I_1247 (I24068,I2859,I23658,I23644,);
nor I_1248 (I24099,I23752,I24034);
nor I_1249 (I23632,I23947,I24099);
nor I_1250 (I23641,I23882,I24017);
nor I_1251 (I23629,I23752,I24017);
not I_1252 (I24185,I2866);
DFFARX1 I_1253 (I514048,I2859,I24185,I24211,);
not I_1254 (I24219,I24211);
nand I_1255 (I24236,I514042,I514063);
and I_1256 (I24253,I24236,I514054);
DFFARX1 I_1257 (I24253,I2859,I24185,I24279,);
DFFARX1 I_1258 (I514045,I2859,I24185,I24296,);
and I_1259 (I24304,I24296,I514057);
nor I_1260 (I24321,I24279,I24304);
DFFARX1 I_1261 (I24321,I2859,I24185,I24153,);
nand I_1262 (I24352,I24296,I514057);
nand I_1263 (I24369,I24219,I24352);
not I_1264 (I24165,I24369);
DFFARX1 I_1265 (I514045,I2859,I24185,I24409,);
DFFARX1 I_1266 (I24409,I2859,I24185,I24174,);
nand I_1267 (I24431,I514066,I514051);
and I_1268 (I24448,I24431,I514042);
DFFARX1 I_1269 (I24448,I2859,I24185,I24474,);
DFFARX1 I_1270 (I24474,I2859,I24185,I24491,);
not I_1271 (I24177,I24491);
not I_1272 (I24513,I24474);
nand I_1273 (I24162,I24513,I24352);
nor I_1274 (I24544,I514060,I514051);
not I_1275 (I24561,I24544);
nor I_1276 (I24578,I24513,I24561);
nor I_1277 (I24595,I24219,I24578);
DFFARX1 I_1278 (I24595,I2859,I24185,I24171,);
nor I_1279 (I24626,I24279,I24561);
nor I_1280 (I24159,I24474,I24626);
nor I_1281 (I24168,I24409,I24544);
nor I_1282 (I24156,I24279,I24544);
not I_1283 (I24712,I2866);
DFFARX1 I_1284 (I102450,I2859,I24712,I24738,);
not I_1285 (I24746,I24738);
nand I_1286 (I24763,I102444,I102438);
and I_1287 (I24780,I24763,I102459);
DFFARX1 I_1288 (I24780,I2859,I24712,I24806,);
DFFARX1 I_1289 (I102456,I2859,I24712,I24823,);
and I_1290 (I24831,I24823,I102453);
nor I_1291 (I24848,I24806,I24831);
DFFARX1 I_1292 (I24848,I2859,I24712,I24680,);
nand I_1293 (I24879,I24823,I102453);
nand I_1294 (I24896,I24746,I24879);
not I_1295 (I24692,I24896);
DFFARX1 I_1296 (I102438,I2859,I24712,I24936,);
DFFARX1 I_1297 (I24936,I2859,I24712,I24701,);
nand I_1298 (I24958,I102441,I102441);
and I_1299 (I24975,I24958,I102462);
DFFARX1 I_1300 (I24975,I2859,I24712,I25001,);
DFFARX1 I_1301 (I25001,I2859,I24712,I25018,);
not I_1302 (I24704,I25018);
not I_1303 (I25040,I25001);
nand I_1304 (I24689,I25040,I24879);
nor I_1305 (I25071,I102447,I102441);
not I_1306 (I25088,I25071);
nor I_1307 (I25105,I25040,I25088);
nor I_1308 (I25122,I24746,I25105);
DFFARX1 I_1309 (I25122,I2859,I24712,I24698,);
nor I_1310 (I25153,I24806,I25088);
nor I_1311 (I24686,I25001,I25153);
nor I_1312 (I24695,I24936,I25071);
nor I_1313 (I24683,I24806,I25071);
not I_1314 (I25239,I2866);
DFFARX1 I_1315 (I2620,I2859,I25239,I25265,);
not I_1316 (I25273,I25265);
nand I_1317 (I25290,I1916,I2820);
and I_1318 (I25307,I25290,I2324);
DFFARX1 I_1319 (I25307,I2859,I25239,I25333,);
DFFARX1 I_1320 (I2700,I2859,I25239,I25350,);
and I_1321 (I25358,I25350,I2284);
nor I_1322 (I25375,I25333,I25358);
DFFARX1 I_1323 (I25375,I2859,I25239,I25207,);
nand I_1324 (I25406,I25350,I2284);
nand I_1325 (I25423,I25273,I25406);
not I_1326 (I25219,I25423);
DFFARX1 I_1327 (I1996,I2859,I25239,I25463,);
DFFARX1 I_1328 (I25463,I2859,I25239,I25228,);
nand I_1329 (I25485,I1644,I2452);
and I_1330 (I25502,I25485,I2388);
DFFARX1 I_1331 (I25502,I2859,I25239,I25528,);
DFFARX1 I_1332 (I25528,I2859,I25239,I25545,);
not I_1333 (I25231,I25545);
not I_1334 (I25567,I25528);
nand I_1335 (I25216,I25567,I25406);
nor I_1336 (I25598,I2404,I2452);
not I_1337 (I25615,I25598);
nor I_1338 (I25632,I25567,I25615);
nor I_1339 (I25649,I25273,I25632);
DFFARX1 I_1340 (I25649,I2859,I25239,I25225,);
nor I_1341 (I25680,I25333,I25615);
nor I_1342 (I25213,I25528,I25680);
nor I_1343 (I25222,I25463,I25598);
nor I_1344 (I25210,I25333,I25598);
not I_1345 (I25766,I2866);
DFFARX1 I_1346 (I366916,I2859,I25766,I25792,);
not I_1347 (I25800,I25792);
nand I_1348 (I25817,I366913,I366928);
and I_1349 (I25834,I25817,I366910);
DFFARX1 I_1350 (I25834,I2859,I25766,I25860,);
DFFARX1 I_1351 (I366907,I2859,I25766,I25877,);
and I_1352 (I25885,I25877,I366907);
nor I_1353 (I25902,I25860,I25885);
DFFARX1 I_1354 (I25902,I2859,I25766,I25734,);
nand I_1355 (I25933,I25877,I366907);
nand I_1356 (I25950,I25800,I25933);
not I_1357 (I25746,I25950);
DFFARX1 I_1358 (I366910,I2859,I25766,I25990,);
DFFARX1 I_1359 (I25990,I2859,I25766,I25755,);
nand I_1360 (I26012,I366922,I366913);
and I_1361 (I26029,I26012,I366925);
DFFARX1 I_1362 (I26029,I2859,I25766,I26055,);
DFFARX1 I_1363 (I26055,I2859,I25766,I26072,);
not I_1364 (I25758,I26072);
not I_1365 (I26094,I26055);
nand I_1366 (I25743,I26094,I25933);
nor I_1367 (I26125,I366919,I366913);
not I_1368 (I26142,I26125);
nor I_1369 (I26159,I26094,I26142);
nor I_1370 (I26176,I25800,I26159);
DFFARX1 I_1371 (I26176,I2859,I25766,I25752,);
nor I_1372 (I26207,I25860,I26142);
nor I_1373 (I25740,I26055,I26207);
nor I_1374 (I25749,I25990,I26125);
nor I_1375 (I25737,I25860,I26125);
not I_1376 (I26293,I2866);
DFFARX1 I_1377 (I373767,I2859,I26293,I26319,);
not I_1378 (I26327,I26319);
nand I_1379 (I26344,I373764,I373779);
and I_1380 (I26361,I26344,I373761);
DFFARX1 I_1381 (I26361,I2859,I26293,I26387,);
DFFARX1 I_1382 (I373758,I2859,I26293,I26404,);
and I_1383 (I26412,I26404,I373758);
nor I_1384 (I26429,I26387,I26412);
DFFARX1 I_1385 (I26429,I2859,I26293,I26261,);
nand I_1386 (I26460,I26404,I373758);
nand I_1387 (I26477,I26327,I26460);
not I_1388 (I26273,I26477);
DFFARX1 I_1389 (I373761,I2859,I26293,I26517,);
DFFARX1 I_1390 (I26517,I2859,I26293,I26282,);
nand I_1391 (I26539,I373773,I373764);
and I_1392 (I26556,I26539,I373776);
DFFARX1 I_1393 (I26556,I2859,I26293,I26582,);
DFFARX1 I_1394 (I26582,I2859,I26293,I26599,);
not I_1395 (I26285,I26599);
not I_1396 (I26621,I26582);
nand I_1397 (I26270,I26621,I26460);
nor I_1398 (I26652,I373770,I373764);
not I_1399 (I26669,I26652);
nor I_1400 (I26686,I26621,I26669);
nor I_1401 (I26703,I26327,I26686);
DFFARX1 I_1402 (I26703,I2859,I26293,I26279,);
nor I_1403 (I26734,I26387,I26669);
nor I_1404 (I26267,I26582,I26734);
nor I_1405 (I26276,I26517,I26652);
nor I_1406 (I26264,I26387,I26652);
not I_1407 (I26820,I2866);
DFFARX1 I_1408 (I535564,I2859,I26820,I26846,);
not I_1409 (I26854,I26846);
nand I_1410 (I26871,I535570,I535588);
and I_1411 (I26888,I26871,I535585);
DFFARX1 I_1412 (I26888,I2859,I26820,I26914,);
DFFARX1 I_1413 (I535582,I2859,I26820,I26931,);
and I_1414 (I26939,I26931,I535576);
nor I_1415 (I26956,I26914,I26939);
DFFARX1 I_1416 (I26956,I2859,I26820,I26788,);
nand I_1417 (I26987,I26931,I535576);
nand I_1418 (I27004,I26854,I26987);
not I_1419 (I26800,I27004);
DFFARX1 I_1420 (I535564,I2859,I26820,I27044,);
DFFARX1 I_1421 (I27044,I2859,I26820,I26809,);
nand I_1422 (I27066,I535579,I535567);
and I_1423 (I27083,I27066,I535591);
DFFARX1 I_1424 (I27083,I2859,I26820,I27109,);
DFFARX1 I_1425 (I27109,I2859,I26820,I27126,);
not I_1426 (I26812,I27126);
not I_1427 (I27148,I27109);
nand I_1428 (I26797,I27148,I26987);
nor I_1429 (I27179,I535573,I535567);
not I_1430 (I27196,I27179);
nor I_1431 (I27213,I27148,I27196);
nor I_1432 (I27230,I26854,I27213);
DFFARX1 I_1433 (I27230,I2859,I26820,I26806,);
nor I_1434 (I27261,I26914,I27196);
nor I_1435 (I26794,I27109,I27261);
nor I_1436 (I26803,I27044,I27179);
nor I_1437 (I26791,I26914,I27179);
not I_1438 (I27347,I2866);
DFFARX1 I_1439 (I83410,I2859,I27347,I27373,);
not I_1440 (I27381,I27373);
nand I_1441 (I27398,I83404,I83398);
and I_1442 (I27415,I27398,I83419);
DFFARX1 I_1443 (I27415,I2859,I27347,I27441,);
DFFARX1 I_1444 (I83416,I2859,I27347,I27458,);
and I_1445 (I27466,I27458,I83413);
nor I_1446 (I27483,I27441,I27466);
DFFARX1 I_1447 (I27483,I2859,I27347,I27315,);
nand I_1448 (I27514,I27458,I83413);
nand I_1449 (I27531,I27381,I27514);
not I_1450 (I27327,I27531);
DFFARX1 I_1451 (I83398,I2859,I27347,I27571,);
DFFARX1 I_1452 (I27571,I2859,I27347,I27336,);
nand I_1453 (I27593,I83401,I83401);
and I_1454 (I27610,I27593,I83422);
DFFARX1 I_1455 (I27610,I2859,I27347,I27636,);
DFFARX1 I_1456 (I27636,I2859,I27347,I27653,);
not I_1457 (I27339,I27653);
not I_1458 (I27675,I27636);
nand I_1459 (I27324,I27675,I27514);
nor I_1460 (I27706,I83407,I83401);
not I_1461 (I27723,I27706);
nor I_1462 (I27740,I27675,I27723);
nor I_1463 (I27757,I27381,I27740);
DFFARX1 I_1464 (I27757,I2859,I27347,I27333,);
nor I_1465 (I27788,I27441,I27723);
nor I_1466 (I27321,I27636,I27788);
nor I_1467 (I27330,I27571,I27706);
nor I_1468 (I27318,I27441,I27706);
not I_1469 (I27874,I2866);
DFFARX1 I_1470 (I544297,I2859,I27874,I27900,);
not I_1471 (I27908,I27900);
nand I_1472 (I27925,I544291,I544312);
and I_1473 (I27942,I27925,I544288);
DFFARX1 I_1474 (I27942,I2859,I27874,I27968,);
DFFARX1 I_1475 (I544309,I2859,I27874,I27985,);
and I_1476 (I27993,I27985,I544306);
nor I_1477 (I28010,I27968,I27993);
DFFARX1 I_1478 (I28010,I2859,I27874,I27842,);
nand I_1479 (I28041,I27985,I544306);
nand I_1480 (I28058,I27908,I28041);
not I_1481 (I27854,I28058);
DFFARX1 I_1482 (I544294,I2859,I27874,I28098,);
DFFARX1 I_1483 (I28098,I2859,I27874,I27863,);
nand I_1484 (I28120,I544303,I544300);
and I_1485 (I28137,I28120,I544285);
DFFARX1 I_1486 (I28137,I2859,I27874,I28163,);
DFFARX1 I_1487 (I28163,I2859,I27874,I28180,);
not I_1488 (I27866,I28180);
not I_1489 (I28202,I28163);
nand I_1490 (I27851,I28202,I28041);
nor I_1491 (I28233,I544285,I544300);
not I_1492 (I28250,I28233);
nor I_1493 (I28267,I28202,I28250);
nor I_1494 (I28284,I27908,I28267);
DFFARX1 I_1495 (I28284,I2859,I27874,I27860,);
nor I_1496 (I28315,I27968,I28250);
nor I_1497 (I27848,I28163,I28315);
nor I_1498 (I27857,I28098,I28233);
nor I_1499 (I27845,I27968,I28233);
not I_1500 (I28401,I2866);
DFFARX1 I_1501 (I115589,I2859,I28401,I28427,);
not I_1502 (I28435,I28427);
nand I_1503 (I28452,I115571,I115586);
and I_1504 (I28469,I28452,I115562);
DFFARX1 I_1505 (I28469,I2859,I28401,I28495,);
DFFARX1 I_1506 (I115565,I2859,I28401,I28512,);
and I_1507 (I28520,I28512,I115580);
nor I_1508 (I28537,I28495,I28520);
DFFARX1 I_1509 (I28537,I2859,I28401,I28369,);
nand I_1510 (I28568,I28512,I115580);
nand I_1511 (I28585,I28435,I28568);
not I_1512 (I28381,I28585);
DFFARX1 I_1513 (I115583,I2859,I28401,I28625,);
DFFARX1 I_1514 (I28625,I2859,I28401,I28390,);
nand I_1515 (I28647,I115562,I115574);
and I_1516 (I28664,I28647,I115568);
DFFARX1 I_1517 (I28664,I2859,I28401,I28690,);
DFFARX1 I_1518 (I28690,I2859,I28401,I28707,);
not I_1519 (I28393,I28707);
not I_1520 (I28729,I28690);
nand I_1521 (I28378,I28729,I28568);
nor I_1522 (I28760,I115577,I115574);
not I_1523 (I28777,I28760);
nor I_1524 (I28794,I28729,I28777);
nor I_1525 (I28811,I28435,I28794);
DFFARX1 I_1526 (I28811,I2859,I28401,I28387,);
nor I_1527 (I28842,I28495,I28777);
nor I_1528 (I28375,I28690,I28842);
nor I_1529 (I28384,I28625,I28760);
nor I_1530 (I28372,I28495,I28760);
not I_1531 (I28928,I2866);
DFFARX1 I_1532 (I306654,I2859,I28928,I28954,);
not I_1533 (I28962,I28954);
nand I_1534 (I28979,I306645,I306663);
and I_1535 (I28996,I28979,I306642);
DFFARX1 I_1536 (I28996,I2859,I28928,I29022,);
DFFARX1 I_1537 (I306645,I2859,I28928,I29039,);
and I_1538 (I29047,I29039,I306648);
nor I_1539 (I29064,I29022,I29047);
DFFARX1 I_1540 (I29064,I2859,I28928,I28896,);
nand I_1541 (I29095,I29039,I306648);
nand I_1542 (I29112,I28962,I29095);
not I_1543 (I28908,I29112);
DFFARX1 I_1544 (I306642,I2859,I28928,I29152,);
DFFARX1 I_1545 (I29152,I2859,I28928,I28917,);
nand I_1546 (I29174,I306660,I306651);
and I_1547 (I29191,I29174,I306666);
DFFARX1 I_1548 (I29191,I2859,I28928,I29217,);
DFFARX1 I_1549 (I29217,I2859,I28928,I29234,);
not I_1550 (I28920,I29234);
not I_1551 (I29256,I29217);
nand I_1552 (I28905,I29256,I29095);
nor I_1553 (I29287,I306657,I306651);
not I_1554 (I29304,I29287);
nor I_1555 (I29321,I29256,I29304);
nor I_1556 (I29338,I28962,I29321);
DFFARX1 I_1557 (I29338,I2859,I28928,I28914,);
nor I_1558 (I29369,I29022,I29304);
nor I_1559 (I28902,I29217,I29369);
nor I_1560 (I28911,I29152,I29287);
nor I_1561 (I28899,I29022,I29287);
not I_1562 (I29455,I2866);
DFFARX1 I_1563 (I121386,I2859,I29455,I29481,);
not I_1564 (I29489,I29481);
nand I_1565 (I29506,I121368,I121383);
and I_1566 (I29523,I29506,I121359);
DFFARX1 I_1567 (I29523,I2859,I29455,I29549,);
DFFARX1 I_1568 (I121362,I2859,I29455,I29566,);
and I_1569 (I29574,I29566,I121377);
nor I_1570 (I29591,I29549,I29574);
DFFARX1 I_1571 (I29591,I2859,I29455,I29423,);
nand I_1572 (I29622,I29566,I121377);
nand I_1573 (I29639,I29489,I29622);
not I_1574 (I29435,I29639);
DFFARX1 I_1575 (I121380,I2859,I29455,I29679,);
DFFARX1 I_1576 (I29679,I2859,I29455,I29444,);
nand I_1577 (I29701,I121359,I121371);
and I_1578 (I29718,I29701,I121365);
DFFARX1 I_1579 (I29718,I2859,I29455,I29744,);
DFFARX1 I_1580 (I29744,I2859,I29455,I29761,);
not I_1581 (I29447,I29761);
not I_1582 (I29783,I29744);
nand I_1583 (I29432,I29783,I29622);
nor I_1584 (I29814,I121374,I121371);
not I_1585 (I29831,I29814);
nor I_1586 (I29848,I29783,I29831);
nor I_1587 (I29865,I29489,I29848);
DFFARX1 I_1588 (I29865,I2859,I29455,I29441,);
nor I_1589 (I29896,I29549,I29831);
nor I_1590 (I29429,I29744,I29896);
nor I_1591 (I29438,I29679,I29814);
nor I_1592 (I29426,I29549,I29814);
not I_1593 (I29982,I2866);
DFFARX1 I_1594 (I127710,I2859,I29982,I30008,);
not I_1595 (I30016,I30008);
nand I_1596 (I30033,I127692,I127707);
and I_1597 (I30050,I30033,I127683);
DFFARX1 I_1598 (I30050,I2859,I29982,I30076,);
DFFARX1 I_1599 (I127686,I2859,I29982,I30093,);
and I_1600 (I30101,I30093,I127701);
nor I_1601 (I30118,I30076,I30101);
DFFARX1 I_1602 (I30118,I2859,I29982,I29950,);
nand I_1603 (I30149,I30093,I127701);
nand I_1604 (I30166,I30016,I30149);
not I_1605 (I29962,I30166);
DFFARX1 I_1606 (I127704,I2859,I29982,I30206,);
DFFARX1 I_1607 (I30206,I2859,I29982,I29971,);
nand I_1608 (I30228,I127683,I127695);
and I_1609 (I30245,I30228,I127689);
DFFARX1 I_1610 (I30245,I2859,I29982,I30271,);
DFFARX1 I_1611 (I30271,I2859,I29982,I30288,);
not I_1612 (I29974,I30288);
not I_1613 (I30310,I30271);
nand I_1614 (I29959,I30310,I30149);
nor I_1615 (I30341,I127698,I127695);
not I_1616 (I30358,I30341);
nor I_1617 (I30375,I30310,I30358);
nor I_1618 (I30392,I30016,I30375);
DFFARX1 I_1619 (I30392,I2859,I29982,I29968,);
nor I_1620 (I30423,I30076,I30358);
nor I_1621 (I29956,I30271,I30423);
nor I_1622 (I29965,I30206,I30341);
nor I_1623 (I29953,I30076,I30341);
not I_1624 (I30509,I2866);
DFFARX1 I_1625 (I314168,I2859,I30509,I30535,);
not I_1626 (I30543,I30535);
nand I_1627 (I30560,I314159,I314177);
and I_1628 (I30577,I30560,I314156);
DFFARX1 I_1629 (I30577,I2859,I30509,I30603,);
DFFARX1 I_1630 (I314159,I2859,I30509,I30620,);
and I_1631 (I30628,I30620,I314162);
nor I_1632 (I30645,I30603,I30628);
DFFARX1 I_1633 (I30645,I2859,I30509,I30477,);
nand I_1634 (I30676,I30620,I314162);
nand I_1635 (I30693,I30543,I30676);
not I_1636 (I30489,I30693);
DFFARX1 I_1637 (I314156,I2859,I30509,I30733,);
DFFARX1 I_1638 (I30733,I2859,I30509,I30498,);
nand I_1639 (I30755,I314174,I314165);
and I_1640 (I30772,I30755,I314180);
DFFARX1 I_1641 (I30772,I2859,I30509,I30798,);
DFFARX1 I_1642 (I30798,I2859,I30509,I30815,);
not I_1643 (I30501,I30815);
not I_1644 (I30837,I30798);
nand I_1645 (I30486,I30837,I30676);
nor I_1646 (I30868,I314171,I314165);
not I_1647 (I30885,I30868);
nor I_1648 (I30902,I30837,I30885);
nor I_1649 (I30919,I30543,I30902);
DFFARX1 I_1650 (I30919,I2859,I30509,I30495,);
nor I_1651 (I30950,I30603,I30885);
nor I_1652 (I30483,I30798,I30950);
nor I_1653 (I30492,I30733,I30868);
nor I_1654 (I30480,I30603,I30868);
not I_1655 (I31036,I2866);
DFFARX1 I_1656 (I468556,I2859,I31036,I31062,);
not I_1657 (I31070,I31062);
nand I_1658 (I31087,I468571,I468550);
and I_1659 (I31104,I31087,I468553);
DFFARX1 I_1660 (I31104,I2859,I31036,I31130,);
DFFARX1 I_1661 (I468574,I2859,I31036,I31147,);
and I_1662 (I31155,I31147,I468553);
nor I_1663 (I31172,I31130,I31155);
DFFARX1 I_1664 (I31172,I2859,I31036,I31004,);
nand I_1665 (I31203,I31147,I468553);
nand I_1666 (I31220,I31070,I31203);
not I_1667 (I31016,I31220);
DFFARX1 I_1668 (I468550,I2859,I31036,I31260,);
DFFARX1 I_1669 (I31260,I2859,I31036,I31025,);
nand I_1670 (I31282,I468562,I468559);
and I_1671 (I31299,I31282,I468565);
DFFARX1 I_1672 (I31299,I2859,I31036,I31325,);
DFFARX1 I_1673 (I31325,I2859,I31036,I31342,);
not I_1674 (I31028,I31342);
not I_1675 (I31364,I31325);
nand I_1676 (I31013,I31364,I31203);
nor I_1677 (I31395,I468568,I468559);
not I_1678 (I31412,I31395);
nor I_1679 (I31429,I31364,I31412);
nor I_1680 (I31446,I31070,I31429);
DFFARX1 I_1681 (I31446,I2859,I31036,I31022,);
nor I_1682 (I31477,I31130,I31412);
nor I_1683 (I31010,I31325,I31477);
nor I_1684 (I31019,I31260,I31395);
nor I_1685 (I31007,I31130,I31395);
not I_1686 (I31563,I2866);
DFFARX1 I_1687 (I192845,I2859,I31563,I31589,);
not I_1688 (I31597,I31589);
nand I_1689 (I31614,I192839,I192830);
and I_1690 (I31631,I31614,I192851);
DFFARX1 I_1691 (I31631,I2859,I31563,I31657,);
DFFARX1 I_1692 (I192833,I2859,I31563,I31674,);
and I_1693 (I31682,I31674,I192827);
nor I_1694 (I31699,I31657,I31682);
DFFARX1 I_1695 (I31699,I2859,I31563,I31531,);
nand I_1696 (I31730,I31674,I192827);
nand I_1697 (I31747,I31597,I31730);
not I_1698 (I31543,I31747);
DFFARX1 I_1699 (I192827,I2859,I31563,I31787,);
DFFARX1 I_1700 (I31787,I2859,I31563,I31552,);
nand I_1701 (I31809,I192854,I192836);
and I_1702 (I31826,I31809,I192842);
DFFARX1 I_1703 (I31826,I2859,I31563,I31852,);
DFFARX1 I_1704 (I31852,I2859,I31563,I31869,);
not I_1705 (I31555,I31869);
not I_1706 (I31891,I31852);
nand I_1707 (I31540,I31891,I31730);
nor I_1708 (I31922,I192848,I192836);
not I_1709 (I31939,I31922);
nor I_1710 (I31956,I31891,I31939);
nor I_1711 (I31973,I31597,I31956);
DFFARX1 I_1712 (I31973,I2859,I31563,I31549,);
nor I_1713 (I32004,I31657,I31939);
nor I_1714 (I31537,I31852,I32004);
nor I_1715 (I31546,I31787,I31922);
nor I_1716 (I31534,I31657,I31922);
not I_1717 (I32090,I2866);
DFFARX1 I_1718 (I78650,I2859,I32090,I32116,);
not I_1719 (I32124,I32116);
nand I_1720 (I32141,I78644,I78638);
and I_1721 (I32158,I32141,I78659);
DFFARX1 I_1722 (I32158,I2859,I32090,I32184,);
DFFARX1 I_1723 (I78656,I2859,I32090,I32201,);
and I_1724 (I32209,I32201,I78653);
nor I_1725 (I32226,I32184,I32209);
DFFARX1 I_1726 (I32226,I2859,I32090,I32058,);
nand I_1727 (I32257,I32201,I78653);
nand I_1728 (I32274,I32124,I32257);
not I_1729 (I32070,I32274);
DFFARX1 I_1730 (I78638,I2859,I32090,I32314,);
DFFARX1 I_1731 (I32314,I2859,I32090,I32079,);
nand I_1732 (I32336,I78641,I78641);
and I_1733 (I32353,I32336,I78662);
DFFARX1 I_1734 (I32353,I2859,I32090,I32379,);
DFFARX1 I_1735 (I32379,I2859,I32090,I32396,);
not I_1736 (I32082,I32396);
not I_1737 (I32418,I32379);
nand I_1738 (I32067,I32418,I32257);
nor I_1739 (I32449,I78647,I78641);
not I_1740 (I32466,I32449);
nor I_1741 (I32483,I32418,I32466);
nor I_1742 (I32500,I32124,I32483);
DFFARX1 I_1743 (I32500,I2859,I32090,I32076,);
nor I_1744 (I32531,I32184,I32466);
nor I_1745 (I32064,I32379,I32531);
nor I_1746 (I32073,I32314,I32449);
nor I_1747 (I32061,I32184,I32449);
not I_1748 (I32617,I2866);
DFFARX1 I_1749 (I335296,I2859,I32617,I32643,);
not I_1750 (I32651,I32643);
nand I_1751 (I32668,I335293,I335308);
and I_1752 (I32685,I32668,I335290);
DFFARX1 I_1753 (I32685,I2859,I32617,I32711,);
DFFARX1 I_1754 (I335287,I2859,I32617,I32728,);
and I_1755 (I32736,I32728,I335287);
nor I_1756 (I32753,I32711,I32736);
DFFARX1 I_1757 (I32753,I2859,I32617,I32585,);
nand I_1758 (I32784,I32728,I335287);
nand I_1759 (I32801,I32651,I32784);
not I_1760 (I32597,I32801);
DFFARX1 I_1761 (I335290,I2859,I32617,I32841,);
DFFARX1 I_1762 (I32841,I2859,I32617,I32606,);
nand I_1763 (I32863,I335302,I335293);
and I_1764 (I32880,I32863,I335305);
DFFARX1 I_1765 (I32880,I2859,I32617,I32906,);
DFFARX1 I_1766 (I32906,I2859,I32617,I32923,);
not I_1767 (I32609,I32923);
not I_1768 (I32945,I32906);
nand I_1769 (I32594,I32945,I32784);
nor I_1770 (I32976,I335299,I335293);
not I_1771 (I32993,I32976);
nor I_1772 (I33010,I32945,I32993);
nor I_1773 (I33027,I32651,I33010);
DFFARX1 I_1774 (I33027,I2859,I32617,I32603,);
nor I_1775 (I33058,I32711,I32993);
nor I_1776 (I32591,I32906,I33058);
nor I_1777 (I32600,I32841,I32976);
nor I_1778 (I32588,I32711,I32976);
not I_1779 (I33144,I2866);
DFFARX1 I_1780 (I281800,I2859,I33144,I33170,);
not I_1781 (I33178,I33170);
nand I_1782 (I33195,I281791,I281809);
and I_1783 (I33212,I33195,I281788);
DFFARX1 I_1784 (I33212,I2859,I33144,I33238,);
DFFARX1 I_1785 (I281791,I2859,I33144,I33255,);
and I_1786 (I33263,I33255,I281794);
nor I_1787 (I33280,I33238,I33263);
DFFARX1 I_1788 (I33280,I2859,I33144,I33112,);
nand I_1789 (I33311,I33255,I281794);
nand I_1790 (I33328,I33178,I33311);
not I_1791 (I33124,I33328);
DFFARX1 I_1792 (I281788,I2859,I33144,I33368,);
DFFARX1 I_1793 (I33368,I2859,I33144,I33133,);
nand I_1794 (I33390,I281806,I281797);
and I_1795 (I33407,I33390,I281812);
DFFARX1 I_1796 (I33407,I2859,I33144,I33433,);
DFFARX1 I_1797 (I33433,I2859,I33144,I33450,);
not I_1798 (I33136,I33450);
not I_1799 (I33472,I33433);
nand I_1800 (I33121,I33472,I33311);
nor I_1801 (I33503,I281803,I281797);
not I_1802 (I33520,I33503);
nor I_1803 (I33537,I33472,I33520);
nor I_1804 (I33554,I33178,I33537);
DFFARX1 I_1805 (I33554,I2859,I33144,I33130,);
nor I_1806 (I33585,I33238,I33520);
nor I_1807 (I33118,I33433,I33585);
nor I_1808 (I33127,I33368,I33503);
nor I_1809 (I33115,I33238,I33503);
not I_1810 (I33671,I2866);
DFFARX1 I_1811 (I100070,I2859,I33671,I33697,);
not I_1812 (I33705,I33697);
nand I_1813 (I33722,I100064,I100058);
and I_1814 (I33739,I33722,I100079);
DFFARX1 I_1815 (I33739,I2859,I33671,I33765,);
DFFARX1 I_1816 (I100076,I2859,I33671,I33782,);
and I_1817 (I33790,I33782,I100073);
nor I_1818 (I33807,I33765,I33790);
DFFARX1 I_1819 (I33807,I2859,I33671,I33639,);
nand I_1820 (I33838,I33782,I100073);
nand I_1821 (I33855,I33705,I33838);
not I_1822 (I33651,I33855);
DFFARX1 I_1823 (I100058,I2859,I33671,I33895,);
DFFARX1 I_1824 (I33895,I2859,I33671,I33660,);
nand I_1825 (I33917,I100061,I100061);
and I_1826 (I33934,I33917,I100082);
DFFARX1 I_1827 (I33934,I2859,I33671,I33960,);
DFFARX1 I_1828 (I33960,I2859,I33671,I33977,);
not I_1829 (I33663,I33977);
not I_1830 (I33999,I33960);
nand I_1831 (I33648,I33999,I33838);
nor I_1832 (I34030,I100067,I100061);
not I_1833 (I34047,I34030);
nor I_1834 (I34064,I33999,I34047);
nor I_1835 (I34081,I33705,I34064);
DFFARX1 I_1836 (I34081,I2859,I33671,I33657,);
nor I_1837 (I34112,I33765,I34047);
nor I_1838 (I33645,I33960,I34112);
nor I_1839 (I33654,I33895,I34030);
nor I_1840 (I33642,I33765,I34030);
not I_1841 (I34198,I2866);
DFFARX1 I_1842 (I469134,I2859,I34198,I34224,);
not I_1843 (I34232,I34224);
nand I_1844 (I34249,I469149,I469128);
and I_1845 (I34266,I34249,I469131);
DFFARX1 I_1846 (I34266,I2859,I34198,I34292,);
DFFARX1 I_1847 (I469152,I2859,I34198,I34309,);
and I_1848 (I34317,I34309,I469131);
nor I_1849 (I34334,I34292,I34317);
DFFARX1 I_1850 (I34334,I2859,I34198,I34166,);
nand I_1851 (I34365,I34309,I469131);
nand I_1852 (I34382,I34232,I34365);
not I_1853 (I34178,I34382);
DFFARX1 I_1854 (I469128,I2859,I34198,I34422,);
DFFARX1 I_1855 (I34422,I2859,I34198,I34187,);
nand I_1856 (I34444,I469140,I469137);
and I_1857 (I34461,I34444,I469143);
DFFARX1 I_1858 (I34461,I2859,I34198,I34487,);
DFFARX1 I_1859 (I34487,I2859,I34198,I34504,);
not I_1860 (I34190,I34504);
not I_1861 (I34526,I34487);
nand I_1862 (I34175,I34526,I34365);
nor I_1863 (I34557,I469146,I469137);
not I_1864 (I34574,I34557);
nor I_1865 (I34591,I34526,I34574);
nor I_1866 (I34608,I34232,I34591);
DFFARX1 I_1867 (I34608,I2859,I34198,I34184,);
nor I_1868 (I34639,I34292,I34574);
nor I_1869 (I34172,I34487,I34639);
nor I_1870 (I34181,I34422,I34557);
nor I_1871 (I34169,I34292,I34557);
not I_1872 (I34725,I2866);
DFFARX1 I_1873 (I402242,I2859,I34725,I34751,);
not I_1874 (I34759,I34751);
nand I_1875 (I34776,I402260,I402254);
and I_1876 (I34793,I34776,I402233);
DFFARX1 I_1877 (I34793,I2859,I34725,I34819,);
DFFARX1 I_1878 (I402251,I2859,I34725,I34836,);
and I_1879 (I34844,I34836,I402236);
nor I_1880 (I34861,I34819,I34844);
DFFARX1 I_1881 (I34861,I2859,I34725,I34693,);
nand I_1882 (I34892,I34836,I402236);
nand I_1883 (I34909,I34759,I34892);
not I_1884 (I34705,I34909);
DFFARX1 I_1885 (I402248,I2859,I34725,I34949,);
DFFARX1 I_1886 (I34949,I2859,I34725,I34714,);
nand I_1887 (I34971,I402257,I402245);
and I_1888 (I34988,I34971,I402239);
DFFARX1 I_1889 (I34988,I2859,I34725,I35014,);
DFFARX1 I_1890 (I35014,I2859,I34725,I35031,);
not I_1891 (I34717,I35031);
not I_1892 (I35053,I35014);
nand I_1893 (I34702,I35053,I34892);
nor I_1894 (I35084,I402233,I402245);
not I_1895 (I35101,I35084);
nor I_1896 (I35118,I35053,I35101);
nor I_1897 (I35135,I34759,I35118);
DFFARX1 I_1898 (I35135,I2859,I34725,I34711,);
nor I_1899 (I35166,I34819,I35101);
nor I_1900 (I34699,I35014,I35166);
nor I_1901 (I34708,I34949,I35084);
nor I_1902 (I34696,I34819,I35084);
not I_1903 (I35252,I2866);
DFFARX1 I_1904 (I213706,I2859,I35252,I35278,);
not I_1905 (I35286,I35278);
nand I_1906 (I35303,I213727,I213721);
and I_1907 (I35320,I35303,I213703);
DFFARX1 I_1908 (I35320,I2859,I35252,I35346,);
DFFARX1 I_1909 (I213706,I2859,I35252,I35363,);
and I_1910 (I35371,I35363,I213715);
nor I_1911 (I35388,I35346,I35371);
DFFARX1 I_1912 (I35388,I2859,I35252,I35220,);
nand I_1913 (I35419,I35363,I213715);
nand I_1914 (I35436,I35286,I35419);
not I_1915 (I35232,I35436);
DFFARX1 I_1916 (I213712,I2859,I35252,I35476,);
DFFARX1 I_1917 (I35476,I2859,I35252,I35241,);
nand I_1918 (I35498,I213718,I213709);
and I_1919 (I35515,I35498,I213703);
DFFARX1 I_1920 (I35515,I2859,I35252,I35541,);
DFFARX1 I_1921 (I35541,I2859,I35252,I35558,);
not I_1922 (I35244,I35558);
not I_1923 (I35580,I35541);
nand I_1924 (I35229,I35580,I35419);
nor I_1925 (I35611,I213724,I213709);
not I_1926 (I35628,I35611);
nor I_1927 (I35645,I35580,I35628);
nor I_1928 (I35662,I35286,I35645);
DFFARX1 I_1929 (I35662,I2859,I35252,I35238,);
nor I_1930 (I35693,I35346,I35628);
nor I_1931 (I35226,I35541,I35693);
nor I_1932 (I35235,I35476,I35611);
nor I_1933 (I35223,I35346,I35611);
not I_1934 (I35779,I2866);
DFFARX1 I_1935 (I503168,I2859,I35779,I35805,);
not I_1936 (I35813,I35805);
nand I_1937 (I35830,I503162,I503183);
and I_1938 (I35847,I35830,I503174);
DFFARX1 I_1939 (I35847,I2859,I35779,I35873,);
DFFARX1 I_1940 (I503165,I2859,I35779,I35890,);
and I_1941 (I35898,I35890,I503177);
nor I_1942 (I35915,I35873,I35898);
DFFARX1 I_1943 (I35915,I2859,I35779,I35747,);
nand I_1944 (I35946,I35890,I503177);
nand I_1945 (I35963,I35813,I35946);
not I_1946 (I35759,I35963);
DFFARX1 I_1947 (I503165,I2859,I35779,I36003,);
DFFARX1 I_1948 (I36003,I2859,I35779,I35768,);
nand I_1949 (I36025,I503186,I503171);
and I_1950 (I36042,I36025,I503162);
DFFARX1 I_1951 (I36042,I2859,I35779,I36068,);
DFFARX1 I_1952 (I36068,I2859,I35779,I36085,);
not I_1953 (I35771,I36085);
not I_1954 (I36107,I36068);
nand I_1955 (I35756,I36107,I35946);
nor I_1956 (I36138,I503180,I503171);
not I_1957 (I36155,I36138);
nor I_1958 (I36172,I36107,I36155);
nor I_1959 (I36189,I35813,I36172);
DFFARX1 I_1960 (I36189,I2859,I35779,I35765,);
nor I_1961 (I36220,I35873,I36155);
nor I_1962 (I35753,I36068,I36220);
nor I_1963 (I35762,I36003,I36138);
nor I_1964 (I35750,I35873,I36138);
not I_1965 (I36306,I2866);
DFFARX1 I_1966 (I367443,I2859,I36306,I36332,);
not I_1967 (I36340,I36332);
nand I_1968 (I36357,I367440,I367455);
and I_1969 (I36374,I36357,I367437);
DFFARX1 I_1970 (I36374,I2859,I36306,I36400,);
DFFARX1 I_1971 (I367434,I2859,I36306,I36417,);
and I_1972 (I36425,I36417,I367434);
nor I_1973 (I36442,I36400,I36425);
DFFARX1 I_1974 (I36442,I2859,I36306,I36274,);
nand I_1975 (I36473,I36417,I367434);
nand I_1976 (I36490,I36340,I36473);
not I_1977 (I36286,I36490);
DFFARX1 I_1978 (I367437,I2859,I36306,I36530,);
DFFARX1 I_1979 (I36530,I2859,I36306,I36295,);
nand I_1980 (I36552,I367449,I367440);
and I_1981 (I36569,I36552,I367452);
DFFARX1 I_1982 (I36569,I2859,I36306,I36595,);
DFFARX1 I_1983 (I36595,I2859,I36306,I36612,);
not I_1984 (I36298,I36612);
not I_1985 (I36634,I36595);
nand I_1986 (I36283,I36634,I36473);
nor I_1987 (I36665,I367446,I367440);
not I_1988 (I36682,I36665);
nor I_1989 (I36699,I36634,I36682);
nor I_1990 (I36716,I36340,I36699);
DFFARX1 I_1991 (I36716,I2859,I36306,I36292,);
nor I_1992 (I36747,I36400,I36682);
nor I_1993 (I36280,I36595,I36747);
nor I_1994 (I36289,I36530,I36665);
nor I_1995 (I36277,I36400,I36665);
not I_1996 (I36833,I2866);
DFFARX1 I_1997 (I340566,I2859,I36833,I36859,);
not I_1998 (I36867,I36859);
nand I_1999 (I36884,I340563,I340578);
and I_2000 (I36901,I36884,I340560);
DFFARX1 I_2001 (I36901,I2859,I36833,I36927,);
DFFARX1 I_2002 (I340557,I2859,I36833,I36944,);
and I_2003 (I36952,I36944,I340557);
nor I_2004 (I36969,I36927,I36952);
DFFARX1 I_2005 (I36969,I2859,I36833,I36801,);
nand I_2006 (I37000,I36944,I340557);
nand I_2007 (I37017,I36867,I37000);
not I_2008 (I36813,I37017);
DFFARX1 I_2009 (I340560,I2859,I36833,I37057,);
DFFARX1 I_2010 (I37057,I2859,I36833,I36822,);
nand I_2011 (I37079,I340572,I340563);
and I_2012 (I37096,I37079,I340575);
DFFARX1 I_2013 (I37096,I2859,I36833,I37122,);
DFFARX1 I_2014 (I37122,I2859,I36833,I37139,);
not I_2015 (I36825,I37139);
not I_2016 (I37161,I37122);
nand I_2017 (I36810,I37161,I37000);
nor I_2018 (I37192,I340569,I340563);
not I_2019 (I37209,I37192);
nor I_2020 (I37226,I37161,I37209);
nor I_2021 (I37243,I36867,I37226);
DFFARX1 I_2022 (I37243,I2859,I36833,I36819,);
nor I_2023 (I37274,I36927,I37209);
nor I_2024 (I36807,I37122,I37274);
nor I_2025 (I36816,I37057,I37192);
nor I_2026 (I36804,I36927,I37192);
not I_2027 (I37360,I2866);
DFFARX1 I_2028 (I418392,I2859,I37360,I37386,);
not I_2029 (I37394,I37386);
nand I_2030 (I37411,I418410,I418404);
and I_2031 (I37428,I37411,I418383);
DFFARX1 I_2032 (I37428,I2859,I37360,I37454,);
DFFARX1 I_2033 (I418401,I2859,I37360,I37471,);
and I_2034 (I37479,I37471,I418386);
nor I_2035 (I37496,I37454,I37479);
DFFARX1 I_2036 (I37496,I2859,I37360,I37328,);
nand I_2037 (I37527,I37471,I418386);
nand I_2038 (I37544,I37394,I37527);
not I_2039 (I37340,I37544);
DFFARX1 I_2040 (I418398,I2859,I37360,I37584,);
DFFARX1 I_2041 (I37584,I2859,I37360,I37349,);
nand I_2042 (I37606,I418407,I418395);
and I_2043 (I37623,I37606,I418389);
DFFARX1 I_2044 (I37623,I2859,I37360,I37649,);
DFFARX1 I_2045 (I37649,I2859,I37360,I37666,);
not I_2046 (I37352,I37666);
not I_2047 (I37688,I37649);
nand I_2048 (I37337,I37688,I37527);
nor I_2049 (I37719,I418383,I418395);
not I_2050 (I37736,I37719);
nor I_2051 (I37753,I37688,I37736);
nor I_2052 (I37770,I37394,I37753);
DFFARX1 I_2053 (I37770,I2859,I37360,I37346,);
nor I_2054 (I37801,I37454,I37736);
nor I_2055 (I37334,I37649,I37801);
nor I_2056 (I37343,I37584,I37719);
nor I_2057 (I37331,I37454,I37719);
not I_2058 (I37887,I2866);
DFFARX1 I_2059 (I243649,I2859,I37887,I37913,);
not I_2060 (I37921,I37913);
nand I_2061 (I37938,I243661,I243646);
and I_2062 (I37955,I37938,I243640);
DFFARX1 I_2063 (I37955,I2859,I37887,I37981,);
DFFARX1 I_2064 (I243655,I2859,I37887,I37998,);
and I_2065 (I38006,I37998,I243643);
nor I_2066 (I38023,I37981,I38006);
DFFARX1 I_2067 (I38023,I2859,I37887,I37855,);
nand I_2068 (I38054,I37998,I243643);
nand I_2069 (I38071,I37921,I38054);
not I_2070 (I37867,I38071);
DFFARX1 I_2071 (I243652,I2859,I37887,I38111,);
DFFARX1 I_2072 (I38111,I2859,I37887,I37876,);
nand I_2073 (I38133,I243658,I243664);
and I_2074 (I38150,I38133,I243640);
DFFARX1 I_2075 (I38150,I2859,I37887,I38176,);
DFFARX1 I_2076 (I38176,I2859,I37887,I38193,);
not I_2077 (I37879,I38193);
not I_2078 (I38215,I38176);
nand I_2079 (I37864,I38215,I38054);
nor I_2080 (I38246,I243643,I243664);
not I_2081 (I38263,I38246);
nor I_2082 (I38280,I38215,I38263);
nor I_2083 (I38297,I37921,I38280);
DFFARX1 I_2084 (I38297,I2859,I37887,I37873,);
nor I_2085 (I38328,I37981,I38263);
nor I_2086 (I37861,I38176,I38328);
nor I_2087 (I37870,I38111,I38246);
nor I_2088 (I37858,I37981,I38246);
not I_2089 (I38414,I2866);
DFFARX1 I_2090 (I439347,I2859,I38414,I38440,);
not I_2091 (I38448,I38440);
nand I_2092 (I38465,I439344,I439350);
and I_2093 (I38482,I38465,I439347);
DFFARX1 I_2094 (I38482,I2859,I38414,I38508,);
DFFARX1 I_2095 (I439350,I2859,I38414,I38525,);
and I_2096 (I38533,I38525,I439344);
nor I_2097 (I38550,I38508,I38533);
DFFARX1 I_2098 (I38550,I2859,I38414,I38382,);
nand I_2099 (I38581,I38525,I439344);
nand I_2100 (I38598,I38448,I38581);
not I_2101 (I38394,I38598);
DFFARX1 I_2102 (I439353,I2859,I38414,I38638,);
DFFARX1 I_2103 (I38638,I2859,I38414,I38403,);
nand I_2104 (I38660,I439356,I439365);
and I_2105 (I38677,I38660,I439359);
DFFARX1 I_2106 (I38677,I2859,I38414,I38703,);
DFFARX1 I_2107 (I38703,I2859,I38414,I38720,);
not I_2108 (I38406,I38720);
not I_2109 (I38742,I38703);
nand I_2110 (I38391,I38742,I38581);
nor I_2111 (I38773,I439362,I439365);
not I_2112 (I38790,I38773);
nor I_2113 (I38807,I38742,I38790);
nor I_2114 (I38824,I38448,I38807);
DFFARX1 I_2115 (I38824,I2859,I38414,I38400,);
nor I_2116 (I38855,I38508,I38790);
nor I_2117 (I38388,I38703,I38855);
nor I_2118 (I38397,I38638,I38773);
nor I_2119 (I38385,I38508,I38773);
not I_2120 (I38941,I2866);
DFFARX1 I_2121 (I557982,I2859,I38941,I38967,);
not I_2122 (I38975,I38967);
nand I_2123 (I38992,I557976,I557997);
and I_2124 (I39009,I38992,I557973);
DFFARX1 I_2125 (I39009,I2859,I38941,I39035,);
DFFARX1 I_2126 (I557994,I2859,I38941,I39052,);
and I_2127 (I39060,I39052,I557991);
nor I_2128 (I39077,I39035,I39060);
DFFARX1 I_2129 (I39077,I2859,I38941,I38909,);
nand I_2130 (I39108,I39052,I557991);
nand I_2131 (I39125,I38975,I39108);
not I_2132 (I38921,I39125);
DFFARX1 I_2133 (I557979,I2859,I38941,I39165,);
DFFARX1 I_2134 (I39165,I2859,I38941,I38930,);
nand I_2135 (I39187,I557988,I557985);
and I_2136 (I39204,I39187,I557970);
DFFARX1 I_2137 (I39204,I2859,I38941,I39230,);
DFFARX1 I_2138 (I39230,I2859,I38941,I39247,);
not I_2139 (I38933,I39247);
not I_2140 (I39269,I39230);
nand I_2141 (I38918,I39269,I39108);
nor I_2142 (I39300,I557970,I557985);
not I_2143 (I39317,I39300);
nor I_2144 (I39334,I39269,I39317);
nor I_2145 (I39351,I38975,I39334);
DFFARX1 I_2146 (I39351,I2859,I38941,I38927,);
nor I_2147 (I39382,I39035,I39317);
nor I_2148 (I38915,I39230,I39382);
nor I_2149 (I38924,I39165,I39300);
nor I_2150 (I38912,I39035,I39300);
not I_2151 (I39468,I2866);
DFFARX1 I_2152 (I403534,I2859,I39468,I39494,);
not I_2153 (I39502,I39494);
nand I_2154 (I39519,I403552,I403546);
and I_2155 (I39536,I39519,I403525);
DFFARX1 I_2156 (I39536,I2859,I39468,I39562,);
DFFARX1 I_2157 (I403543,I2859,I39468,I39579,);
and I_2158 (I39587,I39579,I403528);
nor I_2159 (I39604,I39562,I39587);
DFFARX1 I_2160 (I39604,I2859,I39468,I39436,);
nand I_2161 (I39635,I39579,I403528);
nand I_2162 (I39652,I39502,I39635);
not I_2163 (I39448,I39652);
DFFARX1 I_2164 (I403540,I2859,I39468,I39692,);
DFFARX1 I_2165 (I39692,I2859,I39468,I39457,);
nand I_2166 (I39714,I403549,I403537);
and I_2167 (I39731,I39714,I403531);
DFFARX1 I_2168 (I39731,I2859,I39468,I39757,);
DFFARX1 I_2169 (I39757,I2859,I39468,I39774,);
not I_2170 (I39460,I39774);
not I_2171 (I39796,I39757);
nand I_2172 (I39445,I39796,I39635);
nor I_2173 (I39827,I403525,I403537);
not I_2174 (I39844,I39827);
nor I_2175 (I39861,I39796,I39844);
nor I_2176 (I39878,I39502,I39861);
DFFARX1 I_2177 (I39878,I2859,I39468,I39454,);
nor I_2178 (I39909,I39562,I39844);
nor I_2179 (I39442,I39757,I39909);
nor I_2180 (I39451,I39692,I39827);
nor I_2181 (I39439,I39562,I39827);
not I_2182 (I39995,I2866);
DFFARX1 I_2183 (I16272,I2859,I39995,I40021,);
not I_2184 (I40029,I40021);
nand I_2185 (I40046,I16260,I16266);
and I_2186 (I40063,I40046,I16269);
DFFARX1 I_2187 (I40063,I2859,I39995,I40089,);
DFFARX1 I_2188 (I16251,I2859,I39995,I40106,);
and I_2189 (I40114,I40106,I16257);
nor I_2190 (I40131,I40089,I40114);
DFFARX1 I_2191 (I40131,I2859,I39995,I39963,);
nand I_2192 (I40162,I40106,I16257);
nand I_2193 (I40179,I40029,I40162);
not I_2194 (I39975,I40179);
DFFARX1 I_2195 (I16251,I2859,I39995,I40219,);
DFFARX1 I_2196 (I40219,I2859,I39995,I39984,);
nand I_2197 (I40241,I16254,I16248);
and I_2198 (I40258,I40241,I16263);
DFFARX1 I_2199 (I40258,I2859,I39995,I40284,);
DFFARX1 I_2200 (I40284,I2859,I39995,I40301,);
not I_2201 (I39987,I40301);
not I_2202 (I40323,I40284);
nand I_2203 (I39972,I40323,I40162);
nor I_2204 (I40354,I16248,I16248);
not I_2205 (I40371,I40354);
nor I_2206 (I40388,I40323,I40371);
nor I_2207 (I40405,I40029,I40388);
DFFARX1 I_2208 (I40405,I2859,I39995,I39981,);
nor I_2209 (I40436,I40089,I40371);
nor I_2210 (I39969,I40284,I40436);
nor I_2211 (I39978,I40219,I40354);
nor I_2212 (I39966,I40089,I40354);
not I_2213 (I40522,I2866);
DFFARX1 I_2214 (I271974,I2859,I40522,I40548,);
not I_2215 (I40556,I40548);
nand I_2216 (I40573,I271965,I271983);
and I_2217 (I40590,I40573,I271962);
DFFARX1 I_2218 (I40590,I2859,I40522,I40616,);
DFFARX1 I_2219 (I271965,I2859,I40522,I40633,);
and I_2220 (I40641,I40633,I271968);
nor I_2221 (I40658,I40616,I40641);
DFFARX1 I_2222 (I40658,I2859,I40522,I40490,);
nand I_2223 (I40689,I40633,I271968);
nand I_2224 (I40706,I40556,I40689);
not I_2225 (I40502,I40706);
DFFARX1 I_2226 (I271962,I2859,I40522,I40746,);
DFFARX1 I_2227 (I40746,I2859,I40522,I40511,);
nand I_2228 (I40768,I271980,I271971);
and I_2229 (I40785,I40768,I271986);
DFFARX1 I_2230 (I40785,I2859,I40522,I40811,);
DFFARX1 I_2231 (I40811,I2859,I40522,I40828,);
not I_2232 (I40514,I40828);
not I_2233 (I40850,I40811);
nand I_2234 (I40499,I40850,I40689);
nor I_2235 (I40881,I271977,I271971);
not I_2236 (I40898,I40881);
nor I_2237 (I40915,I40850,I40898);
nor I_2238 (I40932,I40556,I40915);
DFFARX1 I_2239 (I40932,I2859,I40522,I40508,);
nor I_2240 (I40963,I40616,I40898);
nor I_2241 (I40496,I40811,I40963);
nor I_2242 (I40505,I40746,I40881);
nor I_2243 (I40493,I40616,I40881);
not I_2244 (I41049,I2866);
DFFARX1 I_2245 (I497456,I2859,I41049,I41075,);
not I_2246 (I41083,I41075);
nand I_2247 (I41100,I497471,I497450);
and I_2248 (I41117,I41100,I497453);
DFFARX1 I_2249 (I41117,I2859,I41049,I41143,);
DFFARX1 I_2250 (I497474,I2859,I41049,I41160,);
and I_2251 (I41168,I41160,I497453);
nor I_2252 (I41185,I41143,I41168);
DFFARX1 I_2253 (I41185,I2859,I41049,I41017,);
nand I_2254 (I41216,I41160,I497453);
nand I_2255 (I41233,I41083,I41216);
not I_2256 (I41029,I41233);
DFFARX1 I_2257 (I497450,I2859,I41049,I41273,);
DFFARX1 I_2258 (I41273,I2859,I41049,I41038,);
nand I_2259 (I41295,I497462,I497459);
and I_2260 (I41312,I41295,I497465);
DFFARX1 I_2261 (I41312,I2859,I41049,I41338,);
DFFARX1 I_2262 (I41338,I2859,I41049,I41355,);
not I_2263 (I41041,I41355);
not I_2264 (I41377,I41338);
nand I_2265 (I41026,I41377,I41216);
nor I_2266 (I41408,I497468,I497459);
not I_2267 (I41425,I41408);
nor I_2268 (I41442,I41377,I41425);
nor I_2269 (I41459,I41083,I41442);
DFFARX1 I_2270 (I41459,I2859,I41049,I41035,);
nor I_2271 (I41490,I41143,I41425);
nor I_2272 (I41023,I41338,I41490);
nor I_2273 (I41032,I41273,I41408);
nor I_2274 (I41020,I41143,I41408);
not I_2275 (I41576,I2866);
DFFARX1 I_2276 (I557387,I2859,I41576,I41602,);
not I_2277 (I41610,I41602);
nand I_2278 (I41627,I557381,I557402);
and I_2279 (I41644,I41627,I557378);
DFFARX1 I_2280 (I41644,I2859,I41576,I41670,);
DFFARX1 I_2281 (I557399,I2859,I41576,I41687,);
and I_2282 (I41695,I41687,I557396);
nor I_2283 (I41712,I41670,I41695);
DFFARX1 I_2284 (I41712,I2859,I41576,I41544,);
nand I_2285 (I41743,I41687,I557396);
nand I_2286 (I41760,I41610,I41743);
not I_2287 (I41556,I41760);
DFFARX1 I_2288 (I557384,I2859,I41576,I41800,);
DFFARX1 I_2289 (I41800,I2859,I41576,I41565,);
nand I_2290 (I41822,I557393,I557390);
and I_2291 (I41839,I41822,I557375);
DFFARX1 I_2292 (I41839,I2859,I41576,I41865,);
DFFARX1 I_2293 (I41865,I2859,I41576,I41882,);
not I_2294 (I41568,I41882);
not I_2295 (I41904,I41865);
nand I_2296 (I41553,I41904,I41743);
nor I_2297 (I41935,I557375,I557390);
not I_2298 (I41952,I41935);
nor I_2299 (I41969,I41904,I41952);
nor I_2300 (I41986,I41610,I41969);
DFFARX1 I_2301 (I41986,I2859,I41576,I41562,);
nor I_2302 (I42017,I41670,I41952);
nor I_2303 (I41550,I41865,I42017);
nor I_2304 (I41559,I41800,I41935);
nor I_2305 (I41547,I41670,I41935);
not I_2306 (I42103,I2866);
DFFARX1 I_2307 (I261567,I2859,I42103,I42129,);
not I_2308 (I42137,I42129);
nand I_2309 (I42154,I261579,I261564);
and I_2310 (I42171,I42154,I261558);
DFFARX1 I_2311 (I42171,I2859,I42103,I42197,);
DFFARX1 I_2312 (I261573,I2859,I42103,I42214,);
and I_2313 (I42222,I42214,I261561);
nor I_2314 (I42239,I42197,I42222);
DFFARX1 I_2315 (I42239,I2859,I42103,I42071,);
nand I_2316 (I42270,I42214,I261561);
nand I_2317 (I42287,I42137,I42270);
not I_2318 (I42083,I42287);
DFFARX1 I_2319 (I261570,I2859,I42103,I42327,);
DFFARX1 I_2320 (I42327,I2859,I42103,I42092,);
nand I_2321 (I42349,I261576,I261582);
and I_2322 (I42366,I42349,I261558);
DFFARX1 I_2323 (I42366,I2859,I42103,I42392,);
DFFARX1 I_2324 (I42392,I2859,I42103,I42409,);
not I_2325 (I42095,I42409);
not I_2326 (I42431,I42392);
nand I_2327 (I42080,I42431,I42270);
nor I_2328 (I42462,I261561,I261582);
not I_2329 (I42479,I42462);
nor I_2330 (I42496,I42431,I42479);
nor I_2331 (I42513,I42137,I42496);
DFFARX1 I_2332 (I42513,I2859,I42103,I42089,);
nor I_2333 (I42544,I42197,I42479);
nor I_2334 (I42077,I42392,I42544);
nor I_2335 (I42086,I42327,I42462);
nor I_2336 (I42074,I42197,I42462);
not I_2337 (I42630,I2866);
DFFARX1 I_2338 (I369551,I2859,I42630,I42656,);
not I_2339 (I42664,I42656);
nand I_2340 (I42681,I369548,I369563);
and I_2341 (I42698,I42681,I369545);
DFFARX1 I_2342 (I42698,I2859,I42630,I42724,);
DFFARX1 I_2343 (I369542,I2859,I42630,I42741,);
and I_2344 (I42749,I42741,I369542);
nor I_2345 (I42766,I42724,I42749);
DFFARX1 I_2346 (I42766,I2859,I42630,I42598,);
nand I_2347 (I42797,I42741,I369542);
nand I_2348 (I42814,I42664,I42797);
not I_2349 (I42610,I42814);
DFFARX1 I_2350 (I369545,I2859,I42630,I42854,);
DFFARX1 I_2351 (I42854,I2859,I42630,I42619,);
nand I_2352 (I42876,I369557,I369548);
and I_2353 (I42893,I42876,I369560);
DFFARX1 I_2354 (I42893,I2859,I42630,I42919,);
DFFARX1 I_2355 (I42919,I2859,I42630,I42936,);
not I_2356 (I42622,I42936);
not I_2357 (I42958,I42919);
nand I_2358 (I42607,I42958,I42797);
nor I_2359 (I42989,I369554,I369548);
not I_2360 (I43006,I42989);
nor I_2361 (I43023,I42958,I43006);
nor I_2362 (I43040,I42664,I43023);
DFFARX1 I_2363 (I43040,I2859,I42630,I42616,);
nor I_2364 (I43071,I42724,I43006);
nor I_2365 (I42604,I42919,I43071);
nor I_2366 (I42613,I42854,I42989);
nor I_2367 (I42601,I42724,I42989);
not I_2368 (I43157,I2866);
DFFARX1 I_2369 (I2116,I2859,I43157,I43183,);
not I_2370 (I43191,I43183);
nand I_2371 (I43208,I2036,I1788);
and I_2372 (I43225,I43208,I2292);
DFFARX1 I_2373 (I43225,I2859,I43157,I43251,);
DFFARX1 I_2374 (I2132,I2859,I43157,I43268,);
and I_2375 (I43276,I43268,I1468);
nor I_2376 (I43293,I43251,I43276);
DFFARX1 I_2377 (I43293,I2859,I43157,I43125,);
nand I_2378 (I43324,I43268,I1468);
nand I_2379 (I43341,I43191,I43324);
not I_2380 (I43137,I43341);
DFFARX1 I_2381 (I1476,I2859,I43157,I43381,);
DFFARX1 I_2382 (I43381,I2859,I43157,I43146,);
nand I_2383 (I43403,I2020,I2636);
and I_2384 (I43420,I43403,I1540);
DFFARX1 I_2385 (I43420,I2859,I43157,I43446,);
DFFARX1 I_2386 (I43446,I2859,I43157,I43463,);
not I_2387 (I43149,I43463);
not I_2388 (I43485,I43446);
nand I_2389 (I43134,I43485,I43324);
nor I_2390 (I43516,I2348,I2636);
not I_2391 (I43533,I43516);
nor I_2392 (I43550,I43485,I43533);
nor I_2393 (I43567,I43191,I43550);
DFFARX1 I_2394 (I43567,I2859,I43157,I43143,);
nor I_2395 (I43598,I43251,I43533);
nor I_2396 (I43131,I43446,I43598);
nor I_2397 (I43140,I43381,I43516);
nor I_2398 (I43128,I43251,I43516);
not I_2399 (I43684,I2866);
DFFARX1 I_2400 (I151952,I2859,I43684,I43710,);
not I_2401 (I43718,I43710);
nand I_2402 (I43735,I151934,I151949);
and I_2403 (I43752,I43735,I151925);
DFFARX1 I_2404 (I43752,I2859,I43684,I43778,);
DFFARX1 I_2405 (I151928,I2859,I43684,I43795,);
and I_2406 (I43803,I43795,I151943);
nor I_2407 (I43820,I43778,I43803);
DFFARX1 I_2408 (I43820,I2859,I43684,I43652,);
nand I_2409 (I43851,I43795,I151943);
nand I_2410 (I43868,I43718,I43851);
not I_2411 (I43664,I43868);
DFFARX1 I_2412 (I151946,I2859,I43684,I43908,);
DFFARX1 I_2413 (I43908,I2859,I43684,I43673,);
nand I_2414 (I43930,I151925,I151937);
and I_2415 (I43947,I43930,I151931);
DFFARX1 I_2416 (I43947,I2859,I43684,I43973,);
DFFARX1 I_2417 (I43973,I2859,I43684,I43990,);
not I_2418 (I43676,I43990);
not I_2419 (I44012,I43973);
nand I_2420 (I43661,I44012,I43851);
nor I_2421 (I44043,I151940,I151937);
not I_2422 (I44060,I44043);
nor I_2423 (I44077,I44012,I44060);
nor I_2424 (I44094,I43718,I44077);
DFFARX1 I_2425 (I44094,I2859,I43684,I43670,);
nor I_2426 (I44125,I43778,I44060);
nor I_2427 (I43658,I43973,I44125);
nor I_2428 (I43667,I43908,I44043);
nor I_2429 (I43655,I43778,I44043);
not I_2430 (I44211,I2866);
DFFARX1 I_2431 (I406118,I2859,I44211,I44237,);
not I_2432 (I44245,I44237);
nand I_2433 (I44262,I406136,I406130);
and I_2434 (I44279,I44262,I406109);
DFFARX1 I_2435 (I44279,I2859,I44211,I44305,);
DFFARX1 I_2436 (I406127,I2859,I44211,I44322,);
and I_2437 (I44330,I44322,I406112);
nor I_2438 (I44347,I44305,I44330);
DFFARX1 I_2439 (I44347,I2859,I44211,I44179,);
nand I_2440 (I44378,I44322,I406112);
nand I_2441 (I44395,I44245,I44378);
not I_2442 (I44191,I44395);
DFFARX1 I_2443 (I406124,I2859,I44211,I44435,);
DFFARX1 I_2444 (I44435,I2859,I44211,I44200,);
nand I_2445 (I44457,I406133,I406121);
and I_2446 (I44474,I44457,I406115);
DFFARX1 I_2447 (I44474,I2859,I44211,I44500,);
DFFARX1 I_2448 (I44500,I2859,I44211,I44517,);
not I_2449 (I44203,I44517);
not I_2450 (I44539,I44500);
nand I_2451 (I44188,I44539,I44378);
nor I_2452 (I44570,I406109,I406121);
not I_2453 (I44587,I44570);
nor I_2454 (I44604,I44539,I44587);
nor I_2455 (I44621,I44245,I44604);
DFFARX1 I_2456 (I44621,I2859,I44211,I44197,);
nor I_2457 (I44652,I44305,I44587);
nor I_2458 (I44185,I44500,I44652);
nor I_2459 (I44194,I44435,I44570);
nor I_2460 (I44182,I44305,I44570);
not I_2461 (I44738,I2866);
DFFARX1 I_2462 (I164073,I2859,I44738,I44764,);
not I_2463 (I44772,I44764);
nand I_2464 (I44789,I164055,I164070);
and I_2465 (I44806,I44789,I164046);
DFFARX1 I_2466 (I44806,I2859,I44738,I44832,);
DFFARX1 I_2467 (I164049,I2859,I44738,I44849,);
and I_2468 (I44857,I44849,I164064);
nor I_2469 (I44874,I44832,I44857);
DFFARX1 I_2470 (I44874,I2859,I44738,I44706,);
nand I_2471 (I44905,I44849,I164064);
nand I_2472 (I44922,I44772,I44905);
not I_2473 (I44718,I44922);
DFFARX1 I_2474 (I164067,I2859,I44738,I44962,);
DFFARX1 I_2475 (I44962,I2859,I44738,I44727,);
nand I_2476 (I44984,I164046,I164058);
and I_2477 (I45001,I44984,I164052);
DFFARX1 I_2478 (I45001,I2859,I44738,I45027,);
DFFARX1 I_2479 (I45027,I2859,I44738,I45044,);
not I_2480 (I44730,I45044);
not I_2481 (I45066,I45027);
nand I_2482 (I44715,I45066,I44905);
nor I_2483 (I45097,I164061,I164058);
not I_2484 (I45114,I45097);
nor I_2485 (I45131,I45066,I45114);
nor I_2486 (I45148,I44772,I45131);
DFFARX1 I_2487 (I45148,I2859,I44738,I44724,);
nor I_2488 (I45179,I44832,I45114);
nor I_2489 (I44712,I45027,I45179);
nor I_2490 (I44721,I44962,I45097);
nor I_2491 (I44709,I44832,I45097);
not I_2492 (I45265,I2866);
DFFARX1 I_2493 (I441030,I2859,I45265,I45291,);
not I_2494 (I45299,I45291);
nand I_2495 (I45316,I441027,I441033);
and I_2496 (I45333,I45316,I441030);
DFFARX1 I_2497 (I45333,I2859,I45265,I45359,);
DFFARX1 I_2498 (I441033,I2859,I45265,I45376,);
and I_2499 (I45384,I45376,I441027);
nor I_2500 (I45401,I45359,I45384);
DFFARX1 I_2501 (I45401,I2859,I45265,I45233,);
nand I_2502 (I45432,I45376,I441027);
nand I_2503 (I45449,I45299,I45432);
not I_2504 (I45245,I45449);
DFFARX1 I_2505 (I441036,I2859,I45265,I45489,);
DFFARX1 I_2506 (I45489,I2859,I45265,I45254,);
nand I_2507 (I45511,I441039,I441048);
and I_2508 (I45528,I45511,I441042);
DFFARX1 I_2509 (I45528,I2859,I45265,I45554,);
DFFARX1 I_2510 (I45554,I2859,I45265,I45571,);
not I_2511 (I45257,I45571);
not I_2512 (I45593,I45554);
nand I_2513 (I45242,I45593,I45432);
nor I_2514 (I45624,I441045,I441048);
not I_2515 (I45641,I45624);
nor I_2516 (I45658,I45593,I45641);
nor I_2517 (I45675,I45299,I45658);
DFFARX1 I_2518 (I45675,I2859,I45265,I45251,);
nor I_2519 (I45706,I45359,I45641);
nor I_2520 (I45239,I45554,I45706);
nor I_2521 (I45248,I45489,I45624);
nor I_2522 (I45236,I45359,I45624);
not I_2523 (I45792,I2866);
DFFARX1 I_2524 (I481850,I2859,I45792,I45818,);
not I_2525 (I45826,I45818);
nand I_2526 (I45843,I481865,I481844);
and I_2527 (I45860,I45843,I481847);
DFFARX1 I_2528 (I45860,I2859,I45792,I45886,);
DFFARX1 I_2529 (I481868,I2859,I45792,I45903,);
and I_2530 (I45911,I45903,I481847);
nor I_2531 (I45928,I45886,I45911);
DFFARX1 I_2532 (I45928,I2859,I45792,I45760,);
nand I_2533 (I45959,I45903,I481847);
nand I_2534 (I45976,I45826,I45959);
not I_2535 (I45772,I45976);
DFFARX1 I_2536 (I481844,I2859,I45792,I46016,);
DFFARX1 I_2537 (I46016,I2859,I45792,I45781,);
nand I_2538 (I46038,I481856,I481853);
and I_2539 (I46055,I46038,I481859);
DFFARX1 I_2540 (I46055,I2859,I45792,I46081,);
DFFARX1 I_2541 (I46081,I2859,I45792,I46098,);
not I_2542 (I45784,I46098);
not I_2543 (I46120,I46081);
nand I_2544 (I45769,I46120,I45959);
nor I_2545 (I46151,I481862,I481853);
not I_2546 (I46168,I46151);
nor I_2547 (I46185,I46120,I46168);
nor I_2548 (I46202,I45826,I46185);
DFFARX1 I_2549 (I46202,I2859,I45792,I45778,);
nor I_2550 (I46233,I45886,I46168);
nor I_2551 (I45766,I46081,I46233);
nor I_2552 (I45775,I46016,I46151);
nor I_2553 (I45763,I45886,I46151);
not I_2554 (I46319,I2866);
DFFARX1 I_2555 (I569882,I2859,I46319,I46345,);
not I_2556 (I46353,I46345);
nand I_2557 (I46370,I569876,I569897);
and I_2558 (I46387,I46370,I569873);
DFFARX1 I_2559 (I46387,I2859,I46319,I46413,);
DFFARX1 I_2560 (I569894,I2859,I46319,I46430,);
and I_2561 (I46438,I46430,I569891);
nor I_2562 (I46455,I46413,I46438);
DFFARX1 I_2563 (I46455,I2859,I46319,I46287,);
nand I_2564 (I46486,I46430,I569891);
nand I_2565 (I46503,I46353,I46486);
not I_2566 (I46299,I46503);
DFFARX1 I_2567 (I569879,I2859,I46319,I46543,);
DFFARX1 I_2568 (I46543,I2859,I46319,I46308,);
nand I_2569 (I46565,I569888,I569885);
and I_2570 (I46582,I46565,I569870);
DFFARX1 I_2571 (I46582,I2859,I46319,I46608,);
DFFARX1 I_2572 (I46608,I2859,I46319,I46625,);
not I_2573 (I46311,I46625);
not I_2574 (I46647,I46608);
nand I_2575 (I46296,I46647,I46486);
nor I_2576 (I46678,I569870,I569885);
not I_2577 (I46695,I46678);
nor I_2578 (I46712,I46647,I46695);
nor I_2579 (I46729,I46353,I46712);
DFFARX1 I_2580 (I46729,I2859,I46319,I46305,);
nor I_2581 (I46760,I46413,I46695);
nor I_2582 (I46293,I46608,I46760);
nor I_2583 (I46302,I46543,I46678);
nor I_2584 (I46290,I46413,I46678);
not I_2585 (I46846,I2866);
DFFARX1 I_2586 (I566907,I2859,I46846,I46872,);
not I_2587 (I46880,I46872);
nand I_2588 (I46897,I566901,I566922);
and I_2589 (I46914,I46897,I566898);
DFFARX1 I_2590 (I46914,I2859,I46846,I46940,);
DFFARX1 I_2591 (I566919,I2859,I46846,I46957,);
and I_2592 (I46965,I46957,I566916);
nor I_2593 (I46982,I46940,I46965);
DFFARX1 I_2594 (I46982,I2859,I46846,I46814,);
nand I_2595 (I47013,I46957,I566916);
nand I_2596 (I47030,I46880,I47013);
not I_2597 (I46826,I47030);
DFFARX1 I_2598 (I566904,I2859,I46846,I47070,);
DFFARX1 I_2599 (I47070,I2859,I46846,I46835,);
nand I_2600 (I47092,I566913,I566910);
and I_2601 (I47109,I47092,I566895);
DFFARX1 I_2602 (I47109,I2859,I46846,I47135,);
DFFARX1 I_2603 (I47135,I2859,I46846,I47152,);
not I_2604 (I46838,I47152);
not I_2605 (I47174,I47135);
nand I_2606 (I46823,I47174,I47013);
nor I_2607 (I47205,I566895,I566910);
not I_2608 (I47222,I47205);
nor I_2609 (I47239,I47174,I47222);
nor I_2610 (I47256,I46880,I47239);
DFFARX1 I_2611 (I47256,I2859,I46846,I46832,);
nor I_2612 (I47287,I46940,I47222);
nor I_2613 (I46820,I47135,I47287);
nor I_2614 (I46829,I47070,I47205);
nor I_2615 (I46817,I46940,I47205);
not I_2616 (I47373,I2866);
DFFARX1 I_2617 (I357957,I2859,I47373,I47399,);
not I_2618 (I47407,I47399);
nand I_2619 (I47424,I357954,I357969);
and I_2620 (I47441,I47424,I357951);
DFFARX1 I_2621 (I47441,I2859,I47373,I47467,);
DFFARX1 I_2622 (I357948,I2859,I47373,I47484,);
and I_2623 (I47492,I47484,I357948);
nor I_2624 (I47509,I47467,I47492);
DFFARX1 I_2625 (I47509,I2859,I47373,I47341,);
nand I_2626 (I47540,I47484,I357948);
nand I_2627 (I47557,I47407,I47540);
not I_2628 (I47353,I47557);
DFFARX1 I_2629 (I357951,I2859,I47373,I47597,);
DFFARX1 I_2630 (I47597,I2859,I47373,I47362,);
nand I_2631 (I47619,I357963,I357954);
and I_2632 (I47636,I47619,I357966);
DFFARX1 I_2633 (I47636,I2859,I47373,I47662,);
DFFARX1 I_2634 (I47662,I2859,I47373,I47679,);
not I_2635 (I47365,I47679);
not I_2636 (I47701,I47662);
nand I_2637 (I47350,I47701,I47540);
nor I_2638 (I47732,I357960,I357954);
not I_2639 (I47749,I47732);
nor I_2640 (I47766,I47701,I47749);
nor I_2641 (I47783,I47407,I47766);
DFFARX1 I_2642 (I47783,I2859,I47373,I47359,);
nor I_2643 (I47814,I47467,I47749);
nor I_2644 (I47347,I47662,I47814);
nor I_2645 (I47356,I47597,I47732);
nor I_2646 (I47344,I47467,I47732);
not I_2647 (I47900,I2866);
DFFARX1 I_2648 (I397074,I2859,I47900,I47926,);
not I_2649 (I47934,I47926);
nand I_2650 (I47951,I397092,I397086);
and I_2651 (I47968,I47951,I397065);
DFFARX1 I_2652 (I47968,I2859,I47900,I47994,);
DFFARX1 I_2653 (I397083,I2859,I47900,I48011,);
and I_2654 (I48019,I48011,I397068);
nor I_2655 (I48036,I47994,I48019);
DFFARX1 I_2656 (I48036,I2859,I47900,I47868,);
nand I_2657 (I48067,I48011,I397068);
nand I_2658 (I48084,I47934,I48067);
not I_2659 (I47880,I48084);
DFFARX1 I_2660 (I397080,I2859,I47900,I48124,);
DFFARX1 I_2661 (I48124,I2859,I47900,I47889,);
nand I_2662 (I48146,I397089,I397077);
and I_2663 (I48163,I48146,I397071);
DFFARX1 I_2664 (I48163,I2859,I47900,I48189,);
DFFARX1 I_2665 (I48189,I2859,I47900,I48206,);
not I_2666 (I47892,I48206);
not I_2667 (I48228,I48189);
nand I_2668 (I47877,I48228,I48067);
nor I_2669 (I48259,I397065,I397077);
not I_2670 (I48276,I48259);
nor I_2671 (I48293,I48228,I48276);
nor I_2672 (I48310,I47934,I48293);
DFFARX1 I_2673 (I48310,I2859,I47900,I47886,);
nor I_2674 (I48341,I47994,I48276);
nor I_2675 (I47874,I48189,I48341);
nor I_2676 (I47883,I48124,I48259);
nor I_2677 (I47871,I47994,I48259);
not I_2678 (I48427,I2866);
DFFARX1 I_2679 (I258099,I2859,I48427,I48453,);
not I_2680 (I48461,I48453);
nand I_2681 (I48478,I258111,I258096);
and I_2682 (I48495,I48478,I258090);
DFFARX1 I_2683 (I48495,I2859,I48427,I48521,);
DFFARX1 I_2684 (I258105,I2859,I48427,I48538,);
and I_2685 (I48546,I48538,I258093);
nor I_2686 (I48563,I48521,I48546);
DFFARX1 I_2687 (I48563,I2859,I48427,I48395,);
nand I_2688 (I48594,I48538,I258093);
nand I_2689 (I48611,I48461,I48594);
not I_2690 (I48407,I48611);
DFFARX1 I_2691 (I258102,I2859,I48427,I48651,);
DFFARX1 I_2692 (I48651,I2859,I48427,I48416,);
nand I_2693 (I48673,I258108,I258114);
and I_2694 (I48690,I48673,I258090);
DFFARX1 I_2695 (I48690,I2859,I48427,I48716,);
DFFARX1 I_2696 (I48716,I2859,I48427,I48733,);
not I_2697 (I48419,I48733);
not I_2698 (I48755,I48716);
nand I_2699 (I48404,I48755,I48594);
nor I_2700 (I48786,I258093,I258114);
not I_2701 (I48803,I48786);
nor I_2702 (I48820,I48755,I48803);
nor I_2703 (I48837,I48461,I48820);
DFFARX1 I_2704 (I48837,I2859,I48427,I48413,);
nor I_2705 (I48868,I48521,I48803);
nor I_2706 (I48401,I48716,I48868);
nor I_2707 (I48410,I48651,I48786);
nor I_2708 (I48398,I48521,I48786);
not I_2709 (I48954,I2866);
DFFARX1 I_2710 (I488208,I2859,I48954,I48980,);
not I_2711 (I48988,I48980);
nand I_2712 (I49005,I488223,I488202);
and I_2713 (I49022,I49005,I488205);
DFFARX1 I_2714 (I49022,I2859,I48954,I49048,);
DFFARX1 I_2715 (I488226,I2859,I48954,I49065,);
and I_2716 (I49073,I49065,I488205);
nor I_2717 (I49090,I49048,I49073);
DFFARX1 I_2718 (I49090,I2859,I48954,I48922,);
nand I_2719 (I49121,I49065,I488205);
nand I_2720 (I49138,I48988,I49121);
not I_2721 (I48934,I49138);
DFFARX1 I_2722 (I488202,I2859,I48954,I49178,);
DFFARX1 I_2723 (I49178,I2859,I48954,I48943,);
nand I_2724 (I49200,I488214,I488211);
and I_2725 (I49217,I49200,I488217);
DFFARX1 I_2726 (I49217,I2859,I48954,I49243,);
DFFARX1 I_2727 (I49243,I2859,I48954,I49260,);
not I_2728 (I48946,I49260);
not I_2729 (I49282,I49243);
nand I_2730 (I48931,I49282,I49121);
nor I_2731 (I49313,I488220,I488211);
not I_2732 (I49330,I49313);
nor I_2733 (I49347,I49282,I49330);
nor I_2734 (I49364,I48988,I49347);
DFFARX1 I_2735 (I49364,I2859,I48954,I48940,);
nor I_2736 (I49395,I49048,I49330);
nor I_2737 (I48928,I49243,I49395);
nor I_2738 (I48937,I49178,I49313);
nor I_2739 (I48925,I49048,I49313);
not I_2740 (I49481,I2866);
DFFARX1 I_2741 (I106020,I2859,I49481,I49507,);
not I_2742 (I49515,I49507);
nand I_2743 (I49532,I106014,I106008);
and I_2744 (I49549,I49532,I106029);
DFFARX1 I_2745 (I49549,I2859,I49481,I49575,);
DFFARX1 I_2746 (I106026,I2859,I49481,I49592,);
and I_2747 (I49600,I49592,I106023);
nor I_2748 (I49617,I49575,I49600);
DFFARX1 I_2749 (I49617,I2859,I49481,I49449,);
nand I_2750 (I49648,I49592,I106023);
nand I_2751 (I49665,I49515,I49648);
not I_2752 (I49461,I49665);
DFFARX1 I_2753 (I106008,I2859,I49481,I49705,);
DFFARX1 I_2754 (I49705,I2859,I49481,I49470,);
nand I_2755 (I49727,I106011,I106011);
and I_2756 (I49744,I49727,I106032);
DFFARX1 I_2757 (I49744,I2859,I49481,I49770,);
DFFARX1 I_2758 (I49770,I2859,I49481,I49787,);
not I_2759 (I49473,I49787);
not I_2760 (I49809,I49770);
nand I_2761 (I49458,I49809,I49648);
nor I_2762 (I49840,I106017,I106011);
not I_2763 (I49857,I49840);
nor I_2764 (I49874,I49809,I49857);
nor I_2765 (I49891,I49515,I49874);
DFFARX1 I_2766 (I49891,I2859,I49481,I49467,);
nor I_2767 (I49922,I49575,I49857);
nor I_2768 (I49455,I49770,I49922);
nor I_2769 (I49464,I49705,I49840);
nor I_2770 (I49452,I49575,I49840);
not I_2771 (I50008,I2866);
DFFARX1 I_2772 (I199917,I2859,I50008,I50034,);
not I_2773 (I50042,I50034);
nand I_2774 (I50059,I199911,I199902);
and I_2775 (I50076,I50059,I199923);
DFFARX1 I_2776 (I50076,I2859,I50008,I50102,);
DFFARX1 I_2777 (I199905,I2859,I50008,I50119,);
and I_2778 (I50127,I50119,I199899);
nor I_2779 (I50144,I50102,I50127);
DFFARX1 I_2780 (I50144,I2859,I50008,I49976,);
nand I_2781 (I50175,I50119,I199899);
nand I_2782 (I50192,I50042,I50175);
not I_2783 (I49988,I50192);
DFFARX1 I_2784 (I199899,I2859,I50008,I50232,);
DFFARX1 I_2785 (I50232,I2859,I50008,I49997,);
nand I_2786 (I50254,I199926,I199908);
and I_2787 (I50271,I50254,I199914);
DFFARX1 I_2788 (I50271,I2859,I50008,I50297,);
DFFARX1 I_2789 (I50297,I2859,I50008,I50314,);
not I_2790 (I50000,I50314);
not I_2791 (I50336,I50297);
nand I_2792 (I49985,I50336,I50175);
nor I_2793 (I50367,I199920,I199908);
not I_2794 (I50384,I50367);
nor I_2795 (I50401,I50336,I50384);
nor I_2796 (I50418,I50042,I50401);
DFFARX1 I_2797 (I50418,I2859,I50008,I49994,);
nor I_2798 (I50449,I50102,I50384);
nor I_2799 (I49982,I50297,I50449);
nor I_2800 (I49991,I50232,I50367);
nor I_2801 (I49979,I50102,I50367);
not I_2802 (I50535,I2866);
DFFARX1 I_2803 (I565122,I2859,I50535,I50561,);
not I_2804 (I50569,I50561);
nand I_2805 (I50586,I565116,I565137);
and I_2806 (I50603,I50586,I565113);
DFFARX1 I_2807 (I50603,I2859,I50535,I50629,);
DFFARX1 I_2808 (I565134,I2859,I50535,I50646,);
and I_2809 (I50654,I50646,I565131);
nor I_2810 (I50671,I50629,I50654);
DFFARX1 I_2811 (I50671,I2859,I50535,I50503,);
nand I_2812 (I50702,I50646,I565131);
nand I_2813 (I50719,I50569,I50702);
not I_2814 (I50515,I50719);
DFFARX1 I_2815 (I565119,I2859,I50535,I50759,);
DFFARX1 I_2816 (I50759,I2859,I50535,I50524,);
nand I_2817 (I50781,I565128,I565125);
and I_2818 (I50798,I50781,I565110);
DFFARX1 I_2819 (I50798,I2859,I50535,I50824,);
DFFARX1 I_2820 (I50824,I2859,I50535,I50841,);
not I_2821 (I50527,I50841);
not I_2822 (I50863,I50824);
nand I_2823 (I50512,I50863,I50702);
nor I_2824 (I50894,I565110,I565125);
not I_2825 (I50911,I50894);
nor I_2826 (I50928,I50863,I50911);
nor I_2827 (I50945,I50569,I50928);
DFFARX1 I_2828 (I50945,I2859,I50535,I50521,);
nor I_2829 (I50976,I50629,I50911);
nor I_2830 (I50509,I50824,I50976);
nor I_2831 (I50518,I50759,I50894);
nor I_2832 (I50506,I50629,I50894);
not I_2833 (I51062,I2866);
DFFARX1 I_2834 (I399012,I2859,I51062,I51088,);
not I_2835 (I51096,I51088);
nand I_2836 (I51113,I399030,I399024);
and I_2837 (I51130,I51113,I399003);
DFFARX1 I_2838 (I51130,I2859,I51062,I51156,);
DFFARX1 I_2839 (I399021,I2859,I51062,I51173,);
and I_2840 (I51181,I51173,I399006);
nor I_2841 (I51198,I51156,I51181);
DFFARX1 I_2842 (I51198,I2859,I51062,I51030,);
nand I_2843 (I51229,I51173,I399006);
nand I_2844 (I51246,I51096,I51229);
not I_2845 (I51042,I51246);
DFFARX1 I_2846 (I399018,I2859,I51062,I51286,);
DFFARX1 I_2847 (I51286,I2859,I51062,I51051,);
nand I_2848 (I51308,I399027,I399015);
and I_2849 (I51325,I51308,I399009);
DFFARX1 I_2850 (I51325,I2859,I51062,I51351,);
DFFARX1 I_2851 (I51351,I2859,I51062,I51368,);
not I_2852 (I51054,I51368);
not I_2853 (I51390,I51351);
nand I_2854 (I51039,I51390,I51229);
nor I_2855 (I51421,I399003,I399015);
not I_2856 (I51438,I51421);
nor I_2857 (I51455,I51390,I51438);
nor I_2858 (I51472,I51096,I51455);
DFFARX1 I_2859 (I51472,I2859,I51062,I51048,);
nor I_2860 (I51503,I51156,I51438);
nor I_2861 (I51036,I51351,I51503);
nor I_2862 (I51045,I51286,I51421);
nor I_2863 (I51033,I51156,I51421);
not I_2864 (I51589,I2866);
DFFARX1 I_2865 (I489364,I2859,I51589,I51615,);
not I_2866 (I51623,I51615);
nand I_2867 (I51640,I489379,I489358);
and I_2868 (I51657,I51640,I489361);
DFFARX1 I_2869 (I51657,I2859,I51589,I51683,);
DFFARX1 I_2870 (I489382,I2859,I51589,I51700,);
and I_2871 (I51708,I51700,I489361);
nor I_2872 (I51725,I51683,I51708);
DFFARX1 I_2873 (I51725,I2859,I51589,I51557,);
nand I_2874 (I51756,I51700,I489361);
nand I_2875 (I51773,I51623,I51756);
not I_2876 (I51569,I51773);
DFFARX1 I_2877 (I489358,I2859,I51589,I51813,);
DFFARX1 I_2878 (I51813,I2859,I51589,I51578,);
nand I_2879 (I51835,I489370,I489367);
and I_2880 (I51852,I51835,I489373);
DFFARX1 I_2881 (I51852,I2859,I51589,I51878,);
DFFARX1 I_2882 (I51878,I2859,I51589,I51895,);
not I_2883 (I51581,I51895);
not I_2884 (I51917,I51878);
nand I_2885 (I51566,I51917,I51756);
nor I_2886 (I51948,I489376,I489367);
not I_2887 (I51965,I51948);
nor I_2888 (I51982,I51917,I51965);
nor I_2889 (I51999,I51623,I51982);
DFFARX1 I_2890 (I51999,I2859,I51589,I51575,);
nor I_2891 (I52030,I51683,I51965);
nor I_2892 (I51563,I51878,I52030);
nor I_2893 (I51572,I51813,I51948);
nor I_2894 (I51560,I51683,I51948);
not I_2895 (I52116,I2866);
DFFARX1 I_2896 (I287580,I2859,I52116,I52142,);
not I_2897 (I52150,I52142);
nand I_2898 (I52167,I287571,I287589);
and I_2899 (I52184,I52167,I287568);
DFFARX1 I_2900 (I52184,I2859,I52116,I52210,);
DFFARX1 I_2901 (I287571,I2859,I52116,I52227,);
and I_2902 (I52235,I52227,I287574);
nor I_2903 (I52252,I52210,I52235);
DFFARX1 I_2904 (I52252,I2859,I52116,I52084,);
nand I_2905 (I52283,I52227,I287574);
nand I_2906 (I52300,I52150,I52283);
not I_2907 (I52096,I52300);
DFFARX1 I_2908 (I287568,I2859,I52116,I52340,);
DFFARX1 I_2909 (I52340,I2859,I52116,I52105,);
nand I_2910 (I52362,I287586,I287577);
and I_2911 (I52379,I52362,I287592);
DFFARX1 I_2912 (I52379,I2859,I52116,I52405,);
DFFARX1 I_2913 (I52405,I2859,I52116,I52422,);
not I_2914 (I52108,I52422);
not I_2915 (I52444,I52405);
nand I_2916 (I52093,I52444,I52283);
nor I_2917 (I52475,I287583,I287577);
not I_2918 (I52492,I52475);
nor I_2919 (I52509,I52444,I52492);
nor I_2920 (I52526,I52150,I52509);
DFFARX1 I_2921 (I52526,I2859,I52116,I52102,);
nor I_2922 (I52557,I52210,I52492);
nor I_2923 (I52090,I52405,I52557);
nor I_2924 (I52099,I52340,I52475);
nor I_2925 (I52087,I52210,I52475);
not I_2926 (I52643,I2866);
DFFARX1 I_2927 (I297984,I2859,I52643,I52669,);
not I_2928 (I52677,I52669);
nand I_2929 (I52694,I297975,I297993);
and I_2930 (I52711,I52694,I297972);
DFFARX1 I_2931 (I52711,I2859,I52643,I52737,);
DFFARX1 I_2932 (I297975,I2859,I52643,I52754,);
and I_2933 (I52762,I52754,I297978);
nor I_2934 (I52779,I52737,I52762);
DFFARX1 I_2935 (I52779,I2859,I52643,I52611,);
nand I_2936 (I52810,I52754,I297978);
nand I_2937 (I52827,I52677,I52810);
not I_2938 (I52623,I52827);
DFFARX1 I_2939 (I297972,I2859,I52643,I52867,);
DFFARX1 I_2940 (I52867,I2859,I52643,I52632,);
nand I_2941 (I52889,I297990,I297981);
and I_2942 (I52906,I52889,I297996);
DFFARX1 I_2943 (I52906,I2859,I52643,I52932,);
DFFARX1 I_2944 (I52932,I2859,I52643,I52949,);
not I_2945 (I52635,I52949);
not I_2946 (I52971,I52932);
nand I_2947 (I52620,I52971,I52810);
nor I_2948 (I53002,I297987,I297981);
not I_2949 (I53019,I53002);
nor I_2950 (I53036,I52971,I53019);
nor I_2951 (I53053,I52677,I53036);
DFFARX1 I_2952 (I53053,I2859,I52643,I52629,);
nor I_2953 (I53084,I52737,I53019);
nor I_2954 (I52617,I52932,I53084);
nor I_2955 (I52626,I52867,I53002);
nor I_2956 (I52614,I52737,I53002);
not I_2957 (I53170,I2866);
DFFARX1 I_2958 (I506976,I2859,I53170,I53196,);
not I_2959 (I53204,I53196);
nand I_2960 (I53221,I506970,I506991);
and I_2961 (I53238,I53221,I506982);
DFFARX1 I_2962 (I53238,I2859,I53170,I53264,);
DFFARX1 I_2963 (I506973,I2859,I53170,I53281,);
and I_2964 (I53289,I53281,I506985);
nor I_2965 (I53306,I53264,I53289);
DFFARX1 I_2966 (I53306,I2859,I53170,I53138,);
nand I_2967 (I53337,I53281,I506985);
nand I_2968 (I53354,I53204,I53337);
not I_2969 (I53150,I53354);
DFFARX1 I_2970 (I506973,I2859,I53170,I53394,);
DFFARX1 I_2971 (I53394,I2859,I53170,I53159,);
nand I_2972 (I53416,I506994,I506979);
and I_2973 (I53433,I53416,I506970);
DFFARX1 I_2974 (I53433,I2859,I53170,I53459,);
DFFARX1 I_2975 (I53459,I2859,I53170,I53476,);
not I_2976 (I53162,I53476);
not I_2977 (I53498,I53459);
nand I_2978 (I53147,I53498,I53337);
nor I_2979 (I53529,I506988,I506979);
not I_2980 (I53546,I53529);
nor I_2981 (I53563,I53498,I53546);
nor I_2982 (I53580,I53204,I53563);
DFFARX1 I_2983 (I53580,I2859,I53170,I53156,);
nor I_2984 (I53611,I53264,I53546);
nor I_2985 (I53144,I53459,I53611);
nor I_2986 (I53153,I53394,I53529);
nor I_2987 (I53141,I53264,I53529);
not I_2988 (I53697,I2866);
DFFARX1 I_2989 (I323994,I2859,I53697,I53723,);
not I_2990 (I53731,I53723);
nand I_2991 (I53748,I323985,I324003);
and I_2992 (I53765,I53748,I323982);
DFFARX1 I_2993 (I53765,I2859,I53697,I53791,);
DFFARX1 I_2994 (I323985,I2859,I53697,I53808,);
and I_2995 (I53816,I53808,I323988);
nor I_2996 (I53833,I53791,I53816);
DFFARX1 I_2997 (I53833,I2859,I53697,I53665,);
nand I_2998 (I53864,I53808,I323988);
nand I_2999 (I53881,I53731,I53864);
not I_3000 (I53677,I53881);
DFFARX1 I_3001 (I323982,I2859,I53697,I53921,);
DFFARX1 I_3002 (I53921,I2859,I53697,I53686,);
nand I_3003 (I53943,I324000,I323991);
and I_3004 (I53960,I53943,I324006);
DFFARX1 I_3005 (I53960,I2859,I53697,I53986,);
DFFARX1 I_3006 (I53986,I2859,I53697,I54003,);
not I_3007 (I53689,I54003);
not I_3008 (I54025,I53986);
nand I_3009 (I53674,I54025,I53864);
nor I_3010 (I54056,I323997,I323991);
not I_3011 (I54073,I54056);
nor I_3012 (I54090,I54025,I54073);
nor I_3013 (I54107,I53731,I54090);
DFFARX1 I_3014 (I54107,I2859,I53697,I53683,);
nor I_3015 (I54138,I53791,I54073);
nor I_3016 (I53671,I53986,I54138);
nor I_3017 (I53680,I53921,I54056);
nor I_3018 (I53668,I53791,I54056);
not I_3019 (I54224,I2866);
DFFARX1 I_3020 (I2484,I2859,I54224,I54250,);
not I_3021 (I54258,I54250);
nand I_3022 (I54275,I2268,I2572);
and I_3023 (I54292,I54275,I1972);
DFFARX1 I_3024 (I54292,I2859,I54224,I54318,);
DFFARX1 I_3025 (I1868,I2859,I54224,I54335,);
and I_3026 (I54343,I54335,I1860);
nor I_3027 (I54360,I54318,I54343);
DFFARX1 I_3028 (I54360,I2859,I54224,I54192,);
nand I_3029 (I54391,I54335,I1860);
nand I_3030 (I54408,I54258,I54391);
not I_3031 (I54204,I54408);
DFFARX1 I_3032 (I1524,I2859,I54224,I54448,);
DFFARX1 I_3033 (I54448,I2859,I54224,I54213,);
nand I_3034 (I54470,I2060,I2788);
and I_3035 (I54487,I54470,I1580);
DFFARX1 I_3036 (I54487,I2859,I54224,I54513,);
DFFARX1 I_3037 (I54513,I2859,I54224,I54530,);
not I_3038 (I54216,I54530);
not I_3039 (I54552,I54513);
nand I_3040 (I54201,I54552,I54391);
nor I_3041 (I54583,I1460,I2788);
not I_3042 (I54600,I54583);
nor I_3043 (I54617,I54552,I54600);
nor I_3044 (I54634,I54258,I54617);
DFFARX1 I_3045 (I54634,I2859,I54224,I54210,);
nor I_3046 (I54665,I54318,I54600);
nor I_3047 (I54198,I54513,I54665);
nor I_3048 (I54207,I54448,I54583);
nor I_3049 (I54195,I54318,I54583);
not I_3050 (I54751,I2866);
DFFARX1 I_3051 (I162492,I2859,I54751,I54777,);
not I_3052 (I54785,I54777);
nand I_3053 (I54802,I162474,I162489);
and I_3054 (I54819,I54802,I162465);
DFFARX1 I_3055 (I54819,I2859,I54751,I54845,);
DFFARX1 I_3056 (I162468,I2859,I54751,I54862,);
and I_3057 (I54870,I54862,I162483);
nor I_3058 (I54887,I54845,I54870);
DFFARX1 I_3059 (I54887,I2859,I54751,I54719,);
nand I_3060 (I54918,I54862,I162483);
nand I_3061 (I54935,I54785,I54918);
not I_3062 (I54731,I54935);
DFFARX1 I_3063 (I162486,I2859,I54751,I54975,);
DFFARX1 I_3064 (I54975,I2859,I54751,I54740,);
nand I_3065 (I54997,I162465,I162477);
and I_3066 (I55014,I54997,I162471);
DFFARX1 I_3067 (I55014,I2859,I54751,I55040,);
DFFARX1 I_3068 (I55040,I2859,I54751,I55057,);
not I_3069 (I54743,I55057);
not I_3070 (I55079,I55040);
nand I_3071 (I54728,I55079,I54918);
nor I_3072 (I55110,I162480,I162477);
not I_3073 (I55127,I55110);
nor I_3074 (I55144,I55079,I55127);
nor I_3075 (I55161,I54785,I55144);
DFFARX1 I_3076 (I55161,I2859,I54751,I54737,);
nor I_3077 (I55192,I54845,I55127);
nor I_3078 (I54725,I55040,I55192);
nor I_3079 (I54734,I54975,I55110);
nor I_3080 (I54722,I54845,I55110);
not I_3081 (I55278,I2866);
DFFARX1 I_3082 (I454106,I2859,I55278,I55304,);
not I_3083 (I55312,I55304);
nand I_3084 (I55329,I454121,I454100);
and I_3085 (I55346,I55329,I454103);
DFFARX1 I_3086 (I55346,I2859,I55278,I55372,);
DFFARX1 I_3087 (I454124,I2859,I55278,I55389,);
and I_3088 (I55397,I55389,I454103);
nor I_3089 (I55414,I55372,I55397);
DFFARX1 I_3090 (I55414,I2859,I55278,I55246,);
nand I_3091 (I55445,I55389,I454103);
nand I_3092 (I55462,I55312,I55445);
not I_3093 (I55258,I55462);
DFFARX1 I_3094 (I454100,I2859,I55278,I55502,);
DFFARX1 I_3095 (I55502,I2859,I55278,I55267,);
nand I_3096 (I55524,I454112,I454109);
and I_3097 (I55541,I55524,I454115);
DFFARX1 I_3098 (I55541,I2859,I55278,I55567,);
DFFARX1 I_3099 (I55567,I2859,I55278,I55584,);
not I_3100 (I55270,I55584);
not I_3101 (I55606,I55567);
nand I_3102 (I55255,I55606,I55445);
nor I_3103 (I55637,I454118,I454109);
not I_3104 (I55654,I55637);
nor I_3105 (I55671,I55606,I55654);
nor I_3106 (I55688,I55312,I55671);
DFFARX1 I_3107 (I55688,I2859,I55278,I55264,);
nor I_3108 (I55719,I55372,I55654);
nor I_3109 (I55252,I55567,I55719);
nor I_3110 (I55261,I55502,I55637);
nor I_3111 (I55249,I55372,I55637);
not I_3112 (I55805,I2866);
DFFARX1 I_3113 (I374294,I2859,I55805,I55831,);
not I_3114 (I55839,I55831);
nand I_3115 (I55856,I374291,I374306);
and I_3116 (I55873,I55856,I374288);
DFFARX1 I_3117 (I55873,I2859,I55805,I55899,);
DFFARX1 I_3118 (I374285,I2859,I55805,I55916,);
and I_3119 (I55924,I55916,I374285);
nor I_3120 (I55941,I55899,I55924);
DFFARX1 I_3121 (I55941,I2859,I55805,I55773,);
nand I_3122 (I55972,I55916,I374285);
nand I_3123 (I55989,I55839,I55972);
not I_3124 (I55785,I55989);
DFFARX1 I_3125 (I374288,I2859,I55805,I56029,);
DFFARX1 I_3126 (I56029,I2859,I55805,I55794,);
nand I_3127 (I56051,I374300,I374291);
and I_3128 (I56068,I56051,I374303);
DFFARX1 I_3129 (I56068,I2859,I55805,I56094,);
DFFARX1 I_3130 (I56094,I2859,I55805,I56111,);
not I_3131 (I55797,I56111);
not I_3132 (I56133,I56094);
nand I_3133 (I55782,I56133,I55972);
nor I_3134 (I56164,I374297,I374291);
not I_3135 (I56181,I56164);
nor I_3136 (I56198,I56133,I56181);
nor I_3137 (I56215,I55839,I56198);
DFFARX1 I_3138 (I56215,I2859,I55805,I55791,);
nor I_3139 (I56246,I55899,I56181);
nor I_3140 (I55779,I56094,I56246);
nor I_3141 (I55788,I56029,I56164);
nor I_3142 (I55776,I55899,I56164);
not I_3143 (I56332,I2866);
DFFARX1 I_3144 (I561552,I2859,I56332,I56358,);
not I_3145 (I56366,I56358);
nand I_3146 (I56383,I561546,I561567);
and I_3147 (I56400,I56383,I561543);
DFFARX1 I_3148 (I56400,I2859,I56332,I56426,);
DFFARX1 I_3149 (I561564,I2859,I56332,I56443,);
and I_3150 (I56451,I56443,I561561);
nor I_3151 (I56468,I56426,I56451);
DFFARX1 I_3152 (I56468,I2859,I56332,I56300,);
nand I_3153 (I56499,I56443,I561561);
nand I_3154 (I56516,I56366,I56499);
not I_3155 (I56312,I56516);
DFFARX1 I_3156 (I561549,I2859,I56332,I56556,);
DFFARX1 I_3157 (I56556,I2859,I56332,I56321,);
nand I_3158 (I56578,I561558,I561555);
and I_3159 (I56595,I56578,I561540);
DFFARX1 I_3160 (I56595,I2859,I56332,I56621,);
DFFARX1 I_3161 (I56621,I2859,I56332,I56638,);
not I_3162 (I56324,I56638);
not I_3163 (I56660,I56621);
nand I_3164 (I56309,I56660,I56499);
nor I_3165 (I56691,I561540,I561555);
not I_3166 (I56708,I56691);
nor I_3167 (I56725,I56660,I56708);
nor I_3168 (I56742,I56366,I56725);
DFFARX1 I_3169 (I56742,I2859,I56332,I56318,);
nor I_3170 (I56773,I56426,I56708);
nor I_3171 (I56306,I56621,I56773);
nor I_3172 (I56315,I56556,I56691);
nor I_3173 (I56303,I56426,I56691);
not I_3174 (I56859,I2866);
DFFARX1 I_3175 (I14691,I2859,I56859,I56885,);
not I_3176 (I56893,I56885);
nand I_3177 (I56910,I14679,I14685);
and I_3178 (I56927,I56910,I14688);
DFFARX1 I_3179 (I56927,I2859,I56859,I56953,);
DFFARX1 I_3180 (I14670,I2859,I56859,I56970,);
and I_3181 (I56978,I56970,I14676);
nor I_3182 (I56995,I56953,I56978);
DFFARX1 I_3183 (I56995,I2859,I56859,I56827,);
nand I_3184 (I57026,I56970,I14676);
nand I_3185 (I57043,I56893,I57026);
not I_3186 (I56839,I57043);
DFFARX1 I_3187 (I14670,I2859,I56859,I57083,);
DFFARX1 I_3188 (I57083,I2859,I56859,I56848,);
nand I_3189 (I57105,I14673,I14667);
and I_3190 (I57122,I57105,I14682);
DFFARX1 I_3191 (I57122,I2859,I56859,I57148,);
DFFARX1 I_3192 (I57148,I2859,I56859,I57165,);
not I_3193 (I56851,I57165);
not I_3194 (I57187,I57148);
nand I_3195 (I56836,I57187,I57026);
nor I_3196 (I57218,I14667,I14667);
not I_3197 (I57235,I57218);
nor I_3198 (I57252,I57187,I57235);
nor I_3199 (I57269,I56893,I57252);
DFFARX1 I_3200 (I57269,I2859,I56859,I56845,);
nor I_3201 (I57300,I56953,I57235);
nor I_3202 (I56833,I57148,I57300);
nor I_3203 (I56842,I57083,I57218);
nor I_3204 (I56830,I56953,I57218);
not I_3205 (I57386,I2866);
DFFARX1 I_3206 (I365335,I2859,I57386,I57412,);
not I_3207 (I57420,I57412);
nand I_3208 (I57437,I365332,I365347);
and I_3209 (I57454,I57437,I365329);
DFFARX1 I_3210 (I57454,I2859,I57386,I57480,);
DFFARX1 I_3211 (I365326,I2859,I57386,I57497,);
and I_3212 (I57505,I57497,I365326);
nor I_3213 (I57522,I57480,I57505);
DFFARX1 I_3214 (I57522,I2859,I57386,I57354,);
nand I_3215 (I57553,I57497,I365326);
nand I_3216 (I57570,I57420,I57553);
not I_3217 (I57366,I57570);
DFFARX1 I_3218 (I365329,I2859,I57386,I57610,);
DFFARX1 I_3219 (I57610,I2859,I57386,I57375,);
nand I_3220 (I57632,I365341,I365332);
and I_3221 (I57649,I57632,I365344);
DFFARX1 I_3222 (I57649,I2859,I57386,I57675,);
DFFARX1 I_3223 (I57675,I2859,I57386,I57692,);
not I_3224 (I57378,I57692);
not I_3225 (I57714,I57675);
nand I_3226 (I57363,I57714,I57553);
nor I_3227 (I57745,I365338,I365332);
not I_3228 (I57762,I57745);
nor I_3229 (I57779,I57714,I57762);
nor I_3230 (I57796,I57420,I57779);
DFFARX1 I_3231 (I57796,I2859,I57386,I57372,);
nor I_3232 (I57827,I57480,I57762);
nor I_3233 (I57360,I57675,I57827);
nor I_3234 (I57369,I57610,I57745);
nor I_3235 (I57357,I57480,I57745);
not I_3236 (I57913,I2866);
DFFARX1 I_3237 (I236713,I2859,I57913,I57939,);
not I_3238 (I57947,I57939);
nand I_3239 (I57964,I236725,I236710);
and I_3240 (I57981,I57964,I236704);
DFFARX1 I_3241 (I57981,I2859,I57913,I58007,);
DFFARX1 I_3242 (I236719,I2859,I57913,I58024,);
and I_3243 (I58032,I58024,I236707);
nor I_3244 (I58049,I58007,I58032);
DFFARX1 I_3245 (I58049,I2859,I57913,I57881,);
nand I_3246 (I58080,I58024,I236707);
nand I_3247 (I58097,I57947,I58080);
not I_3248 (I57893,I58097);
DFFARX1 I_3249 (I236716,I2859,I57913,I58137,);
DFFARX1 I_3250 (I58137,I2859,I57913,I57902,);
nand I_3251 (I58159,I236722,I236728);
and I_3252 (I58176,I58159,I236704);
DFFARX1 I_3253 (I58176,I2859,I57913,I58202,);
DFFARX1 I_3254 (I58202,I2859,I57913,I58219,);
not I_3255 (I57905,I58219);
not I_3256 (I58241,I58202);
nand I_3257 (I57890,I58241,I58080);
nor I_3258 (I58272,I236707,I236728);
not I_3259 (I58289,I58272);
nor I_3260 (I58306,I58241,I58289);
nor I_3261 (I58323,I57947,I58306);
DFFARX1 I_3262 (I58323,I2859,I57913,I57899,);
nor I_3263 (I58354,I58007,I58289);
nor I_3264 (I57887,I58202,I58354);
nor I_3265 (I57896,I58137,I58272);
nor I_3266 (I57884,I58007,I58272);
not I_3267 (I58443,I2866);
DFFARX1 I_3268 (I144556,I2859,I58443,I58469,);
not I_3269 (I58477,I58469);
DFFARX1 I_3270 (I144553,I2859,I58443,I58503,);
not I_3271 (I58511,I144550);
or I_3272 (I58528,I144562,I144550);
nor I_3273 (I58545,I58503,I144562);
nand I_3274 (I58420,I58511,I58545);
nor I_3275 (I58576,I144571,I144562);
nand I_3276 (I58414,I58576,I58511);
not I_3277 (I58607,I144568);
nand I_3278 (I58624,I58511,I58607);
nor I_3279 (I58641,I144547,I144547);
not I_3280 (I58658,I58641);
nor I_3281 (I58675,I58658,I58624);
nor I_3282 (I58692,I58576,I58675);
DFFARX1 I_3283 (I58692,I2859,I58443,I58429,);
nor I_3284 (I58426,I58641,I58528);
DFFARX1 I_3285 (I58641,I2859,I58443,I58432,);
nor I_3286 (I58751,I58607,I144547);
nor I_3287 (I58768,I58751,I144550);
nor I_3288 (I58785,I144559,I144574);
DFFARX1 I_3289 (I58785,I2859,I58443,I58811,);
nor I_3290 (I58411,I58811,I58768);
DFFARX1 I_3291 (I58811,I2859,I58443,I58842,);
nand I_3292 (I58850,I58842,I144565);
nor I_3293 (I58435,I58477,I58850);
not I_3294 (I58881,I58811);
nand I_3295 (I58898,I58881,I144565);
nor I_3296 (I58915,I58477,I58898);
nor I_3297 (I58417,I58503,I58915);
nor I_3298 (I58946,I144559,I144571);
nor I_3299 (I58963,I58503,I58946);
DFFARX1 I_3300 (I58963,I2859,I58443,I58408,);
and I_3301 (I58423,I58576,I144559);
not I_3302 (I59038,I2866);
DFFARX1 I_3303 (I371129,I2859,I59038,I59064,);
not I_3304 (I59072,I59064);
DFFARX1 I_3305 (I371129,I2859,I59038,I59098,);
not I_3306 (I59106,I371126);
or I_3307 (I59123,I371138,I371126);
nor I_3308 (I59140,I59098,I371138);
nand I_3309 (I59015,I59106,I59140);
nor I_3310 (I59171,I371132,I371138);
nand I_3311 (I59009,I59171,I59106);
not I_3312 (I59202,I371144);
nand I_3313 (I59219,I59106,I59202);
nor I_3314 (I59236,I371135,I371123);
not I_3315 (I59253,I59236);
nor I_3316 (I59270,I59253,I59219);
nor I_3317 (I59287,I59171,I59270);
DFFARX1 I_3318 (I59287,I2859,I59038,I59024,);
nor I_3319 (I59021,I59236,I59123);
DFFARX1 I_3320 (I59236,I2859,I59038,I59027,);
nor I_3321 (I59346,I59202,I371135);
nor I_3322 (I59363,I59346,I371126);
nor I_3323 (I59380,I371126,I371123);
DFFARX1 I_3324 (I59380,I2859,I59038,I59406,);
nor I_3325 (I59006,I59406,I59363);
DFFARX1 I_3326 (I59406,I2859,I59038,I59437,);
nand I_3327 (I59445,I59437,I371141);
nor I_3328 (I59030,I59072,I59445);
not I_3329 (I59476,I59406);
nand I_3330 (I59493,I59476,I371141);
nor I_3331 (I59510,I59072,I59493);
nor I_3332 (I59012,I59098,I59510);
nor I_3333 (I59541,I371126,I371132);
nor I_3334 (I59558,I59098,I59541);
DFFARX1 I_3335 (I59558,I2859,I59038,I59003,);
and I_3336 (I59018,I59171,I371126);
not I_3337 (I59633,I2866);
DFFARX1 I_3338 (I251169,I2859,I59633,I59659,);
not I_3339 (I59667,I59659);
DFFARX1 I_3340 (I251154,I2859,I59633,I59693,);
not I_3341 (I59701,I251178);
or I_3342 (I59718,I251157,I251178);
nor I_3343 (I59735,I59693,I251157);
nand I_3344 (I59610,I59701,I59735);
nor I_3345 (I59766,I251160,I251157);
nand I_3346 (I59604,I59766,I59701);
not I_3347 (I59797,I251163);
nand I_3348 (I59814,I59701,I59797);
nor I_3349 (I59831,I251166,I251172);
not I_3350 (I59848,I59831);
nor I_3351 (I59865,I59848,I59814);
nor I_3352 (I59882,I59766,I59865);
DFFARX1 I_3353 (I59882,I2859,I59633,I59619,);
nor I_3354 (I59616,I59831,I59718);
DFFARX1 I_3355 (I59831,I2859,I59633,I59622,);
nor I_3356 (I59941,I59797,I251166);
nor I_3357 (I59958,I59941,I251178);
nor I_3358 (I59975,I251175,I251157);
DFFARX1 I_3359 (I59975,I2859,I59633,I60001,);
nor I_3360 (I59601,I60001,I59958);
DFFARX1 I_3361 (I60001,I2859,I59633,I60032,);
nand I_3362 (I60040,I60032,I251154);
nor I_3363 (I59625,I59667,I60040);
not I_3364 (I60071,I60001);
nand I_3365 (I60088,I60071,I251154);
nor I_3366 (I60105,I59667,I60088);
nor I_3367 (I59607,I59693,I60105);
nor I_3368 (I60136,I251175,I251160);
nor I_3369 (I60153,I59693,I60136);
DFFARX1 I_3370 (I60153,I2859,I59633,I59598,);
and I_3371 (I59613,I59766,I251175);
not I_3372 (I60228,I2866);
DFFARX1 I_3373 (I284100,I2859,I60228,I60254,);
not I_3374 (I60262,I60254);
DFFARX1 I_3375 (I284121,I2859,I60228,I60288,);
not I_3376 (I60296,I284100);
or I_3377 (I60313,I284112,I284100);
nor I_3378 (I60330,I60288,I284112);
nand I_3379 (I60205,I60296,I60330);
nor I_3380 (I60361,I284109,I284112);
nand I_3381 (I60199,I60361,I60296);
not I_3382 (I60392,I284118);
nand I_3383 (I60409,I60296,I60392);
nor I_3384 (I60426,I284103,I284103);
not I_3385 (I60443,I60426);
nor I_3386 (I60460,I60443,I60409);
nor I_3387 (I60477,I60361,I60460);
DFFARX1 I_3388 (I60477,I2859,I60228,I60214,);
nor I_3389 (I60211,I60426,I60313);
DFFARX1 I_3390 (I60426,I2859,I60228,I60217,);
nor I_3391 (I60536,I60392,I284103);
nor I_3392 (I60553,I60536,I284100);
nor I_3393 (I60570,I284124,I284106);
DFFARX1 I_3394 (I60570,I2859,I60228,I60596,);
nor I_3395 (I60196,I60596,I60553);
DFFARX1 I_3396 (I60596,I2859,I60228,I60627,);
nand I_3397 (I60635,I60627,I284115);
nor I_3398 (I60220,I60262,I60635);
not I_3399 (I60666,I60596);
nand I_3400 (I60683,I60666,I284115);
nor I_3401 (I60700,I60262,I60683);
nor I_3402 (I60202,I60288,I60700);
nor I_3403 (I60731,I284124,I284109);
nor I_3404 (I60748,I60288,I60731);
DFFARX1 I_3405 (I60748,I2859,I60228,I60193,);
and I_3406 (I60208,I60361,I284124);
not I_3407 (I60823,I2866);
DFFARX1 I_3408 (I521117,I2859,I60823,I60849,);
not I_3409 (I60857,I60849);
DFFARX1 I_3410 (I521114,I2859,I60823,I60883,);
not I_3411 (I60891,I521132);
or I_3412 (I60908,I521126,I521132);
nor I_3413 (I60925,I60883,I521126);
nand I_3414 (I60800,I60891,I60925);
nor I_3415 (I60956,I521120,I521126);
nand I_3416 (I60794,I60956,I60891);
not I_3417 (I60987,I521117);
nand I_3418 (I61004,I60891,I60987);
nor I_3419 (I61021,I521123,I521129);
not I_3420 (I61038,I61021);
nor I_3421 (I61055,I61038,I61004);
nor I_3422 (I61072,I60956,I61055);
DFFARX1 I_3423 (I61072,I2859,I60823,I60809,);
nor I_3424 (I60806,I61021,I60908);
DFFARX1 I_3425 (I61021,I2859,I60823,I60812,);
nor I_3426 (I61131,I60987,I521123);
nor I_3427 (I61148,I61131,I521132);
nor I_3428 (I61165,I521135,I521114);
DFFARX1 I_3429 (I61165,I2859,I60823,I61191,);
nor I_3430 (I60791,I61191,I61148);
DFFARX1 I_3431 (I61191,I2859,I60823,I61222,);
nand I_3432 (I61230,I61222,I521138);
nor I_3433 (I60815,I60857,I61230);
not I_3434 (I61261,I61191);
nand I_3435 (I61278,I61261,I521138);
nor I_3436 (I61295,I60857,I61278);
nor I_3437 (I60797,I60883,I61295);
nor I_3438 (I61326,I521135,I521120);
nor I_3439 (I61343,I60883,I61326);
DFFARX1 I_3440 (I61343,I2859,I60823,I60788,);
and I_3441 (I60803,I60956,I521135);
not I_3442 (I61418,I2866);
DFFARX1 I_3443 (I149299,I2859,I61418,I61444,);
not I_3444 (I61452,I61444);
DFFARX1 I_3445 (I149296,I2859,I61418,I61478,);
not I_3446 (I61486,I149293);
or I_3447 (I61503,I149305,I149293);
nor I_3448 (I61520,I61478,I149305);
nand I_3449 (I61395,I61486,I61520);
nor I_3450 (I61551,I149314,I149305);
nand I_3451 (I61389,I61551,I61486);
not I_3452 (I61582,I149311);
nand I_3453 (I61599,I61486,I61582);
nor I_3454 (I61616,I149290,I149290);
not I_3455 (I61633,I61616);
nor I_3456 (I61650,I61633,I61599);
nor I_3457 (I61667,I61551,I61650);
DFFARX1 I_3458 (I61667,I2859,I61418,I61404,);
nor I_3459 (I61401,I61616,I61503);
DFFARX1 I_3460 (I61616,I2859,I61418,I61407,);
nor I_3461 (I61726,I61582,I149290);
nor I_3462 (I61743,I61726,I149293);
nor I_3463 (I61760,I149302,I149317);
DFFARX1 I_3464 (I61760,I2859,I61418,I61786,);
nor I_3465 (I61386,I61786,I61743);
DFFARX1 I_3466 (I61786,I2859,I61418,I61817,);
nand I_3467 (I61825,I61817,I149308);
nor I_3468 (I61410,I61452,I61825);
not I_3469 (I61856,I61786);
nand I_3470 (I61873,I61856,I149308);
nor I_3471 (I61890,I61452,I61873);
nor I_3472 (I61392,I61478,I61890);
nor I_3473 (I61921,I149302,I149314);
nor I_3474 (I61938,I61478,I61921);
DFFARX1 I_3475 (I61938,I2859,I61418,I61383,);
and I_3476 (I61398,I61551,I149302);
not I_3477 (I62013,I2866);
DFFARX1 I_3478 (I41565,I2859,I62013,I62039,);
not I_3479 (I62047,I62039);
DFFARX1 I_3480 (I41559,I2859,I62013,I62073,);
not I_3481 (I62081,I41568);
or I_3482 (I62098,I41553,I41568);
nor I_3483 (I62115,I62073,I41553);
nand I_3484 (I61990,I62081,I62115);
nor I_3485 (I62146,I41544,I41553);
nand I_3486 (I61984,I62146,I62081);
not I_3487 (I62177,I41544);
nand I_3488 (I62194,I62081,I62177);
nor I_3489 (I62211,I41547,I41562);
not I_3490 (I62228,I62211);
nor I_3491 (I62245,I62228,I62194);
nor I_3492 (I62262,I62146,I62245);
DFFARX1 I_3493 (I62262,I2859,I62013,I61999,);
nor I_3494 (I61996,I62211,I62098);
DFFARX1 I_3495 (I62211,I2859,I62013,I62002,);
nor I_3496 (I62321,I62177,I41547);
nor I_3497 (I62338,I62321,I41568);
nor I_3498 (I62355,I41547,I41556);
DFFARX1 I_3499 (I62355,I2859,I62013,I62381,);
nor I_3500 (I61981,I62381,I62338);
DFFARX1 I_3501 (I62381,I2859,I62013,I62412,);
nand I_3502 (I62420,I62412,I41550);
nor I_3503 (I62005,I62047,I62420);
not I_3504 (I62451,I62381);
nand I_3505 (I62468,I62451,I41550);
nor I_3506 (I62485,I62047,I62468);
nor I_3507 (I61987,I62073,I62485);
nor I_3508 (I62516,I41547,I41544);
nor I_3509 (I62533,I62073,I62516);
DFFARX1 I_3510 (I62533,I2859,I62013,I61978,);
and I_3511 (I61993,I62146,I41547);
not I_3512 (I62605,I2866);
DFFARX1 I_3513 (I148763,I2859,I62605,I62631,);
DFFARX1 I_3514 (I62631,I2859,I62605,I62648,);
not I_3515 (I62597,I62648);
not I_3516 (I62670,I62631);
DFFARX1 I_3517 (I148778,I2859,I62605,I62696,);
not I_3518 (I62704,I62696);
and I_3519 (I62721,I62670,I148775);
not I_3520 (I62738,I148763);
nand I_3521 (I62755,I62738,I148775);
not I_3522 (I62772,I148772);
nor I_3523 (I62789,I62772,I148787);
nand I_3524 (I62806,I62789,I148784);
nor I_3525 (I62823,I62806,I62755);
DFFARX1 I_3526 (I62823,I2859,I62605,I62573,);
not I_3527 (I62854,I62806);
not I_3528 (I62871,I148787);
nand I_3529 (I62888,I62871,I148775);
nor I_3530 (I62905,I148787,I148763);
nand I_3531 (I62585,I62721,I62905);
nand I_3532 (I62579,I62670,I148787);
nand I_3533 (I62950,I62772,I148781);
DFFARX1 I_3534 (I62950,I2859,I62605,I62594,);
DFFARX1 I_3535 (I62950,I2859,I62605,I62588,);
not I_3536 (I62995,I148781);
nor I_3537 (I63012,I62995,I148769);
and I_3538 (I63029,I63012,I148790);
or I_3539 (I63046,I63029,I148766);
DFFARX1 I_3540 (I63046,I2859,I62605,I63072,);
nand I_3541 (I63080,I63072,I62738);
nor I_3542 (I62582,I63080,I62888);
nor I_3543 (I62576,I63072,I62704);
DFFARX1 I_3544 (I63072,I2859,I62605,I63134,);
not I_3545 (I63142,I63134);
nor I_3546 (I62591,I63142,I62854);
not I_3547 (I63200,I2866);
DFFARX1 I_3548 (I5732,I2859,I63200,I63226,);
DFFARX1 I_3549 (I63226,I2859,I63200,I63243,);
not I_3550 (I63192,I63243);
not I_3551 (I63265,I63226);
DFFARX1 I_3552 (I5708,I2859,I63200,I63291,);
not I_3553 (I63299,I63291);
and I_3554 (I63316,I63265,I5723);
not I_3555 (I63333,I5711);
nand I_3556 (I63350,I63333,I5723);
not I_3557 (I63367,I5714);
nor I_3558 (I63384,I63367,I5726);
nand I_3559 (I63401,I63384,I5717);
nor I_3560 (I63418,I63401,I63350);
DFFARX1 I_3561 (I63418,I2859,I63200,I63168,);
not I_3562 (I63449,I63401);
not I_3563 (I63466,I5726);
nand I_3564 (I63483,I63466,I5723);
nor I_3565 (I63500,I5726,I5711);
nand I_3566 (I63180,I63316,I63500);
nand I_3567 (I63174,I63265,I5726);
nand I_3568 (I63545,I63367,I5720);
DFFARX1 I_3569 (I63545,I2859,I63200,I63189,);
DFFARX1 I_3570 (I63545,I2859,I63200,I63183,);
not I_3571 (I63590,I5720);
nor I_3572 (I63607,I63590,I5711);
and I_3573 (I63624,I63607,I5708);
or I_3574 (I63641,I63624,I5729);
DFFARX1 I_3575 (I63641,I2859,I63200,I63667,);
nand I_3576 (I63675,I63667,I63333);
nor I_3577 (I63177,I63675,I63483);
nor I_3578 (I63171,I63667,I63299);
DFFARX1 I_3579 (I63667,I2859,I63200,I63729,);
not I_3580 (I63737,I63729);
nor I_3581 (I63186,I63737,I63449);
not I_3582 (I63795,I2866);
DFFARX1 I_3583 (I156141,I2859,I63795,I63821,);
DFFARX1 I_3584 (I63821,I2859,I63795,I63838,);
not I_3585 (I63787,I63838);
not I_3586 (I63860,I63821);
DFFARX1 I_3587 (I156156,I2859,I63795,I63886,);
not I_3588 (I63894,I63886);
and I_3589 (I63911,I63860,I156153);
not I_3590 (I63928,I156141);
nand I_3591 (I63945,I63928,I156153);
not I_3592 (I63962,I156150);
nor I_3593 (I63979,I63962,I156165);
nand I_3594 (I63996,I63979,I156162);
nor I_3595 (I64013,I63996,I63945);
DFFARX1 I_3596 (I64013,I2859,I63795,I63763,);
not I_3597 (I64044,I63996);
not I_3598 (I64061,I156165);
nand I_3599 (I64078,I64061,I156153);
nor I_3600 (I64095,I156165,I156141);
nand I_3601 (I63775,I63911,I64095);
nand I_3602 (I63769,I63860,I156165);
nand I_3603 (I64140,I63962,I156159);
DFFARX1 I_3604 (I64140,I2859,I63795,I63784,);
DFFARX1 I_3605 (I64140,I2859,I63795,I63778,);
not I_3606 (I64185,I156159);
nor I_3607 (I64202,I64185,I156147);
and I_3608 (I64219,I64202,I156168);
or I_3609 (I64236,I64219,I156144);
DFFARX1 I_3610 (I64236,I2859,I63795,I64262,);
nand I_3611 (I64270,I64262,I63928);
nor I_3612 (I63772,I64270,I64078);
nor I_3613 (I63766,I64262,I63894);
DFFARX1 I_3614 (I64262,I2859,I63795,I64324,);
not I_3615 (I64332,I64324);
nor I_3616 (I63781,I64332,I64044);
not I_3617 (I64390,I2866);
DFFARX1 I_3618 (I495138,I2859,I64390,I64416,);
DFFARX1 I_3619 (I64416,I2859,I64390,I64433,);
not I_3620 (I64382,I64433);
not I_3621 (I64455,I64416);
DFFARX1 I_3622 (I495138,I2859,I64390,I64481,);
not I_3623 (I64489,I64481);
and I_3624 (I64506,I64455,I495141);
not I_3625 (I64523,I495153);
nand I_3626 (I64540,I64523,I495141);
not I_3627 (I64557,I495159);
nor I_3628 (I64574,I64557,I495150);
nand I_3629 (I64591,I64574,I495156);
nor I_3630 (I64608,I64591,I64540);
DFFARX1 I_3631 (I64608,I2859,I64390,I64358,);
not I_3632 (I64639,I64591);
not I_3633 (I64656,I495150);
nand I_3634 (I64673,I64656,I495141);
nor I_3635 (I64690,I495150,I495153);
nand I_3636 (I64370,I64506,I64690);
nand I_3637 (I64364,I64455,I495150);
nand I_3638 (I64735,I64557,I495147);
DFFARX1 I_3639 (I64735,I2859,I64390,I64379,);
DFFARX1 I_3640 (I64735,I2859,I64390,I64373,);
not I_3641 (I64780,I495147);
nor I_3642 (I64797,I64780,I495144);
and I_3643 (I64814,I64797,I495162);
or I_3644 (I64831,I64814,I495141);
DFFARX1 I_3645 (I64831,I2859,I64390,I64857,);
nand I_3646 (I64865,I64857,I64523);
nor I_3647 (I64367,I64865,I64673);
nor I_3648 (I64361,I64857,I64489);
DFFARX1 I_3649 (I64857,I2859,I64390,I64919,);
not I_3650 (I64927,I64919);
nor I_3651 (I64376,I64927,I64639);
not I_3652 (I64985,I2866);
DFFARX1 I_3653 (I549661,I2859,I64985,I65011,);
DFFARX1 I_3654 (I65011,I2859,I64985,I65028,);
not I_3655 (I64977,I65028);
not I_3656 (I65050,I65011);
DFFARX1 I_3657 (I549652,I2859,I64985,I65076,);
not I_3658 (I65084,I65076);
and I_3659 (I65101,I65050,I549646);
not I_3660 (I65118,I549640);
nand I_3661 (I65135,I65118,I549646);
not I_3662 (I65152,I549667);
nor I_3663 (I65169,I65152,I549640);
nand I_3664 (I65186,I65169,I549664);
nor I_3665 (I65203,I65186,I65135);
DFFARX1 I_3666 (I65203,I2859,I64985,I64953,);
not I_3667 (I65234,I65186);
not I_3668 (I65251,I549640);
nand I_3669 (I65268,I65251,I549646);
nor I_3670 (I65285,I549640,I549640);
nand I_3671 (I64965,I65101,I65285);
nand I_3672 (I64959,I65050,I549640);
nand I_3673 (I65330,I65152,I549649);
DFFARX1 I_3674 (I65330,I2859,I64985,I64974,);
DFFARX1 I_3675 (I65330,I2859,I64985,I64968,);
not I_3676 (I65375,I549649);
nor I_3677 (I65392,I65375,I549655);
and I_3678 (I65409,I65392,I549658);
or I_3679 (I65426,I65409,I549643);
DFFARX1 I_3680 (I65426,I2859,I64985,I65452,);
nand I_3681 (I65460,I65452,I65118);
nor I_3682 (I64962,I65460,I65268);
nor I_3683 (I64956,I65452,I65084);
DFFARX1 I_3684 (I65452,I2859,I64985,I65514,);
not I_3685 (I65522,I65514);
nor I_3686 (I64971,I65522,I65234);
not I_3687 (I65580,I2866);
DFFARX1 I_3688 (I191219,I2859,I65580,I65606,);
DFFARX1 I_3689 (I65606,I2859,I65580,I65623,);
not I_3690 (I65572,I65623);
not I_3691 (I65645,I65606);
DFFARX1 I_3692 (I191207,I2859,I65580,I65671,);
not I_3693 (I65679,I65671);
and I_3694 (I65696,I65645,I191216);
not I_3695 (I65713,I191213);
nand I_3696 (I65730,I65713,I191216);
not I_3697 (I65747,I191204);
nor I_3698 (I65764,I65747,I191210);
nand I_3699 (I65781,I65764,I191195);
nor I_3700 (I65798,I65781,I65730);
DFFARX1 I_3701 (I65798,I2859,I65580,I65548,);
not I_3702 (I65829,I65781);
not I_3703 (I65846,I191210);
nand I_3704 (I65863,I65846,I191216);
nor I_3705 (I65880,I191210,I191213);
nand I_3706 (I65560,I65696,I65880);
nand I_3707 (I65554,I65645,I191210);
nand I_3708 (I65925,I65747,I191195);
DFFARX1 I_3709 (I65925,I2859,I65580,I65569,);
DFFARX1 I_3710 (I65925,I2859,I65580,I65563,);
not I_3711 (I65970,I191195);
nor I_3712 (I65987,I65970,I191201);
and I_3713 (I66004,I65987,I191198);
or I_3714 (I66021,I66004,I191222);
DFFARX1 I_3715 (I66021,I2859,I65580,I66047,);
nand I_3716 (I66055,I66047,I65713);
nor I_3717 (I65557,I66055,I65863);
nor I_3718 (I65551,I66047,I65679);
DFFARX1 I_3719 (I66047,I2859,I65580,I66109,);
not I_3720 (I66117,I66109);
nor I_3721 (I65566,I66117,I65829);
not I_3722 (I66175,I2866);
DFFARX1 I_3723 (I112400,I2859,I66175,I66201,);
DFFARX1 I_3724 (I66201,I2859,I66175,I66218,);
not I_3725 (I66167,I66218);
not I_3726 (I66240,I66201);
DFFARX1 I_3727 (I112415,I2859,I66175,I66266,);
not I_3728 (I66274,I66266);
and I_3729 (I66291,I66240,I112412);
not I_3730 (I66308,I112400);
nand I_3731 (I66325,I66308,I112412);
not I_3732 (I66342,I112409);
nor I_3733 (I66359,I66342,I112424);
nand I_3734 (I66376,I66359,I112421);
nor I_3735 (I66393,I66376,I66325);
DFFARX1 I_3736 (I66393,I2859,I66175,I66143,);
not I_3737 (I66424,I66376);
not I_3738 (I66441,I112424);
nand I_3739 (I66458,I66441,I112412);
nor I_3740 (I66475,I112424,I112400);
nand I_3741 (I66155,I66291,I66475);
nand I_3742 (I66149,I66240,I112424);
nand I_3743 (I66520,I66342,I112418);
DFFARX1 I_3744 (I66520,I2859,I66175,I66164,);
DFFARX1 I_3745 (I66520,I2859,I66175,I66158,);
not I_3746 (I66565,I112418);
nor I_3747 (I66582,I66565,I112406);
and I_3748 (I66599,I66582,I112427);
or I_3749 (I66616,I66599,I112403);
DFFARX1 I_3750 (I66616,I2859,I66175,I66642,);
nand I_3751 (I66650,I66642,I66308);
nor I_3752 (I66152,I66650,I66458);
nor I_3753 (I66146,I66642,I66274);
DFFARX1 I_3754 (I66642,I2859,I66175,I66704,);
not I_3755 (I66712,I66704);
nor I_3756 (I66161,I66712,I66424);
not I_3757 (I66770,I2866);
DFFARX1 I_3758 (I245389,I2859,I66770,I66796,);
DFFARX1 I_3759 (I66796,I2859,I66770,I66813,);
not I_3760 (I66762,I66813);
not I_3761 (I66835,I66796);
DFFARX1 I_3762 (I245380,I2859,I66770,I66861,);
not I_3763 (I66869,I66861);
and I_3764 (I66886,I66835,I245398);
not I_3765 (I66903,I245395);
nand I_3766 (I66920,I66903,I245398);
not I_3767 (I66937,I245374);
nor I_3768 (I66954,I66937,I245377);
nand I_3769 (I66971,I66954,I245386);
nor I_3770 (I66988,I66971,I66920);
DFFARX1 I_3771 (I66988,I2859,I66770,I66738,);
not I_3772 (I67019,I66971);
not I_3773 (I67036,I245377);
nand I_3774 (I67053,I67036,I245398);
nor I_3775 (I67070,I245377,I245395);
nand I_3776 (I66750,I66886,I67070);
nand I_3777 (I66744,I66835,I245377);
nand I_3778 (I67115,I66937,I245392);
DFFARX1 I_3779 (I67115,I2859,I66770,I66759,);
DFFARX1 I_3780 (I67115,I2859,I66770,I66753,);
not I_3781 (I67160,I245392);
nor I_3782 (I67177,I67160,I245374);
and I_3783 (I67194,I67177,I245383);
or I_3784 (I67211,I67194,I245377);
DFFARX1 I_3785 (I67211,I2859,I66770,I67237,);
nand I_3786 (I67245,I67237,I66903);
nor I_3787 (I66747,I67245,I67053);
nor I_3788 (I66741,I67237,I66869);
DFFARX1 I_3789 (I67237,I2859,I66770,I67299,);
not I_3790 (I67307,I67299);
nor I_3791 (I66756,I67307,I67019);
not I_3792 (I67365,I2866);
DFFARX1 I_3793 (I2252,I2859,I67365,I67391,);
DFFARX1 I_3794 (I67391,I2859,I67365,I67408,);
not I_3795 (I67357,I67408);
not I_3796 (I67430,I67391);
DFFARX1 I_3797 (I2172,I2859,I67365,I67456,);
not I_3798 (I67464,I67456);
and I_3799 (I67481,I67430,I2236);
not I_3800 (I67498,I2092);
nand I_3801 (I67515,I67498,I2236);
not I_3802 (I67532,I2108);
nor I_3803 (I67549,I67532,I1724);
nand I_3804 (I67566,I67549,I2068);
nor I_3805 (I67583,I67566,I67515);
DFFARX1 I_3806 (I67583,I2859,I67365,I67333,);
not I_3807 (I67614,I67566);
not I_3808 (I67631,I1724);
nand I_3809 (I67648,I67631,I2236);
nor I_3810 (I67665,I1724,I2092);
nand I_3811 (I67345,I67481,I67665);
nand I_3812 (I67339,I67430,I1724);
nand I_3813 (I67710,I67532,I2500);
DFFARX1 I_3814 (I67710,I2859,I67365,I67354,);
DFFARX1 I_3815 (I67710,I2859,I67365,I67348,);
not I_3816 (I67755,I2500);
nor I_3817 (I67772,I67755,I1564);
and I_3818 (I67789,I67772,I2444);
or I_3819 (I67806,I67789,I2364);
DFFARX1 I_3820 (I67806,I2859,I67365,I67832,);
nand I_3821 (I67840,I67832,I67498);
nor I_3822 (I67342,I67840,I67648);
nor I_3823 (I67336,I67832,I67464);
DFFARX1 I_3824 (I67832,I2859,I67365,I67894,);
not I_3825 (I67902,I67894);
nor I_3826 (I67351,I67902,I67614);
not I_3827 (I67960,I2866);
DFFARX1 I_3828 (I334239,I2859,I67960,I67986,);
DFFARX1 I_3829 (I67986,I2859,I67960,I68003,);
not I_3830 (I67952,I68003);
not I_3831 (I68025,I67986);
DFFARX1 I_3832 (I334233,I2859,I67960,I68051,);
not I_3833 (I68059,I68051);
and I_3834 (I68076,I68025,I334251);
not I_3835 (I68093,I334239);
nand I_3836 (I68110,I68093,I334251);
not I_3837 (I68127,I334233);
nor I_3838 (I68144,I68127,I334245);
nand I_3839 (I68161,I68144,I334236);
nor I_3840 (I68178,I68161,I68110);
DFFARX1 I_3841 (I68178,I2859,I67960,I67928,);
not I_3842 (I68209,I68161);
not I_3843 (I68226,I334245);
nand I_3844 (I68243,I68226,I334251);
nor I_3845 (I68260,I334245,I334239);
nand I_3846 (I67940,I68076,I68260);
nand I_3847 (I67934,I68025,I334245);
nand I_3848 (I68305,I68127,I334248);
DFFARX1 I_3849 (I68305,I2859,I67960,I67949,);
DFFARX1 I_3850 (I68305,I2859,I67960,I67943,);
not I_3851 (I68350,I334248);
nor I_3852 (I68367,I68350,I334254);
and I_3853 (I68384,I68367,I334236);
or I_3854 (I68401,I68384,I334242);
DFFARX1 I_3855 (I68401,I2859,I67960,I68427,);
nand I_3856 (I68435,I68427,I68093);
nor I_3857 (I67937,I68435,I68243);
nor I_3858 (I67931,I68427,I68059);
DFFARX1 I_3859 (I68427,I2859,I67960,I68489,);
not I_3860 (I68497,I68489);
nor I_3861 (I67946,I68497,I68209);
not I_3862 (I68555,I2866);
DFFARX1 I_3863 (I360062,I2859,I68555,I68581,);
DFFARX1 I_3864 (I68581,I2859,I68555,I68598,);
not I_3865 (I68547,I68598);
not I_3866 (I68620,I68581);
DFFARX1 I_3867 (I360056,I2859,I68555,I68646,);
not I_3868 (I68654,I68646);
and I_3869 (I68671,I68620,I360074);
not I_3870 (I68688,I360062);
nand I_3871 (I68705,I68688,I360074);
not I_3872 (I68722,I360056);
nor I_3873 (I68739,I68722,I360068);
nand I_3874 (I68756,I68739,I360059);
nor I_3875 (I68773,I68756,I68705);
DFFARX1 I_3876 (I68773,I2859,I68555,I68523,);
not I_3877 (I68804,I68756);
not I_3878 (I68821,I360068);
nand I_3879 (I68838,I68821,I360074);
nor I_3880 (I68855,I360068,I360062);
nand I_3881 (I68535,I68671,I68855);
nand I_3882 (I68529,I68620,I360068);
nand I_3883 (I68900,I68722,I360071);
DFFARX1 I_3884 (I68900,I2859,I68555,I68544,);
DFFARX1 I_3885 (I68900,I2859,I68555,I68538,);
not I_3886 (I68945,I360071);
nor I_3887 (I68962,I68945,I360077);
and I_3888 (I68979,I68962,I360059);
or I_3889 (I68996,I68979,I360065);
DFFARX1 I_3890 (I68996,I2859,I68555,I69022,);
nand I_3891 (I69030,I69022,I68688);
nor I_3892 (I68532,I69030,I68838);
nor I_3893 (I68526,I69022,I68654);
DFFARX1 I_3894 (I69022,I2859,I68555,I69084,);
not I_3895 (I69092,I69084);
nor I_3896 (I68541,I69092,I68804);
not I_3897 (I69150,I2866);
DFFARX1 I_3898 (I295094,I2859,I69150,I69176,);
DFFARX1 I_3899 (I69176,I2859,I69150,I69193,);
not I_3900 (I69142,I69193);
not I_3901 (I69215,I69176);
DFFARX1 I_3902 (I295091,I2859,I69150,I69241,);
not I_3903 (I69249,I69241);
and I_3904 (I69266,I69215,I295097);
not I_3905 (I69283,I295082);
nand I_3906 (I69300,I69283,I295097);
not I_3907 (I69317,I295085);
nor I_3908 (I69334,I69317,I295106);
nand I_3909 (I69351,I69334,I295103);
nor I_3910 (I69368,I69351,I69300);
DFFARX1 I_3911 (I69368,I2859,I69150,I69118,);
not I_3912 (I69399,I69351);
not I_3913 (I69416,I295106);
nand I_3914 (I69433,I69416,I295097);
nor I_3915 (I69450,I295106,I295082);
nand I_3916 (I69130,I69266,I69450);
nand I_3917 (I69124,I69215,I295106);
nand I_3918 (I69495,I69317,I295082);
DFFARX1 I_3919 (I69495,I2859,I69150,I69139,);
DFFARX1 I_3920 (I69495,I2859,I69150,I69133,);
not I_3921 (I69540,I295082);
nor I_3922 (I69557,I69540,I295088);
and I_3923 (I69574,I69557,I295100);
or I_3924 (I69591,I69574,I295085);
DFFARX1 I_3925 (I69591,I2859,I69150,I69617,);
nand I_3926 (I69625,I69617,I69283);
nor I_3927 (I69127,I69625,I69433);
nor I_3928 (I69121,I69617,I69249);
DFFARX1 I_3929 (I69617,I2859,I69150,I69679,);
not I_3930 (I69687,I69679);
nor I_3931 (I69136,I69687,I69399);
not I_3932 (I69745,I2866);
DFFARX1 I_3933 (I318214,I2859,I69745,I69771,);
DFFARX1 I_3934 (I69771,I2859,I69745,I69788,);
not I_3935 (I69737,I69788);
not I_3936 (I69810,I69771);
DFFARX1 I_3937 (I318211,I2859,I69745,I69836,);
not I_3938 (I69844,I69836);
and I_3939 (I69861,I69810,I318217);
not I_3940 (I69878,I318202);
nand I_3941 (I69895,I69878,I318217);
not I_3942 (I69912,I318205);
nor I_3943 (I69929,I69912,I318226);
nand I_3944 (I69946,I69929,I318223);
nor I_3945 (I69963,I69946,I69895);
DFFARX1 I_3946 (I69963,I2859,I69745,I69713,);
not I_3947 (I69994,I69946);
not I_3948 (I70011,I318226);
nand I_3949 (I70028,I70011,I318217);
nor I_3950 (I70045,I318226,I318202);
nand I_3951 (I69725,I69861,I70045);
nand I_3952 (I69719,I69810,I318226);
nand I_3953 (I70090,I69912,I318202);
DFFARX1 I_3954 (I70090,I2859,I69745,I69734,);
DFFARX1 I_3955 (I70090,I2859,I69745,I69728,);
not I_3956 (I70135,I318202);
nor I_3957 (I70152,I70135,I318208);
and I_3958 (I70169,I70152,I318220);
or I_3959 (I70186,I70169,I318205);
DFFARX1 I_3960 (I70186,I2859,I69745,I70212,);
nand I_3961 (I70220,I70212,I69878);
nor I_3962 (I69722,I70220,I70028);
nor I_3963 (I69716,I70212,I69844);
DFFARX1 I_3964 (I70212,I2859,I69745,I70274,);
not I_3965 (I70282,I70274);
nor I_3966 (I69731,I70282,I69994);
not I_3967 (I70340,I2866);
DFFARX1 I_3968 (I393204,I2859,I70340,I70366,);
DFFARX1 I_3969 (I70366,I2859,I70340,I70383,);
not I_3970 (I70332,I70383);
not I_3971 (I70405,I70366);
DFFARX1 I_3972 (I393213,I2859,I70340,I70431,);
not I_3973 (I70439,I70431);
and I_3974 (I70456,I70405,I393201);
not I_3975 (I70473,I393192);
nand I_3976 (I70490,I70473,I393201);
not I_3977 (I70507,I393198);
nor I_3978 (I70524,I70507,I393216);
nand I_3979 (I70541,I70524,I393189);
nor I_3980 (I70558,I70541,I70490);
DFFARX1 I_3981 (I70558,I2859,I70340,I70308,);
not I_3982 (I70589,I70541);
not I_3983 (I70606,I393216);
nand I_3984 (I70623,I70606,I393201);
nor I_3985 (I70640,I393216,I393192);
nand I_3986 (I70320,I70456,I70640);
nand I_3987 (I70314,I70405,I393216);
nand I_3988 (I70685,I70507,I393195);
DFFARX1 I_3989 (I70685,I2859,I70340,I70329,);
DFFARX1 I_3990 (I70685,I2859,I70340,I70323,);
not I_3991 (I70730,I393195);
nor I_3992 (I70747,I70730,I393207);
and I_3993 (I70764,I70747,I393189);
or I_3994 (I70781,I70764,I393210);
DFFARX1 I_3995 (I70781,I2859,I70340,I70807,);
nand I_3996 (I70815,I70807,I70473);
nor I_3997 (I70317,I70815,I70623);
nor I_3998 (I70311,I70807,I70439);
DFFARX1 I_3999 (I70807,I2859,I70340,I70869,);
not I_4000 (I70877,I70869);
nor I_4001 (I70326,I70877,I70589);
not I_4002 (I70935,I2866);
DFFARX1 I_4003 (I165100,I2859,I70935,I70961,);
DFFARX1 I_4004 (I70961,I2859,I70935,I70978,);
not I_4005 (I70927,I70978);
not I_4006 (I71000,I70961);
DFFARX1 I_4007 (I165115,I2859,I70935,I71026,);
not I_4008 (I71034,I71026);
and I_4009 (I71051,I71000,I165112);
not I_4010 (I71068,I165100);
nand I_4011 (I71085,I71068,I165112);
not I_4012 (I71102,I165109);
nor I_4013 (I71119,I71102,I165124);
nand I_4014 (I71136,I71119,I165121);
nor I_4015 (I71153,I71136,I71085);
DFFARX1 I_4016 (I71153,I2859,I70935,I70903,);
not I_4017 (I71184,I71136);
not I_4018 (I71201,I165124);
nand I_4019 (I71218,I71201,I165112);
nor I_4020 (I71235,I165124,I165100);
nand I_4021 (I70915,I71051,I71235);
nand I_4022 (I70909,I71000,I165124);
nand I_4023 (I71280,I71102,I165118);
DFFARX1 I_4024 (I71280,I2859,I70935,I70924,);
DFFARX1 I_4025 (I71280,I2859,I70935,I70918,);
not I_4026 (I71325,I165118);
nor I_4027 (I71342,I71325,I165106);
and I_4028 (I71359,I71342,I165127);
or I_4029 (I71376,I71359,I165103);
DFFARX1 I_4030 (I71376,I2859,I70935,I71402,);
nand I_4031 (I71410,I71402,I71068);
nor I_4032 (I70912,I71410,I71218);
nor I_4033 (I70906,I71402,I71034);
DFFARX1 I_4034 (I71402,I2859,I70935,I71464,);
not I_4035 (I71472,I71464);
nor I_4036 (I70921,I71472,I71184);
not I_4037 (I71530,I2866);
DFFARX1 I_4038 (I424200,I2859,I71530,I71556,);
DFFARX1 I_4039 (I71556,I2859,I71530,I71573,);
not I_4040 (I71522,I71573);
not I_4041 (I71595,I71556);
DFFARX1 I_4042 (I424209,I2859,I71530,I71621,);
not I_4043 (I71629,I71621);
and I_4044 (I71646,I71595,I424203);
not I_4045 (I71663,I424197);
nand I_4046 (I71680,I71663,I424203);
not I_4047 (I71697,I424212);
nor I_4048 (I71714,I71697,I424200);
nand I_4049 (I71731,I71714,I424206);
nor I_4050 (I71748,I71731,I71680);
DFFARX1 I_4051 (I71748,I2859,I71530,I71498,);
not I_4052 (I71779,I71731);
not I_4053 (I71796,I424200);
nand I_4054 (I71813,I71796,I424203);
nor I_4055 (I71830,I424200,I424197);
nand I_4056 (I71510,I71646,I71830);
nand I_4057 (I71504,I71595,I424200);
nand I_4058 (I71875,I71697,I424203);
DFFARX1 I_4059 (I71875,I2859,I71530,I71519,);
DFFARX1 I_4060 (I71875,I2859,I71530,I71513,);
not I_4061 (I71920,I424203);
nor I_4062 (I71937,I71920,I424218);
and I_4063 (I71954,I71937,I424215);
or I_4064 (I71971,I71954,I424197);
DFFARX1 I_4065 (I71971,I2859,I71530,I71997,);
nand I_4066 (I72005,I71997,I71663);
nor I_4067 (I71507,I72005,I71813);
nor I_4068 (I71501,I71997,I71629);
DFFARX1 I_4069 (I71997,I2859,I71530,I72059,);
not I_4070 (I72067,I72059);
nor I_4071 (I71516,I72067,I71779);
not I_4072 (I72125,I2866);
DFFARX1 I_4073 (I345833,I2859,I72125,I72151,);
DFFARX1 I_4074 (I72151,I2859,I72125,I72168,);
not I_4075 (I72117,I72168);
not I_4076 (I72190,I72151);
DFFARX1 I_4077 (I345827,I2859,I72125,I72216,);
not I_4078 (I72224,I72216);
and I_4079 (I72241,I72190,I345845);
not I_4080 (I72258,I345833);
nand I_4081 (I72275,I72258,I345845);
not I_4082 (I72292,I345827);
nor I_4083 (I72309,I72292,I345839);
nand I_4084 (I72326,I72309,I345830);
nor I_4085 (I72343,I72326,I72275);
DFFARX1 I_4086 (I72343,I2859,I72125,I72093,);
not I_4087 (I72374,I72326);
not I_4088 (I72391,I345839);
nand I_4089 (I72408,I72391,I345845);
nor I_4090 (I72425,I345839,I345833);
nand I_4091 (I72105,I72241,I72425);
nand I_4092 (I72099,I72190,I345839);
nand I_4093 (I72470,I72292,I345842);
DFFARX1 I_4094 (I72470,I2859,I72125,I72114,);
DFFARX1 I_4095 (I72470,I2859,I72125,I72108,);
not I_4096 (I72515,I345842);
nor I_4097 (I72532,I72515,I345848);
and I_4098 (I72549,I72532,I345830);
or I_4099 (I72566,I72549,I345836);
DFFARX1 I_4100 (I72566,I2859,I72125,I72592,);
nand I_4101 (I72600,I72592,I72258);
nor I_4102 (I72102,I72600,I72408);
nor I_4103 (I72096,I72592,I72224);
DFFARX1 I_4104 (I72592,I2859,I72125,I72654,);
not I_4105 (I72662,I72654);
nor I_4106 (I72111,I72662,I72374);
not I_4107 (I72720,I2866);
DFFARX1 I_4108 (I359008,I2859,I72720,I72746,);
DFFARX1 I_4109 (I72746,I2859,I72720,I72763,);
not I_4110 (I72712,I72763);
not I_4111 (I72785,I72746);
DFFARX1 I_4112 (I359002,I2859,I72720,I72811,);
not I_4113 (I72819,I72811);
and I_4114 (I72836,I72785,I359020);
not I_4115 (I72853,I359008);
nand I_4116 (I72870,I72853,I359020);
not I_4117 (I72887,I359002);
nor I_4118 (I72904,I72887,I359014);
nand I_4119 (I72921,I72904,I359005);
nor I_4120 (I72938,I72921,I72870);
DFFARX1 I_4121 (I72938,I2859,I72720,I72688,);
not I_4122 (I72969,I72921);
not I_4123 (I72986,I359014);
nand I_4124 (I73003,I72986,I359020);
nor I_4125 (I73020,I359014,I359008);
nand I_4126 (I72700,I72836,I73020);
nand I_4127 (I72694,I72785,I359014);
nand I_4128 (I73065,I72887,I359017);
DFFARX1 I_4129 (I73065,I2859,I72720,I72709,);
DFFARX1 I_4130 (I73065,I2859,I72720,I72703,);
not I_4131 (I73110,I359017);
nor I_4132 (I73127,I73110,I359023);
and I_4133 (I73144,I73127,I359005);
or I_4134 (I73161,I73144,I359011);
DFFARX1 I_4135 (I73161,I2859,I72720,I73187,);
nand I_4136 (I73195,I73187,I72853);
nor I_4137 (I72697,I73195,I73003);
nor I_4138 (I72691,I73187,I72819);
DFFARX1 I_4139 (I73187,I2859,I72720,I73249,);
not I_4140 (I73257,I73249);
nor I_4141 (I72706,I73257,I72969);
not I_4142 (I73315,I2866);
DFFARX1 I_4143 (I225615,I2859,I73315,I73341,);
DFFARX1 I_4144 (I73341,I2859,I73315,I73358,);
not I_4145 (I73307,I73358);
not I_4146 (I73380,I73341);
DFFARX1 I_4147 (I225609,I2859,I73315,I73406,);
not I_4148 (I73414,I73406);
and I_4149 (I73431,I73380,I225624);
not I_4150 (I73448,I225621);
nand I_4151 (I73465,I73448,I225624);
not I_4152 (I73482,I225612);
nor I_4153 (I73499,I73482,I225603);
nand I_4154 (I73516,I73499,I225606);
nor I_4155 (I73533,I73516,I73465);
DFFARX1 I_4156 (I73533,I2859,I73315,I73283,);
not I_4157 (I73564,I73516);
not I_4158 (I73581,I225603);
nand I_4159 (I73598,I73581,I225624);
nor I_4160 (I73615,I225603,I225621);
nand I_4161 (I73295,I73431,I73615);
nand I_4162 (I73289,I73380,I225603);
nand I_4163 (I73660,I73482,I225627);
DFFARX1 I_4164 (I73660,I2859,I73315,I73304,);
DFFARX1 I_4165 (I73660,I2859,I73315,I73298,);
not I_4166 (I73705,I225627);
nor I_4167 (I73722,I73705,I225618);
and I_4168 (I73739,I73722,I225603);
or I_4169 (I73756,I73739,I225606);
DFFARX1 I_4170 (I73756,I2859,I73315,I73782,);
nand I_4171 (I73790,I73782,I73448);
nor I_4172 (I73292,I73790,I73598);
nor I_4173 (I73286,I73782,I73414);
DFFARX1 I_4174 (I73782,I2859,I73315,I73844,);
not I_4175 (I73852,I73844);
nor I_4176 (I73301,I73852,I73564);
not I_4177 (I73910,I2866);
DFFARX1 I_4178 (I6259,I2859,I73910,I73936,);
DFFARX1 I_4179 (I73936,I2859,I73910,I73953,);
not I_4180 (I73902,I73953);
not I_4181 (I73975,I73936);
DFFARX1 I_4182 (I6235,I2859,I73910,I74001,);
not I_4183 (I74009,I74001);
and I_4184 (I74026,I73975,I6250);
not I_4185 (I74043,I6238);
nand I_4186 (I74060,I74043,I6250);
not I_4187 (I74077,I6241);
nor I_4188 (I74094,I74077,I6253);
nand I_4189 (I74111,I74094,I6244);
nor I_4190 (I74128,I74111,I74060);
DFFARX1 I_4191 (I74128,I2859,I73910,I73878,);
not I_4192 (I74159,I74111);
not I_4193 (I74176,I6253);
nand I_4194 (I74193,I74176,I6250);
nor I_4195 (I74210,I6253,I6238);
nand I_4196 (I73890,I74026,I74210);
nand I_4197 (I73884,I73975,I6253);
nand I_4198 (I74255,I74077,I6247);
DFFARX1 I_4199 (I74255,I2859,I73910,I73899,);
DFFARX1 I_4200 (I74255,I2859,I73910,I73893,);
not I_4201 (I74300,I6247);
nor I_4202 (I74317,I74300,I6238);
and I_4203 (I74334,I74317,I6235);
or I_4204 (I74351,I74334,I6256);
DFFARX1 I_4205 (I74351,I2859,I73910,I74377,);
nand I_4206 (I74385,I74377,I74043);
nor I_4207 (I73887,I74385,I74193);
nor I_4208 (I73881,I74377,I74009);
DFFARX1 I_4209 (I74377,I2859,I73910,I74439,);
not I_4210 (I74447,I74439);
nor I_4211 (I73896,I74447,I74159);
not I_4212 (I74505,I2866);
DFFARX1 I_4213 (I240187,I2859,I74505,I74531,);
DFFARX1 I_4214 (I74531,I2859,I74505,I74548,);
not I_4215 (I74497,I74548);
not I_4216 (I74570,I74531);
DFFARX1 I_4217 (I240178,I2859,I74505,I74596,);
not I_4218 (I74604,I74596);
and I_4219 (I74621,I74570,I240196);
not I_4220 (I74638,I240193);
nand I_4221 (I74655,I74638,I240196);
not I_4222 (I74672,I240172);
nor I_4223 (I74689,I74672,I240175);
nand I_4224 (I74706,I74689,I240184);
nor I_4225 (I74723,I74706,I74655);
DFFARX1 I_4226 (I74723,I2859,I74505,I74473,);
not I_4227 (I74754,I74706);
not I_4228 (I74771,I240175);
nand I_4229 (I74788,I74771,I240196);
nor I_4230 (I74805,I240175,I240193);
nand I_4231 (I74485,I74621,I74805);
nand I_4232 (I74479,I74570,I240175);
nand I_4233 (I74850,I74672,I240190);
DFFARX1 I_4234 (I74850,I2859,I74505,I74494,);
DFFARX1 I_4235 (I74850,I2859,I74505,I74488,);
not I_4236 (I74895,I240190);
nor I_4237 (I74912,I74895,I240172);
and I_4238 (I74929,I74912,I240181);
or I_4239 (I74946,I74929,I240175);
DFFARX1 I_4240 (I74946,I2859,I74505,I74972,);
nand I_4241 (I74980,I74972,I74638);
nor I_4242 (I74482,I74980,I74788);
nor I_4243 (I74476,I74972,I74604);
DFFARX1 I_4244 (I74972,I2859,I74505,I75034,);
not I_4245 (I75042,I75034);
nor I_4246 (I74491,I75042,I74754);
not I_4247 (I75100,I2866);
DFFARX1 I_4248 (I430371,I2859,I75100,I75126,);
DFFARX1 I_4249 (I75126,I2859,I75100,I75143,);
not I_4250 (I75092,I75143);
not I_4251 (I75165,I75126);
DFFARX1 I_4252 (I430380,I2859,I75100,I75191,);
not I_4253 (I75199,I75191);
and I_4254 (I75216,I75165,I430374);
not I_4255 (I75233,I430368);
nand I_4256 (I75250,I75233,I430374);
not I_4257 (I75267,I430383);
nor I_4258 (I75284,I75267,I430371);
nand I_4259 (I75301,I75284,I430377);
nor I_4260 (I75318,I75301,I75250);
DFFARX1 I_4261 (I75318,I2859,I75100,I75068,);
not I_4262 (I75349,I75301);
not I_4263 (I75366,I430371);
nand I_4264 (I75383,I75366,I430374);
nor I_4265 (I75400,I430371,I430368);
nand I_4266 (I75080,I75216,I75400);
nand I_4267 (I75074,I75165,I430371);
nand I_4268 (I75445,I75267,I430374);
DFFARX1 I_4269 (I75445,I2859,I75100,I75089,);
DFFARX1 I_4270 (I75445,I2859,I75100,I75083,);
not I_4271 (I75490,I430374);
nor I_4272 (I75507,I75490,I430389);
and I_4273 (I75524,I75507,I430386);
or I_4274 (I75541,I75524,I430368);
DFFARX1 I_4275 (I75541,I2859,I75100,I75567,);
nand I_4276 (I75575,I75567,I75233);
nor I_4277 (I75077,I75575,I75383);
nor I_4278 (I75071,I75567,I75199);
DFFARX1 I_4279 (I75567,I2859,I75100,I75629,);
not I_4280 (I75637,I75629);
nor I_4281 (I75086,I75637,I75349);
not I_4282 (I75695,I2866);
DFFARX1 I_4283 (I145601,I2859,I75695,I75721,);
DFFARX1 I_4284 (I75721,I2859,I75695,I75738,);
not I_4285 (I75687,I75738);
not I_4286 (I75760,I75721);
DFFARX1 I_4287 (I145616,I2859,I75695,I75786,);
not I_4288 (I75794,I75786);
and I_4289 (I75811,I75760,I145613);
not I_4290 (I75828,I145601);
nand I_4291 (I75845,I75828,I145613);
not I_4292 (I75862,I145610);
nor I_4293 (I75879,I75862,I145625);
nand I_4294 (I75896,I75879,I145622);
nor I_4295 (I75913,I75896,I75845);
DFFARX1 I_4296 (I75913,I2859,I75695,I75663,);
not I_4297 (I75944,I75896);
not I_4298 (I75961,I145625);
nand I_4299 (I75978,I75961,I145613);
nor I_4300 (I75995,I145625,I145601);
nand I_4301 (I75675,I75811,I75995);
nand I_4302 (I75669,I75760,I145625);
nand I_4303 (I76040,I75862,I145619);
DFFARX1 I_4304 (I76040,I2859,I75695,I75684,);
DFFARX1 I_4305 (I76040,I2859,I75695,I75678,);
not I_4306 (I76085,I145619);
nor I_4307 (I76102,I76085,I145607);
and I_4308 (I76119,I76102,I145628);
or I_4309 (I76136,I76119,I145604);
DFFARX1 I_4310 (I76136,I2859,I75695,I76162,);
nand I_4311 (I76170,I76162,I75828);
nor I_4312 (I75672,I76170,I75978);
nor I_4313 (I75666,I76162,I75794);
DFFARX1 I_4314 (I76162,I2859,I75695,I76224,);
not I_4315 (I76232,I76224);
nor I_4316 (I75681,I76232,I75944);
not I_4317 (I76290,I2866);
DFFARX1 I_4318 (I190131,I2859,I76290,I76316,);
DFFARX1 I_4319 (I76316,I2859,I76290,I76333,);
not I_4320 (I76282,I76333);
not I_4321 (I76355,I76316);
DFFARX1 I_4322 (I190119,I2859,I76290,I76381,);
not I_4323 (I76389,I76381);
and I_4324 (I76406,I76355,I190128);
not I_4325 (I76423,I190125);
nand I_4326 (I76440,I76423,I190128);
not I_4327 (I76457,I190116);
nor I_4328 (I76474,I76457,I190122);
nand I_4329 (I76491,I76474,I190107);
nor I_4330 (I76508,I76491,I76440);
DFFARX1 I_4331 (I76508,I2859,I76290,I76258,);
not I_4332 (I76539,I76491);
not I_4333 (I76556,I190122);
nand I_4334 (I76573,I76556,I190128);
nor I_4335 (I76590,I190122,I190125);
nand I_4336 (I76270,I76406,I76590);
nand I_4337 (I76264,I76355,I190122);
nand I_4338 (I76635,I76457,I190107);
DFFARX1 I_4339 (I76635,I2859,I76290,I76279,);
DFFARX1 I_4340 (I76635,I2859,I76290,I76273,);
not I_4341 (I76680,I190107);
nor I_4342 (I76697,I76680,I190113);
and I_4343 (I76714,I76697,I190110);
or I_4344 (I76731,I76714,I190134);
DFFARX1 I_4345 (I76731,I2859,I76290,I76757,);
nand I_4346 (I76765,I76757,I76423);
nor I_4347 (I76267,I76765,I76573);
nor I_4348 (I76261,I76757,I76389);
DFFARX1 I_4349 (I76757,I2859,I76290,I76819,);
not I_4350 (I76827,I76819);
nor I_4351 (I76276,I76827,I76539);
not I_4352 (I76885,I2866);
DFFARX1 I_4353 (I54728,I2859,I76885,I76911,);
DFFARX1 I_4354 (I76911,I2859,I76885,I76928,);
not I_4355 (I76877,I76928);
not I_4356 (I76950,I76911);
DFFARX1 I_4357 (I54722,I2859,I76885,I76976,);
not I_4358 (I76984,I76976);
and I_4359 (I77001,I76950,I54719);
not I_4360 (I77018,I54740);
nand I_4361 (I77035,I77018,I54719);
not I_4362 (I77052,I54734);
nor I_4363 (I77069,I77052,I54725);
nand I_4364 (I77086,I77069,I54731);
nor I_4365 (I77103,I77086,I77035);
DFFARX1 I_4366 (I77103,I2859,I76885,I76853,);
not I_4367 (I77134,I77086);
not I_4368 (I77151,I54725);
nand I_4369 (I77168,I77151,I54719);
nor I_4370 (I77185,I54725,I54740);
nand I_4371 (I76865,I77001,I77185);
nand I_4372 (I76859,I76950,I54725);
nand I_4373 (I77230,I77052,I54719);
DFFARX1 I_4374 (I77230,I2859,I76885,I76874,);
DFFARX1 I_4375 (I77230,I2859,I76885,I76868,);
not I_4376 (I77275,I54719);
nor I_4377 (I77292,I77275,I54737);
and I_4378 (I77309,I77292,I54743);
or I_4379 (I77326,I77309,I54722);
DFFARX1 I_4380 (I77326,I2859,I76885,I77352,);
nand I_4381 (I77360,I77352,I77018);
nor I_4382 (I76862,I77360,I77168);
nor I_4383 (I76856,I77352,I76984);
DFFARX1 I_4384 (I77352,I2859,I76885,I77414,);
not I_4385 (I77422,I77414);
nor I_4386 (I76871,I77422,I77134);
not I_4387 (I77480,I2866);
DFFARX1 I_4388 (I302608,I2859,I77480,I77506,);
DFFARX1 I_4389 (I77506,I2859,I77480,I77523,);
not I_4390 (I77472,I77523);
not I_4391 (I77545,I77506);
DFFARX1 I_4392 (I302605,I2859,I77480,I77571,);
not I_4393 (I77579,I77571);
and I_4394 (I77596,I77545,I302611);
not I_4395 (I77613,I302596);
nand I_4396 (I77630,I77613,I302611);
not I_4397 (I77647,I302599);
nor I_4398 (I77664,I77647,I302620);
nand I_4399 (I77681,I77664,I302617);
nor I_4400 (I77698,I77681,I77630);
DFFARX1 I_4401 (I77698,I2859,I77480,I77448,);
not I_4402 (I77729,I77681);
not I_4403 (I77746,I302620);
nand I_4404 (I77763,I77746,I302611);
nor I_4405 (I77780,I302620,I302596);
nand I_4406 (I77460,I77596,I77780);
nand I_4407 (I77454,I77545,I302620);
nand I_4408 (I77825,I77647,I302596);
DFFARX1 I_4409 (I77825,I2859,I77480,I77469,);
DFFARX1 I_4410 (I77825,I2859,I77480,I77463,);
not I_4411 (I77870,I302596);
nor I_4412 (I77887,I77870,I302602);
and I_4413 (I77904,I77887,I302614);
or I_4414 (I77921,I77904,I302599);
DFFARX1 I_4415 (I77921,I2859,I77480,I77947,);
nand I_4416 (I77955,I77947,I77613);
nor I_4417 (I77457,I77955,I77763);
nor I_4418 (I77451,I77947,I77579);
DFFARX1 I_4419 (I77947,I2859,I77480,I78009,);
not I_4420 (I78017,I78009);
nor I_4421 (I77466,I78017,I77729);
not I_4422 (I78075,I2866);
DFFARX1 I_4423 (I146128,I2859,I78075,I78101,);
DFFARX1 I_4424 (I78101,I2859,I78075,I78118,);
not I_4425 (I78067,I78118);
not I_4426 (I78140,I78101);
DFFARX1 I_4427 (I146143,I2859,I78075,I78166,);
not I_4428 (I78174,I78166);
and I_4429 (I78191,I78140,I146140);
not I_4430 (I78208,I146128);
nand I_4431 (I78225,I78208,I146140);
not I_4432 (I78242,I146137);
nor I_4433 (I78259,I78242,I146152);
nand I_4434 (I78276,I78259,I146149);
nor I_4435 (I78293,I78276,I78225);
DFFARX1 I_4436 (I78293,I2859,I78075,I78043,);
not I_4437 (I78324,I78276);
not I_4438 (I78341,I146152);
nand I_4439 (I78358,I78341,I146140);
nor I_4440 (I78375,I146152,I146128);
nand I_4441 (I78055,I78191,I78375);
nand I_4442 (I78049,I78140,I146152);
nand I_4443 (I78420,I78242,I146146);
DFFARX1 I_4444 (I78420,I2859,I78075,I78064,);
DFFARX1 I_4445 (I78420,I2859,I78075,I78058,);
not I_4446 (I78465,I146146);
nor I_4447 (I78482,I78465,I146134);
and I_4448 (I78499,I78482,I146155);
or I_4449 (I78516,I78499,I146131);
DFFARX1 I_4450 (I78516,I2859,I78075,I78542,);
nand I_4451 (I78550,I78542,I78208);
nor I_4452 (I78052,I78550,I78358);
nor I_4453 (I78046,I78542,I78174);
DFFARX1 I_4454 (I78542,I2859,I78075,I78604,);
not I_4455 (I78612,I78604);
nor I_4456 (I78061,I78612,I78324);
not I_4457 (I78670,I2866);
DFFARX1 I_4458 (I505900,I2859,I78670,I78696,);
DFFARX1 I_4459 (I78696,I2859,I78670,I78713,);
not I_4460 (I78662,I78713);
not I_4461 (I78735,I78696);
DFFARX1 I_4462 (I505885,I2859,I78670,I78761,);
not I_4463 (I78769,I78761);
and I_4464 (I78786,I78735,I505903);
not I_4465 (I78803,I505885);
nand I_4466 (I78820,I78803,I505903);
not I_4467 (I78837,I505906);
nor I_4468 (I78854,I78837,I505897);
nand I_4469 (I78871,I78854,I505894);
nor I_4470 (I78888,I78871,I78820);
DFFARX1 I_4471 (I78888,I2859,I78670,I78638,);
not I_4472 (I78919,I78871);
not I_4473 (I78936,I505897);
nand I_4474 (I78953,I78936,I505903);
nor I_4475 (I78970,I505897,I505885);
nand I_4476 (I78650,I78786,I78970);
nand I_4477 (I78644,I78735,I505897);
nand I_4478 (I79015,I78837,I505891);
DFFARX1 I_4479 (I79015,I2859,I78670,I78659,);
DFFARX1 I_4480 (I79015,I2859,I78670,I78653,);
not I_4481 (I79060,I505891);
nor I_4482 (I79077,I79060,I505882);
and I_4483 (I79094,I79077,I505888);
or I_4484 (I79111,I79094,I505882);
DFFARX1 I_4485 (I79111,I2859,I78670,I79137,);
nand I_4486 (I79145,I79137,I78803);
nor I_4487 (I78647,I79145,I78953);
nor I_4488 (I78641,I79137,I78769);
DFFARX1 I_4489 (I79137,I2859,I78670,I79199,);
not I_4490 (I79207,I79199);
nor I_4491 (I78656,I79207,I78919);
not I_4492 (I79265,I2866);
DFFARX1 I_4493 (I500340,I2859,I79265,I79291,);
DFFARX1 I_4494 (I79291,I2859,I79265,I79308,);
not I_4495 (I79257,I79308);
not I_4496 (I79330,I79291);
DFFARX1 I_4497 (I500340,I2859,I79265,I79356,);
not I_4498 (I79364,I79356);
and I_4499 (I79381,I79330,I500343);
not I_4500 (I79398,I500355);
nand I_4501 (I79415,I79398,I500343);
not I_4502 (I79432,I500361);
nor I_4503 (I79449,I79432,I500352);
nand I_4504 (I79466,I79449,I500358);
nor I_4505 (I79483,I79466,I79415);
DFFARX1 I_4506 (I79483,I2859,I79265,I79233,);
not I_4507 (I79514,I79466);
not I_4508 (I79531,I500352);
nand I_4509 (I79548,I79531,I500343);
nor I_4510 (I79565,I500352,I500355);
nand I_4511 (I79245,I79381,I79565);
nand I_4512 (I79239,I79330,I500352);
nand I_4513 (I79610,I79432,I500349);
DFFARX1 I_4514 (I79610,I2859,I79265,I79254,);
DFFARX1 I_4515 (I79610,I2859,I79265,I79248,);
not I_4516 (I79655,I500349);
nor I_4517 (I79672,I79655,I500346);
and I_4518 (I79689,I79672,I500364);
or I_4519 (I79706,I79689,I500343);
DFFARX1 I_4520 (I79706,I2859,I79265,I79732,);
nand I_4521 (I79740,I79732,I79398);
nor I_4522 (I79242,I79740,I79548);
nor I_4523 (I79236,I79732,I79364);
DFFARX1 I_4524 (I79732,I2859,I79265,I79794,);
not I_4525 (I79802,I79794);
nor I_4526 (I79251,I79802,I79514);
not I_4527 (I79860,I2866);
DFFARX1 I_4528 (I562751,I2859,I79860,I79886,);
DFFARX1 I_4529 (I79886,I2859,I79860,I79903,);
not I_4530 (I79852,I79903);
not I_4531 (I79925,I79886);
DFFARX1 I_4532 (I562742,I2859,I79860,I79951,);
not I_4533 (I79959,I79951);
and I_4534 (I79976,I79925,I562736);
not I_4535 (I79993,I562730);
nand I_4536 (I80010,I79993,I562736);
not I_4537 (I80027,I562757);
nor I_4538 (I80044,I80027,I562730);
nand I_4539 (I80061,I80044,I562754);
nor I_4540 (I80078,I80061,I80010);
DFFARX1 I_4541 (I80078,I2859,I79860,I79828,);
not I_4542 (I80109,I80061);
not I_4543 (I80126,I562730);
nand I_4544 (I80143,I80126,I562736);
nor I_4545 (I80160,I562730,I562730);
nand I_4546 (I79840,I79976,I80160);
nand I_4547 (I79834,I79925,I562730);
nand I_4548 (I80205,I80027,I562739);
DFFARX1 I_4549 (I80205,I2859,I79860,I79849,);
DFFARX1 I_4550 (I80205,I2859,I79860,I79843,);
not I_4551 (I80250,I562739);
nor I_4552 (I80267,I80250,I562745);
and I_4553 (I80284,I80267,I562748);
or I_4554 (I80301,I80284,I562733);
DFFARX1 I_4555 (I80301,I2859,I79860,I80327,);
nand I_4556 (I80335,I80327,I79993);
nor I_4557 (I79837,I80335,I80143);
nor I_4558 (I79831,I80327,I79959);
DFFARX1 I_4559 (I80327,I2859,I79860,I80389,);
not I_4560 (I80397,I80389);
nor I_4561 (I79846,I80397,I80109);
not I_4562 (I80455,I2866);
DFFARX1 I_4563 (I434859,I2859,I80455,I80481,);
DFFARX1 I_4564 (I80481,I2859,I80455,I80498,);
not I_4565 (I80447,I80498);
not I_4566 (I80520,I80481);
DFFARX1 I_4567 (I434868,I2859,I80455,I80546,);
not I_4568 (I80554,I80546);
and I_4569 (I80571,I80520,I434862);
not I_4570 (I80588,I434856);
nand I_4571 (I80605,I80588,I434862);
not I_4572 (I80622,I434871);
nor I_4573 (I80639,I80622,I434859);
nand I_4574 (I80656,I80639,I434865);
nor I_4575 (I80673,I80656,I80605);
DFFARX1 I_4576 (I80673,I2859,I80455,I80423,);
not I_4577 (I80704,I80656);
not I_4578 (I80721,I434859);
nand I_4579 (I80738,I80721,I434862);
nor I_4580 (I80755,I434859,I434856);
nand I_4581 (I80435,I80571,I80755);
nand I_4582 (I80429,I80520,I434859);
nand I_4583 (I80800,I80622,I434862);
DFFARX1 I_4584 (I80800,I2859,I80455,I80444,);
DFFARX1 I_4585 (I80800,I2859,I80455,I80438,);
not I_4586 (I80845,I434862);
nor I_4587 (I80862,I80845,I434877);
and I_4588 (I80879,I80862,I434874);
or I_4589 (I80896,I80879,I434856);
DFFARX1 I_4590 (I80896,I2859,I80455,I80922,);
nand I_4591 (I80930,I80922,I80588);
nor I_4592 (I80432,I80930,I80738);
nor I_4593 (I80426,I80922,I80554);
DFFARX1 I_4594 (I80922,I2859,I80455,I80984,);
not I_4595 (I80992,I80984);
nor I_4596 (I80441,I80992,I80704);
not I_4597 (I81050,I2866);
DFFARX1 I_4598 (I157195,I2859,I81050,I81076,);
DFFARX1 I_4599 (I81076,I2859,I81050,I81093,);
not I_4600 (I81042,I81093);
not I_4601 (I81115,I81076);
DFFARX1 I_4602 (I157210,I2859,I81050,I81141,);
not I_4603 (I81149,I81141);
and I_4604 (I81166,I81115,I157207);
not I_4605 (I81183,I157195);
nand I_4606 (I81200,I81183,I157207);
not I_4607 (I81217,I157204);
nor I_4608 (I81234,I81217,I157219);
nand I_4609 (I81251,I81234,I157216);
nor I_4610 (I81268,I81251,I81200);
DFFARX1 I_4611 (I81268,I2859,I81050,I81018,);
not I_4612 (I81299,I81251);
not I_4613 (I81316,I157219);
nand I_4614 (I81333,I81316,I157207);
nor I_4615 (I81350,I157219,I157195);
nand I_4616 (I81030,I81166,I81350);
nand I_4617 (I81024,I81115,I157219);
nand I_4618 (I81395,I81217,I157213);
DFFARX1 I_4619 (I81395,I2859,I81050,I81039,);
DFFARX1 I_4620 (I81395,I2859,I81050,I81033,);
not I_4621 (I81440,I157213);
nor I_4622 (I81457,I81440,I157201);
and I_4623 (I81474,I81457,I157222);
or I_4624 (I81491,I81474,I157198);
DFFARX1 I_4625 (I81491,I2859,I81050,I81517,);
nand I_4626 (I81525,I81517,I81183);
nor I_4627 (I81027,I81525,I81333);
nor I_4628 (I81021,I81517,I81149);
DFFARX1 I_4629 (I81517,I2859,I81050,I81579,);
not I_4630 (I81587,I81579);
nor I_4631 (I81036,I81587,I81299);
not I_4632 (I81645,I2866);
DFFARX1 I_4633 (I352157,I2859,I81645,I81671,);
DFFARX1 I_4634 (I81671,I2859,I81645,I81688,);
not I_4635 (I81637,I81688);
not I_4636 (I81710,I81671);
DFFARX1 I_4637 (I352151,I2859,I81645,I81736,);
not I_4638 (I81744,I81736);
and I_4639 (I81761,I81710,I352169);
not I_4640 (I81778,I352157);
nand I_4641 (I81795,I81778,I352169);
not I_4642 (I81812,I352151);
nor I_4643 (I81829,I81812,I352163);
nand I_4644 (I81846,I81829,I352154);
nor I_4645 (I81863,I81846,I81795);
DFFARX1 I_4646 (I81863,I2859,I81645,I81613,);
not I_4647 (I81894,I81846);
not I_4648 (I81911,I352163);
nand I_4649 (I81928,I81911,I352169);
nor I_4650 (I81945,I352163,I352157);
nand I_4651 (I81625,I81761,I81945);
nand I_4652 (I81619,I81710,I352163);
nand I_4653 (I81990,I81812,I352166);
DFFARX1 I_4654 (I81990,I2859,I81645,I81634,);
DFFARX1 I_4655 (I81990,I2859,I81645,I81628,);
not I_4656 (I82035,I352166);
nor I_4657 (I82052,I82035,I352172);
and I_4658 (I82069,I82052,I352154);
or I_4659 (I82086,I82069,I352160);
DFFARX1 I_4660 (I82086,I2859,I81645,I82112,);
nand I_4661 (I82120,I82112,I81778);
nor I_4662 (I81622,I82120,I81928);
nor I_4663 (I81616,I82112,I81744);
DFFARX1 I_4664 (I82112,I2859,I81645,I82174,);
not I_4665 (I82182,I82174);
nor I_4666 (I81631,I82182,I81894);
not I_4667 (I82240,I2866);
DFFARX1 I_4668 (I161411,I2859,I82240,I82266,);
DFFARX1 I_4669 (I82266,I2859,I82240,I82283,);
not I_4670 (I82232,I82283);
not I_4671 (I82305,I82266);
DFFARX1 I_4672 (I161426,I2859,I82240,I82331,);
not I_4673 (I82339,I82331);
and I_4674 (I82356,I82305,I161423);
not I_4675 (I82373,I161411);
nand I_4676 (I82390,I82373,I161423);
not I_4677 (I82407,I161420);
nor I_4678 (I82424,I82407,I161435);
nand I_4679 (I82441,I82424,I161432);
nor I_4680 (I82458,I82441,I82390);
DFFARX1 I_4681 (I82458,I2859,I82240,I82208,);
not I_4682 (I82489,I82441);
not I_4683 (I82506,I161435);
nand I_4684 (I82523,I82506,I161423);
nor I_4685 (I82540,I161435,I161411);
nand I_4686 (I82220,I82356,I82540);
nand I_4687 (I82214,I82305,I161435);
nand I_4688 (I82585,I82407,I161429);
DFFARX1 I_4689 (I82585,I2859,I82240,I82229,);
DFFARX1 I_4690 (I82585,I2859,I82240,I82223,);
not I_4691 (I82630,I161429);
nor I_4692 (I82647,I82630,I161417);
and I_4693 (I82664,I82647,I161438);
or I_4694 (I82681,I82664,I161414);
DFFARX1 I_4695 (I82681,I2859,I82240,I82707,);
nand I_4696 (I82715,I82707,I82373);
nor I_4697 (I82217,I82715,I82523);
nor I_4698 (I82211,I82707,I82339);
DFFARX1 I_4699 (I82707,I2859,I82240,I82769,);
not I_4700 (I82777,I82769);
nor I_4701 (I82226,I82777,I82489);
not I_4702 (I82835,I2866);
DFFARX1 I_4703 (I440469,I2859,I82835,I82861,);
DFFARX1 I_4704 (I82861,I2859,I82835,I82878,);
not I_4705 (I82827,I82878);
not I_4706 (I82900,I82861);
DFFARX1 I_4707 (I440478,I2859,I82835,I82926,);
not I_4708 (I82934,I82926);
and I_4709 (I82951,I82900,I440472);
not I_4710 (I82968,I440466);
nand I_4711 (I82985,I82968,I440472);
not I_4712 (I83002,I440481);
nor I_4713 (I83019,I83002,I440469);
nand I_4714 (I83036,I83019,I440475);
nor I_4715 (I83053,I83036,I82985);
DFFARX1 I_4716 (I83053,I2859,I82835,I82803,);
not I_4717 (I83084,I83036);
not I_4718 (I83101,I440469);
nand I_4719 (I83118,I83101,I440472);
nor I_4720 (I83135,I440469,I440466);
nand I_4721 (I82815,I82951,I83135);
nand I_4722 (I82809,I82900,I440469);
nand I_4723 (I83180,I83002,I440472);
DFFARX1 I_4724 (I83180,I2859,I82835,I82824,);
DFFARX1 I_4725 (I83180,I2859,I82835,I82818,);
not I_4726 (I83225,I440472);
nor I_4727 (I83242,I83225,I440487);
and I_4728 (I83259,I83242,I440484);
or I_4729 (I83276,I83259,I440466);
DFFARX1 I_4730 (I83276,I2859,I82835,I83302,);
nand I_4731 (I83310,I83302,I82968);
nor I_4732 (I82812,I83310,I83118);
nor I_4733 (I82806,I83302,I82934);
DFFARX1 I_4734 (I83302,I2859,I82835,I83364,);
not I_4735 (I83372,I83364);
nor I_4736 (I82821,I83372,I83084);
not I_4737 (I83430,I2866);
DFFARX1 I_4738 (I299140,I2859,I83430,I83456,);
DFFARX1 I_4739 (I83456,I2859,I83430,I83473,);
not I_4740 (I83422,I83473);
not I_4741 (I83495,I83456);
DFFARX1 I_4742 (I299137,I2859,I83430,I83521,);
not I_4743 (I83529,I83521);
and I_4744 (I83546,I83495,I299143);
not I_4745 (I83563,I299128);
nand I_4746 (I83580,I83563,I299143);
not I_4747 (I83597,I299131);
nor I_4748 (I83614,I83597,I299152);
nand I_4749 (I83631,I83614,I299149);
nor I_4750 (I83648,I83631,I83580);
DFFARX1 I_4751 (I83648,I2859,I83430,I83398,);
not I_4752 (I83679,I83631);
not I_4753 (I83696,I299152);
nand I_4754 (I83713,I83696,I299143);
nor I_4755 (I83730,I299152,I299128);
nand I_4756 (I83410,I83546,I83730);
nand I_4757 (I83404,I83495,I299152);
nand I_4758 (I83775,I83597,I299128);
DFFARX1 I_4759 (I83775,I2859,I83430,I83419,);
DFFARX1 I_4760 (I83775,I2859,I83430,I83413,);
not I_4761 (I83820,I299128);
nor I_4762 (I83837,I83820,I299134);
and I_4763 (I83854,I83837,I299146);
or I_4764 (I83871,I83854,I299131);
DFFARX1 I_4765 (I83871,I2859,I83430,I83897,);
nand I_4766 (I83905,I83897,I83563);
nor I_4767 (I83407,I83905,I83713);
nor I_4768 (I83401,I83897,I83529);
DFFARX1 I_4769 (I83897,I2859,I83430,I83959,);
not I_4770 (I83967,I83959);
nor I_4771 (I83416,I83967,I83679);
not I_4772 (I84025,I2866);
DFFARX1 I_4773 (I214905,I2859,I84025,I84051,);
DFFARX1 I_4774 (I84051,I2859,I84025,I84068,);
not I_4775 (I84017,I84068);
not I_4776 (I84090,I84051);
DFFARX1 I_4777 (I214899,I2859,I84025,I84116,);
not I_4778 (I84124,I84116);
and I_4779 (I84141,I84090,I214914);
not I_4780 (I84158,I214911);
nand I_4781 (I84175,I84158,I214914);
not I_4782 (I84192,I214902);
nor I_4783 (I84209,I84192,I214893);
nand I_4784 (I84226,I84209,I214896);
nor I_4785 (I84243,I84226,I84175);
DFFARX1 I_4786 (I84243,I2859,I84025,I83993,);
not I_4787 (I84274,I84226);
not I_4788 (I84291,I214893);
nand I_4789 (I84308,I84291,I214914);
nor I_4790 (I84325,I214893,I214911);
nand I_4791 (I84005,I84141,I84325);
nand I_4792 (I83999,I84090,I214893);
nand I_4793 (I84370,I84192,I214917);
DFFARX1 I_4794 (I84370,I2859,I84025,I84014,);
DFFARX1 I_4795 (I84370,I2859,I84025,I84008,);
not I_4796 (I84415,I214917);
nor I_4797 (I84432,I84415,I214908);
and I_4798 (I84449,I84432,I214893);
or I_4799 (I84466,I84449,I214896);
DFFARX1 I_4800 (I84466,I2859,I84025,I84492,);
nand I_4801 (I84500,I84492,I84158);
nor I_4802 (I84002,I84500,I84308);
nor I_4803 (I83996,I84492,I84124);
DFFARX1 I_4804 (I84492,I2859,I84025,I84554,);
not I_4805 (I84562,I84554);
nor I_4806 (I84011,I84562,I84274);
not I_4807 (I84620,I2866);
DFFARX1 I_4808 (I118197,I2859,I84620,I84646,);
DFFARX1 I_4809 (I84646,I2859,I84620,I84663,);
not I_4810 (I84612,I84663);
not I_4811 (I84685,I84646);
DFFARX1 I_4812 (I118212,I2859,I84620,I84711,);
not I_4813 (I84719,I84711);
and I_4814 (I84736,I84685,I118209);
not I_4815 (I84753,I118197);
nand I_4816 (I84770,I84753,I118209);
not I_4817 (I84787,I118206);
nor I_4818 (I84804,I84787,I118221);
nand I_4819 (I84821,I84804,I118218);
nor I_4820 (I84838,I84821,I84770);
DFFARX1 I_4821 (I84838,I2859,I84620,I84588,);
not I_4822 (I84869,I84821);
not I_4823 (I84886,I118221);
nand I_4824 (I84903,I84886,I118209);
nor I_4825 (I84920,I118221,I118197);
nand I_4826 (I84600,I84736,I84920);
nand I_4827 (I84594,I84685,I118221);
nand I_4828 (I84965,I84787,I118215);
DFFARX1 I_4829 (I84965,I2859,I84620,I84609,);
DFFARX1 I_4830 (I84965,I2859,I84620,I84603,);
not I_4831 (I85010,I118215);
nor I_4832 (I85027,I85010,I118203);
and I_4833 (I85044,I85027,I118224);
or I_4834 (I85061,I85044,I118200);
DFFARX1 I_4835 (I85061,I2859,I84620,I85087,);
nand I_4836 (I85095,I85087,I84753);
nor I_4837 (I84597,I85095,I84903);
nor I_4838 (I84591,I85087,I84719);
DFFARX1 I_4839 (I85087,I2859,I84620,I85149,);
not I_4840 (I85157,I85149);
nor I_4841 (I84606,I85157,I84869);
not I_4842 (I85215,I2866);
DFFARX1 I_4843 (I512428,I2859,I85215,I85241,);
DFFARX1 I_4844 (I85241,I2859,I85215,I85258,);
not I_4845 (I85207,I85258);
not I_4846 (I85280,I85241);
DFFARX1 I_4847 (I512413,I2859,I85215,I85306,);
not I_4848 (I85314,I85306);
and I_4849 (I85331,I85280,I512431);
not I_4850 (I85348,I512413);
nand I_4851 (I85365,I85348,I512431);
not I_4852 (I85382,I512434);
nor I_4853 (I85399,I85382,I512425);
nand I_4854 (I85416,I85399,I512422);
nor I_4855 (I85433,I85416,I85365);
DFFARX1 I_4856 (I85433,I2859,I85215,I85183,);
not I_4857 (I85464,I85416);
not I_4858 (I85481,I512425);
nand I_4859 (I85498,I85481,I512431);
nor I_4860 (I85515,I512425,I512413);
nand I_4861 (I85195,I85331,I85515);
nand I_4862 (I85189,I85280,I512425);
nand I_4863 (I85560,I85382,I512419);
DFFARX1 I_4864 (I85560,I2859,I85215,I85204,);
DFFARX1 I_4865 (I85560,I2859,I85215,I85198,);
not I_4866 (I85605,I512419);
nor I_4867 (I85622,I85605,I512410);
and I_4868 (I85639,I85622,I512416);
or I_4869 (I85656,I85639,I512410);
DFFARX1 I_4870 (I85656,I2859,I85215,I85682,);
nand I_4871 (I85690,I85682,I85348);
nor I_4872 (I85192,I85690,I85498);
nor I_4873 (I85186,I85682,I85314);
DFFARX1 I_4874 (I85682,I2859,I85215,I85744,);
not I_4875 (I85752,I85744);
nor I_4876 (I85201,I85752,I85464);
not I_4877 (I85810,I2866);
DFFARX1 I_4878 (I191763,I2859,I85810,I85836,);
DFFARX1 I_4879 (I85836,I2859,I85810,I85853,);
not I_4880 (I85802,I85853);
not I_4881 (I85875,I85836);
DFFARX1 I_4882 (I191751,I2859,I85810,I85901,);
not I_4883 (I85909,I85901);
and I_4884 (I85926,I85875,I191760);
not I_4885 (I85943,I191757);
nand I_4886 (I85960,I85943,I191760);
not I_4887 (I85977,I191748);
nor I_4888 (I85994,I85977,I191754);
nand I_4889 (I86011,I85994,I191739);
nor I_4890 (I86028,I86011,I85960);
DFFARX1 I_4891 (I86028,I2859,I85810,I85778,);
not I_4892 (I86059,I86011);
not I_4893 (I86076,I191754);
nand I_4894 (I86093,I86076,I191760);
nor I_4895 (I86110,I191754,I191757);
nand I_4896 (I85790,I85926,I86110);
nand I_4897 (I85784,I85875,I191754);
nand I_4898 (I86155,I85977,I191739);
DFFARX1 I_4899 (I86155,I2859,I85810,I85799,);
DFFARX1 I_4900 (I86155,I2859,I85810,I85793,);
not I_4901 (I86200,I191739);
nor I_4902 (I86217,I86200,I191745);
and I_4903 (I86234,I86217,I191742);
or I_4904 (I86251,I86234,I191766);
DFFARX1 I_4905 (I86251,I2859,I85810,I86277,);
nand I_4906 (I86285,I86277,I85943);
nor I_4907 (I85787,I86285,I86093);
nor I_4908 (I85781,I86277,I85909);
DFFARX1 I_4909 (I86277,I2859,I85810,I86339,);
not I_4910 (I86347,I86339);
nor I_4911 (I85796,I86347,I86059);
not I_4912 (I86405,I2866);
DFFARX1 I_4913 (I392558,I2859,I86405,I86431,);
DFFARX1 I_4914 (I86431,I2859,I86405,I86448,);
not I_4915 (I86397,I86448);
not I_4916 (I86470,I86431);
DFFARX1 I_4917 (I392567,I2859,I86405,I86496,);
not I_4918 (I86504,I86496);
and I_4919 (I86521,I86470,I392555);
not I_4920 (I86538,I392546);
nand I_4921 (I86555,I86538,I392555);
not I_4922 (I86572,I392552);
nor I_4923 (I86589,I86572,I392570);
nand I_4924 (I86606,I86589,I392543);
nor I_4925 (I86623,I86606,I86555);
DFFARX1 I_4926 (I86623,I2859,I86405,I86373,);
not I_4927 (I86654,I86606);
not I_4928 (I86671,I392570);
nand I_4929 (I86688,I86671,I392555);
nor I_4930 (I86705,I392570,I392546);
nand I_4931 (I86385,I86521,I86705);
nand I_4932 (I86379,I86470,I392570);
nand I_4933 (I86750,I86572,I392549);
DFFARX1 I_4934 (I86750,I2859,I86405,I86394,);
DFFARX1 I_4935 (I86750,I2859,I86405,I86388,);
not I_4936 (I86795,I392549);
nor I_4937 (I86812,I86795,I392561);
and I_4938 (I86829,I86812,I392543);
or I_4939 (I86846,I86829,I392564);
DFFARX1 I_4940 (I86846,I2859,I86405,I86872,);
nand I_4941 (I86880,I86872,I86538);
nor I_4942 (I86382,I86880,I86688);
nor I_4943 (I86376,I86872,I86504);
DFFARX1 I_4944 (I86872,I2859,I86405,I86934,);
not I_4945 (I86942,I86934);
nor I_4946 (I86391,I86942,I86654);
not I_4947 (I87000,I2866);
DFFARX1 I_4948 (I429249,I2859,I87000,I87026,);
DFFARX1 I_4949 (I87026,I2859,I87000,I87043,);
not I_4950 (I86992,I87043);
not I_4951 (I87065,I87026);
DFFARX1 I_4952 (I429258,I2859,I87000,I87091,);
not I_4953 (I87099,I87091);
and I_4954 (I87116,I87065,I429252);
not I_4955 (I87133,I429246);
nand I_4956 (I87150,I87133,I429252);
not I_4957 (I87167,I429261);
nor I_4958 (I87184,I87167,I429249);
nand I_4959 (I87201,I87184,I429255);
nor I_4960 (I87218,I87201,I87150);
DFFARX1 I_4961 (I87218,I2859,I87000,I86968,);
not I_4962 (I87249,I87201);
not I_4963 (I87266,I429249);
nand I_4964 (I87283,I87266,I429252);
nor I_4965 (I87300,I429249,I429246);
nand I_4966 (I86980,I87116,I87300);
nand I_4967 (I86974,I87065,I429249);
nand I_4968 (I87345,I87167,I429252);
DFFARX1 I_4969 (I87345,I2859,I87000,I86989,);
DFFARX1 I_4970 (I87345,I2859,I87000,I86983,);
not I_4971 (I87390,I429252);
nor I_4972 (I87407,I87390,I429267);
and I_4973 (I87424,I87407,I429264);
or I_4974 (I87441,I87424,I429246);
DFFARX1 I_4975 (I87441,I2859,I87000,I87467,);
nand I_4976 (I87475,I87467,I87133);
nor I_4977 (I86977,I87475,I87283);
nor I_4978 (I86971,I87467,I87099);
DFFARX1 I_4979 (I87467,I2859,I87000,I87529,);
not I_4980 (I87537,I87529);
nor I_4981 (I86986,I87537,I87249);
not I_4982 (I87595,I2866);
DFFARX1 I_4983 (I109765,I2859,I87595,I87621,);
DFFARX1 I_4984 (I87621,I2859,I87595,I87638,);
not I_4985 (I87587,I87638);
not I_4986 (I87660,I87621);
DFFARX1 I_4987 (I109780,I2859,I87595,I87686,);
not I_4988 (I87694,I87686);
and I_4989 (I87711,I87660,I109777);
not I_4990 (I87728,I109765);
nand I_4991 (I87745,I87728,I109777);
not I_4992 (I87762,I109774);
nor I_4993 (I87779,I87762,I109789);
nand I_4994 (I87796,I87779,I109786);
nor I_4995 (I87813,I87796,I87745);
DFFARX1 I_4996 (I87813,I2859,I87595,I87563,);
not I_4997 (I87844,I87796);
not I_4998 (I87861,I109789);
nand I_4999 (I87878,I87861,I109777);
nor I_5000 (I87895,I109789,I109765);
nand I_5001 (I87575,I87711,I87895);
nand I_5002 (I87569,I87660,I109789);
nand I_5003 (I87940,I87762,I109783);
DFFARX1 I_5004 (I87940,I2859,I87595,I87584,);
DFFARX1 I_5005 (I87940,I2859,I87595,I87578,);
not I_5006 (I87985,I109783);
nor I_5007 (I88002,I87985,I109771);
and I_5008 (I88019,I88002,I109792);
or I_5009 (I88036,I88019,I109768);
DFFARX1 I_5010 (I88036,I2859,I87595,I88062,);
nand I_5011 (I88070,I88062,I87728);
nor I_5012 (I87572,I88070,I87878);
nor I_5013 (I87566,I88062,I87694);
DFFARX1 I_5014 (I88062,I2859,I87595,I88124,);
not I_5015 (I88132,I88124);
nor I_5016 (I87581,I88132,I87844);
not I_5017 (I88190,I2866);
DFFARX1 I_5018 (I364805,I2859,I88190,I88216,);
DFFARX1 I_5019 (I88216,I2859,I88190,I88233,);
not I_5020 (I88182,I88233);
not I_5021 (I88255,I88216);
DFFARX1 I_5022 (I364799,I2859,I88190,I88281,);
not I_5023 (I88289,I88281);
and I_5024 (I88306,I88255,I364817);
not I_5025 (I88323,I364805);
nand I_5026 (I88340,I88323,I364817);
not I_5027 (I88357,I364799);
nor I_5028 (I88374,I88357,I364811);
nand I_5029 (I88391,I88374,I364802);
nor I_5030 (I88408,I88391,I88340);
DFFARX1 I_5031 (I88408,I2859,I88190,I88158,);
not I_5032 (I88439,I88391);
not I_5033 (I88456,I364811);
nand I_5034 (I88473,I88456,I364817);
nor I_5035 (I88490,I364811,I364805);
nand I_5036 (I88170,I88306,I88490);
nand I_5037 (I88164,I88255,I364811);
nand I_5038 (I88535,I88357,I364814);
DFFARX1 I_5039 (I88535,I2859,I88190,I88179,);
DFFARX1 I_5040 (I88535,I2859,I88190,I88173,);
not I_5041 (I88580,I364814);
nor I_5042 (I88597,I88580,I364820);
and I_5043 (I88614,I88597,I364802);
or I_5044 (I88631,I88614,I364808);
DFFARX1 I_5045 (I88631,I2859,I88190,I88657,);
nand I_5046 (I88665,I88657,I88323);
nor I_5047 (I88167,I88665,I88473);
nor I_5048 (I88161,I88657,I88289);
DFFARX1 I_5049 (I88657,I2859,I88190,I88719,);
not I_5050 (I88727,I88719);
nor I_5051 (I88176,I88727,I88439);
not I_5052 (I88785,I2866);
DFFARX1 I_5053 (I17326,I2859,I88785,I88811,);
DFFARX1 I_5054 (I88811,I2859,I88785,I88828,);
not I_5055 (I88777,I88828);
not I_5056 (I88850,I88811);
DFFARX1 I_5057 (I17302,I2859,I88785,I88876,);
not I_5058 (I88884,I88876);
and I_5059 (I88901,I88850,I17317);
not I_5060 (I88918,I17305);
nand I_5061 (I88935,I88918,I17317);
not I_5062 (I88952,I17308);
nor I_5063 (I88969,I88952,I17320);
nand I_5064 (I88986,I88969,I17311);
nor I_5065 (I89003,I88986,I88935);
DFFARX1 I_5066 (I89003,I2859,I88785,I88753,);
not I_5067 (I89034,I88986);
not I_5068 (I89051,I17320);
nand I_5069 (I89068,I89051,I17317);
nor I_5070 (I89085,I17320,I17305);
nand I_5071 (I88765,I88901,I89085);
nand I_5072 (I88759,I88850,I17320);
nand I_5073 (I89130,I88952,I17314);
DFFARX1 I_5074 (I89130,I2859,I88785,I88774,);
DFFARX1 I_5075 (I89130,I2859,I88785,I88768,);
not I_5076 (I89175,I17314);
nor I_5077 (I89192,I89175,I17305);
and I_5078 (I89209,I89192,I17302);
or I_5079 (I89226,I89209,I17323);
DFFARX1 I_5080 (I89226,I2859,I88785,I89252,);
nand I_5081 (I89260,I89252,I88918);
nor I_5082 (I88762,I89260,I89068);
nor I_5083 (I88756,I89252,I88884);
DFFARX1 I_5084 (I89252,I2859,I88785,I89314,);
not I_5085 (I89322,I89314);
nor I_5086 (I88771,I89322,I89034);
not I_5087 (I89380,I2866);
DFFARX1 I_5088 (I454678,I2859,I89380,I89406,);
DFFARX1 I_5089 (I89406,I2859,I89380,I89423,);
not I_5090 (I89372,I89423);
not I_5091 (I89445,I89406);
DFFARX1 I_5092 (I454678,I2859,I89380,I89471,);
not I_5093 (I89479,I89471);
and I_5094 (I89496,I89445,I454681);
not I_5095 (I89513,I454693);
nand I_5096 (I89530,I89513,I454681);
not I_5097 (I89547,I454699);
nor I_5098 (I89564,I89547,I454690);
nand I_5099 (I89581,I89564,I454696);
nor I_5100 (I89598,I89581,I89530);
DFFARX1 I_5101 (I89598,I2859,I89380,I89348,);
not I_5102 (I89629,I89581);
not I_5103 (I89646,I454690);
nand I_5104 (I89663,I89646,I454681);
nor I_5105 (I89680,I454690,I454693);
nand I_5106 (I89360,I89496,I89680);
nand I_5107 (I89354,I89445,I454690);
nand I_5108 (I89725,I89547,I454687);
DFFARX1 I_5109 (I89725,I2859,I89380,I89369,);
DFFARX1 I_5110 (I89725,I2859,I89380,I89363,);
not I_5111 (I89770,I454687);
nor I_5112 (I89787,I89770,I454684);
and I_5113 (I89804,I89787,I454702);
or I_5114 (I89821,I89804,I454681);
DFFARX1 I_5115 (I89821,I2859,I89380,I89847,);
nand I_5116 (I89855,I89847,I89513);
nor I_5117 (I89357,I89855,I89663);
nor I_5118 (I89351,I89847,I89479);
DFFARX1 I_5119 (I89847,I2859,I89380,I89909,);
not I_5120 (I89917,I89909);
nor I_5121 (I89366,I89917,I89629);
not I_5122 (I89975,I2866);
DFFARX1 I_5123 (I504812,I2859,I89975,I90001,);
DFFARX1 I_5124 (I90001,I2859,I89975,I90018,);
not I_5125 (I89967,I90018);
not I_5126 (I90040,I90001);
DFFARX1 I_5127 (I504797,I2859,I89975,I90066,);
not I_5128 (I90074,I90066);
and I_5129 (I90091,I90040,I504815);
not I_5130 (I90108,I504797);
nand I_5131 (I90125,I90108,I504815);
not I_5132 (I90142,I504818);
nor I_5133 (I90159,I90142,I504809);
nand I_5134 (I90176,I90159,I504806);
nor I_5135 (I90193,I90176,I90125);
DFFARX1 I_5136 (I90193,I2859,I89975,I89943,);
not I_5137 (I90224,I90176);
not I_5138 (I90241,I504809);
nand I_5139 (I90258,I90241,I504815);
nor I_5140 (I90275,I504809,I504797);
nand I_5141 (I89955,I90091,I90275);
nand I_5142 (I89949,I90040,I504809);
nand I_5143 (I90320,I90142,I504803);
DFFARX1 I_5144 (I90320,I2859,I89975,I89964,);
DFFARX1 I_5145 (I90320,I2859,I89975,I89958,);
not I_5146 (I90365,I504803);
nor I_5147 (I90382,I90365,I504794);
and I_5148 (I90399,I90382,I504800);
or I_5149 (I90416,I90399,I504794);
DFFARX1 I_5150 (I90416,I2859,I89975,I90442,);
nand I_5151 (I90450,I90442,I90108);
nor I_5152 (I89952,I90450,I90258);
nor I_5153 (I89946,I90442,I90074);
DFFARX1 I_5154 (I90442,I2859,I89975,I90504,);
not I_5155 (I90512,I90504);
nor I_5156 (I89961,I90512,I90224);
not I_5157 (I90570,I2866);
DFFARX1 I_5158 (I184691,I2859,I90570,I90596,);
DFFARX1 I_5159 (I90596,I2859,I90570,I90613,);
not I_5160 (I90562,I90613);
not I_5161 (I90635,I90596);
DFFARX1 I_5162 (I184679,I2859,I90570,I90661,);
not I_5163 (I90669,I90661);
and I_5164 (I90686,I90635,I184688);
not I_5165 (I90703,I184685);
nand I_5166 (I90720,I90703,I184688);
not I_5167 (I90737,I184676);
nor I_5168 (I90754,I90737,I184682);
nand I_5169 (I90771,I90754,I184667);
nor I_5170 (I90788,I90771,I90720);
DFFARX1 I_5171 (I90788,I2859,I90570,I90538,);
not I_5172 (I90819,I90771);
not I_5173 (I90836,I184682);
nand I_5174 (I90853,I90836,I184688);
nor I_5175 (I90870,I184682,I184685);
nand I_5176 (I90550,I90686,I90870);
nand I_5177 (I90544,I90635,I184682);
nand I_5178 (I90915,I90737,I184667);
DFFARX1 I_5179 (I90915,I2859,I90570,I90559,);
DFFARX1 I_5180 (I90915,I2859,I90570,I90553,);
not I_5181 (I90960,I184667);
nor I_5182 (I90977,I90960,I184673);
and I_5183 (I90994,I90977,I184670);
or I_5184 (I91011,I90994,I184694);
DFFARX1 I_5185 (I91011,I2859,I90570,I91037,);
nand I_5186 (I91045,I91037,I90703);
nor I_5187 (I90547,I91045,I90853);
nor I_5188 (I90541,I91037,I90669);
DFFARX1 I_5189 (I91037,I2859,I90570,I91099,);
not I_5190 (I91107,I91099);
nor I_5191 (I90556,I91107,I90819);
not I_5192 (I91165,I2866);
DFFARX1 I_5193 (I323416,I2859,I91165,I91191,);
DFFARX1 I_5194 (I91191,I2859,I91165,I91208,);
not I_5195 (I91157,I91208);
not I_5196 (I91230,I91191);
DFFARX1 I_5197 (I323413,I2859,I91165,I91256,);
not I_5198 (I91264,I91256);
and I_5199 (I91281,I91230,I323419);
not I_5200 (I91298,I323404);
nand I_5201 (I91315,I91298,I323419);
not I_5202 (I91332,I323407);
nor I_5203 (I91349,I91332,I323428);
nand I_5204 (I91366,I91349,I323425);
nor I_5205 (I91383,I91366,I91315);
DFFARX1 I_5206 (I91383,I2859,I91165,I91133,);
not I_5207 (I91414,I91366);
not I_5208 (I91431,I323428);
nand I_5209 (I91448,I91431,I323419);
nor I_5210 (I91465,I323428,I323404);
nand I_5211 (I91145,I91281,I91465);
nand I_5212 (I91139,I91230,I323428);
nand I_5213 (I91510,I91332,I323404);
DFFARX1 I_5214 (I91510,I2859,I91165,I91154,);
DFFARX1 I_5215 (I91510,I2859,I91165,I91148,);
not I_5216 (I91555,I323404);
nor I_5217 (I91572,I91555,I323410);
and I_5218 (I91589,I91572,I323422);
or I_5219 (I91606,I91589,I323407);
DFFARX1 I_5220 (I91606,I2859,I91165,I91632,);
nand I_5221 (I91640,I91632,I91298);
nor I_5222 (I91142,I91640,I91448);
nor I_5223 (I91136,I91632,I91264);
DFFARX1 I_5224 (I91632,I2859,I91165,I91694,);
not I_5225 (I91702,I91694);
nor I_5226 (I91151,I91702,I91414);
not I_5227 (I91760,I2866);
DFFARX1 I_5228 (I4077,I2859,I91760,I91786,);
DFFARX1 I_5229 (I91786,I2859,I91760,I91803,);
not I_5230 (I91752,I91803);
not I_5231 (I91825,I91786);
DFFARX1 I_5232 (I4074,I2859,I91760,I91851,);
not I_5233 (I91859,I91851);
and I_5234 (I91876,I91825,I4065);
not I_5235 (I91893,I4062);
nand I_5236 (I91910,I91893,I4065);
not I_5237 (I91927,I4062);
nor I_5238 (I91944,I91927,I4059);
nand I_5239 (I91961,I91944,I4071);
nor I_5240 (I91978,I91961,I91910);
DFFARX1 I_5241 (I91978,I2859,I91760,I91728,);
not I_5242 (I92009,I91961);
not I_5243 (I92026,I4059);
nand I_5244 (I92043,I92026,I4065);
nor I_5245 (I92060,I4059,I4062);
nand I_5246 (I91740,I91876,I92060);
nand I_5247 (I91734,I91825,I4059);
nand I_5248 (I92105,I91927,I4068);
DFFARX1 I_5249 (I92105,I2859,I91760,I91749,);
DFFARX1 I_5250 (I92105,I2859,I91760,I91743,);
not I_5251 (I92150,I4068);
nor I_5252 (I92167,I92150,I4080);
and I_5253 (I92184,I92167,I4065);
or I_5254 (I92201,I92184,I4059);
DFFARX1 I_5255 (I92201,I2859,I91760,I92227,);
nand I_5256 (I92235,I92227,I91893);
nor I_5257 (I91737,I92235,I92043);
nor I_5258 (I91731,I92227,I91859);
DFFARX1 I_5259 (I92227,I2859,I91760,I92289,);
not I_5260 (I92297,I92289);
nor I_5261 (I91746,I92297,I92009);
not I_5262 (I92355,I2866);
DFFARX1 I_5263 (I488780,I2859,I92355,I92381,);
DFFARX1 I_5264 (I92381,I2859,I92355,I92398,);
not I_5265 (I92347,I92398);
not I_5266 (I92420,I92381);
DFFARX1 I_5267 (I488780,I2859,I92355,I92446,);
not I_5268 (I92454,I92446);
and I_5269 (I92471,I92420,I488783);
not I_5270 (I92488,I488795);
nand I_5271 (I92505,I92488,I488783);
not I_5272 (I92522,I488801);
nor I_5273 (I92539,I92522,I488792);
nand I_5274 (I92556,I92539,I488798);
nor I_5275 (I92573,I92556,I92505);
DFFARX1 I_5276 (I92573,I2859,I92355,I92323,);
not I_5277 (I92604,I92556);
not I_5278 (I92621,I488792);
nand I_5279 (I92638,I92621,I488783);
nor I_5280 (I92655,I488792,I488795);
nand I_5281 (I92335,I92471,I92655);
nand I_5282 (I92329,I92420,I488792);
nand I_5283 (I92700,I92522,I488789);
DFFARX1 I_5284 (I92700,I2859,I92355,I92344,);
DFFARX1 I_5285 (I92700,I2859,I92355,I92338,);
not I_5286 (I92745,I488789);
nor I_5287 (I92762,I92745,I488786);
and I_5288 (I92779,I92762,I488804);
or I_5289 (I92796,I92779,I488783);
DFFARX1 I_5290 (I92796,I2859,I92355,I92822,);
nand I_5291 (I92830,I92822,I92488);
nor I_5292 (I92332,I92830,I92638);
nor I_5293 (I92326,I92822,I92454);
DFFARX1 I_5294 (I92822,I2859,I92355,I92884,);
not I_5295 (I92892,I92884);
nor I_5296 (I92341,I92892,I92604);
not I_5297 (I92950,I2866);
DFFARX1 I_5298 (I250591,I2859,I92950,I92976,);
DFFARX1 I_5299 (I92976,I2859,I92950,I92993,);
not I_5300 (I92942,I92993);
not I_5301 (I93015,I92976);
DFFARX1 I_5302 (I250582,I2859,I92950,I93041,);
not I_5303 (I93049,I93041);
and I_5304 (I93066,I93015,I250600);
not I_5305 (I93083,I250597);
nand I_5306 (I93100,I93083,I250600);
not I_5307 (I93117,I250576);
nor I_5308 (I93134,I93117,I250579);
nand I_5309 (I93151,I93134,I250588);
nor I_5310 (I93168,I93151,I93100);
DFFARX1 I_5311 (I93168,I2859,I92950,I92918,);
not I_5312 (I93199,I93151);
not I_5313 (I93216,I250579);
nand I_5314 (I93233,I93216,I250600);
nor I_5315 (I93250,I250579,I250597);
nand I_5316 (I92930,I93066,I93250);
nand I_5317 (I92924,I93015,I250579);
nand I_5318 (I93295,I93117,I250594);
DFFARX1 I_5319 (I93295,I2859,I92950,I92939,);
DFFARX1 I_5320 (I93295,I2859,I92950,I92933,);
not I_5321 (I93340,I250594);
nor I_5322 (I93357,I93340,I250576);
and I_5323 (I93374,I93357,I250585);
or I_5324 (I93391,I93374,I250579);
DFFARX1 I_5325 (I93391,I2859,I92950,I93417,);
nand I_5326 (I93425,I93417,I93083);
nor I_5327 (I92927,I93425,I93233);
nor I_5328 (I92921,I93417,I93049);
DFFARX1 I_5329 (I93417,I2859,I92950,I93479,);
not I_5330 (I93487,I93479);
nor I_5331 (I92936,I93487,I93199);
not I_5332 (I93545,I2866);
DFFARX1 I_5333 (I277754,I2859,I93545,I93571,);
DFFARX1 I_5334 (I93571,I2859,I93545,I93588,);
not I_5335 (I93537,I93588);
not I_5336 (I93610,I93571);
DFFARX1 I_5337 (I277751,I2859,I93545,I93636,);
not I_5338 (I93644,I93636);
and I_5339 (I93661,I93610,I277757);
not I_5340 (I93678,I277742);
nand I_5341 (I93695,I93678,I277757);
not I_5342 (I93712,I277745);
nor I_5343 (I93729,I93712,I277766);
nand I_5344 (I93746,I93729,I277763);
nor I_5345 (I93763,I93746,I93695);
DFFARX1 I_5346 (I93763,I2859,I93545,I93513,);
not I_5347 (I93794,I93746);
not I_5348 (I93811,I277766);
nand I_5349 (I93828,I93811,I277757);
nor I_5350 (I93845,I277766,I277742);
nand I_5351 (I93525,I93661,I93845);
nand I_5352 (I93519,I93610,I277766);
nand I_5353 (I93890,I93712,I277742);
DFFARX1 I_5354 (I93890,I2859,I93545,I93534,);
DFFARX1 I_5355 (I93890,I2859,I93545,I93528,);
not I_5356 (I93935,I277742);
nor I_5357 (I93952,I93935,I277748);
and I_5358 (I93969,I93952,I277760);
or I_5359 (I93986,I93969,I277745);
DFFARX1 I_5360 (I93986,I2859,I93545,I94012,);
nand I_5361 (I94020,I94012,I93678);
nor I_5362 (I93522,I94020,I93828);
nor I_5363 (I93516,I94012,I93644);
DFFARX1 I_5364 (I94012,I2859,I93545,I94074,);
not I_5365 (I94082,I94074);
nor I_5366 (I93531,I94082,I93794);
not I_5367 (I94140,I2866);
DFFARX1 I_5368 (I135061,I2859,I94140,I94166,);
DFFARX1 I_5369 (I94166,I2859,I94140,I94183,);
not I_5370 (I94132,I94183);
not I_5371 (I94205,I94166);
DFFARX1 I_5372 (I135076,I2859,I94140,I94231,);
not I_5373 (I94239,I94231);
and I_5374 (I94256,I94205,I135073);
not I_5375 (I94273,I135061);
nand I_5376 (I94290,I94273,I135073);
not I_5377 (I94307,I135070);
nor I_5378 (I94324,I94307,I135085);
nand I_5379 (I94341,I94324,I135082);
nor I_5380 (I94358,I94341,I94290);
DFFARX1 I_5381 (I94358,I2859,I94140,I94108,);
not I_5382 (I94389,I94341);
not I_5383 (I94406,I135085);
nand I_5384 (I94423,I94406,I135073);
nor I_5385 (I94440,I135085,I135061);
nand I_5386 (I94120,I94256,I94440);
nand I_5387 (I94114,I94205,I135085);
nand I_5388 (I94485,I94307,I135079);
DFFARX1 I_5389 (I94485,I2859,I94140,I94129,);
DFFARX1 I_5390 (I94485,I2859,I94140,I94123,);
not I_5391 (I94530,I135079);
nor I_5392 (I94547,I94530,I135067);
and I_5393 (I94564,I94547,I135088);
or I_5394 (I94581,I94564,I135064);
DFFARX1 I_5395 (I94581,I2859,I94140,I94607,);
nand I_5396 (I94615,I94607,I94273);
nor I_5397 (I94117,I94615,I94423);
nor I_5398 (I94111,I94607,I94239);
DFFARX1 I_5399 (I94607,I2859,I94140,I94669,);
not I_5400 (I94677,I94669);
nor I_5401 (I94126,I94677,I94389);
not I_5402 (I94735,I2866);
DFFARX1 I_5403 (I244811,I2859,I94735,I94761,);
DFFARX1 I_5404 (I94761,I2859,I94735,I94778,);
not I_5405 (I94727,I94778);
not I_5406 (I94800,I94761);
DFFARX1 I_5407 (I244802,I2859,I94735,I94826,);
not I_5408 (I94834,I94826);
and I_5409 (I94851,I94800,I244820);
not I_5410 (I94868,I244817);
nand I_5411 (I94885,I94868,I244820);
not I_5412 (I94902,I244796);
nor I_5413 (I94919,I94902,I244799);
nand I_5414 (I94936,I94919,I244808);
nor I_5415 (I94953,I94936,I94885);
DFFARX1 I_5416 (I94953,I2859,I94735,I94703,);
not I_5417 (I94984,I94936);
not I_5418 (I95001,I244799);
nand I_5419 (I95018,I95001,I244820);
nor I_5420 (I95035,I244799,I244817);
nand I_5421 (I94715,I94851,I95035);
nand I_5422 (I94709,I94800,I244799);
nand I_5423 (I95080,I94902,I244814);
DFFARX1 I_5424 (I95080,I2859,I94735,I94724,);
DFFARX1 I_5425 (I95080,I2859,I94735,I94718,);
not I_5426 (I95125,I244814);
nor I_5427 (I95142,I95125,I244796);
and I_5428 (I95159,I95142,I244805);
or I_5429 (I95176,I95159,I244799);
DFFARX1 I_5430 (I95176,I2859,I94735,I95202,);
nand I_5431 (I95210,I95202,I94868);
nor I_5432 (I94712,I95210,I95018);
nor I_5433 (I94706,I95202,I94834);
DFFARX1 I_5434 (I95202,I2859,I94735,I95264,);
not I_5435 (I95272,I95264);
nor I_5436 (I94721,I95272,I94984);
not I_5437 (I95330,I2866);
DFFARX1 I_5438 (I117670,I2859,I95330,I95356,);
DFFARX1 I_5439 (I95356,I2859,I95330,I95373,);
not I_5440 (I95322,I95373);
not I_5441 (I95395,I95356);
DFFARX1 I_5442 (I117685,I2859,I95330,I95421,);
not I_5443 (I95429,I95421);
and I_5444 (I95446,I95395,I117682);
not I_5445 (I95463,I117670);
nand I_5446 (I95480,I95463,I117682);
not I_5447 (I95497,I117679);
nor I_5448 (I95514,I95497,I117694);
nand I_5449 (I95531,I95514,I117691);
nor I_5450 (I95548,I95531,I95480);
DFFARX1 I_5451 (I95548,I2859,I95330,I95298,);
not I_5452 (I95579,I95531);
not I_5453 (I95596,I117694);
nand I_5454 (I95613,I95596,I117682);
nor I_5455 (I95630,I117694,I117670);
nand I_5456 (I95310,I95446,I95630);
nand I_5457 (I95304,I95395,I117694);
nand I_5458 (I95675,I95497,I117688);
DFFARX1 I_5459 (I95675,I2859,I95330,I95319,);
DFFARX1 I_5460 (I95675,I2859,I95330,I95313,);
not I_5461 (I95720,I117688);
nor I_5462 (I95737,I95720,I117676);
and I_5463 (I95754,I95737,I117697);
or I_5464 (I95771,I95754,I117673);
DFFARX1 I_5465 (I95771,I2859,I95330,I95797,);
nand I_5466 (I95805,I95797,I95463);
nor I_5467 (I95307,I95805,I95613);
nor I_5468 (I95301,I95797,I95429);
DFFARX1 I_5469 (I95797,I2859,I95330,I95859,);
not I_5470 (I95867,I95859);
nor I_5471 (I95316,I95867,I95579);
not I_5472 (I95925,I2866);
DFFARX1 I_5473 (I122940,I2859,I95925,I95951,);
DFFARX1 I_5474 (I95951,I2859,I95925,I95968,);
not I_5475 (I95917,I95968);
not I_5476 (I95990,I95951);
DFFARX1 I_5477 (I122955,I2859,I95925,I96016,);
not I_5478 (I96024,I96016);
and I_5479 (I96041,I95990,I122952);
not I_5480 (I96058,I122940);
nand I_5481 (I96075,I96058,I122952);
not I_5482 (I96092,I122949);
nor I_5483 (I96109,I96092,I122964);
nand I_5484 (I96126,I96109,I122961);
nor I_5485 (I96143,I96126,I96075);
DFFARX1 I_5486 (I96143,I2859,I95925,I95893,);
not I_5487 (I96174,I96126);
not I_5488 (I96191,I122964);
nand I_5489 (I96208,I96191,I122952);
nor I_5490 (I96225,I122964,I122940);
nand I_5491 (I95905,I96041,I96225);
nand I_5492 (I95899,I95990,I122964);
nand I_5493 (I96270,I96092,I122958);
DFFARX1 I_5494 (I96270,I2859,I95925,I95914,);
DFFARX1 I_5495 (I96270,I2859,I95925,I95908,);
not I_5496 (I96315,I122958);
nor I_5497 (I96332,I96315,I122946);
and I_5498 (I96349,I96332,I122967);
or I_5499 (I96366,I96349,I122943);
DFFARX1 I_5500 (I96366,I2859,I95925,I96392,);
nand I_5501 (I96400,I96392,I96058);
nor I_5502 (I95902,I96400,I96208);
nor I_5503 (I95896,I96392,I96024);
DFFARX1 I_5504 (I96392,I2859,I95925,I96454,);
not I_5505 (I96462,I96454);
nor I_5506 (I95911,I96462,I96174);
not I_5507 (I96520,I2866);
DFFARX1 I_5508 (I475486,I2859,I96520,I96546,);
DFFARX1 I_5509 (I96546,I2859,I96520,I96563,);
not I_5510 (I96512,I96563);
not I_5511 (I96585,I96546);
DFFARX1 I_5512 (I475486,I2859,I96520,I96611,);
not I_5513 (I96619,I96611);
and I_5514 (I96636,I96585,I475489);
not I_5515 (I96653,I475501);
nand I_5516 (I96670,I96653,I475489);
not I_5517 (I96687,I475507);
nor I_5518 (I96704,I96687,I475498);
nand I_5519 (I96721,I96704,I475504);
nor I_5520 (I96738,I96721,I96670);
DFFARX1 I_5521 (I96738,I2859,I96520,I96488,);
not I_5522 (I96769,I96721);
not I_5523 (I96786,I475498);
nand I_5524 (I96803,I96786,I475489);
nor I_5525 (I96820,I475498,I475501);
nand I_5526 (I96500,I96636,I96820);
nand I_5527 (I96494,I96585,I475498);
nand I_5528 (I96865,I96687,I475495);
DFFARX1 I_5529 (I96865,I2859,I96520,I96509,);
DFFARX1 I_5530 (I96865,I2859,I96520,I96503,);
not I_5531 (I96910,I475495);
nor I_5532 (I96927,I96910,I475492);
and I_5533 (I96944,I96927,I475510);
or I_5534 (I96961,I96944,I475489);
DFFARX1 I_5535 (I96961,I2859,I96520,I96987,);
nand I_5536 (I96995,I96987,I96653);
nor I_5537 (I96497,I96995,I96803);
nor I_5538 (I96491,I96987,I96619);
DFFARX1 I_5539 (I96987,I2859,I96520,I97049,);
not I_5540 (I97057,I97049);
nor I_5541 (I96506,I97057,I96769);
not I_5542 (I97115,I2866);
DFFARX1 I_5543 (I180883,I2859,I97115,I97141,);
DFFARX1 I_5544 (I97141,I2859,I97115,I97158,);
not I_5545 (I97107,I97158);
not I_5546 (I97180,I97141);
DFFARX1 I_5547 (I180871,I2859,I97115,I97206,);
not I_5548 (I97214,I97206);
and I_5549 (I97231,I97180,I180880);
not I_5550 (I97248,I180877);
nand I_5551 (I97265,I97248,I180880);
not I_5552 (I97282,I180868);
nor I_5553 (I97299,I97282,I180874);
nand I_5554 (I97316,I97299,I180859);
nor I_5555 (I97333,I97316,I97265);
DFFARX1 I_5556 (I97333,I2859,I97115,I97083,);
not I_5557 (I97364,I97316);
not I_5558 (I97381,I180874);
nand I_5559 (I97398,I97381,I180880);
nor I_5560 (I97415,I180874,I180877);
nand I_5561 (I97095,I97231,I97415);
nand I_5562 (I97089,I97180,I180874);
nand I_5563 (I97460,I97282,I180859);
DFFARX1 I_5564 (I97460,I2859,I97115,I97104,);
DFFARX1 I_5565 (I97460,I2859,I97115,I97098,);
not I_5566 (I97505,I180859);
nor I_5567 (I97522,I97505,I180865);
and I_5568 (I97539,I97522,I180862);
or I_5569 (I97556,I97539,I180886);
DFFARX1 I_5570 (I97556,I2859,I97115,I97582,);
nand I_5571 (I97590,I97582,I97248);
nor I_5572 (I97092,I97590,I97398);
nor I_5573 (I97086,I97582,I97214);
DFFARX1 I_5574 (I97582,I2859,I97115,I97644,);
not I_5575 (I97652,I97644);
nor I_5576 (I97101,I97652,I97364);
not I_5577 (I97710,I2866);
DFFARX1 I_5578 (I302030,I2859,I97710,I97736,);
DFFARX1 I_5579 (I97736,I2859,I97710,I97753,);
not I_5580 (I97702,I97753);
not I_5581 (I97775,I97736);
DFFARX1 I_5582 (I302027,I2859,I97710,I97801,);
not I_5583 (I97809,I97801);
and I_5584 (I97826,I97775,I302033);
not I_5585 (I97843,I302018);
nand I_5586 (I97860,I97843,I302033);
not I_5587 (I97877,I302021);
nor I_5588 (I97894,I97877,I302042);
nand I_5589 (I97911,I97894,I302039);
nor I_5590 (I97928,I97911,I97860);
DFFARX1 I_5591 (I97928,I2859,I97710,I97678,);
not I_5592 (I97959,I97911);
not I_5593 (I97976,I302042);
nand I_5594 (I97993,I97976,I302033);
nor I_5595 (I98010,I302042,I302018);
nand I_5596 (I97690,I97826,I98010);
nand I_5597 (I97684,I97775,I302042);
nand I_5598 (I98055,I97877,I302018);
DFFARX1 I_5599 (I98055,I2859,I97710,I97699,);
DFFARX1 I_5600 (I98055,I2859,I97710,I97693,);
not I_5601 (I98100,I302018);
nor I_5602 (I98117,I98100,I302024);
and I_5603 (I98134,I98117,I302036);
or I_5604 (I98151,I98134,I302021);
DFFARX1 I_5605 (I98151,I2859,I97710,I98177,);
nand I_5606 (I98185,I98177,I97843);
nor I_5607 (I97687,I98185,I97993);
nor I_5608 (I97681,I98177,I97809);
DFFARX1 I_5609 (I98177,I2859,I97710,I98239,);
not I_5610 (I98247,I98239);
nor I_5611 (I97696,I98247,I97959);
not I_5612 (I98305,I2866);
DFFARX1 I_5613 (I361643,I2859,I98305,I98331,);
DFFARX1 I_5614 (I98331,I2859,I98305,I98348,);
not I_5615 (I98297,I98348);
not I_5616 (I98370,I98331);
DFFARX1 I_5617 (I361637,I2859,I98305,I98396,);
not I_5618 (I98404,I98396);
and I_5619 (I98421,I98370,I361655);
not I_5620 (I98438,I361643);
nand I_5621 (I98455,I98438,I361655);
not I_5622 (I98472,I361637);
nor I_5623 (I98489,I98472,I361649);
nand I_5624 (I98506,I98489,I361640);
nor I_5625 (I98523,I98506,I98455);
DFFARX1 I_5626 (I98523,I2859,I98305,I98273,);
not I_5627 (I98554,I98506);
not I_5628 (I98571,I361649);
nand I_5629 (I98588,I98571,I361655);
nor I_5630 (I98605,I361649,I361643);
nand I_5631 (I98285,I98421,I98605);
nand I_5632 (I98279,I98370,I361649);
nand I_5633 (I98650,I98472,I361652);
DFFARX1 I_5634 (I98650,I2859,I98305,I98294,);
DFFARX1 I_5635 (I98650,I2859,I98305,I98288,);
not I_5636 (I98695,I361652);
nor I_5637 (I98712,I98695,I361658);
and I_5638 (I98729,I98712,I361640);
or I_5639 (I98746,I98729,I361646);
DFFARX1 I_5640 (I98746,I2859,I98305,I98772,);
nand I_5641 (I98780,I98772,I98438);
nor I_5642 (I98282,I98780,I98588);
nor I_5643 (I98276,I98772,I98404);
DFFARX1 I_5644 (I98772,I2859,I98305,I98834,);
not I_5645 (I98842,I98834);
nor I_5646 (I98291,I98842,I98554);
not I_5647 (I98900,I2866);
DFFARX1 I_5648 (I462192,I2859,I98900,I98926,);
DFFARX1 I_5649 (I98926,I2859,I98900,I98943,);
not I_5650 (I98892,I98943);
not I_5651 (I98965,I98926);
DFFARX1 I_5652 (I462192,I2859,I98900,I98991,);
not I_5653 (I98999,I98991);
and I_5654 (I99016,I98965,I462195);
not I_5655 (I99033,I462207);
nand I_5656 (I99050,I99033,I462195);
not I_5657 (I99067,I462213);
nor I_5658 (I99084,I99067,I462204);
nand I_5659 (I99101,I99084,I462210);
nor I_5660 (I99118,I99101,I99050);
DFFARX1 I_5661 (I99118,I2859,I98900,I98868,);
not I_5662 (I99149,I99101);
not I_5663 (I99166,I462204);
nand I_5664 (I99183,I99166,I462195);
nor I_5665 (I99200,I462204,I462207);
nand I_5666 (I98880,I99016,I99200);
nand I_5667 (I98874,I98965,I462204);
nand I_5668 (I99245,I99067,I462201);
DFFARX1 I_5669 (I99245,I2859,I98900,I98889,);
DFFARX1 I_5670 (I99245,I2859,I98900,I98883,);
not I_5671 (I99290,I462201);
nor I_5672 (I99307,I99290,I462198);
and I_5673 (I99324,I99307,I462216);
or I_5674 (I99341,I99324,I462195);
DFFARX1 I_5675 (I99341,I2859,I98900,I99367,);
nand I_5676 (I99375,I99367,I99033);
nor I_5677 (I98877,I99375,I99183);
nor I_5678 (I98871,I99367,I98999);
DFFARX1 I_5679 (I99367,I2859,I98900,I99429,);
not I_5680 (I99437,I99429);
nor I_5681 (I98886,I99437,I99149);
not I_5682 (I99495,I2866);
DFFARX1 I_5683 (I370075,I2859,I99495,I99521,);
DFFARX1 I_5684 (I99521,I2859,I99495,I99538,);
not I_5685 (I99487,I99538);
not I_5686 (I99560,I99521);
DFFARX1 I_5687 (I370069,I2859,I99495,I99586,);
not I_5688 (I99594,I99586);
and I_5689 (I99611,I99560,I370087);
not I_5690 (I99628,I370075);
nand I_5691 (I99645,I99628,I370087);
not I_5692 (I99662,I370069);
nor I_5693 (I99679,I99662,I370081);
nand I_5694 (I99696,I99679,I370072);
nor I_5695 (I99713,I99696,I99645);
DFFARX1 I_5696 (I99713,I2859,I99495,I99463,);
not I_5697 (I99744,I99696);
not I_5698 (I99761,I370081);
nand I_5699 (I99778,I99761,I370087);
nor I_5700 (I99795,I370081,I370075);
nand I_5701 (I99475,I99611,I99795);
nand I_5702 (I99469,I99560,I370081);
nand I_5703 (I99840,I99662,I370084);
DFFARX1 I_5704 (I99840,I2859,I99495,I99484,);
DFFARX1 I_5705 (I99840,I2859,I99495,I99478,);
not I_5706 (I99885,I370084);
nor I_5707 (I99902,I99885,I370090);
and I_5708 (I99919,I99902,I370072);
or I_5709 (I99936,I99919,I370078);
DFFARX1 I_5710 (I99936,I2859,I99495,I99962,);
nand I_5711 (I99970,I99962,I99628);
nor I_5712 (I99472,I99970,I99778);
nor I_5713 (I99466,I99962,I99594);
DFFARX1 I_5714 (I99962,I2859,I99495,I100024,);
not I_5715 (I100032,I100024);
nor I_5716 (I99481,I100032,I99744);
not I_5717 (I100090,I2866);
DFFARX1 I_5718 (I230939,I2859,I100090,I100116,);
DFFARX1 I_5719 (I100116,I2859,I100090,I100133,);
not I_5720 (I100082,I100133);
not I_5721 (I100155,I100116);
DFFARX1 I_5722 (I230930,I2859,I100090,I100181,);
not I_5723 (I100189,I100181);
and I_5724 (I100206,I100155,I230948);
not I_5725 (I100223,I230945);
nand I_5726 (I100240,I100223,I230948);
not I_5727 (I100257,I230924);
nor I_5728 (I100274,I100257,I230927);
nand I_5729 (I100291,I100274,I230936);
nor I_5730 (I100308,I100291,I100240);
DFFARX1 I_5731 (I100308,I2859,I100090,I100058,);
not I_5732 (I100339,I100291);
not I_5733 (I100356,I230927);
nand I_5734 (I100373,I100356,I230948);
nor I_5735 (I100390,I230927,I230945);
nand I_5736 (I100070,I100206,I100390);
nand I_5737 (I100064,I100155,I230927);
nand I_5738 (I100435,I100257,I230942);
DFFARX1 I_5739 (I100435,I2859,I100090,I100079,);
DFFARX1 I_5740 (I100435,I2859,I100090,I100073,);
not I_5741 (I100480,I230942);
nor I_5742 (I100497,I100480,I230924);
and I_5743 (I100514,I100497,I230933);
or I_5744 (I100531,I100514,I230927);
DFFARX1 I_5745 (I100531,I2859,I100090,I100557,);
nand I_5746 (I100565,I100557,I100223);
nor I_5747 (I100067,I100565,I100373);
nor I_5748 (I100061,I100557,I100189);
DFFARX1 I_5749 (I100557,I2859,I100090,I100619,);
not I_5750 (I100627,I100619);
nor I_5751 (I100076,I100627,I100339);
not I_5752 (I100685,I2866);
DFFARX1 I_5753 (I516780,I2859,I100685,I100711,);
DFFARX1 I_5754 (I100711,I2859,I100685,I100728,);
not I_5755 (I100677,I100728);
not I_5756 (I100750,I100711);
DFFARX1 I_5757 (I516765,I2859,I100685,I100776,);
not I_5758 (I100784,I100776);
and I_5759 (I100801,I100750,I516783);
not I_5760 (I100818,I516765);
nand I_5761 (I100835,I100818,I516783);
not I_5762 (I100852,I516786);
nor I_5763 (I100869,I100852,I516777);
nand I_5764 (I100886,I100869,I516774);
nor I_5765 (I100903,I100886,I100835);
DFFARX1 I_5766 (I100903,I2859,I100685,I100653,);
not I_5767 (I100934,I100886);
not I_5768 (I100951,I516777);
nand I_5769 (I100968,I100951,I516783);
nor I_5770 (I100985,I516777,I516765);
nand I_5771 (I100665,I100801,I100985);
nand I_5772 (I100659,I100750,I516777);
nand I_5773 (I101030,I100852,I516771);
DFFARX1 I_5774 (I101030,I2859,I100685,I100674,);
DFFARX1 I_5775 (I101030,I2859,I100685,I100668,);
not I_5776 (I101075,I516771);
nor I_5777 (I101092,I101075,I516762);
and I_5778 (I101109,I101092,I516768);
or I_5779 (I101126,I101109,I516762);
DFFARX1 I_5780 (I101126,I2859,I100685,I101152,);
nand I_5781 (I101160,I101152,I100818);
nor I_5782 (I100662,I101160,I100968);
nor I_5783 (I100656,I101152,I100784);
DFFARX1 I_5784 (I101152,I2859,I100685,I101214,);
not I_5785 (I101222,I101214);
nor I_5786 (I100671,I101222,I100934);
not I_5787 (I101280,I2866);
DFFARX1 I_5788 (I415814,I2859,I101280,I101306,);
DFFARX1 I_5789 (I101306,I2859,I101280,I101323,);
not I_5790 (I101272,I101323);
not I_5791 (I101345,I101306);
DFFARX1 I_5792 (I415823,I2859,I101280,I101371,);
not I_5793 (I101379,I101371);
and I_5794 (I101396,I101345,I415811);
not I_5795 (I101413,I415802);
nand I_5796 (I101430,I101413,I415811);
not I_5797 (I101447,I415808);
nor I_5798 (I101464,I101447,I415826);
nand I_5799 (I101481,I101464,I415799);
nor I_5800 (I101498,I101481,I101430);
DFFARX1 I_5801 (I101498,I2859,I101280,I101248,);
not I_5802 (I101529,I101481);
not I_5803 (I101546,I415826);
nand I_5804 (I101563,I101546,I415811);
nor I_5805 (I101580,I415826,I415802);
nand I_5806 (I101260,I101396,I101580);
nand I_5807 (I101254,I101345,I415826);
nand I_5808 (I101625,I101447,I415805);
DFFARX1 I_5809 (I101625,I2859,I101280,I101269,);
DFFARX1 I_5810 (I101625,I2859,I101280,I101263,);
not I_5811 (I101670,I415805);
nor I_5812 (I101687,I101670,I415817);
and I_5813 (I101704,I101687,I415799);
or I_5814 (I101721,I101704,I415820);
DFFARX1 I_5815 (I101721,I2859,I101280,I101747,);
nand I_5816 (I101755,I101747,I101413);
nor I_5817 (I101257,I101755,I101563);
nor I_5818 (I101251,I101747,I101379);
DFFARX1 I_5819 (I101747,I2859,I101280,I101809,);
not I_5820 (I101817,I101809);
nor I_5821 (I101266,I101817,I101529);
not I_5822 (I101875,I2866);
DFFARX1 I_5823 (I158776,I2859,I101875,I101901,);
DFFARX1 I_5824 (I101901,I2859,I101875,I101918,);
not I_5825 (I101867,I101918);
not I_5826 (I101940,I101901);
DFFARX1 I_5827 (I158791,I2859,I101875,I101966,);
not I_5828 (I101974,I101966);
and I_5829 (I101991,I101940,I158788);
not I_5830 (I102008,I158776);
nand I_5831 (I102025,I102008,I158788);
not I_5832 (I102042,I158785);
nor I_5833 (I102059,I102042,I158800);
nand I_5834 (I102076,I102059,I158797);
nor I_5835 (I102093,I102076,I102025);
DFFARX1 I_5836 (I102093,I2859,I101875,I101843,);
not I_5837 (I102124,I102076);
not I_5838 (I102141,I158800);
nand I_5839 (I102158,I102141,I158788);
nor I_5840 (I102175,I158800,I158776);
nand I_5841 (I101855,I101991,I102175);
nand I_5842 (I101849,I101940,I158800);
nand I_5843 (I102220,I102042,I158794);
DFFARX1 I_5844 (I102220,I2859,I101875,I101864,);
DFFARX1 I_5845 (I102220,I2859,I101875,I101858,);
not I_5846 (I102265,I158794);
nor I_5847 (I102282,I102265,I158782);
and I_5848 (I102299,I102282,I158803);
or I_5849 (I102316,I102299,I158779);
DFFARX1 I_5850 (I102316,I2859,I101875,I102342,);
nand I_5851 (I102350,I102342,I102008);
nor I_5852 (I101852,I102350,I102158);
nor I_5853 (I101846,I102342,I101974);
DFFARX1 I_5854 (I102342,I2859,I101875,I102404,);
not I_5855 (I102412,I102404);
nor I_5856 (I101861,I102412,I102124);
not I_5857 (I102470,I2866);
DFFARX1 I_5858 (I265616,I2859,I102470,I102496,);
DFFARX1 I_5859 (I102496,I2859,I102470,I102513,);
not I_5860 (I102462,I102513);
not I_5861 (I102535,I102496);
DFFARX1 I_5862 (I265613,I2859,I102470,I102561,);
not I_5863 (I102569,I102561);
and I_5864 (I102586,I102535,I265619);
not I_5865 (I102603,I265604);
nand I_5866 (I102620,I102603,I265619);
not I_5867 (I102637,I265607);
nor I_5868 (I102654,I102637,I265628);
nand I_5869 (I102671,I102654,I265625);
nor I_5870 (I102688,I102671,I102620);
DFFARX1 I_5871 (I102688,I2859,I102470,I102438,);
not I_5872 (I102719,I102671);
not I_5873 (I102736,I265628);
nand I_5874 (I102753,I102736,I265619);
nor I_5875 (I102770,I265628,I265604);
nand I_5876 (I102450,I102586,I102770);
nand I_5877 (I102444,I102535,I265628);
nand I_5878 (I102815,I102637,I265604);
DFFARX1 I_5879 (I102815,I2859,I102470,I102459,);
DFFARX1 I_5880 (I102815,I2859,I102470,I102453,);
not I_5881 (I102860,I265604);
nor I_5882 (I102877,I102860,I265610);
and I_5883 (I102894,I102877,I265622);
or I_5884 (I102911,I102894,I265607);
DFFARX1 I_5885 (I102911,I2859,I102470,I102937,);
nand I_5886 (I102945,I102937,I102603);
nor I_5887 (I102447,I102945,I102753);
nor I_5888 (I102441,I102937,I102569);
DFFARX1 I_5889 (I102937,I2859,I102470,I102999,);
not I_5890 (I103007,I102999);
nor I_5891 (I102456,I103007,I102719);
not I_5892 (I103065,I2866);
DFFARX1 I_5893 (I434298,I2859,I103065,I103091,);
DFFARX1 I_5894 (I103091,I2859,I103065,I103108,);
not I_5895 (I103057,I103108);
not I_5896 (I103130,I103091);
DFFARX1 I_5897 (I434307,I2859,I103065,I103156,);
not I_5898 (I103164,I103156);
and I_5899 (I103181,I103130,I434301);
not I_5900 (I103198,I434295);
nand I_5901 (I103215,I103198,I434301);
not I_5902 (I103232,I434310);
nor I_5903 (I103249,I103232,I434298);
nand I_5904 (I103266,I103249,I434304);
nor I_5905 (I103283,I103266,I103215);
DFFARX1 I_5906 (I103283,I2859,I103065,I103033,);
not I_5907 (I103314,I103266);
not I_5908 (I103331,I434298);
nand I_5909 (I103348,I103331,I434301);
nor I_5910 (I103365,I434298,I434295);
nand I_5911 (I103045,I103181,I103365);
nand I_5912 (I103039,I103130,I434298);
nand I_5913 (I103410,I103232,I434301);
DFFARX1 I_5914 (I103410,I2859,I103065,I103054,);
DFFARX1 I_5915 (I103410,I2859,I103065,I103048,);
not I_5916 (I103455,I434301);
nor I_5917 (I103472,I103455,I434316);
and I_5918 (I103489,I103472,I434313);
or I_5919 (I103506,I103489,I434295);
DFFARX1 I_5920 (I103506,I2859,I103065,I103532,);
nand I_5921 (I103540,I103532,I103198);
nor I_5922 (I103042,I103540,I103348);
nor I_5923 (I103036,I103532,I103164);
DFFARX1 I_5924 (I103532,I2859,I103065,I103594,);
not I_5925 (I103602,I103594);
nor I_5926 (I103051,I103602,I103314);
not I_5927 (I103660,I2866);
DFFARX1 I_5928 (I528631,I2859,I103660,I103686,);
DFFARX1 I_5929 (I103686,I2859,I103660,I103703,);
not I_5930 (I103652,I103703);
not I_5931 (I103725,I103686);
DFFARX1 I_5932 (I528643,I2859,I103660,I103751,);
not I_5933 (I103759,I103751);
and I_5934 (I103776,I103725,I528637);
not I_5935 (I103793,I528649);
nand I_5936 (I103810,I103793,I528637);
not I_5937 (I103827,I528634);
nor I_5938 (I103844,I103827,I528646);
nand I_5939 (I103861,I103844,I528628);
nor I_5940 (I103878,I103861,I103810);
DFFARX1 I_5941 (I103878,I2859,I103660,I103628,);
not I_5942 (I103909,I103861);
not I_5943 (I103926,I528646);
nand I_5944 (I103943,I103926,I528637);
nor I_5945 (I103960,I528646,I528649);
nand I_5946 (I103640,I103776,I103960);
nand I_5947 (I103634,I103725,I528646);
nand I_5948 (I104005,I103827,I528640);
DFFARX1 I_5949 (I104005,I2859,I103660,I103649,);
DFFARX1 I_5950 (I104005,I2859,I103660,I103643,);
not I_5951 (I104050,I528640);
nor I_5952 (I104067,I104050,I528631);
and I_5953 (I104084,I104067,I528628);
or I_5954 (I104101,I104084,I528652);
DFFARX1 I_5955 (I104101,I2859,I103660,I104127,);
nand I_5956 (I104135,I104127,I103793);
nor I_5957 (I103637,I104135,I103943);
nor I_5958 (I103631,I104127,I103759);
DFFARX1 I_5959 (I104127,I2859,I103660,I104189,);
not I_5960 (I104197,I104189);
nor I_5961 (I103646,I104197,I103909);
not I_5962 (I104255,I2866);
DFFARX1 I_5963 (I134007,I2859,I104255,I104281,);
DFFARX1 I_5964 (I104281,I2859,I104255,I104298,);
not I_5965 (I104247,I104298);
not I_5966 (I104320,I104281);
DFFARX1 I_5967 (I134022,I2859,I104255,I104346,);
not I_5968 (I104354,I104346);
and I_5969 (I104371,I104320,I134019);
not I_5970 (I104388,I134007);
nand I_5971 (I104405,I104388,I134019);
not I_5972 (I104422,I134016);
nor I_5973 (I104439,I104422,I134031);
nand I_5974 (I104456,I104439,I134028);
nor I_5975 (I104473,I104456,I104405);
DFFARX1 I_5976 (I104473,I2859,I104255,I104223,);
not I_5977 (I104504,I104456);
not I_5978 (I104521,I134031);
nand I_5979 (I104538,I104521,I134019);
nor I_5980 (I104555,I134031,I134007);
nand I_5981 (I104235,I104371,I104555);
nand I_5982 (I104229,I104320,I134031);
nand I_5983 (I104600,I104422,I134025);
DFFARX1 I_5984 (I104600,I2859,I104255,I104244,);
DFFARX1 I_5985 (I104600,I2859,I104255,I104238,);
not I_5986 (I104645,I134025);
nor I_5987 (I104662,I104645,I134013);
and I_5988 (I104679,I104662,I134034);
or I_5989 (I104696,I104679,I134010);
DFFARX1 I_5990 (I104696,I2859,I104255,I104722,);
nand I_5991 (I104730,I104722,I104388);
nor I_5992 (I104232,I104730,I104538);
nor I_5993 (I104226,I104722,I104354);
DFFARX1 I_5994 (I104722,I2859,I104255,I104784,);
not I_5995 (I104792,I104784);
nor I_5996 (I104241,I104792,I104504);
not I_5997 (I104850,I2866);
DFFARX1 I_5998 (I219070,I2859,I104850,I104876,);
DFFARX1 I_5999 (I104876,I2859,I104850,I104893,);
not I_6000 (I104842,I104893);
not I_6001 (I104915,I104876);
DFFARX1 I_6002 (I219064,I2859,I104850,I104941,);
not I_6003 (I104949,I104941);
and I_6004 (I104966,I104915,I219079);
not I_6005 (I104983,I219076);
nand I_6006 (I105000,I104983,I219079);
not I_6007 (I105017,I219067);
nor I_6008 (I105034,I105017,I219058);
nand I_6009 (I105051,I105034,I219061);
nor I_6010 (I105068,I105051,I105000);
DFFARX1 I_6011 (I105068,I2859,I104850,I104818,);
not I_6012 (I105099,I105051);
not I_6013 (I105116,I219058);
nand I_6014 (I105133,I105116,I219079);
nor I_6015 (I105150,I219058,I219076);
nand I_6016 (I104830,I104966,I105150);
nand I_6017 (I104824,I104915,I219058);
nand I_6018 (I105195,I105017,I219082);
DFFARX1 I_6019 (I105195,I2859,I104850,I104839,);
DFFARX1 I_6020 (I105195,I2859,I104850,I104833,);
not I_6021 (I105240,I219082);
nor I_6022 (I105257,I105240,I219073);
and I_6023 (I105274,I105257,I219058);
or I_6024 (I105291,I105274,I219061);
DFFARX1 I_6025 (I105291,I2859,I104850,I105317,);
nand I_6026 (I105325,I105317,I104983);
nor I_6027 (I104827,I105325,I105133);
nor I_6028 (I104821,I105317,I104949);
DFFARX1 I_6029 (I105317,I2859,I104850,I105379,);
not I_6030 (I105387,I105379);
nor I_6031 (I104836,I105387,I105099);
not I_6032 (I105445,I2866);
DFFARX1 I_6033 (I339509,I2859,I105445,I105471,);
DFFARX1 I_6034 (I105471,I2859,I105445,I105488,);
not I_6035 (I105437,I105488);
not I_6036 (I105510,I105471);
DFFARX1 I_6037 (I339503,I2859,I105445,I105536,);
not I_6038 (I105544,I105536);
and I_6039 (I105561,I105510,I339521);
not I_6040 (I105578,I339509);
nand I_6041 (I105595,I105578,I339521);
not I_6042 (I105612,I339503);
nor I_6043 (I105629,I105612,I339515);
nand I_6044 (I105646,I105629,I339506);
nor I_6045 (I105663,I105646,I105595);
DFFARX1 I_6046 (I105663,I2859,I105445,I105413,);
not I_6047 (I105694,I105646);
not I_6048 (I105711,I339515);
nand I_6049 (I105728,I105711,I339521);
nor I_6050 (I105745,I339515,I339509);
nand I_6051 (I105425,I105561,I105745);
nand I_6052 (I105419,I105510,I339515);
nand I_6053 (I105790,I105612,I339518);
DFFARX1 I_6054 (I105790,I2859,I105445,I105434,);
DFFARX1 I_6055 (I105790,I2859,I105445,I105428,);
not I_6056 (I105835,I339518);
nor I_6057 (I105852,I105835,I339524);
and I_6058 (I105869,I105852,I339506);
or I_6059 (I105886,I105869,I339512);
DFFARX1 I_6060 (I105886,I2859,I105445,I105912,);
nand I_6061 (I105920,I105912,I105578);
nor I_6062 (I105422,I105920,I105728);
nor I_6063 (I105416,I105912,I105544);
DFFARX1 I_6064 (I105912,I2859,I105445,I105974,);
not I_6065 (I105982,I105974);
nor I_6066 (I105431,I105982,I105694);
not I_6067 (I106040,I2866);
DFFARX1 I_6068 (I150344,I2859,I106040,I106066,);
DFFARX1 I_6069 (I106066,I2859,I106040,I106083,);
not I_6070 (I106032,I106083);
not I_6071 (I106105,I106066);
DFFARX1 I_6072 (I150359,I2859,I106040,I106131,);
not I_6073 (I106139,I106131);
and I_6074 (I106156,I106105,I150356);
not I_6075 (I106173,I150344);
nand I_6076 (I106190,I106173,I150356);
not I_6077 (I106207,I150353);
nor I_6078 (I106224,I106207,I150368);
nand I_6079 (I106241,I106224,I150365);
nor I_6080 (I106258,I106241,I106190);
DFFARX1 I_6081 (I106258,I2859,I106040,I106008,);
not I_6082 (I106289,I106241);
not I_6083 (I106306,I150368);
nand I_6084 (I106323,I106306,I150356);
nor I_6085 (I106340,I150368,I150344);
nand I_6086 (I106020,I106156,I106340);
nand I_6087 (I106014,I106105,I150368);
nand I_6088 (I106385,I106207,I150362);
DFFARX1 I_6089 (I106385,I2859,I106040,I106029,);
DFFARX1 I_6090 (I106385,I2859,I106040,I106023,);
not I_6091 (I106430,I150362);
nor I_6092 (I106447,I106430,I150350);
and I_6093 (I106464,I106447,I150371);
or I_6094 (I106481,I106464,I150347);
DFFARX1 I_6095 (I106481,I2859,I106040,I106507,);
nand I_6096 (I106515,I106507,I106173);
nor I_6097 (I106017,I106515,I106323);
nor I_6098 (I106011,I106507,I106139);
DFFARX1 I_6099 (I106507,I2859,I106040,I106569,);
not I_6100 (I106577,I106569);
nor I_6101 (I106026,I106577,I106289);
not I_6102 (I106638,I2866);
DFFARX1 I_6103 (I2676,I2859,I106638,I106664,);
nand I_6104 (I106672,I2612,I2556);
and I_6105 (I106689,I106672,I1388);
DFFARX1 I_6106 (I106689,I2859,I106638,I106715,);
nor I_6107 (I106606,I106715,I106664);
not I_6108 (I106737,I106715);
DFFARX1 I_6109 (I2772,I2859,I106638,I106763,);
nand I_6110 (I106771,I106763,I2548);
not I_6111 (I106788,I106771);
DFFARX1 I_6112 (I106788,I2859,I106638,I106814,);
not I_6113 (I106630,I106814);
nor I_6114 (I106836,I106664,I106771);
nor I_6115 (I106612,I106715,I106836);
DFFARX1 I_6116 (I1804,I2859,I106638,I106876,);
DFFARX1 I_6117 (I106876,I2859,I106638,I106893,);
not I_6118 (I106901,I106893);
not I_6119 (I106918,I106876);
nand I_6120 (I106615,I106918,I106737);
nand I_6121 (I106949,I1780,I1764);
and I_6122 (I106966,I106949,I2140);
DFFARX1 I_6123 (I106966,I2859,I106638,I106992,);
nor I_6124 (I107000,I106992,I106664);
DFFARX1 I_6125 (I107000,I2859,I106638,I106603,);
DFFARX1 I_6126 (I106992,I2859,I106638,I106621,);
nor I_6127 (I107045,I1820,I1764);
not I_6128 (I107062,I107045);
nor I_6129 (I106624,I106901,I107062);
nand I_6130 (I106609,I106918,I107062);
nor I_6131 (I106618,I106664,I107045);
DFFARX1 I_6132 (I107045,I2859,I106638,I106627,);
not I_6133 (I107165,I2866);
DFFARX1 I_6134 (I48925,I2859,I107165,I107191,);
nand I_6135 (I107199,I48937,I48946);
and I_6136 (I107216,I107199,I48925);
DFFARX1 I_6137 (I107216,I2859,I107165,I107242,);
nor I_6138 (I107133,I107242,I107191);
not I_6139 (I107264,I107242);
DFFARX1 I_6140 (I48940,I2859,I107165,I107290,);
nand I_6141 (I107298,I107290,I48928);
not I_6142 (I107315,I107298);
DFFARX1 I_6143 (I107315,I2859,I107165,I107341,);
not I_6144 (I107157,I107341);
nor I_6145 (I107363,I107191,I107298);
nor I_6146 (I107139,I107242,I107363);
DFFARX1 I_6147 (I48931,I2859,I107165,I107403,);
DFFARX1 I_6148 (I107403,I2859,I107165,I107420,);
not I_6149 (I107428,I107420);
not I_6150 (I107445,I107403);
nand I_6151 (I107142,I107445,I107264);
nand I_6152 (I107476,I48922,I48922);
and I_6153 (I107493,I107476,I48934);
DFFARX1 I_6154 (I107493,I2859,I107165,I107519,);
nor I_6155 (I107527,I107519,I107191);
DFFARX1 I_6156 (I107527,I2859,I107165,I107130,);
DFFARX1 I_6157 (I107519,I2859,I107165,I107148,);
nor I_6158 (I107572,I48943,I48922);
not I_6159 (I107589,I107572);
nor I_6160 (I107151,I107428,I107589);
nand I_6161 (I107136,I107445,I107589);
nor I_6162 (I107145,I107191,I107572);
DFFARX1 I_6163 (I107572,I2859,I107165,I107154,);
not I_6164 (I107692,I2866);
DFFARX1 I_6165 (I34169,I2859,I107692,I107718,);
nand I_6166 (I107726,I34181,I34190);
and I_6167 (I107743,I107726,I34169);
DFFARX1 I_6168 (I107743,I2859,I107692,I107769,);
nor I_6169 (I107660,I107769,I107718);
not I_6170 (I107791,I107769);
DFFARX1 I_6171 (I34184,I2859,I107692,I107817,);
nand I_6172 (I107825,I107817,I34172);
not I_6173 (I107842,I107825);
DFFARX1 I_6174 (I107842,I2859,I107692,I107868,);
not I_6175 (I107684,I107868);
nor I_6176 (I107890,I107718,I107825);
nor I_6177 (I107666,I107769,I107890);
DFFARX1 I_6178 (I34175,I2859,I107692,I107930,);
DFFARX1 I_6179 (I107930,I2859,I107692,I107947,);
not I_6180 (I107955,I107947);
not I_6181 (I107972,I107930);
nand I_6182 (I107669,I107972,I107791);
nand I_6183 (I108003,I34166,I34166);
and I_6184 (I108020,I108003,I34178);
DFFARX1 I_6185 (I108020,I2859,I107692,I108046,);
nor I_6186 (I108054,I108046,I107718);
DFFARX1 I_6187 (I108054,I2859,I107692,I107657,);
DFFARX1 I_6188 (I108046,I2859,I107692,I107675,);
nor I_6189 (I108099,I34187,I34166);
not I_6190 (I108116,I108099);
nor I_6191 (I107678,I107955,I108116);
nand I_6192 (I107663,I107972,I108116);
nor I_6193 (I107672,I107718,I108099);
DFFARX1 I_6194 (I108099,I2859,I107692,I107681,);
not I_6195 (I108219,I2866);
DFFARX1 I_6196 (I341087,I2859,I108219,I108245,);
nand I_6197 (I108253,I341090,I341084);
and I_6198 (I108270,I108253,I341096);
DFFARX1 I_6199 (I108270,I2859,I108219,I108296,);
nor I_6200 (I108187,I108296,I108245);
not I_6201 (I108318,I108296);
DFFARX1 I_6202 (I341099,I2859,I108219,I108344,);
nand I_6203 (I108352,I108344,I341090);
not I_6204 (I108369,I108352);
DFFARX1 I_6205 (I108369,I2859,I108219,I108395,);
not I_6206 (I108211,I108395);
nor I_6207 (I108417,I108245,I108352);
nor I_6208 (I108193,I108296,I108417);
DFFARX1 I_6209 (I341102,I2859,I108219,I108457,);
DFFARX1 I_6210 (I108457,I2859,I108219,I108474,);
not I_6211 (I108482,I108474);
not I_6212 (I108499,I108457);
nand I_6213 (I108196,I108499,I108318);
nand I_6214 (I108530,I341084,I341093);
and I_6215 (I108547,I108530,I341087);
DFFARX1 I_6216 (I108547,I2859,I108219,I108573,);
nor I_6217 (I108581,I108573,I108245);
DFFARX1 I_6218 (I108581,I2859,I108219,I108184,);
DFFARX1 I_6219 (I108573,I2859,I108219,I108202,);
nor I_6220 (I108626,I341105,I341093);
not I_6221 (I108643,I108626);
nor I_6222 (I108205,I108482,I108643);
nand I_6223 (I108190,I108499,I108643);
nor I_6224 (I108199,I108245,I108626);
DFFARX1 I_6225 (I108626,I2859,I108219,I108208,);
not I_6226 (I108746,I2866);
DFFARX1 I_6227 (I283534,I2859,I108746,I108772,);
nand I_6228 (I108780,I283525,I283540);
and I_6229 (I108797,I108780,I283546);
DFFARX1 I_6230 (I108797,I2859,I108746,I108823,);
nor I_6231 (I108714,I108823,I108772);
not I_6232 (I108845,I108823);
DFFARX1 I_6233 (I283531,I2859,I108746,I108871,);
nand I_6234 (I108879,I108871,I283525);
not I_6235 (I108896,I108879);
DFFARX1 I_6236 (I108896,I2859,I108746,I108922,);
not I_6237 (I108738,I108922);
nor I_6238 (I108944,I108772,I108879);
nor I_6239 (I108720,I108823,I108944);
DFFARX1 I_6240 (I283528,I2859,I108746,I108984,);
DFFARX1 I_6241 (I108984,I2859,I108746,I109001,);
not I_6242 (I109009,I109001);
not I_6243 (I109026,I108984);
nand I_6244 (I108723,I109026,I108845);
nand I_6245 (I109057,I283522,I283537);
and I_6246 (I109074,I109057,I283522);
DFFARX1 I_6247 (I109074,I2859,I108746,I109100,);
nor I_6248 (I109108,I109100,I108772);
DFFARX1 I_6249 (I109108,I2859,I108746,I108711,);
DFFARX1 I_6250 (I109100,I2859,I108746,I108729,);
nor I_6251 (I109153,I283543,I283537);
not I_6252 (I109170,I109153);
nor I_6253 (I108732,I109009,I109170);
nand I_6254 (I108717,I109026,I109170);
nor I_6255 (I108726,I108772,I109153);
DFFARX1 I_6256 (I109153,I2859,I108746,I108735,);
not I_6257 (I109273,I2866);
DFFARX1 I_6258 (I249435,I2859,I109273,I109299,);
nand I_6259 (I109307,I249420,I249423);
and I_6260 (I109324,I109307,I249438);
DFFARX1 I_6261 (I109324,I2859,I109273,I109350,);
nor I_6262 (I109241,I109350,I109299);
not I_6263 (I109372,I109350);
DFFARX1 I_6264 (I249432,I2859,I109273,I109398,);
nand I_6265 (I109406,I109398,I249423);
not I_6266 (I109423,I109406);
DFFARX1 I_6267 (I109423,I2859,I109273,I109449,);
not I_6268 (I109265,I109449);
nor I_6269 (I109471,I109299,I109406);
nor I_6270 (I109247,I109350,I109471);
DFFARX1 I_6271 (I249429,I2859,I109273,I109511,);
DFFARX1 I_6272 (I109511,I2859,I109273,I109528,);
not I_6273 (I109536,I109528);
not I_6274 (I109553,I109511);
nand I_6275 (I109250,I109553,I109372);
nand I_6276 (I109584,I249444,I249420);
and I_6277 (I109601,I109584,I249441);
DFFARX1 I_6278 (I109601,I2859,I109273,I109627,);
nor I_6279 (I109635,I109627,I109299);
DFFARX1 I_6280 (I109635,I2859,I109273,I109238,);
DFFARX1 I_6281 (I109627,I2859,I109273,I109256,);
nor I_6282 (I109680,I249426,I249420);
not I_6283 (I109697,I109680);
nor I_6284 (I109259,I109536,I109697);
nand I_6285 (I109244,I109553,I109697);
nor I_6286 (I109253,I109299,I109680);
DFFARX1 I_6287 (I109680,I2859,I109273,I109262,);
not I_6288 (I109800,I2866);
DFFARX1 I_6289 (I11505,I2859,I109800,I109826,);
nand I_6290 (I109834,I11529,I11508);
and I_6291 (I109851,I109834,I11505);
DFFARX1 I_6292 (I109851,I2859,I109800,I109877,);
nor I_6293 (I109768,I109877,I109826);
not I_6294 (I109899,I109877);
DFFARX1 I_6295 (I11511,I2859,I109800,I109925,);
nand I_6296 (I109933,I109925,I11520);
not I_6297 (I109950,I109933);
DFFARX1 I_6298 (I109950,I2859,I109800,I109976,);
not I_6299 (I109792,I109976);
nor I_6300 (I109998,I109826,I109933);
nor I_6301 (I109774,I109877,I109998);
DFFARX1 I_6302 (I11514,I2859,I109800,I110038,);
DFFARX1 I_6303 (I110038,I2859,I109800,I110055,);
not I_6304 (I110063,I110055);
not I_6305 (I110080,I110038);
nand I_6306 (I109777,I110080,I109899);
nand I_6307 (I110111,I11526,I11508);
and I_6308 (I110128,I110111,I11517);
DFFARX1 I_6309 (I110128,I2859,I109800,I110154,);
nor I_6310 (I110162,I110154,I109826);
DFFARX1 I_6311 (I110162,I2859,I109800,I109765,);
DFFARX1 I_6312 (I110154,I2859,I109800,I109783,);
nor I_6313 (I110207,I11523,I11508);
not I_6314 (I110224,I110207);
nor I_6315 (I109786,I110063,I110224);
nand I_6316 (I109771,I110080,I110224);
nor I_6317 (I109780,I109826,I110207);
DFFARX1 I_6318 (I110207,I2859,I109800,I109789,);
not I_6319 (I110327,I2866);
DFFARX1 I_6320 (I205895,I2859,I110327,I110353,);
nand I_6321 (I110361,I205907,I205886);
and I_6322 (I110378,I110361,I205910);
DFFARX1 I_6323 (I110378,I2859,I110327,I110404,);
nor I_6324 (I110295,I110404,I110353);
not I_6325 (I110426,I110404);
DFFARX1 I_6326 (I205901,I2859,I110327,I110452,);
nand I_6327 (I110460,I110452,I205883);
not I_6328 (I110477,I110460);
DFFARX1 I_6329 (I110477,I2859,I110327,I110503,);
not I_6330 (I110319,I110503);
nor I_6331 (I110525,I110353,I110460);
nor I_6332 (I110301,I110404,I110525);
DFFARX1 I_6333 (I205898,I2859,I110327,I110565,);
DFFARX1 I_6334 (I110565,I2859,I110327,I110582,);
not I_6335 (I110590,I110582);
not I_6336 (I110607,I110565);
nand I_6337 (I110304,I110607,I110426);
nand I_6338 (I110638,I205883,I205889);
and I_6339 (I110655,I110638,I205892);
DFFARX1 I_6340 (I110655,I2859,I110327,I110681,);
nor I_6341 (I110689,I110681,I110353);
DFFARX1 I_6342 (I110689,I2859,I110327,I110292,);
DFFARX1 I_6343 (I110681,I2859,I110327,I110310,);
nor I_6344 (I110734,I205904,I205889);
not I_6345 (I110751,I110734);
nor I_6346 (I110313,I110590,I110751);
nand I_6347 (I110298,I110607,I110751);
nor I_6348 (I110307,I110353,I110734);
DFFARX1 I_6349 (I110734,I2859,I110327,I110316,);
not I_6350 (I110854,I2866);
DFFARX1 I_6351 (I98868,I2859,I110854,I110880,);
nand I_6352 (I110888,I98868,I98874);
and I_6353 (I110905,I110888,I98892);
DFFARX1 I_6354 (I110905,I2859,I110854,I110931,);
nor I_6355 (I110822,I110931,I110880);
not I_6356 (I110953,I110931);
DFFARX1 I_6357 (I98880,I2859,I110854,I110979,);
nand I_6358 (I110987,I110979,I98877);
not I_6359 (I111004,I110987);
DFFARX1 I_6360 (I111004,I2859,I110854,I111030,);
not I_6361 (I110846,I111030);
nor I_6362 (I111052,I110880,I110987);
nor I_6363 (I110828,I110931,I111052);
DFFARX1 I_6364 (I98886,I2859,I110854,I111092,);
DFFARX1 I_6365 (I111092,I2859,I110854,I111109,);
not I_6366 (I111117,I111109);
not I_6367 (I111134,I111092);
nand I_6368 (I110831,I111134,I110953);
nand I_6369 (I111165,I98871,I98871);
and I_6370 (I111182,I111165,I98883);
DFFARX1 I_6371 (I111182,I2859,I110854,I111208,);
nor I_6372 (I111216,I111208,I110880);
DFFARX1 I_6373 (I111216,I2859,I110854,I110819,);
DFFARX1 I_6374 (I111208,I2859,I110854,I110837,);
nor I_6375 (I111261,I98889,I98871);
not I_6376 (I111278,I111261);
nor I_6377 (I110840,I111117,I111278);
nand I_6378 (I110825,I111134,I111278);
nor I_6379 (I110834,I110880,I111261);
DFFARX1 I_6380 (I111261,I2859,I110854,I110843,);
not I_6381 (I111381,I2866);
DFFARX1 I_6382 (I448898,I2859,I111381,I111407,);
nand I_6383 (I111415,I448913,I448898);
and I_6384 (I111432,I111415,I448916);
DFFARX1 I_6385 (I111432,I2859,I111381,I111458,);
nor I_6386 (I111349,I111458,I111407);
not I_6387 (I111480,I111458);
DFFARX1 I_6388 (I448922,I2859,I111381,I111506,);
nand I_6389 (I111514,I111506,I448904);
not I_6390 (I111531,I111514);
DFFARX1 I_6391 (I111531,I2859,I111381,I111557,);
not I_6392 (I111373,I111557);
nor I_6393 (I111579,I111407,I111514);
nor I_6394 (I111355,I111458,I111579);
DFFARX1 I_6395 (I448901,I2859,I111381,I111619,);
DFFARX1 I_6396 (I111619,I2859,I111381,I111636,);
not I_6397 (I111644,I111636);
not I_6398 (I111661,I111619);
nand I_6399 (I111358,I111661,I111480);
nand I_6400 (I111692,I448901,I448907);
and I_6401 (I111709,I111692,I448919);
DFFARX1 I_6402 (I111709,I2859,I111381,I111735,);
nor I_6403 (I111743,I111735,I111407);
DFFARX1 I_6404 (I111743,I2859,I111381,I111346,);
DFFARX1 I_6405 (I111735,I2859,I111381,I111364,);
nor I_6406 (I111788,I448910,I448907);
not I_6407 (I111805,I111788);
nor I_6408 (I111367,I111644,I111805);
nand I_6409 (I111352,I111661,I111805);
nor I_6410 (I111361,I111407,I111788);
DFFARX1 I_6411 (I111788,I2859,I111381,I111370,);
not I_6412 (I111908,I2866);
DFFARX1 I_6413 (I458146,I2859,I111908,I111934,);
nand I_6414 (I111942,I458161,I458146);
and I_6415 (I111959,I111942,I458164);
DFFARX1 I_6416 (I111959,I2859,I111908,I111985,);
nor I_6417 (I111876,I111985,I111934);
not I_6418 (I112007,I111985);
DFFARX1 I_6419 (I458170,I2859,I111908,I112033,);
nand I_6420 (I112041,I112033,I458152);
not I_6421 (I112058,I112041);
DFFARX1 I_6422 (I112058,I2859,I111908,I112084,);
not I_6423 (I111900,I112084);
nor I_6424 (I112106,I111934,I112041);
nor I_6425 (I111882,I111985,I112106);
DFFARX1 I_6426 (I458149,I2859,I111908,I112146,);
DFFARX1 I_6427 (I112146,I2859,I111908,I112163,);
not I_6428 (I112171,I112163);
not I_6429 (I112188,I112146);
nand I_6430 (I111885,I112188,I112007);
nand I_6431 (I112219,I458149,I458155);
and I_6432 (I112236,I112219,I458167);
DFFARX1 I_6433 (I112236,I2859,I111908,I112262,);
nor I_6434 (I112270,I112262,I111934);
DFFARX1 I_6435 (I112270,I2859,I111908,I111873,);
DFFARX1 I_6436 (I112262,I2859,I111908,I111891,);
nor I_6437 (I112315,I458158,I458155);
not I_6438 (I112332,I112315);
nor I_6439 (I111894,I112171,I112332);
nand I_6440 (I111879,I112188,I112332);
nor I_6441 (I111888,I111934,I112315);
DFFARX1 I_6442 (I112315,I2859,I111908,I111897,);
not I_6443 (I112435,I2866);
DFFARX1 I_6444 (I349519,I2859,I112435,I112461,);
nand I_6445 (I112469,I349522,I349516);
and I_6446 (I112486,I112469,I349528);
DFFARX1 I_6447 (I112486,I2859,I112435,I112512,);
nor I_6448 (I112403,I112512,I112461);
not I_6449 (I112534,I112512);
DFFARX1 I_6450 (I349531,I2859,I112435,I112560,);
nand I_6451 (I112568,I112560,I349522);
not I_6452 (I112585,I112568);
DFFARX1 I_6453 (I112585,I2859,I112435,I112611,);
not I_6454 (I112427,I112611);
nor I_6455 (I112633,I112461,I112568);
nor I_6456 (I112409,I112512,I112633);
DFFARX1 I_6457 (I349534,I2859,I112435,I112673,);
DFFARX1 I_6458 (I112673,I2859,I112435,I112690,);
not I_6459 (I112698,I112690);
not I_6460 (I112715,I112673);
nand I_6461 (I112412,I112715,I112534);
nand I_6462 (I112746,I349516,I349525);
and I_6463 (I112763,I112746,I349519);
DFFARX1 I_6464 (I112763,I2859,I112435,I112789,);
nor I_6465 (I112797,I112789,I112461);
DFFARX1 I_6466 (I112797,I2859,I112435,I112400,);
DFFARX1 I_6467 (I112789,I2859,I112435,I112418,);
nor I_6468 (I112842,I349537,I349525);
not I_6469 (I112859,I112842);
nor I_6470 (I112421,I112698,I112859);
nand I_6471 (I112406,I112715,I112859);
nor I_6472 (I112415,I112461,I112842);
DFFARX1 I_6473 (I112842,I2859,I112435,I112424,);
not I_6474 (I112962,I2866);
DFFARX1 I_6475 (I230361,I2859,I112962,I112988,);
nand I_6476 (I112996,I230346,I230349);
and I_6477 (I113013,I112996,I230364);
DFFARX1 I_6478 (I113013,I2859,I112962,I113039,);
nor I_6479 (I112930,I113039,I112988);
not I_6480 (I113061,I113039);
DFFARX1 I_6481 (I230358,I2859,I112962,I113087,);
nand I_6482 (I113095,I113087,I230349);
not I_6483 (I113112,I113095);
DFFARX1 I_6484 (I113112,I2859,I112962,I113138,);
not I_6485 (I112954,I113138);
nor I_6486 (I113160,I112988,I113095);
nor I_6487 (I112936,I113039,I113160);
DFFARX1 I_6488 (I230355,I2859,I112962,I113200,);
DFFARX1 I_6489 (I113200,I2859,I112962,I113217,);
not I_6490 (I113225,I113217);
not I_6491 (I113242,I113200);
nand I_6492 (I112939,I113242,I113061);
nand I_6493 (I113273,I230370,I230346);
and I_6494 (I113290,I113273,I230367);
DFFARX1 I_6495 (I113290,I2859,I112962,I113316,);
nor I_6496 (I113324,I113316,I112988);
DFFARX1 I_6497 (I113324,I2859,I112962,I112927,);
DFFARX1 I_6498 (I113316,I2859,I112962,I112945,);
nor I_6499 (I113369,I230352,I230346);
not I_6500 (I113386,I113369);
nor I_6501 (I112948,I113225,I113386);
nand I_6502 (I112933,I113242,I113386);
nor I_6503 (I112942,I112988,I113369);
DFFARX1 I_6504 (I113369,I2859,I112962,I112951,);
not I_6505 (I113489,I2866);
DFFARX1 I_6506 (I26791,I2859,I113489,I113515,);
nand I_6507 (I113523,I26803,I26812);
and I_6508 (I113540,I113523,I26791);
DFFARX1 I_6509 (I113540,I2859,I113489,I113566,);
nor I_6510 (I113457,I113566,I113515);
not I_6511 (I113588,I113566);
DFFARX1 I_6512 (I26806,I2859,I113489,I113614,);
nand I_6513 (I113622,I113614,I26794);
not I_6514 (I113639,I113622);
DFFARX1 I_6515 (I113639,I2859,I113489,I113665,);
not I_6516 (I113481,I113665);
nor I_6517 (I113687,I113515,I113622);
nor I_6518 (I113463,I113566,I113687);
DFFARX1 I_6519 (I26797,I2859,I113489,I113727,);
DFFARX1 I_6520 (I113727,I2859,I113489,I113744,);
not I_6521 (I113752,I113744);
not I_6522 (I113769,I113727);
nand I_6523 (I113466,I113769,I113588);
nand I_6524 (I113800,I26788,I26788);
and I_6525 (I113817,I113800,I26800);
DFFARX1 I_6526 (I113817,I2859,I113489,I113843,);
nor I_6527 (I113851,I113843,I113515);
DFFARX1 I_6528 (I113851,I2859,I113489,I113454,);
DFFARX1 I_6529 (I113843,I2859,I113489,I113472,);
nor I_6530 (I113896,I26809,I26788);
not I_6531 (I113913,I113896);
nor I_6532 (I113475,I113752,I113913);
nand I_6533 (I113460,I113769,I113913);
nor I_6534 (I113469,I113515,I113896);
DFFARX1 I_6535 (I113896,I2859,I113489,I113478,);
not I_6536 (I114016,I2866);
DFFARX1 I_6537 (I95893,I2859,I114016,I114042,);
nand I_6538 (I114050,I95893,I95899);
and I_6539 (I114067,I114050,I95917);
DFFARX1 I_6540 (I114067,I2859,I114016,I114093,);
nor I_6541 (I113984,I114093,I114042);
not I_6542 (I114115,I114093);
DFFARX1 I_6543 (I95905,I2859,I114016,I114141,);
nand I_6544 (I114149,I114141,I95902);
not I_6545 (I114166,I114149);
DFFARX1 I_6546 (I114166,I2859,I114016,I114192,);
not I_6547 (I114008,I114192);
nor I_6548 (I114214,I114042,I114149);
nor I_6549 (I113990,I114093,I114214);
DFFARX1 I_6550 (I95911,I2859,I114016,I114254,);
DFFARX1 I_6551 (I114254,I2859,I114016,I114271,);
not I_6552 (I114279,I114271);
not I_6553 (I114296,I114254);
nand I_6554 (I113993,I114296,I114115);
nand I_6555 (I114327,I95896,I95896);
and I_6556 (I114344,I114327,I95908);
DFFARX1 I_6557 (I114344,I2859,I114016,I114370,);
nor I_6558 (I114378,I114370,I114042);
DFFARX1 I_6559 (I114378,I2859,I114016,I113981,);
DFFARX1 I_6560 (I114370,I2859,I114016,I113999,);
nor I_6561 (I114423,I95914,I95896);
not I_6562 (I114440,I114423);
nor I_6563 (I114002,I114279,I114440);
nand I_6564 (I113987,I114296,I114440);
nor I_6565 (I113996,I114042,I114423);
DFFARX1 I_6566 (I114423,I2859,I114016,I114005,);
not I_6567 (I114543,I2866);
DFFARX1 I_6568 (I522863,I2859,I114543,I114569,);
nand I_6569 (I114577,I522860,I522851);
and I_6570 (I114594,I114577,I522848);
DFFARX1 I_6571 (I114594,I2859,I114543,I114620,);
nor I_6572 (I114511,I114620,I114569);
not I_6573 (I114642,I114620);
DFFARX1 I_6574 (I522857,I2859,I114543,I114668,);
nand I_6575 (I114676,I114668,I522866);
not I_6576 (I114693,I114676);
DFFARX1 I_6577 (I114693,I2859,I114543,I114719,);
not I_6578 (I114535,I114719);
nor I_6579 (I114741,I114569,I114676);
nor I_6580 (I114517,I114620,I114741);
DFFARX1 I_6581 (I522869,I2859,I114543,I114781,);
DFFARX1 I_6582 (I114781,I2859,I114543,I114798,);
not I_6583 (I114806,I114798);
not I_6584 (I114823,I114781);
nand I_6585 (I114520,I114823,I114642);
nand I_6586 (I114854,I522848,I522854);
and I_6587 (I114871,I114854,I522872);
DFFARX1 I_6588 (I114871,I2859,I114543,I114897,);
nor I_6589 (I114905,I114897,I114569);
DFFARX1 I_6590 (I114905,I2859,I114543,I114508,);
DFFARX1 I_6591 (I114897,I2859,I114543,I114526,);
nor I_6592 (I114950,I522851,I522854);
not I_6593 (I114967,I114950);
nor I_6594 (I114529,I114806,I114967);
nand I_6595 (I114514,I114823,I114967);
nor I_6596 (I114523,I114569,I114950);
DFFARX1 I_6597 (I114950,I2859,I114543,I114532,);
not I_6598 (I115070,I2866);
DFFARX1 I_6599 (I356370,I2859,I115070,I115096,);
nand I_6600 (I115104,I356373,I356367);
and I_6601 (I115121,I115104,I356379);
DFFARX1 I_6602 (I115121,I2859,I115070,I115147,);
nor I_6603 (I115038,I115147,I115096);
not I_6604 (I115169,I115147);
DFFARX1 I_6605 (I356382,I2859,I115070,I115195,);
nand I_6606 (I115203,I115195,I356373);
not I_6607 (I115220,I115203);
DFFARX1 I_6608 (I115220,I2859,I115070,I115246,);
not I_6609 (I115062,I115246);
nor I_6610 (I115268,I115096,I115203);
nor I_6611 (I115044,I115147,I115268);
DFFARX1 I_6612 (I356385,I2859,I115070,I115308,);
DFFARX1 I_6613 (I115308,I2859,I115070,I115325,);
not I_6614 (I115333,I115325);
not I_6615 (I115350,I115308);
nand I_6616 (I115047,I115350,I115169);
nand I_6617 (I115381,I356367,I356376);
and I_6618 (I115398,I115381,I356370);
DFFARX1 I_6619 (I115398,I2859,I115070,I115424,);
nor I_6620 (I115432,I115424,I115096);
DFFARX1 I_6621 (I115432,I2859,I115070,I115035,);
DFFARX1 I_6622 (I115424,I2859,I115070,I115053,);
nor I_6623 (I115477,I356388,I356376);
not I_6624 (I115494,I115477);
nor I_6625 (I115056,I115333,I115494);
nand I_6626 (I115041,I115350,I115494);
nor I_6627 (I115050,I115096,I115477);
DFFARX1 I_6628 (I115477,I2859,I115070,I115059,);
not I_6629 (I115597,I2866);
DFFARX1 I_6630 (I93513,I2859,I115597,I115623,);
nand I_6631 (I115631,I93513,I93519);
and I_6632 (I115648,I115631,I93537);
DFFARX1 I_6633 (I115648,I2859,I115597,I115674,);
nor I_6634 (I115565,I115674,I115623);
not I_6635 (I115696,I115674);
DFFARX1 I_6636 (I93525,I2859,I115597,I115722,);
nand I_6637 (I115730,I115722,I93522);
not I_6638 (I115747,I115730);
DFFARX1 I_6639 (I115747,I2859,I115597,I115773,);
not I_6640 (I115589,I115773);
nor I_6641 (I115795,I115623,I115730);
nor I_6642 (I115571,I115674,I115795);
DFFARX1 I_6643 (I93531,I2859,I115597,I115835,);
DFFARX1 I_6644 (I115835,I2859,I115597,I115852,);
not I_6645 (I115860,I115852);
not I_6646 (I115877,I115835);
nand I_6647 (I115574,I115877,I115696);
nand I_6648 (I115908,I93516,I93516);
and I_6649 (I115925,I115908,I93528);
DFFARX1 I_6650 (I115925,I2859,I115597,I115951,);
nor I_6651 (I115959,I115951,I115623);
DFFARX1 I_6652 (I115959,I2859,I115597,I115562,);
DFFARX1 I_6653 (I115951,I2859,I115597,I115580,);
nor I_6654 (I116004,I93534,I93516);
not I_6655 (I116021,I116004);
nor I_6656 (I115583,I115860,I116021);
nand I_6657 (I115568,I115877,I116021);
nor I_6658 (I115577,I115623,I116004);
DFFARX1 I_6659 (I116004,I2859,I115597,I115586,);
not I_6660 (I116124,I2866);
DFFARX1 I_6661 (I483000,I2859,I116124,I116150,);
nand I_6662 (I116158,I483015,I483000);
and I_6663 (I116175,I116158,I483018);
DFFARX1 I_6664 (I116175,I2859,I116124,I116201,);
nor I_6665 (I116092,I116201,I116150);
not I_6666 (I116223,I116201);
DFFARX1 I_6667 (I483024,I2859,I116124,I116249,);
nand I_6668 (I116257,I116249,I483006);
not I_6669 (I116274,I116257);
DFFARX1 I_6670 (I116274,I2859,I116124,I116300,);
not I_6671 (I116116,I116300);
nor I_6672 (I116322,I116150,I116257);
nor I_6673 (I116098,I116201,I116322);
DFFARX1 I_6674 (I483003,I2859,I116124,I116362,);
DFFARX1 I_6675 (I116362,I2859,I116124,I116379,);
not I_6676 (I116387,I116379);
not I_6677 (I116404,I116362);
nand I_6678 (I116101,I116404,I116223);
nand I_6679 (I116435,I483003,I483009);
and I_6680 (I116452,I116435,I483021);
DFFARX1 I_6681 (I116452,I2859,I116124,I116478,);
nor I_6682 (I116486,I116478,I116150);
DFFARX1 I_6683 (I116486,I2859,I116124,I116089,);
DFFARX1 I_6684 (I116478,I2859,I116124,I116107,);
nor I_6685 (I116531,I483012,I483009);
not I_6686 (I116548,I116531);
nor I_6687 (I116110,I116387,I116548);
nand I_6688 (I116095,I116404,I116548);
nor I_6689 (I116104,I116150,I116531);
DFFARX1 I_6690 (I116531,I2859,I116124,I116113,);
not I_6691 (I116651,I2866);
DFFARX1 I_6692 (I314746,I2859,I116651,I116677,);
nand I_6693 (I116685,I314737,I314752);
and I_6694 (I116702,I116685,I314758);
DFFARX1 I_6695 (I116702,I2859,I116651,I116728,);
nor I_6696 (I116619,I116728,I116677);
not I_6697 (I116750,I116728);
DFFARX1 I_6698 (I314743,I2859,I116651,I116776,);
nand I_6699 (I116784,I116776,I314737);
not I_6700 (I116801,I116784);
DFFARX1 I_6701 (I116801,I2859,I116651,I116827,);
not I_6702 (I116643,I116827);
nor I_6703 (I116849,I116677,I116784);
nor I_6704 (I116625,I116728,I116849);
DFFARX1 I_6705 (I314740,I2859,I116651,I116889,);
DFFARX1 I_6706 (I116889,I2859,I116651,I116906,);
not I_6707 (I116914,I116906);
not I_6708 (I116931,I116889);
nand I_6709 (I116628,I116931,I116750);
nand I_6710 (I116962,I314734,I314749);
and I_6711 (I116979,I116962,I314734);
DFFARX1 I_6712 (I116979,I2859,I116651,I117005,);
nor I_6713 (I117013,I117005,I116677);
DFFARX1 I_6714 (I117013,I2859,I116651,I116616,);
DFFARX1 I_6715 (I117005,I2859,I116651,I116634,);
nor I_6716 (I117058,I314755,I314749);
not I_6717 (I117075,I117058);
nor I_6718 (I116637,I116914,I117075);
nand I_6719 (I116622,I116931,I117075);
nor I_6720 (I116631,I116677,I117058);
DFFARX1 I_6721 (I117058,I2859,I116651,I116640,);
not I_6722 (I117178,I2866);
DFFARX1 I_6723 (I56830,I2859,I117178,I117204,);
nand I_6724 (I117212,I56842,I56851);
and I_6725 (I117229,I117212,I56830);
DFFARX1 I_6726 (I117229,I2859,I117178,I117255,);
nor I_6727 (I117146,I117255,I117204);
not I_6728 (I117277,I117255);
DFFARX1 I_6729 (I56845,I2859,I117178,I117303,);
nand I_6730 (I117311,I117303,I56833);
not I_6731 (I117328,I117311);
DFFARX1 I_6732 (I117328,I2859,I117178,I117354,);
not I_6733 (I117170,I117354);
nor I_6734 (I117376,I117204,I117311);
nor I_6735 (I117152,I117255,I117376);
DFFARX1 I_6736 (I56836,I2859,I117178,I117416,);
DFFARX1 I_6737 (I117416,I2859,I117178,I117433,);
not I_6738 (I117441,I117433);
not I_6739 (I117458,I117416);
nand I_6740 (I117155,I117458,I117277);
nand I_6741 (I117489,I56827,I56827);
and I_6742 (I117506,I117489,I56839);
DFFARX1 I_6743 (I117506,I2859,I117178,I117532,);
nor I_6744 (I117540,I117532,I117204);
DFFARX1 I_6745 (I117540,I2859,I117178,I117143,);
DFFARX1 I_6746 (I117532,I2859,I117178,I117161,);
nor I_6747 (I117585,I56848,I56827);
not I_6748 (I117602,I117585);
nor I_6749 (I117164,I117441,I117602);
nand I_6750 (I117149,I117458,I117602);
nor I_6751 (I117158,I117204,I117585);
DFFARX1 I_6752 (I117585,I2859,I117178,I117167,);
not I_6753 (I117705,I2866);
DFFARX1 I_6754 (I474330,I2859,I117705,I117731,);
nand I_6755 (I117739,I474345,I474330);
and I_6756 (I117756,I117739,I474348);
DFFARX1 I_6757 (I117756,I2859,I117705,I117782,);
nor I_6758 (I117673,I117782,I117731);
not I_6759 (I117804,I117782);
DFFARX1 I_6760 (I474354,I2859,I117705,I117830,);
nand I_6761 (I117838,I117830,I474336);
not I_6762 (I117855,I117838);
DFFARX1 I_6763 (I117855,I2859,I117705,I117881,);
not I_6764 (I117697,I117881);
nor I_6765 (I117903,I117731,I117838);
nor I_6766 (I117679,I117782,I117903);
DFFARX1 I_6767 (I474333,I2859,I117705,I117943,);
DFFARX1 I_6768 (I117943,I2859,I117705,I117960,);
not I_6769 (I117968,I117960);
not I_6770 (I117985,I117943);
nand I_6771 (I117682,I117985,I117804);
nand I_6772 (I118016,I474333,I474339);
and I_6773 (I118033,I118016,I474351);
DFFARX1 I_6774 (I118033,I2859,I117705,I118059,);
nor I_6775 (I118067,I118059,I117731);
DFFARX1 I_6776 (I118067,I2859,I117705,I117670,);
DFFARX1 I_6777 (I118059,I2859,I117705,I117688,);
nor I_6778 (I118112,I474342,I474339);
not I_6779 (I118129,I118112);
nor I_6780 (I117691,I117968,I118129);
nand I_6781 (I117676,I117985,I118129);
nor I_6782 (I117685,I117731,I118112);
DFFARX1 I_6783 (I118112,I2859,I117705,I117694,);
not I_6784 (I118232,I2866);
DFFARX1 I_6785 (I360586,I2859,I118232,I118258,);
nand I_6786 (I118266,I360589,I360583);
and I_6787 (I118283,I118266,I360595);
DFFARX1 I_6788 (I118283,I2859,I118232,I118309,);
nor I_6789 (I118200,I118309,I118258);
not I_6790 (I118331,I118309);
DFFARX1 I_6791 (I360598,I2859,I118232,I118357,);
nand I_6792 (I118365,I118357,I360589);
not I_6793 (I118382,I118365);
DFFARX1 I_6794 (I118382,I2859,I118232,I118408,);
not I_6795 (I118224,I118408);
nor I_6796 (I118430,I118258,I118365);
nor I_6797 (I118206,I118309,I118430);
DFFARX1 I_6798 (I360601,I2859,I118232,I118470,);
DFFARX1 I_6799 (I118470,I2859,I118232,I118487,);
not I_6800 (I118495,I118487);
not I_6801 (I118512,I118470);
nand I_6802 (I118209,I118512,I118331);
nand I_6803 (I118543,I360583,I360592);
and I_6804 (I118560,I118543,I360586);
DFFARX1 I_6805 (I118560,I2859,I118232,I118586,);
nor I_6806 (I118594,I118586,I118258);
DFFARX1 I_6807 (I118594,I2859,I118232,I118197,);
DFFARX1 I_6808 (I118586,I2859,I118232,I118215,);
nor I_6809 (I118639,I360604,I360592);
not I_6810 (I118656,I118639);
nor I_6811 (I118218,I118495,I118656);
nand I_6812 (I118203,I118512,I118656);
nor I_6813 (I118212,I118258,I118639);
DFFARX1 I_6814 (I118639,I2859,I118232,I118221,);
not I_6815 (I118759,I2866);
DFFARX1 I_6816 (I533845,I2859,I118759,I118785,);
nand I_6817 (I118793,I533842,I533833);
and I_6818 (I118810,I118793,I533830);
DFFARX1 I_6819 (I118810,I2859,I118759,I118836,);
nor I_6820 (I118727,I118836,I118785);
not I_6821 (I118858,I118836);
DFFARX1 I_6822 (I533839,I2859,I118759,I118884,);
nand I_6823 (I118892,I118884,I533848);
not I_6824 (I118909,I118892);
DFFARX1 I_6825 (I118909,I2859,I118759,I118935,);
not I_6826 (I118751,I118935);
nor I_6827 (I118957,I118785,I118892);
nor I_6828 (I118733,I118836,I118957);
DFFARX1 I_6829 (I533851,I2859,I118759,I118997,);
DFFARX1 I_6830 (I118997,I2859,I118759,I119014,);
not I_6831 (I119022,I119014);
not I_6832 (I119039,I118997);
nand I_6833 (I118736,I119039,I118858);
nand I_6834 (I119070,I533830,I533836);
and I_6835 (I119087,I119070,I533854);
DFFARX1 I_6836 (I119087,I2859,I118759,I119113,);
nor I_6837 (I119121,I119113,I118785);
DFFARX1 I_6838 (I119121,I2859,I118759,I118724,);
DFFARX1 I_6839 (I119113,I2859,I118759,I118742,);
nor I_6840 (I119166,I533833,I533836);
not I_6841 (I119183,I119166);
nor I_6842 (I118745,I119022,I119183);
nand I_6843 (I118730,I119039,I119183);
nor I_6844 (I118739,I118785,I119166);
DFFARX1 I_6845 (I119166,I2859,I118759,I118748,);
not I_6846 (I119286,I2866);
DFFARX1 I_6847 (I42601,I2859,I119286,I119312,);
nand I_6848 (I119320,I42613,I42622);
and I_6849 (I119337,I119320,I42601);
DFFARX1 I_6850 (I119337,I2859,I119286,I119363,);
nor I_6851 (I119254,I119363,I119312);
not I_6852 (I119385,I119363);
DFFARX1 I_6853 (I42616,I2859,I119286,I119411,);
nand I_6854 (I119419,I119411,I42604);
not I_6855 (I119436,I119419);
DFFARX1 I_6856 (I119436,I2859,I119286,I119462,);
not I_6857 (I119278,I119462);
nor I_6858 (I119484,I119312,I119419);
nor I_6859 (I119260,I119363,I119484);
DFFARX1 I_6860 (I42607,I2859,I119286,I119524,);
DFFARX1 I_6861 (I119524,I2859,I119286,I119541,);
not I_6862 (I119549,I119541);
not I_6863 (I119566,I119524);
nand I_6864 (I119263,I119566,I119385);
nand I_6865 (I119597,I42598,I42598);
and I_6866 (I119614,I119597,I42610);
DFFARX1 I_6867 (I119614,I2859,I119286,I119640,);
nor I_6868 (I119648,I119640,I119312);
DFFARX1 I_6869 (I119648,I2859,I119286,I119251,);
DFFARX1 I_6870 (I119640,I2859,I119286,I119269,);
nor I_6871 (I119693,I42619,I42598);
not I_6872 (I119710,I119693);
nor I_6873 (I119272,I119549,I119710);
nand I_6874 (I119257,I119566,I119710);
nor I_6875 (I119266,I119312,I119693);
DFFARX1 I_6876 (I119693,I2859,I119286,I119275,);
not I_6877 (I119813,I2866);
DFFARX1 I_6878 (I493982,I2859,I119813,I119839,);
nand I_6879 (I119847,I493997,I493982);
and I_6880 (I119864,I119847,I494000);
DFFARX1 I_6881 (I119864,I2859,I119813,I119890,);
nor I_6882 (I119781,I119890,I119839);
not I_6883 (I119912,I119890);
DFFARX1 I_6884 (I494006,I2859,I119813,I119938,);
nand I_6885 (I119946,I119938,I493988);
not I_6886 (I119963,I119946);
DFFARX1 I_6887 (I119963,I2859,I119813,I119989,);
not I_6888 (I119805,I119989);
nor I_6889 (I120011,I119839,I119946);
nor I_6890 (I119787,I119890,I120011);
DFFARX1 I_6891 (I493985,I2859,I119813,I120051,);
DFFARX1 I_6892 (I120051,I2859,I119813,I120068,);
not I_6893 (I120076,I120068);
not I_6894 (I120093,I120051);
nand I_6895 (I119790,I120093,I119912);
nand I_6896 (I120124,I493985,I493991);
and I_6897 (I120141,I120124,I494003);
DFFARX1 I_6898 (I120141,I2859,I119813,I120167,);
nor I_6899 (I120175,I120167,I119839);
DFFARX1 I_6900 (I120175,I2859,I119813,I119778,);
DFFARX1 I_6901 (I120167,I2859,I119813,I119796,);
nor I_6902 (I120220,I493994,I493991);
not I_6903 (I120237,I120220);
nor I_6904 (I119799,I120076,I120237);
nand I_6905 (I119784,I120093,I120237);
nor I_6906 (I119793,I119839,I120220);
DFFARX1 I_6907 (I120220,I2859,I119813,I119802,);
not I_6908 (I120340,I2866);
DFFARX1 I_6909 (I229783,I2859,I120340,I120366,);
nand I_6910 (I120374,I229768,I229771);
and I_6911 (I120391,I120374,I229786);
DFFARX1 I_6912 (I120391,I2859,I120340,I120417,);
nor I_6913 (I120308,I120417,I120366);
not I_6914 (I120439,I120417);
DFFARX1 I_6915 (I229780,I2859,I120340,I120465,);
nand I_6916 (I120473,I120465,I229771);
not I_6917 (I120490,I120473);
DFFARX1 I_6918 (I120490,I2859,I120340,I120516,);
not I_6919 (I120332,I120516);
nor I_6920 (I120538,I120366,I120473);
nor I_6921 (I120314,I120417,I120538);
DFFARX1 I_6922 (I229777,I2859,I120340,I120578,);
DFFARX1 I_6923 (I120578,I2859,I120340,I120595,);
not I_6924 (I120603,I120595);
not I_6925 (I120620,I120578);
nand I_6926 (I120317,I120620,I120439);
nand I_6927 (I120651,I229792,I229768);
and I_6928 (I120668,I120651,I229789);
DFFARX1 I_6929 (I120668,I2859,I120340,I120694,);
nor I_6930 (I120702,I120694,I120366);
DFFARX1 I_6931 (I120702,I2859,I120340,I120305,);
DFFARX1 I_6932 (I120694,I2859,I120340,I120323,);
nor I_6933 (I120747,I229774,I229768);
not I_6934 (I120764,I120747);
nor I_6935 (I120326,I120603,I120764);
nand I_6936 (I120311,I120620,I120764);
nor I_6937 (I120320,I120366,I120747);
DFFARX1 I_6938 (I120747,I2859,I120340,I120329,);
not I_6939 (I120867,I2866);
DFFARX1 I_6940 (I350046,I2859,I120867,I120893,);
nand I_6941 (I120901,I350049,I350043);
and I_6942 (I120918,I120901,I350055);
DFFARX1 I_6943 (I120918,I2859,I120867,I120944,);
nor I_6944 (I120835,I120944,I120893);
not I_6945 (I120966,I120944);
DFFARX1 I_6946 (I350058,I2859,I120867,I120992,);
nand I_6947 (I121000,I120992,I350049);
not I_6948 (I121017,I121000);
DFFARX1 I_6949 (I121017,I2859,I120867,I121043,);
not I_6950 (I120859,I121043);
nor I_6951 (I121065,I120893,I121000);
nor I_6952 (I120841,I120944,I121065);
DFFARX1 I_6953 (I350061,I2859,I120867,I121105,);
DFFARX1 I_6954 (I121105,I2859,I120867,I121122,);
not I_6955 (I121130,I121122);
not I_6956 (I121147,I121105);
nand I_6957 (I120844,I121147,I120966);
nand I_6958 (I121178,I350043,I350052);
and I_6959 (I121195,I121178,I350046);
DFFARX1 I_6960 (I121195,I2859,I120867,I121221,);
nor I_6961 (I121229,I121221,I120893);
DFFARX1 I_6962 (I121229,I2859,I120867,I120832,);
DFFARX1 I_6963 (I121221,I2859,I120867,I120850,);
nor I_6964 (I121274,I350064,I350052);
not I_6965 (I121291,I121274);
nor I_6966 (I120853,I121130,I121291);
nand I_6967 (I120838,I121147,I121291);
nor I_6968 (I120847,I120893,I121274);
DFFARX1 I_6969 (I121274,I2859,I120867,I120856,);
not I_6970 (I121394,I2866);
DFFARX1 I_6971 (I562156,I2859,I121394,I121420,);
nand I_6972 (I121428,I562135,I562135);
and I_6973 (I121445,I121428,I562162);
DFFARX1 I_6974 (I121445,I2859,I121394,I121471,);
nor I_6975 (I121362,I121471,I121420);
not I_6976 (I121493,I121471);
DFFARX1 I_6977 (I562150,I2859,I121394,I121519,);
nand I_6978 (I121527,I121519,I562153);
not I_6979 (I121544,I121527);
DFFARX1 I_6980 (I121544,I2859,I121394,I121570,);
not I_6981 (I121386,I121570);
nor I_6982 (I121592,I121420,I121527);
nor I_6983 (I121368,I121471,I121592);
DFFARX1 I_6984 (I562144,I2859,I121394,I121632,);
DFFARX1 I_6985 (I121632,I2859,I121394,I121649,);
not I_6986 (I121657,I121649);
not I_6987 (I121674,I121632);
nand I_6988 (I121371,I121674,I121493);
nand I_6989 (I121705,I562141,I562138);
and I_6990 (I121722,I121705,I562159);
DFFARX1 I_6991 (I121722,I2859,I121394,I121748,);
nor I_6992 (I121756,I121748,I121420);
DFFARX1 I_6993 (I121756,I2859,I121394,I121359,);
DFFARX1 I_6994 (I121748,I2859,I121394,I121377,);
nor I_6995 (I121801,I562147,I562138);
not I_6996 (I121818,I121801);
nor I_6997 (I121380,I121657,I121818);
nand I_6998 (I121365,I121674,I121818);
nor I_6999 (I121374,I121420,I121801);
DFFARX1 I_7000 (I121801,I2859,I121394,I121383,);
not I_7001 (I121921,I2866);
DFFARX1 I_7002 (I23629,I2859,I121921,I121947,);
nand I_7003 (I121955,I23641,I23650);
and I_7004 (I121972,I121955,I23629);
DFFARX1 I_7005 (I121972,I2859,I121921,I121998,);
nor I_7006 (I121889,I121998,I121947);
not I_7007 (I122020,I121998);
DFFARX1 I_7008 (I23644,I2859,I121921,I122046,);
nand I_7009 (I122054,I122046,I23632);
not I_7010 (I122071,I122054);
DFFARX1 I_7011 (I122071,I2859,I121921,I122097,);
not I_7012 (I121913,I122097);
nor I_7013 (I122119,I121947,I122054);
nor I_7014 (I121895,I121998,I122119);
DFFARX1 I_7015 (I23635,I2859,I121921,I122159,);
DFFARX1 I_7016 (I122159,I2859,I121921,I122176,);
not I_7017 (I122184,I122176);
not I_7018 (I122201,I122159);
nand I_7019 (I121898,I122201,I122020);
nand I_7020 (I122232,I23626,I23626);
and I_7021 (I122249,I122232,I23638);
DFFARX1 I_7022 (I122249,I2859,I121921,I122275,);
nor I_7023 (I122283,I122275,I121947);
DFFARX1 I_7024 (I122283,I2859,I121921,I121886,);
DFFARX1 I_7025 (I122275,I2859,I121921,I121904,);
nor I_7026 (I122328,I23647,I23626);
not I_7027 (I122345,I122328);
nor I_7028 (I121907,I122184,I122345);
nand I_7029 (I121892,I122201,I122345);
nor I_7030 (I121901,I121947,I122328);
DFFARX1 I_7031 (I122328,I2859,I121921,I121910,);
not I_7032 (I122448,I2866);
DFFARX1 I_7033 (I338979,I2859,I122448,I122474,);
nand I_7034 (I122482,I338982,I338976);
and I_7035 (I122499,I122482,I338988);
DFFARX1 I_7036 (I122499,I2859,I122448,I122525,);
nor I_7037 (I122416,I122525,I122474);
not I_7038 (I122547,I122525);
DFFARX1 I_7039 (I338991,I2859,I122448,I122573,);
nand I_7040 (I122581,I122573,I338982);
not I_7041 (I122598,I122581);
DFFARX1 I_7042 (I122598,I2859,I122448,I122624,);
not I_7043 (I122440,I122624);
nor I_7044 (I122646,I122474,I122581);
nor I_7045 (I122422,I122525,I122646);
DFFARX1 I_7046 (I338994,I2859,I122448,I122686,);
DFFARX1 I_7047 (I122686,I2859,I122448,I122703,);
not I_7048 (I122711,I122703);
not I_7049 (I122728,I122686);
nand I_7050 (I122425,I122728,I122547);
nand I_7051 (I122759,I338976,I338985);
and I_7052 (I122776,I122759,I338979);
DFFARX1 I_7053 (I122776,I2859,I122448,I122802,);
nor I_7054 (I122810,I122802,I122474);
DFFARX1 I_7055 (I122810,I2859,I122448,I122413,);
DFFARX1 I_7056 (I122802,I2859,I122448,I122431,);
nor I_7057 (I122855,I338997,I338985);
not I_7058 (I122872,I122855);
nor I_7059 (I122434,I122711,I122872);
nand I_7060 (I122419,I122728,I122872);
nor I_7061 (I122428,I122474,I122855);
DFFARX1 I_7062 (I122855,I2859,I122448,I122437,);
not I_7063 (I122975,I2866);
DFFARX1 I_7064 (I247701,I2859,I122975,I123001,);
nand I_7065 (I123009,I247686,I247689);
and I_7066 (I123026,I123009,I247704);
DFFARX1 I_7067 (I123026,I2859,I122975,I123052,);
nor I_7068 (I122943,I123052,I123001);
not I_7069 (I123074,I123052);
DFFARX1 I_7070 (I247698,I2859,I122975,I123100,);
nand I_7071 (I123108,I123100,I247689);
not I_7072 (I123125,I123108);
DFFARX1 I_7073 (I123125,I2859,I122975,I123151,);
not I_7074 (I122967,I123151);
nor I_7075 (I123173,I123001,I123108);
nor I_7076 (I122949,I123052,I123173);
DFFARX1 I_7077 (I247695,I2859,I122975,I123213,);
DFFARX1 I_7078 (I123213,I2859,I122975,I123230,);
not I_7079 (I123238,I123230);
not I_7080 (I123255,I123213);
nand I_7081 (I122952,I123255,I123074);
nand I_7082 (I123286,I247710,I247686);
and I_7083 (I123303,I123286,I247707);
DFFARX1 I_7084 (I123303,I2859,I122975,I123329,);
nor I_7085 (I123337,I123329,I123001);
DFFARX1 I_7086 (I123337,I2859,I122975,I122940,);
DFFARX1 I_7087 (I123329,I2859,I122975,I122958,);
nor I_7088 (I123382,I247692,I247686);
not I_7089 (I123399,I123382);
nor I_7090 (I122961,I123238,I123399);
nand I_7091 (I122946,I123255,I123399);
nor I_7092 (I122955,I123001,I123382);
DFFARX1 I_7093 (I123382,I2859,I122975,I122964,);
not I_7094 (I123502,I2866);
DFFARX1 I_7095 (I543711,I2859,I123502,I123528,);
nand I_7096 (I123536,I543690,I543690);
and I_7097 (I123553,I123536,I543717);
DFFARX1 I_7098 (I123553,I2859,I123502,I123579,);
nor I_7099 (I123470,I123579,I123528);
not I_7100 (I123601,I123579);
DFFARX1 I_7101 (I543705,I2859,I123502,I123627,);
nand I_7102 (I123635,I123627,I543708);
not I_7103 (I123652,I123635);
DFFARX1 I_7104 (I123652,I2859,I123502,I123678,);
not I_7105 (I123494,I123678);
nor I_7106 (I123700,I123528,I123635);
nor I_7107 (I123476,I123579,I123700);
DFFARX1 I_7108 (I543699,I2859,I123502,I123740,);
DFFARX1 I_7109 (I123740,I2859,I123502,I123757,);
not I_7110 (I123765,I123757);
not I_7111 (I123782,I123740);
nand I_7112 (I123479,I123782,I123601);
nand I_7113 (I123813,I543696,I543693);
and I_7114 (I123830,I123813,I543714);
DFFARX1 I_7115 (I123830,I2859,I123502,I123856,);
nor I_7116 (I123864,I123856,I123528);
DFFARX1 I_7117 (I123864,I2859,I123502,I123467,);
DFFARX1 I_7118 (I123856,I2859,I123502,I123485,);
nor I_7119 (I123909,I543702,I543693);
not I_7120 (I123926,I123909);
nor I_7121 (I123488,I123765,I123926);
nand I_7122 (I123473,I123782,I123926);
nor I_7123 (I123482,I123528,I123909);
DFFARX1 I_7124 (I123909,I2859,I123502,I123491,);
not I_7125 (I124029,I2866);
DFFARX1 I_7126 (I535001,I2859,I124029,I124055,);
nand I_7127 (I124063,I534998,I534989);
and I_7128 (I124080,I124063,I534986);
DFFARX1 I_7129 (I124080,I2859,I124029,I124106,);
nor I_7130 (I123997,I124106,I124055);
not I_7131 (I124128,I124106);
DFFARX1 I_7132 (I534995,I2859,I124029,I124154,);
nand I_7133 (I124162,I124154,I535004);
not I_7134 (I124179,I124162);
DFFARX1 I_7135 (I124179,I2859,I124029,I124205,);
not I_7136 (I124021,I124205);
nor I_7137 (I124227,I124055,I124162);
nor I_7138 (I124003,I124106,I124227);
DFFARX1 I_7139 (I535007,I2859,I124029,I124267,);
DFFARX1 I_7140 (I124267,I2859,I124029,I124284,);
not I_7141 (I124292,I124284);
not I_7142 (I124309,I124267);
nand I_7143 (I124006,I124309,I124128);
nand I_7144 (I124340,I534986,I534992);
and I_7145 (I124357,I124340,I535010);
DFFARX1 I_7146 (I124357,I2859,I124029,I124383,);
nor I_7147 (I124391,I124383,I124055);
DFFARX1 I_7148 (I124391,I2859,I124029,I123994,);
DFFARX1 I_7149 (I124383,I2859,I124029,I124012,);
nor I_7150 (I124436,I534989,I534992);
not I_7151 (I124453,I124436);
nor I_7152 (I124015,I124292,I124453);
nand I_7153 (I124000,I124309,I124453);
nor I_7154 (I124009,I124055,I124436);
DFFARX1 I_7155 (I124436,I2859,I124029,I124018,);
not I_7156 (I124556,I2866);
DFFARX1 I_7157 (I338452,I2859,I124556,I124582,);
nand I_7158 (I124590,I338455,I338449);
and I_7159 (I124607,I124590,I338461);
DFFARX1 I_7160 (I124607,I2859,I124556,I124633,);
nor I_7161 (I124524,I124633,I124582);
not I_7162 (I124655,I124633);
DFFARX1 I_7163 (I338464,I2859,I124556,I124681,);
nand I_7164 (I124689,I124681,I338455);
not I_7165 (I124706,I124689);
DFFARX1 I_7166 (I124706,I2859,I124556,I124732,);
not I_7167 (I124548,I124732);
nor I_7168 (I124754,I124582,I124689);
nor I_7169 (I124530,I124633,I124754);
DFFARX1 I_7170 (I338467,I2859,I124556,I124794,);
DFFARX1 I_7171 (I124794,I2859,I124556,I124811,);
not I_7172 (I124819,I124811);
not I_7173 (I124836,I124794);
nand I_7174 (I124533,I124836,I124655);
nand I_7175 (I124867,I338449,I338458);
and I_7176 (I124884,I124867,I338452);
DFFARX1 I_7177 (I124884,I2859,I124556,I124910,);
nor I_7178 (I124918,I124910,I124582);
DFFARX1 I_7179 (I124918,I2859,I124556,I124521,);
DFFARX1 I_7180 (I124910,I2859,I124556,I124539,);
nor I_7181 (I124963,I338470,I338458);
not I_7182 (I124980,I124963);
nor I_7183 (I124542,I124819,I124980);
nand I_7184 (I124527,I124836,I124980);
nor I_7185 (I124536,I124582,I124963);
DFFARX1 I_7186 (I124963,I2859,I124556,I124545,);
not I_7187 (I125083,I2866);
DFFARX1 I_7188 (I444396,I2859,I125083,I125109,);
nand I_7189 (I125117,I444393,I444396);
and I_7190 (I125134,I125117,I444405);
DFFARX1 I_7191 (I125134,I2859,I125083,I125160,);
nor I_7192 (I125051,I125160,I125109);
not I_7193 (I125182,I125160);
DFFARX1 I_7194 (I444393,I2859,I125083,I125208,);
nand I_7195 (I125216,I125208,I444411);
not I_7196 (I125233,I125216);
DFFARX1 I_7197 (I125233,I2859,I125083,I125259,);
not I_7198 (I125075,I125259);
nor I_7199 (I125281,I125109,I125216);
nor I_7200 (I125057,I125160,I125281);
DFFARX1 I_7201 (I444399,I2859,I125083,I125321,);
DFFARX1 I_7202 (I125321,I2859,I125083,I125338,);
not I_7203 (I125346,I125338);
not I_7204 (I125363,I125321);
nand I_7205 (I125060,I125363,I125182);
nand I_7206 (I125394,I444408,I444414);
and I_7207 (I125411,I125394,I444399);
DFFARX1 I_7208 (I125411,I2859,I125083,I125437,);
nor I_7209 (I125445,I125437,I125109);
DFFARX1 I_7210 (I125445,I2859,I125083,I125048,);
DFFARX1 I_7211 (I125437,I2859,I125083,I125066,);
nor I_7212 (I125490,I444402,I444414);
not I_7213 (I125507,I125490);
nor I_7214 (I125069,I125346,I125507);
nand I_7215 (I125054,I125363,I125507);
nor I_7216 (I125063,I125109,I125490);
DFFARX1 I_7217 (I125490,I2859,I125083,I125072,);
not I_7218 (I125610,I2866);
DFFARX1 I_7219 (I510796,I2859,I125610,I125636,);
nand I_7220 (I125644,I510778,I510802);
and I_7221 (I125661,I125644,I510793);
DFFARX1 I_7222 (I125661,I2859,I125610,I125687,);
nor I_7223 (I125578,I125687,I125636);
not I_7224 (I125709,I125687);
DFFARX1 I_7225 (I510799,I2859,I125610,I125735,);
nand I_7226 (I125743,I125735,I510787);
not I_7227 (I125760,I125743);
DFFARX1 I_7228 (I125760,I2859,I125610,I125786,);
not I_7229 (I125602,I125786);
nor I_7230 (I125808,I125636,I125743);
nor I_7231 (I125584,I125687,I125808);
DFFARX1 I_7232 (I510778,I2859,I125610,I125848,);
DFFARX1 I_7233 (I125848,I2859,I125610,I125865,);
not I_7234 (I125873,I125865);
not I_7235 (I125890,I125848);
nand I_7236 (I125587,I125890,I125709);
nand I_7237 (I125921,I510784,I510781);
and I_7238 (I125938,I125921,I510790);
DFFARX1 I_7239 (I125938,I2859,I125610,I125964,);
nor I_7240 (I125972,I125964,I125636);
DFFARX1 I_7241 (I125972,I2859,I125610,I125575,);
DFFARX1 I_7242 (I125964,I2859,I125610,I125593,);
nor I_7243 (I126017,I510781,I510781);
not I_7244 (I126034,I126017);
nor I_7245 (I125596,I125873,I126034);
nand I_7246 (I125581,I125890,I126034);
nor I_7247 (I125590,I125636,I126017);
DFFARX1 I_7248 (I126017,I2859,I125610,I125599,);
not I_7249 (I126137,I2866);
DFFARX1 I_7250 (I168903,I2859,I126137,I126163,);
nand I_7251 (I126171,I168915,I168894);
and I_7252 (I126188,I126171,I168918);
DFFARX1 I_7253 (I126188,I2859,I126137,I126214,);
nor I_7254 (I126105,I126214,I126163);
not I_7255 (I126236,I126214);
DFFARX1 I_7256 (I168909,I2859,I126137,I126262,);
nand I_7257 (I126270,I126262,I168891);
not I_7258 (I126287,I126270);
DFFARX1 I_7259 (I126287,I2859,I126137,I126313,);
not I_7260 (I126129,I126313);
nor I_7261 (I126335,I126163,I126270);
nor I_7262 (I126111,I126214,I126335);
DFFARX1 I_7263 (I168906,I2859,I126137,I126375,);
DFFARX1 I_7264 (I126375,I2859,I126137,I126392,);
not I_7265 (I126400,I126392);
not I_7266 (I126417,I126375);
nand I_7267 (I126114,I126417,I126236);
nand I_7268 (I126448,I168891,I168897);
and I_7269 (I126465,I126448,I168900);
DFFARX1 I_7270 (I126465,I2859,I126137,I126491,);
nor I_7271 (I126499,I126491,I126163);
DFFARX1 I_7272 (I126499,I2859,I126137,I126102,);
DFFARX1 I_7273 (I126491,I2859,I126137,I126120,);
nor I_7274 (I126544,I168912,I168897);
not I_7275 (I126561,I126544);
nor I_7276 (I126123,I126400,I126561);
nand I_7277 (I126108,I126417,I126561);
nor I_7278 (I126117,I126163,I126544);
DFFARX1 I_7279 (I126544,I2859,I126137,I126126,);
not I_7280 (I126664,I2866);
DFFARX1 I_7281 (I537247,I2859,I126664,I126690,);
nand I_7282 (I126698,I537274,I537250);
and I_7283 (I126715,I126698,I537259);
DFFARX1 I_7284 (I126715,I2859,I126664,I126741,);
nor I_7285 (I126632,I126741,I126690);
not I_7286 (I126763,I126741);
DFFARX1 I_7287 (I537247,I2859,I126664,I126789,);
nand I_7288 (I126797,I126789,I537271);
not I_7289 (I126814,I126797);
DFFARX1 I_7290 (I126814,I2859,I126664,I126840,);
not I_7291 (I126656,I126840);
nor I_7292 (I126862,I126690,I126797);
nor I_7293 (I126638,I126741,I126862);
DFFARX1 I_7294 (I537253,I2859,I126664,I126902,);
DFFARX1 I_7295 (I126902,I2859,I126664,I126919,);
not I_7296 (I126927,I126919);
not I_7297 (I126944,I126902);
nand I_7298 (I126641,I126944,I126763);
nand I_7299 (I126975,I537268,I537256);
and I_7300 (I126992,I126975,I537262);
DFFARX1 I_7301 (I126992,I2859,I126664,I127018,);
nor I_7302 (I127026,I127018,I126690);
DFFARX1 I_7303 (I127026,I2859,I126664,I126629,);
DFFARX1 I_7304 (I127018,I2859,I126664,I126647,);
nor I_7305 (I127071,I537265,I537256);
not I_7306 (I127088,I127071);
nor I_7307 (I126650,I126927,I127088);
nand I_7308 (I126635,I126944,I127088);
nor I_7309 (I126644,I126690,I127071);
DFFARX1 I_7310 (I127071,I2859,I126664,I126653,);
not I_7311 (I127191,I2866);
DFFARX1 I_7312 (I274864,I2859,I127191,I127217,);
nand I_7313 (I127225,I274855,I274870);
and I_7314 (I127242,I127225,I274876);
DFFARX1 I_7315 (I127242,I2859,I127191,I127268,);
nor I_7316 (I127159,I127268,I127217);
not I_7317 (I127290,I127268);
DFFARX1 I_7318 (I274861,I2859,I127191,I127316,);
nand I_7319 (I127324,I127316,I274855);
not I_7320 (I127341,I127324);
DFFARX1 I_7321 (I127341,I2859,I127191,I127367,);
not I_7322 (I127183,I127367);
nor I_7323 (I127389,I127217,I127324);
nor I_7324 (I127165,I127268,I127389);
DFFARX1 I_7325 (I274858,I2859,I127191,I127429,);
DFFARX1 I_7326 (I127429,I2859,I127191,I127446,);
not I_7327 (I127454,I127446);
not I_7328 (I127471,I127429);
nand I_7329 (I127168,I127471,I127290);
nand I_7330 (I127502,I274852,I274867);
and I_7331 (I127519,I127502,I274852);
DFFARX1 I_7332 (I127519,I2859,I127191,I127545,);
nor I_7333 (I127553,I127545,I127217);
DFFARX1 I_7334 (I127553,I2859,I127191,I127156,);
DFFARX1 I_7335 (I127545,I2859,I127191,I127174,);
nor I_7336 (I127598,I274873,I274867);
not I_7337 (I127615,I127598);
nor I_7338 (I127177,I127454,I127615);
nand I_7339 (I127162,I127471,I127615);
nor I_7340 (I127171,I127217,I127598);
DFFARX1 I_7341 (I127598,I2859,I127191,I127180,);
not I_7342 (I127718,I2866);
DFFARX1 I_7343 (I388024,I2859,I127718,I127744,);
nand I_7344 (I127752,I388021,I388039);
and I_7345 (I127769,I127752,I388030);
DFFARX1 I_7346 (I127769,I2859,I127718,I127795,);
nor I_7347 (I127686,I127795,I127744);
not I_7348 (I127817,I127795);
DFFARX1 I_7349 (I388045,I2859,I127718,I127843,);
nand I_7350 (I127851,I127843,I388027);
not I_7351 (I127868,I127851);
DFFARX1 I_7352 (I127868,I2859,I127718,I127894,);
not I_7353 (I127710,I127894);
nor I_7354 (I127916,I127744,I127851);
nor I_7355 (I127692,I127795,I127916);
DFFARX1 I_7356 (I388033,I2859,I127718,I127956,);
DFFARX1 I_7357 (I127956,I2859,I127718,I127973,);
not I_7358 (I127981,I127973);
not I_7359 (I127998,I127956);
nand I_7360 (I127695,I127998,I127817);
nand I_7361 (I128029,I388021,I388048);
and I_7362 (I128046,I128029,I388036);
DFFARX1 I_7363 (I128046,I2859,I127718,I128072,);
nor I_7364 (I128080,I128072,I127744);
DFFARX1 I_7365 (I128080,I2859,I127718,I127683,);
DFFARX1 I_7366 (I128072,I2859,I127718,I127701,);
nor I_7367 (I128125,I388042,I388048);
not I_7368 (I128142,I128125);
nor I_7369 (I127704,I127981,I128142);
nand I_7370 (I127689,I127998,I128142);
nor I_7371 (I127698,I127744,I128125);
DFFARX1 I_7372 (I128125,I2859,I127718,I127707,);
not I_7373 (I128245,I2866);
DFFARX1 I_7374 (I175431,I2859,I128245,I128271,);
nand I_7375 (I128279,I175443,I175422);
and I_7376 (I128296,I128279,I175446);
DFFARX1 I_7377 (I128296,I2859,I128245,I128322,);
nor I_7378 (I128213,I128322,I128271);
not I_7379 (I128344,I128322);
DFFARX1 I_7380 (I175437,I2859,I128245,I128370,);
nand I_7381 (I128378,I128370,I175419);
not I_7382 (I128395,I128378);
DFFARX1 I_7383 (I128395,I2859,I128245,I128421,);
not I_7384 (I128237,I128421);
nor I_7385 (I128443,I128271,I128378);
nor I_7386 (I128219,I128322,I128443);
DFFARX1 I_7387 (I175434,I2859,I128245,I128483,);
DFFARX1 I_7388 (I128483,I2859,I128245,I128500,);
not I_7389 (I128508,I128500);
not I_7390 (I128525,I128483);
nand I_7391 (I128222,I128525,I128344);
nand I_7392 (I128556,I175419,I175425);
and I_7393 (I128573,I128556,I175428);
DFFARX1 I_7394 (I128573,I2859,I128245,I128599,);
nor I_7395 (I128607,I128599,I128271);
DFFARX1 I_7396 (I128607,I2859,I128245,I128210,);
DFFARX1 I_7397 (I128599,I2859,I128245,I128228,);
nor I_7398 (I128652,I175440,I175425);
not I_7399 (I128669,I128652);
nor I_7400 (I128231,I128508,I128669);
nand I_7401 (I128216,I128525,I128669);
nor I_7402 (I128225,I128271,I128652);
DFFARX1 I_7403 (I128652,I2859,I128245,I128234,);
not I_7404 (I128772,I2866);
DFFARX1 I_7405 (I81018,I2859,I128772,I128798,);
nand I_7406 (I128806,I81018,I81024);
and I_7407 (I128823,I128806,I81042);
DFFARX1 I_7408 (I128823,I2859,I128772,I128849,);
nor I_7409 (I128740,I128849,I128798);
not I_7410 (I128871,I128849);
DFFARX1 I_7411 (I81030,I2859,I128772,I128897,);
nand I_7412 (I128905,I128897,I81027);
not I_7413 (I128922,I128905);
DFFARX1 I_7414 (I128922,I2859,I128772,I128948,);
not I_7415 (I128764,I128948);
nor I_7416 (I128970,I128798,I128905);
nor I_7417 (I128746,I128849,I128970);
DFFARX1 I_7418 (I81036,I2859,I128772,I129010,);
DFFARX1 I_7419 (I129010,I2859,I128772,I129027,);
not I_7420 (I129035,I129027);
not I_7421 (I129052,I129010);
nand I_7422 (I128749,I129052,I128871);
nand I_7423 (I129083,I81021,I81021);
and I_7424 (I129100,I129083,I81033);
DFFARX1 I_7425 (I129100,I2859,I128772,I129126,);
nor I_7426 (I129134,I129126,I128798);
DFFARX1 I_7427 (I129134,I2859,I128772,I128737,);
DFFARX1 I_7428 (I129126,I2859,I128772,I128755,);
nor I_7429 (I129179,I81039,I81021);
not I_7430 (I129196,I129179);
nor I_7431 (I128758,I129035,I129196);
nand I_7432 (I128743,I129052,I129196);
nor I_7433 (I128752,I128798,I129179);
DFFARX1 I_7434 (I129179,I2859,I128772,I128761,);
not I_7435 (I129299,I2866);
DFFARX1 I_7436 (I329774,I2859,I129299,I129325,);
nand I_7437 (I129333,I329765,I329780);
and I_7438 (I129350,I129333,I329786);
DFFARX1 I_7439 (I129350,I2859,I129299,I129376,);
nor I_7440 (I129267,I129376,I129325);
not I_7441 (I129398,I129376);
DFFARX1 I_7442 (I329771,I2859,I129299,I129424,);
nand I_7443 (I129432,I129424,I329765);
not I_7444 (I129449,I129432);
DFFARX1 I_7445 (I129449,I2859,I129299,I129475,);
not I_7446 (I129291,I129475);
nor I_7447 (I129497,I129325,I129432);
nor I_7448 (I129273,I129376,I129497);
DFFARX1 I_7449 (I329768,I2859,I129299,I129537,);
DFFARX1 I_7450 (I129537,I2859,I129299,I129554,);
not I_7451 (I129562,I129554);
not I_7452 (I129579,I129537);
nand I_7453 (I129276,I129579,I129398);
nand I_7454 (I129610,I329762,I329777);
and I_7455 (I129627,I129610,I329762);
DFFARX1 I_7456 (I129627,I2859,I129299,I129653,);
nor I_7457 (I129661,I129653,I129325);
DFFARX1 I_7458 (I129661,I2859,I129299,I129264,);
DFFARX1 I_7459 (I129653,I2859,I129299,I129282,);
nor I_7460 (I129706,I329783,I329777);
not I_7461 (I129723,I129706);
nor I_7462 (I129285,I129562,I129723);
nand I_7463 (I129270,I129579,I129723);
nor I_7464 (I129279,I129325,I129706);
DFFARX1 I_7465 (I129706,I2859,I129299,I129288,);
not I_7466 (I129826,I2866);
DFFARX1 I_7467 (I505356,I2859,I129826,I129852,);
nand I_7468 (I129860,I505338,I505362);
and I_7469 (I129877,I129860,I505353);
DFFARX1 I_7470 (I129877,I2859,I129826,I129903,);
nor I_7471 (I129794,I129903,I129852);
not I_7472 (I129925,I129903);
DFFARX1 I_7473 (I505359,I2859,I129826,I129951,);
nand I_7474 (I129959,I129951,I505347);
not I_7475 (I129976,I129959);
DFFARX1 I_7476 (I129976,I2859,I129826,I130002,);
not I_7477 (I129818,I130002);
nor I_7478 (I130024,I129852,I129959);
nor I_7479 (I129800,I129903,I130024);
DFFARX1 I_7480 (I505338,I2859,I129826,I130064,);
DFFARX1 I_7481 (I130064,I2859,I129826,I130081,);
not I_7482 (I130089,I130081);
not I_7483 (I130106,I130064);
nand I_7484 (I129803,I130106,I129925);
nand I_7485 (I130137,I505344,I505341);
and I_7486 (I130154,I130137,I505350);
DFFARX1 I_7487 (I130154,I2859,I129826,I130180,);
nor I_7488 (I130188,I130180,I129852);
DFFARX1 I_7489 (I130188,I2859,I129826,I129791,);
DFFARX1 I_7490 (I130180,I2859,I129826,I129809,);
nor I_7491 (I130233,I505341,I505341);
not I_7492 (I130250,I130233);
nor I_7493 (I129812,I130089,I130250);
nand I_7494 (I129797,I130106,I130250);
nor I_7495 (I129806,I129852,I130233);
DFFARX1 I_7496 (I130233,I2859,I129826,I129815,);
not I_7497 (I130353,I2866);
DFFARX1 I_7498 (I94108,I2859,I130353,I130379,);
nand I_7499 (I130387,I94108,I94114);
and I_7500 (I130404,I130387,I94132);
DFFARX1 I_7501 (I130404,I2859,I130353,I130430,);
nor I_7502 (I130321,I130430,I130379);
not I_7503 (I130452,I130430);
DFFARX1 I_7504 (I94120,I2859,I130353,I130478,);
nand I_7505 (I130486,I130478,I94117);
not I_7506 (I130503,I130486);
DFFARX1 I_7507 (I130503,I2859,I130353,I130529,);
not I_7508 (I130345,I130529);
nor I_7509 (I130551,I130379,I130486);
nor I_7510 (I130327,I130430,I130551);
DFFARX1 I_7511 (I94126,I2859,I130353,I130591,);
DFFARX1 I_7512 (I130591,I2859,I130353,I130608,);
not I_7513 (I130616,I130608);
not I_7514 (I130633,I130591);
nand I_7515 (I130330,I130633,I130452);
nand I_7516 (I130664,I94111,I94111);
and I_7517 (I130681,I130664,I94123);
DFFARX1 I_7518 (I130681,I2859,I130353,I130707,);
nor I_7519 (I130715,I130707,I130379);
DFFARX1 I_7520 (I130715,I2859,I130353,I130318,);
DFFARX1 I_7521 (I130707,I2859,I130353,I130336,);
nor I_7522 (I130760,I94129,I94111);
not I_7523 (I130777,I130760);
nor I_7524 (I130339,I130616,I130777);
nand I_7525 (I130324,I130633,I130777);
nor I_7526 (I130333,I130379,I130760);
DFFARX1 I_7527 (I130760,I2859,I130353,I130342,);
not I_7528 (I130880,I2866);
DFFARX1 I_7529 (I486468,I2859,I130880,I130906,);
nand I_7530 (I130914,I486483,I486468);
and I_7531 (I130931,I130914,I486486);
DFFARX1 I_7532 (I130931,I2859,I130880,I130957,);
nor I_7533 (I130848,I130957,I130906);
not I_7534 (I130979,I130957);
DFFARX1 I_7535 (I486492,I2859,I130880,I131005,);
nand I_7536 (I131013,I131005,I486474);
not I_7537 (I131030,I131013);
DFFARX1 I_7538 (I131030,I2859,I130880,I131056,);
not I_7539 (I130872,I131056);
nor I_7540 (I131078,I130906,I131013);
nor I_7541 (I130854,I130957,I131078);
DFFARX1 I_7542 (I486471,I2859,I130880,I131118,);
DFFARX1 I_7543 (I131118,I2859,I130880,I131135,);
not I_7544 (I131143,I131135);
not I_7545 (I131160,I131118);
nand I_7546 (I130857,I131160,I130979);
nand I_7547 (I131191,I486471,I486477);
and I_7548 (I131208,I131191,I486489);
DFFARX1 I_7549 (I131208,I2859,I130880,I131234,);
nor I_7550 (I131242,I131234,I130906);
DFFARX1 I_7551 (I131242,I2859,I130880,I130845,);
DFFARX1 I_7552 (I131234,I2859,I130880,I130863,);
nor I_7553 (I131287,I486480,I486477);
not I_7554 (I131304,I131287);
nor I_7555 (I130866,I131143,I131304);
nand I_7556 (I130851,I131160,I131304);
nor I_7557 (I130860,I130906,I131287);
DFFARX1 I_7558 (I131287,I2859,I130880,I130869,);
not I_7559 (I131407,I2866);
DFFARX1 I_7560 (I288158,I2859,I131407,I131433,);
nand I_7561 (I131441,I288149,I288164);
and I_7562 (I131458,I131441,I288170);
DFFARX1 I_7563 (I131458,I2859,I131407,I131484,);
nor I_7564 (I131375,I131484,I131433);
not I_7565 (I131506,I131484);
DFFARX1 I_7566 (I288155,I2859,I131407,I131532,);
nand I_7567 (I131540,I131532,I288149);
not I_7568 (I131557,I131540);
DFFARX1 I_7569 (I131557,I2859,I131407,I131583,);
not I_7570 (I131399,I131583);
nor I_7571 (I131605,I131433,I131540);
nor I_7572 (I131381,I131484,I131605);
DFFARX1 I_7573 (I288152,I2859,I131407,I131645,);
DFFARX1 I_7574 (I131645,I2859,I131407,I131662,);
not I_7575 (I131670,I131662);
not I_7576 (I131687,I131645);
nand I_7577 (I131384,I131687,I131506);
nand I_7578 (I131718,I288146,I288161);
and I_7579 (I131735,I131718,I288146);
DFFARX1 I_7580 (I131735,I2859,I131407,I131761,);
nor I_7581 (I131769,I131761,I131433);
DFFARX1 I_7582 (I131769,I2859,I131407,I131372,);
DFFARX1 I_7583 (I131761,I2859,I131407,I131390,);
nor I_7584 (I131814,I288167,I288161);
not I_7585 (I131831,I131814);
nor I_7586 (I131393,I131670,I131831);
nand I_7587 (I131378,I131687,I131831);
nor I_7588 (I131387,I131433,I131814);
DFFARX1 I_7589 (I131814,I2859,I131407,I131396,);
not I_7590 (I131934,I2866);
DFFARX1 I_7591 (I229176,I2859,I131934,I131960,);
nand I_7592 (I131968,I229176,I229188);
and I_7593 (I131985,I131968,I229173);
DFFARX1 I_7594 (I131985,I2859,I131934,I132011,);
nor I_7595 (I131902,I132011,I131960);
not I_7596 (I132033,I132011);
DFFARX1 I_7597 (I229197,I2859,I131934,I132059,);
nand I_7598 (I132067,I132059,I229194);
not I_7599 (I132084,I132067);
DFFARX1 I_7600 (I132084,I2859,I131934,I132110,);
not I_7601 (I131926,I132110);
nor I_7602 (I132132,I131960,I132067);
nor I_7603 (I131908,I132011,I132132);
DFFARX1 I_7604 (I229185,I2859,I131934,I132172,);
DFFARX1 I_7605 (I132172,I2859,I131934,I132189,);
not I_7606 (I132197,I132189);
not I_7607 (I132214,I132172);
nand I_7608 (I131911,I132214,I132033);
nand I_7609 (I132245,I229173,I229182);
and I_7610 (I132262,I132245,I229191);
DFFARX1 I_7611 (I132262,I2859,I131934,I132288,);
nor I_7612 (I132296,I132288,I131960);
DFFARX1 I_7613 (I132296,I2859,I131934,I131899,);
DFFARX1 I_7614 (I132288,I2859,I131934,I131917,);
nor I_7615 (I132341,I229179,I229182);
not I_7616 (I132358,I132341);
nor I_7617 (I131920,I132197,I132358);
nand I_7618 (I131905,I132214,I132358);
nor I_7619 (I131914,I131960,I132341);
DFFARX1 I_7620 (I132341,I2859,I131934,I131923,);
not I_7621 (I132461,I2866);
DFFARX1 I_7622 (I400298,I2859,I132461,I132487,);
nand I_7623 (I132495,I400295,I400313);
and I_7624 (I132512,I132495,I400304);
DFFARX1 I_7625 (I132512,I2859,I132461,I132538,);
nor I_7626 (I132429,I132538,I132487);
not I_7627 (I132560,I132538);
DFFARX1 I_7628 (I400319,I2859,I132461,I132586,);
nand I_7629 (I132594,I132586,I400301);
not I_7630 (I132611,I132594);
DFFARX1 I_7631 (I132611,I2859,I132461,I132637,);
not I_7632 (I132453,I132637);
nor I_7633 (I132659,I132487,I132594);
nor I_7634 (I132435,I132538,I132659);
DFFARX1 I_7635 (I400307,I2859,I132461,I132699,);
DFFARX1 I_7636 (I132699,I2859,I132461,I132716,);
not I_7637 (I132724,I132716);
not I_7638 (I132741,I132699);
nand I_7639 (I132438,I132741,I132560);
nand I_7640 (I132772,I400295,I400322);
and I_7641 (I132789,I132772,I400310);
DFFARX1 I_7642 (I132789,I2859,I132461,I132815,);
nor I_7643 (I132823,I132815,I132487);
DFFARX1 I_7644 (I132823,I2859,I132461,I132426,);
DFFARX1 I_7645 (I132815,I2859,I132461,I132444,);
nor I_7646 (I132868,I400316,I400322);
not I_7647 (I132885,I132868);
nor I_7648 (I132447,I132724,I132885);
nand I_7649 (I132432,I132741,I132885);
nor I_7650 (I132441,I132487,I132868);
DFFARX1 I_7651 (I132868,I2859,I132461,I132450,);
not I_7652 (I132988,I2866);
DFFARX1 I_7653 (I280644,I2859,I132988,I133014,);
nand I_7654 (I133022,I280635,I280650);
and I_7655 (I133039,I133022,I280656);
DFFARX1 I_7656 (I133039,I2859,I132988,I133065,);
nor I_7657 (I132956,I133065,I133014);
not I_7658 (I133087,I133065);
DFFARX1 I_7659 (I280641,I2859,I132988,I133113,);
nand I_7660 (I133121,I133113,I280635);
not I_7661 (I133138,I133121);
DFFARX1 I_7662 (I133138,I2859,I132988,I133164,);
not I_7663 (I132980,I133164);
nor I_7664 (I133186,I133014,I133121);
nor I_7665 (I132962,I133065,I133186);
DFFARX1 I_7666 (I280638,I2859,I132988,I133226,);
DFFARX1 I_7667 (I133226,I2859,I132988,I133243,);
not I_7668 (I133251,I133243);
not I_7669 (I133268,I133226);
nand I_7670 (I132965,I133268,I133087);
nand I_7671 (I133299,I280632,I280647);
and I_7672 (I133316,I133299,I280632);
DFFARX1 I_7673 (I133316,I2859,I132988,I133342,);
nor I_7674 (I133350,I133342,I133014);
DFFARX1 I_7675 (I133350,I2859,I132988,I132953,);
DFFARX1 I_7676 (I133342,I2859,I132988,I132971,);
nor I_7677 (I133395,I280653,I280647);
not I_7678 (I133412,I133395);
nor I_7679 (I132974,I133251,I133412);
nand I_7680 (I132959,I133268,I133412);
nor I_7681 (I132968,I133014,I133395);
DFFARX1 I_7682 (I133395,I2859,I132988,I132977,);
not I_7683 (I133515,I2866);
DFFARX1 I_7684 (I50506,I2859,I133515,I133541,);
nand I_7685 (I133549,I50518,I50527);
and I_7686 (I133566,I133549,I50506);
DFFARX1 I_7687 (I133566,I2859,I133515,I133592,);
nor I_7688 (I133483,I133592,I133541);
not I_7689 (I133614,I133592);
DFFARX1 I_7690 (I50521,I2859,I133515,I133640,);
nand I_7691 (I133648,I133640,I50509);
not I_7692 (I133665,I133648);
DFFARX1 I_7693 (I133665,I2859,I133515,I133691,);
not I_7694 (I133507,I133691);
nor I_7695 (I133713,I133541,I133648);
nor I_7696 (I133489,I133592,I133713);
DFFARX1 I_7697 (I50512,I2859,I133515,I133753,);
DFFARX1 I_7698 (I133753,I2859,I133515,I133770,);
not I_7699 (I133778,I133770);
not I_7700 (I133795,I133753);
nand I_7701 (I133492,I133795,I133614);
nand I_7702 (I133826,I50503,I50503);
and I_7703 (I133843,I133826,I50515);
DFFARX1 I_7704 (I133843,I2859,I133515,I133869,);
nor I_7705 (I133877,I133869,I133541);
DFFARX1 I_7706 (I133877,I2859,I133515,I133480,);
DFFARX1 I_7707 (I133869,I2859,I133515,I133498,);
nor I_7708 (I133922,I50524,I50503);
not I_7709 (I133939,I133922);
nor I_7710 (I133501,I133778,I133939);
nand I_7711 (I133486,I133795,I133939);
nor I_7712 (I133495,I133541,I133922);
DFFARX1 I_7713 (I133922,I2859,I133515,I133504,);
not I_7714 (I134042,I2866);
DFFARX1 I_7715 (I101843,I2859,I134042,I134068,);
nand I_7716 (I134076,I101843,I101849);
and I_7717 (I134093,I134076,I101867);
DFFARX1 I_7718 (I134093,I2859,I134042,I134119,);
nor I_7719 (I134010,I134119,I134068);
not I_7720 (I134141,I134119);
DFFARX1 I_7721 (I101855,I2859,I134042,I134167,);
nand I_7722 (I134175,I134167,I101852);
not I_7723 (I134192,I134175);
DFFARX1 I_7724 (I134192,I2859,I134042,I134218,);
not I_7725 (I134034,I134218);
nor I_7726 (I134240,I134068,I134175);
nor I_7727 (I134016,I134119,I134240);
DFFARX1 I_7728 (I101861,I2859,I134042,I134280,);
DFFARX1 I_7729 (I134280,I2859,I134042,I134297,);
not I_7730 (I134305,I134297);
not I_7731 (I134322,I134280);
nand I_7732 (I134019,I134322,I134141);
nand I_7733 (I134353,I101846,I101846);
and I_7734 (I134370,I134353,I101858);
DFFARX1 I_7735 (I134370,I2859,I134042,I134396,);
nor I_7736 (I134404,I134396,I134068);
DFFARX1 I_7737 (I134404,I2859,I134042,I134007,);
DFFARX1 I_7738 (I134396,I2859,I134042,I134025,);
nor I_7739 (I134449,I101864,I101846);
not I_7740 (I134466,I134449);
nor I_7741 (I134028,I134305,I134466);
nand I_7742 (I134013,I134322,I134466);
nor I_7743 (I134022,I134068,I134449);
DFFARX1 I_7744 (I134449,I2859,I134042,I134031,);
not I_7745 (I134569,I2866);
DFFARX1 I_7746 (I300874,I2859,I134569,I134595,);
nand I_7747 (I134603,I300865,I300880);
and I_7748 (I134620,I134603,I300886);
DFFARX1 I_7749 (I134620,I2859,I134569,I134646,);
nor I_7750 (I134537,I134646,I134595);
not I_7751 (I134668,I134646);
DFFARX1 I_7752 (I300871,I2859,I134569,I134694,);
nand I_7753 (I134702,I134694,I300865);
not I_7754 (I134719,I134702);
DFFARX1 I_7755 (I134719,I2859,I134569,I134745,);
not I_7756 (I134561,I134745);
nor I_7757 (I134767,I134595,I134702);
nor I_7758 (I134543,I134646,I134767);
DFFARX1 I_7759 (I300868,I2859,I134569,I134807,);
DFFARX1 I_7760 (I134807,I2859,I134569,I134824,);
not I_7761 (I134832,I134824);
not I_7762 (I134849,I134807);
nand I_7763 (I134546,I134849,I134668);
nand I_7764 (I134880,I300862,I300877);
and I_7765 (I134897,I134880,I300862);
DFFARX1 I_7766 (I134897,I2859,I134569,I134923,);
nor I_7767 (I134931,I134923,I134595);
DFFARX1 I_7768 (I134931,I2859,I134569,I134534,);
DFFARX1 I_7769 (I134923,I2859,I134569,I134552,);
nor I_7770 (I134976,I300883,I300877);
not I_7771 (I134993,I134976);
nor I_7772 (I134555,I134832,I134993);
nand I_7773 (I134540,I134849,I134993);
nor I_7774 (I134549,I134595,I134976);
DFFARX1 I_7775 (I134976,I2859,I134569,I134558,);
not I_7776 (I135096,I2866);
DFFARX1 I_7777 (I328040,I2859,I135096,I135122,);
nand I_7778 (I135130,I328031,I328046);
and I_7779 (I135147,I135130,I328052);
DFFARX1 I_7780 (I135147,I2859,I135096,I135173,);
nor I_7781 (I135064,I135173,I135122);
not I_7782 (I135195,I135173);
DFFARX1 I_7783 (I328037,I2859,I135096,I135221,);
nand I_7784 (I135229,I135221,I328031);
not I_7785 (I135246,I135229);
DFFARX1 I_7786 (I135246,I2859,I135096,I135272,);
not I_7787 (I135088,I135272);
nor I_7788 (I135294,I135122,I135229);
nor I_7789 (I135070,I135173,I135294);
DFFARX1 I_7790 (I328034,I2859,I135096,I135334,);
DFFARX1 I_7791 (I135334,I2859,I135096,I135351,);
not I_7792 (I135359,I135351);
not I_7793 (I135376,I135334);
nand I_7794 (I135073,I135376,I135195);
nand I_7795 (I135407,I328028,I328043);
and I_7796 (I135424,I135407,I328028);
DFFARX1 I_7797 (I135424,I2859,I135096,I135450,);
nor I_7798 (I135458,I135450,I135122);
DFFARX1 I_7799 (I135458,I2859,I135096,I135061,);
DFFARX1 I_7800 (I135450,I2859,I135096,I135079,);
nor I_7801 (I135503,I328049,I328043);
not I_7802 (I135520,I135503);
nor I_7803 (I135082,I135359,I135520);
nand I_7804 (I135067,I135376,I135520);
nor I_7805 (I135076,I135122,I135503);
DFFARX1 I_7806 (I135503,I2859,I135096,I135085,);
not I_7807 (I135623,I2866);
DFFARX1 I_7808 (I384794,I2859,I135623,I135649,);
nand I_7809 (I135657,I384791,I384809);
and I_7810 (I135674,I135657,I384800);
DFFARX1 I_7811 (I135674,I2859,I135623,I135700,);
nor I_7812 (I135591,I135700,I135649);
not I_7813 (I135722,I135700);
DFFARX1 I_7814 (I384815,I2859,I135623,I135748,);
nand I_7815 (I135756,I135748,I384797);
not I_7816 (I135773,I135756);
DFFARX1 I_7817 (I135773,I2859,I135623,I135799,);
not I_7818 (I135615,I135799);
nor I_7819 (I135821,I135649,I135756);
nor I_7820 (I135597,I135700,I135821);
DFFARX1 I_7821 (I384803,I2859,I135623,I135861,);
DFFARX1 I_7822 (I135861,I2859,I135623,I135878,);
not I_7823 (I135886,I135878);
not I_7824 (I135903,I135861);
nand I_7825 (I135600,I135903,I135722);
nand I_7826 (I135934,I384791,I384818);
and I_7827 (I135951,I135934,I384806);
DFFARX1 I_7828 (I135951,I2859,I135623,I135977,);
nor I_7829 (I135985,I135977,I135649);
DFFARX1 I_7830 (I135985,I2859,I135623,I135588,);
DFFARX1 I_7831 (I135977,I2859,I135623,I135606,);
nor I_7832 (I136030,I384812,I384818);
not I_7833 (I136047,I136030);
nor I_7834 (I135609,I135886,I136047);
nand I_7835 (I135594,I135903,I136047);
nor I_7836 (I135603,I135649,I136030);
DFFARX1 I_7837 (I136030,I2859,I135623,I135612,);
not I_7838 (I136150,I2866);
DFFARX1 I_7839 (I278332,I2859,I136150,I136176,);
nand I_7840 (I136184,I278323,I278338);
and I_7841 (I136201,I136184,I278344);
DFFARX1 I_7842 (I136201,I2859,I136150,I136227,);
nor I_7843 (I136118,I136227,I136176);
not I_7844 (I136249,I136227);
DFFARX1 I_7845 (I278329,I2859,I136150,I136275,);
nand I_7846 (I136283,I136275,I278323);
not I_7847 (I136300,I136283);
DFFARX1 I_7848 (I136300,I2859,I136150,I136326,);
not I_7849 (I136142,I136326);
nor I_7850 (I136348,I136176,I136283);
nor I_7851 (I136124,I136227,I136348);
DFFARX1 I_7852 (I278326,I2859,I136150,I136388,);
DFFARX1 I_7853 (I136388,I2859,I136150,I136405,);
not I_7854 (I136413,I136405);
not I_7855 (I136430,I136388);
nand I_7856 (I136127,I136430,I136249);
nand I_7857 (I136461,I278320,I278335);
and I_7858 (I136478,I136461,I278320);
DFFARX1 I_7859 (I136478,I2859,I136150,I136504,);
nor I_7860 (I136512,I136504,I136176);
DFFARX1 I_7861 (I136512,I2859,I136150,I136115,);
DFFARX1 I_7862 (I136504,I2859,I136150,I136133,);
nor I_7863 (I136557,I278341,I278335);
not I_7864 (I136574,I136557);
nor I_7865 (I136136,I136413,I136574);
nand I_7866 (I136121,I136430,I136574);
nor I_7867 (I136130,I136176,I136557);
DFFARX1 I_7868 (I136557,I2859,I136150,I136139,);
not I_7869 (I136677,I2866);
DFFARX1 I_7870 (I443835,I2859,I136677,I136703,);
nand I_7871 (I136711,I443832,I443835);
and I_7872 (I136728,I136711,I443844);
DFFARX1 I_7873 (I136728,I2859,I136677,I136754,);
nor I_7874 (I136645,I136754,I136703);
not I_7875 (I136776,I136754);
DFFARX1 I_7876 (I443832,I2859,I136677,I136802,);
nand I_7877 (I136810,I136802,I443850);
not I_7878 (I136827,I136810);
DFFARX1 I_7879 (I136827,I2859,I136677,I136853,);
not I_7880 (I136669,I136853);
nor I_7881 (I136875,I136703,I136810);
nor I_7882 (I136651,I136754,I136875);
DFFARX1 I_7883 (I443838,I2859,I136677,I136915,);
DFFARX1 I_7884 (I136915,I2859,I136677,I136932,);
not I_7885 (I136940,I136932);
not I_7886 (I136957,I136915);
nand I_7887 (I136654,I136957,I136776);
nand I_7888 (I136988,I443847,I443853);
and I_7889 (I137005,I136988,I443838);
DFFARX1 I_7890 (I137005,I2859,I136677,I137031,);
nor I_7891 (I137039,I137031,I136703);
DFFARX1 I_7892 (I137039,I2859,I136677,I136642,);
DFFARX1 I_7893 (I137031,I2859,I136677,I136660,);
nor I_7894 (I137084,I443841,I443853);
not I_7895 (I137101,I137084);
nor I_7896 (I136663,I136940,I137101);
nand I_7897 (I136648,I136957,I137101);
nor I_7898 (I136657,I136703,I137084);
DFFARX1 I_7899 (I137084,I2859,I136677,I136666,);
not I_7900 (I137204,I2866);
DFFARX1 I_7901 (I88753,I2859,I137204,I137230,);
nand I_7902 (I137238,I88753,I88759);
and I_7903 (I137255,I137238,I88777);
DFFARX1 I_7904 (I137255,I2859,I137204,I137281,);
nor I_7905 (I137172,I137281,I137230);
not I_7906 (I137303,I137281);
DFFARX1 I_7907 (I88765,I2859,I137204,I137329,);
nand I_7908 (I137337,I137329,I88762);
not I_7909 (I137354,I137337);
DFFARX1 I_7910 (I137354,I2859,I137204,I137380,);
not I_7911 (I137196,I137380);
nor I_7912 (I137402,I137230,I137337);
nor I_7913 (I137178,I137281,I137402);
DFFARX1 I_7914 (I88771,I2859,I137204,I137442,);
DFFARX1 I_7915 (I137442,I2859,I137204,I137459,);
not I_7916 (I137467,I137459);
not I_7917 (I137484,I137442);
nand I_7918 (I137181,I137484,I137303);
nand I_7919 (I137515,I88756,I88756);
and I_7920 (I137532,I137515,I88768);
DFFARX1 I_7921 (I137532,I2859,I137204,I137558,);
nor I_7922 (I137566,I137558,I137230);
DFFARX1 I_7923 (I137566,I2859,I137204,I137169,);
DFFARX1 I_7924 (I137558,I2859,I137204,I137187,);
nor I_7925 (I137611,I88774,I88756);
not I_7926 (I137628,I137611);
nor I_7927 (I137190,I137467,I137628);
nand I_7928 (I137175,I137484,I137628);
nor I_7929 (I137184,I137230,I137611);
DFFARX1 I_7930 (I137611,I2859,I137204,I137193,);
not I_7931 (I137731,I2866);
DFFARX1 I_7932 (I341614,I2859,I137731,I137757,);
nand I_7933 (I137765,I341617,I341611);
and I_7934 (I137782,I137765,I341623);
DFFARX1 I_7935 (I137782,I2859,I137731,I137808,);
nor I_7936 (I137699,I137808,I137757);
not I_7937 (I137830,I137808);
DFFARX1 I_7938 (I341626,I2859,I137731,I137856,);
nand I_7939 (I137864,I137856,I341617);
not I_7940 (I137881,I137864);
DFFARX1 I_7941 (I137881,I2859,I137731,I137907,);
not I_7942 (I137723,I137907);
nor I_7943 (I137929,I137757,I137864);
nor I_7944 (I137705,I137808,I137929);
DFFARX1 I_7945 (I341629,I2859,I137731,I137969,);
DFFARX1 I_7946 (I137969,I2859,I137731,I137986,);
not I_7947 (I137994,I137986);
not I_7948 (I138011,I137969);
nand I_7949 (I137708,I138011,I137830);
nand I_7950 (I138042,I341611,I341620);
and I_7951 (I138059,I138042,I341614);
DFFARX1 I_7952 (I138059,I2859,I137731,I138085,);
nor I_7953 (I138093,I138085,I137757);
DFFARX1 I_7954 (I138093,I2859,I137731,I137696,);
DFFARX1 I_7955 (I138085,I2859,I137731,I137714,);
nor I_7956 (I138138,I341632,I341620);
not I_7957 (I138155,I138138);
nor I_7958 (I137717,I137994,I138155);
nand I_7959 (I137702,I138011,I138155);
nor I_7960 (I137711,I137757,I138138);
DFFARX1 I_7961 (I138138,I2859,I137731,I137720,);
not I_7962 (I138258,I2866);
DFFARX1 I_7963 (I2668,I2859,I138258,I138284,);
nand I_7964 (I138292,I1964,I2828);
and I_7965 (I138309,I138292,I1836);
DFFARX1 I_7966 (I138309,I2859,I138258,I138335,);
nor I_7967 (I138226,I138335,I138284);
not I_7968 (I138357,I138335);
DFFARX1 I_7969 (I2780,I2859,I138258,I138383,);
nand I_7970 (I138391,I138383,I2212);
not I_7971 (I138408,I138391);
DFFARX1 I_7972 (I138408,I2859,I138258,I138434,);
not I_7973 (I138250,I138434);
nor I_7974 (I138456,I138284,I138391);
nor I_7975 (I138232,I138335,I138456);
DFFARX1 I_7976 (I1732,I2859,I138258,I138496,);
DFFARX1 I_7977 (I138496,I2859,I138258,I138513,);
not I_7978 (I138521,I138513);
not I_7979 (I138538,I138496);
nand I_7980 (I138235,I138538,I138357);
nand I_7981 (I138569,I1484,I2260);
and I_7982 (I138586,I138569,I2220);
DFFARX1 I_7983 (I138586,I2859,I138258,I138612,);
nor I_7984 (I138620,I138612,I138284);
DFFARX1 I_7985 (I138620,I2859,I138258,I138223,);
DFFARX1 I_7986 (I138612,I2859,I138258,I138241,);
nor I_7987 (I138665,I1572,I2260);
not I_7988 (I138682,I138665);
nor I_7989 (I138244,I138521,I138682);
nand I_7990 (I138229,I138538,I138682);
nor I_7991 (I138238,I138284,I138665);
DFFARX1 I_7992 (I138665,I2859,I138258,I138247,);
not I_7993 (I138785,I2866);
DFFARX1 I_7994 (I336344,I2859,I138785,I138811,);
nand I_7995 (I138819,I336347,I336341);
and I_7996 (I138836,I138819,I336353);
DFFARX1 I_7997 (I138836,I2859,I138785,I138862,);
nor I_7998 (I138753,I138862,I138811);
not I_7999 (I138884,I138862);
DFFARX1 I_8000 (I336356,I2859,I138785,I138910,);
nand I_8001 (I138918,I138910,I336347);
not I_8002 (I138935,I138918);
DFFARX1 I_8003 (I138935,I2859,I138785,I138961,);
not I_8004 (I138777,I138961);
nor I_8005 (I138983,I138811,I138918);
nor I_8006 (I138759,I138862,I138983);
DFFARX1 I_8007 (I336359,I2859,I138785,I139023,);
DFFARX1 I_8008 (I139023,I2859,I138785,I139040,);
not I_8009 (I139048,I139040);
not I_8010 (I139065,I139023);
nand I_8011 (I138762,I139065,I138884);
nand I_8012 (I139096,I336341,I336350);
and I_8013 (I139113,I139096,I336344);
DFFARX1 I_8014 (I139113,I2859,I138785,I139139,);
nor I_8015 (I139147,I139139,I138811);
DFFARX1 I_8016 (I139147,I2859,I138785,I138750,);
DFFARX1 I_8017 (I139139,I2859,I138785,I138768,);
nor I_8018 (I139192,I336362,I336350);
not I_8019 (I139209,I139192);
nor I_8020 (I138771,I139048,I139209);
nand I_8021 (I138756,I139065,I139209);
nor I_8022 (I138765,I138811,I139192);
DFFARX1 I_8023 (I139192,I2859,I138785,I138774,);
not I_8024 (I139312,I2866);
DFFARX1 I_8025 (I99463,I2859,I139312,I139338,);
nand I_8026 (I139346,I99463,I99469);
and I_8027 (I139363,I139346,I99487);
DFFARX1 I_8028 (I139363,I2859,I139312,I139389,);
nor I_8029 (I139280,I139389,I139338);
not I_8030 (I139411,I139389);
DFFARX1 I_8031 (I99475,I2859,I139312,I139437,);
nand I_8032 (I139445,I139437,I99472);
not I_8033 (I139462,I139445);
DFFARX1 I_8034 (I139462,I2859,I139312,I139488,);
not I_8035 (I139304,I139488);
nor I_8036 (I139510,I139338,I139445);
nor I_8037 (I139286,I139389,I139510);
DFFARX1 I_8038 (I99481,I2859,I139312,I139550,);
DFFARX1 I_8039 (I139550,I2859,I139312,I139567,);
not I_8040 (I139575,I139567);
not I_8041 (I139592,I139550);
nand I_8042 (I139289,I139592,I139411);
nand I_8043 (I139623,I99466,I99466);
and I_8044 (I139640,I139623,I99478);
DFFARX1 I_8045 (I139640,I2859,I139312,I139666,);
nor I_8046 (I139674,I139666,I139338);
DFFARX1 I_8047 (I139674,I2859,I139312,I139277,);
DFFARX1 I_8048 (I139666,I2859,I139312,I139295,);
nor I_8049 (I139719,I99484,I99466);
not I_8050 (I139736,I139719);
nor I_8051 (I139298,I139575,I139736);
nand I_8052 (I139283,I139592,I139736);
nor I_8053 (I139292,I139338,I139719);
DFFARX1 I_8054 (I139719,I2859,I139312,I139301,);
not I_8055 (I139839,I2866);
DFFARX1 I_8056 (I558586,I2859,I139839,I139865,);
nand I_8057 (I139873,I558565,I558565);
and I_8058 (I139890,I139873,I558592);
DFFARX1 I_8059 (I139890,I2859,I139839,I139916,);
nor I_8060 (I139807,I139916,I139865);
not I_8061 (I139938,I139916);
DFFARX1 I_8062 (I558580,I2859,I139839,I139964,);
nand I_8063 (I139972,I139964,I558583);
not I_8064 (I139989,I139972);
DFFARX1 I_8065 (I139989,I2859,I139839,I140015,);
not I_8066 (I139831,I140015);
nor I_8067 (I140037,I139865,I139972);
nor I_8068 (I139813,I139916,I140037);
DFFARX1 I_8069 (I558574,I2859,I139839,I140077,);
DFFARX1 I_8070 (I140077,I2859,I139839,I140094,);
not I_8071 (I140102,I140094);
not I_8072 (I140119,I140077);
nand I_8073 (I139816,I140119,I139938);
nand I_8074 (I140150,I558571,I558568);
and I_8075 (I140167,I140150,I558589);
DFFARX1 I_8076 (I140167,I2859,I139839,I140193,);
nor I_8077 (I140201,I140193,I139865);
DFFARX1 I_8078 (I140201,I2859,I139839,I139804,);
DFFARX1 I_8079 (I140193,I2859,I139839,I139822,);
nor I_8080 (I140246,I558577,I558568);
not I_8081 (I140263,I140246);
nor I_8082 (I139825,I140102,I140263);
nand I_8083 (I139810,I140119,I140263);
nor I_8084 (I139819,I139865,I140246);
DFFARX1 I_8085 (I140246,I2859,I139839,I139828,);
not I_8086 (I140366,I2866);
DFFARX1 I_8087 (I47344,I2859,I140366,I140392,);
nand I_8088 (I140400,I47356,I47365);
and I_8089 (I140417,I140400,I47344);
DFFARX1 I_8090 (I140417,I2859,I140366,I140443,);
nor I_8091 (I140334,I140443,I140392);
not I_8092 (I140465,I140443);
DFFARX1 I_8093 (I47359,I2859,I140366,I140491,);
nand I_8094 (I140499,I140491,I47347);
not I_8095 (I140516,I140499);
DFFARX1 I_8096 (I140516,I2859,I140366,I140542,);
not I_8097 (I140358,I140542);
nor I_8098 (I140564,I140392,I140499);
nor I_8099 (I140340,I140443,I140564);
DFFARX1 I_8100 (I47350,I2859,I140366,I140604,);
DFFARX1 I_8101 (I140604,I2859,I140366,I140621,);
not I_8102 (I140629,I140621);
not I_8103 (I140646,I140604);
nand I_8104 (I140343,I140646,I140465);
nand I_8105 (I140677,I47341,I47341);
and I_8106 (I140694,I140677,I47353);
DFFARX1 I_8107 (I140694,I2859,I140366,I140720,);
nor I_8108 (I140728,I140720,I140392);
DFFARX1 I_8109 (I140728,I2859,I140366,I140331,);
DFFARX1 I_8110 (I140720,I2859,I140366,I140349,);
nor I_8111 (I140773,I47362,I47341);
not I_8112 (I140790,I140773);
nor I_8113 (I140352,I140629,I140790);
nand I_8114 (I140337,I140646,I140790);
nor I_8115 (I140346,I140392,I140773);
DFFARX1 I_8116 (I140773,I2859,I140366,I140355,);
not I_8117 (I140893,I2866);
DFFARX1 I_8118 (I252903,I2859,I140893,I140919,);
nand I_8119 (I140927,I252888,I252891);
and I_8120 (I140944,I140927,I252906);
DFFARX1 I_8121 (I140944,I2859,I140893,I140970,);
nor I_8122 (I140861,I140970,I140919);
not I_8123 (I140992,I140970);
DFFARX1 I_8124 (I252900,I2859,I140893,I141018,);
nand I_8125 (I141026,I141018,I252891);
not I_8126 (I141043,I141026);
DFFARX1 I_8127 (I141043,I2859,I140893,I141069,);
not I_8128 (I140885,I141069);
nor I_8129 (I141091,I140919,I141026);
nor I_8130 (I140867,I140970,I141091);
DFFARX1 I_8131 (I252897,I2859,I140893,I141131,);
DFFARX1 I_8132 (I141131,I2859,I140893,I141148,);
not I_8133 (I141156,I141148);
not I_8134 (I141173,I141131);
nand I_8135 (I140870,I141173,I140992);
nand I_8136 (I141204,I252912,I252888);
and I_8137 (I141221,I141204,I252909);
DFFARX1 I_8138 (I141221,I2859,I140893,I141247,);
nor I_8139 (I141255,I141247,I140919);
DFFARX1 I_8140 (I141255,I2859,I140893,I140858,);
DFFARX1 I_8141 (I141247,I2859,I140893,I140876,);
nor I_8142 (I141300,I252894,I252888);
not I_8143 (I141317,I141300);
nor I_8144 (I140879,I141156,I141317);
nand I_8145 (I140864,I141173,I141317);
nor I_8146 (I140873,I140919,I141300);
DFFARX1 I_8147 (I141300,I2859,I140893,I140882,);
not I_8148 (I141420,I2866);
DFFARX1 I_8149 (I55776,I2859,I141420,I141446,);
nand I_8150 (I141454,I55788,I55797);
and I_8151 (I141471,I141454,I55776);
DFFARX1 I_8152 (I141471,I2859,I141420,I141497,);
nor I_8153 (I141388,I141497,I141446);
not I_8154 (I141519,I141497);
DFFARX1 I_8155 (I55791,I2859,I141420,I141545,);
nand I_8156 (I141553,I141545,I55779);
not I_8157 (I141570,I141553);
DFFARX1 I_8158 (I141570,I2859,I141420,I141596,);
not I_8159 (I141412,I141596);
nor I_8160 (I141618,I141446,I141553);
nor I_8161 (I141394,I141497,I141618);
DFFARX1 I_8162 (I55782,I2859,I141420,I141658,);
DFFARX1 I_8163 (I141658,I2859,I141420,I141675,);
not I_8164 (I141683,I141675);
not I_8165 (I141700,I141658);
nand I_8166 (I141397,I141700,I141519);
nand I_8167 (I141731,I55773,I55773);
and I_8168 (I141748,I141731,I55785);
DFFARX1 I_8169 (I141748,I2859,I141420,I141774,);
nor I_8170 (I141782,I141774,I141446);
DFFARX1 I_8171 (I141782,I2859,I141420,I141385,);
DFFARX1 I_8172 (I141774,I2859,I141420,I141403,);
nor I_8173 (I141827,I55794,I55773);
not I_8174 (I141844,I141827);
nor I_8175 (I141406,I141683,I141844);
nand I_8176 (I141391,I141700,I141844);
nor I_8177 (I141400,I141446,I141827);
DFFARX1 I_8178 (I141827,I2859,I141420,I141409,);
not I_8179 (I141947,I2866);
DFFARX1 I_8180 (I76258,I2859,I141947,I141973,);
nand I_8181 (I141981,I76258,I76264);
and I_8182 (I141998,I141981,I76282);
DFFARX1 I_8183 (I141998,I2859,I141947,I142024,);
nor I_8184 (I141915,I142024,I141973);
not I_8185 (I142046,I142024);
DFFARX1 I_8186 (I76270,I2859,I141947,I142072,);
nand I_8187 (I142080,I142072,I76267);
not I_8188 (I142097,I142080);
DFFARX1 I_8189 (I142097,I2859,I141947,I142123,);
not I_8190 (I141939,I142123);
nor I_8191 (I142145,I141973,I142080);
nor I_8192 (I141921,I142024,I142145);
DFFARX1 I_8193 (I76276,I2859,I141947,I142185,);
DFFARX1 I_8194 (I142185,I2859,I141947,I142202,);
not I_8195 (I142210,I142202);
not I_8196 (I142227,I142185);
nand I_8197 (I141924,I142227,I142046);
nand I_8198 (I142258,I76261,I76261);
and I_8199 (I142275,I142258,I76273);
DFFARX1 I_8200 (I142275,I2859,I141947,I142301,);
nor I_8201 (I142309,I142301,I141973);
DFFARX1 I_8202 (I142309,I2859,I141947,I141912,);
DFFARX1 I_8203 (I142301,I2859,I141947,I141930,);
nor I_8204 (I142354,I76279,I76261);
not I_8205 (I142371,I142354);
nor I_8206 (I141933,I142210,I142371);
nand I_8207 (I141918,I142227,I142371);
nor I_8208 (I141927,I141973,I142354);
DFFARX1 I_8209 (I142354,I2859,I141947,I141936,);
not I_8210 (I142474,I2866);
DFFARX1 I_8211 (I31007,I2859,I142474,I142500,);
nand I_8212 (I142508,I31019,I31028);
and I_8213 (I142525,I142508,I31007);
DFFARX1 I_8214 (I142525,I2859,I142474,I142551,);
nor I_8215 (I142442,I142551,I142500);
not I_8216 (I142573,I142551);
DFFARX1 I_8217 (I31022,I2859,I142474,I142599,);
nand I_8218 (I142607,I142599,I31010);
not I_8219 (I142624,I142607);
DFFARX1 I_8220 (I142624,I2859,I142474,I142650,);
not I_8221 (I142466,I142650);
nor I_8222 (I142672,I142500,I142607);
nor I_8223 (I142448,I142551,I142672);
DFFARX1 I_8224 (I31013,I2859,I142474,I142712,);
DFFARX1 I_8225 (I142712,I2859,I142474,I142729,);
not I_8226 (I142737,I142729);
not I_8227 (I142754,I142712);
nand I_8228 (I142451,I142754,I142573);
nand I_8229 (I142785,I31004,I31004);
and I_8230 (I142802,I142785,I31016);
DFFARX1 I_8231 (I142802,I2859,I142474,I142828,);
nor I_8232 (I142836,I142828,I142500);
DFFARX1 I_8233 (I142836,I2859,I142474,I142439,);
DFFARX1 I_8234 (I142828,I2859,I142474,I142457,);
nor I_8235 (I142881,I31025,I31004);
not I_8236 (I142898,I142881);
nor I_8237 (I142460,I142737,I142898);
nand I_8238 (I142445,I142754,I142898);
nor I_8239 (I142454,I142500,I142881);
DFFARX1 I_8240 (I142881,I2859,I142474,I142463,);
not I_8241 (I143001,I2866);
DFFARX1 I_8242 (I185223,I2859,I143001,I143027,);
nand I_8243 (I143035,I185235,I185214);
and I_8244 (I143052,I143035,I185238);
DFFARX1 I_8245 (I143052,I2859,I143001,I143078,);
nor I_8246 (I142969,I143078,I143027);
not I_8247 (I143100,I143078);
DFFARX1 I_8248 (I185229,I2859,I143001,I143126,);
nand I_8249 (I143134,I143126,I185211);
not I_8250 (I143151,I143134);
DFFARX1 I_8251 (I143151,I2859,I143001,I143177,);
not I_8252 (I142993,I143177);
nor I_8253 (I143199,I143027,I143134);
nor I_8254 (I142975,I143078,I143199);
DFFARX1 I_8255 (I185226,I2859,I143001,I143239,);
DFFARX1 I_8256 (I143239,I2859,I143001,I143256,);
not I_8257 (I143264,I143256);
not I_8258 (I143281,I143239);
nand I_8259 (I142978,I143281,I143100);
nand I_8260 (I143312,I185211,I185217);
and I_8261 (I143329,I143312,I185220);
DFFARX1 I_8262 (I143329,I2859,I143001,I143355,);
nor I_8263 (I143363,I143355,I143027);
DFFARX1 I_8264 (I143363,I2859,I143001,I142966,);
DFFARX1 I_8265 (I143355,I2859,I143001,I142984,);
nor I_8266 (I143408,I185232,I185217);
not I_8267 (I143425,I143408);
nor I_8268 (I142987,I143264,I143425);
nand I_8269 (I142972,I143281,I143425);
nor I_8270 (I142981,I143027,I143408);
DFFARX1 I_8271 (I143408,I2859,I143001,I142990,);
not I_8272 (I143528,I2866);
DFFARX1 I_8273 (I172167,I2859,I143528,I143554,);
nand I_8274 (I143562,I172179,I172158);
and I_8275 (I143579,I143562,I172182);
DFFARX1 I_8276 (I143579,I2859,I143528,I143605,);
nor I_8277 (I143496,I143605,I143554);
not I_8278 (I143627,I143605);
DFFARX1 I_8279 (I172173,I2859,I143528,I143653,);
nand I_8280 (I143661,I143653,I172155);
not I_8281 (I143678,I143661);
DFFARX1 I_8282 (I143678,I2859,I143528,I143704,);
not I_8283 (I143520,I143704);
nor I_8284 (I143726,I143554,I143661);
nor I_8285 (I143502,I143605,I143726);
DFFARX1 I_8286 (I172170,I2859,I143528,I143766,);
DFFARX1 I_8287 (I143766,I2859,I143528,I143783,);
not I_8288 (I143791,I143783);
not I_8289 (I143808,I143766);
nand I_8290 (I143505,I143808,I143627);
nand I_8291 (I143839,I172155,I172161);
and I_8292 (I143856,I143839,I172164);
DFFARX1 I_8293 (I143856,I2859,I143528,I143882,);
nor I_8294 (I143890,I143882,I143554);
DFFARX1 I_8295 (I143890,I2859,I143528,I143493,);
DFFARX1 I_8296 (I143882,I2859,I143528,I143511,);
nor I_8297 (I143935,I172176,I172161);
not I_8298 (I143952,I143935);
nor I_8299 (I143514,I143791,I143952);
nand I_8300 (I143499,I143808,I143952);
nor I_8301 (I143508,I143554,I143935);
DFFARX1 I_8302 (I143935,I2859,I143528,I143517,);
not I_8303 (I144055,I2866);
DFFARX1 I_8304 (I432615,I2859,I144055,I144081,);
nand I_8305 (I144089,I432612,I432615);
and I_8306 (I144106,I144089,I432624);
DFFARX1 I_8307 (I144106,I2859,I144055,I144132,);
nor I_8308 (I144023,I144132,I144081);
not I_8309 (I144154,I144132);
DFFARX1 I_8310 (I432612,I2859,I144055,I144180,);
nand I_8311 (I144188,I144180,I432630);
not I_8312 (I144205,I144188);
DFFARX1 I_8313 (I144205,I2859,I144055,I144231,);
not I_8314 (I144047,I144231);
nor I_8315 (I144253,I144081,I144188);
nor I_8316 (I144029,I144132,I144253);
DFFARX1 I_8317 (I432618,I2859,I144055,I144293,);
DFFARX1 I_8318 (I144293,I2859,I144055,I144310,);
not I_8319 (I144318,I144310);
not I_8320 (I144335,I144293);
nand I_8321 (I144032,I144335,I144154);
nand I_8322 (I144366,I432627,I432633);
and I_8323 (I144383,I144366,I432618);
DFFARX1 I_8324 (I144383,I2859,I144055,I144409,);
nor I_8325 (I144417,I144409,I144081);
DFFARX1 I_8326 (I144417,I2859,I144055,I144020,);
DFFARX1 I_8327 (I144409,I2859,I144055,I144038,);
nor I_8328 (I144462,I432621,I432633);
not I_8329 (I144479,I144462);
nor I_8330 (I144041,I144318,I144479);
nand I_8331 (I144026,I144335,I144479);
nor I_8332 (I144035,I144081,I144462);
DFFARX1 I_8333 (I144462,I2859,I144055,I144044,);
not I_8334 (I144582,I2866);
DFFARX1 I_8335 (I563941,I2859,I144582,I144608,);
nand I_8336 (I144616,I563920,I563920);
and I_8337 (I144633,I144616,I563947);
DFFARX1 I_8338 (I144633,I2859,I144582,I144659,);
nor I_8339 (I144550,I144659,I144608);
not I_8340 (I144681,I144659);
DFFARX1 I_8341 (I563935,I2859,I144582,I144707,);
nand I_8342 (I144715,I144707,I563938);
not I_8343 (I144732,I144715);
DFFARX1 I_8344 (I144732,I2859,I144582,I144758,);
not I_8345 (I144574,I144758);
nor I_8346 (I144780,I144608,I144715);
nor I_8347 (I144556,I144659,I144780);
DFFARX1 I_8348 (I563929,I2859,I144582,I144820,);
DFFARX1 I_8349 (I144820,I2859,I144582,I144837,);
not I_8350 (I144845,I144837);
not I_8351 (I144862,I144820);
nand I_8352 (I144559,I144862,I144681);
nand I_8353 (I144893,I563926,I563923);
and I_8354 (I144910,I144893,I563944);
DFFARX1 I_8355 (I144910,I2859,I144582,I144936,);
nor I_8356 (I144944,I144936,I144608);
DFFARX1 I_8357 (I144944,I2859,I144582,I144547,);
DFFARX1 I_8358 (I144936,I2859,I144582,I144565,);
nor I_8359 (I144989,I563932,I563923);
not I_8360 (I145006,I144989);
nor I_8361 (I144568,I144845,I145006);
nand I_8362 (I144553,I144862,I145006);
nor I_8363 (I144562,I144608,I144989);
DFFARX1 I_8364 (I144989,I2859,I144582,I144571,);
not I_8365 (I145109,I2866);
DFFARX1 I_8366 (I299718,I2859,I145109,I145135,);
nand I_8367 (I145143,I299709,I299724);
and I_8368 (I145160,I145143,I299730);
DFFARX1 I_8369 (I145160,I2859,I145109,I145186,);
nor I_8370 (I145077,I145186,I145135);
not I_8371 (I145208,I145186);
DFFARX1 I_8372 (I299715,I2859,I145109,I145234,);
nand I_8373 (I145242,I145234,I299709);
not I_8374 (I145259,I145242);
DFFARX1 I_8375 (I145259,I2859,I145109,I145285,);
not I_8376 (I145101,I145285);
nor I_8377 (I145307,I145135,I145242);
nor I_8378 (I145083,I145186,I145307);
DFFARX1 I_8379 (I299712,I2859,I145109,I145347,);
DFFARX1 I_8380 (I145347,I2859,I145109,I145364,);
not I_8381 (I145372,I145364);
not I_8382 (I145389,I145347);
nand I_8383 (I145086,I145389,I145208);
nand I_8384 (I145420,I299706,I299721);
and I_8385 (I145437,I145420,I299706);
DFFARX1 I_8386 (I145437,I2859,I145109,I145463,);
nor I_8387 (I145471,I145463,I145135);
DFFARX1 I_8388 (I145471,I2859,I145109,I145074,);
DFFARX1 I_8389 (I145463,I2859,I145109,I145092,);
nor I_8390 (I145516,I299727,I299721);
not I_8391 (I145533,I145516);
nor I_8392 (I145095,I145372,I145533);
nand I_8393 (I145080,I145389,I145533);
nor I_8394 (I145089,I145135,I145516);
DFFARX1 I_8395 (I145516,I2859,I145109,I145098,);
not I_8396 (I145636,I2866);
DFFARX1 I_8397 (I52087,I2859,I145636,I145662,);
nand I_8398 (I145670,I52099,I52108);
and I_8399 (I145687,I145670,I52087);
DFFARX1 I_8400 (I145687,I2859,I145636,I145713,);
nor I_8401 (I145604,I145713,I145662);
not I_8402 (I145735,I145713);
DFFARX1 I_8403 (I52102,I2859,I145636,I145761,);
nand I_8404 (I145769,I145761,I52090);
not I_8405 (I145786,I145769);
DFFARX1 I_8406 (I145786,I2859,I145636,I145812,);
not I_8407 (I145628,I145812);
nor I_8408 (I145834,I145662,I145769);
nor I_8409 (I145610,I145713,I145834);
DFFARX1 I_8410 (I52093,I2859,I145636,I145874,);
DFFARX1 I_8411 (I145874,I2859,I145636,I145891,);
not I_8412 (I145899,I145891);
not I_8413 (I145916,I145874);
nand I_8414 (I145613,I145916,I145735);
nand I_8415 (I145947,I52084,I52084);
and I_8416 (I145964,I145947,I52096);
DFFARX1 I_8417 (I145964,I2859,I145636,I145990,);
nor I_8418 (I145998,I145990,I145662);
DFFARX1 I_8419 (I145998,I2859,I145636,I145601,);
DFFARX1 I_8420 (I145990,I2859,I145636,I145619,);
nor I_8421 (I146043,I52105,I52084);
not I_8422 (I146060,I146043);
nor I_8423 (I145622,I145899,I146060);
nand I_8424 (I145607,I145916,I146060);
nor I_8425 (I145616,I145662,I146043);
DFFARX1 I_8426 (I146043,I2859,I145636,I145625,);
not I_8427 (I146163,I2866);
DFFARX1 I_8428 (I96488,I2859,I146163,I146189,);
nand I_8429 (I146197,I96488,I96494);
and I_8430 (I146214,I146197,I96512);
DFFARX1 I_8431 (I146214,I2859,I146163,I146240,);
nor I_8432 (I146131,I146240,I146189);
not I_8433 (I146262,I146240);
DFFARX1 I_8434 (I96500,I2859,I146163,I146288,);
nand I_8435 (I146296,I146288,I96497);
not I_8436 (I146313,I146296);
DFFARX1 I_8437 (I146313,I2859,I146163,I146339,);
not I_8438 (I146155,I146339);
nor I_8439 (I146361,I146189,I146296);
nor I_8440 (I146137,I146240,I146361);
DFFARX1 I_8441 (I96506,I2859,I146163,I146401,);
DFFARX1 I_8442 (I146401,I2859,I146163,I146418,);
not I_8443 (I146426,I146418);
not I_8444 (I146443,I146401);
nand I_8445 (I146140,I146443,I146262);
nand I_8446 (I146474,I96491,I96491);
and I_8447 (I146491,I146474,I96503);
DFFARX1 I_8448 (I146491,I2859,I146163,I146517,);
nor I_8449 (I146525,I146517,I146189);
DFFARX1 I_8450 (I146525,I2859,I146163,I146128,);
DFFARX1 I_8451 (I146517,I2859,I146163,I146146,);
nor I_8452 (I146570,I96509,I96491);
not I_8453 (I146587,I146570);
nor I_8454 (I146149,I146426,I146587);
nand I_8455 (I146134,I146443,I146587);
nor I_8456 (I146143,I146189,I146570);
DFFARX1 I_8457 (I146570,I2859,I146163,I146152,);
not I_8458 (I146690,I2866);
DFFARX1 I_8459 (I405466,I2859,I146690,I146716,);
nand I_8460 (I146724,I405463,I405481);
and I_8461 (I146741,I146724,I405472);
DFFARX1 I_8462 (I146741,I2859,I146690,I146767,);
nor I_8463 (I146658,I146767,I146716);
not I_8464 (I146789,I146767);
DFFARX1 I_8465 (I405487,I2859,I146690,I146815,);
nand I_8466 (I146823,I146815,I405469);
not I_8467 (I146840,I146823);
DFFARX1 I_8468 (I146840,I2859,I146690,I146866,);
not I_8469 (I146682,I146866);
nor I_8470 (I146888,I146716,I146823);
nor I_8471 (I146664,I146767,I146888);
DFFARX1 I_8472 (I405475,I2859,I146690,I146928,);
DFFARX1 I_8473 (I146928,I2859,I146690,I146945,);
not I_8474 (I146953,I146945);
not I_8475 (I146970,I146928);
nand I_8476 (I146667,I146970,I146789);
nand I_8477 (I147001,I405463,I405490);
and I_8478 (I147018,I147001,I405478);
DFFARX1 I_8479 (I147018,I2859,I146690,I147044,);
nor I_8480 (I147052,I147044,I146716);
DFFARX1 I_8481 (I147052,I2859,I146690,I146655,);
DFFARX1 I_8482 (I147044,I2859,I146690,I146673,);
nor I_8483 (I147097,I405484,I405490);
not I_8484 (I147114,I147097);
nor I_8485 (I146676,I146953,I147114);
nand I_8486 (I146661,I146970,I147114);
nor I_8487 (I146670,I146716,I147097);
DFFARX1 I_8488 (I147097,I2859,I146690,I146679,);
not I_8489 (I147217,I2866);
DFFARX1 I_8490 (I552041,I2859,I147217,I147243,);
nand I_8491 (I147251,I552020,I552020);
and I_8492 (I147268,I147251,I552047);
DFFARX1 I_8493 (I147268,I2859,I147217,I147294,);
nor I_8494 (I147185,I147294,I147243);
not I_8495 (I147316,I147294);
DFFARX1 I_8496 (I552035,I2859,I147217,I147342,);
nand I_8497 (I147350,I147342,I552038);
not I_8498 (I147367,I147350);
DFFARX1 I_8499 (I147367,I2859,I147217,I147393,);
not I_8500 (I147209,I147393);
nor I_8501 (I147415,I147243,I147350);
nor I_8502 (I147191,I147294,I147415);
DFFARX1 I_8503 (I552029,I2859,I147217,I147455,);
DFFARX1 I_8504 (I147455,I2859,I147217,I147472,);
not I_8505 (I147480,I147472);
not I_8506 (I147497,I147455);
nand I_8507 (I147194,I147497,I147316);
nand I_8508 (I147528,I552026,I552023);
and I_8509 (I147545,I147528,I552044);
DFFARX1 I_8510 (I147545,I2859,I147217,I147571,);
nor I_8511 (I147579,I147571,I147243);
DFFARX1 I_8512 (I147579,I2859,I147217,I147182,);
DFFARX1 I_8513 (I147571,I2859,I147217,I147200,);
nor I_8514 (I147624,I552032,I552023);
not I_8515 (I147641,I147624);
nor I_8516 (I147203,I147480,I147641);
nand I_8517 (I147188,I147497,I147641);
nor I_8518 (I147197,I147243,I147624);
DFFARX1 I_8519 (I147624,I2859,I147217,I147206,);
not I_8520 (I147744,I2866);
DFFARX1 I_8521 (I200999,I2859,I147744,I147770,);
nand I_8522 (I147778,I201011,I200990);
and I_8523 (I147795,I147778,I201014);
DFFARX1 I_8524 (I147795,I2859,I147744,I147821,);
nor I_8525 (I147712,I147821,I147770);
not I_8526 (I147843,I147821);
DFFARX1 I_8527 (I201005,I2859,I147744,I147869,);
nand I_8528 (I147877,I147869,I200987);
not I_8529 (I147894,I147877);
DFFARX1 I_8530 (I147894,I2859,I147744,I147920,);
not I_8531 (I147736,I147920);
nor I_8532 (I147942,I147770,I147877);
nor I_8533 (I147718,I147821,I147942);
DFFARX1 I_8534 (I201002,I2859,I147744,I147982,);
DFFARX1 I_8535 (I147982,I2859,I147744,I147999,);
not I_8536 (I148007,I147999);
not I_8537 (I148024,I147982);
nand I_8538 (I147721,I148024,I147843);
nand I_8539 (I148055,I200987,I200993);
and I_8540 (I148072,I148055,I200996);
DFFARX1 I_8541 (I148072,I2859,I147744,I148098,);
nor I_8542 (I148106,I148098,I147770);
DFFARX1 I_8543 (I148106,I2859,I147744,I147709,);
DFFARX1 I_8544 (I148098,I2859,I147744,I147727,);
nor I_8545 (I148151,I201008,I200993);
not I_8546 (I148168,I148151);
nor I_8547 (I147730,I148007,I148168);
nand I_8548 (I147715,I148024,I148168);
nor I_8549 (I147724,I147770,I148151);
DFFARX1 I_8550 (I148151,I2859,I147744,I147733,);
not I_8551 (I148271,I2866);
DFFARX1 I_8552 (I206983,I2859,I148271,I148297,);
nand I_8553 (I148305,I206995,I206974);
and I_8554 (I148322,I148305,I206998);
DFFARX1 I_8555 (I148322,I2859,I148271,I148348,);
nor I_8556 (I148239,I148348,I148297);
not I_8557 (I148370,I148348);
DFFARX1 I_8558 (I206989,I2859,I148271,I148396,);
nand I_8559 (I148404,I148396,I206971);
not I_8560 (I148421,I148404);
DFFARX1 I_8561 (I148421,I2859,I148271,I148447,);
not I_8562 (I148263,I148447);
nor I_8563 (I148469,I148297,I148404);
nor I_8564 (I148245,I148348,I148469);
DFFARX1 I_8565 (I206986,I2859,I148271,I148509,);
DFFARX1 I_8566 (I148509,I2859,I148271,I148526,);
not I_8567 (I148534,I148526);
not I_8568 (I148551,I148509);
nand I_8569 (I148248,I148551,I148370);
nand I_8570 (I148582,I206971,I206977);
and I_8571 (I148599,I148582,I206980);
DFFARX1 I_8572 (I148599,I2859,I148271,I148625,);
nor I_8573 (I148633,I148625,I148297);
DFFARX1 I_8574 (I148633,I2859,I148271,I148236,);
DFFARX1 I_8575 (I148625,I2859,I148271,I148254,);
nor I_8576 (I148678,I206992,I206977);
not I_8577 (I148695,I148678);
nor I_8578 (I148257,I148534,I148695);
nand I_8579 (I148242,I148551,I148695);
nor I_8580 (I148251,I148297,I148678);
DFFARX1 I_8581 (I148678,I2859,I148271,I148260,);
not I_8582 (I148798,I2866);
DFFARX1 I_8583 (I487624,I2859,I148798,I148824,);
nand I_8584 (I148832,I487639,I487624);
and I_8585 (I148849,I148832,I487642);
DFFARX1 I_8586 (I148849,I2859,I148798,I148875,);
nor I_8587 (I148766,I148875,I148824);
not I_8588 (I148897,I148875);
DFFARX1 I_8589 (I487648,I2859,I148798,I148923,);
nand I_8590 (I148931,I148923,I487630);
not I_8591 (I148948,I148931);
DFFARX1 I_8592 (I148948,I2859,I148798,I148974,);
not I_8593 (I148790,I148974);
nor I_8594 (I148996,I148824,I148931);
nor I_8595 (I148772,I148875,I148996);
DFFARX1 I_8596 (I487627,I2859,I148798,I149036,);
DFFARX1 I_8597 (I149036,I2859,I148798,I149053,);
not I_8598 (I149061,I149053);
not I_8599 (I149078,I149036);
nand I_8600 (I148775,I149078,I148897);
nand I_8601 (I149109,I487627,I487633);
and I_8602 (I149126,I149109,I487645);
DFFARX1 I_8603 (I149126,I2859,I148798,I149152,);
nor I_8604 (I149160,I149152,I148824);
DFFARX1 I_8605 (I149160,I2859,I148798,I148763,);
DFFARX1 I_8606 (I149152,I2859,I148798,I148781,);
nor I_8607 (I149205,I487636,I487633);
not I_8608 (I149222,I149205);
nor I_8609 (I148784,I149061,I149222);
nand I_8610 (I148769,I149078,I149222);
nor I_8611 (I148778,I148824,I149205);
DFFARX1 I_8612 (I149205,I2859,I148798,I148787,);
not I_8613 (I149325,I2866);
DFFARX1 I_8614 (I27318,I2859,I149325,I149351,);
nand I_8615 (I149359,I27330,I27339);
and I_8616 (I149376,I149359,I27318);
DFFARX1 I_8617 (I149376,I2859,I149325,I149402,);
nor I_8618 (I149293,I149402,I149351);
not I_8619 (I149424,I149402);
DFFARX1 I_8620 (I27333,I2859,I149325,I149450,);
nand I_8621 (I149458,I149450,I27321);
not I_8622 (I149475,I149458);
DFFARX1 I_8623 (I149475,I2859,I149325,I149501,);
not I_8624 (I149317,I149501);
nor I_8625 (I149523,I149351,I149458);
nor I_8626 (I149299,I149402,I149523);
DFFARX1 I_8627 (I27324,I2859,I149325,I149563,);
DFFARX1 I_8628 (I149563,I2859,I149325,I149580,);
not I_8629 (I149588,I149580);
not I_8630 (I149605,I149563);
nand I_8631 (I149302,I149605,I149424);
nand I_8632 (I149636,I27315,I27315);
and I_8633 (I149653,I149636,I27327);
DFFARX1 I_8634 (I149653,I2859,I149325,I149679,);
nor I_8635 (I149687,I149679,I149351);
DFFARX1 I_8636 (I149687,I2859,I149325,I149290,);
DFFARX1 I_8637 (I149679,I2859,I149325,I149308,);
nor I_8638 (I149732,I27336,I27315);
not I_8639 (I149749,I149732);
nor I_8640 (I149311,I149588,I149749);
nand I_8641 (I149296,I149605,I149749);
nor I_8642 (I149305,I149351,I149732);
DFFARX1 I_8643 (I149732,I2859,I149325,I149314,);
not I_8644 (I149852,I2866);
DFFARX1 I_8645 (I95298,I2859,I149852,I149878,);
nand I_8646 (I149886,I95298,I95304);
and I_8647 (I149903,I149886,I95322);
DFFARX1 I_8648 (I149903,I2859,I149852,I149929,);
nor I_8649 (I149820,I149929,I149878);
not I_8650 (I149951,I149929);
DFFARX1 I_8651 (I95310,I2859,I149852,I149977,);
nand I_8652 (I149985,I149977,I95307);
not I_8653 (I150002,I149985);
DFFARX1 I_8654 (I150002,I2859,I149852,I150028,);
not I_8655 (I149844,I150028);
nor I_8656 (I150050,I149878,I149985);
nor I_8657 (I149826,I149929,I150050);
DFFARX1 I_8658 (I95316,I2859,I149852,I150090,);
DFFARX1 I_8659 (I150090,I2859,I149852,I150107,);
not I_8660 (I150115,I150107);
not I_8661 (I150132,I150090);
nand I_8662 (I149829,I150132,I149951);
nand I_8663 (I150163,I95301,I95301);
and I_8664 (I150180,I150163,I95313);
DFFARX1 I_8665 (I150180,I2859,I149852,I150206,);
nor I_8666 (I150214,I150206,I149878);
DFFARX1 I_8667 (I150214,I2859,I149852,I149817,);
DFFARX1 I_8668 (I150206,I2859,I149852,I149835,);
nor I_8669 (I150259,I95319,I95301);
not I_8670 (I150276,I150259);
nor I_8671 (I149838,I150115,I150276);
nand I_8672 (I149823,I150132,I150276);
nor I_8673 (I149832,I149878,I150259);
DFFARX1 I_8674 (I150259,I2859,I149852,I149841,);
not I_8675 (I150379,I2866);
DFFARX1 I_8676 (I410634,I2859,I150379,I150405,);
nand I_8677 (I150413,I410631,I410649);
and I_8678 (I150430,I150413,I410640);
DFFARX1 I_8679 (I150430,I2859,I150379,I150456,);
nor I_8680 (I150347,I150456,I150405);
not I_8681 (I150478,I150456);
DFFARX1 I_8682 (I410655,I2859,I150379,I150504,);
nand I_8683 (I150512,I150504,I410637);
not I_8684 (I150529,I150512);
DFFARX1 I_8685 (I150529,I2859,I150379,I150555,);
not I_8686 (I150371,I150555);
nor I_8687 (I150577,I150405,I150512);
nor I_8688 (I150353,I150456,I150577);
DFFARX1 I_8689 (I410643,I2859,I150379,I150617,);
DFFARX1 I_8690 (I150617,I2859,I150379,I150634,);
not I_8691 (I150642,I150634);
not I_8692 (I150659,I150617);
nand I_8693 (I150356,I150659,I150478);
nand I_8694 (I150690,I410631,I410658);
and I_8695 (I150707,I150690,I410646);
DFFARX1 I_8696 (I150707,I2859,I150379,I150733,);
nor I_8697 (I150741,I150733,I150405);
DFFARX1 I_8698 (I150741,I2859,I150379,I150344,);
DFFARX1 I_8699 (I150733,I2859,I150379,I150362,);
nor I_8700 (I150786,I410652,I410658);
not I_8701 (I150803,I150786);
nor I_8702 (I150365,I150642,I150803);
nand I_8703 (I150350,I150659,I150803);
nor I_8704 (I150359,I150405,I150786);
DFFARX1 I_8705 (I150786,I2859,I150379,I150368,);
not I_8706 (I150906,I2866);
DFFARX1 I_8707 (I490514,I2859,I150906,I150932,);
nand I_8708 (I150940,I490529,I490514);
and I_8709 (I150957,I150940,I490532);
DFFARX1 I_8710 (I150957,I2859,I150906,I150983,);
nor I_8711 (I150874,I150983,I150932);
not I_8712 (I151005,I150983);
DFFARX1 I_8713 (I490538,I2859,I150906,I151031,);
nand I_8714 (I151039,I151031,I490520);
not I_8715 (I151056,I151039);
DFFARX1 I_8716 (I151056,I2859,I150906,I151082,);
not I_8717 (I150898,I151082);
nor I_8718 (I151104,I150932,I151039);
nor I_8719 (I150880,I150983,I151104);
DFFARX1 I_8720 (I490517,I2859,I150906,I151144,);
DFFARX1 I_8721 (I151144,I2859,I150906,I151161,);
not I_8722 (I151169,I151161);
not I_8723 (I151186,I151144);
nand I_8724 (I150883,I151186,I151005);
nand I_8725 (I151217,I490517,I490523);
and I_8726 (I151234,I151217,I490535);
DFFARX1 I_8727 (I151234,I2859,I150906,I151260,);
nor I_8728 (I151268,I151260,I150932);
DFFARX1 I_8729 (I151268,I2859,I150906,I150871,);
DFFARX1 I_8730 (I151260,I2859,I150906,I150889,);
nor I_8731 (I151313,I490526,I490523);
not I_8732 (I151330,I151313);
nor I_8733 (I150892,I151169,I151330);
nand I_8734 (I150877,I151186,I151330);
nor I_8735 (I150886,I150932,I151313);
DFFARX1 I_8736 (I151313,I2859,I150906,I150895,);
not I_8737 (I151433,I2866);
DFFARX1 I_8738 (I239031,I2859,I151433,I151459,);
nand I_8739 (I151467,I239016,I239019);
and I_8740 (I151484,I151467,I239034);
DFFARX1 I_8741 (I151484,I2859,I151433,I151510,);
nor I_8742 (I151401,I151510,I151459);
not I_8743 (I151532,I151510);
DFFARX1 I_8744 (I239028,I2859,I151433,I151558,);
nand I_8745 (I151566,I151558,I239019);
not I_8746 (I151583,I151566);
DFFARX1 I_8747 (I151583,I2859,I151433,I151609,);
not I_8748 (I151425,I151609);
nor I_8749 (I151631,I151459,I151566);
nor I_8750 (I151407,I151510,I151631);
DFFARX1 I_8751 (I239025,I2859,I151433,I151671,);
DFFARX1 I_8752 (I151671,I2859,I151433,I151688,);
not I_8753 (I151696,I151688);
not I_8754 (I151713,I151671);
nand I_8755 (I151410,I151713,I151532);
nand I_8756 (I151744,I239040,I239016);
and I_8757 (I151761,I151744,I239037);
DFFARX1 I_8758 (I151761,I2859,I151433,I151787,);
nor I_8759 (I151795,I151787,I151459);
DFFARX1 I_8760 (I151795,I2859,I151433,I151398,);
DFFARX1 I_8761 (I151787,I2859,I151433,I151416,);
nor I_8762 (I151840,I239022,I239016);
not I_8763 (I151857,I151840);
nor I_8764 (I151419,I151696,I151857);
nand I_8765 (I151404,I151713,I151857);
nor I_8766 (I151413,I151459,I151840);
DFFARX1 I_8767 (I151840,I2859,I151433,I151422,);
not I_8768 (I151960,I2866);
DFFARX1 I_8769 (I269084,I2859,I151960,I151986,);
nand I_8770 (I151994,I269075,I269090);
and I_8771 (I152011,I151994,I269096);
DFFARX1 I_8772 (I152011,I2859,I151960,I152037,);
nor I_8773 (I151928,I152037,I151986);
not I_8774 (I152059,I152037);
DFFARX1 I_8775 (I269081,I2859,I151960,I152085,);
nand I_8776 (I152093,I152085,I269075);
not I_8777 (I152110,I152093);
DFFARX1 I_8778 (I152110,I2859,I151960,I152136,);
not I_8779 (I151952,I152136);
nor I_8780 (I152158,I151986,I152093);
nor I_8781 (I151934,I152037,I152158);
DFFARX1 I_8782 (I269078,I2859,I151960,I152198,);
DFFARX1 I_8783 (I152198,I2859,I151960,I152215,);
not I_8784 (I152223,I152215);
not I_8785 (I152240,I152198);
nand I_8786 (I151937,I152240,I152059);
nand I_8787 (I152271,I269072,I269087);
and I_8788 (I152288,I152271,I269072);
DFFARX1 I_8789 (I152288,I2859,I151960,I152314,);
nor I_8790 (I152322,I152314,I151986);
DFFARX1 I_8791 (I152322,I2859,I151960,I151925,);
DFFARX1 I_8792 (I152314,I2859,I151960,I151943,);
nor I_8793 (I152367,I269093,I269087);
not I_8794 (I152384,I152367);
nor I_8795 (I151946,I152223,I152384);
nand I_8796 (I151931,I152240,I152384);
nor I_8797 (I151940,I151986,I152367);
DFFARX1 I_8798 (I152367,I2859,I151960,I151949,);
not I_8799 (I152487,I2866);
DFFARX1 I_8800 (I563346,I2859,I152487,I152513,);
nand I_8801 (I152521,I563325,I563325);
and I_8802 (I152538,I152521,I563352);
DFFARX1 I_8803 (I152538,I2859,I152487,I152564,);
nor I_8804 (I152455,I152564,I152513);
not I_8805 (I152586,I152564);
DFFARX1 I_8806 (I563340,I2859,I152487,I152612,);
nand I_8807 (I152620,I152612,I563343);
not I_8808 (I152637,I152620);
DFFARX1 I_8809 (I152637,I2859,I152487,I152663,);
not I_8810 (I152479,I152663);
nor I_8811 (I152685,I152513,I152620);
nor I_8812 (I152461,I152564,I152685);
DFFARX1 I_8813 (I563334,I2859,I152487,I152725,);
DFFARX1 I_8814 (I152725,I2859,I152487,I152742,);
not I_8815 (I152750,I152742);
not I_8816 (I152767,I152725);
nand I_8817 (I152464,I152767,I152586);
nand I_8818 (I152798,I563331,I563328);
and I_8819 (I152815,I152798,I563349);
DFFARX1 I_8820 (I152815,I2859,I152487,I152841,);
nor I_8821 (I152849,I152841,I152513);
DFFARX1 I_8822 (I152849,I2859,I152487,I152452,);
DFFARX1 I_8823 (I152841,I2859,I152487,I152470,);
nor I_8824 (I152894,I563337,I563328);
not I_8825 (I152911,I152894);
nor I_8826 (I152473,I152750,I152911);
nand I_8827 (I152458,I152767,I152911);
nor I_8828 (I152467,I152513,I152894);
DFFARX1 I_8829 (I152894,I2859,I152487,I152476,);
not I_8830 (I153014,I2866);
DFFARX1 I_8831 (I480110,I2859,I153014,I153040,);
nand I_8832 (I153048,I480125,I480110);
and I_8833 (I153065,I153048,I480128);
DFFARX1 I_8834 (I153065,I2859,I153014,I153091,);
nor I_8835 (I152982,I153091,I153040);
not I_8836 (I153113,I153091);
DFFARX1 I_8837 (I480134,I2859,I153014,I153139,);
nand I_8838 (I153147,I153139,I480116);
not I_8839 (I153164,I153147);
DFFARX1 I_8840 (I153164,I2859,I153014,I153190,);
not I_8841 (I153006,I153190);
nor I_8842 (I153212,I153040,I153147);
nor I_8843 (I152988,I153091,I153212);
DFFARX1 I_8844 (I480113,I2859,I153014,I153252,);
DFFARX1 I_8845 (I153252,I2859,I153014,I153269,);
not I_8846 (I153277,I153269);
not I_8847 (I153294,I153252);
nand I_8848 (I152991,I153294,I153113);
nand I_8849 (I153325,I480113,I480119);
and I_8850 (I153342,I153325,I480131);
DFFARX1 I_8851 (I153342,I2859,I153014,I153368,);
nor I_8852 (I153376,I153368,I153040);
DFFARX1 I_8853 (I153376,I2859,I153014,I152979,);
DFFARX1 I_8854 (I153368,I2859,I153014,I152997,);
nor I_8855 (I153421,I480122,I480119);
not I_8856 (I153438,I153421);
nor I_8857 (I153000,I153277,I153438);
nand I_8858 (I152985,I153294,I153438);
nor I_8859 (I152994,I153040,I153421);
DFFARX1 I_8860 (I153421,I2859,I153014,I153003,);
not I_8861 (I153541,I2866);
DFFARX1 I_8862 (I165639,I2859,I153541,I153567,);
nand I_8863 (I153575,I165651,I165630);
and I_8864 (I153592,I153575,I165654);
DFFARX1 I_8865 (I153592,I2859,I153541,I153618,);
nor I_8866 (I153509,I153618,I153567);
not I_8867 (I153640,I153618);
DFFARX1 I_8868 (I165645,I2859,I153541,I153666,);
nand I_8869 (I153674,I153666,I165627);
not I_8870 (I153691,I153674);
DFFARX1 I_8871 (I153691,I2859,I153541,I153717,);
not I_8872 (I153533,I153717);
nor I_8873 (I153739,I153567,I153674);
nor I_8874 (I153515,I153618,I153739);
DFFARX1 I_8875 (I165642,I2859,I153541,I153779,);
DFFARX1 I_8876 (I153779,I2859,I153541,I153796,);
not I_8877 (I153804,I153796);
not I_8878 (I153821,I153779);
nand I_8879 (I153518,I153821,I153640);
nand I_8880 (I153852,I165627,I165633);
and I_8881 (I153869,I153852,I165636);
DFFARX1 I_8882 (I153869,I2859,I153541,I153895,);
nor I_8883 (I153903,I153895,I153567);
DFFARX1 I_8884 (I153903,I2859,I153541,I153506,);
DFFARX1 I_8885 (I153895,I2859,I153541,I153524,);
nor I_8886 (I153948,I165648,I165633);
not I_8887 (I153965,I153948);
nor I_8888 (I153527,I153804,I153965);
nand I_8889 (I153512,I153821,I153965);
nor I_8890 (I153521,I153567,I153948);
DFFARX1 I_8891 (I153948,I2859,I153541,I153530,);
not I_8892 (I154068,I2866);
DFFARX1 I_8893 (I184135,I2859,I154068,I154094,);
nand I_8894 (I154102,I184147,I184126);
and I_8895 (I154119,I154102,I184150);
DFFARX1 I_8896 (I154119,I2859,I154068,I154145,);
nor I_8897 (I154036,I154145,I154094);
not I_8898 (I154167,I154145);
DFFARX1 I_8899 (I184141,I2859,I154068,I154193,);
nand I_8900 (I154201,I154193,I184123);
not I_8901 (I154218,I154201);
DFFARX1 I_8902 (I154218,I2859,I154068,I154244,);
not I_8903 (I154060,I154244);
nor I_8904 (I154266,I154094,I154201);
nor I_8905 (I154042,I154145,I154266);
DFFARX1 I_8906 (I184138,I2859,I154068,I154306,);
DFFARX1 I_8907 (I154306,I2859,I154068,I154323,);
not I_8908 (I154331,I154323);
not I_8909 (I154348,I154306);
nand I_8910 (I154045,I154348,I154167);
nand I_8911 (I154379,I184123,I184129);
and I_8912 (I154396,I154379,I184132);
DFFARX1 I_8913 (I154396,I2859,I154068,I154422,);
nor I_8914 (I154430,I154422,I154094);
DFFARX1 I_8915 (I154430,I2859,I154068,I154033,);
DFFARX1 I_8916 (I154422,I2859,I154068,I154051,);
nor I_8917 (I154475,I184144,I184129);
not I_8918 (I154492,I154475);
nor I_8919 (I154054,I154331,I154492);
nand I_8920 (I154039,I154348,I154492);
nor I_8921 (I154048,I154094,I154475);
DFFARX1 I_8922 (I154475,I2859,I154068,I154057,);
not I_8923 (I154595,I2866);
DFFARX1 I_8924 (I242499,I2859,I154595,I154621,);
nand I_8925 (I154629,I242484,I242487);
and I_8926 (I154646,I154629,I242502);
DFFARX1 I_8927 (I154646,I2859,I154595,I154672,);
nor I_8928 (I154563,I154672,I154621);
not I_8929 (I154694,I154672);
DFFARX1 I_8930 (I242496,I2859,I154595,I154720,);
nand I_8931 (I154728,I154720,I242487);
not I_8932 (I154745,I154728);
DFFARX1 I_8933 (I154745,I2859,I154595,I154771,);
not I_8934 (I154587,I154771);
nor I_8935 (I154793,I154621,I154728);
nor I_8936 (I154569,I154672,I154793);
DFFARX1 I_8937 (I242493,I2859,I154595,I154833,);
DFFARX1 I_8938 (I154833,I2859,I154595,I154850,);
not I_8939 (I154858,I154850);
not I_8940 (I154875,I154833);
nand I_8941 (I154572,I154875,I154694);
nand I_8942 (I154906,I242508,I242484);
and I_8943 (I154923,I154906,I242505);
DFFARX1 I_8944 (I154923,I2859,I154595,I154949,);
nor I_8945 (I154957,I154949,I154621);
DFFARX1 I_8946 (I154957,I2859,I154595,I154560,);
DFFARX1 I_8947 (I154949,I2859,I154595,I154578,);
nor I_8948 (I155002,I242490,I242484);
not I_8949 (I155019,I155002);
nor I_8950 (I154581,I154858,I155019);
nand I_8951 (I154566,I154875,I155019);
nor I_8952 (I154575,I154621,I155002);
DFFARX1 I_8953 (I155002,I2859,I154595,I154584,);
not I_8954 (I155122,I2866);
DFFARX1 I_8955 (I370599,I2859,I155122,I155148,);
nand I_8956 (I155156,I370602,I370596);
and I_8957 (I155173,I155156,I370608);
DFFARX1 I_8958 (I155173,I2859,I155122,I155199,);
nor I_8959 (I155090,I155199,I155148);
not I_8960 (I155221,I155199);
DFFARX1 I_8961 (I370611,I2859,I155122,I155247,);
nand I_8962 (I155255,I155247,I370602);
not I_8963 (I155272,I155255);
DFFARX1 I_8964 (I155272,I2859,I155122,I155298,);
not I_8965 (I155114,I155298);
nor I_8966 (I155320,I155148,I155255);
nor I_8967 (I155096,I155199,I155320);
DFFARX1 I_8968 (I370614,I2859,I155122,I155360,);
DFFARX1 I_8969 (I155360,I2859,I155122,I155377,);
not I_8970 (I155385,I155377);
not I_8971 (I155402,I155360);
nand I_8972 (I155099,I155402,I155221);
nand I_8973 (I155433,I370596,I370605);
and I_8974 (I155450,I155433,I370599);
DFFARX1 I_8975 (I155450,I2859,I155122,I155476,);
nor I_8976 (I155484,I155476,I155148);
DFFARX1 I_8977 (I155484,I2859,I155122,I155087,);
DFFARX1 I_8978 (I155476,I2859,I155122,I155105,);
nor I_8979 (I155529,I370617,I370605);
not I_8980 (I155546,I155529);
nor I_8981 (I155108,I155385,I155546);
nand I_8982 (I155093,I155402,I155546);
nor I_8983 (I155102,I155148,I155529);
DFFARX1 I_8984 (I155529,I2859,I155122,I155111,);
not I_8985 (I155649,I2866);
DFFARX1 I_8986 (I269662,I2859,I155649,I155675,);
nand I_8987 (I155683,I269653,I269668);
and I_8988 (I155700,I155683,I269674);
DFFARX1 I_8989 (I155700,I2859,I155649,I155726,);
nor I_8990 (I155617,I155726,I155675);
not I_8991 (I155748,I155726);
DFFARX1 I_8992 (I269659,I2859,I155649,I155774,);
nand I_8993 (I155782,I155774,I269653);
not I_8994 (I155799,I155782);
DFFARX1 I_8995 (I155799,I2859,I155649,I155825,);
not I_8996 (I155641,I155825);
nor I_8997 (I155847,I155675,I155782);
nor I_8998 (I155623,I155726,I155847);
DFFARX1 I_8999 (I269656,I2859,I155649,I155887,);
DFFARX1 I_9000 (I155887,I2859,I155649,I155904,);
not I_9001 (I155912,I155904);
not I_9002 (I155929,I155887);
nand I_9003 (I155626,I155929,I155748);
nand I_9004 (I155960,I269650,I269665);
and I_9005 (I155977,I155960,I269650);
DFFARX1 I_9006 (I155977,I2859,I155649,I156003,);
nor I_9007 (I156011,I156003,I155675);
DFFARX1 I_9008 (I156011,I2859,I155649,I155614,);
DFFARX1 I_9009 (I156003,I2859,I155649,I155632,);
nor I_9010 (I156056,I269671,I269665);
not I_9011 (I156073,I156056);
nor I_9012 (I155635,I155912,I156073);
nand I_9013 (I155620,I155929,I156073);
nor I_9014 (I155629,I155675,I156056);
DFFARX1 I_9015 (I156056,I2859,I155649,I155638,);
not I_9016 (I156176,I2866);
DFFARX1 I_9017 (I461036,I2859,I156176,I156202,);
nand I_9018 (I156210,I461051,I461036);
and I_9019 (I156227,I156210,I461054);
DFFARX1 I_9020 (I156227,I2859,I156176,I156253,);
nor I_9021 (I156144,I156253,I156202);
not I_9022 (I156275,I156253);
DFFARX1 I_9023 (I461060,I2859,I156176,I156301,);
nand I_9024 (I156309,I156301,I461042);
not I_9025 (I156326,I156309);
DFFARX1 I_9026 (I156326,I2859,I156176,I156352,);
not I_9027 (I156168,I156352);
nor I_9028 (I156374,I156202,I156309);
nor I_9029 (I156150,I156253,I156374);
DFFARX1 I_9030 (I461039,I2859,I156176,I156414,);
DFFARX1 I_9031 (I156414,I2859,I156176,I156431,);
not I_9032 (I156439,I156431);
not I_9033 (I156456,I156414);
nand I_9034 (I156153,I156456,I156275);
nand I_9035 (I156487,I461039,I461045);
and I_9036 (I156504,I156487,I461057);
DFFARX1 I_9037 (I156504,I2859,I156176,I156530,);
nor I_9038 (I156538,I156530,I156202);
DFFARX1 I_9039 (I156538,I2859,I156176,I156141,);
DFFARX1 I_9040 (I156530,I2859,I156176,I156159,);
nor I_9041 (I156583,I461048,I461045);
not I_9042 (I156600,I156583);
nor I_9043 (I156162,I156439,I156600);
nand I_9044 (I156147,I156456,I156600);
nor I_9045 (I156156,I156202,I156583);
DFFARX1 I_9046 (I156583,I2859,I156176,I156165,);
not I_9047 (I156703,I2866);
DFFARX1 I_9048 (I498606,I2859,I156703,I156729,);
nand I_9049 (I156737,I498621,I498606);
and I_9050 (I156754,I156737,I498624);
DFFARX1 I_9051 (I156754,I2859,I156703,I156780,);
nor I_9052 (I156671,I156780,I156729);
not I_9053 (I156802,I156780);
DFFARX1 I_9054 (I498630,I2859,I156703,I156828,);
nand I_9055 (I156836,I156828,I498612);
not I_9056 (I156853,I156836);
DFFARX1 I_9057 (I156853,I2859,I156703,I156879,);
not I_9058 (I156695,I156879);
nor I_9059 (I156901,I156729,I156836);
nor I_9060 (I156677,I156780,I156901);
DFFARX1 I_9061 (I498609,I2859,I156703,I156941,);
DFFARX1 I_9062 (I156941,I2859,I156703,I156958,);
not I_9063 (I156966,I156958);
not I_9064 (I156983,I156941);
nand I_9065 (I156680,I156983,I156802);
nand I_9066 (I157014,I498609,I498615);
and I_9067 (I157031,I157014,I498627);
DFFARX1 I_9068 (I157031,I2859,I156703,I157057,);
nor I_9069 (I157065,I157057,I156729);
DFFARX1 I_9070 (I157065,I2859,I156703,I156668,);
DFFARX1 I_9071 (I157057,I2859,I156703,I156686,);
nor I_9072 (I157110,I498618,I498615);
not I_9073 (I157127,I157110);
nor I_9074 (I156689,I156966,I157127);
nand I_9075 (I156674,I156983,I157127);
nor I_9076 (I156683,I156729,I157110);
DFFARX1 I_9077 (I157110,I2859,I156703,I156692,);
not I_9078 (I157230,I2866);
DFFARX1 I_9079 (I515148,I2859,I157230,I157256,);
nand I_9080 (I157264,I515130,I515154);
and I_9081 (I157281,I157264,I515145);
DFFARX1 I_9082 (I157281,I2859,I157230,I157307,);
nor I_9083 (I157198,I157307,I157256);
not I_9084 (I157329,I157307);
DFFARX1 I_9085 (I515151,I2859,I157230,I157355,);
nand I_9086 (I157363,I157355,I515139);
not I_9087 (I157380,I157363);
DFFARX1 I_9088 (I157380,I2859,I157230,I157406,);
not I_9089 (I157222,I157406);
nor I_9090 (I157428,I157256,I157363);
nor I_9091 (I157204,I157307,I157428);
DFFARX1 I_9092 (I515130,I2859,I157230,I157468,);
DFFARX1 I_9093 (I157468,I2859,I157230,I157485,);
not I_9094 (I157493,I157485);
not I_9095 (I157510,I157468);
nand I_9096 (I157207,I157510,I157329);
nand I_9097 (I157541,I515136,I515133);
and I_9098 (I157558,I157541,I515142);
DFFARX1 I_9099 (I157558,I2859,I157230,I157584,);
nor I_9100 (I157592,I157584,I157256);
DFFARX1 I_9101 (I157592,I2859,I157230,I157195,);
DFFARX1 I_9102 (I157584,I2859,I157230,I157213,);
nor I_9103 (I157637,I515133,I515133);
not I_9104 (I157654,I157637);
nor I_9105 (I157216,I157493,I157654);
nand I_9106 (I157201,I157510,I157654);
nor I_9107 (I157210,I157256,I157637);
DFFARX1 I_9108 (I157637,I2859,I157230,I157219,);
not I_9109 (I157757,I2866);
DFFARX1 I_9110 (I87563,I2859,I157757,I157783,);
nand I_9111 (I157791,I87563,I87569);
and I_9112 (I157808,I157791,I87587);
DFFARX1 I_9113 (I157808,I2859,I157757,I157834,);
nor I_9114 (I157725,I157834,I157783);
not I_9115 (I157856,I157834);
DFFARX1 I_9116 (I87575,I2859,I157757,I157882,);
nand I_9117 (I157890,I157882,I87572);
not I_9118 (I157907,I157890);
DFFARX1 I_9119 (I157907,I2859,I157757,I157933,);
not I_9120 (I157749,I157933);
nor I_9121 (I157955,I157783,I157890);
nor I_9122 (I157731,I157834,I157955);
DFFARX1 I_9123 (I87581,I2859,I157757,I157995,);
DFFARX1 I_9124 (I157995,I2859,I157757,I158012,);
not I_9125 (I158020,I158012);
not I_9126 (I158037,I157995);
nand I_9127 (I157734,I158037,I157856);
nand I_9128 (I158068,I87566,I87566);
and I_9129 (I158085,I158068,I87578);
DFFARX1 I_9130 (I158085,I2859,I157757,I158111,);
nor I_9131 (I158119,I158111,I157783);
DFFARX1 I_9132 (I158119,I2859,I157757,I157722,);
DFFARX1 I_9133 (I158111,I2859,I157757,I157740,);
nor I_9134 (I158164,I87584,I87566);
not I_9135 (I158181,I158164);
nor I_9136 (I157743,I158020,I158181);
nand I_9137 (I157728,I158037,I158181);
nor I_9138 (I157737,I157783,I158164);
DFFARX1 I_9139 (I158164,I2859,I157757,I157746,);
not I_9140 (I158284,I2866);
DFFARX1 I_9141 (I425883,I2859,I158284,I158310,);
nand I_9142 (I158318,I425880,I425883);
and I_9143 (I158335,I158318,I425892);
DFFARX1 I_9144 (I158335,I2859,I158284,I158361,);
nor I_9145 (I158252,I158361,I158310);
not I_9146 (I158383,I158361);
DFFARX1 I_9147 (I425880,I2859,I158284,I158409,);
nand I_9148 (I158417,I158409,I425898);
not I_9149 (I158434,I158417);
DFFARX1 I_9150 (I158434,I2859,I158284,I158460,);
not I_9151 (I158276,I158460);
nor I_9152 (I158482,I158310,I158417);
nor I_9153 (I158258,I158361,I158482);
DFFARX1 I_9154 (I425886,I2859,I158284,I158522,);
DFFARX1 I_9155 (I158522,I2859,I158284,I158539,);
not I_9156 (I158547,I158539);
not I_9157 (I158564,I158522);
nand I_9158 (I158261,I158564,I158383);
nand I_9159 (I158595,I425895,I425901);
and I_9160 (I158612,I158595,I425886);
DFFARX1 I_9161 (I158612,I2859,I158284,I158638,);
nor I_9162 (I158646,I158638,I158310);
DFFARX1 I_9163 (I158646,I2859,I158284,I158249,);
DFFARX1 I_9164 (I158638,I2859,I158284,I158267,);
nor I_9165 (I158691,I425889,I425901);
not I_9166 (I158708,I158691);
nor I_9167 (I158270,I158547,I158708);
nand I_9168 (I158255,I158564,I158708);
nor I_9169 (I158264,I158310,I158691);
DFFARX1 I_9170 (I158691,I2859,I158284,I158273,);
not I_9171 (I158811,I2866);
DFFARX1 I_9172 (I422262,I2859,I158811,I158837,);
nand I_9173 (I158845,I422259,I422277);
and I_9174 (I158862,I158845,I422268);
DFFARX1 I_9175 (I158862,I2859,I158811,I158888,);
nor I_9176 (I158779,I158888,I158837);
not I_9177 (I158910,I158888);
DFFARX1 I_9178 (I422283,I2859,I158811,I158936,);
nand I_9179 (I158944,I158936,I422265);
not I_9180 (I158961,I158944);
DFFARX1 I_9181 (I158961,I2859,I158811,I158987,);
not I_9182 (I158803,I158987);
nor I_9183 (I159009,I158837,I158944);
nor I_9184 (I158785,I158888,I159009);
DFFARX1 I_9185 (I422271,I2859,I158811,I159049,);
DFFARX1 I_9186 (I159049,I2859,I158811,I159066,);
not I_9187 (I159074,I159066);
not I_9188 (I159091,I159049);
nand I_9189 (I158788,I159091,I158910);
nand I_9190 (I159122,I422259,I422286);
and I_9191 (I159139,I159122,I422274);
DFFARX1 I_9192 (I159139,I2859,I158811,I159165,);
nor I_9193 (I159173,I159165,I158837);
DFFARX1 I_9194 (I159173,I2859,I158811,I158776,);
DFFARX1 I_9195 (I159165,I2859,I158811,I158794,);
nor I_9196 (I159218,I422280,I422286);
not I_9197 (I159235,I159218);
nor I_9198 (I158797,I159074,I159235);
nand I_9199 (I158782,I159091,I159235);
nor I_9200 (I158791,I158837,I159218);
DFFARX1 I_9201 (I159218,I2859,I158811,I158800,);
not I_9202 (I159338,I2866);
DFFARX1 I_9203 (I477798,I2859,I159338,I159364,);
nand I_9204 (I159372,I477813,I477798);
and I_9205 (I159389,I159372,I477816);
DFFARX1 I_9206 (I159389,I2859,I159338,I159415,);
nor I_9207 (I159306,I159415,I159364);
not I_9208 (I159437,I159415);
DFFARX1 I_9209 (I477822,I2859,I159338,I159463,);
nand I_9210 (I159471,I159463,I477804);
not I_9211 (I159488,I159471);
DFFARX1 I_9212 (I159488,I2859,I159338,I159514,);
not I_9213 (I159330,I159514);
nor I_9214 (I159536,I159364,I159471);
nor I_9215 (I159312,I159415,I159536);
DFFARX1 I_9216 (I477801,I2859,I159338,I159576,);
DFFARX1 I_9217 (I159576,I2859,I159338,I159593,);
not I_9218 (I159601,I159593);
not I_9219 (I159618,I159576);
nand I_9220 (I159315,I159618,I159437);
nand I_9221 (I159649,I477801,I477807);
and I_9222 (I159666,I159649,I477819);
DFFARX1 I_9223 (I159666,I2859,I159338,I159692,);
nor I_9224 (I159700,I159692,I159364);
DFFARX1 I_9225 (I159700,I2859,I159338,I159303,);
DFFARX1 I_9226 (I159692,I2859,I159338,I159321,);
nor I_9227 (I159745,I477810,I477807);
not I_9228 (I159762,I159745);
nor I_9229 (I159324,I159601,I159762);
nand I_9230 (I159309,I159618,I159762);
nor I_9231 (I159318,I159364,I159745);
DFFARX1 I_9232 (I159745,I2859,I159338,I159327,);
not I_9233 (I159865,I2866);
DFFARX1 I_9234 (I404820,I2859,I159865,I159891,);
nand I_9235 (I159899,I404817,I404835);
and I_9236 (I159916,I159899,I404826);
DFFARX1 I_9237 (I159916,I2859,I159865,I159942,);
nor I_9238 (I159833,I159942,I159891);
not I_9239 (I159964,I159942);
DFFARX1 I_9240 (I404841,I2859,I159865,I159990,);
nand I_9241 (I159998,I159990,I404823);
not I_9242 (I160015,I159998);
DFFARX1 I_9243 (I160015,I2859,I159865,I160041,);
not I_9244 (I159857,I160041);
nor I_9245 (I160063,I159891,I159998);
nor I_9246 (I159839,I159942,I160063);
DFFARX1 I_9247 (I404829,I2859,I159865,I160103,);
DFFARX1 I_9248 (I160103,I2859,I159865,I160120,);
not I_9249 (I160128,I160120);
not I_9250 (I160145,I160103);
nand I_9251 (I159842,I160145,I159964);
nand I_9252 (I160176,I404817,I404844);
and I_9253 (I160193,I160176,I404832);
DFFARX1 I_9254 (I160193,I2859,I159865,I160219,);
nor I_9255 (I160227,I160219,I159891);
DFFARX1 I_9256 (I160227,I2859,I159865,I159830,);
DFFARX1 I_9257 (I160219,I2859,I159865,I159848,);
nor I_9258 (I160272,I404838,I404844);
not I_9259 (I160289,I160272);
nor I_9260 (I159851,I160128,I160289);
nand I_9261 (I159836,I160145,I160289);
nor I_9262 (I159845,I159891,I160272);
DFFARX1 I_9263 (I160272,I2859,I159865,I159854,);
not I_9264 (I160392,I2866);
DFFARX1 I_9265 (I372180,I2859,I160392,I160418,);
nand I_9266 (I160426,I372183,I372177);
and I_9267 (I160443,I160426,I372189);
DFFARX1 I_9268 (I160443,I2859,I160392,I160469,);
nor I_9269 (I160360,I160469,I160418);
not I_9270 (I160491,I160469);
DFFARX1 I_9271 (I372192,I2859,I160392,I160517,);
nand I_9272 (I160525,I160517,I372183);
not I_9273 (I160542,I160525);
DFFARX1 I_9274 (I160542,I2859,I160392,I160568,);
not I_9275 (I160384,I160568);
nor I_9276 (I160590,I160418,I160525);
nor I_9277 (I160366,I160469,I160590);
DFFARX1 I_9278 (I372195,I2859,I160392,I160630,);
DFFARX1 I_9279 (I160630,I2859,I160392,I160647,);
not I_9280 (I160655,I160647);
not I_9281 (I160672,I160630);
nand I_9282 (I160369,I160672,I160491);
nand I_9283 (I160703,I372177,I372186);
and I_9284 (I160720,I160703,I372180);
DFFARX1 I_9285 (I160720,I2859,I160392,I160746,);
nor I_9286 (I160754,I160746,I160418);
DFFARX1 I_9287 (I160754,I2859,I160392,I160357,);
DFFARX1 I_9288 (I160746,I2859,I160392,I160375,);
nor I_9289 (I160799,I372198,I372186);
not I_9290 (I160816,I160799);
nor I_9291 (I160378,I160655,I160816);
nand I_9292 (I160363,I160672,I160816);
nor I_9293 (I160372,I160418,I160799);
DFFARX1 I_9294 (I160799,I2859,I160392,I160381,);
not I_9295 (I160919,I2866);
DFFARX1 I_9296 (I296828,I2859,I160919,I160945,);
nand I_9297 (I160953,I296819,I296834);
and I_9298 (I160970,I160953,I296840);
DFFARX1 I_9299 (I160970,I2859,I160919,I160996,);
nor I_9300 (I160887,I160996,I160945);
not I_9301 (I161018,I160996);
DFFARX1 I_9302 (I296825,I2859,I160919,I161044,);
nand I_9303 (I161052,I161044,I296819);
not I_9304 (I161069,I161052);
DFFARX1 I_9305 (I161069,I2859,I160919,I161095,);
not I_9306 (I160911,I161095);
nor I_9307 (I161117,I160945,I161052);
nor I_9308 (I160893,I160996,I161117);
DFFARX1 I_9309 (I296822,I2859,I160919,I161157,);
DFFARX1 I_9310 (I161157,I2859,I160919,I161174,);
not I_9311 (I161182,I161174);
not I_9312 (I161199,I161157);
nand I_9313 (I160896,I161199,I161018);
nand I_9314 (I161230,I296816,I296831);
and I_9315 (I161247,I161230,I296816);
DFFARX1 I_9316 (I161247,I2859,I160919,I161273,);
nor I_9317 (I161281,I161273,I160945);
DFFARX1 I_9318 (I161281,I2859,I160919,I160884,);
DFFARX1 I_9319 (I161273,I2859,I160919,I160902,);
nor I_9320 (I161326,I296837,I296831);
not I_9321 (I161343,I161326);
nor I_9322 (I160905,I161182,I161343);
nand I_9323 (I160890,I161199,I161343);
nor I_9324 (I160899,I160945,I161326);
DFFARX1 I_9325 (I161326,I2859,I160919,I160908,);
not I_9326 (I161446,I2866);
DFFARX1 I_9327 (I492826,I2859,I161446,I161472,);
nand I_9328 (I161480,I492841,I492826);
and I_9329 (I161497,I161480,I492844);
DFFARX1 I_9330 (I161497,I2859,I161446,I161523,);
nor I_9331 (I161414,I161523,I161472);
not I_9332 (I161545,I161523);
DFFARX1 I_9333 (I492850,I2859,I161446,I161571,);
nand I_9334 (I161579,I161571,I492832);
not I_9335 (I161596,I161579);
DFFARX1 I_9336 (I161596,I2859,I161446,I161622,);
not I_9337 (I161438,I161622);
nor I_9338 (I161644,I161472,I161579);
nor I_9339 (I161420,I161523,I161644);
DFFARX1 I_9340 (I492829,I2859,I161446,I161684,);
DFFARX1 I_9341 (I161684,I2859,I161446,I161701,);
not I_9342 (I161709,I161701);
not I_9343 (I161726,I161684);
nand I_9344 (I161423,I161726,I161545);
nand I_9345 (I161757,I492829,I492835);
and I_9346 (I161774,I161757,I492847);
DFFARX1 I_9347 (I161774,I2859,I161446,I161800,);
nor I_9348 (I161808,I161800,I161472);
DFFARX1 I_9349 (I161808,I2859,I161446,I161411,);
DFFARX1 I_9350 (I161800,I2859,I161446,I161429,);
nor I_9351 (I161853,I492838,I492835);
not I_9352 (I161870,I161853);
nor I_9353 (I161432,I161709,I161870);
nand I_9354 (I161417,I161726,I161870);
nor I_9355 (I161426,I161472,I161853);
DFFARX1 I_9356 (I161853,I2859,I161446,I161435,);
not I_9357 (I161973,I2866);
DFFARX1 I_9358 (I452944,I2859,I161973,I161999,);
nand I_9359 (I162007,I452959,I452944);
and I_9360 (I162024,I162007,I452962);
DFFARX1 I_9361 (I162024,I2859,I161973,I162050,);
nor I_9362 (I161941,I162050,I161999);
not I_9363 (I162072,I162050);
DFFARX1 I_9364 (I452968,I2859,I161973,I162098,);
nand I_9365 (I162106,I162098,I452950);
not I_9366 (I162123,I162106);
DFFARX1 I_9367 (I162123,I2859,I161973,I162149,);
not I_9368 (I161965,I162149);
nor I_9369 (I162171,I161999,I162106);
nor I_9370 (I161947,I162050,I162171);
DFFARX1 I_9371 (I452947,I2859,I161973,I162211,);
DFFARX1 I_9372 (I162211,I2859,I161973,I162228,);
not I_9373 (I162236,I162228);
not I_9374 (I162253,I162211);
nand I_9375 (I161950,I162253,I162072);
nand I_9376 (I162284,I452947,I452953);
and I_9377 (I162301,I162284,I452965);
DFFARX1 I_9378 (I162301,I2859,I161973,I162327,);
nor I_9379 (I162335,I162327,I161999);
DFFARX1 I_9380 (I162335,I2859,I161973,I161938,);
DFFARX1 I_9381 (I162327,I2859,I161973,I161956,);
nor I_9382 (I162380,I452956,I452953);
not I_9383 (I162397,I162380);
nor I_9384 (I161959,I162236,I162397);
nand I_9385 (I161944,I162253,I162397);
nor I_9386 (I161953,I161999,I162380);
DFFARX1 I_9387 (I162380,I2859,I161973,I161962,);
not I_9388 (I162500,I2866);
DFFARX1 I_9389 (I198279,I2859,I162500,I162526,);
nand I_9390 (I162534,I198291,I198270);
and I_9391 (I162551,I162534,I198294);
DFFARX1 I_9392 (I162551,I2859,I162500,I162577,);
nor I_9393 (I162468,I162577,I162526);
not I_9394 (I162599,I162577);
DFFARX1 I_9395 (I198285,I2859,I162500,I162625,);
nand I_9396 (I162633,I162625,I198267);
not I_9397 (I162650,I162633);
DFFARX1 I_9398 (I162650,I2859,I162500,I162676,);
not I_9399 (I162492,I162676);
nor I_9400 (I162698,I162526,I162633);
nor I_9401 (I162474,I162577,I162698);
DFFARX1 I_9402 (I198282,I2859,I162500,I162738,);
DFFARX1 I_9403 (I162738,I2859,I162500,I162755,);
not I_9404 (I162763,I162755);
not I_9405 (I162780,I162738);
nand I_9406 (I162477,I162780,I162599);
nand I_9407 (I162811,I198267,I198273);
and I_9408 (I162828,I162811,I198276);
DFFARX1 I_9409 (I162828,I2859,I162500,I162854,);
nor I_9410 (I162862,I162854,I162526);
DFFARX1 I_9411 (I162862,I2859,I162500,I162465,);
DFFARX1 I_9412 (I162854,I2859,I162500,I162483,);
nor I_9413 (I162907,I198288,I198273);
not I_9414 (I162924,I162907);
nor I_9415 (I162486,I162763,I162924);
nand I_9416 (I162471,I162780,I162924);
nor I_9417 (I162480,I162526,I162907);
DFFARX1 I_9418 (I162907,I2859,I162500,I162489,);
not I_9419 (I163027,I2866);
DFFARX1 I_9420 (I43655,I2859,I163027,I163053,);
nand I_9421 (I163061,I43667,I43676);
and I_9422 (I163078,I163061,I43655);
DFFARX1 I_9423 (I163078,I2859,I163027,I163104,);
nor I_9424 (I162995,I163104,I163053);
not I_9425 (I163126,I163104);
DFFARX1 I_9426 (I43670,I2859,I163027,I163152,);
nand I_9427 (I163160,I163152,I43658);
not I_9428 (I163177,I163160);
DFFARX1 I_9429 (I163177,I2859,I163027,I163203,);
not I_9430 (I163019,I163203);
nor I_9431 (I163225,I163053,I163160);
nor I_9432 (I163001,I163104,I163225);
DFFARX1 I_9433 (I43661,I2859,I163027,I163265,);
DFFARX1 I_9434 (I163265,I2859,I163027,I163282,);
not I_9435 (I163290,I163282);
not I_9436 (I163307,I163265);
nand I_9437 (I163004,I163307,I163126);
nand I_9438 (I163338,I43652,I43652);
and I_9439 (I163355,I163338,I43664);
DFFARX1 I_9440 (I163355,I2859,I163027,I163381,);
nor I_9441 (I163389,I163381,I163053);
DFFARX1 I_9442 (I163389,I2859,I163027,I162992,);
DFFARX1 I_9443 (I163381,I2859,I163027,I163010,);
nor I_9444 (I163434,I43673,I43652);
not I_9445 (I163451,I163434);
nor I_9446 (I163013,I163290,I163451);
nand I_9447 (I162998,I163307,I163451);
nor I_9448 (I163007,I163053,I163434);
DFFARX1 I_9449 (I163434,I2859,I163027,I163016,);
not I_9450 (I163554,I2866);
DFFARX1 I_9451 (I313012,I2859,I163554,I163580,);
nand I_9452 (I163588,I313003,I313018);
and I_9453 (I163605,I163588,I313024);
DFFARX1 I_9454 (I163605,I2859,I163554,I163631,);
nor I_9455 (I163522,I163631,I163580);
not I_9456 (I163653,I163631);
DFFARX1 I_9457 (I313009,I2859,I163554,I163679,);
nand I_9458 (I163687,I163679,I313003);
not I_9459 (I163704,I163687);
DFFARX1 I_9460 (I163704,I2859,I163554,I163730,);
not I_9461 (I163546,I163730);
nor I_9462 (I163752,I163580,I163687);
nor I_9463 (I163528,I163631,I163752);
DFFARX1 I_9464 (I313006,I2859,I163554,I163792,);
DFFARX1 I_9465 (I163792,I2859,I163554,I163809,);
not I_9466 (I163817,I163809);
not I_9467 (I163834,I163792);
nand I_9468 (I163531,I163834,I163653);
nand I_9469 (I163865,I313000,I313015);
and I_9470 (I163882,I163865,I313000);
DFFARX1 I_9471 (I163882,I2859,I163554,I163908,);
nor I_9472 (I163916,I163908,I163580);
DFFARX1 I_9473 (I163916,I2859,I163554,I163519,);
DFFARX1 I_9474 (I163908,I2859,I163554,I163537,);
nor I_9475 (I163961,I313021,I313015);
not I_9476 (I163978,I163961);
nor I_9477 (I163540,I163817,I163978);
nand I_9478 (I163525,I163834,I163978);
nor I_9479 (I163534,I163580,I163961);
DFFARX1 I_9480 (I163961,I2859,I163554,I163543,);
not I_9481 (I164081,I2866);
DFFARX1 I_9482 (I291048,I2859,I164081,I164107,);
nand I_9483 (I164115,I291039,I291054);
and I_9484 (I164132,I164115,I291060);
DFFARX1 I_9485 (I164132,I2859,I164081,I164158,);
nor I_9486 (I164049,I164158,I164107);
not I_9487 (I164180,I164158);
DFFARX1 I_9488 (I291045,I2859,I164081,I164206,);
nand I_9489 (I164214,I164206,I291039);
not I_9490 (I164231,I164214);
DFFARX1 I_9491 (I164231,I2859,I164081,I164257,);
not I_9492 (I164073,I164257);
nor I_9493 (I164279,I164107,I164214);
nor I_9494 (I164055,I164158,I164279);
DFFARX1 I_9495 (I291042,I2859,I164081,I164319,);
DFFARX1 I_9496 (I164319,I2859,I164081,I164336,);
not I_9497 (I164344,I164336);
not I_9498 (I164361,I164319);
nand I_9499 (I164058,I164361,I164180);
nand I_9500 (I164392,I291036,I291051);
and I_9501 (I164409,I164392,I291036);
DFFARX1 I_9502 (I164409,I2859,I164081,I164435,);
nor I_9503 (I164443,I164435,I164107);
DFFARX1 I_9504 (I164443,I2859,I164081,I164046,);
DFFARX1 I_9505 (I164435,I2859,I164081,I164064,);
nor I_9506 (I164488,I291057,I291051);
not I_9507 (I164505,I164488);
nor I_9508 (I164067,I164344,I164505);
nand I_9509 (I164052,I164361,I164505);
nor I_9510 (I164061,I164107,I164488);
DFFARX1 I_9511 (I164488,I2859,I164081,I164070,);
not I_9512 (I164608,I2866);
DFFARX1 I_9513 (I384148,I2859,I164608,I164634,);
nand I_9514 (I164642,I384145,I384163);
and I_9515 (I164659,I164642,I384154);
DFFARX1 I_9516 (I164659,I2859,I164608,I164685,);
nor I_9517 (I164576,I164685,I164634);
not I_9518 (I164707,I164685);
DFFARX1 I_9519 (I384169,I2859,I164608,I164733,);
nand I_9520 (I164741,I164733,I384151);
not I_9521 (I164758,I164741);
DFFARX1 I_9522 (I164758,I2859,I164608,I164784,);
not I_9523 (I164600,I164784);
nor I_9524 (I164806,I164634,I164741);
nor I_9525 (I164582,I164685,I164806);
DFFARX1 I_9526 (I384157,I2859,I164608,I164846,);
DFFARX1 I_9527 (I164846,I2859,I164608,I164863,);
not I_9528 (I164871,I164863);
not I_9529 (I164888,I164846);
nand I_9530 (I164585,I164888,I164707);
nand I_9531 (I164919,I384145,I384172);
and I_9532 (I164936,I164919,I384160);
DFFARX1 I_9533 (I164936,I2859,I164608,I164962,);
nor I_9534 (I164970,I164962,I164634);
DFFARX1 I_9535 (I164970,I2859,I164608,I164573,);
DFFARX1 I_9536 (I164962,I2859,I164608,I164591,);
nor I_9537 (I165015,I384166,I384172);
not I_9538 (I165032,I165015);
nor I_9539 (I164594,I164871,I165032);
nand I_9540 (I164579,I164888,I165032);
nor I_9541 (I164588,I164634,I165015);
DFFARX1 I_9542 (I165015,I2859,I164608,I164597,);
not I_9543 (I165135,I2866);
DFFARX1 I_9544 (I404174,I2859,I165135,I165161,);
nand I_9545 (I165169,I404171,I404189);
and I_9546 (I165186,I165169,I404180);
DFFARX1 I_9547 (I165186,I2859,I165135,I165212,);
nor I_9548 (I165103,I165212,I165161);
not I_9549 (I165234,I165212);
DFFARX1 I_9550 (I404195,I2859,I165135,I165260,);
nand I_9551 (I165268,I165260,I404177);
not I_9552 (I165285,I165268);
DFFARX1 I_9553 (I165285,I2859,I165135,I165311,);
not I_9554 (I165127,I165311);
nor I_9555 (I165333,I165161,I165268);
nor I_9556 (I165109,I165212,I165333);
DFFARX1 I_9557 (I404183,I2859,I165135,I165373,);
DFFARX1 I_9558 (I165373,I2859,I165135,I165390,);
not I_9559 (I165398,I165390);
not I_9560 (I165415,I165373);
nand I_9561 (I165112,I165415,I165234);
nand I_9562 (I165446,I404171,I404198);
and I_9563 (I165463,I165446,I404186);
DFFARX1 I_9564 (I165463,I2859,I165135,I165489,);
nor I_9565 (I165497,I165489,I165161);
DFFARX1 I_9566 (I165497,I2859,I165135,I165100,);
DFFARX1 I_9567 (I165489,I2859,I165135,I165118,);
nor I_9568 (I165542,I404192,I404198);
not I_9569 (I165559,I165542);
nor I_9570 (I165121,I165398,I165559);
nand I_9571 (I165106,I165415,I165559);
nor I_9572 (I165115,I165161,I165542);
DFFARX1 I_9573 (I165542,I2859,I165135,I165124,);
not I_9574 (I165662,I2866);
DFFARX1 I_9575 (I260405,I2859,I165662,I165688,);
DFFARX1 I_9576 (I165688,I2859,I165662,I165705,);
not I_9577 (I165654,I165705);
not I_9578 (I165727,I165688);
nand I_9579 (I165744,I260402,I260423);
and I_9580 (I165761,I165744,I260426);
DFFARX1 I_9581 (I165761,I2859,I165662,I165787,);
not I_9582 (I165795,I165787);
DFFARX1 I_9583 (I260411,I2859,I165662,I165821,);
and I_9584 (I165829,I165821,I260414);
nand I_9585 (I165846,I165821,I260414);
nand I_9586 (I165633,I165795,I165846);
DFFARX1 I_9587 (I260417,I2859,I165662,I165886,);
nor I_9588 (I165894,I165886,I165829);
DFFARX1 I_9589 (I165894,I2859,I165662,I165627,);
nor I_9590 (I165642,I165886,I165787);
nand I_9591 (I165939,I260402,I260408);
and I_9592 (I165956,I165939,I260420);
DFFARX1 I_9593 (I165956,I2859,I165662,I165982,);
nor I_9594 (I165630,I165982,I165886);
not I_9595 (I166004,I165982);
nor I_9596 (I166021,I166004,I165795);
nor I_9597 (I166038,I165727,I166021);
DFFARX1 I_9598 (I166038,I2859,I165662,I165645,);
nor I_9599 (I166069,I166004,I165886);
nor I_9600 (I166086,I260405,I260408);
nor I_9601 (I165636,I166086,I166069);
not I_9602 (I166117,I166086);
nand I_9603 (I165639,I165846,I166117);
DFFARX1 I_9604 (I166086,I2859,I165662,I165651,);
DFFARX1 I_9605 (I166086,I2859,I165662,I165648,);
not I_9606 (I166206,I2866);
DFFARX1 I_9607 (I215491,I2859,I166206,I166232,);
DFFARX1 I_9608 (I166232,I2859,I166206,I166249,);
not I_9609 (I166198,I166249);
not I_9610 (I166271,I166232);
nand I_9611 (I166288,I215494,I215512);
and I_9612 (I166305,I166288,I215500);
DFFARX1 I_9613 (I166305,I2859,I166206,I166331,);
not I_9614 (I166339,I166331);
DFFARX1 I_9615 (I215491,I2859,I166206,I166365,);
and I_9616 (I166373,I166365,I215509);
nand I_9617 (I166390,I166365,I215509);
nand I_9618 (I166177,I166339,I166390);
DFFARX1 I_9619 (I215503,I2859,I166206,I166430,);
nor I_9620 (I166438,I166430,I166373);
DFFARX1 I_9621 (I166438,I2859,I166206,I166171,);
nor I_9622 (I166186,I166430,I166331);
nand I_9623 (I166483,I215506,I215488);
and I_9624 (I166500,I166483,I215497);
DFFARX1 I_9625 (I166500,I2859,I166206,I166526,);
nor I_9626 (I166174,I166526,I166430);
not I_9627 (I166548,I166526);
nor I_9628 (I166565,I166548,I166339);
nor I_9629 (I166582,I166271,I166565);
DFFARX1 I_9630 (I166582,I2859,I166206,I166189,);
nor I_9631 (I166613,I166548,I166430);
nor I_9632 (I166630,I215488,I215488);
nor I_9633 (I166180,I166630,I166613);
not I_9634 (I166661,I166630);
nand I_9635 (I166183,I166390,I166661);
DFFARX1 I_9636 (I166630,I2859,I166206,I166195,);
DFFARX1 I_9637 (I166630,I2859,I166206,I166192,);
not I_9638 (I166750,I2866);
DFFARX1 I_9639 (I125596,I2859,I166750,I166776,);
DFFARX1 I_9640 (I166776,I2859,I166750,I166793,);
not I_9641 (I166742,I166793);
not I_9642 (I166815,I166776);
nand I_9643 (I166832,I125575,I125599);
and I_9644 (I166849,I166832,I125602);
DFFARX1 I_9645 (I166849,I2859,I166750,I166875,);
not I_9646 (I166883,I166875);
DFFARX1 I_9647 (I125584,I2859,I166750,I166909,);
and I_9648 (I166917,I166909,I125590);
nand I_9649 (I166934,I166909,I125590);
nand I_9650 (I166721,I166883,I166934);
DFFARX1 I_9651 (I125578,I2859,I166750,I166974,);
nor I_9652 (I166982,I166974,I166917);
DFFARX1 I_9653 (I166982,I2859,I166750,I166715,);
nor I_9654 (I166730,I166974,I166875);
nand I_9655 (I167027,I125587,I125575);
and I_9656 (I167044,I167027,I125581);
DFFARX1 I_9657 (I167044,I2859,I166750,I167070,);
nor I_9658 (I166718,I167070,I166974);
not I_9659 (I167092,I167070);
nor I_9660 (I167109,I167092,I166883);
nor I_9661 (I167126,I166815,I167109);
DFFARX1 I_9662 (I167126,I2859,I166750,I166733,);
nor I_9663 (I167157,I167092,I166974);
nor I_9664 (I167174,I125593,I125575);
nor I_9665 (I166724,I167174,I167157);
not I_9666 (I167205,I167174);
nand I_9667 (I166727,I166934,I167205);
DFFARX1 I_9668 (I167174,I2859,I166750,I166739,);
DFFARX1 I_9669 (I167174,I2859,I166750,I166736,);
not I_9670 (I167294,I2866);
DFFARX1 I_9671 (I445515,I2859,I167294,I167320,);
DFFARX1 I_9672 (I167320,I2859,I167294,I167337,);
not I_9673 (I167286,I167337);
not I_9674 (I167359,I167320);
nand I_9675 (I167376,I445515,I445533);
and I_9676 (I167393,I167376,I445527);
DFFARX1 I_9677 (I167393,I2859,I167294,I167419,);
not I_9678 (I167427,I167419);
DFFARX1 I_9679 (I445521,I2859,I167294,I167453,);
and I_9680 (I167461,I167453,I445530);
nand I_9681 (I167478,I167453,I445530);
nand I_9682 (I167265,I167427,I167478);
DFFARX1 I_9683 (I445518,I2859,I167294,I167518,);
nor I_9684 (I167526,I167518,I167461);
DFFARX1 I_9685 (I167526,I2859,I167294,I167259,);
nor I_9686 (I167274,I167518,I167419);
nand I_9687 (I167571,I445518,I445536);
and I_9688 (I167588,I167571,I445521);
DFFARX1 I_9689 (I167588,I2859,I167294,I167614,);
nor I_9690 (I167262,I167614,I167518);
not I_9691 (I167636,I167614);
nor I_9692 (I167653,I167636,I167427);
nor I_9693 (I167670,I167359,I167653);
DFFARX1 I_9694 (I167670,I2859,I167294,I167277,);
nor I_9695 (I167701,I167636,I167518);
nor I_9696 (I167718,I445524,I445536);
nor I_9697 (I167268,I167718,I167701);
not I_9698 (I167749,I167718);
nand I_9699 (I167271,I167478,I167749);
DFFARX1 I_9700 (I167718,I2859,I167294,I167283,);
DFFARX1 I_9701 (I167718,I2859,I167294,I167280,);
not I_9702 (I167838,I2866);
DFFARX1 I_9703 (I484737,I2859,I167838,I167864,);
DFFARX1 I_9704 (I167864,I2859,I167838,I167881,);
not I_9705 (I167830,I167881);
not I_9706 (I167903,I167864);
nand I_9707 (I167920,I484749,I484737);
and I_9708 (I167937,I167920,I484740);
DFFARX1 I_9709 (I167937,I2859,I167838,I167963,);
not I_9710 (I167971,I167963);
DFFARX1 I_9711 (I484758,I2859,I167838,I167997,);
and I_9712 (I168005,I167997,I484734);
nand I_9713 (I168022,I167997,I484734);
nand I_9714 (I167809,I167971,I168022);
DFFARX1 I_9715 (I484752,I2859,I167838,I168062,);
nor I_9716 (I168070,I168062,I168005);
DFFARX1 I_9717 (I168070,I2859,I167838,I167803,);
nor I_9718 (I167818,I168062,I167963);
nand I_9719 (I168115,I484746,I484743);
and I_9720 (I168132,I168115,I484755);
DFFARX1 I_9721 (I168132,I2859,I167838,I168158,);
nor I_9722 (I167806,I168158,I168062);
not I_9723 (I168180,I168158);
nor I_9724 (I168197,I168180,I167971);
nor I_9725 (I168214,I167903,I168197);
DFFARX1 I_9726 (I168214,I2859,I167838,I167821,);
nor I_9727 (I168245,I168180,I168062);
nor I_9728 (I168262,I484734,I484743);
nor I_9729 (I167812,I168262,I168245);
not I_9730 (I168293,I168262);
nand I_9731 (I167815,I168022,I168293);
DFFARX1 I_9732 (I168262,I2859,I167838,I167827,);
DFFARX1 I_9733 (I168262,I2859,I167838,I167824,);
not I_9734 (I168382,I2866);
DFFARX1 I_9735 (I237285,I2859,I168382,I168408,);
DFFARX1 I_9736 (I168408,I2859,I168382,I168425,);
not I_9737 (I168374,I168425);
not I_9738 (I168447,I168408);
nand I_9739 (I168464,I237282,I237303);
and I_9740 (I168481,I168464,I237306);
DFFARX1 I_9741 (I168481,I2859,I168382,I168507,);
not I_9742 (I168515,I168507);
DFFARX1 I_9743 (I237291,I2859,I168382,I168541,);
and I_9744 (I168549,I168541,I237294);
nand I_9745 (I168566,I168541,I237294);
nand I_9746 (I168353,I168515,I168566);
DFFARX1 I_9747 (I237297,I2859,I168382,I168606,);
nor I_9748 (I168614,I168606,I168549);
DFFARX1 I_9749 (I168614,I2859,I168382,I168347,);
nor I_9750 (I168362,I168606,I168507);
nand I_9751 (I168659,I237282,I237288);
and I_9752 (I168676,I168659,I237300);
DFFARX1 I_9753 (I168676,I2859,I168382,I168702,);
nor I_9754 (I168350,I168702,I168606);
not I_9755 (I168724,I168702);
nor I_9756 (I168741,I168724,I168515);
nor I_9757 (I168758,I168447,I168741);
DFFARX1 I_9758 (I168758,I2859,I168382,I168365,);
nor I_9759 (I168789,I168724,I168606);
nor I_9760 (I168806,I237285,I237288);
nor I_9761 (I168356,I168806,I168789);
not I_9762 (I168837,I168806);
nand I_9763 (I168359,I168566,I168837);
DFFARX1 I_9764 (I168806,I2859,I168382,I168371,);
DFFARX1 I_9765 (I168806,I2859,I168382,I168368,);
not I_9766 (I168926,I2866);
DFFARX1 I_9767 (I8355,I2859,I168926,I168952,);
DFFARX1 I_9768 (I168952,I2859,I168926,I168969,);
not I_9769 (I168918,I168969);
not I_9770 (I168991,I168952);
nand I_9771 (I169008,I8343,I8358);
and I_9772 (I169025,I169008,I8346);
DFFARX1 I_9773 (I169025,I2859,I168926,I169051,);
not I_9774 (I169059,I169051);
DFFARX1 I_9775 (I8367,I2859,I168926,I169085,);
and I_9776 (I169093,I169085,I8361);
nand I_9777 (I169110,I169085,I8361);
nand I_9778 (I168897,I169059,I169110);
DFFARX1 I_9779 (I8364,I2859,I168926,I169150,);
nor I_9780 (I169158,I169150,I169093);
DFFARX1 I_9781 (I169158,I2859,I168926,I168891,);
nor I_9782 (I168906,I169150,I169051);
nand I_9783 (I169203,I8343,I8346);
and I_9784 (I169220,I169203,I8349);
DFFARX1 I_9785 (I169220,I2859,I168926,I169246,);
nor I_9786 (I168894,I169246,I169150);
not I_9787 (I169268,I169246);
nor I_9788 (I169285,I169268,I169059);
nor I_9789 (I169302,I168991,I169285);
DFFARX1 I_9790 (I169302,I2859,I168926,I168909,);
nor I_9791 (I169333,I169268,I169150);
nor I_9792 (I169350,I8352,I8346);
nor I_9793 (I168900,I169350,I169333);
not I_9794 (I169381,I169350);
nand I_9795 (I168903,I169110,I169381);
DFFARX1 I_9796 (I169350,I2859,I168926,I168915,);
DFFARX1 I_9797 (I169350,I2859,I168926,I168912,);
not I_9798 (I169470,I2866);
DFFARX1 I_9799 (I256937,I2859,I169470,I169496,);
DFFARX1 I_9800 (I169496,I2859,I169470,I169513,);
not I_9801 (I169462,I169513);
not I_9802 (I169535,I169496);
nand I_9803 (I169552,I256934,I256955);
and I_9804 (I169569,I169552,I256958);
DFFARX1 I_9805 (I169569,I2859,I169470,I169595,);
not I_9806 (I169603,I169595);
DFFARX1 I_9807 (I256943,I2859,I169470,I169629,);
and I_9808 (I169637,I169629,I256946);
nand I_9809 (I169654,I169629,I256946);
nand I_9810 (I169441,I169603,I169654);
DFFARX1 I_9811 (I256949,I2859,I169470,I169694,);
nor I_9812 (I169702,I169694,I169637);
DFFARX1 I_9813 (I169702,I2859,I169470,I169435,);
nor I_9814 (I169450,I169694,I169595);
nand I_9815 (I169747,I256934,I256940);
and I_9816 (I169764,I169747,I256952);
DFFARX1 I_9817 (I169764,I2859,I169470,I169790,);
nor I_9818 (I169438,I169790,I169694);
not I_9819 (I169812,I169790);
nor I_9820 (I169829,I169812,I169603);
nor I_9821 (I169846,I169535,I169829);
DFFARX1 I_9822 (I169846,I2859,I169470,I169453,);
nor I_9823 (I169877,I169812,I169694);
nor I_9824 (I169894,I256937,I256940);
nor I_9825 (I169444,I169894,I169877);
not I_9826 (I169925,I169894);
nand I_9827 (I169447,I169654,I169925);
DFFARX1 I_9828 (I169894,I2859,I169470,I169459,);
DFFARX1 I_9829 (I169894,I2859,I169470,I169456,);
not I_9830 (I170014,I2866);
DFFARX1 I_9831 (I306067,I2859,I170014,I170040,);
DFFARX1 I_9832 (I170040,I2859,I170014,I170057,);
not I_9833 (I170006,I170057);
not I_9834 (I170079,I170040);
nand I_9835 (I170096,I306088,I306079);
and I_9836 (I170113,I170096,I306067);
DFFARX1 I_9837 (I170113,I2859,I170014,I170139,);
not I_9838 (I170147,I170139);
DFFARX1 I_9839 (I306073,I2859,I170014,I170173,);
and I_9840 (I170181,I170173,I306070);
nand I_9841 (I170198,I170173,I306070);
nand I_9842 (I169985,I170147,I170198);
DFFARX1 I_9843 (I306064,I2859,I170014,I170238,);
nor I_9844 (I170246,I170238,I170181);
DFFARX1 I_9845 (I170246,I2859,I170014,I169979,);
nor I_9846 (I169994,I170238,I170139);
nand I_9847 (I170291,I306064,I306076);
and I_9848 (I170308,I170291,I306085);
DFFARX1 I_9849 (I170308,I2859,I170014,I170334,);
nor I_9850 (I169982,I170334,I170238);
not I_9851 (I170356,I170334);
nor I_9852 (I170373,I170356,I170147);
nor I_9853 (I170390,I170079,I170373);
DFFARX1 I_9854 (I170390,I2859,I170014,I169997,);
nor I_9855 (I170421,I170356,I170238);
nor I_9856 (I170438,I306082,I306076);
nor I_9857 (I169988,I170438,I170421);
not I_9858 (I170469,I170438);
nand I_9859 (I169991,I170198,I170469);
DFFARX1 I_9860 (I170438,I2859,I170014,I170003,);
DFFARX1 I_9861 (I170438,I2859,I170014,I170000,);
not I_9862 (I170558,I2866);
DFFARX1 I_9863 (I281213,I2859,I170558,I170584,);
DFFARX1 I_9864 (I170584,I2859,I170558,I170601,);
not I_9865 (I170550,I170601);
not I_9866 (I170623,I170584);
nand I_9867 (I170640,I281234,I281225);
and I_9868 (I170657,I170640,I281213);
DFFARX1 I_9869 (I170657,I2859,I170558,I170683,);
not I_9870 (I170691,I170683);
DFFARX1 I_9871 (I281219,I2859,I170558,I170717,);
and I_9872 (I170725,I170717,I281216);
nand I_9873 (I170742,I170717,I281216);
nand I_9874 (I170529,I170691,I170742);
DFFARX1 I_9875 (I281210,I2859,I170558,I170782,);
nor I_9876 (I170790,I170782,I170725);
DFFARX1 I_9877 (I170790,I2859,I170558,I170523,);
nor I_9878 (I170538,I170782,I170683);
nand I_9879 (I170835,I281210,I281222);
and I_9880 (I170852,I170835,I281231);
DFFARX1 I_9881 (I170852,I2859,I170558,I170878,);
nor I_9882 (I170526,I170878,I170782);
not I_9883 (I170900,I170878);
nor I_9884 (I170917,I170900,I170691);
nor I_9885 (I170934,I170623,I170917);
DFFARX1 I_9886 (I170934,I2859,I170558,I170541,);
nor I_9887 (I170965,I170900,I170782);
nor I_9888 (I170982,I281228,I281222);
nor I_9889 (I170532,I170982,I170965);
not I_9890 (I171013,I170982);
nand I_9891 (I170535,I170742,I171013);
DFFARX1 I_9892 (I170982,I2859,I170558,I170547,);
DFFARX1 I_9893 (I170982,I2859,I170558,I170544,);
not I_9894 (I171102,I2866);
DFFARX1 I_9895 (I40496,I2859,I171102,I171128,);
DFFARX1 I_9896 (I171128,I2859,I171102,I171145,);
not I_9897 (I171094,I171145);
not I_9898 (I171167,I171128);
nand I_9899 (I171184,I40511,I40490);
and I_9900 (I171201,I171184,I40493);
DFFARX1 I_9901 (I171201,I2859,I171102,I171227,);
not I_9902 (I171235,I171227);
DFFARX1 I_9903 (I40499,I2859,I171102,I171261,);
and I_9904 (I171269,I171261,I40493);
nand I_9905 (I171286,I171261,I40493);
nand I_9906 (I171073,I171235,I171286);
DFFARX1 I_9907 (I40508,I2859,I171102,I171326,);
nor I_9908 (I171334,I171326,I171269);
DFFARX1 I_9909 (I171334,I2859,I171102,I171067,);
nor I_9910 (I171082,I171326,I171227);
nand I_9911 (I171379,I40490,I40505);
and I_9912 (I171396,I171379,I40502);
DFFARX1 I_9913 (I171396,I2859,I171102,I171422,);
nor I_9914 (I171070,I171422,I171326);
not I_9915 (I171444,I171422);
nor I_9916 (I171461,I171444,I171235);
nor I_9917 (I171478,I171167,I171461);
DFFARX1 I_9918 (I171478,I2859,I171102,I171085,);
nor I_9919 (I171509,I171444,I171326);
nor I_9920 (I171526,I40514,I40505);
nor I_9921 (I171076,I171526,I171509);
not I_9922 (I171557,I171526);
nand I_9923 (I171079,I171286,I171557);
DFFARX1 I_9924 (I171526,I2859,I171102,I171091,);
DFFARX1 I_9925 (I171526,I2859,I171102,I171088,);
not I_9926 (I171646,I2866);
DFFARX1 I_9927 (I13625,I2859,I171646,I171672,);
DFFARX1 I_9928 (I171672,I2859,I171646,I171689,);
not I_9929 (I171638,I171689);
not I_9930 (I171711,I171672);
nand I_9931 (I171728,I13613,I13628);
and I_9932 (I171745,I171728,I13616);
DFFARX1 I_9933 (I171745,I2859,I171646,I171771,);
not I_9934 (I171779,I171771);
DFFARX1 I_9935 (I13637,I2859,I171646,I171805,);
and I_9936 (I171813,I171805,I13631);
nand I_9937 (I171830,I171805,I13631);
nand I_9938 (I171617,I171779,I171830);
DFFARX1 I_9939 (I13634,I2859,I171646,I171870,);
nor I_9940 (I171878,I171870,I171813);
DFFARX1 I_9941 (I171878,I2859,I171646,I171611,);
nor I_9942 (I171626,I171870,I171771);
nand I_9943 (I171923,I13613,I13616);
and I_9944 (I171940,I171923,I13619);
DFFARX1 I_9945 (I171940,I2859,I171646,I171966,);
nor I_9946 (I171614,I171966,I171870);
not I_9947 (I171988,I171966);
nor I_9948 (I172005,I171988,I171779);
nor I_9949 (I172022,I171711,I172005);
DFFARX1 I_9950 (I172022,I2859,I171646,I171629,);
nor I_9951 (I172053,I171988,I171870);
nor I_9952 (I172070,I13622,I13616);
nor I_9953 (I171620,I172070,I172053);
not I_9954 (I172101,I172070);
nand I_9955 (I171623,I171830,I172101);
DFFARX1 I_9956 (I172070,I2859,I171646,I171635,);
DFFARX1 I_9957 (I172070,I2859,I171646,I171632,);
not I_9958 (I172190,I2866);
DFFARX1 I_9959 (I509149,I2859,I172190,I172216,);
DFFARX1 I_9960 (I172216,I2859,I172190,I172233,);
not I_9961 (I172182,I172233);
not I_9962 (I172255,I172216);
nand I_9963 (I172272,I509161,I509164);
and I_9964 (I172289,I172272,I509167);
DFFARX1 I_9965 (I172289,I2859,I172190,I172315,);
not I_9966 (I172323,I172315);
DFFARX1 I_9967 (I509152,I2859,I172190,I172349,);
and I_9968 (I172357,I172349,I509158);
nand I_9969 (I172374,I172349,I509158);
nand I_9970 (I172161,I172323,I172374);
DFFARX1 I_9971 (I509146,I2859,I172190,I172414,);
nor I_9972 (I172422,I172414,I172357);
DFFARX1 I_9973 (I172422,I2859,I172190,I172155,);
nor I_9974 (I172170,I172414,I172315);
nand I_9975 (I172467,I509149,I509170);
and I_9976 (I172484,I172467,I509155);
DFFARX1 I_9977 (I172484,I2859,I172190,I172510,);
nor I_9978 (I172158,I172510,I172414);
not I_9979 (I172532,I172510);
nor I_9980 (I172549,I172532,I172323);
nor I_9981 (I172566,I172255,I172549);
DFFARX1 I_9982 (I172566,I2859,I172190,I172173,);
nor I_9983 (I172597,I172532,I172414);
nor I_9984 (I172614,I509146,I509170);
nor I_9985 (I172164,I172614,I172597);
not I_9986 (I172645,I172614);
nand I_9987 (I172167,I172374,I172645);
DFFARX1 I_9988 (I172614,I2859,I172190,I172179,);
DFFARX1 I_9989 (I172614,I2859,I172190,I172176,);
not I_9990 (I172734,I2866);
DFFARX1 I_9991 (I491095,I2859,I172734,I172760,);
DFFARX1 I_9992 (I172760,I2859,I172734,I172777,);
not I_9993 (I172726,I172777);
not I_9994 (I172799,I172760);
nand I_9995 (I172816,I491107,I491095);
and I_9996 (I172833,I172816,I491098);
DFFARX1 I_9997 (I172833,I2859,I172734,I172859,);
not I_9998 (I172867,I172859);
DFFARX1 I_9999 (I491116,I2859,I172734,I172893,);
and I_10000 (I172901,I172893,I491092);
nand I_10001 (I172918,I172893,I491092);
nand I_10002 (I172705,I172867,I172918);
DFFARX1 I_10003 (I491110,I2859,I172734,I172958,);
nor I_10004 (I172966,I172958,I172901);
DFFARX1 I_10005 (I172966,I2859,I172734,I172699,);
nor I_10006 (I172714,I172958,I172859);
nand I_10007 (I173011,I491104,I491101);
and I_10008 (I173028,I173011,I491113);
DFFARX1 I_10009 (I173028,I2859,I172734,I173054,);
nor I_10010 (I172702,I173054,I172958);
not I_10011 (I173076,I173054);
nor I_10012 (I173093,I173076,I172867);
nor I_10013 (I173110,I172799,I173093);
DFFARX1 I_10014 (I173110,I2859,I172734,I172717,);
nor I_10015 (I173141,I173076,I172958);
nor I_10016 (I173158,I491092,I491101);
nor I_10017 (I172708,I173158,I173141);
not I_10018 (I173189,I173158);
nand I_10019 (I172711,I172918,I173189);
DFFARX1 I_10020 (I173158,I2859,I172734,I172723,);
DFFARX1 I_10021 (I173158,I2859,I172734,I172720,);
not I_10022 (I173278,I2866);
DFFARX1 I_10023 (I91142,I2859,I173278,I173304,);
DFFARX1 I_10024 (I173304,I2859,I173278,I173321,);
not I_10025 (I173270,I173321);
not I_10026 (I173343,I173304);
nand I_10027 (I173360,I91154,I91133);
and I_10028 (I173377,I173360,I91136);
DFFARX1 I_10029 (I173377,I2859,I173278,I173403,);
not I_10030 (I173411,I173403);
DFFARX1 I_10031 (I91145,I2859,I173278,I173437,);
and I_10032 (I173445,I173437,I91157);
nand I_10033 (I173462,I173437,I91157);
nand I_10034 (I173249,I173411,I173462);
DFFARX1 I_10035 (I91151,I2859,I173278,I173502,);
nor I_10036 (I173510,I173502,I173445);
DFFARX1 I_10037 (I173510,I2859,I173278,I173243,);
nor I_10038 (I173258,I173502,I173403);
nand I_10039 (I173555,I91139,I91136);
and I_10040 (I173572,I173555,I91148);
DFFARX1 I_10041 (I173572,I2859,I173278,I173598,);
nor I_10042 (I173246,I173598,I173502);
not I_10043 (I173620,I173598);
nor I_10044 (I173637,I173620,I173411);
nor I_10045 (I173654,I173343,I173637);
DFFARX1 I_10046 (I173654,I2859,I173278,I173261,);
nor I_10047 (I173685,I173620,I173502);
nor I_10048 (I173702,I91133,I91136);
nor I_10049 (I173252,I173702,I173685);
not I_10050 (I173733,I173702);
nand I_10051 (I173255,I173462,I173733);
DFFARX1 I_10052 (I173702,I2859,I173278,I173267,);
DFFARX1 I_10053 (I173702,I2859,I173278,I173264,);
not I_10054 (I173822,I2866);
DFFARX1 I_10055 (I160905,I2859,I173822,I173848,);
DFFARX1 I_10056 (I173848,I2859,I173822,I173865,);
not I_10057 (I173814,I173865);
not I_10058 (I173887,I173848);
nand I_10059 (I173904,I160884,I160908);
and I_10060 (I173921,I173904,I160911);
DFFARX1 I_10061 (I173921,I2859,I173822,I173947,);
not I_10062 (I173955,I173947);
DFFARX1 I_10063 (I160893,I2859,I173822,I173981,);
and I_10064 (I173989,I173981,I160899);
nand I_10065 (I174006,I173981,I160899);
nand I_10066 (I173793,I173955,I174006);
DFFARX1 I_10067 (I160887,I2859,I173822,I174046,);
nor I_10068 (I174054,I174046,I173989);
DFFARX1 I_10069 (I174054,I2859,I173822,I173787,);
nor I_10070 (I173802,I174046,I173947);
nand I_10071 (I174099,I160896,I160884);
and I_10072 (I174116,I174099,I160890);
DFFARX1 I_10073 (I174116,I2859,I173822,I174142,);
nor I_10074 (I173790,I174142,I174046);
not I_10075 (I174164,I174142);
nor I_10076 (I174181,I174164,I173955);
nor I_10077 (I174198,I173887,I174181);
DFFARX1 I_10078 (I174198,I2859,I173822,I173805,);
nor I_10079 (I174229,I174164,I174046);
nor I_10080 (I174246,I160902,I160884);
nor I_10081 (I173796,I174246,I174229);
not I_10082 (I174277,I174246);
nand I_10083 (I173799,I174006,I174277);
DFFARX1 I_10084 (I174246,I2859,I173822,I173811,);
DFFARX1 I_10085 (I174246,I2859,I173822,I173808,);
not I_10086 (I174366,I2866);
DFFARX1 I_10087 (I408699,I2859,I174366,I174392,);
DFFARX1 I_10088 (I174392,I2859,I174366,I174409,);
not I_10089 (I174358,I174409);
not I_10090 (I174431,I174392);
nand I_10091 (I174448,I408714,I408702);
and I_10092 (I174465,I174448,I408693);
DFFARX1 I_10093 (I174465,I2859,I174366,I174491,);
not I_10094 (I174499,I174491);
DFFARX1 I_10095 (I408705,I2859,I174366,I174525,);
and I_10096 (I174533,I174525,I408696);
nand I_10097 (I174550,I174525,I408696);
nand I_10098 (I174337,I174499,I174550);
DFFARX1 I_10099 (I408711,I2859,I174366,I174590,);
nor I_10100 (I174598,I174590,I174533);
DFFARX1 I_10101 (I174598,I2859,I174366,I174331,);
nor I_10102 (I174346,I174590,I174491);
nand I_10103 (I174643,I408720,I408708);
and I_10104 (I174660,I174643,I408717);
DFFARX1 I_10105 (I174660,I2859,I174366,I174686,);
nor I_10106 (I174334,I174686,I174590);
not I_10107 (I174708,I174686);
nor I_10108 (I174725,I174708,I174499);
nor I_10109 (I174742,I174431,I174725);
DFFARX1 I_10110 (I174742,I2859,I174366,I174349,);
nor I_10111 (I174773,I174708,I174590);
nor I_10112 (I174790,I408693,I408708);
nor I_10113 (I174340,I174790,I174773);
not I_10114 (I174821,I174790);
nand I_10115 (I174343,I174550,I174821);
DFFARX1 I_10116 (I174790,I2859,I174366,I174355,);
DFFARX1 I_10117 (I174790,I2859,I174366,I174352,);
not I_10118 (I174910,I2866);
DFFARX1 I_10119 (I53671,I2859,I174910,I174936,);
DFFARX1 I_10120 (I174936,I2859,I174910,I174953,);
not I_10121 (I174902,I174953);
not I_10122 (I174975,I174936);
nand I_10123 (I174992,I53686,I53665);
and I_10124 (I175009,I174992,I53668);
DFFARX1 I_10125 (I175009,I2859,I174910,I175035,);
not I_10126 (I175043,I175035);
DFFARX1 I_10127 (I53674,I2859,I174910,I175069,);
and I_10128 (I175077,I175069,I53668);
nand I_10129 (I175094,I175069,I53668);
nand I_10130 (I174881,I175043,I175094);
DFFARX1 I_10131 (I53683,I2859,I174910,I175134,);
nor I_10132 (I175142,I175134,I175077);
DFFARX1 I_10133 (I175142,I2859,I174910,I174875,);
nor I_10134 (I174890,I175134,I175035);
nand I_10135 (I175187,I53665,I53680);
and I_10136 (I175204,I175187,I53677);
DFFARX1 I_10137 (I175204,I2859,I174910,I175230,);
nor I_10138 (I174878,I175230,I175134);
not I_10139 (I175252,I175230);
nor I_10140 (I175269,I175252,I175043);
nor I_10141 (I175286,I174975,I175269);
DFFARX1 I_10142 (I175286,I2859,I174910,I174893,);
nor I_10143 (I175317,I175252,I175134);
nor I_10144 (I175334,I53689,I53680);
nor I_10145 (I174884,I175334,I175317);
not I_10146 (I175365,I175334);
nand I_10147 (I174887,I175094,I175365);
DFFARX1 I_10148 (I175334,I2859,I174910,I174899,);
DFFARX1 I_10149 (I175334,I2859,I174910,I174896,);
not I_10150 (I175454,I2866);
DFFARX1 I_10151 (I29956,I2859,I175454,I175480,);
DFFARX1 I_10152 (I175480,I2859,I175454,I175497,);
not I_10153 (I175446,I175497);
not I_10154 (I175519,I175480);
nand I_10155 (I175536,I29971,I29950);
and I_10156 (I175553,I175536,I29953);
DFFARX1 I_10157 (I175553,I2859,I175454,I175579,);
not I_10158 (I175587,I175579);
DFFARX1 I_10159 (I29959,I2859,I175454,I175613,);
and I_10160 (I175621,I175613,I29953);
nand I_10161 (I175638,I175613,I29953);
nand I_10162 (I175425,I175587,I175638);
DFFARX1 I_10163 (I29968,I2859,I175454,I175678,);
nor I_10164 (I175686,I175678,I175621);
DFFARX1 I_10165 (I175686,I2859,I175454,I175419,);
nor I_10166 (I175434,I175678,I175579);
nand I_10167 (I175731,I29950,I29965);
and I_10168 (I175748,I175731,I29962);
DFFARX1 I_10169 (I175748,I2859,I175454,I175774,);
nor I_10170 (I175422,I175774,I175678);
not I_10171 (I175796,I175774);
nor I_10172 (I175813,I175796,I175587);
nor I_10173 (I175830,I175519,I175813);
DFFARX1 I_10174 (I175830,I2859,I175454,I175437,);
nor I_10175 (I175861,I175796,I175678);
nor I_10176 (I175878,I29974,I29965);
nor I_10177 (I175428,I175878,I175861);
not I_10178 (I175909,I175878);
nand I_10179 (I175431,I175638,I175909);
DFFARX1 I_10180 (I175878,I2859,I175454,I175443,);
DFFARX1 I_10181 (I175878,I2859,I175454,I175440,);
not I_10182 (I175998,I2866);
DFFARX1 I_10183 (I517309,I2859,I175998,I176024,);
DFFARX1 I_10184 (I176024,I2859,I175998,I176041,);
not I_10185 (I175990,I176041);
not I_10186 (I176063,I176024);
nand I_10187 (I176080,I517321,I517324);
and I_10188 (I176097,I176080,I517327);
DFFARX1 I_10189 (I176097,I2859,I175998,I176123,);
not I_10190 (I176131,I176123);
DFFARX1 I_10191 (I517312,I2859,I175998,I176157,);
and I_10192 (I176165,I176157,I517318);
nand I_10193 (I176182,I176157,I517318);
nand I_10194 (I175969,I176131,I176182);
DFFARX1 I_10195 (I517306,I2859,I175998,I176222,);
nor I_10196 (I176230,I176222,I176165);
DFFARX1 I_10197 (I176230,I2859,I175998,I175963,);
nor I_10198 (I175978,I176222,I176123);
nand I_10199 (I176275,I517309,I517330);
and I_10200 (I176292,I176275,I517315);
DFFARX1 I_10201 (I176292,I2859,I175998,I176318,);
nor I_10202 (I175966,I176318,I176222);
not I_10203 (I176340,I176318);
nor I_10204 (I176357,I176340,I176131);
nor I_10205 (I176374,I176063,I176357);
DFFARX1 I_10206 (I176374,I2859,I175998,I175981,);
nor I_10207 (I176405,I176340,I176222);
nor I_10208 (I176422,I517306,I517330);
nor I_10209 (I175972,I176422,I176405);
not I_10210 (I176453,I176422);
nand I_10211 (I175975,I176182,I176453);
DFFARX1 I_10212 (I176422,I2859,I175998,I175987,);
DFFARX1 I_10213 (I176422,I2859,I175998,I175984,);
not I_10214 (I176542,I2866);
DFFARX1 I_10215 (I450635,I2859,I176542,I176568,);
DFFARX1 I_10216 (I176568,I2859,I176542,I176585,);
not I_10217 (I176534,I176585);
not I_10218 (I176607,I176568);
nand I_10219 (I176624,I450647,I450635);
and I_10220 (I176641,I176624,I450638);
DFFARX1 I_10221 (I176641,I2859,I176542,I176667,);
not I_10222 (I176675,I176667);
DFFARX1 I_10223 (I450656,I2859,I176542,I176701,);
and I_10224 (I176709,I176701,I450632);
nand I_10225 (I176726,I176701,I450632);
nand I_10226 (I176513,I176675,I176726);
DFFARX1 I_10227 (I450650,I2859,I176542,I176766,);
nor I_10228 (I176774,I176766,I176709);
DFFARX1 I_10229 (I176774,I2859,I176542,I176507,);
nor I_10230 (I176522,I176766,I176667);
nand I_10231 (I176819,I450644,I450641);
and I_10232 (I176836,I176819,I450653);
DFFARX1 I_10233 (I176836,I2859,I176542,I176862,);
nor I_10234 (I176510,I176862,I176766);
not I_10235 (I176884,I176862);
nor I_10236 (I176901,I176884,I176675);
nor I_10237 (I176918,I176607,I176901);
DFFARX1 I_10238 (I176918,I2859,I176542,I176525,);
nor I_10239 (I176949,I176884,I176766);
nor I_10240 (I176966,I450632,I450641);
nor I_10241 (I176516,I176966,I176949);
not I_10242 (I176997,I176966);
nand I_10243 (I176519,I176726,I176997);
DFFARX1 I_10244 (I176966,I2859,I176542,I176531,);
DFFARX1 I_10245 (I176966,I2859,I176542,I176528,);
not I_10246 (I177086,I2866);
DFFARX1 I_10247 (I496297,I2859,I177086,I177112,);
DFFARX1 I_10248 (I177112,I2859,I177086,I177129,);
not I_10249 (I177078,I177129);
not I_10250 (I177151,I177112);
nand I_10251 (I177168,I496309,I496297);
and I_10252 (I177185,I177168,I496300);
DFFARX1 I_10253 (I177185,I2859,I177086,I177211,);
not I_10254 (I177219,I177211);
DFFARX1 I_10255 (I496318,I2859,I177086,I177245,);
and I_10256 (I177253,I177245,I496294);
nand I_10257 (I177270,I177245,I496294);
nand I_10258 (I177057,I177219,I177270);
DFFARX1 I_10259 (I496312,I2859,I177086,I177310,);
nor I_10260 (I177318,I177310,I177253);
DFFARX1 I_10261 (I177318,I2859,I177086,I177051,);
nor I_10262 (I177066,I177310,I177211);
nand I_10263 (I177363,I496306,I496303);
and I_10264 (I177380,I177363,I496315);
DFFARX1 I_10265 (I177380,I2859,I177086,I177406,);
nor I_10266 (I177054,I177406,I177310);
not I_10267 (I177428,I177406);
nor I_10268 (I177445,I177428,I177219);
nor I_10269 (I177462,I177151,I177445);
DFFARX1 I_10270 (I177462,I2859,I177086,I177069,);
nor I_10271 (I177493,I177428,I177310);
nor I_10272 (I177510,I496294,I496303);
nor I_10273 (I177060,I177510,I177493);
not I_10274 (I177541,I177510);
nand I_10275 (I177063,I177270,I177541);
DFFARX1 I_10276 (I177510,I2859,I177086,I177075,);
DFFARX1 I_10277 (I177510,I2859,I177086,I177072,);
not I_10278 (I177630,I2866);
DFFARX1 I_10279 (I525178,I2859,I177630,I177656,);
DFFARX1 I_10280 (I177656,I2859,I177630,I177673,);
not I_10281 (I177622,I177673);
not I_10282 (I177695,I177656);
nand I_10283 (I177712,I525175,I525172);
and I_10284 (I177729,I177712,I525160);
DFFARX1 I_10285 (I177729,I2859,I177630,I177755,);
not I_10286 (I177763,I177755);
DFFARX1 I_10287 (I525184,I2859,I177630,I177789,);
and I_10288 (I177797,I177789,I525169);
nand I_10289 (I177814,I177789,I525169);
nand I_10290 (I177601,I177763,I177814);
DFFARX1 I_10291 (I525163,I2859,I177630,I177854,);
nor I_10292 (I177862,I177854,I177797);
DFFARX1 I_10293 (I177862,I2859,I177630,I177595,);
nor I_10294 (I177610,I177854,I177755);
nand I_10295 (I177907,I525160,I525166);
and I_10296 (I177924,I177907,I525181);
DFFARX1 I_10297 (I177924,I2859,I177630,I177950,);
nor I_10298 (I177598,I177950,I177854);
not I_10299 (I177972,I177950);
nor I_10300 (I177989,I177972,I177763);
nor I_10301 (I178006,I177695,I177989);
DFFARX1 I_10302 (I178006,I2859,I177630,I177613,);
nor I_10303 (I178037,I177972,I177854);
nor I_10304 (I178054,I525163,I525166);
nor I_10305 (I177604,I178054,I178037);
not I_10306 (I178085,I178054);
nand I_10307 (I177607,I177814,I178085);
DFFARX1 I_10308 (I178054,I2859,I177630,I177619,);
DFFARX1 I_10309 (I178054,I2859,I177630,I177616,);
not I_10310 (I178174,I2866);
DFFARX1 I_10311 (I56306,I2859,I178174,I178200,);
DFFARX1 I_10312 (I178200,I2859,I178174,I178217,);
not I_10313 (I178166,I178217);
not I_10314 (I178239,I178200);
nand I_10315 (I178256,I56321,I56300);
and I_10316 (I178273,I178256,I56303);
DFFARX1 I_10317 (I178273,I2859,I178174,I178299,);
not I_10318 (I178307,I178299);
DFFARX1 I_10319 (I56309,I2859,I178174,I178333,);
and I_10320 (I178341,I178333,I56303);
nand I_10321 (I178358,I178333,I56303);
nand I_10322 (I178145,I178307,I178358);
DFFARX1 I_10323 (I56318,I2859,I178174,I178398,);
nor I_10324 (I178406,I178398,I178341);
DFFARX1 I_10325 (I178406,I2859,I178174,I178139,);
nor I_10326 (I178154,I178398,I178299);
nand I_10327 (I178451,I56300,I56315);
and I_10328 (I178468,I178451,I56312);
DFFARX1 I_10329 (I178468,I2859,I178174,I178494,);
nor I_10330 (I178142,I178494,I178398);
not I_10331 (I178516,I178494);
nor I_10332 (I178533,I178516,I178307);
nor I_10333 (I178550,I178239,I178533);
DFFARX1 I_10334 (I178550,I2859,I178174,I178157,);
nor I_10335 (I178581,I178516,I178398);
nor I_10336 (I178598,I56324,I56315);
nor I_10337 (I178148,I178598,I178581);
not I_10338 (I178629,I178598);
nand I_10339 (I178151,I178358,I178629);
DFFARX1 I_10340 (I178598,I2859,I178174,I178163,);
DFFARX1 I_10341 (I178598,I2859,I178174,I178160,);
not I_10342 (I178718,I2866);
DFFARX1 I_10343 (I322251,I2859,I178718,I178744,);
DFFARX1 I_10344 (I178744,I2859,I178718,I178761,);
not I_10345 (I178710,I178761);
not I_10346 (I178783,I178744);
nand I_10347 (I178800,I322272,I322263);
and I_10348 (I178817,I178800,I322251);
DFFARX1 I_10349 (I178817,I2859,I178718,I178843,);
not I_10350 (I178851,I178843);
DFFARX1 I_10351 (I322257,I2859,I178718,I178877,);
and I_10352 (I178885,I178877,I322254);
nand I_10353 (I178902,I178877,I322254);
nand I_10354 (I178689,I178851,I178902);
DFFARX1 I_10355 (I322248,I2859,I178718,I178942,);
nor I_10356 (I178950,I178942,I178885);
DFFARX1 I_10357 (I178950,I2859,I178718,I178683,);
nor I_10358 (I178698,I178942,I178843);
nand I_10359 (I178995,I322248,I322260);
and I_10360 (I179012,I178995,I322269);
DFFARX1 I_10361 (I179012,I2859,I178718,I179038,);
nor I_10362 (I178686,I179038,I178942);
not I_10363 (I179060,I179038);
nor I_10364 (I179077,I179060,I178851);
nor I_10365 (I179094,I178783,I179077);
DFFARX1 I_10366 (I179094,I2859,I178718,I178701,);
nor I_10367 (I179125,I179060,I178942);
nor I_10368 (I179142,I322266,I322260);
nor I_10369 (I178692,I179142,I179125);
not I_10370 (I179173,I179142);
nand I_10371 (I178695,I178902,I179173);
DFFARX1 I_10372 (I179142,I2859,I178718,I178707,);
DFFARX1 I_10373 (I179142,I2859,I178718,I178704,);
not I_10374 (I179262,I2866);
DFFARX1 I_10375 (I10990,I2859,I179262,I179288,);
DFFARX1 I_10376 (I179288,I2859,I179262,I179305,);
not I_10377 (I179254,I179305);
not I_10378 (I179327,I179288);
nand I_10379 (I179344,I10978,I10993);
and I_10380 (I179361,I179344,I10981);
DFFARX1 I_10381 (I179361,I2859,I179262,I179387,);
not I_10382 (I179395,I179387);
DFFARX1 I_10383 (I11002,I2859,I179262,I179421,);
and I_10384 (I179429,I179421,I10996);
nand I_10385 (I179446,I179421,I10996);
nand I_10386 (I179233,I179395,I179446);
DFFARX1 I_10387 (I10999,I2859,I179262,I179486,);
nor I_10388 (I179494,I179486,I179429);
DFFARX1 I_10389 (I179494,I2859,I179262,I179227,);
nor I_10390 (I179242,I179486,I179387);
nand I_10391 (I179539,I10978,I10981);
and I_10392 (I179556,I179539,I10984);
DFFARX1 I_10393 (I179556,I2859,I179262,I179582,);
nor I_10394 (I179230,I179582,I179486);
not I_10395 (I179604,I179582);
nor I_10396 (I179621,I179604,I179395);
nor I_10397 (I179638,I179327,I179621);
DFFARX1 I_10398 (I179638,I2859,I179262,I179245,);
nor I_10399 (I179669,I179604,I179486);
nor I_10400 (I179686,I10987,I10981);
nor I_10401 (I179236,I179686,I179669);
not I_10402 (I179717,I179686);
nand I_10403 (I179239,I179446,I179717);
DFFARX1 I_10404 (I179686,I2859,I179262,I179251,);
DFFARX1 I_10405 (I179686,I2859,I179262,I179248,);
not I_10406 (I179806,I2866);
DFFARX1 I_10407 (I289883,I2859,I179806,I179832,);
DFFARX1 I_10408 (I179832,I2859,I179806,I179849,);
not I_10409 (I179798,I179849);
not I_10410 (I179871,I179832);
nand I_10411 (I179888,I289904,I289895);
and I_10412 (I179905,I179888,I289883);
DFFARX1 I_10413 (I179905,I2859,I179806,I179931,);
not I_10414 (I179939,I179931);
DFFARX1 I_10415 (I289889,I2859,I179806,I179965,);
and I_10416 (I179973,I179965,I289886);
nand I_10417 (I179990,I179965,I289886);
nand I_10418 (I179777,I179939,I179990);
DFFARX1 I_10419 (I289880,I2859,I179806,I180030,);
nor I_10420 (I180038,I180030,I179973);
DFFARX1 I_10421 (I180038,I2859,I179806,I179771,);
nor I_10422 (I179786,I180030,I179931);
nand I_10423 (I180083,I289880,I289892);
and I_10424 (I180100,I180083,I289901);
DFFARX1 I_10425 (I180100,I2859,I179806,I180126,);
nor I_10426 (I179774,I180126,I180030);
not I_10427 (I180148,I180126);
nor I_10428 (I180165,I180148,I179939);
nor I_10429 (I180182,I179871,I180165);
DFFARX1 I_10430 (I180182,I2859,I179806,I179789,);
nor I_10431 (I180213,I180148,I180030);
nor I_10432 (I180230,I289898,I289892);
nor I_10433 (I179780,I180230,I180213);
not I_10434 (I180261,I180230);
nand I_10435 (I179783,I179990,I180261);
DFFARX1 I_10436 (I180230,I2859,I179806,I179795,);
DFFARX1 I_10437 (I180230,I2859,I179806,I179792,);
not I_10438 (I180350,I2866);
DFFARX1 I_10439 (I411283,I2859,I180350,I180376,);
DFFARX1 I_10440 (I180376,I2859,I180350,I180393,);
not I_10441 (I180342,I180393);
not I_10442 (I180415,I180376);
nand I_10443 (I180432,I411298,I411286);
and I_10444 (I180449,I180432,I411277);
DFFARX1 I_10445 (I180449,I2859,I180350,I180475,);
not I_10446 (I180483,I180475);
DFFARX1 I_10447 (I411289,I2859,I180350,I180509,);
and I_10448 (I180517,I180509,I411280);
nand I_10449 (I180534,I180509,I411280);
nand I_10450 (I180321,I180483,I180534);
DFFARX1 I_10451 (I411295,I2859,I180350,I180574,);
nor I_10452 (I180582,I180574,I180517);
DFFARX1 I_10453 (I180582,I2859,I180350,I180315,);
nor I_10454 (I180330,I180574,I180475);
nand I_10455 (I180627,I411304,I411292);
and I_10456 (I180644,I180627,I411301);
DFFARX1 I_10457 (I180644,I2859,I180350,I180670,);
nor I_10458 (I180318,I180670,I180574);
not I_10459 (I180692,I180670);
nor I_10460 (I180709,I180692,I180483);
nor I_10461 (I180726,I180415,I180709);
DFFARX1 I_10462 (I180726,I2859,I180350,I180333,);
nor I_10463 (I180757,I180692,I180574);
nor I_10464 (I180774,I411277,I411292);
nor I_10465 (I180324,I180774,I180757);
not I_10466 (I180805,I180774);
nand I_10467 (I180327,I180534,I180805);
DFFARX1 I_10468 (I180774,I2859,I180350,I180339,);
DFFARX1 I_10469 (I180774,I2859,I180350,I180336,);
not I_10470 (I180894,I2866);
DFFARX1 I_10471 (I391903,I2859,I180894,I180920,);
DFFARX1 I_10472 (I180920,I2859,I180894,I180937,);
not I_10473 (I180886,I180937);
not I_10474 (I180959,I180920);
nand I_10475 (I180976,I391918,I391906);
and I_10476 (I180993,I180976,I391897);
DFFARX1 I_10477 (I180993,I2859,I180894,I181019,);
not I_10478 (I181027,I181019);
DFFARX1 I_10479 (I391909,I2859,I180894,I181053,);
and I_10480 (I181061,I181053,I391900);
nand I_10481 (I181078,I181053,I391900);
nand I_10482 (I180865,I181027,I181078);
DFFARX1 I_10483 (I391915,I2859,I180894,I181118,);
nor I_10484 (I181126,I181118,I181061);
DFFARX1 I_10485 (I181126,I2859,I180894,I180859,);
nor I_10486 (I180874,I181118,I181019);
nand I_10487 (I181171,I391924,I391912);
and I_10488 (I181188,I181171,I391921);
DFFARX1 I_10489 (I181188,I2859,I180894,I181214,);
nor I_10490 (I180862,I181214,I181118);
not I_10491 (I181236,I181214);
nor I_10492 (I181253,I181236,I181027);
nor I_10493 (I181270,I180959,I181253);
DFFARX1 I_10494 (I181270,I2859,I180894,I180877,);
nor I_10495 (I181301,I181236,I181118);
nor I_10496 (I181318,I391897,I391912);
nor I_10497 (I180868,I181318,I181301);
not I_10498 (I181349,I181318);
nand I_10499 (I180871,I181078,I181349);
DFFARX1 I_10500 (I181318,I2859,I180894,I180883,);
DFFARX1 I_10501 (I181318,I2859,I180894,I180880,);
not I_10502 (I181438,I2866);
DFFARX1 I_10503 (I450057,I2859,I181438,I181464,);
DFFARX1 I_10504 (I181464,I2859,I181438,I181481,);
not I_10505 (I181430,I181481);
not I_10506 (I181503,I181464);
nand I_10507 (I181520,I450069,I450057);
and I_10508 (I181537,I181520,I450060);
DFFARX1 I_10509 (I181537,I2859,I181438,I181563,);
not I_10510 (I181571,I181563);
DFFARX1 I_10511 (I450078,I2859,I181438,I181597,);
and I_10512 (I181605,I181597,I450054);
nand I_10513 (I181622,I181597,I450054);
nand I_10514 (I181409,I181571,I181622);
DFFARX1 I_10515 (I450072,I2859,I181438,I181662,);
nor I_10516 (I181670,I181662,I181605);
DFFARX1 I_10517 (I181670,I2859,I181438,I181403,);
nor I_10518 (I181418,I181662,I181563);
nand I_10519 (I181715,I450066,I450063);
and I_10520 (I181732,I181715,I450075);
DFFARX1 I_10521 (I181732,I2859,I181438,I181758,);
nor I_10522 (I181406,I181758,I181662);
not I_10523 (I181780,I181758);
nor I_10524 (I181797,I181780,I181571);
nor I_10525 (I181814,I181503,I181797);
DFFARX1 I_10526 (I181814,I2859,I181438,I181421,);
nor I_10527 (I181845,I181780,I181662);
nor I_10528 (I181862,I450054,I450063);
nor I_10529 (I181412,I181862,I181845);
not I_10530 (I181893,I181862);
nand I_10531 (I181415,I181622,I181893);
DFFARX1 I_10532 (I181862,I2859,I181438,I181427,);
DFFARX1 I_10533 (I181862,I2859,I181438,I181424,);
not I_10534 (I181982,I2866);
DFFARX1 I_10535 (I489939,I2859,I181982,I182008,);
DFFARX1 I_10536 (I182008,I2859,I181982,I182025,);
not I_10537 (I181974,I182025);
not I_10538 (I182047,I182008);
nand I_10539 (I182064,I489951,I489939);
and I_10540 (I182081,I182064,I489942);
DFFARX1 I_10541 (I182081,I2859,I181982,I182107,);
not I_10542 (I182115,I182107);
DFFARX1 I_10543 (I489960,I2859,I181982,I182141,);
and I_10544 (I182149,I182141,I489936);
nand I_10545 (I182166,I182141,I489936);
nand I_10546 (I181953,I182115,I182166);
DFFARX1 I_10547 (I489954,I2859,I181982,I182206,);
nor I_10548 (I182214,I182206,I182149);
DFFARX1 I_10549 (I182214,I2859,I181982,I181947,);
nor I_10550 (I181962,I182206,I182107);
nand I_10551 (I182259,I489948,I489945);
and I_10552 (I182276,I182259,I489957);
DFFARX1 I_10553 (I182276,I2859,I181982,I182302,);
nor I_10554 (I181950,I182302,I182206);
not I_10555 (I182324,I182302);
nor I_10556 (I182341,I182324,I182115);
nor I_10557 (I182358,I182047,I182341);
DFFARX1 I_10558 (I182358,I2859,I181982,I181965,);
nor I_10559 (I182389,I182324,I182206);
nor I_10560 (I182406,I489936,I489945);
nor I_10561 (I181956,I182406,I182389);
not I_10562 (I182437,I182406);
nand I_10563 (I181959,I182166,I182437);
DFFARX1 I_10564 (I182406,I2859,I181982,I181971,);
DFFARX1 I_10565 (I182406,I2859,I181982,I181968,);
not I_10566 (I182526,I2866);
DFFARX1 I_10567 (I35226,I2859,I182526,I182552,);
DFFARX1 I_10568 (I182552,I2859,I182526,I182569,);
not I_10569 (I182518,I182569);
not I_10570 (I182591,I182552);
nand I_10571 (I182608,I35241,I35220);
and I_10572 (I182625,I182608,I35223);
DFFARX1 I_10573 (I182625,I2859,I182526,I182651,);
not I_10574 (I182659,I182651);
DFFARX1 I_10575 (I35229,I2859,I182526,I182685,);
and I_10576 (I182693,I182685,I35223);
nand I_10577 (I182710,I182685,I35223);
nand I_10578 (I182497,I182659,I182710);
DFFARX1 I_10579 (I35238,I2859,I182526,I182750,);
nor I_10580 (I182758,I182750,I182693);
DFFARX1 I_10581 (I182758,I2859,I182526,I182491,);
nor I_10582 (I182506,I182750,I182651);
nand I_10583 (I182803,I35220,I35235);
and I_10584 (I182820,I182803,I35232);
DFFARX1 I_10585 (I182820,I2859,I182526,I182846,);
nor I_10586 (I182494,I182846,I182750);
not I_10587 (I182868,I182846);
nor I_10588 (I182885,I182868,I182659);
nor I_10589 (I182902,I182591,I182885);
DFFARX1 I_10590 (I182902,I2859,I182526,I182509,);
nor I_10591 (I182933,I182868,I182750);
nor I_10592 (I182950,I35244,I35235);
nor I_10593 (I182500,I182950,I182933);
not I_10594 (I182981,I182950);
nand I_10595 (I182503,I182710,I182981);
DFFARX1 I_10596 (I182950,I2859,I182526,I182515,);
DFFARX1 I_10597 (I182950,I2859,I182526,I182512,);
not I_10598 (I183070,I2866);
DFFARX1 I_10599 (I301443,I2859,I183070,I183096,);
DFFARX1 I_10600 (I183096,I2859,I183070,I183113,);
not I_10601 (I183062,I183113);
not I_10602 (I183135,I183096);
nand I_10603 (I183152,I301464,I301455);
and I_10604 (I183169,I183152,I301443);
DFFARX1 I_10605 (I183169,I2859,I183070,I183195,);
not I_10606 (I183203,I183195);
DFFARX1 I_10607 (I301449,I2859,I183070,I183229,);
and I_10608 (I183237,I183229,I301446);
nand I_10609 (I183254,I183229,I301446);
nand I_10610 (I183041,I183203,I183254);
DFFARX1 I_10611 (I301440,I2859,I183070,I183294,);
nor I_10612 (I183302,I183294,I183237);
DFFARX1 I_10613 (I183302,I2859,I183070,I183035,);
nor I_10614 (I183050,I183294,I183195);
nand I_10615 (I183347,I301440,I301452);
and I_10616 (I183364,I183347,I301461);
DFFARX1 I_10617 (I183364,I2859,I183070,I183390,);
nor I_10618 (I183038,I183390,I183294);
not I_10619 (I183412,I183390);
nor I_10620 (I183429,I183412,I183203);
nor I_10621 (I183446,I183135,I183429);
DFFARX1 I_10622 (I183446,I2859,I183070,I183053,);
nor I_10623 (I183477,I183412,I183294);
nor I_10624 (I183494,I301458,I301452);
nor I_10625 (I183044,I183494,I183477);
not I_10626 (I183525,I183494);
nand I_10627 (I183047,I183254,I183525);
DFFARX1 I_10628 (I183494,I2859,I183070,I183059,);
DFFARX1 I_10629 (I183494,I2859,I183070,I183056,);
not I_10630 (I183614,I2866);
DFFARX1 I_10631 (I226201,I2859,I183614,I183640,);
DFFARX1 I_10632 (I183640,I2859,I183614,I183657,);
not I_10633 (I183606,I183657);
not I_10634 (I183679,I183640);
nand I_10635 (I183696,I226204,I226222);
and I_10636 (I183713,I183696,I226210);
DFFARX1 I_10637 (I183713,I2859,I183614,I183739,);
not I_10638 (I183747,I183739);
DFFARX1 I_10639 (I226201,I2859,I183614,I183773,);
and I_10640 (I183781,I183773,I226219);
nand I_10641 (I183798,I183773,I226219);
nand I_10642 (I183585,I183747,I183798);
DFFARX1 I_10643 (I226213,I2859,I183614,I183838,);
nor I_10644 (I183846,I183838,I183781);
DFFARX1 I_10645 (I183846,I2859,I183614,I183579,);
nor I_10646 (I183594,I183838,I183739);
nand I_10647 (I183891,I226216,I226198);
and I_10648 (I183908,I183891,I226207);
DFFARX1 I_10649 (I183908,I2859,I183614,I183934,);
nor I_10650 (I183582,I183934,I183838);
not I_10651 (I183956,I183934);
nor I_10652 (I183973,I183956,I183747);
nor I_10653 (I183990,I183679,I183973);
DFFARX1 I_10654 (I183990,I2859,I183614,I183597,);
nor I_10655 (I184021,I183956,I183838);
nor I_10656 (I184038,I226198,I226198);
nor I_10657 (I183588,I184038,I184021);
not I_10658 (I184069,I184038);
nand I_10659 (I183591,I183798,I184069);
DFFARX1 I_10660 (I184038,I2859,I183614,I183603,);
DFFARX1 I_10661 (I184038,I2859,I183614,I183600,);
not I_10662 (I184158,I2866);
DFFARX1 I_10663 (I214301,I2859,I184158,I184184,);
DFFARX1 I_10664 (I184184,I2859,I184158,I184201,);
not I_10665 (I184150,I184201);
not I_10666 (I184223,I184184);
nand I_10667 (I184240,I214304,I214322);
and I_10668 (I184257,I184240,I214310);
DFFARX1 I_10669 (I184257,I2859,I184158,I184283,);
not I_10670 (I184291,I184283);
DFFARX1 I_10671 (I214301,I2859,I184158,I184317,);
and I_10672 (I184325,I184317,I214319);
nand I_10673 (I184342,I184317,I214319);
nand I_10674 (I184129,I184291,I184342);
DFFARX1 I_10675 (I214313,I2859,I184158,I184382,);
nor I_10676 (I184390,I184382,I184325);
DFFARX1 I_10677 (I184390,I2859,I184158,I184123,);
nor I_10678 (I184138,I184382,I184283);
nand I_10679 (I184435,I214316,I214298);
and I_10680 (I184452,I184435,I214307);
DFFARX1 I_10681 (I184452,I2859,I184158,I184478,);
nor I_10682 (I184126,I184478,I184382);
not I_10683 (I184500,I184478);
nor I_10684 (I184517,I184500,I184291);
nor I_10685 (I184534,I184223,I184517);
DFFARX1 I_10686 (I184534,I2859,I184158,I184141,);
nor I_10687 (I184565,I184500,I184382);
nor I_10688 (I184582,I214298,I214298);
nor I_10689 (I184132,I184582,I184565);
not I_10690 (I184613,I184582);
nand I_10691 (I184135,I184342,I184613);
DFFARX1 I_10692 (I184582,I2859,I184158,I184147,);
DFFARX1 I_10693 (I184582,I2859,I184158,I184144,);
not I_10694 (I184702,I2866);
DFFARX1 I_10695 (I81622,I2859,I184702,I184728,);
DFFARX1 I_10696 (I184728,I2859,I184702,I184745,);
not I_10697 (I184694,I184745);
not I_10698 (I184767,I184728);
nand I_10699 (I184784,I81634,I81613);
and I_10700 (I184801,I184784,I81616);
DFFARX1 I_10701 (I184801,I2859,I184702,I184827,);
not I_10702 (I184835,I184827);
DFFARX1 I_10703 (I81625,I2859,I184702,I184861,);
and I_10704 (I184869,I184861,I81637);
nand I_10705 (I184886,I184861,I81637);
nand I_10706 (I184673,I184835,I184886);
DFFARX1 I_10707 (I81631,I2859,I184702,I184926,);
nor I_10708 (I184934,I184926,I184869);
DFFARX1 I_10709 (I184934,I2859,I184702,I184667,);
nor I_10710 (I184682,I184926,I184827);
nand I_10711 (I184979,I81619,I81616);
and I_10712 (I184996,I184979,I81628);
DFFARX1 I_10713 (I184996,I2859,I184702,I185022,);
nor I_10714 (I184670,I185022,I184926);
not I_10715 (I185044,I185022);
nor I_10716 (I185061,I185044,I184835);
nor I_10717 (I185078,I184767,I185061);
DFFARX1 I_10718 (I185078,I2859,I184702,I184685,);
nor I_10719 (I185109,I185044,I184926);
nor I_10720 (I185126,I81613,I81616);
nor I_10721 (I184676,I185126,I185109);
not I_10722 (I185157,I185126);
nand I_10723 (I184679,I184886,I185157);
DFFARX1 I_10724 (I185126,I2859,I184702,I184691,);
DFFARX1 I_10725 (I185126,I2859,I184702,I184688,);
not I_10726 (I185246,I2866);
DFFARX1 I_10727 (I142460,I2859,I185246,I185272,);
DFFARX1 I_10728 (I185272,I2859,I185246,I185289,);
not I_10729 (I185238,I185289);
not I_10730 (I185311,I185272);
nand I_10731 (I185328,I142439,I142463);
and I_10732 (I185345,I185328,I142466);
DFFARX1 I_10733 (I185345,I2859,I185246,I185371,);
not I_10734 (I185379,I185371);
DFFARX1 I_10735 (I142448,I2859,I185246,I185405,);
and I_10736 (I185413,I185405,I142454);
nand I_10737 (I185430,I185405,I142454);
nand I_10738 (I185217,I185379,I185430);
DFFARX1 I_10739 (I142442,I2859,I185246,I185470,);
nor I_10740 (I185478,I185470,I185413);
DFFARX1 I_10741 (I185478,I2859,I185246,I185211,);
nor I_10742 (I185226,I185470,I185371);
nand I_10743 (I185523,I142451,I142439);
and I_10744 (I185540,I185523,I142445);
DFFARX1 I_10745 (I185540,I2859,I185246,I185566,);
nor I_10746 (I185214,I185566,I185470);
not I_10747 (I185588,I185566);
nor I_10748 (I185605,I185588,I185379);
nor I_10749 (I185622,I185311,I185605);
DFFARX1 I_10750 (I185622,I2859,I185246,I185229,);
nor I_10751 (I185653,I185588,I185470);
nor I_10752 (I185670,I142457,I142439);
nor I_10753 (I185220,I185670,I185653);
not I_10754 (I185701,I185670);
nand I_10755 (I185223,I185430,I185701);
DFFARX1 I_10756 (I185670,I2859,I185246,I185235,);
DFFARX1 I_10757 (I185670,I2859,I185246,I185232,);
not I_10758 (I185790,I2866);
DFFARX1 I_10759 (I395133,I2859,I185790,I185816,);
DFFARX1 I_10760 (I185816,I2859,I185790,I185833,);
not I_10761 (I185782,I185833);
not I_10762 (I185855,I185816);
nand I_10763 (I185872,I395148,I395136);
and I_10764 (I185889,I185872,I395127);
DFFARX1 I_10765 (I185889,I2859,I185790,I185915,);
not I_10766 (I185923,I185915);
DFFARX1 I_10767 (I395139,I2859,I185790,I185949,);
and I_10768 (I185957,I185949,I395130);
nand I_10769 (I185974,I185949,I395130);
nand I_10770 (I185761,I185923,I185974);
DFFARX1 I_10771 (I395145,I2859,I185790,I186014,);
nor I_10772 (I186022,I186014,I185957);
DFFARX1 I_10773 (I186022,I2859,I185790,I185755,);
nor I_10774 (I185770,I186014,I185915);
nand I_10775 (I186067,I395154,I395142);
and I_10776 (I186084,I186067,I395151);
DFFARX1 I_10777 (I186084,I2859,I185790,I186110,);
nor I_10778 (I185758,I186110,I186014);
not I_10779 (I186132,I186110);
nor I_10780 (I186149,I186132,I185923);
nor I_10781 (I186166,I185855,I186149);
DFFARX1 I_10782 (I186166,I2859,I185790,I185773,);
nor I_10783 (I186197,I186132,I186014);
nor I_10784 (I186214,I395127,I395142);
nor I_10785 (I185764,I186214,I186197);
not I_10786 (I186245,I186214);
nand I_10787 (I185767,I185974,I186245);
DFFARX1 I_10788 (I186214,I2859,I185790,I185779,);
DFFARX1 I_10789 (I186214,I2859,I185790,I185776,);
not I_10790 (I186334,I2866);
DFFARX1 I_10791 (I378983,I2859,I186334,I186360,);
DFFARX1 I_10792 (I186360,I2859,I186334,I186377,);
not I_10793 (I186326,I186377);
not I_10794 (I186399,I186360);
nand I_10795 (I186416,I378998,I378986);
and I_10796 (I186433,I186416,I378977);
DFFARX1 I_10797 (I186433,I2859,I186334,I186459,);
not I_10798 (I186467,I186459);
DFFARX1 I_10799 (I378989,I2859,I186334,I186493,);
and I_10800 (I186501,I186493,I378980);
nand I_10801 (I186518,I186493,I378980);
nand I_10802 (I186305,I186467,I186518);
DFFARX1 I_10803 (I378995,I2859,I186334,I186558,);
nor I_10804 (I186566,I186558,I186501);
DFFARX1 I_10805 (I186566,I2859,I186334,I186299,);
nor I_10806 (I186314,I186558,I186459);
nand I_10807 (I186611,I379004,I378992);
and I_10808 (I186628,I186611,I379001);
DFFARX1 I_10809 (I186628,I2859,I186334,I186654,);
nor I_10810 (I186302,I186654,I186558);
not I_10811 (I186676,I186654);
nor I_10812 (I186693,I186676,I186467);
nor I_10813 (I186710,I186399,I186693);
DFFARX1 I_10814 (I186710,I2859,I186334,I186317,);
nor I_10815 (I186741,I186676,I186558);
nor I_10816 (I186758,I378977,I378992);
nor I_10817 (I186308,I186758,I186741);
not I_10818 (I186789,I186758);
nand I_10819 (I186311,I186518,I186789);
DFFARX1 I_10820 (I186758,I2859,I186334,I186323,);
DFFARX1 I_10821 (I186758,I2859,I186334,I186320,);
not I_10822 (I186878,I2866);
DFFARX1 I_10823 (I82812,I2859,I186878,I186904,);
DFFARX1 I_10824 (I186904,I2859,I186878,I186921,);
not I_10825 (I186870,I186921);
not I_10826 (I186943,I186904);
nand I_10827 (I186960,I82824,I82803);
and I_10828 (I186977,I186960,I82806);
DFFARX1 I_10829 (I186977,I2859,I186878,I187003,);
not I_10830 (I187011,I187003);
DFFARX1 I_10831 (I82815,I2859,I186878,I187037,);
and I_10832 (I187045,I187037,I82827);
nand I_10833 (I187062,I187037,I82827);
nand I_10834 (I186849,I187011,I187062);
DFFARX1 I_10835 (I82821,I2859,I186878,I187102,);
nor I_10836 (I187110,I187102,I187045);
DFFARX1 I_10837 (I187110,I2859,I186878,I186843,);
nor I_10838 (I186858,I187102,I187003);
nand I_10839 (I187155,I82809,I82806);
and I_10840 (I187172,I187155,I82818);
DFFARX1 I_10841 (I187172,I2859,I186878,I187198,);
nor I_10842 (I186846,I187198,I187102);
not I_10843 (I187220,I187198);
nor I_10844 (I187237,I187220,I187011);
nor I_10845 (I187254,I186943,I187237);
DFFARX1 I_10846 (I187254,I2859,I186878,I186861,);
nor I_10847 (I187285,I187220,I187102);
nor I_10848 (I187302,I82803,I82806);
nor I_10849 (I186852,I187302,I187285);
not I_10850 (I187333,I187302);
nand I_10851 (I186855,I187062,I187333);
DFFARX1 I_10852 (I187302,I2859,I186878,I186867,);
DFFARX1 I_10853 (I187302,I2859,I186878,I186864,);
not I_10854 (I187422,I2866);
DFFARX1 I_10855 (I57360,I2859,I187422,I187448,);
DFFARX1 I_10856 (I187448,I2859,I187422,I187465,);
not I_10857 (I187414,I187465);
not I_10858 (I187487,I187448);
nand I_10859 (I187504,I57375,I57354);
and I_10860 (I187521,I187504,I57357);
DFFARX1 I_10861 (I187521,I2859,I187422,I187547,);
not I_10862 (I187555,I187547);
DFFARX1 I_10863 (I57363,I2859,I187422,I187581,);
and I_10864 (I187589,I187581,I57357);
nand I_10865 (I187606,I187581,I57357);
nand I_10866 (I187393,I187555,I187606);
DFFARX1 I_10867 (I57372,I2859,I187422,I187646,);
nor I_10868 (I187654,I187646,I187589);
DFFARX1 I_10869 (I187654,I2859,I187422,I187387,);
nor I_10870 (I187402,I187646,I187547);
nand I_10871 (I187699,I57354,I57369);
and I_10872 (I187716,I187699,I57366);
DFFARX1 I_10873 (I187716,I2859,I187422,I187742,);
nor I_10874 (I187390,I187742,I187646);
not I_10875 (I187764,I187742);
nor I_10876 (I187781,I187764,I187555);
nor I_10877 (I187798,I187487,I187781);
DFFARX1 I_10878 (I187798,I2859,I187422,I187405,);
nor I_10879 (I187829,I187764,I187646);
nor I_10880 (I187846,I57378,I57369);
nor I_10881 (I187396,I187846,I187829);
not I_10882 (I187877,I187846);
nand I_10883 (I187399,I187606,I187877);
DFFARX1 I_10884 (I187846,I2859,I187422,I187411,);
DFFARX1 I_10885 (I187846,I2859,I187422,I187408,);
not I_10886 (I187966,I2866);
DFFARX1 I_10887 (I18895,I2859,I187966,I187992,);
DFFARX1 I_10888 (I187992,I2859,I187966,I188009,);
not I_10889 (I187958,I188009);
not I_10890 (I188031,I187992);
nand I_10891 (I188048,I18883,I18898);
and I_10892 (I188065,I188048,I18886);
DFFARX1 I_10893 (I188065,I2859,I187966,I188091,);
not I_10894 (I188099,I188091);
DFFARX1 I_10895 (I18907,I2859,I187966,I188125,);
and I_10896 (I188133,I188125,I18901);
nand I_10897 (I188150,I188125,I18901);
nand I_10898 (I187937,I188099,I188150);
DFFARX1 I_10899 (I18904,I2859,I187966,I188190,);
nor I_10900 (I188198,I188190,I188133);
DFFARX1 I_10901 (I188198,I2859,I187966,I187931,);
nor I_10902 (I187946,I188190,I188091);
nand I_10903 (I188243,I18883,I18886);
and I_10904 (I188260,I188243,I18889);
DFFARX1 I_10905 (I188260,I2859,I187966,I188286,);
nor I_10906 (I187934,I188286,I188190);
not I_10907 (I188308,I188286);
nor I_10908 (I188325,I188308,I188099);
nor I_10909 (I188342,I188031,I188325);
DFFARX1 I_10910 (I188342,I2859,I187966,I187949,);
nor I_10911 (I188373,I188308,I188190);
nor I_10912 (I188390,I18892,I18886);
nor I_10913 (I187940,I188390,I188373);
not I_10914 (I188421,I188390);
nand I_10915 (I187943,I188150,I188421);
DFFARX1 I_10916 (I188390,I2859,I187966,I187955,);
DFFARX1 I_10917 (I188390,I2859,I187966,I187952,);
not I_10918 (I188510,I2866);
DFFARX1 I_10919 (I111367,I2859,I188510,I188536,);
DFFARX1 I_10920 (I188536,I2859,I188510,I188553,);
not I_10921 (I188502,I188553);
not I_10922 (I188575,I188536);
nand I_10923 (I188592,I111346,I111370);
and I_10924 (I188609,I188592,I111373);
DFFARX1 I_10925 (I188609,I2859,I188510,I188635,);
not I_10926 (I188643,I188635);
DFFARX1 I_10927 (I111355,I2859,I188510,I188669,);
and I_10928 (I188677,I188669,I111361);
nand I_10929 (I188694,I188669,I111361);
nand I_10930 (I188481,I188643,I188694);
DFFARX1 I_10931 (I111349,I2859,I188510,I188734,);
nor I_10932 (I188742,I188734,I188677);
DFFARX1 I_10933 (I188742,I2859,I188510,I188475,);
nor I_10934 (I188490,I188734,I188635);
nand I_10935 (I188787,I111358,I111346);
and I_10936 (I188804,I188787,I111352);
DFFARX1 I_10937 (I188804,I2859,I188510,I188830,);
nor I_10938 (I188478,I188830,I188734);
not I_10939 (I188852,I188830);
nor I_10940 (I188869,I188852,I188643);
nor I_10941 (I188886,I188575,I188869);
DFFARX1 I_10942 (I188886,I2859,I188510,I188493,);
nor I_10943 (I188917,I188852,I188734);
nor I_10944 (I188934,I111364,I111346);
nor I_10945 (I188484,I188934,I188917);
not I_10946 (I188965,I188934);
nand I_10947 (I188487,I188694,I188965);
DFFARX1 I_10948 (I188934,I2859,I188510,I188499,);
DFFARX1 I_10949 (I188934,I2859,I188510,I188496,);
not I_10950 (I189054,I2866);
DFFARX1 I_10951 (I60800,I2859,I189054,I189080,);
DFFARX1 I_10952 (I189080,I2859,I189054,I189097,);
not I_10953 (I189046,I189097);
not I_10954 (I189119,I189080);
nand I_10955 (I189136,I60809,I60812);
and I_10956 (I189153,I189136,I60791);
DFFARX1 I_10957 (I189153,I2859,I189054,I189179,);
not I_10958 (I189187,I189179);
DFFARX1 I_10959 (I60806,I2859,I189054,I189213,);
and I_10960 (I189221,I189213,I60794);
nand I_10961 (I189238,I189213,I60794);
nand I_10962 (I189025,I189187,I189238);
DFFARX1 I_10963 (I60788,I2859,I189054,I189278,);
nor I_10964 (I189286,I189278,I189221);
DFFARX1 I_10965 (I189286,I2859,I189054,I189019,);
nor I_10966 (I189034,I189278,I189179);
nand I_10967 (I189331,I60803,I60797);
and I_10968 (I189348,I189331,I60788);
DFFARX1 I_10969 (I189348,I2859,I189054,I189374,);
nor I_10970 (I189022,I189374,I189278);
not I_10971 (I189396,I189374);
nor I_10972 (I189413,I189396,I189187);
nor I_10973 (I189430,I189119,I189413);
DFFARX1 I_10974 (I189430,I2859,I189054,I189037,);
nor I_10975 (I189461,I189396,I189278);
nor I_10976 (I189478,I60815,I60797);
nor I_10977 (I189028,I189478,I189461);
not I_10978 (I189509,I189478);
nand I_10979 (I189031,I189238,I189509);
DFFARX1 I_10980 (I189478,I2859,I189054,I189043,);
DFFARX1 I_10981 (I189478,I2859,I189054,I189040,);
not I_10982 (I189598,I2866);
DFFARX1 I_10983 (I402885,I2859,I189598,I189624,);
DFFARX1 I_10984 (I189624,I2859,I189598,I189641,);
not I_10985 (I189590,I189641);
not I_10986 (I189663,I189624);
nand I_10987 (I189680,I402900,I402888);
and I_10988 (I189697,I189680,I402879);
DFFARX1 I_10989 (I189697,I2859,I189598,I189723,);
not I_10990 (I189731,I189723);
DFFARX1 I_10991 (I402891,I2859,I189598,I189757,);
and I_10992 (I189765,I189757,I402882);
nand I_10993 (I189782,I189757,I402882);
nand I_10994 (I189569,I189731,I189782);
DFFARX1 I_10995 (I402897,I2859,I189598,I189822,);
nor I_10996 (I189830,I189822,I189765);
DFFARX1 I_10997 (I189830,I2859,I189598,I189563,);
nor I_10998 (I189578,I189822,I189723);
nand I_10999 (I189875,I402906,I402894);
and I_11000 (I189892,I189875,I402903);
DFFARX1 I_11001 (I189892,I2859,I189598,I189918,);
nor I_11002 (I189566,I189918,I189822);
not I_11003 (I189940,I189918);
nor I_11004 (I189957,I189940,I189731);
nor I_11005 (I189974,I189663,I189957);
DFFARX1 I_11006 (I189974,I2859,I189598,I189581,);
nor I_11007 (I190005,I189940,I189822);
nor I_11008 (I190022,I402879,I402894);
nor I_11009 (I189572,I190022,I190005);
not I_11010 (I190053,I190022);
nand I_11011 (I189575,I189782,I190053);
DFFARX1 I_11012 (I190022,I2859,I189598,I189587,);
DFFARX1 I_11013 (I190022,I2859,I189598,I189584,);
not I_11014 (I190142,I2866);
DFFARX1 I_11015 (I220251,I2859,I190142,I190168,);
DFFARX1 I_11016 (I190168,I2859,I190142,I190185,);
not I_11017 (I190134,I190185);
not I_11018 (I190207,I190168);
nand I_11019 (I190224,I220254,I220272);
and I_11020 (I190241,I190224,I220260);
DFFARX1 I_11021 (I190241,I2859,I190142,I190267,);
not I_11022 (I190275,I190267);
DFFARX1 I_11023 (I220251,I2859,I190142,I190301,);
and I_11024 (I190309,I190301,I220269);
nand I_11025 (I190326,I190301,I220269);
nand I_11026 (I190113,I190275,I190326);
DFFARX1 I_11027 (I220263,I2859,I190142,I190366,);
nor I_11028 (I190374,I190366,I190309);
DFFARX1 I_11029 (I190374,I2859,I190142,I190107,);
nor I_11030 (I190122,I190366,I190267);
nand I_11031 (I190419,I220266,I220248);
and I_11032 (I190436,I190419,I220257);
DFFARX1 I_11033 (I190436,I2859,I190142,I190462,);
nor I_11034 (I190110,I190462,I190366);
not I_11035 (I190484,I190462);
nor I_11036 (I190501,I190484,I190275);
nor I_11037 (I190518,I190207,I190501);
DFFARX1 I_11038 (I190518,I2859,I190142,I190125,);
nor I_11039 (I190549,I190484,I190366);
nor I_11040 (I190566,I220248,I220248);
nor I_11041 (I190116,I190566,I190549);
not I_11042 (I190597,I190566);
nand I_11043 (I190119,I190326,I190597);
DFFARX1 I_11044 (I190566,I2859,I190142,I190131,);
DFFARX1 I_11045 (I190566,I2859,I190142,I190128,);
not I_11046 (I190686,I2866);
DFFARX1 I_11047 (I541337,I2859,I190686,I190712,);
DFFARX1 I_11048 (I190712,I2859,I190686,I190729,);
not I_11049 (I190678,I190729);
not I_11050 (I190751,I190712);
nand I_11051 (I190768,I541313,I541334);
and I_11052 (I190785,I190768,I541331);
DFFARX1 I_11053 (I190785,I2859,I190686,I190811,);
not I_11054 (I190819,I190811);
DFFARX1 I_11055 (I541310,I2859,I190686,I190845,);
and I_11056 (I190853,I190845,I541322);
nand I_11057 (I190870,I190845,I541322);
nand I_11058 (I190657,I190819,I190870);
DFFARX1 I_11059 (I541325,I2859,I190686,I190910,);
nor I_11060 (I190918,I190910,I190853);
DFFARX1 I_11061 (I190918,I2859,I190686,I190651,);
nor I_11062 (I190666,I190910,I190811);
nand I_11063 (I190963,I541328,I541316);
and I_11064 (I190980,I190963,I541319);
DFFARX1 I_11065 (I190980,I2859,I190686,I191006,);
nor I_11066 (I190654,I191006,I190910);
not I_11067 (I191028,I191006);
nor I_11068 (I191045,I191028,I190819);
nor I_11069 (I191062,I190751,I191045);
DFFARX1 I_11070 (I191062,I2859,I190686,I190669,);
nor I_11071 (I191093,I191028,I190910);
nor I_11072 (I191110,I541310,I541316);
nor I_11073 (I190660,I191110,I191093);
not I_11074 (I191141,I191110);
nand I_11075 (I190663,I190870,I191141);
DFFARX1 I_11076 (I191110,I2859,I190686,I190675,);
DFFARX1 I_11077 (I191110,I2859,I190686,I190672,);
not I_11078 (I191230,I2866);
DFFARX1 I_11079 (I523444,I2859,I191230,I191256,);
DFFARX1 I_11080 (I191256,I2859,I191230,I191273,);
not I_11081 (I191222,I191273);
not I_11082 (I191295,I191256);
nand I_11083 (I191312,I523441,I523438);
and I_11084 (I191329,I191312,I523426);
DFFARX1 I_11085 (I191329,I2859,I191230,I191355,);
not I_11086 (I191363,I191355);
DFFARX1 I_11087 (I523450,I2859,I191230,I191389,);
and I_11088 (I191397,I191389,I523435);
nand I_11089 (I191414,I191389,I523435);
nand I_11090 (I191201,I191363,I191414);
DFFARX1 I_11091 (I523429,I2859,I191230,I191454,);
nor I_11092 (I191462,I191454,I191397);
DFFARX1 I_11093 (I191462,I2859,I191230,I191195,);
nor I_11094 (I191210,I191454,I191355);
nand I_11095 (I191507,I523426,I523432);
and I_11096 (I191524,I191507,I523447);
DFFARX1 I_11097 (I191524,I2859,I191230,I191550,);
nor I_11098 (I191198,I191550,I191454);
not I_11099 (I191572,I191550);
nor I_11100 (I191589,I191572,I191363);
nor I_11101 (I191606,I191295,I191589);
DFFARX1 I_11102 (I191606,I2859,I191230,I191213,);
nor I_11103 (I191637,I191572,I191454);
nor I_11104 (I191654,I523429,I523432);
nor I_11105 (I191204,I191654,I191637);
not I_11106 (I191685,I191654);
nand I_11107 (I191207,I191414,I191685);
DFFARX1 I_11108 (I191654,I2859,I191230,I191219,);
DFFARX1 I_11109 (I191654,I2859,I191230,I191216,);
not I_11110 (I191774,I2866);
DFFARX1 I_11111 (I409991,I2859,I191774,I191800,);
DFFARX1 I_11112 (I191800,I2859,I191774,I191817,);
not I_11113 (I191766,I191817);
not I_11114 (I191839,I191800);
nand I_11115 (I191856,I410006,I409994);
and I_11116 (I191873,I191856,I409985);
DFFARX1 I_11117 (I191873,I2859,I191774,I191899,);
not I_11118 (I191907,I191899);
DFFARX1 I_11119 (I409997,I2859,I191774,I191933,);
and I_11120 (I191941,I191933,I409988);
nand I_11121 (I191958,I191933,I409988);
nand I_11122 (I191745,I191907,I191958);
DFFARX1 I_11123 (I410003,I2859,I191774,I191998,);
nor I_11124 (I192006,I191998,I191941);
DFFARX1 I_11125 (I192006,I2859,I191774,I191739,);
nor I_11126 (I191754,I191998,I191899);
nand I_11127 (I192051,I410012,I410000);
and I_11128 (I192068,I192051,I410009);
DFFARX1 I_11129 (I192068,I2859,I191774,I192094,);
nor I_11130 (I191742,I192094,I191998);
not I_11131 (I192116,I192094);
nor I_11132 (I192133,I192116,I191907);
nor I_11133 (I192150,I191839,I192133);
DFFARX1 I_11134 (I192150,I2859,I191774,I191757,);
nor I_11135 (I192181,I192116,I191998);
nor I_11136 (I192198,I409985,I410000);
nor I_11137 (I191748,I192198,I192181);
not I_11138 (I192229,I192198);
nand I_11139 (I191751,I191958,I192229);
DFFARX1 I_11140 (I192198,I2859,I191774,I191763,);
DFFARX1 I_11141 (I192198,I2859,I191774,I191760,);
not I_11142 (I192318,I2866);
DFFARX1 I_11143 (I130339,I2859,I192318,I192344,);
DFFARX1 I_11144 (I192344,I2859,I192318,I192361,);
not I_11145 (I192310,I192361);
not I_11146 (I192383,I192344);
nand I_11147 (I192400,I130318,I130342);
and I_11148 (I192417,I192400,I130345);
DFFARX1 I_11149 (I192417,I2859,I192318,I192443,);
not I_11150 (I192451,I192443);
DFFARX1 I_11151 (I130327,I2859,I192318,I192477,);
and I_11152 (I192485,I192477,I130333);
nand I_11153 (I192502,I192477,I130333);
nand I_11154 (I192289,I192451,I192502);
DFFARX1 I_11155 (I130321,I2859,I192318,I192542,);
nor I_11156 (I192550,I192542,I192485);
DFFARX1 I_11157 (I192550,I2859,I192318,I192283,);
nor I_11158 (I192298,I192542,I192443);
nand I_11159 (I192595,I130330,I130318);
and I_11160 (I192612,I192595,I130324);
DFFARX1 I_11161 (I192612,I2859,I192318,I192638,);
nor I_11162 (I192286,I192638,I192542);
not I_11163 (I192660,I192638);
nor I_11164 (I192677,I192660,I192451);
nor I_11165 (I192694,I192383,I192677);
DFFARX1 I_11166 (I192694,I2859,I192318,I192301,);
nor I_11167 (I192725,I192660,I192542);
nor I_11168 (I192742,I130336,I130318);
nor I_11169 (I192292,I192742,I192725);
not I_11170 (I192773,I192742);
nand I_11171 (I192295,I192502,I192773);
DFFARX1 I_11172 (I192742,I2859,I192318,I192307,);
DFFARX1 I_11173 (I192742,I2859,I192318,I192304,);
not I_11174 (I192862,I2866);
DFFARX1 I_11175 (I32064,I2859,I192862,I192888,);
DFFARX1 I_11176 (I192888,I2859,I192862,I192905,);
not I_11177 (I192854,I192905);
not I_11178 (I192927,I192888);
nand I_11179 (I192944,I32079,I32058);
and I_11180 (I192961,I192944,I32061);
DFFARX1 I_11181 (I192961,I2859,I192862,I192987,);
not I_11182 (I192995,I192987);
DFFARX1 I_11183 (I32067,I2859,I192862,I193021,);
and I_11184 (I193029,I193021,I32061);
nand I_11185 (I193046,I193021,I32061);
nand I_11186 (I192833,I192995,I193046);
DFFARX1 I_11187 (I32076,I2859,I192862,I193086,);
nor I_11188 (I193094,I193086,I193029);
DFFARX1 I_11189 (I193094,I2859,I192862,I192827,);
nor I_11190 (I192842,I193086,I192987);
nand I_11191 (I193139,I32058,I32073);
and I_11192 (I193156,I193139,I32070);
DFFARX1 I_11193 (I193156,I2859,I192862,I193182,);
nor I_11194 (I192830,I193182,I193086);
not I_11195 (I193204,I193182);
nor I_11196 (I193221,I193204,I192995);
nor I_11197 (I193238,I192927,I193221);
DFFARX1 I_11198 (I193238,I2859,I192862,I192845,);
nor I_11199 (I193269,I193204,I193086);
nor I_11200 (I193286,I32082,I32073);
nor I_11201 (I192836,I193286,I193269);
not I_11202 (I193317,I193286);
nand I_11203 (I192839,I193046,I193317);
DFFARX1 I_11204 (I193286,I2859,I192862,I192851,);
DFFARX1 I_11205 (I193286,I2859,I192862,I192848,);
not I_11206 (I193406,I2866);
DFFARX1 I_11207 (I252313,I2859,I193406,I193432,);
DFFARX1 I_11208 (I193432,I2859,I193406,I193449,);
not I_11209 (I193398,I193449);
not I_11210 (I193471,I193432);
nand I_11211 (I193488,I252310,I252331);
and I_11212 (I193505,I193488,I252334);
DFFARX1 I_11213 (I193505,I2859,I193406,I193531,);
not I_11214 (I193539,I193531);
DFFARX1 I_11215 (I252319,I2859,I193406,I193565,);
and I_11216 (I193573,I193565,I252322);
nand I_11217 (I193590,I193565,I252322);
nand I_11218 (I193377,I193539,I193590);
DFFARX1 I_11219 (I252325,I2859,I193406,I193630,);
nor I_11220 (I193638,I193630,I193573);
DFFARX1 I_11221 (I193638,I2859,I193406,I193371,);
nor I_11222 (I193386,I193630,I193531);
nand I_11223 (I193683,I252310,I252316);
and I_11224 (I193700,I193683,I252328);
DFFARX1 I_11225 (I193700,I2859,I193406,I193726,);
nor I_11226 (I193374,I193726,I193630);
not I_11227 (I193748,I193726);
nor I_11228 (I193765,I193748,I193539);
nor I_11229 (I193782,I193471,I193765);
DFFARX1 I_11230 (I193782,I2859,I193406,I193389,);
nor I_11231 (I193813,I193748,I193630);
nor I_11232 (I193830,I252313,I252316);
nor I_11233 (I193380,I193830,I193813);
not I_11234 (I193861,I193830);
nand I_11235 (I193383,I193590,I193861);
DFFARX1 I_11236 (I193830,I2859,I193406,I193395,);
DFFARX1 I_11237 (I193830,I2859,I193406,I193392,);
not I_11238 (I193950,I2866);
DFFARX1 I_11239 (I395779,I2859,I193950,I193976,);
DFFARX1 I_11240 (I193976,I2859,I193950,I193993,);
not I_11241 (I193942,I193993);
not I_11242 (I194015,I193976);
nand I_11243 (I194032,I395794,I395782);
and I_11244 (I194049,I194032,I395773);
DFFARX1 I_11245 (I194049,I2859,I193950,I194075,);
not I_11246 (I194083,I194075);
DFFARX1 I_11247 (I395785,I2859,I193950,I194109,);
and I_11248 (I194117,I194109,I395776);
nand I_11249 (I194134,I194109,I395776);
nand I_11250 (I193921,I194083,I194134);
DFFARX1 I_11251 (I395791,I2859,I193950,I194174,);
nor I_11252 (I194182,I194174,I194117);
DFFARX1 I_11253 (I194182,I2859,I193950,I193915,);
nor I_11254 (I193930,I194174,I194075);
nand I_11255 (I194227,I395800,I395788);
and I_11256 (I194244,I194227,I395797);
DFFARX1 I_11257 (I194244,I2859,I193950,I194270,);
nor I_11258 (I193918,I194270,I194174);
not I_11259 (I194292,I194270);
nor I_11260 (I194309,I194292,I194083);
nor I_11261 (I194326,I194015,I194309);
DFFARX1 I_11262 (I194326,I2859,I193950,I193933,);
nor I_11263 (I194357,I194292,I194174);
nor I_11264 (I194374,I395773,I395788);
nor I_11265 (I193924,I194374,I194357);
not I_11266 (I194405,I194374);
nand I_11267 (I193927,I194134,I194405);
DFFARX1 I_11268 (I194374,I2859,I193950,I193939,);
DFFARX1 I_11269 (I194374,I2859,I193950,I193936,);
not I_11270 (I194494,I2866);
DFFARX1 I_11271 (I241909,I2859,I194494,I194520,);
DFFARX1 I_11272 (I194520,I2859,I194494,I194537,);
not I_11273 (I194486,I194537);
not I_11274 (I194559,I194520);
nand I_11275 (I194576,I241906,I241927);
and I_11276 (I194593,I194576,I241930);
DFFARX1 I_11277 (I194593,I2859,I194494,I194619,);
not I_11278 (I194627,I194619);
DFFARX1 I_11279 (I241915,I2859,I194494,I194653,);
and I_11280 (I194661,I194653,I241918);
nand I_11281 (I194678,I194653,I241918);
nand I_11282 (I194465,I194627,I194678);
DFFARX1 I_11283 (I241921,I2859,I194494,I194718,);
nor I_11284 (I194726,I194718,I194661);
DFFARX1 I_11285 (I194726,I2859,I194494,I194459,);
nor I_11286 (I194474,I194718,I194619);
nand I_11287 (I194771,I241906,I241912);
and I_11288 (I194788,I194771,I241924);
DFFARX1 I_11289 (I194788,I2859,I194494,I194814,);
nor I_11290 (I194462,I194814,I194718);
not I_11291 (I194836,I194814);
nor I_11292 (I194853,I194836,I194627);
nor I_11293 (I194870,I194559,I194853);
DFFARX1 I_11294 (I194870,I2859,I194494,I194477,);
nor I_11295 (I194901,I194836,I194718);
nor I_11296 (I194918,I241909,I241912);
nor I_11297 (I194468,I194918,I194901);
not I_11298 (I194949,I194918);
nand I_11299 (I194471,I194678,I194949);
DFFARX1 I_11300 (I194918,I2859,I194494,I194483,);
DFFARX1 I_11301 (I194918,I2859,I194494,I194480,);
not I_11302 (I195038,I2866);
DFFARX1 I_11303 (I346893,I2859,I195038,I195064,);
DFFARX1 I_11304 (I195064,I2859,I195038,I195081,);
not I_11305 (I195030,I195081);
not I_11306 (I195103,I195064);
nand I_11307 (I195120,I346887,I346884);
and I_11308 (I195137,I195120,I346899);
DFFARX1 I_11309 (I195137,I2859,I195038,I195163,);
not I_11310 (I195171,I195163);
DFFARX1 I_11311 (I346887,I2859,I195038,I195197,);
and I_11312 (I195205,I195197,I346881);
nand I_11313 (I195222,I195197,I346881);
nand I_11314 (I195009,I195171,I195222);
DFFARX1 I_11315 (I346881,I2859,I195038,I195262,);
nor I_11316 (I195270,I195262,I195205);
DFFARX1 I_11317 (I195270,I2859,I195038,I195003,);
nor I_11318 (I195018,I195262,I195163);
nand I_11319 (I195315,I346896,I346890);
and I_11320 (I195332,I195315,I346884);
DFFARX1 I_11321 (I195332,I2859,I195038,I195358,);
nor I_11322 (I195006,I195358,I195262);
not I_11323 (I195380,I195358);
nor I_11324 (I195397,I195380,I195171);
nor I_11325 (I195414,I195103,I195397);
DFFARX1 I_11326 (I195414,I2859,I195038,I195021,);
nor I_11327 (I195445,I195380,I195262);
nor I_11328 (I195462,I346902,I346890);
nor I_11329 (I195012,I195462,I195445);
not I_11330 (I195493,I195462);
nand I_11331 (I195015,I195222,I195493);
DFFARX1 I_11332 (I195462,I2859,I195038,I195027,);
DFFARX1 I_11333 (I195462,I2859,I195038,I195024,);
not I_11334 (I195582,I2866);
DFFARX1 I_11335 (I294507,I2859,I195582,I195608,);
DFFARX1 I_11336 (I195608,I2859,I195582,I195625,);
not I_11337 (I195574,I195625);
not I_11338 (I195647,I195608);
nand I_11339 (I195664,I294528,I294519);
and I_11340 (I195681,I195664,I294507);
DFFARX1 I_11341 (I195681,I2859,I195582,I195707,);
not I_11342 (I195715,I195707);
DFFARX1 I_11343 (I294513,I2859,I195582,I195741,);
and I_11344 (I195749,I195741,I294510);
nand I_11345 (I195766,I195741,I294510);
nand I_11346 (I195553,I195715,I195766);
DFFARX1 I_11347 (I294504,I2859,I195582,I195806,);
nor I_11348 (I195814,I195806,I195749);
DFFARX1 I_11349 (I195814,I2859,I195582,I195547,);
nor I_11350 (I195562,I195806,I195707);
nand I_11351 (I195859,I294504,I294516);
and I_11352 (I195876,I195859,I294525);
DFFARX1 I_11353 (I195876,I2859,I195582,I195902,);
nor I_11354 (I195550,I195902,I195806);
not I_11355 (I195924,I195902);
nor I_11356 (I195941,I195924,I195715);
nor I_11357 (I195958,I195647,I195941);
DFFARX1 I_11358 (I195958,I2859,I195582,I195565,);
nor I_11359 (I195989,I195924,I195806);
nor I_11360 (I196006,I294522,I294516);
nor I_11361 (I195556,I196006,I195989);
not I_11362 (I196037,I196006);
nand I_11363 (I195559,I195766,I196037);
DFFARX1 I_11364 (I196006,I2859,I195582,I195571,);
DFFARX1 I_11365 (I196006,I2859,I195582,I195568,);
not I_11366 (I196126,I2866);
DFFARX1 I_11367 (I467975,I2859,I196126,I196152,);
DFFARX1 I_11368 (I196152,I2859,I196126,I196169,);
not I_11369 (I196118,I196169);
not I_11370 (I196191,I196152);
nand I_11371 (I196208,I467987,I467975);
and I_11372 (I196225,I196208,I467978);
DFFARX1 I_11373 (I196225,I2859,I196126,I196251,);
not I_11374 (I196259,I196251);
DFFARX1 I_11375 (I467996,I2859,I196126,I196285,);
and I_11376 (I196293,I196285,I467972);
nand I_11377 (I196310,I196285,I467972);
nand I_11378 (I196097,I196259,I196310);
DFFARX1 I_11379 (I467990,I2859,I196126,I196350,);
nor I_11380 (I196358,I196350,I196293);
DFFARX1 I_11381 (I196358,I2859,I196126,I196091,);
nor I_11382 (I196106,I196350,I196251);
nand I_11383 (I196403,I467984,I467981);
and I_11384 (I196420,I196403,I467993);
DFFARX1 I_11385 (I196420,I2859,I196126,I196446,);
nor I_11386 (I196094,I196446,I196350);
not I_11387 (I196468,I196446);
nor I_11388 (I196485,I196468,I196259);
nor I_11389 (I196502,I196191,I196485);
DFFARX1 I_11390 (I196502,I2859,I196126,I196109,);
nor I_11391 (I196533,I196468,I196350);
nor I_11392 (I196550,I467972,I467981);
nor I_11393 (I196100,I196550,I196533);
not I_11394 (I196581,I196550);
nand I_11395 (I196103,I196310,I196581);
DFFARX1 I_11396 (I196550,I2859,I196126,I196115,);
DFFARX1 I_11397 (I196550,I2859,I196126,I196112,);
not I_11398 (I196670,I2866);
DFFARX1 I_11399 (I111894,I2859,I196670,I196696,);
DFFARX1 I_11400 (I196696,I2859,I196670,I196713,);
not I_11401 (I196662,I196713);
not I_11402 (I196735,I196696);
nand I_11403 (I196752,I111873,I111897);
and I_11404 (I196769,I196752,I111900);
DFFARX1 I_11405 (I196769,I2859,I196670,I196795,);
not I_11406 (I196803,I196795);
DFFARX1 I_11407 (I111882,I2859,I196670,I196829,);
and I_11408 (I196837,I196829,I111888);
nand I_11409 (I196854,I196829,I111888);
nand I_11410 (I196641,I196803,I196854);
DFFARX1 I_11411 (I111876,I2859,I196670,I196894,);
nor I_11412 (I196902,I196894,I196837);
DFFARX1 I_11413 (I196902,I2859,I196670,I196635,);
nor I_11414 (I196650,I196894,I196795);
nand I_11415 (I196947,I111885,I111873);
and I_11416 (I196964,I196947,I111879);
DFFARX1 I_11417 (I196964,I2859,I196670,I196990,);
nor I_11418 (I196638,I196990,I196894);
not I_11419 (I197012,I196990);
nor I_11420 (I197029,I197012,I196803);
nor I_11421 (I197046,I196735,I197029);
DFFARX1 I_11422 (I197046,I2859,I196670,I196653,);
nor I_11423 (I197077,I197012,I196894);
nor I_11424 (I197094,I111891,I111873);
nor I_11425 (I196644,I197094,I197077);
not I_11426 (I197125,I197094);
nand I_11427 (I196647,I196854,I197125);
DFFARX1 I_11428 (I197094,I2859,I196670,I196659,);
DFFARX1 I_11429 (I197094,I2859,I196670,I196656,);
not I_11430 (I197214,I2866);
DFFARX1 I_11431 (I531536,I2859,I197214,I197240,);
DFFARX1 I_11432 (I197240,I2859,I197214,I197257,);
not I_11433 (I197206,I197257);
not I_11434 (I197279,I197240);
nand I_11435 (I197296,I531533,I531530);
and I_11436 (I197313,I197296,I531518);
DFFARX1 I_11437 (I197313,I2859,I197214,I197339,);
not I_11438 (I197347,I197339);
DFFARX1 I_11439 (I531542,I2859,I197214,I197373,);
and I_11440 (I197381,I197373,I531527);
nand I_11441 (I197398,I197373,I531527);
nand I_11442 (I197185,I197347,I197398);
DFFARX1 I_11443 (I531521,I2859,I197214,I197438,);
nor I_11444 (I197446,I197438,I197381);
DFFARX1 I_11445 (I197446,I2859,I197214,I197179,);
nor I_11446 (I197194,I197438,I197339);
nand I_11447 (I197491,I531518,I531524);
and I_11448 (I197508,I197491,I531539);
DFFARX1 I_11449 (I197508,I2859,I197214,I197534,);
nor I_11450 (I197182,I197534,I197438);
not I_11451 (I197556,I197534);
nor I_11452 (I197573,I197556,I197347);
nor I_11453 (I197590,I197279,I197573);
DFFARX1 I_11454 (I197590,I2859,I197214,I197197,);
nor I_11455 (I197621,I197556,I197438);
nor I_11456 (I197638,I531521,I531524);
nor I_11457 (I197188,I197638,I197621);
not I_11458 (I197669,I197638);
nand I_11459 (I197191,I197398,I197669);
DFFARX1 I_11460 (I197638,I2859,I197214,I197203,);
DFFARX1 I_11461 (I197638,I2859,I197214,I197200,);
not I_11462 (I197758,I2866);
DFFARX1 I_11463 (I350582,I2859,I197758,I197784,);
DFFARX1 I_11464 (I197784,I2859,I197758,I197801,);
not I_11465 (I197750,I197801);
not I_11466 (I197823,I197784);
nand I_11467 (I197840,I350576,I350573);
and I_11468 (I197857,I197840,I350588);
DFFARX1 I_11469 (I197857,I2859,I197758,I197883,);
not I_11470 (I197891,I197883);
DFFARX1 I_11471 (I350576,I2859,I197758,I197917,);
and I_11472 (I197925,I197917,I350570);
nand I_11473 (I197942,I197917,I350570);
nand I_11474 (I197729,I197891,I197942);
DFFARX1 I_11475 (I350570,I2859,I197758,I197982,);
nor I_11476 (I197990,I197982,I197925);
DFFARX1 I_11477 (I197990,I2859,I197758,I197723,);
nor I_11478 (I197738,I197982,I197883);
nand I_11479 (I198035,I350585,I350579);
and I_11480 (I198052,I198035,I350573);
DFFARX1 I_11481 (I198052,I2859,I197758,I198078,);
nor I_11482 (I197726,I198078,I197982);
not I_11483 (I198100,I198078);
nor I_11484 (I198117,I198100,I197891);
nor I_11485 (I198134,I197823,I198117);
DFFARX1 I_11486 (I198134,I2859,I197758,I197741,);
nor I_11487 (I198165,I198100,I197982);
nor I_11488 (I198182,I350591,I350579);
nor I_11489 (I197732,I198182,I198165);
not I_11490 (I198213,I198182);
nand I_11491 (I197735,I197942,I198213);
DFFARX1 I_11492 (I198182,I2859,I197758,I197747,);
DFFARX1 I_11493 (I198182,I2859,I197758,I197744,);
not I_11494 (I198302,I2866);
DFFARX1 I_11495 (I322829,I2859,I198302,I198328,);
DFFARX1 I_11496 (I198328,I2859,I198302,I198345,);
not I_11497 (I198294,I198345);
not I_11498 (I198367,I198328);
nand I_11499 (I198384,I322850,I322841);
and I_11500 (I198401,I198384,I322829);
DFFARX1 I_11501 (I198401,I2859,I198302,I198427,);
not I_11502 (I198435,I198427);
DFFARX1 I_11503 (I322835,I2859,I198302,I198461,);
and I_11504 (I198469,I198461,I322832);
nand I_11505 (I198486,I198461,I322832);
nand I_11506 (I198273,I198435,I198486);
DFFARX1 I_11507 (I322826,I2859,I198302,I198526,);
nor I_11508 (I198534,I198526,I198469);
DFFARX1 I_11509 (I198534,I2859,I198302,I198267,);
nor I_11510 (I198282,I198526,I198427);
nand I_11511 (I198579,I322826,I322838);
and I_11512 (I198596,I198579,I322847);
DFFARX1 I_11513 (I198596,I2859,I198302,I198622,);
nor I_11514 (I198270,I198622,I198526);
not I_11515 (I198644,I198622);
nor I_11516 (I198661,I198644,I198435);
nor I_11517 (I198678,I198367,I198661);
DFFARX1 I_11518 (I198678,I2859,I198302,I198285,);
nor I_11519 (I198709,I198644,I198526);
nor I_11520 (I198726,I322844,I322838);
nor I_11521 (I198276,I198726,I198709);
not I_11522 (I198757,I198726);
nand I_11523 (I198279,I198486,I198757);
DFFARX1 I_11524 (I198726,I2859,I198302,I198291,);
DFFARX1 I_11525 (I198726,I2859,I198302,I198288,);
not I_11526 (I198846,I2866);
DFFARX1 I_11527 (I79837,I2859,I198846,I198872,);
DFFARX1 I_11528 (I198872,I2859,I198846,I198889,);
not I_11529 (I198838,I198889);
not I_11530 (I198911,I198872);
nand I_11531 (I198928,I79849,I79828);
and I_11532 (I198945,I198928,I79831);
DFFARX1 I_11533 (I198945,I2859,I198846,I198971,);
not I_11534 (I198979,I198971);
DFFARX1 I_11535 (I79840,I2859,I198846,I199005,);
and I_11536 (I199013,I199005,I79852);
nand I_11537 (I199030,I199005,I79852);
nand I_11538 (I198817,I198979,I199030);
DFFARX1 I_11539 (I79846,I2859,I198846,I199070,);
nor I_11540 (I199078,I199070,I199013);
DFFARX1 I_11541 (I199078,I2859,I198846,I198811,);
nor I_11542 (I198826,I199070,I198971);
nand I_11543 (I199123,I79834,I79831);
and I_11544 (I199140,I199123,I79843);
DFFARX1 I_11545 (I199140,I2859,I198846,I199166,);
nor I_11546 (I198814,I199166,I199070);
not I_11547 (I199188,I199166);
nor I_11548 (I199205,I199188,I198979);
nor I_11549 (I199222,I198911,I199205);
DFFARX1 I_11550 (I199222,I2859,I198846,I198829,);
nor I_11551 (I199253,I199188,I199070);
nor I_11552 (I199270,I79828,I79831);
nor I_11553 (I198820,I199270,I199253);
not I_11554 (I199301,I199270);
nand I_11555 (I198823,I199030,I199301);
DFFARX1 I_11556 (I199270,I2859,I198846,I198835,);
DFFARX1 I_11557 (I199270,I2859,I198846,I198832,);
not I_11558 (I199390,I2866);
DFFARX1 I_11559 (I27848,I2859,I199390,I199416,);
DFFARX1 I_11560 (I199416,I2859,I199390,I199433,);
not I_11561 (I199382,I199433);
not I_11562 (I199455,I199416);
nand I_11563 (I199472,I27863,I27842);
and I_11564 (I199489,I199472,I27845);
DFFARX1 I_11565 (I199489,I2859,I199390,I199515,);
not I_11566 (I199523,I199515);
DFFARX1 I_11567 (I27851,I2859,I199390,I199549,);
and I_11568 (I199557,I199549,I27845);
nand I_11569 (I199574,I199549,I27845);
nand I_11570 (I199361,I199523,I199574);
DFFARX1 I_11571 (I27860,I2859,I199390,I199614,);
nor I_11572 (I199622,I199614,I199557);
DFFARX1 I_11573 (I199622,I2859,I199390,I199355,);
nor I_11574 (I199370,I199614,I199515);
nand I_11575 (I199667,I27842,I27857);
and I_11576 (I199684,I199667,I27854);
DFFARX1 I_11577 (I199684,I2859,I199390,I199710,);
nor I_11578 (I199358,I199710,I199614);
not I_11579 (I199732,I199710);
nor I_11580 (I199749,I199732,I199523);
nor I_11581 (I199766,I199455,I199749);
DFFARX1 I_11582 (I199766,I2859,I199390,I199373,);
nor I_11583 (I199797,I199732,I199614);
nor I_11584 (I199814,I27866,I27857);
nor I_11585 (I199364,I199814,I199797);
not I_11586 (I199845,I199814);
nand I_11587 (I199367,I199574,I199845);
DFFARX1 I_11588 (I199814,I2859,I199390,I199379,);
DFFARX1 I_11589 (I199814,I2859,I199390,I199376,);
not I_11590 (I199934,I2866);
DFFARX1 I_11591 (I52617,I2859,I199934,I199960,);
DFFARX1 I_11592 (I199960,I2859,I199934,I199977,);
not I_11593 (I199926,I199977);
not I_11594 (I199999,I199960);
nand I_11595 (I200016,I52632,I52611);
and I_11596 (I200033,I200016,I52614);
DFFARX1 I_11597 (I200033,I2859,I199934,I200059,);
not I_11598 (I200067,I200059);
DFFARX1 I_11599 (I52620,I2859,I199934,I200093,);
and I_11600 (I200101,I200093,I52614);
nand I_11601 (I200118,I200093,I52614);
nand I_11602 (I199905,I200067,I200118);
DFFARX1 I_11603 (I52629,I2859,I199934,I200158,);
nor I_11604 (I200166,I200158,I200101);
DFFARX1 I_11605 (I200166,I2859,I199934,I199899,);
nor I_11606 (I199914,I200158,I200059);
nand I_11607 (I200211,I52611,I52626);
and I_11608 (I200228,I200211,I52623);
DFFARX1 I_11609 (I200228,I2859,I199934,I200254,);
nor I_11610 (I199902,I200254,I200158);
not I_11611 (I200276,I200254);
nor I_11612 (I200293,I200276,I200067);
nor I_11613 (I200310,I199999,I200293);
DFFARX1 I_11614 (I200310,I2859,I199934,I199917,);
nor I_11615 (I200341,I200276,I200158);
nor I_11616 (I200358,I52635,I52626);
nor I_11617 (I199908,I200358,I200341);
not I_11618 (I200389,I200358);
nand I_11619 (I199911,I200118,I200389);
DFFARX1 I_11620 (I200358,I2859,I199934,I199923,);
DFFARX1 I_11621 (I200358,I2859,I199934,I199920,);
not I_11622 (I200478,I2866);
DFFARX1 I_11623 (I443271,I2859,I200478,I200504,);
DFFARX1 I_11624 (I200504,I2859,I200478,I200521,);
not I_11625 (I200470,I200521);
not I_11626 (I200543,I200504);
nand I_11627 (I200560,I443271,I443289);
and I_11628 (I200577,I200560,I443283);
DFFARX1 I_11629 (I200577,I2859,I200478,I200603,);
not I_11630 (I200611,I200603);
DFFARX1 I_11631 (I443277,I2859,I200478,I200637,);
and I_11632 (I200645,I200637,I443286);
nand I_11633 (I200662,I200637,I443286);
nand I_11634 (I200449,I200611,I200662);
DFFARX1 I_11635 (I443274,I2859,I200478,I200702,);
nor I_11636 (I200710,I200702,I200645);
DFFARX1 I_11637 (I200710,I2859,I200478,I200443,);
nor I_11638 (I200458,I200702,I200603);
nand I_11639 (I200755,I443274,I443292);
and I_11640 (I200772,I200755,I443277);
DFFARX1 I_11641 (I200772,I2859,I200478,I200798,);
nor I_11642 (I200446,I200798,I200702);
not I_11643 (I200820,I200798);
nor I_11644 (I200837,I200820,I200611);
nor I_11645 (I200854,I200543,I200837);
DFFARX1 I_11646 (I200854,I2859,I200478,I200461,);
nor I_11647 (I200885,I200820,I200702);
nor I_11648 (I200902,I443280,I443292);
nor I_11649 (I200452,I200902,I200885);
not I_11650 (I200933,I200902);
nand I_11651 (I200455,I200662,I200933);
DFFARX1 I_11652 (I200902,I2859,I200478,I200467,);
DFFARX1 I_11653 (I200902,I2859,I200478,I200464,);
not I_11654 (I201022,I2866);
DFFARX1 I_11655 (I415159,I2859,I201022,I201048,);
DFFARX1 I_11656 (I201048,I2859,I201022,I201065,);
not I_11657 (I201014,I201065);
not I_11658 (I201087,I201048);
nand I_11659 (I201104,I415174,I415162);
and I_11660 (I201121,I201104,I415153);
DFFARX1 I_11661 (I201121,I2859,I201022,I201147,);
not I_11662 (I201155,I201147);
DFFARX1 I_11663 (I415165,I2859,I201022,I201181,);
and I_11664 (I201189,I201181,I415156);
nand I_11665 (I201206,I201181,I415156);
nand I_11666 (I200993,I201155,I201206);
DFFARX1 I_11667 (I415171,I2859,I201022,I201246,);
nor I_11668 (I201254,I201246,I201189);
DFFARX1 I_11669 (I201254,I2859,I201022,I200987,);
nor I_11670 (I201002,I201246,I201147);
nand I_11671 (I201299,I415180,I415168);
and I_11672 (I201316,I201299,I415177);
DFFARX1 I_11673 (I201316,I2859,I201022,I201342,);
nor I_11674 (I200990,I201342,I201246);
not I_11675 (I201364,I201342);
nor I_11676 (I201381,I201364,I201155);
nor I_11677 (I201398,I201087,I201381);
DFFARX1 I_11678 (I201398,I2859,I201022,I201005,);
nor I_11679 (I201429,I201364,I201246);
nor I_11680 (I201446,I415153,I415168);
nor I_11681 (I200996,I201446,I201429);
not I_11682 (I201477,I201446);
nand I_11683 (I200999,I201206,I201477);
DFFARX1 I_11684 (I201446,I2859,I201022,I201011,);
DFFARX1 I_11685 (I201446,I2859,I201022,I201008,);
not I_11686 (I201566,I2866);
DFFARX1 I_11687 (I263295,I2859,I201566,I201592,);
DFFARX1 I_11688 (I201592,I2859,I201566,I201609,);
not I_11689 (I201558,I201609);
not I_11690 (I201631,I201592);
nand I_11691 (I201648,I263292,I263313);
and I_11692 (I201665,I201648,I263316);
DFFARX1 I_11693 (I201665,I2859,I201566,I201691,);
not I_11694 (I201699,I201691);
DFFARX1 I_11695 (I263301,I2859,I201566,I201725,);
and I_11696 (I201733,I201725,I263304);
nand I_11697 (I201750,I201725,I263304);
nand I_11698 (I201537,I201699,I201750);
DFFARX1 I_11699 (I263307,I2859,I201566,I201790,);
nor I_11700 (I201798,I201790,I201733);
DFFARX1 I_11701 (I201798,I2859,I201566,I201531,);
nor I_11702 (I201546,I201790,I201691);
nand I_11703 (I201843,I263292,I263298);
and I_11704 (I201860,I201843,I263310);
DFFARX1 I_11705 (I201860,I2859,I201566,I201886,);
nor I_11706 (I201534,I201886,I201790);
not I_11707 (I201908,I201886);
nor I_11708 (I201925,I201908,I201699);
nor I_11709 (I201942,I201631,I201925);
DFFARX1 I_11710 (I201942,I2859,I201566,I201549,);
nor I_11711 (I201973,I201908,I201790);
nor I_11712 (I201990,I263295,I263298);
nor I_11713 (I201540,I201990,I201973);
not I_11714 (I202021,I201990);
nand I_11715 (I201543,I201750,I202021);
DFFARX1 I_11716 (I201990,I2859,I201566,I201555,);
DFFARX1 I_11717 (I201990,I2859,I201566,I201552,);
not I_11718 (I202110,I2866);
DFFARX1 I_11719 (I136136,I2859,I202110,I202136,);
DFFARX1 I_11720 (I202136,I2859,I202110,I202153,);
not I_11721 (I202102,I202153);
not I_11722 (I202175,I202136);
nand I_11723 (I202192,I136115,I136139);
and I_11724 (I202209,I202192,I136142);
DFFARX1 I_11725 (I202209,I2859,I202110,I202235,);
not I_11726 (I202243,I202235);
DFFARX1 I_11727 (I136124,I2859,I202110,I202269,);
and I_11728 (I202277,I202269,I136130);
nand I_11729 (I202294,I202269,I136130);
nand I_11730 (I202081,I202243,I202294);
DFFARX1 I_11731 (I136118,I2859,I202110,I202334,);
nor I_11732 (I202342,I202334,I202277);
DFFARX1 I_11733 (I202342,I2859,I202110,I202075,);
nor I_11734 (I202090,I202334,I202235);
nand I_11735 (I202387,I136127,I136115);
and I_11736 (I202404,I202387,I136121);
DFFARX1 I_11737 (I202404,I2859,I202110,I202430,);
nor I_11738 (I202078,I202430,I202334);
not I_11739 (I202452,I202430);
nor I_11740 (I202469,I202452,I202243);
nor I_11741 (I202486,I202175,I202469);
DFFARX1 I_11742 (I202486,I2859,I202110,I202093,);
nor I_11743 (I202517,I202452,I202334);
nor I_11744 (I202534,I136133,I136115);
nor I_11745 (I202084,I202534,I202517);
not I_11746 (I202565,I202534);
nand I_11747 (I202087,I202294,I202565);
DFFARX1 I_11748 (I202534,I2859,I202110,I202099,);
DFFARX1 I_11749 (I202534,I2859,I202110,I202096,);
not I_11750 (I202654,I2866);
DFFARX1 I_11751 (I29429,I2859,I202654,I202680,);
DFFARX1 I_11752 (I202680,I2859,I202654,I202697,);
not I_11753 (I202646,I202697);
not I_11754 (I202719,I202680);
nand I_11755 (I202736,I29444,I29423);
and I_11756 (I202753,I202736,I29426);
DFFARX1 I_11757 (I202753,I2859,I202654,I202779,);
not I_11758 (I202787,I202779);
DFFARX1 I_11759 (I29432,I2859,I202654,I202813,);
and I_11760 (I202821,I202813,I29426);
nand I_11761 (I202838,I202813,I29426);
nand I_11762 (I202625,I202787,I202838);
DFFARX1 I_11763 (I29441,I2859,I202654,I202878,);
nor I_11764 (I202886,I202878,I202821);
DFFARX1 I_11765 (I202886,I2859,I202654,I202619,);
nor I_11766 (I202634,I202878,I202779);
nand I_11767 (I202931,I29423,I29438);
and I_11768 (I202948,I202931,I29435);
DFFARX1 I_11769 (I202948,I2859,I202654,I202974,);
nor I_11770 (I202622,I202974,I202878);
not I_11771 (I202996,I202974);
nor I_11772 (I203013,I202996,I202787);
nor I_11773 (I203030,I202719,I203013);
DFFARX1 I_11774 (I203030,I2859,I202654,I202637,);
nor I_11775 (I203061,I202996,I202878);
nor I_11776 (I203078,I29447,I29438);
nor I_11777 (I202628,I203078,I203061);
not I_11778 (I203109,I203078);
nand I_11779 (I202631,I202838,I203109);
DFFARX1 I_11780 (I203078,I2859,I202654,I202643,);
DFFARX1 I_11781 (I203078,I2859,I202654,I202640,);
not I_11782 (I203198,I2866);
DFFARX1 I_11783 (I260983,I2859,I203198,I203224,);
DFFARX1 I_11784 (I203224,I2859,I203198,I203241,);
not I_11785 (I203190,I203241);
not I_11786 (I203263,I203224);
nand I_11787 (I203280,I260980,I261001);
and I_11788 (I203297,I203280,I261004);
DFFARX1 I_11789 (I203297,I2859,I203198,I203323,);
not I_11790 (I203331,I203323);
DFFARX1 I_11791 (I260989,I2859,I203198,I203357,);
and I_11792 (I203365,I203357,I260992);
nand I_11793 (I203382,I203357,I260992);
nand I_11794 (I203169,I203331,I203382);
DFFARX1 I_11795 (I260995,I2859,I203198,I203422,);
nor I_11796 (I203430,I203422,I203365);
DFFARX1 I_11797 (I203430,I2859,I203198,I203163,);
nor I_11798 (I203178,I203422,I203323);
nand I_11799 (I203475,I260980,I260986);
and I_11800 (I203492,I203475,I260998);
DFFARX1 I_11801 (I203492,I2859,I203198,I203518,);
nor I_11802 (I203166,I203518,I203422);
not I_11803 (I203540,I203518);
nor I_11804 (I203557,I203540,I203331);
nor I_11805 (I203574,I203263,I203557);
DFFARX1 I_11806 (I203574,I2859,I203198,I203181,);
nor I_11807 (I203605,I203540,I203422);
nor I_11808 (I203622,I260983,I260986);
nor I_11809 (I203172,I203622,I203605);
not I_11810 (I203653,I203622);
nand I_11811 (I203175,I203382,I203653);
DFFARX1 I_11812 (I203622,I2859,I203198,I203187,);
DFFARX1 I_11813 (I203622,I2859,I203198,I203184,);
not I_11814 (I203742,I2866);
DFFARX1 I_11815 (I464507,I2859,I203742,I203768,);
DFFARX1 I_11816 (I203768,I2859,I203742,I203785,);
not I_11817 (I203734,I203785);
not I_11818 (I203807,I203768);
nand I_11819 (I203824,I464519,I464507);
and I_11820 (I203841,I203824,I464510);
DFFARX1 I_11821 (I203841,I2859,I203742,I203867,);
not I_11822 (I203875,I203867);
DFFARX1 I_11823 (I464528,I2859,I203742,I203901,);
and I_11824 (I203909,I203901,I464504);
nand I_11825 (I203926,I203901,I464504);
nand I_11826 (I203713,I203875,I203926);
DFFARX1 I_11827 (I464522,I2859,I203742,I203966,);
nor I_11828 (I203974,I203966,I203909);
DFFARX1 I_11829 (I203974,I2859,I203742,I203707,);
nor I_11830 (I203722,I203966,I203867);
nand I_11831 (I204019,I464516,I464513);
and I_11832 (I204036,I204019,I464525);
DFFARX1 I_11833 (I204036,I2859,I203742,I204062,);
nor I_11834 (I203710,I204062,I203966);
not I_11835 (I204084,I204062);
nor I_11836 (I204101,I204084,I203875);
nor I_11837 (I204118,I203807,I204101);
DFFARX1 I_11838 (I204118,I2859,I203742,I203725,);
nor I_11839 (I204149,I204084,I203966);
nor I_11840 (I204166,I464504,I464513);
nor I_11841 (I203716,I204166,I204149);
not I_11842 (I204197,I204166);
nand I_11843 (I203719,I203926,I204197);
DFFARX1 I_11844 (I204166,I2859,I203742,I203731,);
DFFARX1 I_11845 (I204166,I2859,I203742,I203728,);
not I_11846 (I204286,I2866);
DFFARX1 I_11847 (I26267,I2859,I204286,I204312,);
DFFARX1 I_11848 (I204312,I2859,I204286,I204329,);
not I_11849 (I204278,I204329);
not I_11850 (I204351,I204312);
nand I_11851 (I204368,I26282,I26261);
and I_11852 (I204385,I204368,I26264);
DFFARX1 I_11853 (I204385,I2859,I204286,I204411,);
not I_11854 (I204419,I204411);
DFFARX1 I_11855 (I26270,I2859,I204286,I204445,);
and I_11856 (I204453,I204445,I26264);
nand I_11857 (I204470,I204445,I26264);
nand I_11858 (I204257,I204419,I204470);
DFFARX1 I_11859 (I26279,I2859,I204286,I204510,);
nor I_11860 (I204518,I204510,I204453);
DFFARX1 I_11861 (I204518,I2859,I204286,I204251,);
nor I_11862 (I204266,I204510,I204411);
nand I_11863 (I204563,I26261,I26276);
and I_11864 (I204580,I204563,I26273);
DFFARX1 I_11865 (I204580,I2859,I204286,I204606,);
nor I_11866 (I204254,I204606,I204510);
not I_11867 (I204628,I204606);
nor I_11868 (I204645,I204628,I204419);
nor I_11869 (I204662,I204351,I204645);
DFFARX1 I_11870 (I204662,I2859,I204286,I204269,);
nor I_11871 (I204693,I204628,I204510);
nor I_11872 (I204710,I26285,I26276);
nor I_11873 (I204260,I204710,I204693);
not I_11874 (I204741,I204710);
nand I_11875 (I204263,I204470,I204741);
DFFARX1 I_11876 (I204710,I2859,I204286,I204275,);
DFFARX1 I_11877 (I204710,I2859,I204286,I204272,);
not I_11878 (I204830,I2866);
DFFARX1 I_11879 (I495719,I2859,I204830,I204856,);
DFFARX1 I_11880 (I204856,I2859,I204830,I204873,);
not I_11881 (I204822,I204873);
not I_11882 (I204895,I204856);
nand I_11883 (I204912,I495731,I495719);
and I_11884 (I204929,I204912,I495722);
DFFARX1 I_11885 (I204929,I2859,I204830,I204955,);
not I_11886 (I204963,I204955);
DFFARX1 I_11887 (I495740,I2859,I204830,I204989,);
and I_11888 (I204997,I204989,I495716);
nand I_11889 (I205014,I204989,I495716);
nand I_11890 (I204801,I204963,I205014);
DFFARX1 I_11891 (I495734,I2859,I204830,I205054,);
nor I_11892 (I205062,I205054,I204997);
DFFARX1 I_11893 (I205062,I2859,I204830,I204795,);
nor I_11894 (I204810,I205054,I204955);
nand I_11895 (I205107,I495728,I495725);
and I_11896 (I205124,I205107,I495737);
DFFARX1 I_11897 (I205124,I2859,I204830,I205150,);
nor I_11898 (I204798,I205150,I205054);
not I_11899 (I205172,I205150);
nor I_11900 (I205189,I205172,I204963);
nor I_11901 (I205206,I204895,I205189);
DFFARX1 I_11902 (I205206,I2859,I204830,I204813,);
nor I_11903 (I205237,I205172,I205054);
nor I_11904 (I205254,I495716,I495725);
nor I_11905 (I204804,I205254,I205237);
not I_11906 (I205285,I205254);
nand I_11907 (I204807,I205014,I205285);
DFFARX1 I_11908 (I205254,I2859,I204830,I204819,);
DFFARX1 I_11909 (I205254,I2859,I204830,I204816,);
not I_11910 (I205374,I2866);
DFFARX1 I_11911 (I444954,I2859,I205374,I205400,);
DFFARX1 I_11912 (I205400,I2859,I205374,I205417,);
not I_11913 (I205366,I205417);
not I_11914 (I205439,I205400);
nand I_11915 (I205456,I444954,I444972);
and I_11916 (I205473,I205456,I444966);
DFFARX1 I_11917 (I205473,I2859,I205374,I205499,);
not I_11918 (I205507,I205499);
DFFARX1 I_11919 (I444960,I2859,I205374,I205533,);
and I_11920 (I205541,I205533,I444969);
nand I_11921 (I205558,I205533,I444969);
nand I_11922 (I205345,I205507,I205558);
DFFARX1 I_11923 (I444957,I2859,I205374,I205598,);
nor I_11924 (I205606,I205598,I205541);
DFFARX1 I_11925 (I205606,I2859,I205374,I205339,);
nor I_11926 (I205354,I205598,I205499);
nand I_11927 (I205651,I444957,I444975);
and I_11928 (I205668,I205651,I444960);
DFFARX1 I_11929 (I205668,I2859,I205374,I205694,);
nor I_11930 (I205342,I205694,I205598);
not I_11931 (I205716,I205694);
nor I_11932 (I205733,I205716,I205507);
nor I_11933 (I205750,I205439,I205733);
DFFARX1 I_11934 (I205750,I2859,I205374,I205357,);
nor I_11935 (I205781,I205716,I205598);
nor I_11936 (I205798,I444963,I444975);
nor I_11937 (I205348,I205798,I205781);
not I_11938 (I205829,I205798);
nand I_11939 (I205351,I205558,I205829);
DFFARX1 I_11940 (I205798,I2859,I205374,I205363,);
DFFARX1 I_11941 (I205798,I2859,I205374,I205360,);
not I_11942 (I205918,I2866);
DFFARX1 I_11943 (I432051,I2859,I205918,I205944,);
DFFARX1 I_11944 (I205944,I2859,I205918,I205961,);
not I_11945 (I205910,I205961);
not I_11946 (I205983,I205944);
nand I_11947 (I206000,I432051,I432069);
and I_11948 (I206017,I206000,I432063);
DFFARX1 I_11949 (I206017,I2859,I205918,I206043,);
not I_11950 (I206051,I206043);
DFFARX1 I_11951 (I432057,I2859,I205918,I206077,);
and I_11952 (I206085,I206077,I432066);
nand I_11953 (I206102,I206077,I432066);
nand I_11954 (I205889,I206051,I206102);
DFFARX1 I_11955 (I432054,I2859,I205918,I206142,);
nor I_11956 (I206150,I206142,I206085);
DFFARX1 I_11957 (I206150,I2859,I205918,I205883,);
nor I_11958 (I205898,I206142,I206043);
nand I_11959 (I206195,I432054,I432072);
and I_11960 (I206212,I206195,I432057);
DFFARX1 I_11961 (I206212,I2859,I205918,I206238,);
nor I_11962 (I205886,I206238,I206142);
not I_11963 (I206260,I206238);
nor I_11964 (I206277,I206260,I206051);
nor I_11965 (I206294,I205983,I206277);
DFFARX1 I_11966 (I206294,I2859,I205918,I205901,);
nor I_11967 (I206325,I206260,I206142);
nor I_11968 (I206342,I432060,I432072);
nor I_11969 (I205892,I206342,I206325);
not I_11970 (I206373,I206342);
nand I_11971 (I205895,I206102,I206373);
DFFARX1 I_11972 (I206342,I2859,I205918,I205907,);
DFFARX1 I_11973 (I206342,I2859,I205918,I205904,);
not I_11974 (I206462,I2866);
DFFARX1 I_11975 (I216681,I2859,I206462,I206488,);
DFFARX1 I_11976 (I206488,I2859,I206462,I206505,);
not I_11977 (I206454,I206505);
not I_11978 (I206527,I206488);
nand I_11979 (I206544,I216684,I216702);
and I_11980 (I206561,I206544,I216690);
DFFARX1 I_11981 (I206561,I2859,I206462,I206587,);
not I_11982 (I206595,I206587);
DFFARX1 I_11983 (I216681,I2859,I206462,I206621,);
and I_11984 (I206629,I206621,I216699);
nand I_11985 (I206646,I206621,I216699);
nand I_11986 (I206433,I206595,I206646);
DFFARX1 I_11987 (I216693,I2859,I206462,I206686,);
nor I_11988 (I206694,I206686,I206629);
DFFARX1 I_11989 (I206694,I2859,I206462,I206427,);
nor I_11990 (I206442,I206686,I206587);
nand I_11991 (I206739,I216696,I216678);
and I_11992 (I206756,I206739,I216687);
DFFARX1 I_11993 (I206756,I2859,I206462,I206782,);
nor I_11994 (I206430,I206782,I206686);
not I_11995 (I206804,I206782);
nor I_11996 (I206821,I206804,I206595);
nor I_11997 (I206838,I206527,I206821);
DFFARX1 I_11998 (I206838,I2859,I206462,I206445,);
nor I_11999 (I206869,I206804,I206686);
nor I_12000 (I206886,I216678,I216678);
nor I_12001 (I206436,I206886,I206869);
not I_12002 (I206917,I206886);
nand I_12003 (I206439,I206646,I206917);
DFFARX1 I_12004 (I206886,I2859,I206462,I206451,);
DFFARX1 I_12005 (I206886,I2859,I206462,I206448,);
not I_12006 (I207006,I2866);
DFFARX1 I_12007 (I5193,I2859,I207006,I207032,);
DFFARX1 I_12008 (I207032,I2859,I207006,I207049,);
not I_12009 (I206998,I207049);
not I_12010 (I207071,I207032);
nand I_12011 (I207088,I5181,I5196);
and I_12012 (I207105,I207088,I5184);
DFFARX1 I_12013 (I207105,I2859,I207006,I207131,);
not I_12014 (I207139,I207131);
DFFARX1 I_12015 (I5205,I2859,I207006,I207165,);
and I_12016 (I207173,I207165,I5199);
nand I_12017 (I207190,I207165,I5199);
nand I_12018 (I206977,I207139,I207190);
DFFARX1 I_12019 (I5202,I2859,I207006,I207230,);
nor I_12020 (I207238,I207230,I207173);
DFFARX1 I_12021 (I207238,I2859,I207006,I206971,);
nor I_12022 (I206986,I207230,I207131);
nand I_12023 (I207283,I5181,I5184);
and I_12024 (I207300,I207283,I5187);
DFFARX1 I_12025 (I207300,I2859,I207006,I207326,);
nor I_12026 (I206974,I207326,I207230);
not I_12027 (I207348,I207326);
nor I_12028 (I207365,I207348,I207139);
nor I_12029 (I207382,I207071,I207365);
DFFARX1 I_12030 (I207382,I2859,I207006,I206989,);
nor I_12031 (I207413,I207348,I207230);
nor I_12032 (I207430,I5190,I5184);
nor I_12033 (I206980,I207430,I207413);
not I_12034 (I207461,I207430);
nand I_12035 (I206983,I207190,I207461);
DFFARX1 I_12036 (I207430,I2859,I207006,I206995,);
DFFARX1 I_12037 (I207430,I2859,I207006,I206992,);
not I_12038 (I207550,I2866);
DFFARX1 I_12039 (I156689,I2859,I207550,I207576,);
DFFARX1 I_12040 (I207576,I2859,I207550,I207593,);
not I_12041 (I207542,I207593);
not I_12042 (I207615,I207576);
nand I_12043 (I207632,I156668,I156692);
and I_12044 (I207649,I207632,I156695);
DFFARX1 I_12045 (I207649,I2859,I207550,I207675,);
not I_12046 (I207683,I207675);
DFFARX1 I_12047 (I156677,I2859,I207550,I207709,);
and I_12048 (I207717,I207709,I156683);
nand I_12049 (I207734,I207709,I156683);
nand I_12050 (I207521,I207683,I207734);
DFFARX1 I_12051 (I156671,I2859,I207550,I207774,);
nor I_12052 (I207782,I207774,I207717);
DFFARX1 I_12053 (I207782,I2859,I207550,I207515,);
nor I_12054 (I207530,I207774,I207675);
nand I_12055 (I207827,I156680,I156668);
and I_12056 (I207844,I207827,I156674);
DFFARX1 I_12057 (I207844,I2859,I207550,I207870,);
nor I_12058 (I207518,I207870,I207774);
not I_12059 (I207892,I207870);
nor I_12060 (I207909,I207892,I207683);
nor I_12061 (I207926,I207615,I207909);
DFFARX1 I_12062 (I207926,I2859,I207550,I207533,);
nor I_12063 (I207957,I207892,I207774);
nor I_12064 (I207974,I156686,I156668);
nor I_12065 (I207524,I207974,I207957);
not I_12066 (I208005,I207974);
nand I_12067 (I207527,I207734,I208005);
DFFARX1 I_12068 (I207974,I2859,I207550,I207539,);
DFFARX1 I_12069 (I207974,I2859,I207550,I207536,);
not I_12070 (I208094,I2866);
DFFARX1 I_12071 (I262717,I2859,I208094,I208120,);
DFFARX1 I_12072 (I208120,I2859,I208094,I208137,);
not I_12073 (I208086,I208137);
not I_12074 (I208159,I208120);
nand I_12075 (I208176,I262714,I262735);
and I_12076 (I208193,I208176,I262738);
DFFARX1 I_12077 (I208193,I2859,I208094,I208219,);
not I_12078 (I208227,I208219);
DFFARX1 I_12079 (I262723,I2859,I208094,I208253,);
and I_12080 (I208261,I208253,I262726);
nand I_12081 (I208278,I208253,I262726);
nand I_12082 (I208065,I208227,I208278);
DFFARX1 I_12083 (I262729,I2859,I208094,I208318,);
nor I_12084 (I208326,I208318,I208261);
DFFARX1 I_12085 (I208326,I2859,I208094,I208059,);
nor I_12086 (I208074,I208318,I208219);
nand I_12087 (I208371,I262714,I262720);
and I_12088 (I208388,I208371,I262732);
DFFARX1 I_12089 (I208388,I2859,I208094,I208414,);
nor I_12090 (I208062,I208414,I208318);
not I_12091 (I208436,I208414);
nor I_12092 (I208453,I208436,I208227);
nor I_12093 (I208470,I208159,I208453);
DFFARX1 I_12094 (I208470,I2859,I208094,I208077,);
nor I_12095 (I208501,I208436,I208318);
nor I_12096 (I208518,I262717,I262720);
nor I_12097 (I208068,I208518,I208501);
not I_12098 (I208549,I208518);
nand I_12099 (I208071,I208278,I208549);
DFFARX1 I_12100 (I208518,I2859,I208094,I208083,);
DFFARX1 I_12101 (I208518,I2859,I208094,I208080,);
not I_12102 (I208638,I2866);
DFFARX1 I_12103 (I248845,I2859,I208638,I208664,);
DFFARX1 I_12104 (I208664,I2859,I208638,I208681,);
not I_12105 (I208630,I208681);
not I_12106 (I208703,I208664);
nand I_12107 (I208720,I248842,I248863);
and I_12108 (I208737,I208720,I248866);
DFFARX1 I_12109 (I208737,I2859,I208638,I208763,);
not I_12110 (I208771,I208763);
DFFARX1 I_12111 (I248851,I2859,I208638,I208797,);
and I_12112 (I208805,I208797,I248854);
nand I_12113 (I208822,I208797,I248854);
nand I_12114 (I208609,I208771,I208822);
DFFARX1 I_12115 (I248857,I2859,I208638,I208862,);
nor I_12116 (I208870,I208862,I208805);
DFFARX1 I_12117 (I208870,I2859,I208638,I208603,);
nor I_12118 (I208618,I208862,I208763);
nand I_12119 (I208915,I248842,I248848);
and I_12120 (I208932,I208915,I248860);
DFFARX1 I_12121 (I208932,I2859,I208638,I208958,);
nor I_12122 (I208606,I208958,I208862);
not I_12123 (I208980,I208958);
nor I_12124 (I208997,I208980,I208771);
nor I_12125 (I209014,I208703,I208997);
DFFARX1 I_12126 (I209014,I2859,I208638,I208621,);
nor I_12127 (I209045,I208980,I208862);
nor I_12128 (I209062,I248845,I248848);
nor I_12129 (I208612,I209062,I209045);
not I_12130 (I209093,I209062);
nand I_12131 (I208615,I208822,I209093);
DFFARX1 I_12132 (I209062,I2859,I208638,I208627,);
DFFARX1 I_12133 (I209062,I2859,I208638,I208624,);
not I_12134 (I209182,I2866);
DFFARX1 I_12135 (I511325,I2859,I209182,I209208,);
DFFARX1 I_12136 (I209208,I2859,I209182,I209225,);
not I_12137 (I209174,I209225);
not I_12138 (I209247,I209208);
nand I_12139 (I209264,I511337,I511340);
and I_12140 (I209281,I209264,I511343);
DFFARX1 I_12141 (I209281,I2859,I209182,I209307,);
not I_12142 (I209315,I209307);
DFFARX1 I_12143 (I511328,I2859,I209182,I209341,);
and I_12144 (I209349,I209341,I511334);
nand I_12145 (I209366,I209341,I511334);
nand I_12146 (I209153,I209315,I209366);
DFFARX1 I_12147 (I511322,I2859,I209182,I209406,);
nor I_12148 (I209414,I209406,I209349);
DFFARX1 I_12149 (I209414,I2859,I209182,I209147,);
nor I_12150 (I209162,I209406,I209307);
nand I_12151 (I209459,I511325,I511346);
and I_12152 (I209476,I209459,I511331);
DFFARX1 I_12153 (I209476,I2859,I209182,I209502,);
nor I_12154 (I209150,I209502,I209406);
not I_12155 (I209524,I209502);
nor I_12156 (I209541,I209524,I209315);
nor I_12157 (I209558,I209247,I209541);
DFFARX1 I_12158 (I209558,I2859,I209182,I209165,);
nor I_12159 (I209589,I209524,I209406);
nor I_12160 (I209606,I511322,I511346);
nor I_12161 (I209156,I209606,I209589);
not I_12162 (I209637,I209606);
nand I_12163 (I209159,I209366,I209637);
DFFARX1 I_12164 (I209606,I2859,I209182,I209171,);
DFFARX1 I_12165 (I209606,I2859,I209182,I209168,);
not I_12166 (I209726,I2866);
DFFARX1 I_12167 (I354798,I2859,I209726,I209752,);
DFFARX1 I_12168 (I209752,I2859,I209726,I209769,);
not I_12169 (I209718,I209769);
not I_12170 (I209791,I209752);
nand I_12171 (I209808,I354792,I354789);
and I_12172 (I209825,I209808,I354804);
DFFARX1 I_12173 (I209825,I2859,I209726,I209851,);
not I_12174 (I209859,I209851);
DFFARX1 I_12175 (I354792,I2859,I209726,I209885,);
and I_12176 (I209893,I209885,I354786);
nand I_12177 (I209910,I209885,I354786);
nand I_12178 (I209697,I209859,I209910);
DFFARX1 I_12179 (I354786,I2859,I209726,I209950,);
nor I_12180 (I209958,I209950,I209893);
DFFARX1 I_12181 (I209958,I2859,I209726,I209691,);
nor I_12182 (I209706,I209950,I209851);
nand I_12183 (I210003,I354801,I354795);
and I_12184 (I210020,I210003,I354789);
DFFARX1 I_12185 (I210020,I2859,I209726,I210046,);
nor I_12186 (I209694,I210046,I209950);
not I_12187 (I210068,I210046);
nor I_12188 (I210085,I210068,I209859);
nor I_12189 (I210102,I209791,I210085);
DFFARX1 I_12190 (I210102,I2859,I209726,I209709,);
nor I_12191 (I210133,I210068,I209950);
nor I_12192 (I210150,I354807,I354795);
nor I_12193 (I209700,I210150,I210133);
not I_12194 (I210181,I210150);
nand I_12195 (I209703,I209910,I210181);
DFFARX1 I_12196 (I210150,I2859,I209726,I209715,);
DFFARX1 I_12197 (I210150,I2859,I209726,I209712,);
not I_12198 (I210270,I2866);
DFFARX1 I_12199 (I387381,I2859,I210270,I210296,);
DFFARX1 I_12200 (I210296,I2859,I210270,I210313,);
not I_12201 (I210262,I210313);
not I_12202 (I210335,I210296);
nand I_12203 (I210352,I387396,I387384);
and I_12204 (I210369,I210352,I387375);
DFFARX1 I_12205 (I210369,I2859,I210270,I210395,);
not I_12206 (I210403,I210395);
DFFARX1 I_12207 (I387387,I2859,I210270,I210429,);
and I_12208 (I210437,I210429,I387378);
nand I_12209 (I210454,I210429,I387378);
nand I_12210 (I210241,I210403,I210454);
DFFARX1 I_12211 (I387393,I2859,I210270,I210494,);
nor I_12212 (I210502,I210494,I210437);
DFFARX1 I_12213 (I210502,I2859,I210270,I210235,);
nor I_12214 (I210250,I210494,I210395);
nand I_12215 (I210547,I387402,I387390);
and I_12216 (I210564,I210547,I387399);
DFFARX1 I_12217 (I210564,I2859,I210270,I210590,);
nor I_12218 (I210238,I210590,I210494);
not I_12219 (I210612,I210590);
nor I_12220 (I210629,I210612,I210403);
nor I_12221 (I210646,I210335,I210629);
DFFARX1 I_12222 (I210646,I2859,I210270,I210253,);
nor I_12223 (I210677,I210612,I210494);
nor I_12224 (I210694,I387375,I387390);
nor I_12225 (I210244,I210694,I210677);
not I_12226 (I210725,I210694);
nand I_12227 (I210247,I210454,I210725);
DFFARX1 I_12228 (I210694,I2859,I210270,I210259,);
DFFARX1 I_12229 (I210694,I2859,I210270,I210256,);
not I_12230 (I210814,I2866);
DFFARX1 I_12231 (I13098,I2859,I210814,I210840,);
DFFARX1 I_12232 (I210840,I2859,I210814,I210857,);
not I_12233 (I210806,I210857);
not I_12234 (I210879,I210840);
nand I_12235 (I210896,I13086,I13101);
and I_12236 (I210913,I210896,I13089);
DFFARX1 I_12237 (I210913,I2859,I210814,I210939,);
not I_12238 (I210947,I210939);
DFFARX1 I_12239 (I13110,I2859,I210814,I210973,);
and I_12240 (I210981,I210973,I13104);
nand I_12241 (I210998,I210973,I13104);
nand I_12242 (I210785,I210947,I210998);
DFFARX1 I_12243 (I13107,I2859,I210814,I211038,);
nor I_12244 (I211046,I211038,I210981);
DFFARX1 I_12245 (I211046,I2859,I210814,I210779,);
nor I_12246 (I210794,I211038,I210939);
nand I_12247 (I211091,I13086,I13089);
and I_12248 (I211108,I211091,I13092);
DFFARX1 I_12249 (I211108,I2859,I210814,I211134,);
nor I_12250 (I210782,I211134,I211038);
not I_12251 (I211156,I211134);
nor I_12252 (I211173,I211156,I210947);
nor I_12253 (I211190,I210879,I211173);
DFFARX1 I_12254 (I211190,I2859,I210814,I210797,);
nor I_12255 (I211221,I211156,I211038);
nor I_12256 (I211238,I13095,I13089);
nor I_12257 (I210788,I211238,I211221);
not I_12258 (I211269,I211238);
nand I_12259 (I210791,I210998,I211269);
DFFARX1 I_12260 (I211238,I2859,I210814,I210803,);
DFFARX1 I_12261 (I211238,I2859,I210814,I210800,);
not I_12262 (I211355,I2866);
DFFARX1 I_12263 (I317055,I2859,I211355,I211381,);
DFFARX1 I_12264 (I211381,I2859,I211355,I211398,);
not I_12265 (I211347,I211398);
DFFARX1 I_12266 (I317049,I2859,I211355,I211429,);
not I_12267 (I211437,I317046);
nor I_12268 (I211454,I211381,I211437);
not I_12269 (I211471,I317058);
not I_12270 (I211488,I317061);
nand I_12271 (I211505,I211488,I317058);
nor I_12272 (I211522,I211437,I211505);
nor I_12273 (I211539,I211429,I211522);
DFFARX1 I_12274 (I211488,I2859,I211355,I211344,);
nor I_12275 (I211570,I317061,I317070);
nand I_12276 (I211587,I211570,I317064);
nor I_12277 (I211604,I211587,I211471);
nand I_12278 (I211329,I211604,I317046);
DFFARX1 I_12279 (I211587,I2859,I211355,I211341,);
nand I_12280 (I211649,I211471,I317061);
nor I_12281 (I211666,I211471,I317061);
nand I_12282 (I211335,I211454,I211666);
not I_12283 (I211697,I317052);
nor I_12284 (I211714,I211697,I211649);
DFFARX1 I_12285 (I211714,I2859,I211355,I211323,);
nor I_12286 (I211745,I211697,I317067);
and I_12287 (I211762,I211745,I317046);
or I_12288 (I211779,I211762,I317049);
DFFARX1 I_12289 (I211779,I2859,I211355,I211805,);
nor I_12290 (I211813,I211805,I211429);
nor I_12291 (I211332,I211381,I211813);
not I_12292 (I211844,I211805);
nor I_12293 (I211861,I211844,I211539);
DFFARX1 I_12294 (I211861,I2859,I211355,I211338,);
nand I_12295 (I211892,I211844,I211471);
nor I_12296 (I211326,I211697,I211892);
not I_12297 (I211950,I2866);
DFFARX1 I_12298 (I67333,I2859,I211950,I211976,);
DFFARX1 I_12299 (I211976,I2859,I211950,I211993,);
not I_12300 (I211942,I211993);
DFFARX1 I_12301 (I67357,I2859,I211950,I212024,);
not I_12302 (I212032,I67351);
nor I_12303 (I212049,I211976,I212032);
not I_12304 (I212066,I67345);
not I_12305 (I212083,I67342);
nand I_12306 (I212100,I212083,I67345);
nor I_12307 (I212117,I212032,I212100);
nor I_12308 (I212134,I212024,I212117);
DFFARX1 I_12309 (I212083,I2859,I211950,I211939,);
nor I_12310 (I212165,I67342,I67336);
nand I_12311 (I212182,I212165,I67354);
nor I_12312 (I212199,I212182,I212066);
nand I_12313 (I211924,I212199,I67351);
DFFARX1 I_12314 (I212182,I2859,I211950,I211936,);
nand I_12315 (I212244,I212066,I67342);
nor I_12316 (I212261,I212066,I67342);
nand I_12317 (I211930,I212049,I212261);
not I_12318 (I212292,I67348);
nor I_12319 (I212309,I212292,I212244);
DFFARX1 I_12320 (I212309,I2859,I211950,I211918,);
nor I_12321 (I212340,I212292,I67333);
and I_12322 (I212357,I212340,I67339);
or I_12323 (I212374,I212357,I67336);
DFFARX1 I_12324 (I212374,I2859,I211950,I212400,);
nor I_12325 (I212408,I212400,I212024);
nor I_12326 (I211927,I211976,I212408);
not I_12327 (I212439,I212400);
nor I_12328 (I212456,I212439,I212134);
DFFARX1 I_12329 (I212456,I2859,I211950,I211933,);
nand I_12330 (I212487,I212439,I212066);
nor I_12331 (I211921,I212292,I212487);
not I_12332 (I212545,I2866);
DFFARX1 I_12333 (I247111,I2859,I212545,I212571,);
DFFARX1 I_12334 (I212571,I2859,I212545,I212588,);
not I_12335 (I212537,I212588);
DFFARX1 I_12336 (I247123,I2859,I212545,I212619,);
not I_12337 (I212627,I247108);
nor I_12338 (I212644,I212571,I212627);
not I_12339 (I212661,I247126);
not I_12340 (I212678,I247117);
nand I_12341 (I212695,I212678,I247126);
nor I_12342 (I212712,I212627,I212695);
nor I_12343 (I212729,I212619,I212712);
DFFARX1 I_12344 (I212678,I2859,I212545,I212534,);
nor I_12345 (I212760,I247117,I247129);
nand I_12346 (I212777,I212760,I247132);
nor I_12347 (I212794,I212777,I212661);
nand I_12348 (I212519,I212794,I247108);
DFFARX1 I_12349 (I212777,I2859,I212545,I212531,);
nand I_12350 (I212839,I212661,I247117);
nor I_12351 (I212856,I212661,I247117);
nand I_12352 (I212525,I212644,I212856);
not I_12353 (I212887,I247108);
nor I_12354 (I212904,I212887,I212839);
DFFARX1 I_12355 (I212904,I2859,I212545,I212513,);
nor I_12356 (I212935,I212887,I247120);
and I_12357 (I212952,I212935,I247114);
or I_12358 (I212969,I212952,I247111);
DFFARX1 I_12359 (I212969,I2859,I212545,I212995,);
nor I_12360 (I213003,I212995,I212619);
nor I_12361 (I212522,I212571,I213003);
not I_12362 (I213034,I212995);
nor I_12363 (I213051,I213034,I212729);
DFFARX1 I_12364 (I213051,I2859,I212545,I212528,);
nand I_12365 (I213082,I213034,I212661);
nor I_12366 (I212516,I212887,I213082);
not I_12367 (I213140,I2866);
DFFARX1 I_12368 (I76853,I2859,I213140,I213166,);
DFFARX1 I_12369 (I213166,I2859,I213140,I213183,);
not I_12370 (I213132,I213183);
DFFARX1 I_12371 (I76877,I2859,I213140,I213214,);
not I_12372 (I213222,I76871);
nor I_12373 (I213239,I213166,I213222);
not I_12374 (I213256,I76865);
not I_12375 (I213273,I76862);
nand I_12376 (I213290,I213273,I76865);
nor I_12377 (I213307,I213222,I213290);
nor I_12378 (I213324,I213214,I213307);
DFFARX1 I_12379 (I213273,I2859,I213140,I213129,);
nor I_12380 (I213355,I76862,I76856);
nand I_12381 (I213372,I213355,I76874);
nor I_12382 (I213389,I213372,I213256);
nand I_12383 (I213114,I213389,I76871);
DFFARX1 I_12384 (I213372,I2859,I213140,I213126,);
nand I_12385 (I213434,I213256,I76862);
nor I_12386 (I213451,I213256,I76862);
nand I_12387 (I213120,I213239,I213451);
not I_12388 (I213482,I76868);
nor I_12389 (I213499,I213482,I213434);
DFFARX1 I_12390 (I213499,I2859,I213140,I213108,);
nor I_12391 (I213530,I213482,I76853);
and I_12392 (I213547,I213530,I76859);
or I_12393 (I213564,I213547,I76856);
DFFARX1 I_12394 (I213564,I2859,I213140,I213590,);
nor I_12395 (I213598,I213590,I213214);
nor I_12396 (I213117,I213166,I213598);
not I_12397 (I213629,I213590);
nor I_12398 (I213646,I213629,I213324);
DFFARX1 I_12399 (I213646,I2859,I213140,I213123,);
nand I_12400 (I213677,I213629,I213256);
nor I_12401 (I213111,I213482,I213677);
not I_12402 (I213735,I2866);
DFFARX1 I_12403 (I376408,I2859,I213735,I213761,);
DFFARX1 I_12404 (I213761,I2859,I213735,I213778,);
not I_12405 (I213727,I213778);
DFFARX1 I_12406 (I376396,I2859,I213735,I213809,);
not I_12407 (I213817,I376393);
nor I_12408 (I213834,I213761,I213817);
not I_12409 (I213851,I376405);
not I_12410 (I213868,I376402);
nand I_12411 (I213885,I213868,I376405);
nor I_12412 (I213902,I213817,I213885);
nor I_12413 (I213919,I213809,I213902);
DFFARX1 I_12414 (I213868,I2859,I213735,I213724,);
nor I_12415 (I213950,I376402,I376411);
nand I_12416 (I213967,I213950,I376414);
nor I_12417 (I213984,I213967,I213851);
nand I_12418 (I213709,I213984,I376393);
DFFARX1 I_12419 (I213967,I2859,I213735,I213721,);
nand I_12420 (I214029,I213851,I376402);
nor I_12421 (I214046,I213851,I376402);
nand I_12422 (I213715,I213834,I214046);
not I_12423 (I214077,I376417);
nor I_12424 (I214094,I214077,I214029);
DFFARX1 I_12425 (I214094,I2859,I213735,I213703,);
nor I_12426 (I214125,I214077,I376420);
and I_12427 (I214142,I214125,I376399);
or I_12428 (I214159,I214142,I376393);
DFFARX1 I_12429 (I214159,I2859,I213735,I214185,);
nor I_12430 (I214193,I214185,I213809);
nor I_12431 (I213712,I213761,I214193);
not I_12432 (I214224,I214185);
nor I_12433 (I214241,I214224,I213919);
DFFARX1 I_12434 (I214241,I2859,I213735,I213718,);
nand I_12435 (I214272,I214224,I213851);
nor I_12436 (I213706,I214077,I214272);
not I_12437 (I214330,I2866);
DFFARX1 I_12438 (I92918,I2859,I214330,I214356,);
DFFARX1 I_12439 (I214356,I2859,I214330,I214373,);
not I_12440 (I214322,I214373);
DFFARX1 I_12441 (I92942,I2859,I214330,I214404,);
not I_12442 (I214412,I92936);
nor I_12443 (I214429,I214356,I214412);
not I_12444 (I214446,I92930);
not I_12445 (I214463,I92927);
nand I_12446 (I214480,I214463,I92930);
nor I_12447 (I214497,I214412,I214480);
nor I_12448 (I214514,I214404,I214497);
DFFARX1 I_12449 (I214463,I2859,I214330,I214319,);
nor I_12450 (I214545,I92927,I92921);
nand I_12451 (I214562,I214545,I92939);
nor I_12452 (I214579,I214562,I214446);
nand I_12453 (I214304,I214579,I92936);
DFFARX1 I_12454 (I214562,I2859,I214330,I214316,);
nand I_12455 (I214624,I214446,I92927);
nor I_12456 (I214641,I214446,I92927);
nand I_12457 (I214310,I214429,I214641);
not I_12458 (I214672,I92933);
nor I_12459 (I214689,I214672,I214624);
DFFARX1 I_12460 (I214689,I2859,I214330,I214298,);
nor I_12461 (I214720,I214672,I92918);
and I_12462 (I214737,I214720,I92924);
or I_12463 (I214754,I214737,I92921);
DFFARX1 I_12464 (I214754,I2859,I214330,I214780,);
nor I_12465 (I214788,I214780,I214404);
nor I_12466 (I214307,I214356,I214788);
not I_12467 (I214819,I214780);
nor I_12468 (I214836,I214819,I214514);
DFFARX1 I_12469 (I214836,I2859,I214330,I214313,);
nand I_12470 (I214867,I214819,I214446);
nor I_12471 (I214301,I214672,I214867);
not I_12472 (I214925,I2866);
DFFARX1 I_12473 (I393850,I2859,I214925,I214951,);
DFFARX1 I_12474 (I214951,I2859,I214925,I214968,);
not I_12475 (I214917,I214968);
DFFARX1 I_12476 (I393838,I2859,I214925,I214999,);
not I_12477 (I215007,I393835);
nor I_12478 (I215024,I214951,I215007);
not I_12479 (I215041,I393847);
not I_12480 (I215058,I393844);
nand I_12481 (I215075,I215058,I393847);
nor I_12482 (I215092,I215007,I215075);
nor I_12483 (I215109,I214999,I215092);
DFFARX1 I_12484 (I215058,I2859,I214925,I214914,);
nor I_12485 (I215140,I393844,I393853);
nand I_12486 (I215157,I215140,I393856);
nor I_12487 (I215174,I215157,I215041);
nand I_12488 (I214899,I215174,I393835);
DFFARX1 I_12489 (I215157,I2859,I214925,I214911,);
nand I_12490 (I215219,I215041,I393844);
nor I_12491 (I215236,I215041,I393844);
nand I_12492 (I214905,I215024,I215236);
not I_12493 (I215267,I393859);
nor I_12494 (I215284,I215267,I215219);
DFFARX1 I_12495 (I215284,I2859,I214925,I214893,);
nor I_12496 (I215315,I215267,I393862);
and I_12497 (I215332,I215315,I393841);
or I_12498 (I215349,I215332,I393835);
DFFARX1 I_12499 (I215349,I2859,I214925,I215375,);
nor I_12500 (I215383,I215375,I214999);
nor I_12501 (I214902,I214951,I215383);
not I_12502 (I215414,I215375);
nor I_12503 (I215431,I215414,I215109);
DFFARX1 I_12504 (I215431,I2859,I214925,I214908,);
nand I_12505 (I215462,I215414,I215041);
nor I_12506 (I214896,I215267,I215462);
not I_12507 (I215520,I2866);
DFFARX1 I_12508 (I101248,I2859,I215520,I215546,);
DFFARX1 I_12509 (I215546,I2859,I215520,I215563,);
not I_12510 (I215512,I215563);
DFFARX1 I_12511 (I101272,I2859,I215520,I215594,);
not I_12512 (I215602,I101266);
nor I_12513 (I215619,I215546,I215602);
not I_12514 (I215636,I101260);
not I_12515 (I215653,I101257);
nand I_12516 (I215670,I215653,I101260);
nor I_12517 (I215687,I215602,I215670);
nor I_12518 (I215704,I215594,I215687);
DFFARX1 I_12519 (I215653,I2859,I215520,I215509,);
nor I_12520 (I215735,I101257,I101251);
nand I_12521 (I215752,I215735,I101269);
nor I_12522 (I215769,I215752,I215636);
nand I_12523 (I215494,I215769,I101266);
DFFARX1 I_12524 (I215752,I2859,I215520,I215506,);
nand I_12525 (I215814,I215636,I101257);
nor I_12526 (I215831,I215636,I101257);
nand I_12527 (I215500,I215619,I215831);
not I_12528 (I215862,I101263);
nor I_12529 (I215879,I215862,I215814);
DFFARX1 I_12530 (I215879,I2859,I215520,I215488,);
nor I_12531 (I215910,I215862,I101248);
and I_12532 (I215927,I215910,I101254);
or I_12533 (I215944,I215927,I101251);
DFFARX1 I_12534 (I215944,I2859,I215520,I215970,);
nor I_12535 (I215978,I215970,I215594);
nor I_12536 (I215497,I215546,I215978);
not I_12537 (I216009,I215970);
nor I_12538 (I216026,I216009,I215704);
DFFARX1 I_12539 (I216026,I2859,I215520,I215503,);
nand I_12540 (I216057,I216009,I215636);
nor I_12541 (I215491,I215862,I216057);
not I_12542 (I216115,I2866);
DFFARX1 I_12543 (I58426,I2859,I216115,I216141,);
DFFARX1 I_12544 (I216141,I2859,I216115,I216158,);
not I_12545 (I216107,I216158);
DFFARX1 I_12546 (I58414,I2859,I216115,I216189,);
not I_12547 (I216197,I58420);
nor I_12548 (I216214,I216141,I216197);
not I_12549 (I216231,I58411);
not I_12550 (I216248,I58429);
nand I_12551 (I216265,I216248,I58411);
nor I_12552 (I216282,I216197,I216265);
nor I_12553 (I216299,I216189,I216282);
DFFARX1 I_12554 (I216248,I2859,I216115,I216104,);
nor I_12555 (I216330,I58429,I58408);
nand I_12556 (I216347,I216330,I58435);
nor I_12557 (I216364,I216347,I216231);
nand I_12558 (I216089,I216364,I58420);
DFFARX1 I_12559 (I216347,I2859,I216115,I216101,);
nand I_12560 (I216409,I216231,I58429);
nor I_12561 (I216426,I216231,I58429);
nand I_12562 (I216095,I216214,I216426);
not I_12563 (I216457,I58423);
nor I_12564 (I216474,I216457,I216409);
DFFARX1 I_12565 (I216474,I2859,I216115,I216083,);
nor I_12566 (I216505,I216457,I58408);
and I_12567 (I216522,I216505,I58432);
or I_12568 (I216539,I216522,I58417);
DFFARX1 I_12569 (I216539,I2859,I216115,I216565,);
nor I_12570 (I216573,I216565,I216189);
nor I_12571 (I216092,I216141,I216573);
not I_12572 (I216604,I216565);
nor I_12573 (I216621,I216604,I216299);
DFFARX1 I_12574 (I216621,I2859,I216115,I216098,);
nand I_12575 (I216652,I216604,I216231);
nor I_12576 (I216086,I216457,I216652);
not I_12577 (I216710,I2866);
DFFARX1 I_12578 (I526325,I2859,I216710,I216736,);
DFFARX1 I_12579 (I216736,I2859,I216710,I216753,);
not I_12580 (I216702,I216753);
DFFARX1 I_12581 (I526331,I2859,I216710,I216784,);
not I_12582 (I216792,I526319);
nor I_12583 (I216809,I216736,I216792);
not I_12584 (I216826,I526322);
not I_12585 (I216843,I526328);
nand I_12586 (I216860,I216843,I526322);
nor I_12587 (I216877,I216792,I216860);
nor I_12588 (I216894,I216784,I216877);
DFFARX1 I_12589 (I216843,I2859,I216710,I216699,);
nor I_12590 (I216925,I526328,I526319);
nand I_12591 (I216942,I216925,I526337);
nor I_12592 (I216959,I216942,I216826);
nand I_12593 (I216684,I216959,I526319);
DFFARX1 I_12594 (I216942,I2859,I216710,I216696,);
nand I_12595 (I217004,I216826,I526328);
nor I_12596 (I217021,I216826,I526328);
nand I_12597 (I216690,I216809,I217021);
not I_12598 (I217052,I526316);
nor I_12599 (I217069,I217052,I217004);
DFFARX1 I_12600 (I217069,I2859,I216710,I216678,);
nor I_12601 (I217100,I217052,I526340);
and I_12602 (I217117,I217100,I526316);
or I_12603 (I217134,I217117,I526334);
DFFARX1 I_12604 (I217134,I2859,I216710,I217160,);
nor I_12605 (I217168,I217160,I216784);
nor I_12606 (I216687,I216736,I217168);
not I_12607 (I217199,I217160);
nor I_12608 (I217216,I217199,I216894);
DFFARX1 I_12609 (I217216,I2859,I216710,I216693,);
nand I_12610 (I217247,I217199,I216826);
nor I_12611 (I216681,I217052,I217247);
not I_12612 (I217305,I2866);
DFFARX1 I_12613 (I291623,I2859,I217305,I217331,);
DFFARX1 I_12614 (I217331,I2859,I217305,I217348,);
not I_12615 (I217297,I217348);
DFFARX1 I_12616 (I291617,I2859,I217305,I217379,);
not I_12617 (I217387,I291614);
nor I_12618 (I217404,I217331,I217387);
not I_12619 (I217421,I291626);
not I_12620 (I217438,I291629);
nand I_12621 (I217455,I217438,I291626);
nor I_12622 (I217472,I217387,I217455);
nor I_12623 (I217489,I217379,I217472);
DFFARX1 I_12624 (I217438,I2859,I217305,I217294,);
nor I_12625 (I217520,I291629,I291638);
nand I_12626 (I217537,I217520,I291632);
nor I_12627 (I217554,I217537,I217421);
nand I_12628 (I217279,I217554,I291614);
DFFARX1 I_12629 (I217537,I2859,I217305,I217291,);
nand I_12630 (I217599,I217421,I291629);
nor I_12631 (I217616,I217421,I291629);
nand I_12632 (I217285,I217404,I217616);
not I_12633 (I217647,I291620);
nor I_12634 (I217664,I217647,I217599);
DFFARX1 I_12635 (I217664,I2859,I217305,I217273,);
nor I_12636 (I217695,I217647,I291635);
and I_12637 (I217712,I217695,I291614);
or I_12638 (I217729,I217712,I291617);
DFFARX1 I_12639 (I217729,I2859,I217305,I217755,);
nor I_12640 (I217763,I217755,I217379);
nor I_12641 (I217282,I217331,I217763);
not I_12642 (I217794,I217755);
nor I_12643 (I217811,I217794,I217489);
DFFARX1 I_12644 (I217811,I2859,I217305,I217288,);
nand I_12645 (I217842,I217794,I217421);
nor I_12646 (I217276,I217647,I217842);
not I_12647 (I217900,I2866);
DFFARX1 I_12648 (I236129,I2859,I217900,I217926,);
DFFARX1 I_12649 (I217926,I2859,I217900,I217943,);
not I_12650 (I217892,I217943);
DFFARX1 I_12651 (I236141,I2859,I217900,I217974,);
not I_12652 (I217982,I236126);
nor I_12653 (I217999,I217926,I217982);
not I_12654 (I218016,I236144);
not I_12655 (I218033,I236135);
nand I_12656 (I218050,I218033,I236144);
nor I_12657 (I218067,I217982,I218050);
nor I_12658 (I218084,I217974,I218067);
DFFARX1 I_12659 (I218033,I2859,I217900,I217889,);
nor I_12660 (I218115,I236135,I236147);
nand I_12661 (I218132,I218115,I236150);
nor I_12662 (I218149,I218132,I218016);
nand I_12663 (I217874,I218149,I236126);
DFFARX1 I_12664 (I218132,I2859,I217900,I217886,);
nand I_12665 (I218194,I218016,I236135);
nor I_12666 (I218211,I218016,I236135);
nand I_12667 (I217880,I217999,I218211);
not I_12668 (I218242,I236126);
nor I_12669 (I218259,I218242,I218194);
DFFARX1 I_12670 (I218259,I2859,I217900,I217868,);
nor I_12671 (I218290,I218242,I236138);
and I_12672 (I218307,I218290,I236132);
or I_12673 (I218324,I218307,I236129);
DFFARX1 I_12674 (I218324,I2859,I217900,I218350,);
nor I_12675 (I218358,I218350,I217974);
nor I_12676 (I217877,I217926,I218358);
not I_12677 (I218389,I218350);
nor I_12678 (I218406,I218389,I218084);
DFFARX1 I_12679 (I218406,I2859,I217900,I217883,);
nand I_12680 (I218437,I218389,I218016);
nor I_12681 (I217871,I218242,I218437);
not I_12682 (I218495,I2866);
DFFARX1 I_12683 (I175963,I2859,I218495,I218521,);
DFFARX1 I_12684 (I218521,I2859,I218495,I218538,);
not I_12685 (I218487,I218538);
DFFARX1 I_12686 (I175987,I2859,I218495,I218569,);
not I_12687 (I218577,I175966);
nor I_12688 (I218594,I218521,I218577);
not I_12689 (I218611,I175972);
not I_12690 (I218628,I175978);
nand I_12691 (I218645,I218628,I175972);
nor I_12692 (I218662,I218577,I218645);
nor I_12693 (I218679,I218569,I218662);
DFFARX1 I_12694 (I218628,I2859,I218495,I218484,);
nor I_12695 (I218710,I175978,I175990);
nand I_12696 (I218727,I218710,I175984);
nor I_12697 (I218744,I218727,I218611);
nand I_12698 (I218469,I218744,I175966);
DFFARX1 I_12699 (I218727,I2859,I218495,I218481,);
nand I_12700 (I218789,I218611,I175978);
nor I_12701 (I218806,I218611,I175978);
nand I_12702 (I218475,I218594,I218806);
not I_12703 (I218837,I175969);
nor I_12704 (I218854,I218837,I218789);
DFFARX1 I_12705 (I218854,I2859,I218495,I218463,);
nor I_12706 (I218885,I218837,I175963);
and I_12707 (I218902,I218885,I175981);
or I_12708 (I218919,I218902,I175975);
DFFARX1 I_12709 (I218919,I2859,I218495,I218945,);
nor I_12710 (I218953,I218945,I218569);
nor I_12711 (I218472,I218521,I218953);
not I_12712 (I218984,I218945);
nor I_12713 (I219001,I218984,I218679);
DFFARX1 I_12714 (I219001,I2859,I218495,I218478,);
nand I_12715 (I219032,I218984,I218611);
nor I_12716 (I218466,I218837,I219032);
not I_12717 (I219090,I2866);
DFFARX1 I_12718 (I501514,I2859,I219090,I219116,);
DFFARX1 I_12719 (I219116,I2859,I219090,I219133,);
not I_12720 (I219082,I219133);
DFFARX1 I_12721 (I501496,I2859,I219090,I219164,);
not I_12722 (I219172,I501502);
nor I_12723 (I219189,I219116,I219172);
not I_12724 (I219206,I501517);
not I_12725 (I219223,I501508);
nand I_12726 (I219240,I219223,I501517);
nor I_12727 (I219257,I219172,I219240);
nor I_12728 (I219274,I219164,I219257);
DFFARX1 I_12729 (I219223,I2859,I219090,I219079,);
nor I_12730 (I219305,I501508,I501520);
nand I_12731 (I219322,I219305,I501499);
nor I_12732 (I219339,I219322,I219206);
nand I_12733 (I219064,I219339,I501502);
DFFARX1 I_12734 (I219322,I2859,I219090,I219076,);
nand I_12735 (I219384,I219206,I501508);
nor I_12736 (I219401,I219206,I501508);
nand I_12737 (I219070,I219189,I219401);
not I_12738 (I219432,I501505);
nor I_12739 (I219449,I219432,I219384);
DFFARX1 I_12740 (I219449,I2859,I219090,I219058,);
nor I_12741 (I219480,I219432,I501511);
and I_12742 (I219497,I219480,I501496);
or I_12743 (I219514,I219497,I501499);
DFFARX1 I_12744 (I219514,I2859,I219090,I219540,);
nor I_12745 (I219548,I219540,I219164);
nor I_12746 (I219067,I219116,I219548);
not I_12747 (I219579,I219540);
nor I_12748 (I219596,I219579,I219274);
DFFARX1 I_12749 (I219596,I2859,I219090,I219073,);
nand I_12750 (I219627,I219579,I219206);
nor I_12751 (I219061,I219432,I219627);
not I_12752 (I219685,I2866);
DFFARX1 I_12753 (I104818,I2859,I219685,I219711,);
DFFARX1 I_12754 (I219711,I2859,I219685,I219728,);
not I_12755 (I219677,I219728);
DFFARX1 I_12756 (I104842,I2859,I219685,I219759,);
not I_12757 (I219767,I104836);
nor I_12758 (I219784,I219711,I219767);
not I_12759 (I219801,I104830);
not I_12760 (I219818,I104827);
nand I_12761 (I219835,I219818,I104830);
nor I_12762 (I219852,I219767,I219835);
nor I_12763 (I219869,I219759,I219852);
DFFARX1 I_12764 (I219818,I2859,I219685,I219674,);
nor I_12765 (I219900,I104827,I104821);
nand I_12766 (I219917,I219900,I104839);
nor I_12767 (I219934,I219917,I219801);
nand I_12768 (I219659,I219934,I104836);
DFFARX1 I_12769 (I219917,I2859,I219685,I219671,);
nand I_12770 (I219979,I219801,I104827);
nor I_12771 (I219996,I219801,I104827);
nand I_12772 (I219665,I219784,I219996);
not I_12773 (I220027,I104833);
nor I_12774 (I220044,I220027,I219979);
DFFARX1 I_12775 (I220044,I2859,I219685,I219653,);
nor I_12776 (I220075,I220027,I104818);
and I_12777 (I220092,I220075,I104824);
or I_12778 (I220109,I220092,I104821);
DFFARX1 I_12779 (I220109,I2859,I219685,I220135,);
nor I_12780 (I220143,I220135,I219759);
nor I_12781 (I219662,I219711,I220143);
not I_12782 (I220174,I220135);
nor I_12783 (I220191,I220174,I219869);
DFFARX1 I_12784 (I220191,I2859,I219685,I219668,);
nand I_12785 (I220222,I220174,I219801);
nor I_12786 (I219656,I220027,I220222);
not I_12787 (I220280,I2866);
DFFARX1 I_12788 (I304917,I2859,I220280,I220306,);
DFFARX1 I_12789 (I220306,I2859,I220280,I220323,);
not I_12790 (I220272,I220323);
DFFARX1 I_12791 (I304911,I2859,I220280,I220354,);
not I_12792 (I220362,I304908);
nor I_12793 (I220379,I220306,I220362);
not I_12794 (I220396,I304920);
not I_12795 (I220413,I304923);
nand I_12796 (I220430,I220413,I304920);
nor I_12797 (I220447,I220362,I220430);
nor I_12798 (I220464,I220354,I220447);
DFFARX1 I_12799 (I220413,I2859,I220280,I220269,);
nor I_12800 (I220495,I304923,I304932);
nand I_12801 (I220512,I220495,I304926);
nor I_12802 (I220529,I220512,I220396);
nand I_12803 (I220254,I220529,I304908);
DFFARX1 I_12804 (I220512,I2859,I220280,I220266,);
nand I_12805 (I220574,I220396,I304923);
nor I_12806 (I220591,I220396,I304923);
nand I_12807 (I220260,I220379,I220591);
not I_12808 (I220622,I304914);
nor I_12809 (I220639,I220622,I220574);
DFFARX1 I_12810 (I220639,I2859,I220280,I220248,);
nor I_12811 (I220670,I220622,I304929);
and I_12812 (I220687,I220670,I304908);
or I_12813 (I220704,I220687,I304911);
DFFARX1 I_12814 (I220704,I2859,I220280,I220730,);
nor I_12815 (I220738,I220730,I220354);
nor I_12816 (I220257,I220306,I220738);
not I_12817 (I220769,I220730);
nor I_12818 (I220786,I220769,I220464);
DFFARX1 I_12819 (I220786,I2859,I220280,I220263,);
nand I_12820 (I220817,I220769,I220396);
nor I_12821 (I220251,I220622,I220817);
not I_12822 (I220875,I2866);
DFFARX1 I_12823 (I347417,I2859,I220875,I220901,);
DFFARX1 I_12824 (I220901,I2859,I220875,I220918,);
not I_12825 (I220867,I220918);
DFFARX1 I_12826 (I347414,I2859,I220875,I220949,);
not I_12827 (I220957,I347414);
nor I_12828 (I220974,I220901,I220957);
not I_12829 (I220991,I347411);
not I_12830 (I221008,I347426);
nand I_12831 (I221025,I221008,I347411);
nor I_12832 (I221042,I220957,I221025);
nor I_12833 (I221059,I220949,I221042);
DFFARX1 I_12834 (I221008,I2859,I220875,I220864,);
nor I_12835 (I221090,I347426,I347420);
nand I_12836 (I221107,I221090,I347408);
nor I_12837 (I221124,I221107,I220991);
nand I_12838 (I220849,I221124,I347414);
DFFARX1 I_12839 (I221107,I2859,I220875,I220861,);
nand I_12840 (I221169,I220991,I347426);
nor I_12841 (I221186,I220991,I347426);
nand I_12842 (I220855,I220974,I221186);
not I_12843 (I221217,I347429);
nor I_12844 (I221234,I221217,I221169);
DFFARX1 I_12845 (I221234,I2859,I220875,I220843,);
nor I_12846 (I221265,I221217,I347408);
and I_12847 (I221282,I221265,I347423);
or I_12848 (I221299,I221282,I347411);
DFFARX1 I_12849 (I221299,I2859,I220875,I221325,);
nor I_12850 (I221333,I221325,I220949);
nor I_12851 (I220852,I220901,I221333);
not I_12852 (I221364,I221325);
nor I_12853 (I221381,I221364,I221059);
DFFARX1 I_12854 (I221381,I2859,I220875,I220858,);
nand I_12855 (I221412,I221364,I220991);
nor I_12856 (I220846,I221217,I221412);
not I_12857 (I221470,I2866);
DFFARX1 I_12858 (I69713,I2859,I221470,I221496,);
DFFARX1 I_12859 (I221496,I2859,I221470,I221513,);
not I_12860 (I221462,I221513);
DFFARX1 I_12861 (I69737,I2859,I221470,I221544,);
not I_12862 (I221552,I69731);
nor I_12863 (I221569,I221496,I221552);
not I_12864 (I221586,I69725);
not I_12865 (I221603,I69722);
nand I_12866 (I221620,I221603,I69725);
nor I_12867 (I221637,I221552,I221620);
nor I_12868 (I221654,I221544,I221637);
DFFARX1 I_12869 (I221603,I2859,I221470,I221459,);
nor I_12870 (I221685,I69722,I69716);
nand I_12871 (I221702,I221685,I69734);
nor I_12872 (I221719,I221702,I221586);
nand I_12873 (I221444,I221719,I69731);
DFFARX1 I_12874 (I221702,I2859,I221470,I221456,);
nand I_12875 (I221764,I221586,I69722);
nor I_12876 (I221781,I221586,I69722);
nand I_12877 (I221450,I221569,I221781);
not I_12878 (I221812,I69728);
nor I_12879 (I221829,I221812,I221764);
DFFARX1 I_12880 (I221829,I2859,I221470,I221438,);
nor I_12881 (I221860,I221812,I69713);
and I_12882 (I221877,I221860,I69719);
or I_12883 (I221894,I221877,I69716);
DFFARX1 I_12884 (I221894,I2859,I221470,I221920,);
nor I_12885 (I221928,I221920,I221544);
nor I_12886 (I221447,I221496,I221928);
not I_12887 (I221959,I221920);
nor I_12888 (I221976,I221959,I221654);
DFFARX1 I_12889 (I221976,I2859,I221470,I221453,);
nand I_12890 (I222007,I221959,I221586);
nor I_12891 (I221441,I221812,I222007);
not I_12892 (I222065,I2866);
DFFARX1 I_12893 (I235551,I2859,I222065,I222091,);
DFFARX1 I_12894 (I222091,I2859,I222065,I222108,);
not I_12895 (I222057,I222108);
DFFARX1 I_12896 (I235563,I2859,I222065,I222139,);
not I_12897 (I222147,I235548);
nor I_12898 (I222164,I222091,I222147);
not I_12899 (I222181,I235566);
not I_12900 (I222198,I235557);
nand I_12901 (I222215,I222198,I235566);
nor I_12902 (I222232,I222147,I222215);
nor I_12903 (I222249,I222139,I222232);
DFFARX1 I_12904 (I222198,I2859,I222065,I222054,);
nor I_12905 (I222280,I235557,I235569);
nand I_12906 (I222297,I222280,I235572);
nor I_12907 (I222314,I222297,I222181);
nand I_12908 (I222039,I222314,I235548);
DFFARX1 I_12909 (I222297,I2859,I222065,I222051,);
nand I_12910 (I222359,I222181,I235557);
nor I_12911 (I222376,I222181,I235557);
nand I_12912 (I222045,I222164,I222376);
not I_12913 (I222407,I235548);
nor I_12914 (I222424,I222407,I222359);
DFFARX1 I_12915 (I222424,I2859,I222065,I222033,);
nor I_12916 (I222455,I222407,I235560);
and I_12917 (I222472,I222455,I235554);
or I_12918 (I222489,I222472,I235551);
DFFARX1 I_12919 (I222489,I2859,I222065,I222515,);
nor I_12920 (I222523,I222515,I222139);
nor I_12921 (I222042,I222091,I222523);
not I_12922 (I222554,I222515);
nor I_12923 (I222571,I222554,I222249);
DFFARX1 I_12924 (I222571,I2859,I222065,I222048,);
nand I_12925 (I222602,I222554,I222181);
nor I_12926 (I222036,I222407,I222602);
not I_12927 (I222660,I2866);
DFFARX1 I_12928 (I90538,I2859,I222660,I222686,);
DFFARX1 I_12929 (I222686,I2859,I222660,I222703,);
not I_12930 (I222652,I222703);
DFFARX1 I_12931 (I90562,I2859,I222660,I222734,);
not I_12932 (I222742,I90556);
nor I_12933 (I222759,I222686,I222742);
not I_12934 (I222776,I90550);
not I_12935 (I222793,I90547);
nand I_12936 (I222810,I222793,I90550);
nor I_12937 (I222827,I222742,I222810);
nor I_12938 (I222844,I222734,I222827);
DFFARX1 I_12939 (I222793,I2859,I222660,I222649,);
nor I_12940 (I222875,I90547,I90541);
nand I_12941 (I222892,I222875,I90559);
nor I_12942 (I222909,I222892,I222776);
nand I_12943 (I222634,I222909,I90556);
DFFARX1 I_12944 (I222892,I2859,I222660,I222646,);
nand I_12945 (I222954,I222776,I90547);
nor I_12946 (I222971,I222776,I90547);
nand I_12947 (I222640,I222759,I222971);
not I_12948 (I223002,I90553);
nor I_12949 (I223019,I223002,I222954);
DFFARX1 I_12950 (I223019,I2859,I222660,I222628,);
nor I_12951 (I223050,I223002,I90538);
and I_12952 (I223067,I223050,I90544);
or I_12953 (I223084,I223067,I90541);
DFFARX1 I_12954 (I223084,I2859,I222660,I223110,);
nor I_12955 (I223118,I223110,I222734);
nor I_12956 (I222637,I222686,I223118);
not I_12957 (I223149,I223110);
nor I_12958 (I223166,I223149,I222844);
DFFARX1 I_12959 (I223166,I2859,I222660,I222643,);
nand I_12960 (I223197,I223149,I222776);
nor I_12961 (I222631,I223002,I223197);
not I_12962 (I223255,I2866);
DFFARX1 I_12963 (I255781,I2859,I223255,I223281,);
DFFARX1 I_12964 (I223281,I2859,I223255,I223298,);
not I_12965 (I223247,I223298);
DFFARX1 I_12966 (I255793,I2859,I223255,I223329,);
not I_12967 (I223337,I255778);
nor I_12968 (I223354,I223281,I223337);
not I_12969 (I223371,I255796);
not I_12970 (I223388,I255787);
nand I_12971 (I223405,I223388,I255796);
nor I_12972 (I223422,I223337,I223405);
nor I_12973 (I223439,I223329,I223422);
DFFARX1 I_12974 (I223388,I2859,I223255,I223244,);
nor I_12975 (I223470,I255787,I255799);
nand I_12976 (I223487,I223470,I255802);
nor I_12977 (I223504,I223487,I223371);
nand I_12978 (I223229,I223504,I255778);
DFFARX1 I_12979 (I223487,I2859,I223255,I223241,);
nand I_12980 (I223549,I223371,I255787);
nor I_12981 (I223566,I223371,I255787);
nand I_12982 (I223235,I223354,I223566);
not I_12983 (I223597,I255778);
nor I_12984 (I223614,I223597,I223549);
DFFARX1 I_12985 (I223614,I2859,I223255,I223223,);
nor I_12986 (I223645,I223597,I255790);
and I_12987 (I223662,I223645,I255784);
or I_12988 (I223679,I223662,I255781);
DFFARX1 I_12989 (I223679,I2859,I223255,I223705,);
nor I_12990 (I223713,I223705,I223329);
nor I_12991 (I223232,I223281,I223713);
not I_12992 (I223744,I223705);
nor I_12993 (I223761,I223744,I223439);
DFFARX1 I_12994 (I223761,I2859,I223255,I223238,);
nand I_12995 (I223792,I223744,I223371);
nor I_12996 (I223226,I223597,I223792);
not I_12997 (I223850,I2866);
DFFARX1 I_12998 (I446076,I2859,I223850,I223876,);
DFFARX1 I_12999 (I223876,I2859,I223850,I223893,);
not I_13000 (I223842,I223893);
DFFARX1 I_13001 (I446079,I2859,I223850,I223924,);
not I_13002 (I223932,I446082);
nor I_13003 (I223949,I223876,I223932);
not I_13004 (I223966,I446094);
not I_13005 (I223983,I446085);
nand I_13006 (I224000,I223983,I446094);
nor I_13007 (I224017,I223932,I224000);
nor I_13008 (I224034,I223924,I224017);
DFFARX1 I_13009 (I223983,I2859,I223850,I223839,);
nor I_13010 (I224065,I446085,I446091);
nand I_13011 (I224082,I224065,I446079);
nor I_13012 (I224099,I224082,I223966);
nand I_13013 (I223824,I224099,I446082);
DFFARX1 I_13014 (I224082,I2859,I223850,I223836,);
nand I_13015 (I224144,I223966,I446085);
nor I_13016 (I224161,I223966,I446085);
nand I_13017 (I223830,I223949,I224161);
not I_13018 (I224192,I446082);
nor I_13019 (I224209,I224192,I224144);
DFFARX1 I_13020 (I224209,I2859,I223850,I223818,);
nor I_13021 (I224240,I224192,I446088);
and I_13022 (I224257,I224240,I446076);
or I_13023 (I224274,I224257,I446097);
DFFARX1 I_13024 (I224274,I2859,I223850,I224300,);
nor I_13025 (I224308,I224300,I223924);
nor I_13026 (I223827,I223876,I224308);
not I_13027 (I224339,I224300);
nor I_13028 (I224356,I224339,I224034);
DFFARX1 I_13029 (I224356,I2859,I223850,I223833,);
nand I_13030 (I224387,I224339,I223966);
nor I_13031 (I223821,I224192,I224387);
not I_13032 (I224445,I2866);
DFFARX1 I_13033 (I367970,I2859,I224445,I224471,);
DFFARX1 I_13034 (I224471,I2859,I224445,I224488,);
not I_13035 (I224437,I224488);
DFFARX1 I_13036 (I367967,I2859,I224445,I224519,);
not I_13037 (I224527,I367967);
nor I_13038 (I224544,I224471,I224527);
not I_13039 (I224561,I367964);
not I_13040 (I224578,I367979);
nand I_13041 (I224595,I224578,I367964);
nor I_13042 (I224612,I224527,I224595);
nor I_13043 (I224629,I224519,I224612);
DFFARX1 I_13044 (I224578,I2859,I224445,I224434,);
nor I_13045 (I224660,I367979,I367973);
nand I_13046 (I224677,I224660,I367961);
nor I_13047 (I224694,I224677,I224561);
nand I_13048 (I224419,I224694,I367967);
DFFARX1 I_13049 (I224677,I2859,I224445,I224431,);
nand I_13050 (I224739,I224561,I367979);
nor I_13051 (I224756,I224561,I367979);
nand I_13052 (I224425,I224544,I224756);
not I_13053 (I224787,I367982);
nor I_13054 (I224804,I224787,I224739);
DFFARX1 I_13055 (I224804,I2859,I224445,I224413,);
nor I_13056 (I224835,I224787,I367961);
and I_13057 (I224852,I224835,I367976);
or I_13058 (I224869,I224852,I367964);
DFFARX1 I_13059 (I224869,I2859,I224445,I224895,);
nor I_13060 (I224903,I224895,I224519);
nor I_13061 (I224422,I224471,I224903);
not I_13062 (I224934,I224895);
nor I_13063 (I224951,I224934,I224629);
DFFARX1 I_13064 (I224951,I2859,I224445,I224428,);
nand I_13065 (I224982,I224934,I224561);
nor I_13066 (I224416,I224787,I224982);
not I_13067 (I225040,I2866);
DFFARX1 I_13068 (I292779,I2859,I225040,I225066,);
DFFARX1 I_13069 (I225066,I2859,I225040,I225083,);
not I_13070 (I225032,I225083);
DFFARX1 I_13071 (I292773,I2859,I225040,I225114,);
not I_13072 (I225122,I292770);
nor I_13073 (I225139,I225066,I225122);
not I_13074 (I225156,I292782);
not I_13075 (I225173,I292785);
nand I_13076 (I225190,I225173,I292782);
nor I_13077 (I225207,I225122,I225190);
nor I_13078 (I225224,I225114,I225207);
DFFARX1 I_13079 (I225173,I2859,I225040,I225029,);
nor I_13080 (I225255,I292785,I292794);
nand I_13081 (I225272,I225255,I292788);
nor I_13082 (I225289,I225272,I225156);
nand I_13083 (I225014,I225289,I292770);
DFFARX1 I_13084 (I225272,I2859,I225040,I225026,);
nand I_13085 (I225334,I225156,I292785);
nor I_13086 (I225351,I225156,I292785);
nand I_13087 (I225020,I225139,I225351);
not I_13088 (I225382,I292776);
nor I_13089 (I225399,I225382,I225334);
DFFARX1 I_13090 (I225399,I2859,I225040,I225008,);
nor I_13091 (I225430,I225382,I292791);
and I_13092 (I225447,I225430,I292770);
or I_13093 (I225464,I225447,I292773);
DFFARX1 I_13094 (I225464,I2859,I225040,I225490,);
nor I_13095 (I225498,I225490,I225114);
nor I_13096 (I225017,I225066,I225498);
not I_13097 (I225529,I225490);
nor I_13098 (I225546,I225529,I225224);
DFFARX1 I_13099 (I225546,I2859,I225040,I225023,);
nand I_13100 (I225577,I225529,I225156);
nor I_13101 (I225011,I225382,I225577);
not I_13102 (I225635,I2866);
DFFARX1 I_13103 (I437661,I2859,I225635,I225661,);
DFFARX1 I_13104 (I225661,I2859,I225635,I225678,);
not I_13105 (I225627,I225678);
DFFARX1 I_13106 (I437664,I2859,I225635,I225709,);
not I_13107 (I225717,I437667);
nor I_13108 (I225734,I225661,I225717);
not I_13109 (I225751,I437679);
not I_13110 (I225768,I437670);
nand I_13111 (I225785,I225768,I437679);
nor I_13112 (I225802,I225717,I225785);
nor I_13113 (I225819,I225709,I225802);
DFFARX1 I_13114 (I225768,I2859,I225635,I225624,);
nor I_13115 (I225850,I437670,I437676);
nand I_13116 (I225867,I225850,I437664);
nor I_13117 (I225884,I225867,I225751);
nand I_13118 (I225609,I225884,I437667);
DFFARX1 I_13119 (I225867,I2859,I225635,I225621,);
nand I_13120 (I225929,I225751,I437670);
nor I_13121 (I225946,I225751,I437670);
nand I_13122 (I225615,I225734,I225946);
not I_13123 (I225977,I437667);
nor I_13124 (I225994,I225977,I225929);
DFFARX1 I_13125 (I225994,I2859,I225635,I225603,);
nor I_13126 (I226025,I225977,I437673);
and I_13127 (I226042,I226025,I437661);
or I_13128 (I226059,I226042,I437682);
DFFARX1 I_13129 (I226059,I2859,I225635,I226085,);
nor I_13130 (I226093,I226085,I225709);
nor I_13131 (I225612,I225661,I226093);
not I_13132 (I226124,I226085);
nor I_13133 (I226141,I226124,I225819);
DFFARX1 I_13134 (I226141,I2859,I225635,I225618,);
nand I_13135 (I226172,I226124,I225751);
nor I_13136 (I225606,I225977,I226172);
not I_13137 (I226230,I2866);
DFFARX1 I_13138 (I375348,I2859,I226230,I226256,);
DFFARX1 I_13139 (I226256,I2859,I226230,I226273,);
not I_13140 (I226222,I226273);
DFFARX1 I_13141 (I375345,I2859,I226230,I226304,);
not I_13142 (I226312,I375345);
nor I_13143 (I226329,I226256,I226312);
not I_13144 (I226346,I375342);
not I_13145 (I226363,I375357);
nand I_13146 (I226380,I226363,I375342);
nor I_13147 (I226397,I226312,I226380);
nor I_13148 (I226414,I226304,I226397);
DFFARX1 I_13149 (I226363,I2859,I226230,I226219,);
nor I_13150 (I226445,I375357,I375351);
nand I_13151 (I226462,I226445,I375339);
nor I_13152 (I226479,I226462,I226346);
nand I_13153 (I226204,I226479,I375345);
DFFARX1 I_13154 (I226462,I2859,I226230,I226216,);
nand I_13155 (I226524,I226346,I375357);
nor I_13156 (I226541,I226346,I375357);
nand I_13157 (I226210,I226329,I226541);
not I_13158 (I226572,I375360);
nor I_13159 (I226589,I226572,I226524);
DFFARX1 I_13160 (I226589,I2859,I226230,I226198,);
nor I_13161 (I226620,I226572,I375339);
and I_13162 (I226637,I226620,I375354);
or I_13163 (I226654,I226637,I375342);
DFFARX1 I_13164 (I226654,I2859,I226230,I226680,);
nor I_13165 (I226688,I226680,I226304);
nor I_13166 (I226207,I226256,I226688);
not I_13167 (I226719,I226680);
nor I_13168 (I226736,I226719,I226414);
DFFARX1 I_13169 (I226736,I2859,I226230,I226213,);
nand I_13170 (I226767,I226719,I226346);
nor I_13171 (I226201,I226572,I226767);
not I_13172 (I226825,I2866);
DFFARX1 I_13173 (I538384,I2859,I226825,I226851,);
DFFARX1 I_13174 (I226851,I2859,I226825,I226868,);
not I_13175 (I226817,I226868);
DFFARX1 I_13176 (I538390,I2859,I226825,I226899,);
not I_13177 (I226907,I538393);
nor I_13178 (I226924,I226851,I226907);
not I_13179 (I226941,I538396);
not I_13180 (I226958,I538381);
nand I_13181 (I226975,I226958,I538396);
nor I_13182 (I226992,I226907,I226975);
nor I_13183 (I227009,I226899,I226992);
DFFARX1 I_13184 (I226958,I2859,I226825,I226814,);
nor I_13185 (I227040,I538381,I538387);
nand I_13186 (I227057,I227040,I538369);
nor I_13187 (I227074,I227057,I226941);
nand I_13188 (I226799,I227074,I538393);
DFFARX1 I_13189 (I227057,I2859,I226825,I226811,);
nand I_13190 (I227119,I226941,I538381);
nor I_13191 (I227136,I226941,I538381);
nand I_13192 (I226805,I226924,I227136);
not I_13193 (I227167,I538369);
nor I_13194 (I227184,I227167,I227119);
DFFARX1 I_13195 (I227184,I2859,I226825,I226793,);
nor I_13196 (I227215,I227167,I538378);
and I_13197 (I227232,I227215,I538375);
or I_13198 (I227249,I227232,I538372);
DFFARX1 I_13199 (I227249,I2859,I226825,I227275,);
nor I_13200 (I227283,I227275,I226899);
nor I_13201 (I226802,I226851,I227283);
not I_13202 (I227314,I227275);
nor I_13203 (I227331,I227314,I227009);
DFFARX1 I_13204 (I227331,I2859,I226825,I226808,);
nand I_13205 (I227362,I227314,I226941);
nor I_13206 (I226796,I227167,I227362);
not I_13207 (I227420,I2866);
DFFARX1 I_13208 (I59616,I2859,I227420,I227446,);
DFFARX1 I_13209 (I227446,I2859,I227420,I227463,);
not I_13210 (I227412,I227463);
DFFARX1 I_13211 (I59604,I2859,I227420,I227494,);
not I_13212 (I227502,I59610);
nor I_13213 (I227519,I227446,I227502);
not I_13214 (I227536,I59601);
not I_13215 (I227553,I59619);
nand I_13216 (I227570,I227553,I59601);
nor I_13217 (I227587,I227502,I227570);
nor I_13218 (I227604,I227494,I227587);
DFFARX1 I_13219 (I227553,I2859,I227420,I227409,);
nor I_13220 (I227635,I59619,I59598);
nand I_13221 (I227652,I227635,I59625);
nor I_13222 (I227669,I227652,I227536);
nand I_13223 (I227394,I227669,I59610);
DFFARX1 I_13224 (I227652,I2859,I227420,I227406,);
nand I_13225 (I227714,I227536,I59619);
nor I_13226 (I227731,I227536,I59619);
nand I_13227 (I227400,I227519,I227731);
not I_13228 (I227762,I59613);
nor I_13229 (I227779,I227762,I227714);
DFFARX1 I_13230 (I227779,I2859,I227420,I227388,);
nor I_13231 (I227810,I227762,I59598);
and I_13232 (I227827,I227810,I59622);
or I_13233 (I227844,I227827,I59607);
DFFARX1 I_13234 (I227844,I2859,I227420,I227870,);
nor I_13235 (I227878,I227870,I227494);
nor I_13236 (I227397,I227446,I227878);
not I_13237 (I227909,I227870);
nor I_13238 (I227926,I227909,I227604);
DFFARX1 I_13239 (I227926,I2859,I227420,I227403,);
nand I_13240 (I227957,I227909,I227536);
nor I_13241 (I227391,I227762,I227957);
not I_13242 (I228015,I2866);
DFFARX1 I_13243 (I147724,I2859,I228015,I228041,);
DFFARX1 I_13244 (I228041,I2859,I228015,I228058,);
not I_13245 (I228007,I228058);
DFFARX1 I_13246 (I147712,I2859,I228015,I228089,);
not I_13247 (I228097,I147715);
nor I_13248 (I228114,I228041,I228097);
not I_13249 (I228131,I147718);
not I_13250 (I228148,I147730);
nand I_13251 (I228165,I228148,I147718);
nor I_13252 (I228182,I228097,I228165);
nor I_13253 (I228199,I228089,I228182);
DFFARX1 I_13254 (I228148,I2859,I228015,I228004,);
nor I_13255 (I228230,I147730,I147721);
nand I_13256 (I228247,I228230,I147709);
nor I_13257 (I228264,I228247,I228131);
nand I_13258 (I227989,I228264,I147715);
DFFARX1 I_13259 (I228247,I2859,I228015,I228001,);
nand I_13260 (I228309,I228131,I147730);
nor I_13261 (I228326,I228131,I147730);
nand I_13262 (I227995,I228114,I228326);
not I_13263 (I228357,I147727);
nor I_13264 (I228374,I228357,I228309);
DFFARX1 I_13265 (I228374,I2859,I228015,I227983,);
nor I_13266 (I228405,I228357,I147733);
and I_13267 (I228422,I228405,I147736);
or I_13268 (I228439,I228422,I147709);
DFFARX1 I_13269 (I228439,I2859,I228015,I228465,);
nor I_13270 (I228473,I228465,I228089);
nor I_13271 (I227992,I228041,I228473);
not I_13272 (I228504,I228465);
nor I_13273 (I228521,I228504,I228199);
DFFARX1 I_13274 (I228521,I2859,I228015,I227998,);
nand I_13275 (I228552,I228504,I228131);
nor I_13276 (I227986,I228357,I228552);
not I_13277 (I228610,I2866);
DFFARX1 I_13278 (I2836,I2859,I228610,I228636,);
DFFARX1 I_13279 (I228636,I2859,I228610,I228653,);
not I_13280 (I228602,I228653);
DFFARX1 I_13281 (I2804,I2859,I228610,I228684,);
not I_13282 (I228692,I2588);
nor I_13283 (I228709,I228636,I228692);
not I_13284 (I228726,I2028);
not I_13285 (I228743,I2356);
nand I_13286 (I228760,I228743,I2028);
nor I_13287 (I228777,I228692,I228760);
nor I_13288 (I228794,I228684,I228777);
DFFARX1 I_13289 (I228743,I2859,I228610,I228599,);
nor I_13290 (I228825,I2356,I1980);
nand I_13291 (I228842,I228825,I2300);
nor I_13292 (I228859,I228842,I228726);
nand I_13293 (I228584,I228859,I2588);
DFFARX1 I_13294 (I228842,I2859,I228610,I228596,);
nand I_13295 (I228904,I228726,I2356);
nor I_13296 (I228921,I228726,I2356);
nand I_13297 (I228590,I228709,I228921);
not I_13298 (I228952,I2724);
nor I_13299 (I228969,I228952,I228904);
DFFARX1 I_13300 (I228969,I2859,I228610,I228578,);
nor I_13301 (I229000,I228952,I1884);
and I_13302 (I229017,I229000,I1412);
or I_13303 (I229034,I229017,I1492);
DFFARX1 I_13304 (I229034,I2859,I228610,I229060,);
nor I_13305 (I229068,I229060,I228684);
nor I_13306 (I228587,I228636,I229068);
not I_13307 (I229099,I229060);
nor I_13308 (I229116,I229099,I228794);
DFFARX1 I_13309 (I229116,I2859,I228610,I228593,);
nand I_13310 (I229147,I229099,I228726);
nor I_13311 (I228581,I228952,I229147);
not I_13312 (I229205,I2866);
DFFARX1 I_13313 (I458742,I2859,I229205,I229231,);
DFFARX1 I_13314 (I229231,I2859,I229205,I229248,);
not I_13315 (I229197,I229248);
DFFARX1 I_13316 (I458724,I2859,I229205,I229279,);
not I_13317 (I229287,I458730);
nor I_13318 (I229304,I229231,I229287);
not I_13319 (I229321,I458745);
not I_13320 (I229338,I458736);
nand I_13321 (I229355,I229338,I458745);
nor I_13322 (I229372,I229287,I229355);
nor I_13323 (I229389,I229279,I229372);
DFFARX1 I_13324 (I229338,I2859,I229205,I229194,);
nor I_13325 (I229420,I458736,I458748);
nand I_13326 (I229437,I229420,I458727);
nor I_13327 (I229454,I229437,I229321);
nand I_13328 (I229179,I229454,I458730);
DFFARX1 I_13329 (I229437,I2859,I229205,I229191,);
nand I_13330 (I229499,I229321,I458736);
nor I_13331 (I229516,I229321,I458736);
nand I_13332 (I229185,I229304,I229516);
not I_13333 (I229547,I458733);
nor I_13334 (I229564,I229547,I229499);
DFFARX1 I_13335 (I229564,I2859,I229205,I229173,);
nor I_13336 (I229595,I229547,I458739);
and I_13337 (I229612,I229595,I458724);
or I_13338 (I229629,I229612,I458727);
DFFARX1 I_13339 (I229629,I2859,I229205,I229655,);
nor I_13340 (I229663,I229655,I229279);
nor I_13341 (I229182,I229231,I229663);
not I_13342 (I229694,I229655);
nor I_13343 (I229711,I229694,I229389);
DFFARX1 I_13344 (I229711,I2859,I229205,I229188,);
nand I_13345 (I229742,I229694,I229321);
nor I_13346 (I229176,I229547,I229742);
not I_13347 (I229800,I2866);
DFFARX1 I_13348 (I463348,I2859,I229800,I229826,);
not I_13349 (I229834,I229826);
DFFARX1 I_13350 (I463354,I2859,I229800,I229860,);
not I_13351 (I229868,I463348);
nand I_13352 (I229885,I229868,I463351);
not I_13353 (I229902,I229885);
nor I_13354 (I229919,I229902,I463369);
nor I_13355 (I229936,I229834,I229919);
DFFARX1 I_13356 (I229936,I2859,I229800,I229786,);
not I_13357 (I229967,I463369);
nand I_13358 (I229984,I229967,I229902);
and I_13359 (I230001,I229967,I463372);
nand I_13360 (I230018,I230001,I463351);
nor I_13361 (I229783,I230018,I229967);
and I_13362 (I229774,I229860,I230018);
not I_13363 (I230063,I230018);
nand I_13364 (I229777,I229860,I230063);
nor I_13365 (I229771,I229826,I230018);
not I_13366 (I230108,I463357);
nor I_13367 (I230125,I230108,I463372);
nand I_13368 (I230142,I230125,I229967);
nor I_13369 (I229780,I229885,I230142);
nor I_13370 (I230173,I230108,I463363);
and I_13371 (I230190,I230173,I463360);
or I_13372 (I230207,I230190,I463366);
DFFARX1 I_13373 (I230207,I2859,I229800,I230233,);
nor I_13374 (I230241,I230233,I229984);
DFFARX1 I_13375 (I230241,I2859,I229800,I229768,);
DFFARX1 I_13376 (I230233,I2859,I229800,I229792,);
not I_13377 (I230286,I230233);
nor I_13378 (I230303,I230286,I229860);
nor I_13379 (I230320,I230125,I230303);
DFFARX1 I_13380 (I230320,I2859,I229800,I229789,);
not I_13381 (I230378,I2866);
DFFARX1 I_13382 (I122419,I2859,I230378,I230404,);
not I_13383 (I230412,I230404);
DFFARX1 I_13384 (I122434,I2859,I230378,I230438,);
not I_13385 (I230446,I122437);
nand I_13386 (I230463,I230446,I122416);
not I_13387 (I230480,I230463);
nor I_13388 (I230497,I230480,I122440);
nor I_13389 (I230514,I230412,I230497);
DFFARX1 I_13390 (I230514,I2859,I230378,I230364,);
not I_13391 (I230545,I122440);
nand I_13392 (I230562,I230545,I230480);
and I_13393 (I230579,I230545,I122422);
nand I_13394 (I230596,I230579,I122413);
nor I_13395 (I230361,I230596,I230545);
and I_13396 (I230352,I230438,I230596);
not I_13397 (I230641,I230596);
nand I_13398 (I230355,I230438,I230641);
nor I_13399 (I230349,I230404,I230596);
not I_13400 (I230686,I122413);
nor I_13401 (I230703,I230686,I122422);
nand I_13402 (I230720,I230703,I230545);
nor I_13403 (I230358,I230463,I230720);
nor I_13404 (I230751,I230686,I122428);
and I_13405 (I230768,I230751,I122431);
or I_13406 (I230785,I230768,I122425);
DFFARX1 I_13407 (I230785,I2859,I230378,I230811,);
nor I_13408 (I230819,I230811,I230562);
DFFARX1 I_13409 (I230819,I2859,I230378,I230346,);
DFFARX1 I_13410 (I230811,I2859,I230378,I230370,);
not I_13411 (I230864,I230811);
nor I_13412 (I230881,I230864,I230438);
nor I_13413 (I230898,I230703,I230881);
DFFARX1 I_13414 (I230898,I2859,I230378,I230367,);
not I_13415 (I230956,I2866);
DFFARX1 I_13416 (I423557,I2859,I230956,I230982,);
not I_13417 (I230990,I230982);
DFFARX1 I_13418 (I423554,I2859,I230956,I231016,);
not I_13419 (I231024,I423551);
nand I_13420 (I231041,I231024,I423578);
not I_13421 (I231058,I231041);
nor I_13422 (I231075,I231058,I423566);
nor I_13423 (I231092,I230990,I231075);
DFFARX1 I_13424 (I231092,I2859,I230956,I230942,);
not I_13425 (I231123,I423566);
nand I_13426 (I231140,I231123,I231058);
and I_13427 (I231157,I231123,I423572);
nand I_13428 (I231174,I231157,I423563);
nor I_13429 (I230939,I231174,I231123);
and I_13430 (I230930,I231016,I231174);
not I_13431 (I231219,I231174);
nand I_13432 (I230933,I231016,I231219);
nor I_13433 (I230927,I230982,I231174);
not I_13434 (I231264,I423560);
nor I_13435 (I231281,I231264,I423572);
nand I_13436 (I231298,I231281,I231123);
nor I_13437 (I230936,I231041,I231298);
nor I_13438 (I231329,I231264,I423575);
and I_13439 (I231346,I231329,I423569);
or I_13440 (I231363,I231346,I423551);
DFFARX1 I_13441 (I231363,I2859,I230956,I231389,);
nor I_13442 (I231397,I231389,I231140);
DFFARX1 I_13443 (I231397,I2859,I230956,I230924,);
DFFARX1 I_13444 (I231389,I2859,I230956,I230948,);
not I_13445 (I231442,I231389);
nor I_13446 (I231459,I231442,I231016);
nor I_13447 (I231476,I231281,I231459);
DFFARX1 I_13448 (I231476,I2859,I230956,I230945,);
not I_13449 (I231534,I2866);
DFFARX1 I_13450 (I124527,I2859,I231534,I231560,);
not I_13451 (I231568,I231560);
DFFARX1 I_13452 (I124542,I2859,I231534,I231594,);
not I_13453 (I231602,I124545);
nand I_13454 (I231619,I231602,I124524);
not I_13455 (I231636,I231619);
nor I_13456 (I231653,I231636,I124548);
nor I_13457 (I231670,I231568,I231653);
DFFARX1 I_13458 (I231670,I2859,I231534,I231520,);
not I_13459 (I231701,I124548);
nand I_13460 (I231718,I231701,I231636);
and I_13461 (I231735,I231701,I124530);
nand I_13462 (I231752,I231735,I124521);
nor I_13463 (I231517,I231752,I231701);
and I_13464 (I231508,I231594,I231752);
not I_13465 (I231797,I231752);
nand I_13466 (I231511,I231594,I231797);
nor I_13467 (I231505,I231560,I231752);
not I_13468 (I231842,I124521);
nor I_13469 (I231859,I231842,I124530);
nand I_13470 (I231876,I231859,I231701);
nor I_13471 (I231514,I231619,I231876);
nor I_13472 (I231907,I231842,I124536);
and I_13473 (I231924,I231907,I124539);
or I_13474 (I231941,I231924,I124533);
DFFARX1 I_13475 (I231941,I2859,I231534,I231967,);
nor I_13476 (I231975,I231967,I231718);
DFFARX1 I_13477 (I231975,I2859,I231534,I231502,);
DFFARX1 I_13478 (I231967,I2859,I231534,I231526,);
not I_13479 (I232020,I231967);
nor I_13480 (I232037,I232020,I231594);
nor I_13481 (I232054,I231859,I232037);
DFFARX1 I_13482 (I232054,I2859,I231534,I231523,);
not I_13483 (I232112,I2866);
DFFARX1 I_13484 (I151404,I2859,I232112,I232138,);
not I_13485 (I232146,I232138);
DFFARX1 I_13486 (I151419,I2859,I232112,I232172,);
not I_13487 (I232180,I151422);
nand I_13488 (I232197,I232180,I151401);
not I_13489 (I232214,I232197);
nor I_13490 (I232231,I232214,I151425);
nor I_13491 (I232248,I232146,I232231);
DFFARX1 I_13492 (I232248,I2859,I232112,I232098,);
not I_13493 (I232279,I151425);
nand I_13494 (I232296,I232279,I232214);
and I_13495 (I232313,I232279,I151407);
nand I_13496 (I232330,I232313,I151398);
nor I_13497 (I232095,I232330,I232279);
and I_13498 (I232086,I232172,I232330);
not I_13499 (I232375,I232330);
nand I_13500 (I232089,I232172,I232375);
nor I_13501 (I232083,I232138,I232330);
not I_13502 (I232420,I151398);
nor I_13503 (I232437,I232420,I151407);
nand I_13504 (I232454,I232437,I232279);
nor I_13505 (I232092,I232197,I232454);
nor I_13506 (I232485,I232420,I151413);
and I_13507 (I232502,I232485,I151416);
or I_13508 (I232519,I232502,I151410);
DFFARX1 I_13509 (I232519,I2859,I232112,I232545,);
nor I_13510 (I232553,I232545,I232296);
DFFARX1 I_13511 (I232553,I2859,I232112,I232080,);
DFFARX1 I_13512 (I232545,I2859,I232112,I232104,);
not I_13513 (I232598,I232545);
nor I_13514 (I232615,I232598,I232172);
nor I_13515 (I232632,I232437,I232615);
DFFARX1 I_13516 (I232632,I2859,I232112,I232101,);
not I_13517 (I232690,I2866);
DFFARX1 I_13518 (I114514,I2859,I232690,I232716,);
not I_13519 (I232724,I232716);
DFFARX1 I_13520 (I114529,I2859,I232690,I232750,);
not I_13521 (I232758,I114532);
nand I_13522 (I232775,I232758,I114511);
not I_13523 (I232792,I232775);
nor I_13524 (I232809,I232792,I114535);
nor I_13525 (I232826,I232724,I232809);
DFFARX1 I_13526 (I232826,I2859,I232690,I232676,);
not I_13527 (I232857,I114535);
nand I_13528 (I232874,I232857,I232792);
and I_13529 (I232891,I232857,I114517);
nand I_13530 (I232908,I232891,I114508);
nor I_13531 (I232673,I232908,I232857);
and I_13532 (I232664,I232750,I232908);
not I_13533 (I232953,I232908);
nand I_13534 (I232667,I232750,I232953);
nor I_13535 (I232661,I232716,I232908);
not I_13536 (I232998,I114508);
nor I_13537 (I233015,I232998,I114517);
nand I_13538 (I233032,I233015,I232857);
nor I_13539 (I232670,I232775,I233032);
nor I_13540 (I233063,I232998,I114523);
and I_13541 (I233080,I233063,I114526);
or I_13542 (I233097,I233080,I114520);
DFFARX1 I_13543 (I233097,I2859,I232690,I233123,);
nor I_13544 (I233131,I233123,I232874);
DFFARX1 I_13545 (I233131,I2859,I232690,I232658,);
DFFARX1 I_13546 (I233123,I2859,I232690,I232682,);
not I_13547 (I233176,I233123);
nor I_13548 (I233193,I233176,I232750);
nor I_13549 (I233210,I233015,I233193);
DFFARX1 I_13550 (I233210,I2859,I232690,I232679,);
not I_13551 (I233268,I2866);
DFFARX1 I_13552 (I391257,I2859,I233268,I233294,);
not I_13553 (I233302,I233294);
DFFARX1 I_13554 (I391254,I2859,I233268,I233328,);
not I_13555 (I233336,I391251);
nand I_13556 (I233353,I233336,I391278);
not I_13557 (I233370,I233353);
nor I_13558 (I233387,I233370,I391266);
nor I_13559 (I233404,I233302,I233387);
DFFARX1 I_13560 (I233404,I2859,I233268,I233254,);
not I_13561 (I233435,I391266);
nand I_13562 (I233452,I233435,I233370);
and I_13563 (I233469,I233435,I391272);
nand I_13564 (I233486,I233469,I391263);
nor I_13565 (I233251,I233486,I233435);
and I_13566 (I233242,I233328,I233486);
not I_13567 (I233531,I233486);
nand I_13568 (I233245,I233328,I233531);
nor I_13569 (I233239,I233294,I233486);
not I_13570 (I233576,I391260);
nor I_13571 (I233593,I233576,I391272);
nand I_13572 (I233610,I233593,I233435);
nor I_13573 (I233248,I233353,I233610);
nor I_13574 (I233641,I233576,I391275);
and I_13575 (I233658,I233641,I391269);
or I_13576 (I233675,I233658,I391251);
DFFARX1 I_13577 (I233675,I2859,I233268,I233701,);
nor I_13578 (I233709,I233701,I233452);
DFFARX1 I_13579 (I233709,I2859,I233268,I233236,);
DFFARX1 I_13580 (I233701,I2859,I233268,I233260,);
not I_13581 (I233754,I233701);
nor I_13582 (I233771,I233754,I233328);
nor I_13583 (I233788,I233593,I233771);
DFFARX1 I_13584 (I233788,I2859,I233268,I233257,);
not I_13585 (I233846,I2866);
DFFARX1 I_13586 (I436560,I2859,I233846,I233872,);
not I_13587 (I233880,I233872);
DFFARX1 I_13588 (I436551,I2859,I233846,I233906,);
not I_13589 (I233914,I436545);
nand I_13590 (I233931,I233914,I436557);
not I_13591 (I233948,I233931);
nor I_13592 (I233965,I233948,I436548);
nor I_13593 (I233982,I233880,I233965);
DFFARX1 I_13594 (I233982,I2859,I233846,I233832,);
not I_13595 (I234013,I436548);
nand I_13596 (I234030,I234013,I233948);
and I_13597 (I234047,I234013,I436554);
nand I_13598 (I234064,I234047,I436539);
nor I_13599 (I233829,I234064,I234013);
and I_13600 (I233820,I233906,I234064);
not I_13601 (I234109,I234064);
nand I_13602 (I233823,I233906,I234109);
nor I_13603 (I233817,I233872,I234064);
not I_13604 (I234154,I436539);
nor I_13605 (I234171,I234154,I436554);
nand I_13606 (I234188,I234171,I234013);
nor I_13607 (I233826,I233931,I234188);
nor I_13608 (I234219,I234154,I436542);
and I_13609 (I234236,I234219,I436545);
or I_13610 (I234253,I234236,I436542);
DFFARX1 I_13611 (I234253,I2859,I233846,I234279,);
nor I_13612 (I234287,I234279,I234030);
DFFARX1 I_13613 (I234287,I2859,I233846,I233814,);
DFFARX1 I_13614 (I234279,I2859,I233846,I233838,);
not I_13615 (I234332,I234279);
nor I_13616 (I234349,I234332,I233906);
nor I_13617 (I234366,I234171,I234349);
DFFARX1 I_13618 (I234366,I2859,I233846,I233835,);
not I_13619 (I234424,I2866);
DFFARX1 I_13620 (I442170,I2859,I234424,I234450,);
not I_13621 (I234458,I234450);
DFFARX1 I_13622 (I442161,I2859,I234424,I234484,);
not I_13623 (I234492,I442155);
nand I_13624 (I234509,I234492,I442167);
not I_13625 (I234526,I234509);
nor I_13626 (I234543,I234526,I442158);
nor I_13627 (I234560,I234458,I234543);
DFFARX1 I_13628 (I234560,I2859,I234424,I234410,);
not I_13629 (I234591,I442158);
nand I_13630 (I234608,I234591,I234526);
and I_13631 (I234625,I234591,I442164);
nand I_13632 (I234642,I234625,I442149);
nor I_13633 (I234407,I234642,I234591);
and I_13634 (I234398,I234484,I234642);
not I_13635 (I234687,I234642);
nand I_13636 (I234401,I234484,I234687);
nor I_13637 (I234395,I234450,I234642);
not I_13638 (I234732,I442149);
nor I_13639 (I234749,I234732,I442164);
nand I_13640 (I234766,I234749,I234591);
nor I_13641 (I234404,I234509,I234766);
nor I_13642 (I234797,I234732,I442152);
and I_13643 (I234814,I234797,I442155);
or I_13644 (I234831,I234814,I442152);
DFFARX1 I_13645 (I234831,I2859,I234424,I234857,);
nor I_13646 (I234865,I234857,I234608);
DFFARX1 I_13647 (I234865,I2859,I234424,I234392,);
DFFARX1 I_13648 (I234857,I2859,I234424,I234416,);
not I_13649 (I234910,I234857);
nor I_13650 (I234927,I234910,I234484);
nor I_13651 (I234944,I234749,I234927);
DFFARX1 I_13652 (I234944,I2859,I234424,I234413,);
not I_13653 (I235002,I2866);
DFFARX1 I_13654 (I221441,I2859,I235002,I235028,);
not I_13655 (I235036,I235028);
DFFARX1 I_13656 (I221453,I2859,I235002,I235062,);
not I_13657 (I235070,I221459);
nand I_13658 (I235087,I235070,I221450);
not I_13659 (I235104,I235087);
nor I_13660 (I235121,I235104,I221456);
nor I_13661 (I235138,I235036,I235121);
DFFARX1 I_13662 (I235138,I2859,I235002,I234988,);
not I_13663 (I235169,I221456);
nand I_13664 (I235186,I235169,I235104);
and I_13665 (I235203,I235169,I221447);
nand I_13666 (I235220,I235203,I221438);
nor I_13667 (I234985,I235220,I235169);
and I_13668 (I234976,I235062,I235220);
not I_13669 (I235265,I235220);
nand I_13670 (I234979,I235062,I235265);
nor I_13671 (I234973,I235028,I235220);
not I_13672 (I235310,I221444);
nor I_13673 (I235327,I235310,I221447);
nand I_13674 (I235344,I235327,I235169);
nor I_13675 (I234982,I235087,I235344);
nor I_13676 (I235375,I235310,I221441);
and I_13677 (I235392,I235375,I221438);
or I_13678 (I235409,I235392,I221462);
DFFARX1 I_13679 (I235409,I2859,I235002,I235435,);
nor I_13680 (I235443,I235435,I235186);
DFFARX1 I_13681 (I235443,I2859,I235002,I234970,);
DFFARX1 I_13682 (I235435,I2859,I235002,I234994,);
not I_13683 (I235488,I235435);
nor I_13684 (I235505,I235488,I235062);
nor I_13685 (I235522,I235327,I235505);
DFFARX1 I_13686 (I235522,I2859,I235002,I234991,);
not I_13687 (I235580,I2866);
DFFARX1 I_13688 (I174343,I2859,I235580,I235606,);
not I_13689 (I235614,I235606);
DFFARX1 I_13690 (I174355,I2859,I235580,I235640,);
not I_13691 (I235648,I174331);
nand I_13692 (I235665,I235648,I174358);
not I_13693 (I235682,I235665);
nor I_13694 (I235699,I235682,I174346);
nor I_13695 (I235716,I235614,I235699);
DFFARX1 I_13696 (I235716,I2859,I235580,I235566,);
not I_13697 (I235747,I174346);
nand I_13698 (I235764,I235747,I235682);
and I_13699 (I235781,I235747,I174331);
nand I_13700 (I235798,I235781,I174334);
nor I_13701 (I235563,I235798,I235747);
and I_13702 (I235554,I235640,I235798);
not I_13703 (I235843,I235798);
nand I_13704 (I235557,I235640,I235843);
nor I_13705 (I235551,I235606,I235798);
not I_13706 (I235888,I174340);
nor I_13707 (I235905,I235888,I174331);
nand I_13708 (I235922,I235905,I235747);
nor I_13709 (I235560,I235665,I235922);
nor I_13710 (I235953,I235888,I174349);
and I_13711 (I235970,I235953,I174337);
or I_13712 (I235987,I235970,I174352);
DFFARX1 I_13713 (I235987,I2859,I235580,I236013,);
nor I_13714 (I236021,I236013,I235764);
DFFARX1 I_13715 (I236021,I2859,I235580,I235548,);
DFFARX1 I_13716 (I236013,I2859,I235580,I235572,);
not I_13717 (I236066,I236013);
nor I_13718 (I236083,I236066,I235640);
nor I_13719 (I236100,I235905,I236083);
DFFARX1 I_13720 (I236100,I2859,I235580,I235569,);
not I_13721 (I236158,I2866);
DFFARX1 I_13722 (I67943,I2859,I236158,I236184,);
not I_13723 (I236192,I236184);
DFFARX1 I_13724 (I67928,I2859,I236158,I236218,);
not I_13725 (I236226,I67946);
nand I_13726 (I236243,I236226,I67931);
not I_13727 (I236260,I236243);
nor I_13728 (I236277,I236260,I67928);
nor I_13729 (I236294,I236192,I236277);
DFFARX1 I_13730 (I236294,I2859,I236158,I236144,);
not I_13731 (I236325,I67928);
nand I_13732 (I236342,I236325,I236260);
and I_13733 (I236359,I236325,I67931);
nand I_13734 (I236376,I236359,I67952);
nor I_13735 (I236141,I236376,I236325);
and I_13736 (I236132,I236218,I236376);
not I_13737 (I236421,I236376);
nand I_13738 (I236135,I236218,I236421);
nor I_13739 (I236129,I236184,I236376);
not I_13740 (I236466,I67940);
nor I_13741 (I236483,I236466,I67931);
nand I_13742 (I236500,I236483,I236325);
nor I_13743 (I236138,I236243,I236500);
nor I_13744 (I236531,I236466,I67934);
and I_13745 (I236548,I236531,I67949);
or I_13746 (I236565,I236548,I67937);
DFFARX1 I_13747 (I236565,I2859,I236158,I236591,);
nor I_13748 (I236599,I236591,I236342);
DFFARX1 I_13749 (I236599,I2859,I236158,I236126,);
DFFARX1 I_13750 (I236591,I2859,I236158,I236150,);
not I_13751 (I236644,I236591);
nor I_13752 (I236661,I236644,I236218);
nor I_13753 (I236678,I236483,I236661);
DFFARX1 I_13754 (I236678,I2859,I236158,I236147,);
not I_13755 (I236736,I2866);
DFFARX1 I_13756 (I183047,I2859,I236736,I236762,);
not I_13757 (I236770,I236762);
DFFARX1 I_13758 (I183059,I2859,I236736,I236796,);
not I_13759 (I236804,I183035);
nand I_13760 (I236821,I236804,I183062);
not I_13761 (I236838,I236821);
nor I_13762 (I236855,I236838,I183050);
nor I_13763 (I236872,I236770,I236855);
DFFARX1 I_13764 (I236872,I2859,I236736,I236722,);
not I_13765 (I236903,I183050);
nand I_13766 (I236920,I236903,I236838);
and I_13767 (I236937,I236903,I183035);
nand I_13768 (I236954,I236937,I183038);
nor I_13769 (I236719,I236954,I236903);
and I_13770 (I236710,I236796,I236954);
not I_13771 (I236999,I236954);
nand I_13772 (I236713,I236796,I236999);
nor I_13773 (I236707,I236762,I236954);
not I_13774 (I237044,I183044);
nor I_13775 (I237061,I237044,I183035);
nand I_13776 (I237078,I237061,I236903);
nor I_13777 (I236716,I236821,I237078);
nor I_13778 (I237109,I237044,I183053);
and I_13779 (I237126,I237109,I183041);
or I_13780 (I237143,I237126,I183056);
DFFARX1 I_13781 (I237143,I2859,I236736,I237169,);
nor I_13782 (I237177,I237169,I236920);
DFFARX1 I_13783 (I237177,I2859,I236736,I236704,);
DFFARX1 I_13784 (I237169,I2859,I236736,I236728,);
not I_13785 (I237222,I237169);
nor I_13786 (I237239,I237222,I236796);
nor I_13787 (I237256,I237061,I237239);
DFFARX1 I_13788 (I237256,I2859,I236736,I236725,);
not I_13789 (I237314,I2866);
DFFARX1 I_13790 (I112933,I2859,I237314,I237340,);
not I_13791 (I237348,I237340);
DFFARX1 I_13792 (I112948,I2859,I237314,I237374,);
not I_13793 (I237382,I112951);
nand I_13794 (I237399,I237382,I112930);
not I_13795 (I237416,I237399);
nor I_13796 (I237433,I237416,I112954);
nor I_13797 (I237450,I237348,I237433);
DFFARX1 I_13798 (I237450,I2859,I237314,I237300,);
not I_13799 (I237481,I112954);
nand I_13800 (I237498,I237481,I237416);
and I_13801 (I237515,I237481,I112936);
nand I_13802 (I237532,I237515,I112927);
nor I_13803 (I237297,I237532,I237481);
and I_13804 (I237288,I237374,I237532);
not I_13805 (I237577,I237532);
nand I_13806 (I237291,I237374,I237577);
nor I_13807 (I237285,I237340,I237532);
not I_13808 (I237622,I112927);
nor I_13809 (I237639,I237622,I112936);
nand I_13810 (I237656,I237639,I237481);
nor I_13811 (I237294,I237399,I237656);
nor I_13812 (I237687,I237622,I112942);
and I_13813 (I237704,I237687,I112945);
or I_13814 (I237721,I237704,I112939);
DFFARX1 I_13815 (I237721,I2859,I237314,I237747,);
nor I_13816 (I237755,I237747,I237498);
DFFARX1 I_13817 (I237755,I2859,I237314,I237282,);
DFFARX1 I_13818 (I237747,I2859,I237314,I237306,);
not I_13819 (I237800,I237747);
nor I_13820 (I237817,I237800,I237374);
nor I_13821 (I237834,I237639,I237817);
DFFARX1 I_13822 (I237834,I2859,I237314,I237303,);
not I_13823 (I237892,I2866);
DFFARX1 I_13824 (I435438,I2859,I237892,I237918,);
not I_13825 (I237926,I237918);
DFFARX1 I_13826 (I435429,I2859,I237892,I237952,);
not I_13827 (I237960,I435423);
nand I_13828 (I237977,I237960,I435435);
not I_13829 (I237994,I237977);
nor I_13830 (I238011,I237994,I435426);
nor I_13831 (I238028,I237926,I238011);
DFFARX1 I_13832 (I238028,I2859,I237892,I237878,);
not I_13833 (I238059,I435426);
nand I_13834 (I238076,I238059,I237994);
and I_13835 (I238093,I238059,I435432);
nand I_13836 (I238110,I238093,I435417);
nor I_13837 (I237875,I238110,I238059);
and I_13838 (I237866,I237952,I238110);
not I_13839 (I238155,I238110);
nand I_13840 (I237869,I237952,I238155);
nor I_13841 (I237863,I237918,I238110);
not I_13842 (I238200,I435417);
nor I_13843 (I238217,I238200,I435432);
nand I_13844 (I238234,I238217,I238059);
nor I_13845 (I237872,I237977,I238234);
nor I_13846 (I238265,I238200,I435420);
and I_13847 (I238282,I238265,I435423);
or I_13848 (I238299,I238282,I435420);
DFFARX1 I_13849 (I238299,I2859,I237892,I238325,);
nor I_13850 (I238333,I238325,I238076);
DFFARX1 I_13851 (I238333,I2859,I237892,I237860,);
DFFARX1 I_13852 (I238325,I2859,I237892,I237884,);
not I_13853 (I238378,I238325);
nor I_13854 (I238395,I238378,I237952);
nor I_13855 (I238412,I238217,I238395);
DFFARX1 I_13856 (I238412,I2859,I237892,I237881,);
not I_13857 (I238470,I2866);
DFFARX1 I_13858 (I159309,I2859,I238470,I238496,);
not I_13859 (I238504,I238496);
DFFARX1 I_13860 (I159324,I2859,I238470,I238530,);
not I_13861 (I238538,I159327);
nand I_13862 (I238555,I238538,I159306);
not I_13863 (I238572,I238555);
nor I_13864 (I238589,I238572,I159330);
nor I_13865 (I238606,I238504,I238589);
DFFARX1 I_13866 (I238606,I2859,I238470,I238456,);
not I_13867 (I238637,I159330);
nand I_13868 (I238654,I238637,I238572);
and I_13869 (I238671,I238637,I159312);
nand I_13870 (I238688,I238671,I159303);
nor I_13871 (I238453,I238688,I238637);
and I_13872 (I238444,I238530,I238688);
not I_13873 (I238733,I238688);
nand I_13874 (I238447,I238530,I238733);
nor I_13875 (I238441,I238496,I238688);
not I_13876 (I238778,I159303);
nor I_13877 (I238795,I238778,I159312);
nand I_13878 (I238812,I238795,I238637);
nor I_13879 (I238450,I238555,I238812);
nor I_13880 (I238843,I238778,I159318);
and I_13881 (I238860,I238843,I159321);
or I_13882 (I238877,I238860,I159315);
DFFARX1 I_13883 (I238877,I2859,I238470,I238903,);
nor I_13884 (I238911,I238903,I238654);
DFFARX1 I_13885 (I238911,I2859,I238470,I238438,);
DFFARX1 I_13886 (I238903,I2859,I238470,I238462,);
not I_13887 (I238956,I238903);
nor I_13888 (I238973,I238956,I238530);
nor I_13889 (I238990,I238795,I238973);
DFFARX1 I_13890 (I238990,I2859,I238470,I238459,);
not I_13891 (I239048,I2866);
DFFARX1 I_13892 (I203719,I2859,I239048,I239074,);
not I_13893 (I239082,I239074);
DFFARX1 I_13894 (I203731,I2859,I239048,I239108,);
not I_13895 (I239116,I203707);
nand I_13896 (I239133,I239116,I203734);
not I_13897 (I239150,I239133);
nor I_13898 (I239167,I239150,I203722);
nor I_13899 (I239184,I239082,I239167);
DFFARX1 I_13900 (I239184,I2859,I239048,I239034,);
not I_13901 (I239215,I203722);
nand I_13902 (I239232,I239215,I239150);
and I_13903 (I239249,I239215,I203707);
nand I_13904 (I239266,I239249,I203710);
nor I_13905 (I239031,I239266,I239215);
and I_13906 (I239022,I239108,I239266);
not I_13907 (I239311,I239266);
nand I_13908 (I239025,I239108,I239311);
nor I_13909 (I239019,I239074,I239266);
not I_13910 (I239356,I203716);
nor I_13911 (I239373,I239356,I203707);
nand I_13912 (I239390,I239373,I239215);
nor I_13913 (I239028,I239133,I239390);
nor I_13914 (I239421,I239356,I203725);
and I_13915 (I239438,I239421,I203713);
or I_13916 (I239455,I239438,I203728);
DFFARX1 I_13917 (I239455,I2859,I239048,I239481,);
nor I_13918 (I239489,I239481,I239232);
DFFARX1 I_13919 (I239489,I2859,I239048,I239016,);
DFFARX1 I_13920 (I239481,I2859,I239048,I239040,);
not I_13921 (I239534,I239481);
nor I_13922 (I239551,I239534,I239108);
nor I_13923 (I239568,I239373,I239551);
DFFARX1 I_13924 (I239568,I2859,I239048,I239037,);
not I_13925 (I239626,I2866);
DFFARX1 I_13926 (I271384,I2859,I239626,I239652,);
not I_13927 (I239660,I239652);
DFFARX1 I_13928 (I271396,I2859,I239626,I239686,);
not I_13929 (I239694,I271387);
nand I_13930 (I239711,I239694,I271390);
not I_13931 (I239728,I239711);
nor I_13932 (I239745,I239728,I271393);
nor I_13933 (I239762,I239660,I239745);
DFFARX1 I_13934 (I239762,I2859,I239626,I239612,);
not I_13935 (I239793,I271393);
nand I_13936 (I239810,I239793,I239728);
and I_13937 (I239827,I239793,I271387);
nand I_13938 (I239844,I239827,I271399);
nor I_13939 (I239609,I239844,I239793);
and I_13940 (I239600,I239686,I239844);
not I_13941 (I239889,I239844);
nand I_13942 (I239603,I239686,I239889);
nor I_13943 (I239597,I239652,I239844);
not I_13944 (I239934,I271405);
nor I_13945 (I239951,I239934,I271387);
nand I_13946 (I239968,I239951,I239793);
nor I_13947 (I239606,I239711,I239968);
nor I_13948 (I239999,I239934,I271384);
and I_13949 (I240016,I239999,I271402);
or I_13950 (I240033,I240016,I271408);
DFFARX1 I_13951 (I240033,I2859,I239626,I240059,);
nor I_13952 (I240067,I240059,I239810);
DFFARX1 I_13953 (I240067,I2859,I239626,I239594,);
DFFARX1 I_13954 (I240059,I2859,I239626,I239618,);
not I_13955 (I240112,I240059);
nor I_13956 (I240129,I240112,I239686);
nor I_13957 (I240146,I239951,I240129);
DFFARX1 I_13958 (I240146,I2859,I239626,I239615,);
not I_13959 (I240204,I2866);
DFFARX1 I_13960 (I478954,I2859,I240204,I240230,);
not I_13961 (I240238,I240230);
DFFARX1 I_13962 (I478960,I2859,I240204,I240264,);
not I_13963 (I240272,I478954);
nand I_13964 (I240289,I240272,I478957);
not I_13965 (I240306,I240289);
nor I_13966 (I240323,I240306,I478975);
nor I_13967 (I240340,I240238,I240323);
DFFARX1 I_13968 (I240340,I2859,I240204,I240190,);
not I_13969 (I240371,I478975);
nand I_13970 (I240388,I240371,I240306);
and I_13971 (I240405,I240371,I478978);
nand I_13972 (I240422,I240405,I478957);
nor I_13973 (I240187,I240422,I240371);
and I_13974 (I240178,I240264,I240422);
not I_13975 (I240467,I240422);
nand I_13976 (I240181,I240264,I240467);
nor I_13977 (I240175,I240230,I240422);
not I_13978 (I240512,I478963);
nor I_13979 (I240529,I240512,I478978);
nand I_13980 (I240546,I240529,I240371);
nor I_13981 (I240184,I240289,I240546);
nor I_13982 (I240577,I240512,I478969);
and I_13983 (I240594,I240577,I478966);
or I_13984 (I240611,I240594,I478972);
DFFARX1 I_13985 (I240611,I2859,I240204,I240637,);
nor I_13986 (I240645,I240637,I240388);
DFFARX1 I_13987 (I240645,I2859,I240204,I240172,);
DFFARX1 I_13988 (I240637,I2859,I240204,I240196,);
not I_13989 (I240690,I240637);
nor I_13990 (I240707,I240690,I240264);
nor I_13991 (I240724,I240529,I240707);
DFFARX1 I_13992 (I240724,I2859,I240204,I240193,);
not I_13993 (I240782,I2866);
DFFARX1 I_13994 (I14143,I2859,I240782,I240808,);
not I_13995 (I240816,I240808);
DFFARX1 I_13996 (I14146,I2859,I240782,I240842,);
not I_13997 (I240850,I14140);
nand I_13998 (I240867,I240850,I14164);
not I_13999 (I240884,I240867);
nor I_14000 (I240901,I240884,I14143);
nor I_14001 (I240918,I240816,I240901);
DFFARX1 I_14002 (I240918,I2859,I240782,I240768,);
not I_14003 (I240949,I14143);
nand I_14004 (I240966,I240949,I240884);
and I_14005 (I240983,I240949,I14158);
nand I_14006 (I241000,I240983,I14152);
nor I_14007 (I240765,I241000,I240949);
and I_14008 (I240756,I240842,I241000);
not I_14009 (I241045,I241000);
nand I_14010 (I240759,I240842,I241045);
nor I_14011 (I240753,I240808,I241000);
not I_14012 (I241090,I14161);
nor I_14013 (I241107,I241090,I14158);
nand I_14014 (I241124,I241107,I240949);
nor I_14015 (I240762,I240867,I241124);
nor I_14016 (I241155,I241090,I14140);
and I_14017 (I241172,I241155,I14149);
or I_14018 (I241189,I241172,I14155);
DFFARX1 I_14019 (I241189,I2859,I240782,I241215,);
nor I_14020 (I241223,I241215,I240966);
DFFARX1 I_14021 (I241223,I2859,I240782,I240750,);
DFFARX1 I_14022 (I241215,I2859,I240782,I240774,);
not I_14023 (I241268,I241215);
nor I_14024 (I241285,I241268,I240842);
nor I_14025 (I241302,I241107,I241285);
DFFARX1 I_14026 (I241302,I2859,I240782,I240771,);
not I_14027 (I241360,I2866);
DFFARX1 I_14028 (I506444,I2859,I241360,I241386,);
not I_14029 (I241394,I241386);
DFFARX1 I_14030 (I506438,I2859,I241360,I241420,);
not I_14031 (I241428,I506447);
nand I_14032 (I241445,I241428,I506426);
not I_14033 (I241462,I241445);
nor I_14034 (I241479,I241462,I506435);
nor I_14035 (I241496,I241394,I241479);
DFFARX1 I_14036 (I241496,I2859,I241360,I241346,);
not I_14037 (I241527,I506435);
nand I_14038 (I241544,I241527,I241462);
and I_14039 (I241561,I241527,I506450);
nand I_14040 (I241578,I241561,I506429);
nor I_14041 (I241343,I241578,I241527);
and I_14042 (I241334,I241420,I241578);
not I_14043 (I241623,I241578);
nand I_14044 (I241337,I241420,I241623);
nor I_14045 (I241331,I241386,I241578);
not I_14046 (I241668,I506432);
nor I_14047 (I241685,I241668,I506450);
nand I_14048 (I241702,I241685,I241527);
nor I_14049 (I241340,I241445,I241702);
nor I_14050 (I241733,I241668,I506441);
and I_14051 (I241750,I241733,I506429);
or I_14052 (I241767,I241750,I506426);
DFFARX1 I_14053 (I241767,I2859,I241360,I241793,);
nor I_14054 (I241801,I241793,I241544);
DFFARX1 I_14055 (I241801,I2859,I241360,I241328,);
DFFARX1 I_14056 (I241793,I2859,I241360,I241352,);
not I_14057 (I241846,I241793);
nor I_14058 (I241863,I241846,I241420);
nor I_14059 (I241880,I241685,I241863);
DFFARX1 I_14060 (I241880,I2859,I241360,I241349,);
not I_14061 (I241938,I2866);
DFFARX1 I_14062 (I60214,I2859,I241938,I241964,);
not I_14063 (I241972,I241964);
DFFARX1 I_14064 (I60193,I2859,I241938,I241998,);
not I_14065 (I242006,I60193);
nand I_14066 (I242023,I242006,I60220);
not I_14067 (I242040,I242023);
nor I_14068 (I242057,I242040,I60196);
nor I_14069 (I242074,I241972,I242057);
DFFARX1 I_14070 (I242074,I2859,I241938,I241924,);
not I_14071 (I242105,I60196);
nand I_14072 (I242122,I242105,I242040);
and I_14073 (I242139,I242105,I60217);
nand I_14074 (I242156,I242139,I60199);
nor I_14075 (I241921,I242156,I242105);
and I_14076 (I241912,I241998,I242156);
not I_14077 (I242201,I242156);
nand I_14078 (I241915,I241998,I242201);
nor I_14079 (I241909,I241964,I242156);
not I_14080 (I242246,I60202);
nor I_14081 (I242263,I242246,I60217);
nand I_14082 (I242280,I242263,I242105);
nor I_14083 (I241918,I242023,I242280);
nor I_14084 (I242311,I242246,I60208);
and I_14085 (I242328,I242311,I60205);
or I_14086 (I242345,I242328,I60211);
DFFARX1 I_14087 (I242345,I2859,I241938,I242371,);
nor I_14088 (I242379,I242371,I242122);
DFFARX1 I_14089 (I242379,I2859,I241938,I241906,);
DFFARX1 I_14090 (I242371,I2859,I241938,I241930,);
not I_14091 (I242424,I242371);
nor I_14092 (I242441,I242424,I241998);
nor I_14093 (I242458,I242263,I242441);
DFFARX1 I_14094 (I242458,I2859,I241938,I241927,);
not I_14095 (I242516,I2866);
DFFARX1 I_14096 (I189575,I2859,I242516,I242542,);
not I_14097 (I242550,I242542);
DFFARX1 I_14098 (I189587,I2859,I242516,I242576,);
not I_14099 (I242584,I189563);
nand I_14100 (I242601,I242584,I189590);
not I_14101 (I242618,I242601);
nor I_14102 (I242635,I242618,I189578);
nor I_14103 (I242652,I242550,I242635);
DFFARX1 I_14104 (I242652,I2859,I242516,I242502,);
not I_14105 (I242683,I189578);
nand I_14106 (I242700,I242683,I242618);
and I_14107 (I242717,I242683,I189563);
nand I_14108 (I242734,I242717,I189566);
nor I_14109 (I242499,I242734,I242683);
and I_14110 (I242490,I242576,I242734);
not I_14111 (I242779,I242734);
nand I_14112 (I242493,I242576,I242779);
nor I_14113 (I242487,I242542,I242734);
not I_14114 (I242824,I189572);
nor I_14115 (I242841,I242824,I189563);
nand I_14116 (I242858,I242841,I242683);
nor I_14117 (I242496,I242601,I242858);
nor I_14118 (I242889,I242824,I189581);
and I_14119 (I242906,I242889,I189569);
or I_14120 (I242923,I242906,I189584);
DFFARX1 I_14121 (I242923,I2859,I242516,I242949,);
nor I_14122 (I242957,I242949,I242700);
DFFARX1 I_14123 (I242957,I2859,I242516,I242484,);
DFFARX1 I_14124 (I242949,I2859,I242516,I242508,);
not I_14125 (I243002,I242949);
nor I_14126 (I243019,I243002,I242576);
nor I_14127 (I243036,I242841,I243019);
DFFARX1 I_14128 (I243036,I2859,I242516,I242505,);
not I_14129 (I243094,I2866);
DFFARX1 I_14130 (I61404,I2859,I243094,I243120,);
not I_14131 (I243128,I243120);
DFFARX1 I_14132 (I61383,I2859,I243094,I243154,);
not I_14133 (I243162,I61383);
nand I_14134 (I243179,I243162,I61410);
not I_14135 (I243196,I243179);
nor I_14136 (I243213,I243196,I61386);
nor I_14137 (I243230,I243128,I243213);
DFFARX1 I_14138 (I243230,I2859,I243094,I243080,);
not I_14139 (I243261,I61386);
nand I_14140 (I243278,I243261,I243196);
and I_14141 (I243295,I243261,I61407);
nand I_14142 (I243312,I243295,I61389);
nor I_14143 (I243077,I243312,I243261);
and I_14144 (I243068,I243154,I243312);
not I_14145 (I243357,I243312);
nand I_14146 (I243071,I243154,I243357);
nor I_14147 (I243065,I243120,I243312);
not I_14148 (I243402,I61392);
nor I_14149 (I243419,I243402,I61407);
nand I_14150 (I243436,I243419,I243261);
nor I_14151 (I243074,I243179,I243436);
nor I_14152 (I243467,I243402,I61398);
and I_14153 (I243484,I243467,I61395);
or I_14154 (I243501,I243484,I61401);
DFFARX1 I_14155 (I243501,I2859,I243094,I243527,);
nor I_14156 (I243535,I243527,I243278);
DFFARX1 I_14157 (I243535,I2859,I243094,I243062,);
DFFARX1 I_14158 (I243527,I2859,I243094,I243086,);
not I_14159 (I243580,I243527);
nor I_14160 (I243597,I243580,I243154);
nor I_14161 (I243614,I243419,I243597);
DFFARX1 I_14162 (I243614,I2859,I243094,I243083,);
not I_14163 (I243672,I2866);
DFFARX1 I_14164 (I378337,I2859,I243672,I243698,);
not I_14165 (I243706,I243698);
DFFARX1 I_14166 (I378334,I2859,I243672,I243732,);
not I_14167 (I243740,I378331);
nand I_14168 (I243757,I243740,I378358);
not I_14169 (I243774,I243757);
nor I_14170 (I243791,I243774,I378346);
nor I_14171 (I243808,I243706,I243791);
DFFARX1 I_14172 (I243808,I2859,I243672,I243658,);
not I_14173 (I243839,I378346);
nand I_14174 (I243856,I243839,I243774);
and I_14175 (I243873,I243839,I378352);
nand I_14176 (I243890,I243873,I378343);
nor I_14177 (I243655,I243890,I243839);
and I_14178 (I243646,I243732,I243890);
not I_14179 (I243935,I243890);
nand I_14180 (I243649,I243732,I243935);
nor I_14181 (I243643,I243698,I243890);
not I_14182 (I243980,I378340);
nor I_14183 (I243997,I243980,I378352);
nand I_14184 (I244014,I243997,I243839);
nor I_14185 (I243652,I243757,I244014);
nor I_14186 (I244045,I243980,I378355);
and I_14187 (I244062,I244045,I378349);
or I_14188 (I244079,I244062,I378331);
DFFARX1 I_14189 (I244079,I2859,I243672,I244105,);
nor I_14190 (I244113,I244105,I243856);
DFFARX1 I_14191 (I244113,I2859,I243672,I243640,);
DFFARX1 I_14192 (I244105,I2859,I243672,I243664,);
not I_14193 (I244158,I244105);
nor I_14194 (I244175,I244158,I243732);
nor I_14195 (I244192,I243997,I244175);
DFFARX1 I_14196 (I244192,I2859,I243672,I243661,);
not I_14197 (I244250,I2866);
DFFARX1 I_14198 (I359535,I2859,I244250,I244276,);
not I_14199 (I244284,I244276);
DFFARX1 I_14200 (I359535,I2859,I244250,I244310,);
not I_14201 (I244318,I359532);
nand I_14202 (I244335,I244318,I359547);
not I_14203 (I244352,I244335);
nor I_14204 (I244369,I244352,I359541);
nor I_14205 (I244386,I244284,I244369);
DFFARX1 I_14206 (I244386,I2859,I244250,I244236,);
not I_14207 (I244417,I359541);
nand I_14208 (I244434,I244417,I244352);
and I_14209 (I244451,I244417,I359538);
nand I_14210 (I244468,I244451,I359529);
nor I_14211 (I244233,I244468,I244417);
and I_14212 (I244224,I244310,I244468);
not I_14213 (I244513,I244468);
nand I_14214 (I244227,I244310,I244513);
nor I_14215 (I244221,I244276,I244468);
not I_14216 (I244558,I359550);
nor I_14217 (I244575,I244558,I359538);
nand I_14218 (I244592,I244575,I244417);
nor I_14219 (I244230,I244335,I244592);
nor I_14220 (I244623,I244558,I359529);
and I_14221 (I244640,I244623,I359532);
or I_14222 (I244657,I244640,I359544);
DFFARX1 I_14223 (I244657,I2859,I244250,I244683,);
nor I_14224 (I244691,I244683,I244434);
DFFARX1 I_14225 (I244691,I2859,I244250,I244218,);
DFFARX1 I_14226 (I244683,I2859,I244250,I244242,);
not I_14227 (I244736,I244683);
nor I_14228 (I244753,I244736,I244310);
nor I_14229 (I244770,I244575,I244753);
DFFARX1 I_14230 (I244770,I2859,I244250,I244239,);
not I_14231 (I244828,I2866);
DFFARX1 I_14232 (I435999,I2859,I244828,I244854,);
not I_14233 (I244862,I244854);
DFFARX1 I_14234 (I435990,I2859,I244828,I244888,);
not I_14235 (I244896,I435984);
nand I_14236 (I244913,I244896,I435996);
not I_14237 (I244930,I244913);
nor I_14238 (I244947,I244930,I435987);
nor I_14239 (I244964,I244862,I244947);
DFFARX1 I_14240 (I244964,I2859,I244828,I244814,);
not I_14241 (I244995,I435987);
nand I_14242 (I245012,I244995,I244930);
and I_14243 (I245029,I244995,I435993);
nand I_14244 (I245046,I245029,I435978);
nor I_14245 (I244811,I245046,I244995);
and I_14246 (I244802,I244888,I245046);
not I_14247 (I245091,I245046);
nand I_14248 (I244805,I244888,I245091);
nor I_14249 (I244799,I244854,I245046);
not I_14250 (I245136,I435978);
nor I_14251 (I245153,I245136,I435993);
nand I_14252 (I245170,I245153,I244995);
nor I_14253 (I244808,I244913,I245170);
nor I_14254 (I245201,I245136,I435981);
and I_14255 (I245218,I245201,I435984);
or I_14256 (I245235,I245218,I435981);
DFFARX1 I_14257 (I245235,I2859,I244828,I245261,);
nor I_14258 (I245269,I245261,I245012);
DFFARX1 I_14259 (I245269,I2859,I244828,I244796,);
DFFARX1 I_14260 (I245261,I2859,I244828,I244820,);
not I_14261 (I245314,I245261);
nor I_14262 (I245331,I245314,I244888);
nor I_14263 (I245348,I245153,I245331);
DFFARX1 I_14264 (I245348,I2859,I244828,I244817,);
not I_14265 (I245406,I2866);
DFFARX1 I_14266 (I530374,I2859,I245406,I245432,);
not I_14267 (I245440,I245432);
DFFARX1 I_14268 (I530386,I2859,I245406,I245466,);
not I_14269 (I245474,I530377);
nand I_14270 (I245491,I245474,I530365);
not I_14271 (I245508,I245491);
nor I_14272 (I245525,I245508,I530362);
nor I_14273 (I245542,I245440,I245525);
DFFARX1 I_14274 (I245542,I2859,I245406,I245392,);
not I_14275 (I245573,I530362);
nand I_14276 (I245590,I245573,I245508);
and I_14277 (I245607,I245573,I530368);
nand I_14278 (I245624,I245607,I530365);
nor I_14279 (I245389,I245624,I245573);
and I_14280 (I245380,I245466,I245624);
not I_14281 (I245669,I245624);
nand I_14282 (I245383,I245466,I245669);
nor I_14283 (I245377,I245432,I245624);
not I_14284 (I245714,I530383);
nor I_14285 (I245731,I245714,I530368);
nand I_14286 (I245748,I245731,I245573);
nor I_14287 (I245386,I245491,I245748);
nor I_14288 (I245779,I245714,I530371);
and I_14289 (I245796,I245779,I530362);
or I_14290 (I245813,I245796,I530380);
DFFARX1 I_14291 (I245813,I2859,I245406,I245839,);
nor I_14292 (I245847,I245839,I245590);
DFFARX1 I_14293 (I245847,I2859,I245406,I245374,);
DFFARX1 I_14294 (I245839,I2859,I245406,I245398,);
not I_14295 (I245892,I245839);
nor I_14296 (I245909,I245892,I245466);
nor I_14297 (I245926,I245731,I245909);
DFFARX1 I_14298 (I245926,I2859,I245406,I245395,);
not I_14299 (I245984,I2866);
DFFARX1 I_14300 (I548450,I2859,I245984,I246010,);
not I_14301 (I246018,I246010);
DFFARX1 I_14302 (I548450,I2859,I245984,I246044,);
not I_14303 (I246052,I548474);
nand I_14304 (I246069,I246052,I548456);
not I_14305 (I246086,I246069);
nor I_14306 (I246103,I246086,I548471);
nor I_14307 (I246120,I246018,I246103);
DFFARX1 I_14308 (I246120,I2859,I245984,I245970,);
not I_14309 (I246151,I548471);
nand I_14310 (I246168,I246151,I246086);
and I_14311 (I246185,I246151,I548453);
nand I_14312 (I246202,I246185,I548462);
nor I_14313 (I245967,I246202,I246151);
and I_14314 (I245958,I246044,I246202);
not I_14315 (I246247,I246202);
nand I_14316 (I245961,I246044,I246247);
nor I_14317 (I245955,I246010,I246202);
not I_14318 (I246292,I548459);
nor I_14319 (I246309,I246292,I548453);
nand I_14320 (I246326,I246309,I246151);
nor I_14321 (I245964,I246069,I246326);
nor I_14322 (I246357,I246292,I548468);
and I_14323 (I246374,I246357,I548477);
or I_14324 (I246391,I246374,I548465);
DFFARX1 I_14325 (I246391,I2859,I245984,I246417,);
nor I_14326 (I246425,I246417,I246168);
DFFARX1 I_14327 (I246425,I2859,I245984,I245952,);
DFFARX1 I_14328 (I246417,I2859,I245984,I245976,);
not I_14329 (I246470,I246417);
nor I_14330 (I246487,I246470,I246044);
nor I_14331 (I246504,I246309,I246487);
DFFARX1 I_14332 (I246504,I2859,I245984,I245973,);
not I_14333 (I246562,I2866);
DFFARX1 I_14334 (I332658,I2859,I246562,I246588,);
not I_14335 (I246596,I246588);
DFFARX1 I_14336 (I332658,I2859,I246562,I246622,);
not I_14337 (I246630,I332655);
nand I_14338 (I246647,I246630,I332670);
not I_14339 (I246664,I246647);
nor I_14340 (I246681,I246664,I332664);
nor I_14341 (I246698,I246596,I246681);
DFFARX1 I_14342 (I246698,I2859,I246562,I246548,);
not I_14343 (I246729,I332664);
nand I_14344 (I246746,I246729,I246664);
and I_14345 (I246763,I246729,I332661);
nand I_14346 (I246780,I246763,I332652);
nor I_14347 (I246545,I246780,I246729);
and I_14348 (I246536,I246622,I246780);
not I_14349 (I246825,I246780);
nand I_14350 (I246539,I246622,I246825);
nor I_14351 (I246533,I246588,I246780);
not I_14352 (I246870,I332673);
nor I_14353 (I246887,I246870,I332661);
nand I_14354 (I246904,I246887,I246729);
nor I_14355 (I246542,I246647,I246904);
nor I_14356 (I246935,I246870,I332652);
and I_14357 (I246952,I246935,I332655);
or I_14358 (I246969,I246952,I332667);
DFFARX1 I_14359 (I246969,I2859,I246562,I246995,);
nor I_14360 (I247003,I246995,I246746);
DFFARX1 I_14361 (I247003,I2859,I246562,I246530,);
DFFARX1 I_14362 (I246995,I2859,I246562,I246554,);
not I_14363 (I247048,I246995);
nor I_14364 (I247065,I247048,I246622);
nor I_14365 (I247082,I246887,I247065);
DFFARX1 I_14366 (I247082,I2859,I246562,I246551,);
not I_14367 (I247140,I2866);
DFFARX1 I_14368 (I310688,I2859,I247140,I247166,);
not I_14369 (I247174,I247166);
DFFARX1 I_14370 (I310700,I2859,I247140,I247200,);
not I_14371 (I247208,I310691);
nand I_14372 (I247225,I247208,I310694);
not I_14373 (I247242,I247225);
nor I_14374 (I247259,I247242,I310697);
nor I_14375 (I247276,I247174,I247259);
DFFARX1 I_14376 (I247276,I2859,I247140,I247126,);
not I_14377 (I247307,I310697);
nand I_14378 (I247324,I247307,I247242);
and I_14379 (I247341,I247307,I310691);
nand I_14380 (I247358,I247341,I310703);
nor I_14381 (I247123,I247358,I247307);
and I_14382 (I247114,I247200,I247358);
not I_14383 (I247403,I247358);
nand I_14384 (I247117,I247200,I247403);
nor I_14385 (I247111,I247166,I247358);
not I_14386 (I247448,I310709);
nor I_14387 (I247465,I247448,I310691);
nand I_14388 (I247482,I247465,I247307);
nor I_14389 (I247120,I247225,I247482);
nor I_14390 (I247513,I247448,I310688);
and I_14391 (I247530,I247513,I310706);
or I_14392 (I247547,I247530,I310712);
DFFARX1 I_14393 (I247547,I2859,I247140,I247573,);
nor I_14394 (I247581,I247573,I247324);
DFFARX1 I_14395 (I247581,I2859,I247140,I247108,);
DFFARX1 I_14396 (I247573,I2859,I247140,I247132,);
not I_14397 (I247626,I247573);
nor I_14398 (I247643,I247626,I247200);
nor I_14399 (I247660,I247465,I247643);
DFFARX1 I_14400 (I247660,I2859,I247140,I247129,);
not I_14401 (I247718,I2866);
DFFARX1 I_14402 (I285834,I2859,I247718,I247744,);
not I_14403 (I247752,I247744);
DFFARX1 I_14404 (I285846,I2859,I247718,I247778,);
not I_14405 (I247786,I285837);
nand I_14406 (I247803,I247786,I285840);
not I_14407 (I247820,I247803);
nor I_14408 (I247837,I247820,I285843);
nor I_14409 (I247854,I247752,I247837);
DFFARX1 I_14410 (I247854,I2859,I247718,I247704,);
not I_14411 (I247885,I285843);
nand I_14412 (I247902,I247885,I247820);
and I_14413 (I247919,I247885,I285837);
nand I_14414 (I247936,I247919,I285849);
nor I_14415 (I247701,I247936,I247885);
and I_14416 (I247692,I247778,I247936);
not I_14417 (I247981,I247936);
nand I_14418 (I247695,I247778,I247981);
nor I_14419 (I247689,I247744,I247936);
not I_14420 (I248026,I285855);
nor I_14421 (I248043,I248026,I285837);
nand I_14422 (I248060,I248043,I247885);
nor I_14423 (I247698,I247803,I248060);
nor I_14424 (I248091,I248026,I285834);
and I_14425 (I248108,I248091,I285852);
or I_14426 (I248125,I248108,I285858);
DFFARX1 I_14427 (I248125,I2859,I247718,I248151,);
nor I_14428 (I248159,I248151,I247902);
DFFARX1 I_14429 (I248159,I2859,I247718,I247686,);
DFFARX1 I_14430 (I248151,I2859,I247718,I247710,);
not I_14431 (I248204,I248151);
nor I_14432 (I248221,I248204,I247778);
nor I_14433 (I248238,I248043,I248221);
DFFARX1 I_14434 (I248238,I2859,I247718,I247707,);
not I_14435 (I248296,I2866);
DFFARX1 I_14436 (I564515,I2859,I248296,I248322,);
not I_14437 (I248330,I248322);
DFFARX1 I_14438 (I564515,I2859,I248296,I248356,);
not I_14439 (I248364,I564539);
nand I_14440 (I248381,I248364,I564521);
not I_14441 (I248398,I248381);
nor I_14442 (I248415,I248398,I564536);
nor I_14443 (I248432,I248330,I248415);
DFFARX1 I_14444 (I248432,I2859,I248296,I248282,);
not I_14445 (I248463,I564536);
nand I_14446 (I248480,I248463,I248398);
and I_14447 (I248497,I248463,I564518);
nand I_14448 (I248514,I248497,I564527);
nor I_14449 (I248279,I248514,I248463);
and I_14450 (I248270,I248356,I248514);
not I_14451 (I248559,I248514);
nand I_14452 (I248273,I248356,I248559);
nor I_14453 (I248267,I248322,I248514);
not I_14454 (I248604,I564524);
nor I_14455 (I248621,I248604,I564518);
nand I_14456 (I248638,I248621,I248463);
nor I_14457 (I248276,I248381,I248638);
nor I_14458 (I248669,I248604,I564533);
and I_14459 (I248686,I248669,I564542);
or I_14460 (I248703,I248686,I564530);
DFFARX1 I_14461 (I248703,I2859,I248296,I248729,);
nor I_14462 (I248737,I248729,I248480);
DFFARX1 I_14463 (I248737,I2859,I248296,I248264,);
DFFARX1 I_14464 (I248729,I2859,I248296,I248288,);
not I_14465 (I248782,I248729);
nor I_14466 (I248799,I248782,I248356);
nor I_14467 (I248816,I248621,I248799);
DFFARX1 I_14468 (I248816,I2859,I248296,I248285,);
not I_14469 (I248874,I2866);
DFFARX1 I_14470 (I419035,I2859,I248874,I248900,);
not I_14471 (I248908,I248900);
DFFARX1 I_14472 (I419032,I2859,I248874,I248934,);
not I_14473 (I248942,I419029);
nand I_14474 (I248959,I248942,I419056);
not I_14475 (I248976,I248959);
nor I_14476 (I248993,I248976,I419044);
nor I_14477 (I249010,I248908,I248993);
DFFARX1 I_14478 (I249010,I2859,I248874,I248860,);
not I_14479 (I249041,I419044);
nand I_14480 (I249058,I249041,I248976);
and I_14481 (I249075,I249041,I419050);
nand I_14482 (I249092,I249075,I419041);
nor I_14483 (I248857,I249092,I249041);
and I_14484 (I248848,I248934,I249092);
not I_14485 (I249137,I249092);
nand I_14486 (I248851,I248934,I249137);
nor I_14487 (I248845,I248900,I249092);
not I_14488 (I249182,I419038);
nor I_14489 (I249199,I249182,I419050);
nand I_14490 (I249216,I249199,I249041);
nor I_14491 (I248854,I248959,I249216);
nor I_14492 (I249247,I249182,I419053);
and I_14493 (I249264,I249247,I419047);
or I_14494 (I249281,I249264,I419029);
DFFARX1 I_14495 (I249281,I2859,I248874,I249307,);
nor I_14496 (I249315,I249307,I249058);
DFFARX1 I_14497 (I249315,I2859,I248874,I248842,);
DFFARX1 I_14498 (I249307,I2859,I248874,I248866,);
not I_14499 (I249360,I249307);
nor I_14500 (I249377,I249360,I248934);
nor I_14501 (I249394,I249199,I249377);
DFFARX1 I_14502 (I249394,I2859,I248874,I248863,);
not I_14503 (I249452,I2866);
DFFARX1 I_14504 (I342144,I2859,I249452,I249478,);
not I_14505 (I249486,I249478);
DFFARX1 I_14506 (I342144,I2859,I249452,I249512,);
not I_14507 (I249520,I342141);
nand I_14508 (I249537,I249520,I342156);
not I_14509 (I249554,I249537);
nor I_14510 (I249571,I249554,I342150);
nor I_14511 (I249588,I249486,I249571);
DFFARX1 I_14512 (I249588,I2859,I249452,I249438,);
not I_14513 (I249619,I342150);
nand I_14514 (I249636,I249619,I249554);
and I_14515 (I249653,I249619,I342147);
nand I_14516 (I249670,I249653,I342138);
nor I_14517 (I249435,I249670,I249619);
and I_14518 (I249426,I249512,I249670);
not I_14519 (I249715,I249670);
nand I_14520 (I249429,I249512,I249715);
nor I_14521 (I249423,I249478,I249670);
not I_14522 (I249760,I342159);
nor I_14523 (I249777,I249760,I342147);
nand I_14524 (I249794,I249777,I249619);
nor I_14525 (I249432,I249537,I249794);
nor I_14526 (I249825,I249760,I342138);
and I_14527 (I249842,I249825,I342141);
or I_14528 (I249859,I249842,I342153);
DFFARX1 I_14529 (I249859,I2859,I249452,I249885,);
nor I_14530 (I249893,I249885,I249636);
DFFARX1 I_14531 (I249893,I2859,I249452,I249420,);
DFFARX1 I_14532 (I249885,I2859,I249452,I249444,);
not I_14533 (I249938,I249885);
nor I_14534 (I249955,I249938,I249512);
nor I_14535 (I249972,I249777,I249955);
DFFARX1 I_14536 (I249972,I2859,I249452,I249441,);
not I_14537 (I250030,I2866);
DFFARX1 I_14538 (I16778,I2859,I250030,I250056,);
not I_14539 (I250064,I250056);
DFFARX1 I_14540 (I16781,I2859,I250030,I250090,);
not I_14541 (I250098,I16775);
nand I_14542 (I250115,I250098,I16799);
not I_14543 (I250132,I250115);
nor I_14544 (I250149,I250132,I16778);
nor I_14545 (I250166,I250064,I250149);
DFFARX1 I_14546 (I250166,I2859,I250030,I250016,);
not I_14547 (I250197,I16778);
nand I_14548 (I250214,I250197,I250132);
and I_14549 (I250231,I250197,I16793);
nand I_14550 (I250248,I250231,I16787);
nor I_14551 (I250013,I250248,I250197);
and I_14552 (I250004,I250090,I250248);
not I_14553 (I250293,I250248);
nand I_14554 (I250007,I250090,I250293);
nor I_14555 (I250001,I250056,I250248);
not I_14556 (I250338,I16796);
nor I_14557 (I250355,I250338,I16793);
nand I_14558 (I250372,I250355,I250197);
nor I_14559 (I250010,I250115,I250372);
nor I_14560 (I250403,I250338,I16775);
and I_14561 (I250420,I250403,I16784);
or I_14562 (I250437,I250420,I16790);
DFFARX1 I_14563 (I250437,I2859,I250030,I250463,);
nor I_14564 (I250471,I250463,I250214);
DFFARX1 I_14565 (I250471,I2859,I250030,I249998,);
DFFARX1 I_14566 (I250463,I2859,I250030,I250022,);
not I_14567 (I250516,I250463);
nor I_14568 (I250533,I250516,I250090);
nor I_14569 (I250550,I250355,I250533);
DFFARX1 I_14570 (I250550,I2859,I250030,I250019,);
not I_14571 (I250608,I2866);
DFFARX1 I_14572 (I19940,I2859,I250608,I250634,);
not I_14573 (I250642,I250634);
DFFARX1 I_14574 (I19943,I2859,I250608,I250668,);
not I_14575 (I250676,I19937);
nand I_14576 (I250693,I250676,I19961);
not I_14577 (I250710,I250693);
nor I_14578 (I250727,I250710,I19940);
nor I_14579 (I250744,I250642,I250727);
DFFARX1 I_14580 (I250744,I2859,I250608,I250594,);
not I_14581 (I250775,I19940);
nand I_14582 (I250792,I250775,I250710);
and I_14583 (I250809,I250775,I19955);
nand I_14584 (I250826,I250809,I19949);
nor I_14585 (I250591,I250826,I250775);
and I_14586 (I250582,I250668,I250826);
not I_14587 (I250871,I250826);
nand I_14588 (I250585,I250668,I250871);
nor I_14589 (I250579,I250634,I250826);
not I_14590 (I250916,I19958);
nor I_14591 (I250933,I250916,I19955);
nand I_14592 (I250950,I250933,I250775);
nor I_14593 (I250588,I250693,I250950);
nor I_14594 (I250981,I250916,I19937);
and I_14595 (I250998,I250981,I19946);
or I_14596 (I251015,I250998,I19952);
DFFARX1 I_14597 (I251015,I2859,I250608,I251041,);
nor I_14598 (I251049,I251041,I250792);
DFFARX1 I_14599 (I251049,I2859,I250608,I250576,);
DFFARX1 I_14600 (I251041,I2859,I250608,I250600,);
not I_14601 (I251094,I251041);
nor I_14602 (I251111,I251094,I250668);
nor I_14603 (I251128,I250933,I251111);
DFFARX1 I_14604 (I251128,I2859,I250608,I250597,);
not I_14605 (I251186,I2866);
DFFARX1 I_14606 (I355319,I2859,I251186,I251212,);
not I_14607 (I251220,I251212);
DFFARX1 I_14608 (I355319,I2859,I251186,I251246,);
not I_14609 (I251254,I355316);
nand I_14610 (I251271,I251254,I355331);
not I_14611 (I251288,I251271);
nor I_14612 (I251305,I251288,I355325);
nor I_14613 (I251322,I251220,I251305);
DFFARX1 I_14614 (I251322,I2859,I251186,I251172,);
not I_14615 (I251353,I355325);
nand I_14616 (I251370,I251353,I251288);
and I_14617 (I251387,I251353,I355322);
nand I_14618 (I251404,I251387,I355313);
nor I_14619 (I251169,I251404,I251353);
and I_14620 (I251160,I251246,I251404);
not I_14621 (I251449,I251404);
nand I_14622 (I251163,I251246,I251449);
nor I_14623 (I251157,I251212,I251404);
not I_14624 (I251494,I355334);
nor I_14625 (I251511,I251494,I355322);
nand I_14626 (I251528,I251511,I251353);
nor I_14627 (I251166,I251271,I251528);
nor I_14628 (I251559,I251494,I355313);
and I_14629 (I251576,I251559,I355316);
or I_14630 (I251593,I251576,I355328);
DFFARX1 I_14631 (I251593,I2859,I251186,I251619,);
nor I_14632 (I251627,I251619,I251370);
DFFARX1 I_14633 (I251627,I2859,I251186,I251154,);
DFFARX1 I_14634 (I251619,I2859,I251186,I251178,);
not I_14635 (I251672,I251619);
nor I_14636 (I251689,I251672,I251246);
nor I_14637 (I251706,I251511,I251689);
DFFARX1 I_14638 (I251706,I2859,I251186,I251175,);
not I_14639 (I251764,I2866);
DFFARX1 I_14640 (I180327,I2859,I251764,I251790,);
not I_14641 (I251798,I251790);
DFFARX1 I_14642 (I180339,I2859,I251764,I251824,);
not I_14643 (I251832,I180315);
nand I_14644 (I251849,I251832,I180342);
not I_14645 (I251866,I251849);
nor I_14646 (I251883,I251866,I180330);
nor I_14647 (I251900,I251798,I251883);
DFFARX1 I_14648 (I251900,I2859,I251764,I251750,);
not I_14649 (I251931,I180330);
nand I_14650 (I251948,I251931,I251866);
and I_14651 (I251965,I251931,I180315);
nand I_14652 (I251982,I251965,I180318);
nor I_14653 (I251747,I251982,I251931);
and I_14654 (I251738,I251824,I251982);
not I_14655 (I252027,I251982);
nand I_14656 (I251741,I251824,I252027);
nor I_14657 (I251735,I251790,I251982);
not I_14658 (I252072,I180324);
nor I_14659 (I252089,I252072,I180315);
nand I_14660 (I252106,I252089,I251931);
nor I_14661 (I251744,I251849,I252106);
nor I_14662 (I252137,I252072,I180333);
and I_14663 (I252154,I252137,I180321);
or I_14664 (I252171,I252154,I180336);
DFFARX1 I_14665 (I252171,I2859,I251764,I252197,);
nor I_14666 (I252205,I252197,I251948);
DFFARX1 I_14667 (I252205,I2859,I251764,I251732,);
DFFARX1 I_14668 (I252197,I2859,I251764,I251756,);
not I_14669 (I252250,I252197);
nor I_14670 (I252267,I252250,I251824);
nor I_14671 (I252284,I252089,I252267);
DFFARX1 I_14672 (I252284,I2859,I251764,I251753,);
not I_14673 (I252342,I2866);
DFFARX1 I_14674 (I152458,I2859,I252342,I252368,);
not I_14675 (I252376,I252368);
DFFARX1 I_14676 (I152473,I2859,I252342,I252402,);
not I_14677 (I252410,I152476);
nand I_14678 (I252427,I252410,I152455);
not I_14679 (I252444,I252427);
nor I_14680 (I252461,I252444,I152479);
nor I_14681 (I252478,I252376,I252461);
DFFARX1 I_14682 (I252478,I2859,I252342,I252328,);
not I_14683 (I252509,I152479);
nand I_14684 (I252526,I252509,I252444);
and I_14685 (I252543,I252509,I152461);
nand I_14686 (I252560,I252543,I152452);
nor I_14687 (I252325,I252560,I252509);
and I_14688 (I252316,I252402,I252560);
not I_14689 (I252605,I252560);
nand I_14690 (I252319,I252402,I252605);
nor I_14691 (I252313,I252368,I252560);
not I_14692 (I252650,I152452);
nor I_14693 (I252667,I252650,I152461);
nand I_14694 (I252684,I252667,I252509);
nor I_14695 (I252322,I252427,I252684);
nor I_14696 (I252715,I252650,I152467);
and I_14697 (I252732,I252715,I152470);
or I_14698 (I252749,I252732,I152464);
DFFARX1 I_14699 (I252749,I2859,I252342,I252775,);
nor I_14700 (I252783,I252775,I252526);
DFFARX1 I_14701 (I252783,I2859,I252342,I252310,);
DFFARX1 I_14702 (I252775,I2859,I252342,I252334,);
not I_14703 (I252828,I252775);
nor I_14704 (I252845,I252828,I252402);
nor I_14705 (I252862,I252667,I252845);
DFFARX1 I_14706 (I252862,I2859,I252342,I252331,);
not I_14707 (I252920,I2866);
DFFARX1 I_14708 (I162998,I2859,I252920,I252946,);
not I_14709 (I252954,I252946);
DFFARX1 I_14710 (I163013,I2859,I252920,I252980,);
not I_14711 (I252988,I163016);
nand I_14712 (I253005,I252988,I162995);
not I_14713 (I253022,I253005);
nor I_14714 (I253039,I253022,I163019);
nor I_14715 (I253056,I252954,I253039);
DFFARX1 I_14716 (I253056,I2859,I252920,I252906,);
not I_14717 (I253087,I163019);
nand I_14718 (I253104,I253087,I253022);
and I_14719 (I253121,I253087,I163001);
nand I_14720 (I253138,I253121,I162992);
nor I_14721 (I252903,I253138,I253087);
and I_14722 (I252894,I252980,I253138);
not I_14723 (I253183,I253138);
nand I_14724 (I252897,I252980,I253183);
nor I_14725 (I252891,I252946,I253138);
not I_14726 (I253228,I162992);
nor I_14727 (I253245,I253228,I163001);
nand I_14728 (I253262,I253245,I253087);
nor I_14729 (I252900,I253005,I253262);
nor I_14730 (I253293,I253228,I163007);
and I_14731 (I253310,I253293,I163010);
or I_14732 (I253327,I253310,I163004);
DFFARX1 I_14733 (I253327,I2859,I252920,I253353,);
nor I_14734 (I253361,I253353,I253104);
DFFARX1 I_14735 (I253361,I2859,I252920,I252888,);
DFFARX1 I_14736 (I253353,I2859,I252920,I252912,);
not I_14737 (I253406,I253353);
nor I_14738 (I253423,I253406,I252980);
nor I_14739 (I253440,I253245,I253423);
DFFARX1 I_14740 (I253440,I2859,I252920,I252909,);
not I_14741 (I253498,I2866);
DFFARX1 I_14742 (I293348,I2859,I253498,I253524,);
not I_14743 (I253532,I253524);
DFFARX1 I_14744 (I293360,I2859,I253498,I253558,);
not I_14745 (I253566,I293351);
nand I_14746 (I253583,I253566,I293354);
not I_14747 (I253600,I253583);
nor I_14748 (I253617,I253600,I293357);
nor I_14749 (I253634,I253532,I253617);
DFFARX1 I_14750 (I253634,I2859,I253498,I253484,);
not I_14751 (I253665,I293357);
nand I_14752 (I253682,I253665,I253600);
and I_14753 (I253699,I253665,I293351);
nand I_14754 (I253716,I253699,I293363);
nor I_14755 (I253481,I253716,I253665);
and I_14756 (I253472,I253558,I253716);
not I_14757 (I253761,I253716);
nand I_14758 (I253475,I253558,I253761);
nor I_14759 (I253469,I253524,I253716);
not I_14760 (I253806,I293369);
nor I_14761 (I253823,I253806,I293351);
nand I_14762 (I253840,I253823,I253665);
nor I_14763 (I253478,I253583,I253840);
nor I_14764 (I253871,I253806,I293348);
and I_14765 (I253888,I253871,I293366);
or I_14766 (I253905,I253888,I293372);
DFFARX1 I_14767 (I253905,I2859,I253498,I253931,);
nor I_14768 (I253939,I253931,I253682);
DFFARX1 I_14769 (I253939,I2859,I253498,I253466,);
DFFARX1 I_14770 (I253931,I2859,I253498,I253490,);
not I_14771 (I253984,I253931);
nor I_14772 (I254001,I253984,I253558);
nor I_14773 (I254018,I253823,I254001);
DFFARX1 I_14774 (I254018,I2859,I253498,I253487,);
not I_14775 (I254076,I2866);
DFFARX1 I_14776 (I420327,I2859,I254076,I254102,);
not I_14777 (I254110,I254102);
DFFARX1 I_14778 (I420324,I2859,I254076,I254136,);
not I_14779 (I254144,I420321);
nand I_14780 (I254161,I254144,I420348);
not I_14781 (I254178,I254161);
nor I_14782 (I254195,I254178,I420336);
nor I_14783 (I254212,I254110,I254195);
DFFARX1 I_14784 (I254212,I2859,I254076,I254062,);
not I_14785 (I254243,I420336);
nand I_14786 (I254260,I254243,I254178);
and I_14787 (I254277,I254243,I420342);
nand I_14788 (I254294,I254277,I420333);
nor I_14789 (I254059,I254294,I254243);
and I_14790 (I254050,I254136,I254294);
not I_14791 (I254339,I254294);
nand I_14792 (I254053,I254136,I254339);
nor I_14793 (I254047,I254102,I254294);
not I_14794 (I254384,I420330);
nor I_14795 (I254401,I254384,I420342);
nand I_14796 (I254418,I254401,I254243);
nor I_14797 (I254056,I254161,I254418);
nor I_14798 (I254449,I254384,I420345);
and I_14799 (I254466,I254449,I420339);
or I_14800 (I254483,I254466,I420321);
DFFARX1 I_14801 (I254483,I2859,I254076,I254509,);
nor I_14802 (I254517,I254509,I254260);
DFFARX1 I_14803 (I254517,I2859,I254076,I254044,);
DFFARX1 I_14804 (I254509,I2859,I254076,I254068,);
not I_14805 (I254562,I254509);
nor I_14806 (I254579,I254562,I254136);
nor I_14807 (I254596,I254401,I254579);
DFFARX1 I_14808 (I254596,I2859,I254076,I254065,);
not I_14809 (I254654,I2866);
DFFARX1 I_14810 (I455834,I2859,I254654,I254680,);
not I_14811 (I254688,I254680);
DFFARX1 I_14812 (I455840,I2859,I254654,I254714,);
not I_14813 (I254722,I455834);
nand I_14814 (I254739,I254722,I455837);
not I_14815 (I254756,I254739);
nor I_14816 (I254773,I254756,I455855);
nor I_14817 (I254790,I254688,I254773);
DFFARX1 I_14818 (I254790,I2859,I254654,I254640,);
not I_14819 (I254821,I455855);
nand I_14820 (I254838,I254821,I254756);
and I_14821 (I254855,I254821,I455858);
nand I_14822 (I254872,I254855,I455837);
nor I_14823 (I254637,I254872,I254821);
and I_14824 (I254628,I254714,I254872);
not I_14825 (I254917,I254872);
nand I_14826 (I254631,I254714,I254917);
nor I_14827 (I254625,I254680,I254872);
not I_14828 (I254962,I455843);
nor I_14829 (I254979,I254962,I455858);
nand I_14830 (I254996,I254979,I254821);
nor I_14831 (I254634,I254739,I254996);
nor I_14832 (I255027,I254962,I455849);
and I_14833 (I255044,I255027,I455846);
or I_14834 (I255061,I255044,I455852);
DFFARX1 I_14835 (I255061,I2859,I254654,I255087,);
nor I_14836 (I255095,I255087,I254838);
DFFARX1 I_14837 (I255095,I2859,I254654,I254622,);
DFFARX1 I_14838 (I255087,I2859,I254654,I254646,);
not I_14839 (I255140,I255087);
nor I_14840 (I255157,I255140,I254714);
nor I_14841 (I255174,I254979,I255157);
DFFARX1 I_14842 (I255174,I2859,I254654,I254643,);
not I_14843 (I255232,I2866);
DFFARX1 I_14844 (I108190,I2859,I255232,I255258,);
not I_14845 (I255266,I255258);
DFFARX1 I_14846 (I108205,I2859,I255232,I255292,);
not I_14847 (I255300,I108208);
nand I_14848 (I255317,I255300,I108187);
not I_14849 (I255334,I255317);
nor I_14850 (I255351,I255334,I108211);
nor I_14851 (I255368,I255266,I255351);
DFFARX1 I_14852 (I255368,I2859,I255232,I255218,);
not I_14853 (I255399,I108211);
nand I_14854 (I255416,I255399,I255334);
and I_14855 (I255433,I255399,I108193);
nand I_14856 (I255450,I255433,I108184);
nor I_14857 (I255215,I255450,I255399);
and I_14858 (I255206,I255292,I255450);
not I_14859 (I255495,I255450);
nand I_14860 (I255209,I255292,I255495);
nor I_14861 (I255203,I255258,I255450);
not I_14862 (I255540,I108184);
nor I_14863 (I255557,I255540,I108193);
nand I_14864 (I255574,I255557,I255399);
nor I_14865 (I255212,I255317,I255574);
nor I_14866 (I255605,I255540,I108199);
and I_14867 (I255622,I255605,I108202);
or I_14868 (I255639,I255622,I108196);
DFFARX1 I_14869 (I255639,I2859,I255232,I255665,);
nor I_14870 (I255673,I255665,I255416);
DFFARX1 I_14871 (I255673,I2859,I255232,I255200,);
DFFARX1 I_14872 (I255665,I2859,I255232,I255224,);
not I_14873 (I255718,I255665);
nor I_14874 (I255735,I255718,I255292);
nor I_14875 (I255752,I255557,I255735);
DFFARX1 I_14876 (I255752,I2859,I255232,I255221,);
not I_14877 (I255810,I2866);
DFFARX1 I_14878 (I69133,I2859,I255810,I255836,);
not I_14879 (I255844,I255836);
DFFARX1 I_14880 (I69118,I2859,I255810,I255870,);
not I_14881 (I255878,I69136);
nand I_14882 (I255895,I255878,I69121);
not I_14883 (I255912,I255895);
nor I_14884 (I255929,I255912,I69118);
nor I_14885 (I255946,I255844,I255929);
DFFARX1 I_14886 (I255946,I2859,I255810,I255796,);
not I_14887 (I255977,I69118);
nand I_14888 (I255994,I255977,I255912);
and I_14889 (I256011,I255977,I69121);
nand I_14890 (I256028,I256011,I69142);
nor I_14891 (I255793,I256028,I255977);
and I_14892 (I255784,I255870,I256028);
not I_14893 (I256073,I256028);
nand I_14894 (I255787,I255870,I256073);
nor I_14895 (I255781,I255836,I256028);
not I_14896 (I256118,I69130);
nor I_14897 (I256135,I256118,I69121);
nand I_14898 (I256152,I256135,I255977);
nor I_14899 (I255790,I255895,I256152);
nor I_14900 (I256183,I256118,I69124);
and I_14901 (I256200,I256183,I69139);
or I_14902 (I256217,I256200,I69127);
DFFARX1 I_14903 (I256217,I2859,I255810,I256243,);
nor I_14904 (I256251,I256243,I255994);
DFFARX1 I_14905 (I256251,I2859,I255810,I255778,);
DFFARX1 I_14906 (I256243,I2859,I255810,I255802,);
not I_14907 (I256296,I256243);
nor I_14908 (I256313,I256296,I255870);
nor I_14909 (I256330,I256135,I256313);
DFFARX1 I_14910 (I256330,I2859,I255810,I255799,);
not I_14911 (I256388,I2866);
DFFARX1 I_14912 (I354265,I2859,I256388,I256414,);
not I_14913 (I256422,I256414);
DFFARX1 I_14914 (I354265,I2859,I256388,I256448,);
not I_14915 (I256456,I354262);
nand I_14916 (I256473,I256456,I354277);
not I_14917 (I256490,I256473);
nor I_14918 (I256507,I256490,I354271);
nor I_14919 (I256524,I256422,I256507);
DFFARX1 I_14920 (I256524,I2859,I256388,I256374,);
not I_14921 (I256555,I354271);
nand I_14922 (I256572,I256555,I256490);
and I_14923 (I256589,I256555,I354268);
nand I_14924 (I256606,I256589,I354259);
nor I_14925 (I256371,I256606,I256555);
and I_14926 (I256362,I256448,I256606);
not I_14927 (I256651,I256606);
nand I_14928 (I256365,I256448,I256651);
nor I_14929 (I256359,I256414,I256606);
not I_14930 (I256696,I354280);
nor I_14931 (I256713,I256696,I354268);
nand I_14932 (I256730,I256713,I256555);
nor I_14933 (I256368,I256473,I256730);
nor I_14934 (I256761,I256696,I354259);
and I_14935 (I256778,I256761,I354262);
or I_14936 (I256795,I256778,I354274);
DFFARX1 I_14937 (I256795,I2859,I256388,I256821,);
nor I_14938 (I256829,I256821,I256572);
DFFARX1 I_14939 (I256829,I2859,I256388,I256356,);
DFFARX1 I_14940 (I256821,I2859,I256388,I256380,);
not I_14941 (I256874,I256821);
nor I_14942 (I256891,I256874,I256448);
nor I_14943 (I256908,I256713,I256891);
DFFARX1 I_14944 (I256908,I2859,I256388,I256377,);
not I_14945 (I256966,I2866);
DFFARX1 I_14946 (I64968,I2859,I256966,I256992,);
not I_14947 (I257000,I256992);
DFFARX1 I_14948 (I64953,I2859,I256966,I257026,);
not I_14949 (I257034,I64971);
nand I_14950 (I257051,I257034,I64956);
not I_14951 (I257068,I257051);
nor I_14952 (I257085,I257068,I64953);
nor I_14953 (I257102,I257000,I257085);
DFFARX1 I_14954 (I257102,I2859,I256966,I256952,);
not I_14955 (I257133,I64953);
nand I_14956 (I257150,I257133,I257068);
and I_14957 (I257167,I257133,I64956);
nand I_14958 (I257184,I257167,I64977);
nor I_14959 (I256949,I257184,I257133);
and I_14960 (I256940,I257026,I257184);
not I_14961 (I257229,I257184);
nand I_14962 (I256943,I257026,I257229);
nor I_14963 (I256937,I256992,I257184);
not I_14964 (I257274,I64965);
nor I_14965 (I257291,I257274,I64956);
nand I_14966 (I257308,I257291,I257133);
nor I_14967 (I256946,I257051,I257308);
nor I_14968 (I257339,I257274,I64959);
and I_14969 (I257356,I257339,I64974);
or I_14970 (I257373,I257356,I64962);
DFFARX1 I_14971 (I257373,I2859,I256966,I257399,);
nor I_14972 (I257407,I257399,I257150);
DFFARX1 I_14973 (I257407,I2859,I256966,I256934,);
DFFARX1 I_14974 (I257399,I2859,I256966,I256958,);
not I_14975 (I257452,I257399);
nor I_14976 (I257469,I257452,I257026);
nor I_14977 (I257486,I257291,I257469);
DFFARX1 I_14978 (I257486,I2859,I256966,I256955,);
not I_14979 (I257544,I2866);
DFFARX1 I_14980 (I325138,I2859,I257544,I257570,);
not I_14981 (I257578,I257570);
DFFARX1 I_14982 (I325150,I2859,I257544,I257604,);
not I_14983 (I257612,I325141);
nand I_14984 (I257629,I257612,I325144);
not I_14985 (I257646,I257629);
nor I_14986 (I257663,I257646,I325147);
nor I_14987 (I257680,I257578,I257663);
DFFARX1 I_14988 (I257680,I2859,I257544,I257530,);
not I_14989 (I257711,I325147);
nand I_14990 (I257728,I257711,I257646);
and I_14991 (I257745,I257711,I325141);
nand I_14992 (I257762,I257745,I325153);
nor I_14993 (I257527,I257762,I257711);
and I_14994 (I257518,I257604,I257762);
not I_14995 (I257807,I257762);
nand I_14996 (I257521,I257604,I257807);
nor I_14997 (I257515,I257570,I257762);
not I_14998 (I257852,I325159);
nor I_14999 (I257869,I257852,I325141);
nand I_15000 (I257886,I257869,I257711);
nor I_15001 (I257524,I257629,I257886);
nor I_15002 (I257917,I257852,I325138);
and I_15003 (I257934,I257917,I325156);
or I_15004 (I257951,I257934,I325162);
DFFARX1 I_15005 (I257951,I2859,I257544,I257977,);
nor I_15006 (I257985,I257977,I257728);
DFFARX1 I_15007 (I257985,I2859,I257544,I257512,);
DFFARX1 I_15008 (I257977,I2859,I257544,I257536,);
not I_15009 (I258030,I257977);
nor I_15010 (I258047,I258030,I257604);
nor I_15011 (I258064,I257869,I258047);
DFFARX1 I_15012 (I258064,I2859,I257544,I257533,);
not I_15013 (I258122,I2866);
DFFARX1 I_15014 (I173799,I2859,I258122,I258148,);
not I_15015 (I258156,I258148);
DFFARX1 I_15016 (I173811,I2859,I258122,I258182,);
not I_15017 (I258190,I173787);
nand I_15018 (I258207,I258190,I173814);
not I_15019 (I258224,I258207);
nor I_15020 (I258241,I258224,I173802);
nor I_15021 (I258258,I258156,I258241);
DFFARX1 I_15022 (I258258,I2859,I258122,I258108,);
not I_15023 (I258289,I173802);
nand I_15024 (I258306,I258289,I258224);
and I_15025 (I258323,I258289,I173787);
nand I_15026 (I258340,I258323,I173790);
nor I_15027 (I258105,I258340,I258289);
and I_15028 (I258096,I258182,I258340);
not I_15029 (I258385,I258340);
nand I_15030 (I258099,I258182,I258385);
nor I_15031 (I258093,I258148,I258340);
not I_15032 (I258430,I173796);
nor I_15033 (I258447,I258430,I173787);
nand I_15034 (I258464,I258447,I258289);
nor I_15035 (I258102,I258207,I258464);
nor I_15036 (I258495,I258430,I173805);
and I_15037 (I258512,I258495,I173793);
or I_15038 (I258529,I258512,I173808);
DFFARX1 I_15039 (I258529,I2859,I258122,I258555,);
nor I_15040 (I258563,I258555,I258306);
DFFARX1 I_15041 (I258563,I2859,I258122,I258090,);
DFFARX1 I_15042 (I258555,I2859,I258122,I258114,);
not I_15043 (I258608,I258555);
nor I_15044 (I258625,I258608,I258182);
nor I_15045 (I258642,I258447,I258625);
DFFARX1 I_15046 (I258642,I2859,I258122,I258111,);
not I_15047 (I258700,I2866);
DFFARX1 I_15048 (I307798,I2859,I258700,I258726,);
not I_15049 (I258734,I258726);
DFFARX1 I_15050 (I307810,I2859,I258700,I258760,);
not I_15051 (I258768,I307801);
nand I_15052 (I258785,I258768,I307804);
not I_15053 (I258802,I258785);
nor I_15054 (I258819,I258802,I307807);
nor I_15055 (I258836,I258734,I258819);
DFFARX1 I_15056 (I258836,I2859,I258700,I258686,);
not I_15057 (I258867,I307807);
nand I_15058 (I258884,I258867,I258802);
and I_15059 (I258901,I258867,I307801);
nand I_15060 (I258918,I258901,I307813);
nor I_15061 (I258683,I258918,I258867);
and I_15062 (I258674,I258760,I258918);
not I_15063 (I258963,I258918);
nand I_15064 (I258677,I258760,I258963);
nor I_15065 (I258671,I258726,I258918);
not I_15066 (I259008,I307819);
nor I_15067 (I259025,I259008,I307801);
nand I_15068 (I259042,I259025,I258867);
nor I_15069 (I258680,I258785,I259042);
nor I_15070 (I259073,I259008,I307798);
and I_15071 (I259090,I259073,I307816);
or I_15072 (I259107,I259090,I307822);
DFFARX1 I_15073 (I259107,I2859,I258700,I259133,);
nor I_15074 (I259141,I259133,I258884);
DFFARX1 I_15075 (I259141,I2859,I258700,I258668,);
DFFARX1 I_15076 (I259133,I2859,I258700,I258692,);
not I_15077 (I259186,I259133);
nor I_15078 (I259203,I259186,I258760);
nor I_15079 (I259220,I259025,I259203);
DFFARX1 I_15080 (I259220,I2859,I258700,I258689,);
not I_15081 (I259278,I2866);
DFFARX1 I_15082 (I374818,I2859,I259278,I259304,);
not I_15083 (I259312,I259304);
DFFARX1 I_15084 (I374818,I2859,I259278,I259338,);
not I_15085 (I259346,I374815);
nand I_15086 (I259363,I259346,I374830);
not I_15087 (I259380,I259363);
nor I_15088 (I259397,I259380,I374824);
nor I_15089 (I259414,I259312,I259397);
DFFARX1 I_15090 (I259414,I2859,I259278,I259264,);
not I_15091 (I259445,I374824);
nand I_15092 (I259462,I259445,I259380);
and I_15093 (I259479,I259445,I374821);
nand I_15094 (I259496,I259479,I374812);
nor I_15095 (I259261,I259496,I259445);
and I_15096 (I259252,I259338,I259496);
not I_15097 (I259541,I259496);
nand I_15098 (I259255,I259338,I259541);
nor I_15099 (I259249,I259304,I259496);
not I_15100 (I259586,I374833);
nor I_15101 (I259603,I259586,I374821);
nand I_15102 (I259620,I259603,I259445);
nor I_15103 (I259258,I259363,I259620);
nor I_15104 (I259651,I259586,I374812);
and I_15105 (I259668,I259651,I374815);
or I_15106 (I259685,I259668,I374827);
DFFARX1 I_15107 (I259685,I2859,I259278,I259711,);
nor I_15108 (I259719,I259711,I259462);
DFFARX1 I_15109 (I259719,I2859,I259278,I259246,);
DFFARX1 I_15110 (I259711,I2859,I259278,I259270,);
not I_15111 (I259764,I259711);
nor I_15112 (I259781,I259764,I259338);
nor I_15113 (I259798,I259603,I259781);
DFFARX1 I_15114 (I259798,I2859,I259278,I259267,);
not I_15115 (I259856,I2866);
DFFARX1 I_15116 (I152985,I2859,I259856,I259882,);
not I_15117 (I259890,I259882);
DFFARX1 I_15118 (I153000,I2859,I259856,I259916,);
not I_15119 (I259924,I153003);
nand I_15120 (I259941,I259924,I152982);
not I_15121 (I259958,I259941);
nor I_15122 (I259975,I259958,I153006);
nor I_15123 (I259992,I259890,I259975);
DFFARX1 I_15124 (I259992,I2859,I259856,I259842,);
not I_15125 (I260023,I153006);
nand I_15126 (I260040,I260023,I259958);
and I_15127 (I260057,I260023,I152988);
nand I_15128 (I260074,I260057,I152979);
nor I_15129 (I259839,I260074,I260023);
and I_15130 (I259830,I259916,I260074);
not I_15131 (I260119,I260074);
nand I_15132 (I259833,I259916,I260119);
nor I_15133 (I259827,I259882,I260074);
not I_15134 (I260164,I152979);
nor I_15135 (I260181,I260164,I152988);
nand I_15136 (I260198,I260181,I260023);
nor I_15137 (I259836,I259941,I260198);
nor I_15138 (I260229,I260164,I152994);
and I_15139 (I260246,I260229,I152997);
or I_15140 (I260263,I260246,I152991);
DFFARX1 I_15141 (I260263,I2859,I259856,I260289,);
nor I_15142 (I260297,I260289,I260040);
DFFARX1 I_15143 (I260297,I2859,I259856,I259824,);
DFFARX1 I_15144 (I260289,I2859,I259856,I259848,);
not I_15145 (I260342,I260289);
nor I_15146 (I260359,I260342,I259916);
nor I_15147 (I260376,I260181,I260359);
DFFARX1 I_15148 (I260376,I2859,I259856,I259845,);
not I_15149 (I260434,I2866);
DFFARX1 I_15150 (I187399,I2859,I260434,I260460,);
not I_15151 (I260468,I260460);
DFFARX1 I_15152 (I187411,I2859,I260434,I260494,);
not I_15153 (I260502,I187387);
nand I_15154 (I260519,I260502,I187414);
not I_15155 (I260536,I260519);
nor I_15156 (I260553,I260536,I187402);
nor I_15157 (I260570,I260468,I260553);
DFFARX1 I_15158 (I260570,I2859,I260434,I260420,);
not I_15159 (I260601,I187402);
nand I_15160 (I260618,I260601,I260536);
and I_15161 (I260635,I260601,I187387);
nand I_15162 (I260652,I260635,I187390);
nor I_15163 (I260417,I260652,I260601);
and I_15164 (I260408,I260494,I260652);
not I_15165 (I260697,I260652);
nand I_15166 (I260411,I260494,I260697);
nor I_15167 (I260405,I260460,I260652);
not I_15168 (I260742,I187396);
nor I_15169 (I260759,I260742,I187387);
nand I_15170 (I260776,I260759,I260601);
nor I_15171 (I260414,I260519,I260776);
nor I_15172 (I260807,I260742,I187405);
and I_15173 (I260824,I260807,I187393);
or I_15174 (I260841,I260824,I187408);
DFFARX1 I_15175 (I260841,I2859,I260434,I260867,);
nor I_15176 (I260875,I260867,I260618);
DFFARX1 I_15177 (I260875,I2859,I260434,I260402,);
DFFARX1 I_15178 (I260867,I2859,I260434,I260426,);
not I_15179 (I260920,I260867);
nor I_15180 (I260937,I260920,I260494);
nor I_15181 (I260954,I260759,I260937);
DFFARX1 I_15182 (I260954,I2859,I260434,I260423,);
not I_15183 (I261012,I2866);
DFFARX1 I_15184 (I543095,I2859,I261012,I261038,);
not I_15185 (I261046,I261038);
DFFARX1 I_15186 (I543095,I2859,I261012,I261072,);
not I_15187 (I261080,I543119);
nand I_15188 (I261097,I261080,I543101);
not I_15189 (I261114,I261097);
nor I_15190 (I261131,I261114,I543116);
nor I_15191 (I261148,I261046,I261131);
DFFARX1 I_15192 (I261148,I2859,I261012,I260998,);
not I_15193 (I261179,I543116);
nand I_15194 (I261196,I261179,I261114);
and I_15195 (I261213,I261179,I543098);
nand I_15196 (I261230,I261213,I543107);
nor I_15197 (I260995,I261230,I261179);
and I_15198 (I260986,I261072,I261230);
not I_15199 (I261275,I261230);
nand I_15200 (I260989,I261072,I261275);
nor I_15201 (I260983,I261038,I261230);
not I_15202 (I261320,I543104);
nor I_15203 (I261337,I261320,I543098);
nand I_15204 (I261354,I261337,I261179);
nor I_15205 (I260992,I261097,I261354);
nor I_15206 (I261385,I261320,I543113);
and I_15207 (I261402,I261385,I543122);
or I_15208 (I261419,I261402,I543110);
DFFARX1 I_15209 (I261419,I2859,I261012,I261445,);
nor I_15210 (I261453,I261445,I261196);
DFFARX1 I_15211 (I261453,I2859,I261012,I260980,);
DFFARX1 I_15212 (I261445,I2859,I261012,I261004,);
not I_15213 (I261498,I261445);
nor I_15214 (I261515,I261498,I261072);
nor I_15215 (I261532,I261337,I261515);
DFFARX1 I_15216 (I261532,I2859,I261012,I261001,);
not I_15217 (I261590,I2866);
DFFARX1 I_15218 (I75083,I2859,I261590,I261616,);
not I_15219 (I261624,I261616);
DFFARX1 I_15220 (I75068,I2859,I261590,I261650,);
not I_15221 (I261658,I75086);
nand I_15222 (I261675,I261658,I75071);
not I_15223 (I261692,I261675);
nor I_15224 (I261709,I261692,I75068);
nor I_15225 (I261726,I261624,I261709);
DFFARX1 I_15226 (I261726,I2859,I261590,I261576,);
not I_15227 (I261757,I75068);
nand I_15228 (I261774,I261757,I261692);
and I_15229 (I261791,I261757,I75071);
nand I_15230 (I261808,I261791,I75092);
nor I_15231 (I261573,I261808,I261757);
and I_15232 (I261564,I261650,I261808);
not I_15233 (I261853,I261808);
nand I_15234 (I261567,I261650,I261853);
nor I_15235 (I261561,I261616,I261808);
not I_15236 (I261898,I75080);
nor I_15237 (I261915,I261898,I75071);
nand I_15238 (I261932,I261915,I261757);
nor I_15239 (I261570,I261675,I261932);
nor I_15240 (I261963,I261898,I75074);
and I_15241 (I261980,I261963,I75089);
or I_15242 (I261997,I261980,I75077);
DFFARX1 I_15243 (I261997,I2859,I261590,I262023,);
nor I_15244 (I262031,I262023,I261774);
DFFARX1 I_15245 (I262031,I2859,I261590,I261558,);
DFFARX1 I_15246 (I262023,I2859,I261590,I261582,);
not I_15247 (I262076,I262023);
nor I_15248 (I262093,I262076,I261650);
nor I_15249 (I262110,I261915,I262093);
DFFARX1 I_15250 (I262110,I2859,I261590,I261579,);
not I_15251 (I262168,I2866);
DFFARX1 I_15252 (I556185,I2859,I262168,I262194,);
not I_15253 (I262202,I262194);
DFFARX1 I_15254 (I556185,I2859,I262168,I262228,);
not I_15255 (I262236,I556209);
nand I_15256 (I262253,I262236,I556191);
not I_15257 (I262270,I262253);
nor I_15258 (I262287,I262270,I556206);
nor I_15259 (I262304,I262202,I262287);
DFFARX1 I_15260 (I262304,I2859,I262168,I262154,);
not I_15261 (I262335,I556206);
nand I_15262 (I262352,I262335,I262270);
and I_15263 (I262369,I262335,I556188);
nand I_15264 (I262386,I262369,I556197);
nor I_15265 (I262151,I262386,I262335);
and I_15266 (I262142,I262228,I262386);
not I_15267 (I262431,I262386);
nand I_15268 (I262145,I262228,I262431);
nor I_15269 (I262139,I262194,I262386);
not I_15270 (I262476,I556194);
nor I_15271 (I262493,I262476,I556188);
nand I_15272 (I262510,I262493,I262335);
nor I_15273 (I262148,I262253,I262510);
nor I_15274 (I262541,I262476,I556203);
and I_15275 (I262558,I262541,I556212);
or I_15276 (I262575,I262558,I556200);
DFFARX1 I_15277 (I262575,I2859,I262168,I262601,);
nor I_15278 (I262609,I262601,I262352);
DFFARX1 I_15279 (I262609,I2859,I262168,I262136,);
DFFARX1 I_15280 (I262601,I2859,I262168,I262160,);
not I_15281 (I262654,I262601);
nor I_15282 (I262671,I262654,I262228);
nor I_15283 (I262688,I262493,I262671);
DFFARX1 I_15284 (I262688,I2859,I262168,I262157,);
not I_15285 (I262746,I2866);
DFFARX1 I_15286 (I39987,I2859,I262746,I262772,);
not I_15287 (I262780,I262772);
DFFARX1 I_15288 (I39966,I2859,I262746,I262806,);
not I_15289 (I262814,I39963);
nand I_15290 (I262831,I262814,I39978);
not I_15291 (I262848,I262831);
nor I_15292 (I262865,I262848,I39966);
nor I_15293 (I262882,I262780,I262865);
DFFARX1 I_15294 (I262882,I2859,I262746,I262732,);
not I_15295 (I262913,I39966);
nand I_15296 (I262930,I262913,I262848);
and I_15297 (I262947,I262913,I39969);
nand I_15298 (I262964,I262947,I39984);
nor I_15299 (I262729,I262964,I262913);
and I_15300 (I262720,I262806,I262964);
not I_15301 (I263009,I262964);
nand I_15302 (I262723,I262806,I263009);
nor I_15303 (I262717,I262772,I262964);
not I_15304 (I263054,I39975);
nor I_15305 (I263071,I263054,I39969);
nand I_15306 (I263088,I263071,I262913);
nor I_15307 (I262726,I262831,I263088);
nor I_15308 (I263119,I263054,I39963);
and I_15309 (I263136,I263119,I39972);
or I_15310 (I263153,I263136,I39981);
DFFARX1 I_15311 (I263153,I2859,I262746,I263179,);
nor I_15312 (I263187,I263179,I262930);
DFFARX1 I_15313 (I263187,I2859,I262746,I262714,);
DFFARX1 I_15314 (I263179,I2859,I262746,I262738,);
not I_15315 (I263232,I263179);
nor I_15316 (I263249,I263232,I262806);
nor I_15317 (I263266,I263071,I263249);
DFFARX1 I_15318 (I263266,I2859,I262746,I262735,);
not I_15319 (I263324,I2866);
DFFARX1 I_15320 (I499762,I2859,I263324,I263350,);
not I_15321 (I263358,I263350);
DFFARX1 I_15322 (I499768,I2859,I263324,I263384,);
not I_15323 (I263392,I499762);
nand I_15324 (I263409,I263392,I499765);
not I_15325 (I263426,I263409);
nor I_15326 (I263443,I263426,I499783);
nor I_15327 (I263460,I263358,I263443);
DFFARX1 I_15328 (I263460,I2859,I263324,I263310,);
not I_15329 (I263491,I499783);
nand I_15330 (I263508,I263491,I263426);
and I_15331 (I263525,I263491,I499786);
nand I_15332 (I263542,I263525,I499765);
nor I_15333 (I263307,I263542,I263491);
and I_15334 (I263298,I263384,I263542);
not I_15335 (I263587,I263542);
nand I_15336 (I263301,I263384,I263587);
nor I_15337 (I263295,I263350,I263542);
not I_15338 (I263632,I499771);
nor I_15339 (I263649,I263632,I499786);
nand I_15340 (I263666,I263649,I263491);
nor I_15341 (I263304,I263409,I263666);
nor I_15342 (I263697,I263632,I499777);
and I_15343 (I263714,I263697,I499774);
or I_15344 (I263731,I263714,I499780);
DFFARX1 I_15345 (I263731,I2859,I263324,I263757,);
nor I_15346 (I263765,I263757,I263508);
DFFARX1 I_15347 (I263765,I2859,I263324,I263292,);
DFFARX1 I_15348 (I263757,I2859,I263324,I263316,);
not I_15349 (I263810,I263757);
nor I_15350 (I263827,I263810,I263384);
nor I_15351 (I263844,I263649,I263827);
DFFARX1 I_15352 (I263844,I2859,I263324,I263313,);
not I_15353 (I263902,I2866);
DFFARX1 I_15354 (I315890,I2859,I263902,I263928,);
not I_15355 (I263936,I263928);
DFFARX1 I_15356 (I315902,I2859,I263902,I263962,);
not I_15357 (I263970,I315893);
nand I_15358 (I263987,I263970,I315896);
not I_15359 (I264004,I263987);
nor I_15360 (I264021,I264004,I315899);
nor I_15361 (I264038,I263936,I264021);
DFFARX1 I_15362 (I264038,I2859,I263902,I263888,);
not I_15363 (I264069,I315899);
nand I_15364 (I264086,I264069,I264004);
and I_15365 (I264103,I264069,I315893);
nand I_15366 (I264120,I264103,I315905);
nor I_15367 (I263885,I264120,I264069);
and I_15368 (I263876,I263962,I264120);
not I_15369 (I264165,I264120);
nand I_15370 (I263879,I263962,I264165);
nor I_15371 (I263873,I263928,I264120);
not I_15372 (I264210,I315911);
nor I_15373 (I264227,I264210,I315893);
nand I_15374 (I264244,I264227,I264069);
nor I_15375 (I263882,I263987,I264244);
nor I_15376 (I264275,I264210,I315890);
and I_15377 (I264292,I264275,I315908);
or I_15378 (I264309,I264292,I315914);
DFFARX1 I_15379 (I264309,I2859,I263902,I264335,);
nor I_15380 (I264343,I264335,I264086);
DFFARX1 I_15381 (I264343,I2859,I263902,I263870,);
DFFARX1 I_15382 (I264335,I2859,I263902,I263894,);
not I_15383 (I264388,I264335);
nor I_15384 (I264405,I264388,I263962);
nor I_15385 (I264422,I264227,I264405);
DFFARX1 I_15386 (I264422,I2859,I263902,I263891,);
not I_15387 (I264480,I2866);
DFFARX1 I_15388 (I353738,I2859,I264480,I264506,);
not I_15389 (I264514,I264506);
DFFARX1 I_15390 (I353738,I2859,I264480,I264540,);
not I_15391 (I264548,I353735);
nand I_15392 (I264565,I264548,I353750);
not I_15393 (I264582,I264565);
nor I_15394 (I264599,I264582,I353744);
nor I_15395 (I264616,I264514,I264599);
DFFARX1 I_15396 (I264616,I2859,I264480,I264466,);
not I_15397 (I264647,I353744);
nand I_15398 (I264664,I264647,I264582);
and I_15399 (I264681,I264647,I353741);
nand I_15400 (I264698,I264681,I353732);
nor I_15401 (I264463,I264698,I264647);
and I_15402 (I264454,I264540,I264698);
not I_15403 (I264743,I264698);
nand I_15404 (I264457,I264540,I264743);
nor I_15405 (I264451,I264506,I264698);
not I_15406 (I264788,I353753);
nor I_15407 (I264805,I264788,I353741);
nand I_15408 (I264822,I264805,I264647);
nor I_15409 (I264460,I264565,I264822);
nor I_15410 (I264853,I264788,I353732);
and I_15411 (I264870,I264853,I353735);
or I_15412 (I264887,I264870,I353747);
DFFARX1 I_15413 (I264887,I2859,I264480,I264913,);
nor I_15414 (I264921,I264913,I264664);
DFFARX1 I_15415 (I264921,I2859,I264480,I264448,);
DFFARX1 I_15416 (I264913,I2859,I264480,I264472,);
not I_15417 (I264966,I264913);
nor I_15418 (I264983,I264966,I264540);
nor I_15419 (I265000,I264805,I264983);
DFFARX1 I_15420 (I265000,I2859,I264480,I264469,);
not I_15421 (I265058,I2866);
DFFARX1 I_15422 (I73283,I2859,I265058,I265084,);
not I_15423 (I265092,I265084);
nand I_15424 (I265109,I73286,I73307);
and I_15425 (I265126,I265109,I73295);
DFFARX1 I_15426 (I265126,I2859,I265058,I265152,);
not I_15427 (I265160,I73292);
DFFARX1 I_15428 (I73283,I2859,I265058,I265186,);
not I_15429 (I265194,I265186);
nor I_15430 (I265211,I265194,I265092);
and I_15431 (I265228,I265211,I73292);
nor I_15432 (I265245,I265194,I265160);
nor I_15433 (I265041,I265152,I265245);
DFFARX1 I_15434 (I73301,I2859,I265058,I265285,);
nor I_15435 (I265293,I265285,I265152);
not I_15436 (I265310,I265293);
not I_15437 (I265327,I265285);
nor I_15438 (I265344,I265327,I265228);
DFFARX1 I_15439 (I265344,I2859,I265058,I265044,);
nand I_15440 (I265375,I73286,I73289);
and I_15441 (I265392,I265375,I73298);
DFFARX1 I_15442 (I265392,I2859,I265058,I265418,);
nor I_15443 (I265426,I265418,I265285);
DFFARX1 I_15444 (I265426,I2859,I265058,I265026,);
nand I_15445 (I265457,I265418,I265327);
nand I_15446 (I265035,I265310,I265457);
not I_15447 (I265488,I265418);
nor I_15448 (I265505,I265488,I265228);
DFFARX1 I_15449 (I265505,I2859,I265058,I265047,);
nor I_15450 (I265536,I73304,I73289);
or I_15451 (I265038,I265285,I265536);
nor I_15452 (I265029,I265418,I265536);
or I_15453 (I265032,I265152,I265536);
DFFARX1 I_15454 (I265536,I2859,I265058,I265050,);
not I_15455 (I265636,I2866);
DFFARX1 I_15456 (I459320,I2859,I265636,I265662,);
not I_15457 (I265670,I265662);
nand I_15458 (I265687,I459302,I459314);
and I_15459 (I265704,I265687,I459317);
DFFARX1 I_15460 (I265704,I2859,I265636,I265730,);
not I_15461 (I265738,I459311);
DFFARX1 I_15462 (I459308,I2859,I265636,I265764,);
not I_15463 (I265772,I265764);
nor I_15464 (I265789,I265772,I265670);
and I_15465 (I265806,I265789,I459311);
nor I_15466 (I265823,I265772,I265738);
nor I_15467 (I265619,I265730,I265823);
DFFARX1 I_15468 (I459326,I2859,I265636,I265863,);
nor I_15469 (I265871,I265863,I265730);
not I_15470 (I265888,I265871);
not I_15471 (I265905,I265863);
nor I_15472 (I265922,I265905,I265806);
DFFARX1 I_15473 (I265922,I2859,I265636,I265622,);
nand I_15474 (I265953,I459305,I459305);
and I_15475 (I265970,I265953,I459302);
DFFARX1 I_15476 (I265970,I2859,I265636,I265996,);
nor I_15477 (I266004,I265996,I265863);
DFFARX1 I_15478 (I266004,I2859,I265636,I265604,);
nand I_15479 (I266035,I265996,I265905);
nand I_15480 (I265613,I265888,I266035);
not I_15481 (I266066,I265996);
nor I_15482 (I266083,I266066,I265806);
DFFARX1 I_15483 (I266083,I2859,I265636,I265625,);
nor I_15484 (I266114,I459323,I459305);
or I_15485 (I265616,I265863,I266114);
nor I_15486 (I265607,I265996,I266114);
or I_15487 (I265610,I265730,I266114);
DFFARX1 I_15488 (I266114,I2859,I265636,I265628,);
not I_15489 (I266214,I2866);
DFFARX1 I_15490 (I234392,I2859,I266214,I266240,);
not I_15491 (I266248,I266240);
nand I_15492 (I266265,I234401,I234410);
and I_15493 (I266282,I266265,I234416);
DFFARX1 I_15494 (I266282,I2859,I266214,I266308,);
not I_15495 (I266316,I234413);
DFFARX1 I_15496 (I234398,I2859,I266214,I266342,);
not I_15497 (I266350,I266342);
nor I_15498 (I266367,I266350,I266248);
and I_15499 (I266384,I266367,I234413);
nor I_15500 (I266401,I266350,I266316);
nor I_15501 (I266197,I266308,I266401);
DFFARX1 I_15502 (I234407,I2859,I266214,I266441,);
nor I_15503 (I266449,I266441,I266308);
not I_15504 (I266466,I266449);
not I_15505 (I266483,I266441);
nor I_15506 (I266500,I266483,I266384);
DFFARX1 I_15507 (I266500,I2859,I266214,I266200,);
nand I_15508 (I266531,I234404,I234395);
and I_15509 (I266548,I266531,I234392);
DFFARX1 I_15510 (I266548,I2859,I266214,I266574,);
nor I_15511 (I266582,I266574,I266441);
DFFARX1 I_15512 (I266582,I2859,I266214,I266182,);
nand I_15513 (I266613,I266574,I266483);
nand I_15514 (I266191,I266466,I266613);
not I_15515 (I266644,I266574);
nor I_15516 (I266661,I266644,I266384);
DFFARX1 I_15517 (I266661,I2859,I266214,I266203,);
nor I_15518 (I266692,I234395,I234395);
or I_15519 (I266194,I266441,I266692);
nor I_15520 (I266185,I266574,I266692);
or I_15521 (I266188,I266308,I266692);
DFFARX1 I_15522 (I266692,I2859,I266214,I266206,);
not I_15523 (I266792,I2866);
DFFARX1 I_15524 (I46290,I2859,I266792,I266818,);
not I_15525 (I266826,I266818);
nand I_15526 (I266843,I46299,I46308);
and I_15527 (I266860,I266843,I46287);
DFFARX1 I_15528 (I266860,I2859,I266792,I266886,);
not I_15529 (I266894,I46290);
DFFARX1 I_15530 (I46305,I2859,I266792,I266920,);
not I_15531 (I266928,I266920);
nor I_15532 (I266945,I266928,I266826);
and I_15533 (I266962,I266945,I46290);
nor I_15534 (I266979,I266928,I266894);
nor I_15535 (I266775,I266886,I266979);
DFFARX1 I_15536 (I46296,I2859,I266792,I267019,);
nor I_15537 (I267027,I267019,I266886);
not I_15538 (I267044,I267027);
not I_15539 (I267061,I267019);
nor I_15540 (I267078,I267061,I266962);
DFFARX1 I_15541 (I267078,I2859,I266792,I266778,);
nand I_15542 (I267109,I46311,I46287);
and I_15543 (I267126,I267109,I46293);
DFFARX1 I_15544 (I267126,I2859,I266792,I267152,);
nor I_15545 (I267160,I267152,I267019);
DFFARX1 I_15546 (I267160,I2859,I266792,I266760,);
nand I_15547 (I267191,I267152,I267061);
nand I_15548 (I266769,I267044,I267191);
not I_15549 (I267222,I267152);
nor I_15550 (I267239,I267222,I266962);
DFFARX1 I_15551 (I267239,I2859,I266792,I266781,);
nor I_15552 (I267270,I46302,I46287);
or I_15553 (I266772,I267019,I267270);
nor I_15554 (I266763,I267152,I267270);
or I_15555 (I266766,I266886,I267270);
DFFARX1 I_15556 (I267270,I2859,I266792,I266784,);
not I_15557 (I267370,I2866);
DFFARX1 I_15558 (I22575,I2859,I267370,I267396,);
not I_15559 (I267404,I267396);
nand I_15560 (I267421,I22584,I22593);
and I_15561 (I267438,I267421,I22572);
DFFARX1 I_15562 (I267438,I2859,I267370,I267464,);
not I_15563 (I267472,I22575);
DFFARX1 I_15564 (I22590,I2859,I267370,I267498,);
not I_15565 (I267506,I267498);
nor I_15566 (I267523,I267506,I267404);
and I_15567 (I267540,I267523,I22575);
nor I_15568 (I267557,I267506,I267472);
nor I_15569 (I267353,I267464,I267557);
DFFARX1 I_15570 (I22581,I2859,I267370,I267597,);
nor I_15571 (I267605,I267597,I267464);
not I_15572 (I267622,I267605);
not I_15573 (I267639,I267597);
nor I_15574 (I267656,I267639,I267540);
DFFARX1 I_15575 (I267656,I2859,I267370,I267356,);
nand I_15576 (I267687,I22596,I22572);
and I_15577 (I267704,I267687,I22578);
DFFARX1 I_15578 (I267704,I2859,I267370,I267730,);
nor I_15579 (I267738,I267730,I267597);
DFFARX1 I_15580 (I267738,I2859,I267370,I267338,);
nand I_15581 (I267769,I267730,I267639);
nand I_15582 (I267347,I267622,I267769);
not I_15583 (I267800,I267730);
nor I_15584 (I267817,I267800,I267540);
DFFARX1 I_15585 (I267817,I2859,I267370,I267359,);
nor I_15586 (I267848,I22587,I22572);
or I_15587 (I267350,I267597,I267848);
nor I_15588 (I267341,I267730,I267848);
or I_15589 (I267344,I267464,I267848);
DFFARX1 I_15590 (I267848,I2859,I267370,I267362,);
not I_15591 (I267948,I2866);
DFFARX1 I_15592 (I544907,I2859,I267948,I267974,);
not I_15593 (I267982,I267974);
nand I_15594 (I267999,I544892,I544880);
and I_15595 (I268016,I267999,I544895);
DFFARX1 I_15596 (I268016,I2859,I267948,I268042,);
not I_15597 (I268050,I544880);
DFFARX1 I_15598 (I544898,I2859,I267948,I268076,);
not I_15599 (I268084,I268076);
nor I_15600 (I268101,I268084,I267982);
and I_15601 (I268118,I268101,I544880);
nor I_15602 (I268135,I268084,I268050);
nor I_15603 (I267931,I268042,I268135);
DFFARX1 I_15604 (I544886,I2859,I267948,I268175,);
nor I_15605 (I268183,I268175,I268042);
not I_15606 (I268200,I268183);
not I_15607 (I268217,I268175);
nor I_15608 (I268234,I268217,I268118);
DFFARX1 I_15609 (I268234,I2859,I267948,I267934,);
nand I_15610 (I268265,I544883,I544889);
and I_15611 (I268282,I268265,I544904);
DFFARX1 I_15612 (I268282,I2859,I267948,I268308,);
nor I_15613 (I268316,I268308,I268175);
DFFARX1 I_15614 (I268316,I2859,I267948,I267916,);
nand I_15615 (I268347,I268308,I268217);
nand I_15616 (I267925,I268200,I268347);
not I_15617 (I268378,I268308);
nor I_15618 (I268395,I268378,I268118);
DFFARX1 I_15619 (I268395,I2859,I267948,I267937,);
nor I_15620 (I268426,I544901,I544889);
or I_15621 (I267928,I268175,I268426);
nor I_15622 (I267919,I268308,I268426);
or I_15623 (I267922,I268042,I268426);
DFFARX1 I_15624 (I268426,I2859,I267948,I267940,);
not I_15625 (I268526,I2866);
DFFARX1 I_15626 (I228578,I2859,I268526,I268552,);
not I_15627 (I268560,I268552);
nand I_15628 (I268577,I228593,I228578);
and I_15629 (I268594,I268577,I228581);
DFFARX1 I_15630 (I268594,I2859,I268526,I268620,);
not I_15631 (I268628,I228581);
DFFARX1 I_15632 (I228590,I2859,I268526,I268654,);
not I_15633 (I268662,I268654);
nor I_15634 (I268679,I268662,I268560);
and I_15635 (I268696,I268679,I228581);
nor I_15636 (I268713,I268662,I268628);
nor I_15637 (I268509,I268620,I268713);
DFFARX1 I_15638 (I228584,I2859,I268526,I268753,);
nor I_15639 (I268761,I268753,I268620);
not I_15640 (I268778,I268761);
not I_15641 (I268795,I268753);
nor I_15642 (I268812,I268795,I268696);
DFFARX1 I_15643 (I268812,I2859,I268526,I268512,);
nand I_15644 (I268843,I228587,I228596);
and I_15645 (I268860,I268843,I228602);
DFFARX1 I_15646 (I268860,I2859,I268526,I268886,);
nor I_15647 (I268894,I268886,I268753);
DFFARX1 I_15648 (I268894,I2859,I268526,I268494,);
nand I_15649 (I268925,I268886,I268795);
nand I_15650 (I268503,I268778,I268925);
not I_15651 (I268956,I268886);
nor I_15652 (I268973,I268956,I268696);
DFFARX1 I_15653 (I268973,I2859,I268526,I268515,);
nor I_15654 (I269004,I228599,I228596);
or I_15655 (I268506,I268753,I269004);
nor I_15656 (I268497,I268886,I269004);
or I_15657 (I268500,I268620,I269004);
DFFARX1 I_15658 (I269004,I2859,I268526,I268518,);
not I_15659 (I269104,I2866);
DFFARX1 I_15660 (I130869,I2859,I269104,I269130,);
not I_15661 (I269138,I269130);
nand I_15662 (I269155,I130872,I130848);
and I_15663 (I269172,I269155,I130845);
DFFARX1 I_15664 (I269172,I2859,I269104,I269198,);
not I_15665 (I269206,I130851);
DFFARX1 I_15666 (I130845,I2859,I269104,I269232,);
not I_15667 (I269240,I269232);
nor I_15668 (I269257,I269240,I269138);
and I_15669 (I269274,I269257,I130851);
nor I_15670 (I269291,I269240,I269206);
nor I_15671 (I269087,I269198,I269291);
DFFARX1 I_15672 (I130854,I2859,I269104,I269331,);
nor I_15673 (I269339,I269331,I269198);
not I_15674 (I269356,I269339);
not I_15675 (I269373,I269331);
nor I_15676 (I269390,I269373,I269274);
DFFARX1 I_15677 (I269390,I2859,I269104,I269090,);
nand I_15678 (I269421,I130857,I130866);
and I_15679 (I269438,I269421,I130863);
DFFARX1 I_15680 (I269438,I2859,I269104,I269464,);
nor I_15681 (I269472,I269464,I269331);
DFFARX1 I_15682 (I269472,I2859,I269104,I269072,);
nand I_15683 (I269503,I269464,I269373);
nand I_15684 (I269081,I269356,I269503);
not I_15685 (I269534,I269464);
nor I_15686 (I269551,I269534,I269274);
DFFARX1 I_15687 (I269551,I2859,I269104,I269093,);
nor I_15688 (I269582,I130860,I130866);
or I_15689 (I269084,I269331,I269582);
nor I_15690 (I269075,I269464,I269582);
or I_15691 (I269078,I269198,I269582);
DFFARX1 I_15692 (I269582,I2859,I269104,I269096,);
not I_15693 (I269682,I2866);
DFFARX1 I_15694 (I211918,I2859,I269682,I269708,);
not I_15695 (I269716,I269708);
nand I_15696 (I269733,I211933,I211918);
and I_15697 (I269750,I269733,I211921);
DFFARX1 I_15698 (I269750,I2859,I269682,I269776,);
not I_15699 (I269784,I211921);
DFFARX1 I_15700 (I211930,I2859,I269682,I269810,);
not I_15701 (I269818,I269810);
nor I_15702 (I269835,I269818,I269716);
and I_15703 (I269852,I269835,I211921);
nor I_15704 (I269869,I269818,I269784);
nor I_15705 (I269665,I269776,I269869);
DFFARX1 I_15706 (I211924,I2859,I269682,I269909,);
nor I_15707 (I269917,I269909,I269776);
not I_15708 (I269934,I269917);
not I_15709 (I269951,I269909);
nor I_15710 (I269968,I269951,I269852);
DFFARX1 I_15711 (I269968,I2859,I269682,I269668,);
nand I_15712 (I269999,I211927,I211936);
and I_15713 (I270016,I269999,I211942);
DFFARX1 I_15714 (I270016,I2859,I269682,I270042,);
nor I_15715 (I270050,I270042,I269909);
DFFARX1 I_15716 (I270050,I2859,I269682,I269650,);
nand I_15717 (I270081,I270042,I269951);
nand I_15718 (I269659,I269934,I270081);
not I_15719 (I270112,I270042);
nor I_15720 (I270129,I270112,I269852);
DFFARX1 I_15721 (I270129,I2859,I269682,I269671,);
nor I_15722 (I270160,I211939,I211936);
or I_15723 (I269662,I269909,I270160);
nor I_15724 (I269653,I270042,I270160);
or I_15725 (I269656,I269776,I270160);
DFFARX1 I_15726 (I270160,I2859,I269682,I269674,);
not I_15727 (I270260,I2866);
DFFARX1 I_15728 (I529206,I2859,I270260,I270286,);
not I_15729 (I270294,I270286);
nand I_15730 (I270311,I529230,I529212);
and I_15731 (I270328,I270311,I529218);
DFFARX1 I_15732 (I270328,I2859,I270260,I270354,);
not I_15733 (I270362,I529224);
DFFARX1 I_15734 (I529209,I2859,I270260,I270388,);
not I_15735 (I270396,I270388);
nor I_15736 (I270413,I270396,I270294);
and I_15737 (I270430,I270413,I529224);
nor I_15738 (I270447,I270396,I270362);
nor I_15739 (I270243,I270354,I270447);
DFFARX1 I_15740 (I529221,I2859,I270260,I270487,);
nor I_15741 (I270495,I270487,I270354);
not I_15742 (I270512,I270495);
not I_15743 (I270529,I270487);
nor I_15744 (I270546,I270529,I270430);
DFFARX1 I_15745 (I270546,I2859,I270260,I270246,);
nand I_15746 (I270577,I529227,I529215);
and I_15747 (I270594,I270577,I529209);
DFFARX1 I_15748 (I270594,I2859,I270260,I270620,);
nor I_15749 (I270628,I270620,I270487);
DFFARX1 I_15750 (I270628,I2859,I270260,I270228,);
nand I_15751 (I270659,I270620,I270529);
nand I_15752 (I270237,I270512,I270659);
not I_15753 (I270690,I270620);
nor I_15754 (I270707,I270690,I270430);
DFFARX1 I_15755 (I270707,I2859,I270260,I270249,);
nor I_15756 (I270738,I529206,I529215);
or I_15757 (I270240,I270487,I270738);
nor I_15758 (I270231,I270620,I270738);
or I_15759 (I270234,I270354,I270738);
DFFARX1 I_15760 (I270738,I2859,I270260,I270252,);
not I_15761 (I270838,I2866);
DFFARX1 I_15762 (I511866,I2859,I270838,I270864,);
not I_15763 (I270872,I270864);
nand I_15764 (I270889,I511869,I511878);
and I_15765 (I270906,I270889,I511881);
DFFARX1 I_15766 (I270906,I2859,I270838,I270932,);
not I_15767 (I270940,I511890);
DFFARX1 I_15768 (I511872,I2859,I270838,I270966,);
not I_15769 (I270974,I270966);
nor I_15770 (I270991,I270974,I270872);
and I_15771 (I271008,I270991,I511890);
nor I_15772 (I271025,I270974,I270940);
nor I_15773 (I270821,I270932,I271025);
DFFARX1 I_15774 (I511869,I2859,I270838,I271065,);
nor I_15775 (I271073,I271065,I270932);
not I_15776 (I271090,I271073);
not I_15777 (I271107,I271065);
nor I_15778 (I271124,I271107,I271008);
DFFARX1 I_15779 (I271124,I2859,I270838,I270824,);
nand I_15780 (I271155,I511887,I511866);
and I_15781 (I271172,I271155,I511884);
DFFARX1 I_15782 (I271172,I2859,I270838,I271198,);
nor I_15783 (I271206,I271198,I271065);
DFFARX1 I_15784 (I271206,I2859,I270838,I270806,);
nand I_15785 (I271237,I271198,I271107);
nand I_15786 (I270815,I271090,I271237);
not I_15787 (I271268,I271198);
nor I_15788 (I271285,I271268,I271008);
DFFARX1 I_15789 (I271285,I2859,I270838,I270827,);
nor I_15790 (I271316,I511875,I511866);
or I_15791 (I270818,I271065,I271316);
nor I_15792 (I270809,I271198,I271316);
or I_15793 (I270812,I270932,I271316);
DFFARX1 I_15794 (I271316,I2859,I270838,I270830,);
not I_15795 (I271416,I2866);
DFFARX1 I_15796 (I470302,I2859,I271416,I271442,);
not I_15797 (I271450,I271442);
nand I_15798 (I271467,I470284,I470296);
and I_15799 (I271484,I271467,I470299);
DFFARX1 I_15800 (I271484,I2859,I271416,I271510,);
not I_15801 (I271518,I470293);
DFFARX1 I_15802 (I470290,I2859,I271416,I271544,);
not I_15803 (I271552,I271544);
nor I_15804 (I271569,I271552,I271450);
and I_15805 (I271586,I271569,I470293);
nor I_15806 (I271603,I271552,I271518);
nor I_15807 (I271399,I271510,I271603);
DFFARX1 I_15808 (I470308,I2859,I271416,I271643,);
nor I_15809 (I271651,I271643,I271510);
not I_15810 (I271668,I271651);
not I_15811 (I271685,I271643);
nor I_15812 (I271702,I271685,I271586);
DFFARX1 I_15813 (I271702,I2859,I271416,I271402,);
nand I_15814 (I271733,I470287,I470287);
and I_15815 (I271750,I271733,I470284);
DFFARX1 I_15816 (I271750,I2859,I271416,I271776,);
nor I_15817 (I271784,I271776,I271643);
DFFARX1 I_15818 (I271784,I2859,I271416,I271384,);
nand I_15819 (I271815,I271776,I271685);
nand I_15820 (I271393,I271668,I271815);
not I_15821 (I271846,I271776);
nor I_15822 (I271863,I271846,I271586);
DFFARX1 I_15823 (I271863,I2859,I271416,I271405,);
nor I_15824 (I271894,I470305,I470287);
or I_15825 (I271396,I271643,I271894);
nor I_15826 (I271387,I271776,I271894);
or I_15827 (I271390,I271510,I271894);
DFFARX1 I_15828 (I271894,I2859,I271416,I271408,);
not I_15829 (I271994,I2866);
DFFARX1 I_15830 (I238438,I2859,I271994,I272020,);
not I_15831 (I272028,I272020);
nand I_15832 (I272045,I238447,I238456);
and I_15833 (I272062,I272045,I238462);
DFFARX1 I_15834 (I272062,I2859,I271994,I272088,);
not I_15835 (I272096,I238459);
DFFARX1 I_15836 (I238444,I2859,I271994,I272122,);
not I_15837 (I272130,I272122);
nor I_15838 (I272147,I272130,I272028);
and I_15839 (I272164,I272147,I238459);
nor I_15840 (I272181,I272130,I272096);
nor I_15841 (I271977,I272088,I272181);
DFFARX1 I_15842 (I238453,I2859,I271994,I272221,);
nor I_15843 (I272229,I272221,I272088);
not I_15844 (I272246,I272229);
not I_15845 (I272263,I272221);
nor I_15846 (I272280,I272263,I272164);
DFFARX1 I_15847 (I272280,I2859,I271994,I271980,);
nand I_15848 (I272311,I238450,I238441);
and I_15849 (I272328,I272311,I238438);
DFFARX1 I_15850 (I272328,I2859,I271994,I272354,);
nor I_15851 (I272362,I272354,I272221);
DFFARX1 I_15852 (I272362,I2859,I271994,I271962,);
nand I_15853 (I272393,I272354,I272263);
nand I_15854 (I271971,I272246,I272393);
not I_15855 (I272424,I272354);
nor I_15856 (I272441,I272424,I272164);
DFFARX1 I_15857 (I272441,I2859,I271994,I271983,);
nor I_15858 (I272472,I238441,I238441);
or I_15859 (I271974,I272221,I272472);
nor I_15860 (I271965,I272354,I272472);
or I_15861 (I271968,I272088,I272472);
DFFARX1 I_15862 (I272472,I2859,I271994,I271986,);
not I_15863 (I272572,I2866);
DFFARX1 I_15864 (I107681,I2859,I272572,I272598,);
not I_15865 (I272606,I272598);
nand I_15866 (I272623,I107684,I107660);
and I_15867 (I272640,I272623,I107657);
DFFARX1 I_15868 (I272640,I2859,I272572,I272666,);
not I_15869 (I272674,I107663);
DFFARX1 I_15870 (I107657,I2859,I272572,I272700,);
not I_15871 (I272708,I272700);
nor I_15872 (I272725,I272708,I272606);
and I_15873 (I272742,I272725,I107663);
nor I_15874 (I272759,I272708,I272674);
nor I_15875 (I272555,I272666,I272759);
DFFARX1 I_15876 (I107666,I2859,I272572,I272799,);
nor I_15877 (I272807,I272799,I272666);
not I_15878 (I272824,I272807);
not I_15879 (I272841,I272799);
nor I_15880 (I272858,I272841,I272742);
DFFARX1 I_15881 (I272858,I2859,I272572,I272558,);
nand I_15882 (I272889,I107669,I107678);
and I_15883 (I272906,I272889,I107675);
DFFARX1 I_15884 (I272906,I2859,I272572,I272932,);
nor I_15885 (I272940,I272932,I272799);
DFFARX1 I_15886 (I272940,I2859,I272572,I272540,);
nand I_15887 (I272971,I272932,I272841);
nand I_15888 (I272549,I272824,I272971);
not I_15889 (I273002,I272932);
nor I_15890 (I273019,I273002,I272742);
DFFARX1 I_15891 (I273019,I2859,I272572,I272561,);
nor I_15892 (I273050,I107672,I107678);
or I_15893 (I272552,I272799,I273050);
nor I_15894 (I272543,I272932,I273050);
or I_15895 (I272546,I272666,I273050);
DFFARX1 I_15896 (I273050,I2859,I272572,I272564,);
not I_15897 (I273150,I2866);
DFFARX1 I_15898 (I481284,I2859,I273150,I273176,);
not I_15899 (I273184,I273176);
nand I_15900 (I273201,I481266,I481278);
and I_15901 (I273218,I273201,I481281);
DFFARX1 I_15902 (I273218,I2859,I273150,I273244,);
not I_15903 (I273252,I481275);
DFFARX1 I_15904 (I481272,I2859,I273150,I273278,);
not I_15905 (I273286,I273278);
nor I_15906 (I273303,I273286,I273184);
and I_15907 (I273320,I273303,I481275);
nor I_15908 (I273337,I273286,I273252);
nor I_15909 (I273133,I273244,I273337);
DFFARX1 I_15910 (I481290,I2859,I273150,I273377,);
nor I_15911 (I273385,I273377,I273244);
not I_15912 (I273402,I273385);
not I_15913 (I273419,I273377);
nor I_15914 (I273436,I273419,I273320);
DFFARX1 I_15915 (I273436,I2859,I273150,I273136,);
nand I_15916 (I273467,I481269,I481269);
and I_15917 (I273484,I273467,I481266);
DFFARX1 I_15918 (I273484,I2859,I273150,I273510,);
nor I_15919 (I273518,I273510,I273377);
DFFARX1 I_15920 (I273518,I2859,I273150,I273118,);
nand I_15921 (I273549,I273510,I273419);
nand I_15922 (I273127,I273402,I273549);
not I_15923 (I273580,I273510);
nor I_15924 (I273597,I273580,I273320);
DFFARX1 I_15925 (I273597,I2859,I273150,I273139,);
nor I_15926 (I273628,I481287,I481269);
or I_15927 (I273130,I273377,I273628);
nor I_15928 (I273121,I273510,I273628);
or I_15929 (I273124,I273244,I273628);
DFFARX1 I_15930 (I273628,I2859,I273150,I273142,);
not I_15931 (I273728,I2866);
DFFARX1 I_15932 (I257512,I2859,I273728,I273754,);
not I_15933 (I273762,I273754);
nand I_15934 (I273779,I257521,I257530);
and I_15935 (I273796,I273779,I257536);
DFFARX1 I_15936 (I273796,I2859,I273728,I273822,);
not I_15937 (I273830,I257533);
DFFARX1 I_15938 (I257518,I2859,I273728,I273856,);
not I_15939 (I273864,I273856);
nor I_15940 (I273881,I273864,I273762);
and I_15941 (I273898,I273881,I257533);
nor I_15942 (I273915,I273864,I273830);
nor I_15943 (I273711,I273822,I273915);
DFFARX1 I_15944 (I257527,I2859,I273728,I273955,);
nor I_15945 (I273963,I273955,I273822);
not I_15946 (I273980,I273963);
not I_15947 (I273997,I273955);
nor I_15948 (I274014,I273997,I273898);
DFFARX1 I_15949 (I274014,I2859,I273728,I273714,);
nand I_15950 (I274045,I257524,I257515);
and I_15951 (I274062,I274045,I257512);
DFFARX1 I_15952 (I274062,I2859,I273728,I274088,);
nor I_15953 (I274096,I274088,I273955);
DFFARX1 I_15954 (I274096,I2859,I273728,I273696,);
nand I_15955 (I274127,I274088,I273997);
nand I_15956 (I273705,I273980,I274127);
not I_15957 (I274158,I274088);
nor I_15958 (I274175,I274158,I273898);
DFFARX1 I_15959 (I274175,I2859,I273728,I273717,);
nor I_15960 (I274206,I257515,I257515);
or I_15961 (I273708,I273955,I274206);
nor I_15962 (I273699,I274088,I274206);
or I_15963 (I273702,I273822,I274206);
DFFARX1 I_15964 (I274206,I2859,I273728,I273720,);
not I_15965 (I274306,I2866);
DFFARX1 I_15966 (I427008,I2859,I274306,I274332,);
not I_15967 (I274340,I274332);
nand I_15968 (I274357,I427005,I427023);
and I_15969 (I274374,I274357,I427020);
DFFARX1 I_15970 (I274374,I2859,I274306,I274400,);
not I_15971 (I274408,I427002);
DFFARX1 I_15972 (I427005,I2859,I274306,I274434,);
not I_15973 (I274442,I274434);
nor I_15974 (I274459,I274442,I274340);
and I_15975 (I274476,I274459,I427002);
nor I_15976 (I274493,I274442,I274408);
nor I_15977 (I274289,I274400,I274493);
DFFARX1 I_15978 (I427014,I2859,I274306,I274533,);
nor I_15979 (I274541,I274533,I274400);
not I_15980 (I274558,I274541);
not I_15981 (I274575,I274533);
nor I_15982 (I274592,I274575,I274476);
DFFARX1 I_15983 (I274592,I2859,I274306,I274292,);
nand I_15984 (I274623,I427017,I427002);
and I_15985 (I274640,I274623,I427008);
DFFARX1 I_15986 (I274640,I2859,I274306,I274666,);
nor I_15987 (I274674,I274666,I274533);
DFFARX1 I_15988 (I274674,I2859,I274306,I274274,);
nand I_15989 (I274705,I274666,I274575);
nand I_15990 (I274283,I274558,I274705);
not I_15991 (I274736,I274666);
nor I_15992 (I274753,I274736,I274476);
DFFARX1 I_15993 (I274753,I2859,I274306,I274295,);
nor I_15994 (I274784,I427011,I427002);
or I_15995 (I274286,I274533,I274784);
nor I_15996 (I274277,I274666,I274784);
or I_15997 (I274280,I274400,I274784);
DFFARX1 I_15998 (I274784,I2859,I274306,I274298,);
not I_15999 (I274884,I2866);
DFFARX1 I_16000 (I75663,I2859,I274884,I274910,);
not I_16001 (I274918,I274910);
nand I_16002 (I274935,I75666,I75687);
and I_16003 (I274952,I274935,I75675);
DFFARX1 I_16004 (I274952,I2859,I274884,I274978,);
not I_16005 (I274986,I75672);
DFFARX1 I_16006 (I75663,I2859,I274884,I275012,);
not I_16007 (I275020,I275012);
nor I_16008 (I275037,I275020,I274918);
and I_16009 (I275054,I275037,I75672);
nor I_16010 (I275071,I275020,I274986);
nor I_16011 (I274867,I274978,I275071);
DFFARX1 I_16012 (I75681,I2859,I274884,I275111,);
nor I_16013 (I275119,I275111,I274978);
not I_16014 (I275136,I275119);
not I_16015 (I275153,I275111);
nor I_16016 (I275170,I275153,I275054);
DFFARX1 I_16017 (I275170,I2859,I274884,I274870,);
nand I_16018 (I275201,I75666,I75669);
and I_16019 (I275218,I275201,I75678);
DFFARX1 I_16020 (I275218,I2859,I274884,I275244,);
nor I_16021 (I275252,I275244,I275111);
DFFARX1 I_16022 (I275252,I2859,I274884,I274852,);
nand I_16023 (I275283,I275244,I275153);
nand I_16024 (I274861,I275136,I275283);
not I_16025 (I275314,I275244);
nor I_16026 (I275331,I275314,I275054);
DFFARX1 I_16027 (I275331,I2859,I274884,I274873,);
nor I_16028 (I275362,I75684,I75669);
or I_16029 (I274864,I275111,I275362);
nor I_16030 (I274855,I275244,I275362);
or I_16031 (I274858,I274978,I275362);
DFFARX1 I_16032 (I275362,I2859,I274884,I274876,);
not I_16033 (I275462,I2866);
DFFARX1 I_16034 (I18368,I2859,I275462,I275488,);
not I_16035 (I275496,I275488);
nand I_16036 (I275513,I18365,I18356);
and I_16037 (I275530,I275513,I18356);
DFFARX1 I_16038 (I275530,I2859,I275462,I275556,);
not I_16039 (I275564,I18359);
DFFARX1 I_16040 (I18374,I2859,I275462,I275590,);
not I_16041 (I275598,I275590);
nor I_16042 (I275615,I275598,I275496);
and I_16043 (I275632,I275615,I18359);
nor I_16044 (I275649,I275598,I275564);
nor I_16045 (I275445,I275556,I275649);
DFFARX1 I_16046 (I18359,I2859,I275462,I275689,);
nor I_16047 (I275697,I275689,I275556);
not I_16048 (I275714,I275697);
not I_16049 (I275731,I275689);
nor I_16050 (I275748,I275731,I275632);
DFFARX1 I_16051 (I275748,I2859,I275462,I275448,);
nand I_16052 (I275779,I18377,I18362);
and I_16053 (I275796,I275779,I18380);
DFFARX1 I_16054 (I275796,I2859,I275462,I275822,);
nor I_16055 (I275830,I275822,I275689);
DFFARX1 I_16056 (I275830,I2859,I275462,I275430,);
nand I_16057 (I275861,I275822,I275731);
nand I_16058 (I275439,I275714,I275861);
not I_16059 (I275892,I275822);
nor I_16060 (I275909,I275892,I275632);
DFFARX1 I_16061 (I275909,I2859,I275462,I275451,);
nor I_16062 (I275940,I18371,I18362);
or I_16063 (I275442,I275689,I275940);
nor I_16064 (I275433,I275822,I275940);
or I_16065 (I275436,I275556,I275940);
DFFARX1 I_16066 (I275940,I2859,I275462,I275454,);
not I_16067 (I276040,I2866);
DFFARX1 I_16068 (I211323,I2859,I276040,I276066,);
not I_16069 (I276074,I276066);
nand I_16070 (I276091,I211338,I211323);
and I_16071 (I276108,I276091,I211326);
DFFARX1 I_16072 (I276108,I2859,I276040,I276134,);
not I_16073 (I276142,I211326);
DFFARX1 I_16074 (I211335,I2859,I276040,I276168,);
not I_16075 (I276176,I276168);
nor I_16076 (I276193,I276176,I276074);
and I_16077 (I276210,I276193,I211326);
nor I_16078 (I276227,I276176,I276142);
nor I_16079 (I276023,I276134,I276227);
DFFARX1 I_16080 (I211329,I2859,I276040,I276267,);
nor I_16081 (I276275,I276267,I276134);
not I_16082 (I276292,I276275);
not I_16083 (I276309,I276267);
nor I_16084 (I276326,I276309,I276210);
DFFARX1 I_16085 (I276326,I2859,I276040,I276026,);
nand I_16086 (I276357,I211332,I211341);
and I_16087 (I276374,I276357,I211347);
DFFARX1 I_16088 (I276374,I2859,I276040,I276400,);
nor I_16089 (I276408,I276400,I276267);
DFFARX1 I_16090 (I276408,I2859,I276040,I276008,);
nand I_16091 (I276439,I276400,I276309);
nand I_16092 (I276017,I276292,I276439);
not I_16093 (I276470,I276400);
nor I_16094 (I276487,I276470,I276210);
DFFARX1 I_16095 (I276487,I2859,I276040,I276029,);
nor I_16096 (I276518,I211344,I211341);
or I_16097 (I276020,I276267,I276518);
nor I_16098 (I276011,I276400,I276518);
or I_16099 (I276014,I276134,I276518);
DFFARX1 I_16100 (I276518,I2859,I276040,I276032,);
not I_16101 (I276618,I2866);
DFFARX1 I_16102 (I206436,I2859,I276618,I276644,);
not I_16103 (I276652,I276644);
nand I_16104 (I276669,I206427,I206445);
and I_16105 (I276686,I276669,I206448);
DFFARX1 I_16106 (I276686,I2859,I276618,I276712,);
not I_16107 (I276720,I206442);
DFFARX1 I_16108 (I206430,I2859,I276618,I276746,);
not I_16109 (I276754,I276746);
nor I_16110 (I276771,I276754,I276652);
and I_16111 (I276788,I276771,I206442);
nor I_16112 (I276805,I276754,I276720);
nor I_16113 (I276601,I276712,I276805);
DFFARX1 I_16114 (I206439,I2859,I276618,I276845,);
nor I_16115 (I276853,I276845,I276712);
not I_16116 (I276870,I276853);
not I_16117 (I276887,I276845);
nor I_16118 (I276904,I276887,I276788);
DFFARX1 I_16119 (I276904,I2859,I276618,I276604,);
nand I_16120 (I276935,I206454,I206451);
and I_16121 (I276952,I276935,I206433);
DFFARX1 I_16122 (I276952,I2859,I276618,I276978,);
nor I_16123 (I276986,I276978,I276845);
DFFARX1 I_16124 (I276986,I2859,I276618,I276586,);
nand I_16125 (I277017,I276978,I276887);
nand I_16126 (I276595,I276870,I277017);
not I_16127 (I277048,I276978);
nor I_16128 (I277065,I277048,I276788);
DFFARX1 I_16129 (I277065,I2859,I276618,I276607,);
nor I_16130 (I277096,I206427,I206451);
or I_16131 (I276598,I276845,I277096);
nor I_16132 (I276589,I276978,I277096);
or I_16133 (I276592,I276712,I277096);
DFFARX1 I_16134 (I277096,I2859,I276618,I276610,);
not I_16135 (I277196,I2866);
DFFARX1 I_16136 (I522270,I2859,I277196,I277222,);
not I_16137 (I277230,I277222);
nand I_16138 (I277247,I522294,I522276);
and I_16139 (I277264,I277247,I522282);
DFFARX1 I_16140 (I277264,I2859,I277196,I277290,);
not I_16141 (I277298,I522288);
DFFARX1 I_16142 (I522273,I2859,I277196,I277324,);
not I_16143 (I277332,I277324);
nor I_16144 (I277349,I277332,I277230);
and I_16145 (I277366,I277349,I522288);
nor I_16146 (I277383,I277332,I277298);
nor I_16147 (I277179,I277290,I277383);
DFFARX1 I_16148 (I522285,I2859,I277196,I277423,);
nor I_16149 (I277431,I277423,I277290);
not I_16150 (I277448,I277431);
not I_16151 (I277465,I277423);
nor I_16152 (I277482,I277465,I277366);
DFFARX1 I_16153 (I277482,I2859,I277196,I277182,);
nand I_16154 (I277513,I522291,I522279);
and I_16155 (I277530,I277513,I522273);
DFFARX1 I_16156 (I277530,I2859,I277196,I277556,);
nor I_16157 (I277564,I277556,I277423);
DFFARX1 I_16158 (I277564,I2859,I277196,I277164,);
nand I_16159 (I277595,I277556,I277465);
nand I_16160 (I277173,I277448,I277595);
not I_16161 (I277626,I277556);
nor I_16162 (I277643,I277626,I277366);
DFFARX1 I_16163 (I277643,I2859,I277196,I277185,);
nor I_16164 (I277674,I522270,I522279);
or I_16165 (I277176,I277423,I277674);
nor I_16166 (I277167,I277556,I277674);
or I_16167 (I277170,I277290,I277674);
DFFARX1 I_16168 (I277674,I2859,I277196,I277188,);
not I_16169 (I277774,I2866);
DFFARX1 I_16170 (I386107,I2859,I277774,I277800,);
not I_16171 (I277808,I277800);
nand I_16172 (I277825,I386083,I386098);
and I_16173 (I277842,I277825,I386110);
DFFARX1 I_16174 (I277842,I2859,I277774,I277868,);
not I_16175 (I277876,I386095);
DFFARX1 I_16176 (I386086,I2859,I277774,I277902,);
not I_16177 (I277910,I277902);
nor I_16178 (I277927,I277910,I277808);
and I_16179 (I277944,I277927,I386095);
nor I_16180 (I277961,I277910,I277876);
nor I_16181 (I277757,I277868,I277961);
DFFARX1 I_16182 (I386083,I2859,I277774,I278001,);
nor I_16183 (I278009,I278001,I277868);
not I_16184 (I278026,I278009);
not I_16185 (I278043,I278001);
nor I_16186 (I278060,I278043,I277944);
DFFARX1 I_16187 (I278060,I2859,I277774,I277760,);
nand I_16188 (I278091,I386101,I386092);
and I_16189 (I278108,I278091,I386104);
DFFARX1 I_16190 (I278108,I2859,I277774,I278134,);
nor I_16191 (I278142,I278134,I278001);
DFFARX1 I_16192 (I278142,I2859,I277774,I277742,);
nand I_16193 (I278173,I278134,I278043);
nand I_16194 (I277751,I278026,I278173);
not I_16195 (I278204,I278134);
nor I_16196 (I278221,I278204,I277944);
DFFARX1 I_16197 (I278221,I2859,I277774,I277763,);
nor I_16198 (I278252,I386089,I386092);
or I_16199 (I277754,I278001,I278252);
nor I_16200 (I277745,I278134,I278252);
or I_16201 (I277748,I277868,I278252);
DFFARX1 I_16202 (I278252,I2859,I277774,I277766,);
not I_16203 (I278352,I2866);
DFFARX1 I_16204 (I182500,I2859,I278352,I278378,);
not I_16205 (I278386,I278378);
nand I_16206 (I278403,I182491,I182509);
and I_16207 (I278420,I278403,I182512);
DFFARX1 I_16208 (I278420,I2859,I278352,I278446,);
not I_16209 (I278454,I182506);
DFFARX1 I_16210 (I182494,I2859,I278352,I278480,);
not I_16211 (I278488,I278480);
nor I_16212 (I278505,I278488,I278386);
and I_16213 (I278522,I278505,I182506);
nor I_16214 (I278539,I278488,I278454);
nor I_16215 (I278335,I278446,I278539);
DFFARX1 I_16216 (I182503,I2859,I278352,I278579,);
nor I_16217 (I278587,I278579,I278446);
not I_16218 (I278604,I278587);
not I_16219 (I278621,I278579);
nor I_16220 (I278638,I278621,I278522);
DFFARX1 I_16221 (I278638,I2859,I278352,I278338,);
nand I_16222 (I278669,I182518,I182515);
and I_16223 (I278686,I278669,I182497);
DFFARX1 I_16224 (I278686,I2859,I278352,I278712,);
nor I_16225 (I278720,I278712,I278579);
DFFARX1 I_16226 (I278720,I2859,I278352,I278320,);
nand I_16227 (I278751,I278712,I278621);
nand I_16228 (I278329,I278604,I278751);
not I_16229 (I278782,I278712);
nor I_16230 (I278799,I278782,I278522);
DFFARX1 I_16231 (I278799,I2859,I278352,I278341,);
nor I_16232 (I278830,I182491,I182515);
or I_16233 (I278332,I278579,I278830);
nor I_16234 (I278323,I278712,I278830);
or I_16235 (I278326,I278446,I278830);
DFFARX1 I_16236 (I278830,I2859,I278352,I278344,);
not I_16237 (I278930,I2866);
DFFARX1 I_16238 (I222628,I2859,I278930,I278956,);
not I_16239 (I278964,I278956);
nand I_16240 (I278981,I222643,I222628);
and I_16241 (I278998,I278981,I222631);
DFFARX1 I_16242 (I278998,I2859,I278930,I279024,);
not I_16243 (I279032,I222631);
DFFARX1 I_16244 (I222640,I2859,I278930,I279058,);
not I_16245 (I279066,I279058);
nor I_16246 (I279083,I279066,I278964);
and I_16247 (I279100,I279083,I222631);
nor I_16248 (I279117,I279066,I279032);
nor I_16249 (I278913,I279024,I279117);
DFFARX1 I_16250 (I222634,I2859,I278930,I279157,);
nor I_16251 (I279165,I279157,I279024);
not I_16252 (I279182,I279165);
not I_16253 (I279199,I279157);
nor I_16254 (I279216,I279199,I279100);
DFFARX1 I_16255 (I279216,I2859,I278930,I278916,);
nand I_16256 (I279247,I222637,I222646);
and I_16257 (I279264,I279247,I222652);
DFFARX1 I_16258 (I279264,I2859,I278930,I279290,);
nor I_16259 (I279298,I279290,I279157);
DFFARX1 I_16260 (I279298,I2859,I278930,I278898,);
nand I_16261 (I279329,I279290,I279199);
nand I_16262 (I278907,I279182,I279329);
not I_16263 (I279360,I279290);
nor I_16264 (I279377,I279360,I279100);
DFFARX1 I_16265 (I279377,I2859,I278930,I278919,);
nor I_16266 (I279408,I222649,I222646);
or I_16267 (I278910,I279157,I279408);
nor I_16268 (I278901,I279290,I279408);
or I_16269 (I278904,I279024,I279408);
DFFARX1 I_16270 (I279408,I2859,I278930,I278922,);
not I_16271 (I279508,I2866);
DFFARX1 I_16272 (I201540,I2859,I279508,I279534,);
not I_16273 (I279542,I279534);
nand I_16274 (I279559,I201531,I201549);
and I_16275 (I279576,I279559,I201552);
DFFARX1 I_16276 (I279576,I2859,I279508,I279602,);
not I_16277 (I279610,I201546);
DFFARX1 I_16278 (I201534,I2859,I279508,I279636,);
not I_16279 (I279644,I279636);
nor I_16280 (I279661,I279644,I279542);
and I_16281 (I279678,I279661,I201546);
nor I_16282 (I279695,I279644,I279610);
nor I_16283 (I279491,I279602,I279695);
DFFARX1 I_16284 (I201543,I2859,I279508,I279735,);
nor I_16285 (I279743,I279735,I279602);
not I_16286 (I279760,I279743);
not I_16287 (I279777,I279735);
nor I_16288 (I279794,I279777,I279678);
DFFARX1 I_16289 (I279794,I2859,I279508,I279494,);
nand I_16290 (I279825,I201558,I201555);
and I_16291 (I279842,I279825,I201537);
DFFARX1 I_16292 (I279842,I2859,I279508,I279868,);
nor I_16293 (I279876,I279868,I279735);
DFFARX1 I_16294 (I279876,I2859,I279508,I279476,);
nand I_16295 (I279907,I279868,I279777);
nand I_16296 (I279485,I279760,I279907);
not I_16297 (I279938,I279868);
nor I_16298 (I279955,I279938,I279678);
DFFARX1 I_16299 (I279955,I2859,I279508,I279497,);
nor I_16300 (I279986,I201531,I201555);
or I_16301 (I279488,I279735,I279986);
nor I_16302 (I279479,I279868,I279986);
or I_16303 (I279482,I279602,I279986);
DFFARX1 I_16304 (I279986,I2859,I279508,I279500,);
not I_16305 (I280086,I2866);
DFFARX1 I_16306 (I179236,I2859,I280086,I280112,);
not I_16307 (I280120,I280112);
nand I_16308 (I280137,I179227,I179245);
and I_16309 (I280154,I280137,I179248);
DFFARX1 I_16310 (I280154,I2859,I280086,I280180,);
not I_16311 (I280188,I179242);
DFFARX1 I_16312 (I179230,I2859,I280086,I280214,);
not I_16313 (I280222,I280214);
nor I_16314 (I280239,I280222,I280120);
and I_16315 (I280256,I280239,I179242);
nor I_16316 (I280273,I280222,I280188);
nor I_16317 (I280069,I280180,I280273);
DFFARX1 I_16318 (I179239,I2859,I280086,I280313,);
nor I_16319 (I280321,I280313,I280180);
not I_16320 (I280338,I280321);
not I_16321 (I280355,I280313);
nor I_16322 (I280372,I280355,I280256);
DFFARX1 I_16323 (I280372,I2859,I280086,I280072,);
nand I_16324 (I280403,I179254,I179251);
and I_16325 (I280420,I280403,I179233);
DFFARX1 I_16326 (I280420,I2859,I280086,I280446,);
nor I_16327 (I280454,I280446,I280313);
DFFARX1 I_16328 (I280454,I2859,I280086,I280054,);
nand I_16329 (I280485,I280446,I280355);
nand I_16330 (I280063,I280338,I280485);
not I_16331 (I280516,I280446);
nor I_16332 (I280533,I280516,I280256);
DFFARX1 I_16333 (I280533,I2859,I280086,I280075,);
nor I_16334 (I280564,I179227,I179251);
or I_16335 (I280066,I280313,I280564);
nor I_16336 (I280057,I280446,I280564);
or I_16337 (I280060,I280180,I280564);
DFFARX1 I_16338 (I280564,I2859,I280086,I280078,);
not I_16339 (I280664,I2866);
DFFARX1 I_16340 (I437106,I2859,I280664,I280690,);
not I_16341 (I280698,I280690);
nand I_16342 (I280715,I437103,I437121);
and I_16343 (I280732,I280715,I437118);
DFFARX1 I_16344 (I280732,I2859,I280664,I280758,);
not I_16345 (I280766,I437100);
DFFARX1 I_16346 (I437103,I2859,I280664,I280792,);
not I_16347 (I280800,I280792);
nor I_16348 (I280817,I280800,I280698);
and I_16349 (I280834,I280817,I437100);
nor I_16350 (I280851,I280800,I280766);
nor I_16351 (I280647,I280758,I280851);
DFFARX1 I_16352 (I437112,I2859,I280664,I280891,);
nor I_16353 (I280899,I280891,I280758);
not I_16354 (I280916,I280899);
not I_16355 (I280933,I280891);
nor I_16356 (I280950,I280933,I280834);
DFFARX1 I_16357 (I280950,I2859,I280664,I280650,);
nand I_16358 (I280981,I437115,I437100);
and I_16359 (I280998,I280981,I437106);
DFFARX1 I_16360 (I280998,I2859,I280664,I281024,);
nor I_16361 (I281032,I281024,I280891);
DFFARX1 I_16362 (I281032,I2859,I280664,I280632,);
nand I_16363 (I281063,I281024,I280933);
nand I_16364 (I280641,I280916,I281063);
not I_16365 (I281094,I281024);
nor I_16366 (I281111,I281094,I280834);
DFFARX1 I_16367 (I281111,I2859,I280664,I280653,);
nor I_16368 (I281142,I437109,I437100);
or I_16369 (I280644,I280891,I281142);
nor I_16370 (I280635,I281024,I281142);
or I_16371 (I280638,I280758,I281142);
DFFARX1 I_16372 (I281142,I2859,I280664,I280656,);
not I_16373 (I281242,I2866);
DFFARX1 I_16374 (I105413,I2859,I281242,I281268,);
not I_16375 (I281276,I281268);
nand I_16376 (I281293,I105416,I105437);
and I_16377 (I281310,I281293,I105425);
DFFARX1 I_16378 (I281310,I2859,I281242,I281336,);
not I_16379 (I281344,I105422);
DFFARX1 I_16380 (I105413,I2859,I281242,I281370,);
not I_16381 (I281378,I281370);
nor I_16382 (I281395,I281378,I281276);
and I_16383 (I281412,I281395,I105422);
nor I_16384 (I281429,I281378,I281344);
nor I_16385 (I281225,I281336,I281429);
DFFARX1 I_16386 (I105431,I2859,I281242,I281469,);
nor I_16387 (I281477,I281469,I281336);
not I_16388 (I281494,I281477);
not I_16389 (I281511,I281469);
nor I_16390 (I281528,I281511,I281412);
DFFARX1 I_16391 (I281528,I2859,I281242,I281228,);
nand I_16392 (I281559,I105416,I105419);
and I_16393 (I281576,I281559,I105428);
DFFARX1 I_16394 (I281576,I2859,I281242,I281602,);
nor I_16395 (I281610,I281602,I281469);
DFFARX1 I_16396 (I281610,I2859,I281242,I281210,);
nand I_16397 (I281641,I281602,I281511);
nand I_16398 (I281219,I281494,I281641);
not I_16399 (I281672,I281602);
nor I_16400 (I281689,I281672,I281412);
DFFARX1 I_16401 (I281689,I2859,I281242,I281231,);
nor I_16402 (I281720,I105434,I105419);
or I_16403 (I281222,I281469,I281720);
nor I_16404 (I281213,I281602,I281720);
or I_16405 (I281216,I281336,I281720);
DFFARX1 I_16406 (I281720,I2859,I281242,I281234,);
not I_16407 (I281820,I2866);
DFFARX1 I_16408 (I36277,I2859,I281820,I281846,);
not I_16409 (I281854,I281846);
nand I_16410 (I281871,I36286,I36295);
and I_16411 (I281888,I281871,I36274);
DFFARX1 I_16412 (I281888,I2859,I281820,I281914,);
not I_16413 (I281922,I36277);
DFFARX1 I_16414 (I36292,I2859,I281820,I281948,);
not I_16415 (I281956,I281948);
nor I_16416 (I281973,I281956,I281854);
and I_16417 (I281990,I281973,I36277);
nor I_16418 (I282007,I281956,I281922);
nor I_16419 (I281803,I281914,I282007);
DFFARX1 I_16420 (I36283,I2859,I281820,I282047,);
nor I_16421 (I282055,I282047,I281914);
not I_16422 (I282072,I282055);
not I_16423 (I282089,I282047);
nor I_16424 (I282106,I282089,I281990);
DFFARX1 I_16425 (I282106,I2859,I281820,I281806,);
nand I_16426 (I282137,I36298,I36274);
and I_16427 (I282154,I282137,I36280);
DFFARX1 I_16428 (I282154,I2859,I281820,I282180,);
nor I_16429 (I282188,I282180,I282047);
DFFARX1 I_16430 (I282188,I2859,I281820,I281788,);
nand I_16431 (I282219,I282180,I282089);
nand I_16432 (I281797,I282072,I282219);
not I_16433 (I282250,I282180);
nor I_16434 (I282267,I282250,I281990);
DFFARX1 I_16435 (I282267,I2859,I281820,I281809,);
nor I_16436 (I282298,I36289,I36274);
or I_16437 (I281800,I282047,I282298);
nor I_16438 (I281791,I282180,I282298);
or I_16439 (I281794,I281914,I282298);
DFFARX1 I_16440 (I282298,I2859,I281820,I281812,);
not I_16441 (I282398,I2866);
DFFARX1 I_16442 (I362706,I2859,I282398,I282424,);
not I_16443 (I282432,I282424);
nand I_16444 (I282449,I362694,I362712);
and I_16445 (I282466,I282449,I362709);
DFFARX1 I_16446 (I282466,I2859,I282398,I282492,);
not I_16447 (I282500,I362700);
DFFARX1 I_16448 (I362697,I2859,I282398,I282526,);
not I_16449 (I282534,I282526);
nor I_16450 (I282551,I282534,I282432);
and I_16451 (I282568,I282551,I362700);
nor I_16452 (I282585,I282534,I282500);
nor I_16453 (I282381,I282492,I282585);
DFFARX1 I_16454 (I362691,I2859,I282398,I282625,);
nor I_16455 (I282633,I282625,I282492);
not I_16456 (I282650,I282633);
not I_16457 (I282667,I282625);
nor I_16458 (I282684,I282667,I282568);
DFFARX1 I_16459 (I282684,I2859,I282398,I282384,);
nand I_16460 (I282715,I362691,I362694);
and I_16461 (I282732,I282715,I362697);
DFFARX1 I_16462 (I282732,I2859,I282398,I282758,);
nor I_16463 (I282766,I282758,I282625);
DFFARX1 I_16464 (I282766,I2859,I282398,I282366,);
nand I_16465 (I282797,I282758,I282667);
nand I_16466 (I282375,I282650,I282797);
not I_16467 (I282828,I282758);
nor I_16468 (I282845,I282828,I282568);
DFFARX1 I_16469 (I282845,I2859,I282398,I282387,);
nor I_16470 (I282876,I362703,I362694);
or I_16471 (I282378,I282625,I282876);
nor I_16472 (I282369,I282758,I282876);
or I_16473 (I282372,I282492,I282876);
DFFARX1 I_16474 (I282876,I2859,I282398,I282390,);
not I_16475 (I282976,I2866);
DFFARX1 I_16476 (I414531,I2859,I282976,I283002,);
not I_16477 (I283010,I283002);
nand I_16478 (I283027,I414507,I414522);
and I_16479 (I283044,I283027,I414534);
DFFARX1 I_16480 (I283044,I2859,I282976,I283070,);
not I_16481 (I283078,I414519);
DFFARX1 I_16482 (I414510,I2859,I282976,I283104,);
not I_16483 (I283112,I283104);
nor I_16484 (I283129,I283112,I283010);
and I_16485 (I283146,I283129,I414519);
nor I_16486 (I283163,I283112,I283078);
nor I_16487 (I282959,I283070,I283163);
DFFARX1 I_16488 (I414507,I2859,I282976,I283203,);
nor I_16489 (I283211,I283203,I283070);
not I_16490 (I283228,I283211);
not I_16491 (I283245,I283203);
nor I_16492 (I283262,I283245,I283146);
DFFARX1 I_16493 (I283262,I2859,I282976,I282962,);
nand I_16494 (I283293,I414525,I414516);
and I_16495 (I283310,I283293,I414528);
DFFARX1 I_16496 (I283310,I2859,I282976,I283336,);
nor I_16497 (I283344,I283336,I283203);
DFFARX1 I_16498 (I283344,I2859,I282976,I282944,);
nand I_16499 (I283375,I283336,I283245);
nand I_16500 (I282953,I283228,I283375);
not I_16501 (I283406,I283336);
nor I_16502 (I283423,I283406,I283146);
DFFARX1 I_16503 (I283423,I2859,I282976,I282965,);
nor I_16504 (I283454,I414513,I414516);
or I_16505 (I282956,I283203,I283454);
nor I_16506 (I282947,I283336,I283454);
or I_16507 (I282950,I283070,I283454);
DFFARX1 I_16508 (I283454,I2859,I282976,I282968,);
not I_16509 (I283554,I2866);
DFFARX1 I_16510 (I178148,I2859,I283554,I283580,);
not I_16511 (I283588,I283580);
nand I_16512 (I283605,I178139,I178157);
and I_16513 (I283622,I283605,I178160);
DFFARX1 I_16514 (I283622,I2859,I283554,I283648,);
not I_16515 (I283656,I178154);
DFFARX1 I_16516 (I178142,I2859,I283554,I283682,);
not I_16517 (I283690,I283682);
nor I_16518 (I283707,I283690,I283588);
and I_16519 (I283724,I283707,I178154);
nor I_16520 (I283741,I283690,I283656);
nor I_16521 (I283537,I283648,I283741);
DFFARX1 I_16522 (I178151,I2859,I283554,I283781,);
nor I_16523 (I283789,I283781,I283648);
not I_16524 (I283806,I283789);
not I_16525 (I283823,I283781);
nor I_16526 (I283840,I283823,I283724);
DFFARX1 I_16527 (I283840,I2859,I283554,I283540,);
nand I_16528 (I283871,I178166,I178163);
and I_16529 (I283888,I283871,I178145);
DFFARX1 I_16530 (I283888,I2859,I283554,I283914,);
nor I_16531 (I283922,I283914,I283781);
DFFARX1 I_16532 (I283922,I2859,I283554,I283522,);
nand I_16533 (I283953,I283914,I283823);
nand I_16534 (I283531,I283806,I283953);
not I_16535 (I283984,I283914);
nor I_16536 (I284001,I283984,I283724);
DFFARX1 I_16537 (I284001,I2859,I283554,I283543,);
nor I_16538 (I284032,I178139,I178163);
or I_16539 (I283534,I283781,I284032);
nor I_16540 (I283525,I283914,I284032);
or I_16541 (I283528,I283648,I284032);
DFFARX1 I_16542 (I284032,I2859,I283554,I283546,);
not I_16543 (I284132,I2866);
DFFARX1 I_16544 (I262136,I2859,I284132,I284158,);
not I_16545 (I284166,I284158);
nand I_16546 (I284183,I262145,I262154);
and I_16547 (I284200,I284183,I262160);
DFFARX1 I_16548 (I284200,I2859,I284132,I284226,);
not I_16549 (I284234,I262157);
DFFARX1 I_16550 (I262142,I2859,I284132,I284260,);
not I_16551 (I284268,I284260);
nor I_16552 (I284285,I284268,I284166);
and I_16553 (I284302,I284285,I262157);
nor I_16554 (I284319,I284268,I284234);
nor I_16555 (I284115,I284226,I284319);
DFFARX1 I_16556 (I262151,I2859,I284132,I284359,);
nor I_16557 (I284367,I284359,I284226);
not I_16558 (I284384,I284367);
not I_16559 (I284401,I284359);
nor I_16560 (I284418,I284401,I284302);
DFFARX1 I_16561 (I284418,I2859,I284132,I284118,);
nand I_16562 (I284449,I262148,I262139);
and I_16563 (I284466,I284449,I262136);
DFFARX1 I_16564 (I284466,I2859,I284132,I284492,);
nor I_16565 (I284500,I284492,I284359);
DFFARX1 I_16566 (I284500,I2859,I284132,I284100,);
nand I_16567 (I284531,I284492,I284401);
nand I_16568 (I284109,I284384,I284531);
not I_16569 (I284562,I284492);
nor I_16570 (I284579,I284562,I284302);
DFFARX1 I_16571 (I284579,I2859,I284132,I284121,);
nor I_16572 (I284610,I262139,I262139);
or I_16573 (I284112,I284359,I284610);
nor I_16574 (I284103,I284492,I284610);
or I_16575 (I284106,I284226,I284610);
DFFARX1 I_16576 (I284610,I2859,I284132,I284124,);
not I_16577 (I284710,I2866);
DFFARX1 I_16578 (I407425,I2859,I284710,I284736,);
not I_16579 (I284744,I284736);
nand I_16580 (I284761,I407401,I407416);
and I_16581 (I284778,I284761,I407428);
DFFARX1 I_16582 (I284778,I2859,I284710,I284804,);
not I_16583 (I284812,I407413);
DFFARX1 I_16584 (I407404,I2859,I284710,I284838,);
not I_16585 (I284846,I284838);
nor I_16586 (I284863,I284846,I284744);
and I_16587 (I284880,I284863,I407413);
nor I_16588 (I284897,I284846,I284812);
nor I_16589 (I284693,I284804,I284897);
DFFARX1 I_16590 (I407401,I2859,I284710,I284937,);
nor I_16591 (I284945,I284937,I284804);
not I_16592 (I284962,I284945);
not I_16593 (I284979,I284937);
nor I_16594 (I284996,I284979,I284880);
DFFARX1 I_16595 (I284996,I2859,I284710,I284696,);
nand I_16596 (I285027,I407419,I407410);
and I_16597 (I285044,I285027,I407422);
DFFARX1 I_16598 (I285044,I2859,I284710,I285070,);
nor I_16599 (I285078,I285070,I284937);
DFFARX1 I_16600 (I285078,I2859,I284710,I284678,);
nand I_16601 (I285109,I285070,I284979);
nand I_16602 (I284687,I284962,I285109);
not I_16603 (I285140,I285070);
nor I_16604 (I285157,I285140,I284880);
DFFARX1 I_16605 (I285157,I2859,I284710,I284699,);
nor I_16606 (I285188,I407407,I407410);
or I_16607 (I284690,I284937,I285188);
nor I_16608 (I284681,I285070,I285188);
or I_16609 (I284684,I284804,I285188);
DFFARX1 I_16610 (I285188,I2859,I284710,I284702,);
not I_16611 (I285288,I2866);
DFFARX1 I_16612 (I202084,I2859,I285288,I285314,);
not I_16613 (I285322,I285314);
nand I_16614 (I285339,I202075,I202093);
and I_16615 (I285356,I285339,I202096);
DFFARX1 I_16616 (I285356,I2859,I285288,I285382,);
not I_16617 (I285390,I202090);
DFFARX1 I_16618 (I202078,I2859,I285288,I285416,);
not I_16619 (I285424,I285416);
nor I_16620 (I285441,I285424,I285322);
and I_16621 (I285458,I285441,I202090);
nor I_16622 (I285475,I285424,I285390);
nor I_16623 (I285271,I285382,I285475);
DFFARX1 I_16624 (I202087,I2859,I285288,I285515,);
nor I_16625 (I285523,I285515,I285382);
not I_16626 (I285540,I285523);
not I_16627 (I285557,I285515);
nor I_16628 (I285574,I285557,I285458);
DFFARX1 I_16629 (I285574,I2859,I285288,I285274,);
nand I_16630 (I285605,I202102,I202099);
and I_16631 (I285622,I285605,I202081);
DFFARX1 I_16632 (I285622,I2859,I285288,I285648,);
nor I_16633 (I285656,I285648,I285515);
DFFARX1 I_16634 (I285656,I2859,I285288,I285256,);
nand I_16635 (I285687,I285648,I285557);
nand I_16636 (I285265,I285540,I285687);
not I_16637 (I285718,I285648);
nor I_16638 (I285735,I285718,I285458);
DFFARX1 I_16639 (I285735,I2859,I285288,I285277,);
nor I_16640 (I285766,I202075,I202099);
or I_16641 (I285268,I285515,I285766);
nor I_16642 (I285259,I285648,I285766);
or I_16643 (I285262,I285382,I285766);
DFFARX1 I_16644 (I285766,I2859,I285288,I285280,);
not I_16645 (I285866,I2866);
DFFARX1 I_16646 (I55249,I2859,I285866,I285892,);
not I_16647 (I285900,I285892);
nand I_16648 (I285917,I55258,I55267);
and I_16649 (I285934,I285917,I55246);
DFFARX1 I_16650 (I285934,I2859,I285866,I285960,);
not I_16651 (I285968,I55249);
DFFARX1 I_16652 (I55264,I2859,I285866,I285994,);
not I_16653 (I286002,I285994);
nor I_16654 (I286019,I286002,I285900);
and I_16655 (I286036,I286019,I55249);
nor I_16656 (I286053,I286002,I285968);
nor I_16657 (I285849,I285960,I286053);
DFFARX1 I_16658 (I55255,I2859,I285866,I286093,);
nor I_16659 (I286101,I286093,I285960);
not I_16660 (I286118,I286101);
not I_16661 (I286135,I286093);
nor I_16662 (I286152,I286135,I286036);
DFFARX1 I_16663 (I286152,I2859,I285866,I285852,);
nand I_16664 (I286183,I55270,I55246);
and I_16665 (I286200,I286183,I55252);
DFFARX1 I_16666 (I286200,I2859,I285866,I286226,);
nor I_16667 (I286234,I286226,I286093);
DFFARX1 I_16668 (I286234,I2859,I285866,I285834,);
nand I_16669 (I286265,I286226,I286135);
nand I_16670 (I285843,I286118,I286265);
not I_16671 (I286296,I286226);
nor I_16672 (I286313,I286296,I286036);
DFFARX1 I_16673 (I286313,I2859,I285866,I285855,);
nor I_16674 (I286344,I55261,I55246);
or I_16675 (I285846,I286093,I286344);
nor I_16676 (I285837,I286226,I286344);
or I_16677 (I285840,I285960,I286344);
DFFARX1 I_16678 (I286344,I2859,I285866,I285858,);
not I_16679 (I286444,I2866);
DFFARX1 I_16680 (I89943,I2859,I286444,I286470,);
not I_16681 (I286478,I286470);
nand I_16682 (I286495,I89946,I89967);
and I_16683 (I286512,I286495,I89955);
DFFARX1 I_16684 (I286512,I2859,I286444,I286538,);
not I_16685 (I286546,I89952);
DFFARX1 I_16686 (I89943,I2859,I286444,I286572,);
not I_16687 (I286580,I286572);
nor I_16688 (I286597,I286580,I286478);
and I_16689 (I286614,I286597,I89952);
nor I_16690 (I286631,I286580,I286546);
nor I_16691 (I286427,I286538,I286631);
DFFARX1 I_16692 (I89961,I2859,I286444,I286671,);
nor I_16693 (I286679,I286671,I286538);
not I_16694 (I286696,I286679);
not I_16695 (I286713,I286671);
nor I_16696 (I286730,I286713,I286614);
DFFARX1 I_16697 (I286730,I2859,I286444,I286430,);
nand I_16698 (I286761,I89946,I89949);
and I_16699 (I286778,I286761,I89958);
DFFARX1 I_16700 (I286778,I2859,I286444,I286804,);
nor I_16701 (I286812,I286804,I286671);
DFFARX1 I_16702 (I286812,I2859,I286444,I286412,);
nand I_16703 (I286843,I286804,I286713);
nand I_16704 (I286421,I286696,I286843);
not I_16705 (I286874,I286804);
nor I_16706 (I286891,I286874,I286614);
DFFARX1 I_16707 (I286891,I2859,I286444,I286433,);
nor I_16708 (I286922,I89964,I89949);
or I_16709 (I286424,I286671,I286922);
nor I_16710 (I286415,I286804,I286922);
or I_16711 (I286418,I286538,I286922);
DFFARX1 I_16712 (I286922,I2859,I286444,I286436,);
not I_16713 (I287022,I2866);
DFFARX1 I_16714 (I128761,I2859,I287022,I287048,);
not I_16715 (I287056,I287048);
nand I_16716 (I287073,I128764,I128740);
and I_16717 (I287090,I287073,I128737);
DFFARX1 I_16718 (I287090,I2859,I287022,I287116,);
not I_16719 (I287124,I128743);
DFFARX1 I_16720 (I128737,I2859,I287022,I287150,);
not I_16721 (I287158,I287150);
nor I_16722 (I287175,I287158,I287056);
and I_16723 (I287192,I287175,I128743);
nor I_16724 (I287209,I287158,I287124);
nor I_16725 (I287005,I287116,I287209);
DFFARX1 I_16726 (I128746,I2859,I287022,I287249,);
nor I_16727 (I287257,I287249,I287116);
not I_16728 (I287274,I287257);
not I_16729 (I287291,I287249);
nor I_16730 (I287308,I287291,I287192);
DFFARX1 I_16731 (I287308,I2859,I287022,I287008,);
nand I_16732 (I287339,I128749,I128758);
and I_16733 (I287356,I287339,I128755);
DFFARX1 I_16734 (I287356,I2859,I287022,I287382,);
nor I_16735 (I287390,I287382,I287249);
DFFARX1 I_16736 (I287390,I2859,I287022,I286990,);
nand I_16737 (I287421,I287382,I287291);
nand I_16738 (I286999,I287274,I287421);
not I_16739 (I287452,I287382);
nor I_16740 (I287469,I287452,I287192);
DFFARX1 I_16741 (I287469,I2859,I287022,I287011,);
nor I_16742 (I287500,I128752,I128758);
or I_16743 (I287002,I287249,I287500);
nor I_16744 (I286993,I287382,I287500);
or I_16745 (I286996,I287116,I287500);
DFFARX1 I_16746 (I287500,I2859,I287022,I287014,);
not I_16747 (I287600,I2866);
DFFARX1 I_16748 (I88158,I2859,I287600,I287626,);
not I_16749 (I287634,I287626);
nand I_16750 (I287651,I88161,I88182);
and I_16751 (I287668,I287651,I88170);
DFFARX1 I_16752 (I287668,I2859,I287600,I287694,);
not I_16753 (I287702,I88167);
DFFARX1 I_16754 (I88158,I2859,I287600,I287728,);
not I_16755 (I287736,I287728);
nor I_16756 (I287753,I287736,I287634);
and I_16757 (I287770,I287753,I88167);
nor I_16758 (I287787,I287736,I287702);
nor I_16759 (I287583,I287694,I287787);
DFFARX1 I_16760 (I88176,I2859,I287600,I287827,);
nor I_16761 (I287835,I287827,I287694);
not I_16762 (I287852,I287835);
not I_16763 (I287869,I287827);
nor I_16764 (I287886,I287869,I287770);
DFFARX1 I_16765 (I287886,I2859,I287600,I287586,);
nand I_16766 (I287917,I88161,I88164);
and I_16767 (I287934,I287917,I88173);
DFFARX1 I_16768 (I287934,I2859,I287600,I287960,);
nor I_16769 (I287968,I287960,I287827);
DFFARX1 I_16770 (I287968,I2859,I287600,I287568,);
nand I_16771 (I287999,I287960,I287869);
nand I_16772 (I287577,I287852,I287999);
not I_16773 (I288030,I287960);
nor I_16774 (I288047,I288030,I287770);
DFFARX1 I_16775 (I288047,I2859,I287600,I287589,);
nor I_16776 (I288078,I88179,I88164);
or I_16777 (I287580,I287827,I288078);
nor I_16778 (I287571,I287960,I288078);
or I_16779 (I287574,I287694,I288078);
DFFARX1 I_16780 (I288078,I2859,I287600,I287592,);
not I_16781 (I288178,I2866);
DFFARX1 I_16782 (I218463,I2859,I288178,I288204,);
not I_16783 (I288212,I288204);
nand I_16784 (I288229,I218478,I218463);
and I_16785 (I288246,I288229,I218466);
DFFARX1 I_16786 (I288246,I2859,I288178,I288272,);
not I_16787 (I288280,I218466);
DFFARX1 I_16788 (I218475,I2859,I288178,I288306,);
not I_16789 (I288314,I288306);
nor I_16790 (I288331,I288314,I288212);
and I_16791 (I288348,I288331,I218466);
nor I_16792 (I288365,I288314,I288280);
nor I_16793 (I288161,I288272,I288365);
DFFARX1 I_16794 (I218469,I2859,I288178,I288405,);
nor I_16795 (I288413,I288405,I288272);
not I_16796 (I288430,I288413);
not I_16797 (I288447,I288405);
nor I_16798 (I288464,I288447,I288348);
DFFARX1 I_16799 (I288464,I2859,I288178,I288164,);
nand I_16800 (I288495,I218472,I218481);
and I_16801 (I288512,I288495,I218487);
DFFARX1 I_16802 (I288512,I2859,I288178,I288538,);
nor I_16803 (I288546,I288538,I288405);
DFFARX1 I_16804 (I288546,I2859,I288178,I288146,);
nand I_16805 (I288577,I288538,I288447);
nand I_16806 (I288155,I288430,I288577);
not I_16807 (I288608,I288538);
nor I_16808 (I288625,I288608,I288348);
DFFARX1 I_16809 (I288625,I2859,I288178,I288167,);
nor I_16810 (I288656,I218484,I218481);
or I_16811 (I288158,I288405,I288656);
nor I_16812 (I288149,I288538,I288656);
or I_16813 (I288152,I288272,I288656);
DFFARX1 I_16814 (I288656,I2859,I288178,I288170,);
not I_16815 (I288756,I2866);
DFFARX1 I_16816 (I178692,I2859,I288756,I288782,);
not I_16817 (I288790,I288782);
nand I_16818 (I288807,I178683,I178701);
and I_16819 (I288824,I288807,I178704);
DFFARX1 I_16820 (I288824,I2859,I288756,I288850,);
not I_16821 (I288858,I178698);
DFFARX1 I_16822 (I178686,I2859,I288756,I288884,);
not I_16823 (I288892,I288884);
nor I_16824 (I288909,I288892,I288790);
and I_16825 (I288926,I288909,I178698);
nor I_16826 (I288943,I288892,I288858);
nor I_16827 (I288739,I288850,I288943);
DFFARX1 I_16828 (I178695,I2859,I288756,I288983,);
nor I_16829 (I288991,I288983,I288850);
not I_16830 (I289008,I288991);
not I_16831 (I289025,I288983);
nor I_16832 (I289042,I289025,I288926);
DFFARX1 I_16833 (I289042,I2859,I288756,I288742,);
nand I_16834 (I289073,I178710,I178707);
and I_16835 (I289090,I289073,I178689);
DFFARX1 I_16836 (I289090,I2859,I288756,I289116,);
nor I_16837 (I289124,I289116,I288983);
DFFARX1 I_16838 (I289124,I2859,I288756,I288724,);
nand I_16839 (I289155,I289116,I289025);
nand I_16840 (I288733,I289008,I289155);
not I_16841 (I289186,I289116);
nor I_16842 (I289203,I289186,I288926);
DFFARX1 I_16843 (I289203,I2859,I288756,I288745,);
nor I_16844 (I289234,I178683,I178707);
or I_16845 (I288736,I288983,I289234);
nor I_16846 (I288727,I289116,I289234);
or I_16847 (I288730,I288850,I289234);
DFFARX1 I_16848 (I289234,I2859,I288756,I288748,);
not I_16849 (I289334,I2866);
DFFARX1 I_16850 (I254044,I2859,I289334,I289360,);
not I_16851 (I289368,I289360);
nand I_16852 (I289385,I254053,I254062);
and I_16853 (I289402,I289385,I254068);
DFFARX1 I_16854 (I289402,I2859,I289334,I289428,);
not I_16855 (I289436,I254065);
DFFARX1 I_16856 (I254050,I2859,I289334,I289462,);
not I_16857 (I289470,I289462);
nor I_16858 (I289487,I289470,I289368);
and I_16859 (I289504,I289487,I254065);
nor I_16860 (I289521,I289470,I289436);
nor I_16861 (I289317,I289428,I289521);
DFFARX1 I_16862 (I254059,I2859,I289334,I289561,);
nor I_16863 (I289569,I289561,I289428);
not I_16864 (I289586,I289569);
not I_16865 (I289603,I289561);
nor I_16866 (I289620,I289603,I289504);
DFFARX1 I_16867 (I289620,I2859,I289334,I289320,);
nand I_16868 (I289651,I254056,I254047);
and I_16869 (I289668,I289651,I254044);
DFFARX1 I_16870 (I289668,I2859,I289334,I289694,);
nor I_16871 (I289702,I289694,I289561);
DFFARX1 I_16872 (I289702,I2859,I289334,I289302,);
nand I_16873 (I289733,I289694,I289603);
nand I_16874 (I289311,I289586,I289733);
not I_16875 (I289764,I289694);
nor I_16876 (I289781,I289764,I289504);
DFFARX1 I_16877 (I289781,I2859,I289334,I289323,);
nor I_16878 (I289812,I254047,I254047);
or I_16879 (I289314,I289561,I289812);
nor I_16880 (I289305,I289694,I289812);
or I_16881 (I289308,I289428,I289812);
DFFARX1 I_16882 (I289812,I2859,I289334,I289326,);
not I_16883 (I289912,I2866);
DFFARX1 I_16884 (I49452,I2859,I289912,I289938,);
not I_16885 (I289946,I289938);
nand I_16886 (I289963,I49461,I49470);
and I_16887 (I289980,I289963,I49449);
DFFARX1 I_16888 (I289980,I2859,I289912,I290006,);
not I_16889 (I290014,I49452);
DFFARX1 I_16890 (I49467,I2859,I289912,I290040,);
not I_16891 (I290048,I290040);
nor I_16892 (I290065,I290048,I289946);
and I_16893 (I290082,I290065,I49452);
nor I_16894 (I290099,I290048,I290014);
nor I_16895 (I289895,I290006,I290099);
DFFARX1 I_16896 (I49458,I2859,I289912,I290139,);
nor I_16897 (I290147,I290139,I290006);
not I_16898 (I290164,I290147);
not I_16899 (I290181,I290139);
nor I_16900 (I290198,I290181,I290082);
DFFARX1 I_16901 (I290198,I2859,I289912,I289898,);
nand I_16902 (I290229,I49473,I49449);
and I_16903 (I290246,I290229,I49455);
DFFARX1 I_16904 (I290246,I2859,I289912,I290272,);
nor I_16905 (I290280,I290272,I290139);
DFFARX1 I_16906 (I290280,I2859,I289912,I289880,);
nand I_16907 (I290311,I290272,I290181);
nand I_16908 (I289889,I290164,I290311);
not I_16909 (I290342,I290272);
nor I_16910 (I290359,I290342,I290082);
DFFARX1 I_16911 (I290359,I2859,I289912,I289901,);
nor I_16912 (I290390,I49464,I49449);
or I_16913 (I289892,I290139,I290390);
nor I_16914 (I289883,I290272,I290390);
or I_16915 (I289886,I290006,I290390);
DFFARX1 I_16916 (I290390,I2859,I289912,I289904,);
not I_16917 (I290490,I2866);
DFFARX1 I_16918 (I100653,I2859,I290490,I290516,);
not I_16919 (I290524,I290516);
nand I_16920 (I290541,I100656,I100677);
and I_16921 (I290558,I290541,I100665);
DFFARX1 I_16922 (I290558,I2859,I290490,I290584,);
not I_16923 (I290592,I100662);
DFFARX1 I_16924 (I100653,I2859,I290490,I290618,);
not I_16925 (I290626,I290618);
nor I_16926 (I290643,I290626,I290524);
and I_16927 (I290660,I290643,I100662);
nor I_16928 (I290677,I290626,I290592);
nor I_16929 (I290473,I290584,I290677);
DFFARX1 I_16930 (I100671,I2859,I290490,I290717,);
nor I_16931 (I290725,I290717,I290584);
not I_16932 (I290742,I290725);
not I_16933 (I290759,I290717);
nor I_16934 (I290776,I290759,I290660);
DFFARX1 I_16935 (I290776,I2859,I290490,I290476,);
nand I_16936 (I290807,I100656,I100659);
and I_16937 (I290824,I290807,I100668);
DFFARX1 I_16938 (I290824,I2859,I290490,I290850,);
nor I_16939 (I290858,I290850,I290717);
DFFARX1 I_16940 (I290858,I2859,I290490,I290458,);
nand I_16941 (I290889,I290850,I290759);
nand I_16942 (I290467,I290742,I290889);
not I_16943 (I290920,I290850);
nor I_16944 (I290937,I290920,I290660);
DFFARX1 I_16945 (I290937,I2859,I290490,I290479,);
nor I_16946 (I290968,I100674,I100659);
or I_16947 (I290470,I290717,I290968);
nor I_16948 (I290461,I290850,I290968);
or I_16949 (I290464,I290584,I290968);
DFFARX1 I_16950 (I290968,I2859,I290490,I290482,);
not I_16951 (I291068,I2866);
DFFARX1 I_16952 (I92323,I2859,I291068,I291094,);
not I_16953 (I291102,I291094);
nand I_16954 (I291119,I92326,I92347);
and I_16955 (I291136,I291119,I92335);
DFFARX1 I_16956 (I291136,I2859,I291068,I291162,);
not I_16957 (I291170,I92332);
DFFARX1 I_16958 (I92323,I2859,I291068,I291196,);
not I_16959 (I291204,I291196);
nor I_16960 (I291221,I291204,I291102);
and I_16961 (I291238,I291221,I92332);
nor I_16962 (I291255,I291204,I291170);
nor I_16963 (I291051,I291162,I291255);
DFFARX1 I_16964 (I92341,I2859,I291068,I291295,);
nor I_16965 (I291303,I291295,I291162);
not I_16966 (I291320,I291303);
not I_16967 (I291337,I291295);
nor I_16968 (I291354,I291337,I291238);
DFFARX1 I_16969 (I291354,I2859,I291068,I291054,);
nand I_16970 (I291385,I92326,I92329);
and I_16971 (I291402,I291385,I92338);
DFFARX1 I_16972 (I291402,I2859,I291068,I291428,);
nor I_16973 (I291436,I291428,I291295);
DFFARX1 I_16974 (I291436,I2859,I291068,I291036,);
nand I_16975 (I291467,I291428,I291337);
nand I_16976 (I291045,I291320,I291467);
not I_16977 (I291498,I291428);
nor I_16978 (I291515,I291498,I291238);
DFFARX1 I_16979 (I291515,I2859,I291068,I291057,);
nor I_16980 (I291546,I92344,I92329);
or I_16981 (I291048,I291295,I291546);
nor I_16982 (I291039,I291428,I291546);
or I_16983 (I291042,I291162,I291546);
DFFARX1 I_16984 (I291546,I2859,I291068,I291060,);
not I_16985 (I291646,I2866);
DFFARX1 I_16986 (I539552,I2859,I291646,I291672,);
not I_16987 (I291680,I291672);
nand I_16988 (I291697,I539537,I539525);
and I_16989 (I291714,I291697,I539540);
DFFARX1 I_16990 (I291714,I2859,I291646,I291740,);
not I_16991 (I291748,I539525);
DFFARX1 I_16992 (I539543,I2859,I291646,I291774,);
not I_16993 (I291782,I291774);
nor I_16994 (I291799,I291782,I291680);
and I_16995 (I291816,I291799,I539525);
nor I_16996 (I291833,I291782,I291748);
nor I_16997 (I291629,I291740,I291833);
DFFARX1 I_16998 (I539531,I2859,I291646,I291873,);
nor I_16999 (I291881,I291873,I291740);
not I_17000 (I291898,I291881);
not I_17001 (I291915,I291873);
nor I_17002 (I291932,I291915,I291816);
DFFARX1 I_17003 (I291932,I2859,I291646,I291632,);
nand I_17004 (I291963,I539528,I539534);
and I_17005 (I291980,I291963,I539549);
DFFARX1 I_17006 (I291980,I2859,I291646,I292006,);
nor I_17007 (I292014,I292006,I291873);
DFFARX1 I_17008 (I292014,I2859,I291646,I291614,);
nand I_17009 (I292045,I292006,I291915);
nand I_17010 (I291623,I291898,I292045);
not I_17011 (I292076,I292006);
nor I_17012 (I292093,I292076,I291816);
DFFARX1 I_17013 (I292093,I2859,I291646,I291635,);
nor I_17014 (I292124,I539546,I539534);
or I_17015 (I291626,I291873,I292124);
nor I_17016 (I291617,I292006,I292124);
or I_17017 (I291620,I291740,I292124);
DFFARX1 I_17018 (I292124,I2859,I291646,I291638,);
not I_17019 (I292224,I2866);
DFFARX1 I_17020 (I193380,I2859,I292224,I292250,);
not I_17021 (I292258,I292250);
nand I_17022 (I292275,I193371,I193389);
and I_17023 (I292292,I292275,I193392);
DFFARX1 I_17024 (I292292,I2859,I292224,I292318,);
not I_17025 (I292326,I193386);
DFFARX1 I_17026 (I193374,I2859,I292224,I292352,);
not I_17027 (I292360,I292352);
nor I_17028 (I292377,I292360,I292258);
and I_17029 (I292394,I292377,I193386);
nor I_17030 (I292411,I292360,I292326);
nor I_17031 (I292207,I292318,I292411);
DFFARX1 I_17032 (I193383,I2859,I292224,I292451,);
nor I_17033 (I292459,I292451,I292318);
not I_17034 (I292476,I292459);
not I_17035 (I292493,I292451);
nor I_17036 (I292510,I292493,I292394);
DFFARX1 I_17037 (I292510,I2859,I292224,I292210,);
nand I_17038 (I292541,I193398,I193395);
and I_17039 (I292558,I292541,I193377);
DFFARX1 I_17040 (I292558,I2859,I292224,I292584,);
nor I_17041 (I292592,I292584,I292451);
DFFARX1 I_17042 (I292592,I2859,I292224,I292192,);
nand I_17043 (I292623,I292584,I292493);
nand I_17044 (I292201,I292476,I292623);
not I_17045 (I292654,I292584);
nor I_17046 (I292671,I292654,I292394);
DFFARX1 I_17047 (I292671,I2859,I292224,I292213,);
nor I_17048 (I292702,I193371,I193395);
or I_17049 (I292204,I292451,I292702);
nor I_17050 (I292195,I292584,I292702);
or I_17051 (I292198,I292318,I292702);
DFFARX1 I_17052 (I292702,I2859,I292224,I292216,);
not I_17053 (I292802,I2866);
DFFARX1 I_17054 (I372719,I2859,I292802,I292828,);
not I_17055 (I292836,I292828);
nand I_17056 (I292853,I372707,I372725);
and I_17057 (I292870,I292853,I372722);
DFFARX1 I_17058 (I292870,I2859,I292802,I292896,);
not I_17059 (I292904,I372713);
DFFARX1 I_17060 (I372710,I2859,I292802,I292930,);
not I_17061 (I292938,I292930);
nor I_17062 (I292955,I292938,I292836);
and I_17063 (I292972,I292955,I372713);
nor I_17064 (I292989,I292938,I292904);
nor I_17065 (I292785,I292896,I292989);
DFFARX1 I_17066 (I372704,I2859,I292802,I293029,);
nor I_17067 (I293037,I293029,I292896);
not I_17068 (I293054,I293037);
not I_17069 (I293071,I293029);
nor I_17070 (I293088,I293071,I292972);
DFFARX1 I_17071 (I293088,I2859,I292802,I292788,);
nand I_17072 (I293119,I372704,I372707);
and I_17073 (I293136,I293119,I372710);
DFFARX1 I_17074 (I293136,I2859,I292802,I293162,);
nor I_17075 (I293170,I293162,I293029);
DFFARX1 I_17076 (I293170,I2859,I292802,I292770,);
nand I_17077 (I293201,I293162,I293071);
nand I_17078 (I292779,I293054,I293201);
not I_17079 (I293232,I293162);
nor I_17080 (I293249,I293232,I292972);
DFFARX1 I_17081 (I293249,I2859,I292802,I292791,);
nor I_17082 (I293280,I372716,I372707);
or I_17083 (I292782,I293029,I293280);
nor I_17084 (I292773,I293162,I293280);
or I_17085 (I292776,I292896,I293280);
DFFARX1 I_17086 (I293280,I2859,I292802,I292794,);
not I_17087 (I293380,I2866);
DFFARX1 I_17088 (I213108,I2859,I293380,I293406,);
not I_17089 (I293414,I293406);
nand I_17090 (I293431,I213123,I213108);
and I_17091 (I293448,I293431,I213111);
DFFARX1 I_17092 (I293448,I2859,I293380,I293474,);
not I_17093 (I293482,I213111);
DFFARX1 I_17094 (I213120,I2859,I293380,I293508,);
not I_17095 (I293516,I293508);
nor I_17096 (I293533,I293516,I293414);
and I_17097 (I293550,I293533,I213111);
nor I_17098 (I293567,I293516,I293482);
nor I_17099 (I293363,I293474,I293567);
DFFARX1 I_17100 (I213114,I2859,I293380,I293607,);
nor I_17101 (I293615,I293607,I293474);
not I_17102 (I293632,I293615);
not I_17103 (I293649,I293607);
nor I_17104 (I293666,I293649,I293550);
DFFARX1 I_17105 (I293666,I2859,I293380,I293366,);
nand I_17106 (I293697,I213117,I213126);
and I_17107 (I293714,I293697,I213132);
DFFARX1 I_17108 (I293714,I2859,I293380,I293740,);
nor I_17109 (I293748,I293740,I293607);
DFFARX1 I_17110 (I293748,I2859,I293380,I293348,);
nand I_17111 (I293779,I293740,I293649);
nand I_17112 (I293357,I293632,I293779);
not I_17113 (I293810,I293740);
nor I_17114 (I293827,I293810,I293550);
DFFARX1 I_17115 (I293827,I2859,I293380,I293369,);
nor I_17116 (I293858,I213129,I213126);
or I_17117 (I293360,I293607,I293858);
nor I_17118 (I293351,I293740,I293858);
or I_17119 (I293354,I293474,I293858);
DFFARX1 I_17120 (I293858,I2859,I293380,I293372,);
not I_17121 (I293958,I2866);
DFFARX1 I_17122 (I15733,I2859,I293958,I293984,);
not I_17123 (I293992,I293984);
nand I_17124 (I294009,I15730,I15721);
and I_17125 (I294026,I294009,I15721);
DFFARX1 I_17126 (I294026,I2859,I293958,I294052,);
not I_17127 (I294060,I15724);
DFFARX1 I_17128 (I15739,I2859,I293958,I294086,);
not I_17129 (I294094,I294086);
nor I_17130 (I294111,I294094,I293992);
and I_17131 (I294128,I294111,I15724);
nor I_17132 (I294145,I294094,I294060);
nor I_17133 (I293941,I294052,I294145);
DFFARX1 I_17134 (I15724,I2859,I293958,I294185,);
nor I_17135 (I294193,I294185,I294052);
not I_17136 (I294210,I294193);
not I_17137 (I294227,I294185);
nor I_17138 (I294244,I294227,I294128);
DFFARX1 I_17139 (I294244,I2859,I293958,I293944,);
nand I_17140 (I294275,I15742,I15727);
and I_17141 (I294292,I294275,I15745);
DFFARX1 I_17142 (I294292,I2859,I293958,I294318,);
nor I_17143 (I294326,I294318,I294185);
DFFARX1 I_17144 (I294326,I2859,I293958,I293926,);
nand I_17145 (I294357,I294318,I294227);
nand I_17146 (I293935,I294210,I294357);
not I_17147 (I294388,I294318);
nor I_17148 (I294405,I294388,I294128);
DFFARX1 I_17149 (I294405,I2859,I293958,I293947,);
nor I_17150 (I294436,I15736,I15727);
or I_17151 (I293938,I294185,I294436);
nor I_17152 (I293929,I294318,I294436);
or I_17153 (I293932,I294052,I294436);
DFFARX1 I_17154 (I294436,I2859,I293958,I293950,);
not I_17155 (I294536,I2866);
DFFARX1 I_17156 (I28372,I2859,I294536,I294562,);
not I_17157 (I294570,I294562);
nand I_17158 (I294587,I28381,I28390);
and I_17159 (I294604,I294587,I28369);
DFFARX1 I_17160 (I294604,I2859,I294536,I294630,);
not I_17161 (I294638,I28372);
DFFARX1 I_17162 (I28387,I2859,I294536,I294664,);
not I_17163 (I294672,I294664);
nor I_17164 (I294689,I294672,I294570);
and I_17165 (I294706,I294689,I28372);
nor I_17166 (I294723,I294672,I294638);
nor I_17167 (I294519,I294630,I294723);
DFFARX1 I_17168 (I28378,I2859,I294536,I294763,);
nor I_17169 (I294771,I294763,I294630);
not I_17170 (I294788,I294771);
not I_17171 (I294805,I294763);
nor I_17172 (I294822,I294805,I294706);
DFFARX1 I_17173 (I294822,I2859,I294536,I294522,);
nand I_17174 (I294853,I28393,I28369);
and I_17175 (I294870,I294853,I28375);
DFFARX1 I_17176 (I294870,I2859,I294536,I294896,);
nor I_17177 (I294904,I294896,I294763);
DFFARX1 I_17178 (I294904,I2859,I294536,I294504,);
nand I_17179 (I294935,I294896,I294805);
nand I_17180 (I294513,I294788,I294935);
not I_17181 (I294966,I294896);
nor I_17182 (I294983,I294966,I294706);
DFFARX1 I_17183 (I294983,I2859,I294536,I294525,);
nor I_17184 (I295014,I28384,I28369);
or I_17185 (I294516,I294763,I295014);
nor I_17186 (I294507,I294896,I295014);
or I_17187 (I294510,I294630,I295014);
DFFARX1 I_17188 (I295014,I2859,I294536,I294528,);
not I_17189 (I295114,I2866);
DFFARX1 I_17190 (I340045,I2859,I295114,I295140,);
not I_17191 (I295148,I295140);
nand I_17192 (I295165,I340033,I340051);
and I_17193 (I295182,I295165,I340048);
DFFARX1 I_17194 (I295182,I2859,I295114,I295208,);
not I_17195 (I295216,I340039);
DFFARX1 I_17196 (I340036,I2859,I295114,I295242,);
not I_17197 (I295250,I295242);
nor I_17198 (I295267,I295250,I295148);
and I_17199 (I295284,I295267,I340039);
nor I_17200 (I295301,I295250,I295216);
nor I_17201 (I295097,I295208,I295301);
DFFARX1 I_17202 (I340030,I2859,I295114,I295341,);
nor I_17203 (I295349,I295341,I295208);
not I_17204 (I295366,I295349);
not I_17205 (I295383,I295341);
nor I_17206 (I295400,I295383,I295284);
DFFARX1 I_17207 (I295400,I2859,I295114,I295100,);
nand I_17208 (I295431,I340030,I340033);
and I_17209 (I295448,I295431,I340036);
DFFARX1 I_17210 (I295448,I2859,I295114,I295474,);
nor I_17211 (I295482,I295474,I295341);
DFFARX1 I_17212 (I295482,I2859,I295114,I295082,);
nand I_17213 (I295513,I295474,I295383);
nand I_17214 (I295091,I295366,I295513);
not I_17215 (I295544,I295474);
nor I_17216 (I295561,I295544,I295284);
DFFARX1 I_17217 (I295561,I2859,I295114,I295103,);
nor I_17218 (I295592,I340042,I340033);
or I_17219 (I295094,I295341,I295592);
nor I_17220 (I295085,I295474,I295592);
or I_17221 (I295088,I295208,I295592);
DFFARX1 I_17222 (I295592,I2859,I295114,I295106,);
not I_17223 (I295692,I2866);
DFFARX1 I_17224 (I518394,I2859,I295692,I295718,);
not I_17225 (I295726,I295718);
nand I_17226 (I295743,I518397,I518406);
and I_17227 (I295760,I295743,I518409);
DFFARX1 I_17228 (I295760,I2859,I295692,I295786,);
not I_17229 (I295794,I518418);
DFFARX1 I_17230 (I518400,I2859,I295692,I295820,);
not I_17231 (I295828,I295820);
nor I_17232 (I295845,I295828,I295726);
and I_17233 (I295862,I295845,I518418);
nor I_17234 (I295879,I295828,I295794);
nor I_17235 (I295675,I295786,I295879);
DFFARX1 I_17236 (I518397,I2859,I295692,I295919,);
nor I_17237 (I295927,I295919,I295786);
not I_17238 (I295944,I295927);
not I_17239 (I295961,I295919);
nor I_17240 (I295978,I295961,I295862);
DFFARX1 I_17241 (I295978,I2859,I295692,I295678,);
nand I_17242 (I296009,I518415,I518394);
and I_17243 (I296026,I296009,I518412);
DFFARX1 I_17244 (I296026,I2859,I295692,I296052,);
nor I_17245 (I296060,I296052,I295919);
DFFARX1 I_17246 (I296060,I2859,I295692,I295660,);
nand I_17247 (I296091,I296052,I295961);
nand I_17248 (I295669,I295944,I296091);
not I_17249 (I296122,I296052);
nor I_17250 (I296139,I296122,I295862);
DFFARX1 I_17251 (I296139,I2859,I295692,I295681,);
nor I_17252 (I296170,I518403,I518394);
or I_17253 (I295672,I295919,I296170);
nor I_17254 (I295663,I296052,I296170);
or I_17255 (I295666,I295786,I296170);
DFFARX1 I_17256 (I296170,I2859,I295692,I295684,);
not I_17257 (I296270,I2866);
DFFARX1 I_17258 (I547882,I2859,I296270,I296296,);
not I_17259 (I296304,I296296);
nand I_17260 (I296321,I547867,I547855);
and I_17261 (I296338,I296321,I547870);
DFFARX1 I_17262 (I296338,I2859,I296270,I296364,);
not I_17263 (I296372,I547855);
DFFARX1 I_17264 (I547873,I2859,I296270,I296398,);
not I_17265 (I296406,I296398);
nor I_17266 (I296423,I296406,I296304);
and I_17267 (I296440,I296423,I547855);
nor I_17268 (I296457,I296406,I296372);
nor I_17269 (I296253,I296364,I296457);
DFFARX1 I_17270 (I547861,I2859,I296270,I296497,);
nor I_17271 (I296505,I296497,I296364);
not I_17272 (I296522,I296505);
not I_17273 (I296539,I296497);
nor I_17274 (I296556,I296539,I296440);
DFFARX1 I_17275 (I296556,I2859,I296270,I296256,);
nand I_17276 (I296587,I547858,I547864);
and I_17277 (I296604,I296587,I547879);
DFFARX1 I_17278 (I296604,I2859,I296270,I296630,);
nor I_17279 (I296638,I296630,I296497);
DFFARX1 I_17280 (I296638,I2859,I296270,I296238,);
nand I_17281 (I296669,I296630,I296539);
nand I_17282 (I296247,I296522,I296669);
not I_17283 (I296700,I296630);
nor I_17284 (I296717,I296700,I296440);
DFFARX1 I_17285 (I296717,I2859,I296270,I296259,);
nor I_17286 (I296748,I547876,I547864);
or I_17287 (I296250,I296497,I296748);
nor I_17288 (I296241,I296630,I296748);
or I_17289 (I296244,I296364,I296748);
DFFARX1 I_17290 (I296748,I2859,I296270,I296262,);
not I_17291 (I296848,I2866);
DFFARX1 I_17292 (I45236,I2859,I296848,I296874,);
not I_17293 (I296882,I296874);
nand I_17294 (I296899,I45245,I45254);
and I_17295 (I296916,I296899,I45233);
DFFARX1 I_17296 (I296916,I2859,I296848,I296942,);
not I_17297 (I296950,I45236);
DFFARX1 I_17298 (I45251,I2859,I296848,I296976,);
not I_17299 (I296984,I296976);
nor I_17300 (I297001,I296984,I296882);
and I_17301 (I297018,I297001,I45236);
nor I_17302 (I297035,I296984,I296950);
nor I_17303 (I296831,I296942,I297035);
DFFARX1 I_17304 (I45242,I2859,I296848,I297075,);
nor I_17305 (I297083,I297075,I296942);
not I_17306 (I297100,I297083);
not I_17307 (I297117,I297075);
nor I_17308 (I297134,I297117,I297018);
DFFARX1 I_17309 (I297134,I2859,I296848,I296834,);
nand I_17310 (I297165,I45257,I45233);
and I_17311 (I297182,I297165,I45239);
DFFARX1 I_17312 (I297182,I2859,I296848,I297208,);
nor I_17313 (I297216,I297208,I297075);
DFFARX1 I_17314 (I297216,I2859,I296848,I296816,);
nand I_17315 (I297247,I297208,I297117);
nand I_17316 (I296825,I297100,I297247);
not I_17317 (I297278,I297208);
nor I_17318 (I297295,I297278,I297018);
DFFARX1 I_17319 (I297295,I2859,I296848,I296837,);
nor I_17320 (I297326,I45248,I45233);
or I_17321 (I296828,I297075,I297326);
nor I_17322 (I296819,I297208,I297326);
or I_17323 (I296822,I296942,I297326);
DFFARX1 I_17324 (I297326,I2859,I296848,I296840,);
not I_17325 (I297426,I2866);
DFFARX1 I_17326 (I366395,I2859,I297426,I297452,);
not I_17327 (I297460,I297452);
nand I_17328 (I297477,I366383,I366401);
and I_17329 (I297494,I297477,I366398);
DFFARX1 I_17330 (I297494,I2859,I297426,I297520,);
not I_17331 (I297528,I366389);
DFFARX1 I_17332 (I366386,I2859,I297426,I297554,);
not I_17333 (I297562,I297554);
nor I_17334 (I297579,I297562,I297460);
and I_17335 (I297596,I297579,I366389);
nor I_17336 (I297613,I297562,I297528);
nor I_17337 (I297409,I297520,I297613);
DFFARX1 I_17338 (I366380,I2859,I297426,I297653,);
nor I_17339 (I297661,I297653,I297520);
not I_17340 (I297678,I297661);
not I_17341 (I297695,I297653);
nor I_17342 (I297712,I297695,I297596);
DFFARX1 I_17343 (I297712,I2859,I297426,I297412,);
nand I_17344 (I297743,I366380,I366383);
and I_17345 (I297760,I297743,I366386);
DFFARX1 I_17346 (I297760,I2859,I297426,I297786,);
nor I_17347 (I297794,I297786,I297653);
DFFARX1 I_17348 (I297794,I2859,I297426,I297394,);
nand I_17349 (I297825,I297786,I297695);
nand I_17350 (I297403,I297678,I297825);
not I_17351 (I297856,I297786);
nor I_17352 (I297873,I297856,I297596);
DFFARX1 I_17353 (I297873,I2859,I297426,I297415,);
nor I_17354 (I297904,I366392,I366383);
or I_17355 (I297406,I297653,I297904);
nor I_17356 (I297397,I297786,I297904);
or I_17357 (I297400,I297520,I297904);
DFFARX1 I_17358 (I297904,I2859,I297426,I297418,);
not I_17359 (I298004,I2866);
DFFARX1 I_17360 (I516218,I2859,I298004,I298030,);
not I_17361 (I298038,I298030);
nand I_17362 (I298055,I516221,I516230);
and I_17363 (I298072,I298055,I516233);
DFFARX1 I_17364 (I298072,I2859,I298004,I298098,);
not I_17365 (I298106,I516242);
DFFARX1 I_17366 (I516224,I2859,I298004,I298132,);
not I_17367 (I298140,I298132);
nor I_17368 (I298157,I298140,I298038);
and I_17369 (I298174,I298157,I516242);
nor I_17370 (I298191,I298140,I298106);
nor I_17371 (I297987,I298098,I298191);
DFFARX1 I_17372 (I516221,I2859,I298004,I298231,);
nor I_17373 (I298239,I298231,I298098);
not I_17374 (I298256,I298239);
not I_17375 (I298273,I298231);
nor I_17376 (I298290,I298273,I298174);
DFFARX1 I_17377 (I298290,I2859,I298004,I297990,);
nand I_17378 (I298321,I516239,I516218);
and I_17379 (I298338,I298321,I516236);
DFFARX1 I_17380 (I298338,I2859,I298004,I298364,);
nor I_17381 (I298372,I298364,I298231);
DFFARX1 I_17382 (I298372,I2859,I298004,I297972,);
nand I_17383 (I298403,I298364,I298273);
nand I_17384 (I297981,I298256,I298403);
not I_17385 (I298434,I298364);
nor I_17386 (I298451,I298434,I298174);
DFFARX1 I_17387 (I298451,I2859,I298004,I297993,);
nor I_17388 (I298482,I516227,I516218);
or I_17389 (I297984,I298231,I298482);
nor I_17390 (I297975,I298364,I298482);
or I_17391 (I297978,I298098,I298482);
DFFARX1 I_17392 (I298482,I2859,I298004,I297996,);
not I_17393 (I298582,I2866);
DFFARX1 I_17394 (I157746,I2859,I298582,I298608,);
not I_17395 (I298616,I298608);
nand I_17396 (I298633,I157749,I157725);
and I_17397 (I298650,I298633,I157722);
DFFARX1 I_17398 (I298650,I2859,I298582,I298676,);
not I_17399 (I298684,I157728);
DFFARX1 I_17400 (I157722,I2859,I298582,I298710,);
not I_17401 (I298718,I298710);
nor I_17402 (I298735,I298718,I298616);
and I_17403 (I298752,I298735,I157728);
nor I_17404 (I298769,I298718,I298684);
nor I_17405 (I298565,I298676,I298769);
DFFARX1 I_17406 (I157731,I2859,I298582,I298809,);
nor I_17407 (I298817,I298809,I298676);
not I_17408 (I298834,I298817);
not I_17409 (I298851,I298809);
nor I_17410 (I298868,I298851,I298752);
DFFARX1 I_17411 (I298868,I2859,I298582,I298568,);
nand I_17412 (I298899,I157734,I157743);
and I_17413 (I298916,I298899,I157740);
DFFARX1 I_17414 (I298916,I2859,I298582,I298942,);
nor I_17415 (I298950,I298942,I298809);
DFFARX1 I_17416 (I298950,I2859,I298582,I298550,);
nand I_17417 (I298981,I298942,I298851);
nand I_17418 (I298559,I298834,I298981);
not I_17419 (I299012,I298942);
nor I_17420 (I299029,I299012,I298752);
DFFARX1 I_17421 (I299029,I2859,I298582,I298571,);
nor I_17422 (I299060,I157737,I157743);
or I_17423 (I298562,I298809,I299060);
nor I_17424 (I298553,I298942,I299060);
or I_17425 (I298556,I298676,I299060);
DFFARX1 I_17426 (I299060,I2859,I298582,I298574,);
not I_17427 (I299160,I2866);
DFFARX1 I_17428 (I553832,I2859,I299160,I299186,);
not I_17429 (I299194,I299186);
nand I_17430 (I299211,I553817,I553805);
and I_17431 (I299228,I299211,I553820);
DFFARX1 I_17432 (I299228,I2859,I299160,I299254,);
not I_17433 (I299262,I553805);
DFFARX1 I_17434 (I553823,I2859,I299160,I299288,);
not I_17435 (I299296,I299288);
nor I_17436 (I299313,I299296,I299194);
and I_17437 (I299330,I299313,I553805);
nor I_17438 (I299347,I299296,I299262);
nor I_17439 (I299143,I299254,I299347);
DFFARX1 I_17440 (I553811,I2859,I299160,I299387,);
nor I_17441 (I299395,I299387,I299254);
not I_17442 (I299412,I299395);
not I_17443 (I299429,I299387);
nor I_17444 (I299446,I299429,I299330);
DFFARX1 I_17445 (I299446,I2859,I299160,I299146,);
nand I_17446 (I299477,I553808,I553814);
and I_17447 (I299494,I299477,I553829);
DFFARX1 I_17448 (I299494,I2859,I299160,I299520,);
nor I_17449 (I299528,I299520,I299387);
DFFARX1 I_17450 (I299528,I2859,I299160,I299128,);
nand I_17451 (I299559,I299520,I299429);
nand I_17452 (I299137,I299412,I299559);
not I_17453 (I299590,I299520);
nor I_17454 (I299607,I299590,I299330);
DFFARX1 I_17455 (I299607,I2859,I299160,I299149,);
nor I_17456 (I299638,I553826,I553814);
or I_17457 (I299140,I299387,I299638);
nor I_17458 (I299131,I299520,I299638);
or I_17459 (I299134,I299254,I299638);
DFFARX1 I_17460 (I299638,I2859,I299160,I299152,);
not I_17461 (I299738,I2866);
DFFARX1 I_17462 (I232080,I2859,I299738,I299764,);
not I_17463 (I299772,I299764);
nand I_17464 (I299789,I232089,I232098);
and I_17465 (I299806,I299789,I232104);
DFFARX1 I_17466 (I299806,I2859,I299738,I299832,);
not I_17467 (I299840,I232101);
DFFARX1 I_17468 (I232086,I2859,I299738,I299866,);
not I_17469 (I299874,I299866);
nor I_17470 (I299891,I299874,I299772);
and I_17471 (I299908,I299891,I232101);
nor I_17472 (I299925,I299874,I299840);
nor I_17473 (I299721,I299832,I299925);
DFFARX1 I_17474 (I232095,I2859,I299738,I299965,);
nor I_17475 (I299973,I299965,I299832);
not I_17476 (I299990,I299973);
not I_17477 (I300007,I299965);
nor I_17478 (I300024,I300007,I299908);
DFFARX1 I_17479 (I300024,I2859,I299738,I299724,);
nand I_17480 (I300055,I232092,I232083);
and I_17481 (I300072,I300055,I232080);
DFFARX1 I_17482 (I300072,I2859,I299738,I300098,);
nor I_17483 (I300106,I300098,I299965);
DFFARX1 I_17484 (I300106,I2859,I299738,I299706,);
nand I_17485 (I300137,I300098,I300007);
nand I_17486 (I299715,I299990,I300137);
not I_17487 (I300168,I300098);
nor I_17488 (I300185,I300168,I299908);
DFFARX1 I_17489 (I300185,I2859,I299738,I299727,);
nor I_17490 (I300216,I232083,I232083);
or I_17491 (I299718,I299965,I300216);
nor I_17492 (I299709,I300098,I300216);
or I_17493 (I299712,I299832,I300216);
DFFARX1 I_17494 (I300216,I2859,I299738,I299730,);
not I_17495 (I300316,I2866);
DFFARX1 I_17496 (I524004,I2859,I300316,I300342,);
not I_17497 (I300350,I300342);
nand I_17498 (I300367,I524028,I524010);
and I_17499 (I300384,I300367,I524016);
DFFARX1 I_17500 (I300384,I2859,I300316,I300410,);
not I_17501 (I300418,I524022);
DFFARX1 I_17502 (I524007,I2859,I300316,I300444,);
not I_17503 (I300452,I300444);
nor I_17504 (I300469,I300452,I300350);
and I_17505 (I300486,I300469,I524022);
nor I_17506 (I300503,I300452,I300418);
nor I_17507 (I300299,I300410,I300503);
DFFARX1 I_17508 (I524019,I2859,I300316,I300543,);
nor I_17509 (I300551,I300543,I300410);
not I_17510 (I300568,I300551);
not I_17511 (I300585,I300543);
nor I_17512 (I300602,I300585,I300486);
DFFARX1 I_17513 (I300602,I2859,I300316,I300302,);
nand I_17514 (I300633,I524025,I524013);
and I_17515 (I300650,I300633,I524007);
DFFARX1 I_17516 (I300650,I2859,I300316,I300676,);
nor I_17517 (I300684,I300676,I300543);
DFFARX1 I_17518 (I300684,I2859,I300316,I300284,);
nand I_17519 (I300715,I300676,I300585);
nand I_17520 (I300293,I300568,I300715);
not I_17521 (I300746,I300676);
nor I_17522 (I300763,I300746,I300486);
DFFARX1 I_17523 (I300763,I2859,I300316,I300305,);
nor I_17524 (I300794,I524004,I524013);
or I_17525 (I300296,I300543,I300794);
nor I_17526 (I300287,I300676,I300794);
or I_17527 (I300290,I300410,I300794);
DFFARX1 I_17528 (I300794,I2859,I300316,I300308,);
not I_17529 (I300894,I2866);
DFFARX1 I_17530 (I482440,I2859,I300894,I300920,);
not I_17531 (I300928,I300920);
nand I_17532 (I300945,I482422,I482434);
and I_17533 (I300962,I300945,I482437);
DFFARX1 I_17534 (I300962,I2859,I300894,I300988,);
not I_17535 (I300996,I482431);
DFFARX1 I_17536 (I482428,I2859,I300894,I301022,);
not I_17537 (I301030,I301022);
nor I_17538 (I301047,I301030,I300928);
and I_17539 (I301064,I301047,I482431);
nor I_17540 (I301081,I301030,I300996);
nor I_17541 (I300877,I300988,I301081);
DFFARX1 I_17542 (I482446,I2859,I300894,I301121,);
nor I_17543 (I301129,I301121,I300988);
not I_17544 (I301146,I301129);
not I_17545 (I301163,I301121);
nor I_17546 (I301180,I301163,I301064);
DFFARX1 I_17547 (I301180,I2859,I300894,I300880,);
nand I_17548 (I301211,I482425,I482425);
and I_17549 (I301228,I301211,I482422);
DFFARX1 I_17550 (I301228,I2859,I300894,I301254,);
nor I_17551 (I301262,I301254,I301121);
DFFARX1 I_17552 (I301262,I2859,I300894,I300862,);
nand I_17553 (I301293,I301254,I301163);
nand I_17554 (I300871,I301146,I301293);
not I_17555 (I301324,I301254);
nor I_17556 (I301341,I301324,I301064);
DFFARX1 I_17557 (I301341,I2859,I300894,I300883,);
nor I_17558 (I301372,I482443,I482425);
or I_17559 (I300874,I301121,I301372);
nor I_17560 (I300865,I301254,I301372);
or I_17561 (I300868,I300988,I301372);
DFFARX1 I_17562 (I301372,I2859,I300894,I300886,);
not I_17563 (I301472,I2866);
DFFARX1 I_17564 (I447204,I2859,I301472,I301498,);
not I_17565 (I301506,I301498);
nand I_17566 (I301523,I447201,I447219);
and I_17567 (I301540,I301523,I447216);
DFFARX1 I_17568 (I301540,I2859,I301472,I301566,);
not I_17569 (I301574,I447198);
DFFARX1 I_17570 (I447201,I2859,I301472,I301600,);
not I_17571 (I301608,I301600);
nor I_17572 (I301625,I301608,I301506);
and I_17573 (I301642,I301625,I447198);
nor I_17574 (I301659,I301608,I301574);
nor I_17575 (I301455,I301566,I301659);
DFFARX1 I_17576 (I447210,I2859,I301472,I301699,);
nor I_17577 (I301707,I301699,I301566);
not I_17578 (I301724,I301707);
not I_17579 (I301741,I301699);
nor I_17580 (I301758,I301741,I301642);
DFFARX1 I_17581 (I301758,I2859,I301472,I301458,);
nand I_17582 (I301789,I447213,I447198);
and I_17583 (I301806,I301789,I447204);
DFFARX1 I_17584 (I301806,I2859,I301472,I301832,);
nor I_17585 (I301840,I301832,I301699);
DFFARX1 I_17586 (I301840,I2859,I301472,I301440,);
nand I_17587 (I301871,I301832,I301741);
nand I_17588 (I301449,I301724,I301871);
not I_17589 (I301902,I301832);
nor I_17590 (I301919,I301902,I301642);
DFFARX1 I_17591 (I301919,I2859,I301472,I301461,);
nor I_17592 (I301950,I447207,I447198);
or I_17593 (I301452,I301699,I301950);
nor I_17594 (I301443,I301832,I301950);
or I_17595 (I301446,I301566,I301950);
DFFARX1 I_17596 (I301950,I2859,I301472,I301464,);
not I_17597 (I302050,I2866);
DFFARX1 I_17598 (I530940,I2859,I302050,I302076,);
not I_17599 (I302084,I302076);
nand I_17600 (I302101,I530964,I530946);
and I_17601 (I302118,I302101,I530952);
DFFARX1 I_17602 (I302118,I2859,I302050,I302144,);
not I_17603 (I302152,I530958);
DFFARX1 I_17604 (I530943,I2859,I302050,I302178,);
not I_17605 (I302186,I302178);
nor I_17606 (I302203,I302186,I302084);
and I_17607 (I302220,I302203,I530958);
nor I_17608 (I302237,I302186,I302152);
nor I_17609 (I302033,I302144,I302237);
DFFARX1 I_17610 (I530955,I2859,I302050,I302277,);
nor I_17611 (I302285,I302277,I302144);
not I_17612 (I302302,I302285);
not I_17613 (I302319,I302277);
nor I_17614 (I302336,I302319,I302220);
DFFARX1 I_17615 (I302336,I2859,I302050,I302036,);
nand I_17616 (I302367,I530961,I530949);
and I_17617 (I302384,I302367,I530943);
DFFARX1 I_17618 (I302384,I2859,I302050,I302410,);
nor I_17619 (I302418,I302410,I302277);
DFFARX1 I_17620 (I302418,I2859,I302050,I302018,);
nand I_17621 (I302449,I302410,I302319);
nand I_17622 (I302027,I302302,I302449);
not I_17623 (I302480,I302410);
nor I_17624 (I302497,I302480,I302220);
DFFARX1 I_17625 (I302497,I2859,I302050,I302039,);
nor I_17626 (I302528,I530940,I530949);
or I_17627 (I302030,I302277,I302528);
nor I_17628 (I302021,I302410,I302528);
or I_17629 (I302024,I302144,I302528);
DFFARX1 I_17630 (I302528,I2859,I302050,I302042,);
not I_17631 (I302628,I2866);
DFFARX1 I_17632 (I365868,I2859,I302628,I302654,);
not I_17633 (I302662,I302654);
nand I_17634 (I302679,I365856,I365874);
and I_17635 (I302696,I302679,I365871);
DFFARX1 I_17636 (I302696,I2859,I302628,I302722,);
not I_17637 (I302730,I365862);
DFFARX1 I_17638 (I365859,I2859,I302628,I302756,);
not I_17639 (I302764,I302756);
nor I_17640 (I302781,I302764,I302662);
and I_17641 (I302798,I302781,I365862);
nor I_17642 (I302815,I302764,I302730);
nor I_17643 (I302611,I302722,I302815);
DFFARX1 I_17644 (I365853,I2859,I302628,I302855,);
nor I_17645 (I302863,I302855,I302722);
not I_17646 (I302880,I302863);
not I_17647 (I302897,I302855);
nor I_17648 (I302914,I302897,I302798);
DFFARX1 I_17649 (I302914,I2859,I302628,I302614,);
nand I_17650 (I302945,I365853,I365856);
and I_17651 (I302962,I302945,I365859);
DFFARX1 I_17652 (I302962,I2859,I302628,I302988,);
nor I_17653 (I302996,I302988,I302855);
DFFARX1 I_17654 (I302996,I2859,I302628,I302596,);
nand I_17655 (I303027,I302988,I302897);
nand I_17656 (I302605,I302880,I303027);
not I_17657 (I303058,I302988);
nor I_17658 (I303075,I303058,I302798);
DFFARX1 I_17659 (I303075,I2859,I302628,I302617,);
nor I_17660 (I303106,I365865,I365856);
or I_17661 (I302608,I302855,I303106);
nor I_17662 (I302599,I302988,I303106);
or I_17663 (I302602,I302722,I303106);
DFFARX1 I_17664 (I303106,I2859,I302628,I302620,);
not I_17665 (I303206,I2866);
DFFARX1 I_17666 (I485330,I2859,I303206,I303232,);
not I_17667 (I303240,I303232);
nand I_17668 (I303257,I485312,I485324);
and I_17669 (I303274,I303257,I485327);
DFFARX1 I_17670 (I303274,I2859,I303206,I303300,);
not I_17671 (I303308,I485321);
DFFARX1 I_17672 (I485318,I2859,I303206,I303334,);
not I_17673 (I303342,I303334);
nor I_17674 (I303359,I303342,I303240);
and I_17675 (I303376,I303359,I485321);
nor I_17676 (I303393,I303342,I303308);
nor I_17677 (I303189,I303300,I303393);
DFFARX1 I_17678 (I485336,I2859,I303206,I303433,);
nor I_17679 (I303441,I303433,I303300);
not I_17680 (I303458,I303441);
not I_17681 (I303475,I303433);
nor I_17682 (I303492,I303475,I303376);
DFFARX1 I_17683 (I303492,I2859,I303206,I303192,);
nand I_17684 (I303523,I485315,I485315);
and I_17685 (I303540,I303523,I485312);
DFFARX1 I_17686 (I303540,I2859,I303206,I303566,);
nor I_17687 (I303574,I303566,I303433);
DFFARX1 I_17688 (I303574,I2859,I303206,I303174,);
nand I_17689 (I303605,I303566,I303475);
nand I_17690 (I303183,I303458,I303605);
not I_17691 (I303636,I303566);
nor I_17692 (I303653,I303636,I303376);
DFFARX1 I_17693 (I303653,I2859,I303206,I303195,);
nor I_17694 (I303684,I485333,I485315);
or I_17695 (I303186,I303433,I303684);
nor I_17696 (I303177,I303566,I303684);
or I_17697 (I303180,I303300,I303684);
DFFARX1 I_17698 (I303684,I2859,I303206,I303198,);
not I_17699 (I303784,I2866);
DFFARX1 I_17700 (I357436,I2859,I303784,I303810,);
not I_17701 (I303818,I303810);
nand I_17702 (I303835,I357424,I357442);
and I_17703 (I303852,I303835,I357439);
DFFARX1 I_17704 (I303852,I2859,I303784,I303878,);
not I_17705 (I303886,I357430);
DFFARX1 I_17706 (I357427,I2859,I303784,I303912,);
not I_17707 (I303920,I303912);
nor I_17708 (I303937,I303920,I303818);
and I_17709 (I303954,I303937,I357430);
nor I_17710 (I303971,I303920,I303886);
nor I_17711 (I303767,I303878,I303971);
DFFARX1 I_17712 (I357421,I2859,I303784,I304011,);
nor I_17713 (I304019,I304011,I303878);
not I_17714 (I304036,I304019);
not I_17715 (I304053,I304011);
nor I_17716 (I304070,I304053,I303954);
DFFARX1 I_17717 (I304070,I2859,I303784,I303770,);
nand I_17718 (I304101,I357421,I357424);
and I_17719 (I304118,I304101,I357427);
DFFARX1 I_17720 (I304118,I2859,I303784,I304144,);
nor I_17721 (I304152,I304144,I304011);
DFFARX1 I_17722 (I304152,I2859,I303784,I303752,);
nand I_17723 (I304183,I304144,I304053);
nand I_17724 (I303761,I304036,I304183);
not I_17725 (I304214,I304144);
nor I_17726 (I304231,I304214,I303954);
DFFARX1 I_17727 (I304231,I2859,I303784,I303773,);
nor I_17728 (I304262,I357433,I357424);
or I_17729 (I303764,I304011,I304262);
nor I_17730 (I303755,I304144,I304262);
or I_17731 (I303758,I303878,I304262);
DFFARX1 I_17732 (I304262,I2859,I303784,I303776,);
not I_17733 (I304362,I2866);
DFFARX1 I_17734 (I333721,I2859,I304362,I304388,);
not I_17735 (I304396,I304388);
nand I_17736 (I304413,I333709,I333727);
and I_17737 (I304430,I304413,I333724);
DFFARX1 I_17738 (I304430,I2859,I304362,I304456,);
not I_17739 (I304464,I333715);
DFFARX1 I_17740 (I333712,I2859,I304362,I304490,);
not I_17741 (I304498,I304490);
nor I_17742 (I304515,I304498,I304396);
and I_17743 (I304532,I304515,I333715);
nor I_17744 (I304549,I304498,I304464);
nor I_17745 (I304345,I304456,I304549);
DFFARX1 I_17746 (I333706,I2859,I304362,I304589,);
nor I_17747 (I304597,I304589,I304456);
not I_17748 (I304614,I304597);
not I_17749 (I304631,I304589);
nor I_17750 (I304648,I304631,I304532);
DFFARX1 I_17751 (I304648,I2859,I304362,I304348,);
nand I_17752 (I304679,I333706,I333709);
and I_17753 (I304696,I304679,I333712);
DFFARX1 I_17754 (I304696,I2859,I304362,I304722,);
nor I_17755 (I304730,I304722,I304589);
DFFARX1 I_17756 (I304730,I2859,I304362,I304330,);
nand I_17757 (I304761,I304722,I304631);
nand I_17758 (I304339,I304614,I304761);
not I_17759 (I304792,I304722);
nor I_17760 (I304809,I304792,I304532);
DFFARX1 I_17761 (I304809,I2859,I304362,I304351,);
nor I_17762 (I304840,I333718,I333709);
or I_17763 (I304342,I304589,I304840);
nor I_17764 (I304333,I304722,I304840);
or I_17765 (I304336,I304456,I304840);
DFFARX1 I_17766 (I304840,I2859,I304362,I304354,);
not I_17767 (I304940,I2866);
DFFARX1 I_17768 (I192292,I2859,I304940,I304966,);
not I_17769 (I304974,I304966);
nand I_17770 (I304991,I192283,I192301);
and I_17771 (I305008,I304991,I192304);
DFFARX1 I_17772 (I305008,I2859,I304940,I305034,);
not I_17773 (I305042,I192298);
DFFARX1 I_17774 (I192286,I2859,I304940,I305068,);
not I_17775 (I305076,I305068);
nor I_17776 (I305093,I305076,I304974);
and I_17777 (I305110,I305093,I192298);
nor I_17778 (I305127,I305076,I305042);
nor I_17779 (I304923,I305034,I305127);
DFFARX1 I_17780 (I192295,I2859,I304940,I305167,);
nor I_17781 (I305175,I305167,I305034);
not I_17782 (I305192,I305175);
not I_17783 (I305209,I305167);
nor I_17784 (I305226,I305209,I305110);
DFFARX1 I_17785 (I305226,I2859,I304940,I304926,);
nand I_17786 (I305257,I192310,I192307);
and I_17787 (I305274,I305257,I192289);
DFFARX1 I_17788 (I305274,I2859,I304940,I305300,);
nor I_17789 (I305308,I305300,I305167);
DFFARX1 I_17790 (I305308,I2859,I304940,I304908,);
nand I_17791 (I305339,I305300,I305209);
nand I_17792 (I304917,I305192,I305339);
not I_17793 (I305370,I305300);
nor I_17794 (I305387,I305370,I305110);
DFFARX1 I_17795 (I305387,I2859,I304940,I304929,);
nor I_17796 (I305418,I192283,I192307);
or I_17797 (I304920,I305167,I305418);
nor I_17798 (I304911,I305300,I305418);
or I_17799 (I304914,I305034,I305418);
DFFARX1 I_17800 (I305418,I2859,I304940,I304932,);
not I_17801 (I305518,I2866);
DFFARX1 I_17802 (I380293,I2859,I305518,I305544,);
not I_17803 (I305552,I305544);
nand I_17804 (I305569,I380269,I380284);
and I_17805 (I305586,I305569,I380296);
DFFARX1 I_17806 (I305586,I2859,I305518,I305612,);
not I_17807 (I305620,I380281);
DFFARX1 I_17808 (I380272,I2859,I305518,I305646,);
not I_17809 (I305654,I305646);
nor I_17810 (I305671,I305654,I305552);
and I_17811 (I305688,I305671,I380281);
nor I_17812 (I305705,I305654,I305620);
nor I_17813 (I305501,I305612,I305705);
DFFARX1 I_17814 (I380269,I2859,I305518,I305745,);
nor I_17815 (I305753,I305745,I305612);
not I_17816 (I305770,I305753);
not I_17817 (I305787,I305745);
nor I_17818 (I305804,I305787,I305688);
DFFARX1 I_17819 (I305804,I2859,I305518,I305504,);
nand I_17820 (I305835,I380287,I380278);
and I_17821 (I305852,I305835,I380290);
DFFARX1 I_17822 (I305852,I2859,I305518,I305878,);
nor I_17823 (I305886,I305878,I305745);
DFFARX1 I_17824 (I305886,I2859,I305518,I305486,);
nand I_17825 (I305917,I305878,I305787);
nand I_17826 (I305495,I305770,I305917);
not I_17827 (I305948,I305878);
nor I_17828 (I305965,I305948,I305688);
DFFARX1 I_17829 (I305965,I2859,I305518,I305507,);
nor I_17830 (I305996,I380275,I380278);
or I_17831 (I305498,I305745,I305996);
nor I_17832 (I305489,I305878,I305996);
or I_17833 (I305492,I305612,I305996);
DFFARX1 I_17834 (I305996,I2859,I305518,I305510,);
not I_17835 (I306096,I2866);
DFFARX1 I_17836 (I33115,I2859,I306096,I306122,);
not I_17837 (I306130,I306122);
nand I_17838 (I306147,I33124,I33133);
and I_17839 (I306164,I306147,I33112);
DFFARX1 I_17840 (I306164,I2859,I306096,I306190,);
not I_17841 (I306198,I33115);
DFFARX1 I_17842 (I33130,I2859,I306096,I306224,);
not I_17843 (I306232,I306224);
nor I_17844 (I306249,I306232,I306130);
and I_17845 (I306266,I306249,I33115);
nor I_17846 (I306283,I306232,I306198);
nor I_17847 (I306079,I306190,I306283);
DFFARX1 I_17848 (I33121,I2859,I306096,I306323,);
nor I_17849 (I306331,I306323,I306190);
not I_17850 (I306348,I306331);
not I_17851 (I306365,I306323);
nor I_17852 (I306382,I306365,I306266);
DFFARX1 I_17853 (I306382,I2859,I306096,I306082,);
nand I_17854 (I306413,I33136,I33112);
and I_17855 (I306430,I306413,I33118);
DFFARX1 I_17856 (I306430,I2859,I306096,I306456,);
nor I_17857 (I306464,I306456,I306323);
DFFARX1 I_17858 (I306464,I2859,I306096,I306064,);
nand I_17859 (I306495,I306456,I306365);
nand I_17860 (I306073,I306348,I306495);
not I_17861 (I306526,I306456);
nor I_17862 (I306543,I306526,I306266);
DFFARX1 I_17863 (I306543,I2859,I306096,I306085,);
nor I_17864 (I306574,I33127,I33112);
or I_17865 (I306076,I306323,I306574);
nor I_17866 (I306067,I306456,I306574);
or I_17867 (I306070,I306190,I306574);
DFFARX1 I_17868 (I306574,I2859,I306096,I306088,);
not I_17869 (I306674,I2866);
DFFARX1 I_17870 (I110316,I2859,I306674,I306700,);
not I_17871 (I306708,I306700);
nand I_17872 (I306725,I110319,I110295);
and I_17873 (I306742,I306725,I110292);
DFFARX1 I_17874 (I306742,I2859,I306674,I306768,);
not I_17875 (I306776,I110298);
DFFARX1 I_17876 (I110292,I2859,I306674,I306802,);
not I_17877 (I306810,I306802);
nor I_17878 (I306827,I306810,I306708);
and I_17879 (I306844,I306827,I110298);
nor I_17880 (I306861,I306810,I306776);
nor I_17881 (I306657,I306768,I306861);
DFFARX1 I_17882 (I110301,I2859,I306674,I306901,);
nor I_17883 (I306909,I306901,I306768);
not I_17884 (I306926,I306909);
not I_17885 (I306943,I306901);
nor I_17886 (I306960,I306943,I306844);
DFFARX1 I_17887 (I306960,I2859,I306674,I306660,);
nand I_17888 (I306991,I110304,I110313);
and I_17889 (I307008,I306991,I110310);
DFFARX1 I_17890 (I307008,I2859,I306674,I307034,);
nor I_17891 (I307042,I307034,I306901);
DFFARX1 I_17892 (I307042,I2859,I306674,I306642,);
nand I_17893 (I307073,I307034,I306943);
nand I_17894 (I306651,I306926,I307073);
not I_17895 (I307104,I307034);
nor I_17896 (I307121,I307104,I306844);
DFFARX1 I_17897 (I307121,I2859,I306674,I306663,);
nor I_17898 (I307152,I110307,I110313);
or I_17899 (I306654,I306901,I307152);
nor I_17900 (I306645,I307034,I307152);
or I_17901 (I306648,I306768,I307152);
DFFARX1 I_17902 (I307152,I2859,I306674,I306666,);
not I_17903 (I307252,I2866);
DFFARX1 I_17904 (I465100,I2859,I307252,I307278,);
not I_17905 (I307286,I307278);
nand I_17906 (I307303,I465082,I465094);
and I_17907 (I307320,I307303,I465097);
DFFARX1 I_17908 (I307320,I2859,I307252,I307346,);
not I_17909 (I307354,I465091);
DFFARX1 I_17910 (I465088,I2859,I307252,I307380,);
not I_17911 (I307388,I307380);
nor I_17912 (I307405,I307388,I307286);
and I_17913 (I307422,I307405,I465091);
nor I_17914 (I307439,I307388,I307354);
nor I_17915 (I307235,I307346,I307439);
DFFARX1 I_17916 (I465106,I2859,I307252,I307479,);
nor I_17917 (I307487,I307479,I307346);
not I_17918 (I307504,I307487);
not I_17919 (I307521,I307479);
nor I_17920 (I307538,I307521,I307422);
DFFARX1 I_17921 (I307538,I2859,I307252,I307238,);
nand I_17922 (I307569,I465085,I465085);
and I_17923 (I307586,I307569,I465082);
DFFARX1 I_17924 (I307586,I2859,I307252,I307612,);
nor I_17925 (I307620,I307612,I307479);
DFFARX1 I_17926 (I307620,I2859,I307252,I307220,);
nand I_17927 (I307651,I307612,I307521);
nand I_17928 (I307229,I307504,I307651);
not I_17929 (I307682,I307612);
nor I_17930 (I307699,I307682,I307422);
DFFARX1 I_17931 (I307699,I2859,I307252,I307241,);
nor I_17932 (I307730,I465103,I465085);
or I_17933 (I307232,I307479,I307730);
nor I_17934 (I307223,I307612,I307730);
or I_17935 (I307226,I307346,I307730);
DFFARX1 I_17936 (I307730,I2859,I307252,I307244,);
not I_17937 (I307830,I2866);
DFFARX1 I_17938 (I220843,I2859,I307830,I307856,);
not I_17939 (I307864,I307856);
nand I_17940 (I307881,I220858,I220843);
and I_17941 (I307898,I307881,I220846);
DFFARX1 I_17942 (I307898,I2859,I307830,I307924,);
not I_17943 (I307932,I220846);
DFFARX1 I_17944 (I220855,I2859,I307830,I307958,);
not I_17945 (I307966,I307958);
nor I_17946 (I307983,I307966,I307864);
and I_17947 (I308000,I307983,I220846);
nor I_17948 (I308017,I307966,I307932);
nor I_17949 (I307813,I307924,I308017);
DFFARX1 I_17950 (I220849,I2859,I307830,I308057,);
nor I_17951 (I308065,I308057,I307924);
not I_17952 (I308082,I308065);
not I_17953 (I308099,I308057);
nor I_17954 (I308116,I308099,I308000);
DFFARX1 I_17955 (I308116,I2859,I307830,I307816,);
nand I_17956 (I308147,I220852,I220861);
and I_17957 (I308164,I308147,I220867);
DFFARX1 I_17958 (I308164,I2859,I307830,I308190,);
nor I_17959 (I308198,I308190,I308057);
DFFARX1 I_17960 (I308198,I2859,I307830,I307798,);
nand I_17961 (I308229,I308190,I308099);
nand I_17962 (I307807,I308082,I308229);
not I_17963 (I308260,I308190);
nor I_17964 (I308277,I308260,I308000);
DFFARX1 I_17965 (I308277,I2859,I307830,I307819,);
nor I_17966 (I308308,I220864,I220861);
or I_17967 (I307810,I308057,I308308);
nor I_17968 (I307801,I308190,I308308);
or I_17969 (I307804,I307924,I308308);
DFFARX1 I_17970 (I308308,I2859,I307830,I307822,);
not I_17971 (I308408,I2866);
DFFARX1 I_17972 (I351639,I2859,I308408,I308434,);
not I_17973 (I308442,I308434);
nand I_17974 (I308459,I351627,I351645);
and I_17975 (I308476,I308459,I351642);
DFFARX1 I_17976 (I308476,I2859,I308408,I308502,);
not I_17977 (I308510,I351633);
DFFARX1 I_17978 (I351630,I2859,I308408,I308536,);
not I_17979 (I308544,I308536);
nor I_17980 (I308561,I308544,I308442);
and I_17981 (I308578,I308561,I351633);
nor I_17982 (I308595,I308544,I308510);
nor I_17983 (I308391,I308502,I308595);
DFFARX1 I_17984 (I351624,I2859,I308408,I308635,);
nor I_17985 (I308643,I308635,I308502);
not I_17986 (I308660,I308643);
not I_17987 (I308677,I308635);
nor I_17988 (I308694,I308677,I308578);
DFFARX1 I_17989 (I308694,I2859,I308408,I308394,);
nand I_17990 (I308725,I351624,I351627);
and I_17991 (I308742,I308725,I351630);
DFFARX1 I_17992 (I308742,I2859,I308408,I308768,);
nor I_17993 (I308776,I308768,I308635);
DFFARX1 I_17994 (I308776,I2859,I308408,I308376,);
nand I_17995 (I308807,I308768,I308677);
nand I_17996 (I308385,I308660,I308807);
not I_17997 (I308838,I308768);
nor I_17998 (I308855,I308838,I308578);
DFFARX1 I_17999 (I308855,I2859,I308408,I308397,);
nor I_18000 (I308886,I351636,I351627);
or I_18001 (I308388,I308635,I308886);
nor I_18002 (I308379,I308768,I308886);
or I_18003 (I308382,I308502,I308886);
DFFARX1 I_18004 (I308886,I2859,I308408,I308400,);
not I_18005 (I308986,I2866);
DFFARX1 I_18006 (I534408,I2859,I308986,I309012,);
not I_18007 (I309020,I309012);
nand I_18008 (I309037,I534432,I534414);
and I_18009 (I309054,I309037,I534420);
DFFARX1 I_18010 (I309054,I2859,I308986,I309080,);
not I_18011 (I309088,I534426);
DFFARX1 I_18012 (I534411,I2859,I308986,I309114,);
not I_18013 (I309122,I309114);
nor I_18014 (I309139,I309122,I309020);
and I_18015 (I309156,I309139,I534426);
nor I_18016 (I309173,I309122,I309088);
nor I_18017 (I308969,I309080,I309173);
DFFARX1 I_18018 (I534423,I2859,I308986,I309213,);
nor I_18019 (I309221,I309213,I309080);
not I_18020 (I309238,I309221);
not I_18021 (I309255,I309213);
nor I_18022 (I309272,I309255,I309156);
DFFARX1 I_18023 (I309272,I2859,I308986,I308972,);
nand I_18024 (I309303,I534429,I534417);
and I_18025 (I309320,I309303,I534411);
DFFARX1 I_18026 (I309320,I2859,I308986,I309346,);
nor I_18027 (I309354,I309346,I309213);
DFFARX1 I_18028 (I309354,I2859,I308986,I308954,);
nand I_18029 (I309385,I309346,I309255);
nand I_18030 (I308963,I309238,I309385);
not I_18031 (I309416,I309346);
nor I_18032 (I309433,I309416,I309156);
DFFARX1 I_18033 (I309433,I2859,I308986,I308975,);
nor I_18034 (I309464,I534408,I534417);
or I_18035 (I308966,I309213,I309464);
nor I_18036 (I308957,I309346,I309464);
or I_18037 (I308960,I309080,I309464);
DFFARX1 I_18038 (I309464,I2859,I308986,I308978,);
not I_18039 (I309564,I2866);
DFFARX1 I_18040 (I79233,I2859,I309564,I309590,);
not I_18041 (I309598,I309590);
nand I_18042 (I309615,I79236,I79257);
and I_18043 (I309632,I309615,I79245);
DFFARX1 I_18044 (I309632,I2859,I309564,I309658,);
not I_18045 (I309666,I79242);
DFFARX1 I_18046 (I79233,I2859,I309564,I309692,);
not I_18047 (I309700,I309692);
nor I_18048 (I309717,I309700,I309598);
and I_18049 (I309734,I309717,I79242);
nor I_18050 (I309751,I309700,I309666);
nor I_18051 (I309547,I309658,I309751);
DFFARX1 I_18052 (I79251,I2859,I309564,I309791,);
nor I_18053 (I309799,I309791,I309658);
not I_18054 (I309816,I309799);
not I_18055 (I309833,I309791);
nor I_18056 (I309850,I309833,I309734);
DFFARX1 I_18057 (I309850,I2859,I309564,I309550,);
nand I_18058 (I309881,I79236,I79239);
and I_18059 (I309898,I309881,I79248);
DFFARX1 I_18060 (I309898,I2859,I309564,I309924,);
nor I_18061 (I309932,I309924,I309791);
DFFARX1 I_18062 (I309932,I2859,I309564,I309532,);
nand I_18063 (I309963,I309924,I309833);
nand I_18064 (I309541,I309816,I309963);
not I_18065 (I309994,I309924);
nor I_18066 (I310011,I309994,I309734);
DFFARX1 I_18067 (I310011,I2859,I309564,I309553,);
nor I_18068 (I310042,I79254,I79239);
or I_18069 (I309544,I309791,I310042);
nor I_18070 (I309535,I309924,I310042);
or I_18071 (I309538,I309658,I310042);
DFFARX1 I_18072 (I310042,I2859,I309564,I309556,);
not I_18073 (I310142,I2866);
DFFARX1 I_18074 (I188484,I2859,I310142,I310168,);
not I_18075 (I310176,I310168);
nand I_18076 (I310193,I188475,I188493);
and I_18077 (I310210,I310193,I188496);
DFFARX1 I_18078 (I310210,I2859,I310142,I310236,);
not I_18079 (I310244,I188490);
DFFARX1 I_18080 (I188478,I2859,I310142,I310270,);
not I_18081 (I310278,I310270);
nor I_18082 (I310295,I310278,I310176);
and I_18083 (I310312,I310295,I188490);
nor I_18084 (I310329,I310278,I310244);
nor I_18085 (I310125,I310236,I310329);
DFFARX1 I_18086 (I188487,I2859,I310142,I310369,);
nor I_18087 (I310377,I310369,I310236);
not I_18088 (I310394,I310377);
not I_18089 (I310411,I310369);
nor I_18090 (I310428,I310411,I310312);
DFFARX1 I_18091 (I310428,I2859,I310142,I310128,);
nand I_18092 (I310459,I188502,I188499);
and I_18093 (I310476,I310459,I188481);
DFFARX1 I_18094 (I310476,I2859,I310142,I310502,);
nor I_18095 (I310510,I310502,I310369);
DFFARX1 I_18096 (I310510,I2859,I310142,I310110,);
nand I_18097 (I310541,I310502,I310411);
nand I_18098 (I310119,I310394,I310541);
not I_18099 (I310572,I310502);
nor I_18100 (I310589,I310572,I310312);
DFFARX1 I_18101 (I310589,I2859,I310142,I310131,);
nor I_18102 (I310620,I188475,I188499);
or I_18103 (I310122,I310369,I310620);
nor I_18104 (I310113,I310502,I310620);
or I_18105 (I310116,I310236,I310620);
DFFARX1 I_18106 (I310620,I2859,I310142,I310134,);
not I_18107 (I310720,I2866);
DFFARX1 I_18108 (I12571,I2859,I310720,I310746,);
not I_18109 (I310754,I310746);
nand I_18110 (I310771,I12568,I12559);
and I_18111 (I310788,I310771,I12559);
DFFARX1 I_18112 (I310788,I2859,I310720,I310814,);
not I_18113 (I310822,I12562);
DFFARX1 I_18114 (I12577,I2859,I310720,I310848,);
not I_18115 (I310856,I310848);
nor I_18116 (I310873,I310856,I310754);
and I_18117 (I310890,I310873,I12562);
nor I_18118 (I310907,I310856,I310822);
nor I_18119 (I310703,I310814,I310907);
DFFARX1 I_18120 (I12562,I2859,I310720,I310947,);
nor I_18121 (I310955,I310947,I310814);
not I_18122 (I310972,I310955);
not I_18123 (I310989,I310947);
nor I_18124 (I311006,I310989,I310890);
DFFARX1 I_18125 (I311006,I2859,I310720,I310706,);
nand I_18126 (I311037,I12580,I12565);
and I_18127 (I311054,I311037,I12583);
DFFARX1 I_18128 (I311054,I2859,I310720,I311080,);
nor I_18129 (I311088,I311080,I310947);
DFFARX1 I_18130 (I311088,I2859,I310720,I310688,);
nand I_18131 (I311119,I311080,I310989);
nand I_18132 (I310697,I310972,I311119);
not I_18133 (I311150,I311080);
nor I_18134 (I311167,I311150,I310890);
DFFARX1 I_18135 (I311167,I2859,I310720,I310709,);
nor I_18136 (I311198,I12574,I12565);
or I_18137 (I310700,I310947,I311198);
nor I_18138 (I310691,I311080,I311198);
or I_18139 (I310694,I310814,I311198);
DFFARX1 I_18140 (I311198,I2859,I310720,I310712,);
not I_18141 (I311298,I2866);
DFFARX1 I_18142 (I455274,I2859,I311298,I311324,);
not I_18143 (I311332,I311324);
nand I_18144 (I311349,I455256,I455268);
and I_18145 (I311366,I311349,I455271);
DFFARX1 I_18146 (I311366,I2859,I311298,I311392,);
not I_18147 (I311400,I455265);
DFFARX1 I_18148 (I455262,I2859,I311298,I311426,);
not I_18149 (I311434,I311426);
nor I_18150 (I311451,I311434,I311332);
and I_18151 (I311468,I311451,I455265);
nor I_18152 (I311485,I311434,I311400);
nor I_18153 (I311281,I311392,I311485);
DFFARX1 I_18154 (I455280,I2859,I311298,I311525,);
nor I_18155 (I311533,I311525,I311392);
not I_18156 (I311550,I311533);
not I_18157 (I311567,I311525);
nor I_18158 (I311584,I311567,I311468);
DFFARX1 I_18159 (I311584,I2859,I311298,I311284,);
nand I_18160 (I311615,I455259,I455259);
and I_18161 (I311632,I311615,I455256);
DFFARX1 I_18162 (I311632,I2859,I311298,I311658,);
nor I_18163 (I311666,I311658,I311525);
DFFARX1 I_18164 (I311666,I2859,I311298,I311266,);
nand I_18165 (I311697,I311658,I311567);
nand I_18166 (I311275,I311550,I311697);
not I_18167 (I311728,I311658);
nor I_18168 (I311745,I311728,I311468);
DFFARX1 I_18169 (I311745,I2859,I311298,I311287,);
nor I_18170 (I311776,I455277,I455259);
or I_18171 (I311278,I311525,I311776);
nor I_18172 (I311269,I311658,I311776);
or I_18173 (I311272,I311392,I311776);
DFFARX1 I_18174 (I311776,I2859,I311298,I311290,);
not I_18175 (I311876,I2866);
DFFARX1 I_18176 (I243062,I2859,I311876,I311902,);
not I_18177 (I311910,I311902);
nand I_18178 (I311927,I243071,I243080);
and I_18179 (I311944,I311927,I243086);
DFFARX1 I_18180 (I311944,I2859,I311876,I311970,);
not I_18181 (I311978,I243083);
DFFARX1 I_18182 (I243068,I2859,I311876,I312004,);
not I_18183 (I312012,I312004);
nor I_18184 (I312029,I312012,I311910);
and I_18185 (I312046,I312029,I243083);
nor I_18186 (I312063,I312012,I311978);
nor I_18187 (I311859,I311970,I312063);
DFFARX1 I_18188 (I243077,I2859,I311876,I312103,);
nor I_18189 (I312111,I312103,I311970);
not I_18190 (I312128,I312111);
not I_18191 (I312145,I312103);
nor I_18192 (I312162,I312145,I312046);
DFFARX1 I_18193 (I312162,I2859,I311876,I311862,);
nand I_18194 (I312193,I243074,I243065);
and I_18195 (I312210,I312193,I243062);
DFFARX1 I_18196 (I312210,I2859,I311876,I312236,);
nor I_18197 (I312244,I312236,I312103);
DFFARX1 I_18198 (I312244,I2859,I311876,I311844,);
nand I_18199 (I312275,I312236,I312145);
nand I_18200 (I311853,I312128,I312275);
not I_18201 (I312306,I312236);
nor I_18202 (I312323,I312306,I312046);
DFFARX1 I_18203 (I312323,I2859,I311876,I311865,);
nor I_18204 (I312354,I243065,I243065);
or I_18205 (I311856,I312103,I312354);
nor I_18206 (I311847,I312236,I312354);
or I_18207 (I311850,I311970,I312354);
DFFARX1 I_18208 (I312354,I2859,I311876,I311868,);
not I_18209 (I312454,I2866);
DFFARX1 I_18210 (I499202,I2859,I312454,I312480,);
not I_18211 (I312488,I312480);
nand I_18212 (I312505,I499184,I499196);
and I_18213 (I312522,I312505,I499199);
DFFARX1 I_18214 (I312522,I2859,I312454,I312548,);
not I_18215 (I312556,I499193);
DFFARX1 I_18216 (I499190,I2859,I312454,I312582,);
not I_18217 (I312590,I312582);
nor I_18218 (I312607,I312590,I312488);
and I_18219 (I312624,I312607,I499193);
nor I_18220 (I312641,I312590,I312556);
nor I_18221 (I312437,I312548,I312641);
DFFARX1 I_18222 (I499208,I2859,I312454,I312681,);
nor I_18223 (I312689,I312681,I312548);
not I_18224 (I312706,I312689);
not I_18225 (I312723,I312681);
nor I_18226 (I312740,I312723,I312624);
DFFARX1 I_18227 (I312740,I2859,I312454,I312440,);
nand I_18228 (I312771,I499187,I499187);
and I_18229 (I312788,I312771,I499184);
DFFARX1 I_18230 (I312788,I2859,I312454,I312814,);
nor I_18231 (I312822,I312814,I312681);
DFFARX1 I_18232 (I312822,I2859,I312454,I312422,);
nand I_18233 (I312853,I312814,I312723);
nand I_18234 (I312431,I312706,I312853);
not I_18235 (I312884,I312814);
nor I_18236 (I312901,I312884,I312624);
DFFARX1 I_18237 (I312901,I2859,I312454,I312443,);
nor I_18238 (I312932,I499205,I499187);
or I_18239 (I312434,I312681,I312932);
nor I_18240 (I312425,I312814,I312932);
or I_18241 (I312428,I312548,I312932);
DFFARX1 I_18242 (I312932,I2859,I312454,I312446,);
not I_18243 (I313032,I2866);
DFFARX1 I_18244 (I536140,I2859,I313032,I313058,);
not I_18245 (I313066,I313058);
nand I_18246 (I313083,I536128,I536146);
and I_18247 (I313100,I313083,I536137);
DFFARX1 I_18248 (I313100,I2859,I313032,I313126,);
not I_18249 (I313134,I536152);
DFFARX1 I_18250 (I536149,I2859,I313032,I313160,);
not I_18251 (I313168,I313160);
nor I_18252 (I313185,I313168,I313066);
and I_18253 (I313202,I313185,I536152);
nor I_18254 (I313219,I313168,I313134);
nor I_18255 (I313015,I313126,I313219);
DFFARX1 I_18256 (I536131,I2859,I313032,I313259,);
nor I_18257 (I313267,I313259,I313126);
not I_18258 (I313284,I313267);
not I_18259 (I313301,I313259);
nor I_18260 (I313318,I313301,I313202);
DFFARX1 I_18261 (I313318,I2859,I313032,I313018,);
nand I_18262 (I313349,I536125,I536125);
and I_18263 (I313366,I313349,I536134);
DFFARX1 I_18264 (I313366,I2859,I313032,I313392,);
nor I_18265 (I313400,I313392,I313259);
DFFARX1 I_18266 (I313400,I2859,I313032,I313000,);
nand I_18267 (I313431,I313392,I313301);
nand I_18268 (I313009,I313284,I313431);
not I_18269 (I313462,I313392);
nor I_18270 (I313479,I313462,I313202);
DFFARX1 I_18271 (I313479,I2859,I313032,I313021,);
nor I_18272 (I313510,I536143,I536125);
or I_18273 (I313012,I313259,I313510);
nor I_18274 (I313003,I313392,I313510);
or I_18275 (I313006,I313126,I313510);
DFFARX1 I_18276 (I313510,I2859,I313032,I313024,);
not I_18277 (I313610,I2866);
DFFARX1 I_18278 (I169988,I2859,I313610,I313636,);
not I_18279 (I313644,I313636);
nand I_18280 (I313661,I169979,I169997);
and I_18281 (I313678,I313661,I170000);
DFFARX1 I_18282 (I313678,I2859,I313610,I313704,);
not I_18283 (I313712,I169994);
DFFARX1 I_18284 (I169982,I2859,I313610,I313738,);
not I_18285 (I313746,I313738);
nor I_18286 (I313763,I313746,I313644);
and I_18287 (I313780,I313763,I169994);
nor I_18288 (I313797,I313746,I313712);
nor I_18289 (I313593,I313704,I313797);
DFFARX1 I_18290 (I169991,I2859,I313610,I313837,);
nor I_18291 (I313845,I313837,I313704);
not I_18292 (I313862,I313845);
not I_18293 (I313879,I313837);
nor I_18294 (I313896,I313879,I313780);
DFFARX1 I_18295 (I313896,I2859,I313610,I313596,);
nand I_18296 (I313927,I170006,I170003);
and I_18297 (I313944,I313927,I169985);
DFFARX1 I_18298 (I313944,I2859,I313610,I313970,);
nor I_18299 (I313978,I313970,I313837);
DFFARX1 I_18300 (I313978,I2859,I313610,I313578,);
nand I_18301 (I314009,I313970,I313879);
nand I_18302 (I313587,I313862,I314009);
not I_18303 (I314040,I313970);
nor I_18304 (I314057,I314040,I313780);
DFFARX1 I_18305 (I314057,I2859,I313610,I313599,);
nor I_18306 (I314088,I169979,I170003);
or I_18307 (I313590,I313837,I314088);
nor I_18308 (I313581,I313970,I314088);
or I_18309 (I313584,I313704,I314088);
DFFARX1 I_18310 (I314088,I2859,I313610,I313602,);
not I_18311 (I314188,I2866);
DFFARX1 I_18312 (I153530,I2859,I314188,I314214,);
not I_18313 (I314222,I314214);
nand I_18314 (I314239,I153533,I153509);
and I_18315 (I314256,I314239,I153506);
DFFARX1 I_18316 (I314256,I2859,I314188,I314282,);
not I_18317 (I314290,I153512);
DFFARX1 I_18318 (I153506,I2859,I314188,I314316,);
not I_18319 (I314324,I314316);
nor I_18320 (I314341,I314324,I314222);
and I_18321 (I314358,I314341,I153512);
nor I_18322 (I314375,I314324,I314290);
nor I_18323 (I314171,I314282,I314375);
DFFARX1 I_18324 (I153515,I2859,I314188,I314415,);
nor I_18325 (I314423,I314415,I314282);
not I_18326 (I314440,I314423);
not I_18327 (I314457,I314415);
nor I_18328 (I314474,I314457,I314358);
DFFARX1 I_18329 (I314474,I2859,I314188,I314174,);
nand I_18330 (I314505,I153518,I153527);
and I_18331 (I314522,I314505,I153524);
DFFARX1 I_18332 (I314522,I2859,I314188,I314548,);
nor I_18333 (I314556,I314548,I314415);
DFFARX1 I_18334 (I314556,I2859,I314188,I314156,);
nand I_18335 (I314587,I314548,I314457);
nand I_18336 (I314165,I314440,I314587);
not I_18337 (I314618,I314548);
nor I_18338 (I314635,I314618,I314358);
DFFARX1 I_18339 (I314635,I2859,I314188,I314177,);
nor I_18340 (I314666,I153521,I153527);
or I_18341 (I314168,I314415,I314666);
nor I_18342 (I314159,I314548,I314666);
or I_18343 (I314162,I314282,I314666);
DFFARX1 I_18344 (I314666,I2859,I314188,I314180,);
not I_18345 (I314766,I2866);
DFFARX1 I_18346 (I420991,I2859,I314766,I314792,);
not I_18347 (I314800,I314792);
nand I_18348 (I314817,I420967,I420982);
and I_18349 (I314834,I314817,I420994);
DFFARX1 I_18350 (I314834,I2859,I314766,I314860,);
not I_18351 (I314868,I420979);
DFFARX1 I_18352 (I420970,I2859,I314766,I314894,);
not I_18353 (I314902,I314894);
nor I_18354 (I314919,I314902,I314800);
and I_18355 (I314936,I314919,I420979);
nor I_18356 (I314953,I314902,I314868);
nor I_18357 (I314749,I314860,I314953);
DFFARX1 I_18358 (I420967,I2859,I314766,I314993,);
nor I_18359 (I315001,I314993,I314860);
not I_18360 (I315018,I315001);
not I_18361 (I315035,I314993);
nor I_18362 (I315052,I315035,I314936);
DFFARX1 I_18363 (I315052,I2859,I314766,I314752,);
nand I_18364 (I315083,I420985,I420976);
and I_18365 (I315100,I315083,I420988);
DFFARX1 I_18366 (I315100,I2859,I314766,I315126,);
nor I_18367 (I315134,I315126,I314993);
DFFARX1 I_18368 (I315134,I2859,I314766,I314734,);
nand I_18369 (I315165,I315126,I315035);
nand I_18370 (I314743,I315018,I315165);
not I_18371 (I315196,I315126);
nor I_18372 (I315213,I315196,I314936);
DFFARX1 I_18373 (I315213,I2859,I314766,I314755,);
nor I_18374 (I315244,I420973,I420976);
or I_18375 (I314746,I314993,I315244);
nor I_18376 (I314737,I315126,I315244);
or I_18377 (I314740,I314860,I315244);
DFFARX1 I_18378 (I315244,I2859,I314766,I314758,);
not I_18379 (I315344,I2866);
DFFARX1 I_18380 (I245952,I2859,I315344,I315370,);
not I_18381 (I315378,I315370);
nand I_18382 (I315395,I245961,I245970);
and I_18383 (I315412,I315395,I245976);
DFFARX1 I_18384 (I315412,I2859,I315344,I315438,);
not I_18385 (I315446,I245973);
DFFARX1 I_18386 (I245958,I2859,I315344,I315472,);
not I_18387 (I315480,I315472);
nor I_18388 (I315497,I315480,I315378);
and I_18389 (I315514,I315497,I245973);
nor I_18390 (I315531,I315480,I315446);
nor I_18391 (I315327,I315438,I315531);
DFFARX1 I_18392 (I245967,I2859,I315344,I315571,);
nor I_18393 (I315579,I315571,I315438);
not I_18394 (I315596,I315579);
not I_18395 (I315613,I315571);
nor I_18396 (I315630,I315613,I315514);
DFFARX1 I_18397 (I315630,I2859,I315344,I315330,);
nand I_18398 (I315661,I245964,I245955);
and I_18399 (I315678,I315661,I245952);
DFFARX1 I_18400 (I315678,I2859,I315344,I315704,);
nor I_18401 (I315712,I315704,I315571);
DFFARX1 I_18402 (I315712,I2859,I315344,I315312,);
nand I_18403 (I315743,I315704,I315613);
nand I_18404 (I315321,I315596,I315743);
not I_18405 (I315774,I315704);
nor I_18406 (I315791,I315774,I315514);
DFFARX1 I_18407 (I315791,I2859,I315344,I315333,);
nor I_18408 (I315822,I245955,I245955);
or I_18409 (I315324,I315571,I315822);
nor I_18410 (I315315,I315704,I315822);
or I_18411 (I315318,I315438,I315822);
DFFARX1 I_18412 (I315822,I2859,I315344,I315336,);
not I_18413 (I315922,I2866);
DFFARX1 I_18414 (I7301,I2859,I315922,I315948,);
not I_18415 (I315956,I315948);
nand I_18416 (I315973,I7298,I7289);
and I_18417 (I315990,I315973,I7289);
DFFARX1 I_18418 (I315990,I2859,I315922,I316016,);
not I_18419 (I316024,I7292);
DFFARX1 I_18420 (I7307,I2859,I315922,I316050,);
not I_18421 (I316058,I316050);
nor I_18422 (I316075,I316058,I315956);
and I_18423 (I316092,I316075,I7292);
nor I_18424 (I316109,I316058,I316024);
nor I_18425 (I315905,I316016,I316109);
DFFARX1 I_18426 (I7292,I2859,I315922,I316149,);
nor I_18427 (I316157,I316149,I316016);
not I_18428 (I316174,I316157);
not I_18429 (I316191,I316149);
nor I_18430 (I316208,I316191,I316092);
DFFARX1 I_18431 (I316208,I2859,I315922,I315908,);
nand I_18432 (I316239,I7310,I7295);
and I_18433 (I316256,I316239,I7313);
DFFARX1 I_18434 (I316256,I2859,I315922,I316282,);
nor I_18435 (I316290,I316282,I316149);
DFFARX1 I_18436 (I316290,I2859,I315922,I315890,);
nand I_18437 (I316321,I316282,I316191);
nand I_18438 (I315899,I316174,I316321);
not I_18439 (I316352,I316282);
nor I_18440 (I316369,I316352,I316092);
DFFARX1 I_18441 (I316369,I2859,I315922,I315911,);
nor I_18442 (I316400,I7304,I7295);
or I_18443 (I315902,I316149,I316400);
nor I_18444 (I315893,I316282,I316400);
or I_18445 (I315896,I316016,I316400);
DFFARX1 I_18446 (I316400,I2859,I315922,I315914,);
not I_18447 (I316500,I2866);
DFFARX1 I_18448 (I117167,I2859,I316500,I316526,);
not I_18449 (I316534,I316526);
nand I_18450 (I316551,I117170,I117146);
and I_18451 (I316568,I316551,I117143);
DFFARX1 I_18452 (I316568,I2859,I316500,I316594,);
not I_18453 (I316602,I117149);
DFFARX1 I_18454 (I117143,I2859,I316500,I316628,);
not I_18455 (I316636,I316628);
nor I_18456 (I316653,I316636,I316534);
and I_18457 (I316670,I316653,I117149);
nor I_18458 (I316687,I316636,I316602);
nor I_18459 (I316483,I316594,I316687);
DFFARX1 I_18460 (I117152,I2859,I316500,I316727,);
nor I_18461 (I316735,I316727,I316594);
not I_18462 (I316752,I316735);
not I_18463 (I316769,I316727);
nor I_18464 (I316786,I316769,I316670);
DFFARX1 I_18465 (I316786,I2859,I316500,I316486,);
nand I_18466 (I316817,I117155,I117164);
and I_18467 (I316834,I316817,I117161);
DFFARX1 I_18468 (I316834,I2859,I316500,I316860,);
nor I_18469 (I316868,I316860,I316727);
DFFARX1 I_18470 (I316868,I2859,I316500,I316468,);
nand I_18471 (I316899,I316860,I316769);
nand I_18472 (I316477,I316752,I316899);
not I_18473 (I316930,I316860);
nor I_18474 (I316947,I316930,I316670);
DFFARX1 I_18475 (I316947,I2859,I316500,I316489,);
nor I_18476 (I316978,I117158,I117164);
or I_18477 (I316480,I316727,I316978);
nor I_18478 (I316471,I316860,I316978);
or I_18479 (I316474,I316594,I316978);
DFFARX1 I_18480 (I316978,I2859,I316500,I316492,);
not I_18481 (I317078,I2866);
DFFARX1 I_18482 (I208612,I2859,I317078,I317104,);
not I_18483 (I317112,I317104);
nand I_18484 (I317129,I208603,I208621);
and I_18485 (I317146,I317129,I208624);
DFFARX1 I_18486 (I317146,I2859,I317078,I317172,);
not I_18487 (I317180,I208618);
DFFARX1 I_18488 (I208606,I2859,I317078,I317206,);
not I_18489 (I317214,I317206);
nor I_18490 (I317231,I317214,I317112);
and I_18491 (I317248,I317231,I208618);
nor I_18492 (I317265,I317214,I317180);
nor I_18493 (I317061,I317172,I317265);
DFFARX1 I_18494 (I208615,I2859,I317078,I317305,);
nor I_18495 (I317313,I317305,I317172);
not I_18496 (I317330,I317313);
not I_18497 (I317347,I317305);
nor I_18498 (I317364,I317347,I317248);
DFFARX1 I_18499 (I317364,I2859,I317078,I317064,);
nand I_18500 (I317395,I208630,I208627);
and I_18501 (I317412,I317395,I208609);
DFFARX1 I_18502 (I317412,I2859,I317078,I317438,);
nor I_18503 (I317446,I317438,I317305);
DFFARX1 I_18504 (I317446,I2859,I317078,I317046,);
nand I_18505 (I317477,I317438,I317347);
nand I_18506 (I317055,I317330,I317477);
not I_18507 (I317508,I317438);
nor I_18508 (I317525,I317508,I317248);
DFFARX1 I_18509 (I317525,I2859,I317078,I317067,);
nor I_18510 (I317556,I208603,I208627);
or I_18511 (I317058,I317305,I317556);
nor I_18512 (I317049,I317438,I317556);
or I_18513 (I317052,I317172,I317556);
DFFARX1 I_18514 (I317556,I2859,I317078,I317070,);
not I_18515 (I317656,I2866);
DFFARX1 I_18516 (I508058,I2859,I317656,I317682,);
not I_18517 (I317690,I317682);
nand I_18518 (I317707,I508061,I508070);
and I_18519 (I317724,I317707,I508073);
DFFARX1 I_18520 (I317724,I2859,I317656,I317750,);
not I_18521 (I317758,I508082);
DFFARX1 I_18522 (I508064,I2859,I317656,I317784,);
not I_18523 (I317792,I317784);
nor I_18524 (I317809,I317792,I317690);
and I_18525 (I317826,I317809,I508082);
nor I_18526 (I317843,I317792,I317758);
nor I_18527 (I317639,I317750,I317843);
DFFARX1 I_18528 (I508061,I2859,I317656,I317883,);
nor I_18529 (I317891,I317883,I317750);
not I_18530 (I317908,I317891);
not I_18531 (I317925,I317883);
nor I_18532 (I317942,I317925,I317826);
DFFARX1 I_18533 (I317942,I2859,I317656,I317642,);
nand I_18534 (I317973,I508079,I508058);
and I_18535 (I317990,I317973,I508076);
DFFARX1 I_18536 (I317990,I2859,I317656,I318016,);
nor I_18537 (I318024,I318016,I317883);
DFFARX1 I_18538 (I318024,I2859,I317656,I317624,);
nand I_18539 (I318055,I318016,I317925);
nand I_18540 (I317633,I317908,I318055);
not I_18541 (I318086,I318016);
nor I_18542 (I318103,I318086,I317826);
DFFARX1 I_18543 (I318103,I2859,I317656,I317645,);
nor I_18544 (I318134,I508067,I508058);
or I_18545 (I317636,I317883,I318134);
nor I_18546 (I317627,I318016,I318134);
or I_18547 (I317630,I317750,I318134);
DFFARX1 I_18548 (I318134,I2859,I317656,I317648,);
not I_18549 (I318234,I2866);
DFFARX1 I_18550 (I568112,I2859,I318234,I318260,);
not I_18551 (I318268,I318260);
nand I_18552 (I318285,I568097,I568085);
and I_18553 (I318302,I318285,I568100);
DFFARX1 I_18554 (I318302,I2859,I318234,I318328,);
not I_18555 (I318336,I568085);
DFFARX1 I_18556 (I568103,I2859,I318234,I318362,);
not I_18557 (I318370,I318362);
nor I_18558 (I318387,I318370,I318268);
and I_18559 (I318404,I318387,I568085);
nor I_18560 (I318421,I318370,I318336);
nor I_18561 (I318217,I318328,I318421);
DFFARX1 I_18562 (I568091,I2859,I318234,I318461,);
nor I_18563 (I318469,I318461,I318328);
not I_18564 (I318486,I318469);
not I_18565 (I318503,I318461);
nor I_18566 (I318520,I318503,I318404);
DFFARX1 I_18567 (I318520,I2859,I318234,I318220,);
nand I_18568 (I318551,I568088,I568094);
and I_18569 (I318568,I318551,I568109);
DFFARX1 I_18570 (I318568,I2859,I318234,I318594,);
nor I_18571 (I318602,I318594,I318461);
DFFARX1 I_18572 (I318602,I2859,I318234,I318202,);
nand I_18573 (I318633,I318594,I318503);
nand I_18574 (I318211,I318486,I318633);
not I_18575 (I318664,I318594);
nor I_18576 (I318681,I318664,I318404);
DFFARX1 I_18577 (I318681,I2859,I318234,I318223,);
nor I_18578 (I318712,I568106,I568094);
or I_18579 (I318214,I318461,I318712);
nor I_18580 (I318205,I318594,I318712);
or I_18581 (I318208,I318328,I318712);
DFFARX1 I_18582 (I318712,I2859,I318234,I318226,);
not I_18583 (I318812,I2866);
DFFARX1 I_18584 (I115059,I2859,I318812,I318838,);
not I_18585 (I318846,I318838);
nand I_18586 (I318863,I115062,I115038);
and I_18587 (I318880,I318863,I115035);
DFFARX1 I_18588 (I318880,I2859,I318812,I318906,);
not I_18589 (I318914,I115041);
DFFARX1 I_18590 (I115035,I2859,I318812,I318940,);
not I_18591 (I318948,I318940);
nor I_18592 (I318965,I318948,I318846);
and I_18593 (I318982,I318965,I115041);
nor I_18594 (I318999,I318948,I318914);
nor I_18595 (I318795,I318906,I318999);
DFFARX1 I_18596 (I115044,I2859,I318812,I319039,);
nor I_18597 (I319047,I319039,I318906);
not I_18598 (I319064,I319047);
not I_18599 (I319081,I319039);
nor I_18600 (I319098,I319081,I318982);
DFFARX1 I_18601 (I319098,I2859,I318812,I318798,);
nand I_18602 (I319129,I115047,I115056);
and I_18603 (I319146,I319129,I115053);
DFFARX1 I_18604 (I319146,I2859,I318812,I319172,);
nor I_18605 (I319180,I319172,I319039);
DFFARX1 I_18606 (I319180,I2859,I318812,I318780,);
nand I_18607 (I319211,I319172,I319081);
nand I_18608 (I318789,I319064,I319211);
not I_18609 (I319242,I319172);
nor I_18610 (I319259,I319242,I318982);
DFFARX1 I_18611 (I319259,I2859,I318812,I318801,);
nor I_18612 (I319290,I115050,I115056);
or I_18613 (I318792,I319039,I319290);
nor I_18614 (I318783,I319172,I319290);
or I_18615 (I318786,I318906,I319290);
DFFARX1 I_18616 (I319290,I2859,I318812,I318804,);
not I_18617 (I319390,I2866);
DFFARX1 I_18618 (I54195,I2859,I319390,I319416,);
not I_18619 (I319424,I319416);
nand I_18620 (I319441,I54204,I54213);
and I_18621 (I319458,I319441,I54192);
DFFARX1 I_18622 (I319458,I2859,I319390,I319484,);
not I_18623 (I319492,I54195);
DFFARX1 I_18624 (I54210,I2859,I319390,I319518,);
not I_18625 (I319526,I319518);
nor I_18626 (I319543,I319526,I319424);
and I_18627 (I319560,I319543,I54195);
nor I_18628 (I319577,I319526,I319492);
nor I_18629 (I319373,I319484,I319577);
DFFARX1 I_18630 (I54201,I2859,I319390,I319617,);
nor I_18631 (I319625,I319617,I319484);
not I_18632 (I319642,I319625);
not I_18633 (I319659,I319617);
nor I_18634 (I319676,I319659,I319560);
DFFARX1 I_18635 (I319676,I2859,I319390,I319376,);
nand I_18636 (I319707,I54216,I54192);
and I_18637 (I319724,I319707,I54198);
DFFARX1 I_18638 (I319724,I2859,I319390,I319750,);
nor I_18639 (I319758,I319750,I319617);
DFFARX1 I_18640 (I319758,I2859,I319390,I319358,);
nand I_18641 (I319789,I319750,I319659);
nand I_18642 (I319367,I319642,I319789);
not I_18643 (I319820,I319750);
nor I_18644 (I319837,I319820,I319560);
DFFARX1 I_18645 (I319837,I2859,I319390,I319379,);
nor I_18646 (I319868,I54207,I54192);
or I_18647 (I319370,I319617,I319868);
nor I_18648 (I319361,I319750,I319868);
or I_18649 (I319364,I319484,I319868);
DFFARX1 I_18650 (I319868,I2859,I319390,I319382,);
not I_18651 (I319968,I2866);
DFFARX1 I_18652 (I532096,I2859,I319968,I319994,);
not I_18653 (I320002,I319994);
nand I_18654 (I320019,I532120,I532102);
and I_18655 (I320036,I320019,I532108);
DFFARX1 I_18656 (I320036,I2859,I319968,I320062,);
not I_18657 (I320070,I532114);
DFFARX1 I_18658 (I532099,I2859,I319968,I320096,);
not I_18659 (I320104,I320096);
nor I_18660 (I320121,I320104,I320002);
and I_18661 (I320138,I320121,I532114);
nor I_18662 (I320155,I320104,I320070);
nor I_18663 (I319951,I320062,I320155);
DFFARX1 I_18664 (I532111,I2859,I319968,I320195,);
nor I_18665 (I320203,I320195,I320062);
not I_18666 (I320220,I320203);
not I_18667 (I320237,I320195);
nor I_18668 (I320254,I320237,I320138);
DFFARX1 I_18669 (I320254,I2859,I319968,I319954,);
nand I_18670 (I320285,I532117,I532105);
and I_18671 (I320302,I320285,I532099);
DFFARX1 I_18672 (I320302,I2859,I319968,I320328,);
nor I_18673 (I320336,I320328,I320195);
DFFARX1 I_18674 (I320336,I2859,I319968,I319936,);
nand I_18675 (I320367,I320328,I320237);
nand I_18676 (I319945,I320220,I320367);
not I_18677 (I320398,I320328);
nor I_18678 (I320415,I320398,I320138);
DFFARX1 I_18679 (I320415,I2859,I319968,I319957,);
nor I_18680 (I320446,I532096,I532105);
or I_18681 (I319948,I320195,I320446);
nor I_18682 (I319939,I320328,I320446);
or I_18683 (I319942,I320062,I320446);
DFFARX1 I_18684 (I320446,I2859,I319968,I319960,);
not I_18685 (I320546,I2866);
DFFARX1 I_18686 (I136666,I2859,I320546,I320572,);
not I_18687 (I320580,I320572);
nand I_18688 (I320597,I136669,I136645);
and I_18689 (I320614,I320597,I136642);
DFFARX1 I_18690 (I320614,I2859,I320546,I320640,);
not I_18691 (I320648,I136648);
DFFARX1 I_18692 (I136642,I2859,I320546,I320674,);
not I_18693 (I320682,I320674);
nor I_18694 (I320699,I320682,I320580);
and I_18695 (I320716,I320699,I136648);
nor I_18696 (I320733,I320682,I320648);
nor I_18697 (I320529,I320640,I320733);
DFFARX1 I_18698 (I136651,I2859,I320546,I320773,);
nor I_18699 (I320781,I320773,I320640);
not I_18700 (I320798,I320781);
not I_18701 (I320815,I320773);
nor I_18702 (I320832,I320815,I320716);
DFFARX1 I_18703 (I320832,I2859,I320546,I320532,);
nand I_18704 (I320863,I136654,I136663);
and I_18705 (I320880,I320863,I136660);
DFFARX1 I_18706 (I320880,I2859,I320546,I320906,);
nor I_18707 (I320914,I320906,I320773);
DFFARX1 I_18708 (I320914,I2859,I320546,I320514,);
nand I_18709 (I320945,I320906,I320815);
nand I_18710 (I320523,I320798,I320945);
not I_18711 (I320976,I320906);
nor I_18712 (I320993,I320976,I320716);
DFFARX1 I_18713 (I320993,I2859,I320546,I320535,);
nor I_18714 (I321024,I136657,I136663);
or I_18715 (I320526,I320773,I321024);
nor I_18716 (I320517,I320906,I321024);
or I_18717 (I320520,I320640,I321024);
DFFARX1 I_18718 (I321024,I2859,I320546,I320538,);
not I_18719 (I321124,I2866);
DFFARX1 I_18720 (I467412,I2859,I321124,I321150,);
not I_18721 (I321158,I321150);
nand I_18722 (I321175,I467394,I467406);
and I_18723 (I321192,I321175,I467409);
DFFARX1 I_18724 (I321192,I2859,I321124,I321218,);
not I_18725 (I321226,I467403);
DFFARX1 I_18726 (I467400,I2859,I321124,I321252,);
not I_18727 (I321260,I321252);
nor I_18728 (I321277,I321260,I321158);
and I_18729 (I321294,I321277,I467403);
nor I_18730 (I321311,I321260,I321226);
nor I_18731 (I321107,I321218,I321311);
DFFARX1 I_18732 (I467418,I2859,I321124,I321351,);
nor I_18733 (I321359,I321351,I321218);
not I_18734 (I321376,I321359);
not I_18735 (I321393,I321351);
nor I_18736 (I321410,I321393,I321294);
DFFARX1 I_18737 (I321410,I2859,I321124,I321110,);
nand I_18738 (I321441,I467397,I467397);
and I_18739 (I321458,I321441,I467394);
DFFARX1 I_18740 (I321458,I2859,I321124,I321484,);
nor I_18741 (I321492,I321484,I321351);
DFFARX1 I_18742 (I321492,I2859,I321124,I321092,);
nand I_18743 (I321523,I321484,I321393);
nand I_18744 (I321101,I321376,I321523);
not I_18745 (I321554,I321484);
nor I_18746 (I321571,I321554,I321294);
DFFARX1 I_18747 (I321571,I2859,I321124,I321113,);
nor I_18748 (I321602,I467415,I467397);
or I_18749 (I321104,I321351,I321602);
nor I_18750 (I321095,I321484,I321602);
or I_18751 (I321098,I321218,I321602);
DFFARX1 I_18752 (I321602,I2859,I321124,I321116,);
not I_18753 (I321702,I2866);
DFFARX1 I_18754 (I466834,I2859,I321702,I321728,);
not I_18755 (I321736,I321728);
nand I_18756 (I321753,I466816,I466828);
and I_18757 (I321770,I321753,I466831);
DFFARX1 I_18758 (I321770,I2859,I321702,I321796,);
not I_18759 (I321804,I466825);
DFFARX1 I_18760 (I466822,I2859,I321702,I321830,);
not I_18761 (I321838,I321830);
nor I_18762 (I321855,I321838,I321736);
and I_18763 (I321872,I321855,I466825);
nor I_18764 (I321889,I321838,I321804);
nor I_18765 (I321685,I321796,I321889);
DFFARX1 I_18766 (I466840,I2859,I321702,I321929,);
nor I_18767 (I321937,I321929,I321796);
not I_18768 (I321954,I321937);
not I_18769 (I321971,I321929);
nor I_18770 (I321988,I321971,I321872);
DFFARX1 I_18771 (I321988,I2859,I321702,I321688,);
nand I_18772 (I322019,I466819,I466819);
and I_18773 (I322036,I322019,I466816);
DFFARX1 I_18774 (I322036,I2859,I321702,I322062,);
nor I_18775 (I322070,I322062,I321929);
DFFARX1 I_18776 (I322070,I2859,I321702,I321670,);
nand I_18777 (I322101,I322062,I321971);
nand I_18778 (I321679,I321954,I322101);
not I_18779 (I322132,I322062);
nor I_18780 (I322149,I322132,I321872);
DFFARX1 I_18781 (I322149,I2859,I321702,I321691,);
nor I_18782 (I322180,I466837,I466819);
or I_18783 (I321682,I321929,I322180);
nor I_18784 (I321673,I322062,I322180);
or I_18785 (I321676,I321796,I322180);
DFFARX1 I_18786 (I322180,I2859,I321702,I321694,);
not I_18787 (I322280,I2866);
DFFARX1 I_18788 (I143517,I2859,I322280,I322306,);
not I_18789 (I322314,I322306);
nand I_18790 (I322331,I143520,I143496);
and I_18791 (I322348,I322331,I143493);
DFFARX1 I_18792 (I322348,I2859,I322280,I322374,);
not I_18793 (I322382,I143499);
DFFARX1 I_18794 (I143493,I2859,I322280,I322408,);
not I_18795 (I322416,I322408);
nor I_18796 (I322433,I322416,I322314);
and I_18797 (I322450,I322433,I143499);
nor I_18798 (I322467,I322416,I322382);
nor I_18799 (I322263,I322374,I322467);
DFFARX1 I_18800 (I143502,I2859,I322280,I322507,);
nor I_18801 (I322515,I322507,I322374);
not I_18802 (I322532,I322515);
not I_18803 (I322549,I322507);
nor I_18804 (I322566,I322549,I322450);
DFFARX1 I_18805 (I322566,I2859,I322280,I322266,);
nand I_18806 (I322597,I143505,I143514);
and I_18807 (I322614,I322597,I143511);
DFFARX1 I_18808 (I322614,I2859,I322280,I322640,);
nor I_18809 (I322648,I322640,I322507);
DFFARX1 I_18810 (I322648,I2859,I322280,I322248,);
nand I_18811 (I322679,I322640,I322549);
nand I_18812 (I322257,I322532,I322679);
not I_18813 (I322710,I322640);
nor I_18814 (I322727,I322710,I322450);
DFFARX1 I_18815 (I322727,I2859,I322280,I322269,);
nor I_18816 (I322758,I143508,I143514);
or I_18817 (I322260,I322507,I322758);
nor I_18818 (I322251,I322640,I322758);
or I_18819 (I322254,I322374,I322758);
DFFARX1 I_18820 (I322758,I2859,I322280,I322272,);
not I_18821 (I322858,I2866);
DFFARX1 I_18822 (I15206,I2859,I322858,I322884,);
not I_18823 (I322892,I322884);
nand I_18824 (I322909,I15203,I15194);
and I_18825 (I322926,I322909,I15194);
DFFARX1 I_18826 (I322926,I2859,I322858,I322952,);
not I_18827 (I322960,I15197);
DFFARX1 I_18828 (I15212,I2859,I322858,I322986,);
not I_18829 (I322994,I322986);
nor I_18830 (I323011,I322994,I322892);
and I_18831 (I323028,I323011,I15197);
nor I_18832 (I323045,I322994,I322960);
nor I_18833 (I322841,I322952,I323045);
DFFARX1 I_18834 (I15197,I2859,I322858,I323085,);
nor I_18835 (I323093,I323085,I322952);
not I_18836 (I323110,I323093);
not I_18837 (I323127,I323085);
nor I_18838 (I323144,I323127,I323028);
DFFARX1 I_18839 (I323144,I2859,I322858,I322844,);
nand I_18840 (I323175,I15215,I15200);
and I_18841 (I323192,I323175,I15218);
DFFARX1 I_18842 (I323192,I2859,I322858,I323218,);
nor I_18843 (I323226,I323218,I323085);
DFFARX1 I_18844 (I323226,I2859,I322858,I322826,);
nand I_18845 (I323257,I323218,I323127);
nand I_18846 (I322835,I323110,I323257);
not I_18847 (I323288,I323218);
nor I_18848 (I323305,I323288,I323028);
DFFARX1 I_18849 (I323305,I2859,I322858,I322847,);
nor I_18850 (I323336,I15209,I15200);
or I_18851 (I322838,I323085,I323336);
nor I_18852 (I322829,I323218,I323336);
or I_18853 (I322832,I322952,I323336);
DFFARX1 I_18854 (I323336,I2859,I322858,I322850,);
not I_18855 (I323436,I2866);
DFFARX1 I_18856 (I233236,I2859,I323436,I323462,);
not I_18857 (I323470,I323462);
nand I_18858 (I323487,I233245,I233254);
and I_18859 (I323504,I323487,I233260);
DFFARX1 I_18860 (I323504,I2859,I323436,I323530,);
not I_18861 (I323538,I233257);
DFFARX1 I_18862 (I233242,I2859,I323436,I323564,);
not I_18863 (I323572,I323564);
nor I_18864 (I323589,I323572,I323470);
and I_18865 (I323606,I323589,I233257);
nor I_18866 (I323623,I323572,I323538);
nor I_18867 (I323419,I323530,I323623);
DFFARX1 I_18868 (I233251,I2859,I323436,I323663,);
nor I_18869 (I323671,I323663,I323530);
not I_18870 (I323688,I323671);
not I_18871 (I323705,I323663);
nor I_18872 (I323722,I323705,I323606);
DFFARX1 I_18873 (I323722,I2859,I323436,I323422,);
nand I_18874 (I323753,I233248,I233239);
and I_18875 (I323770,I323753,I233236);
DFFARX1 I_18876 (I323770,I2859,I323436,I323796,);
nor I_18877 (I323804,I323796,I323663);
DFFARX1 I_18878 (I323804,I2859,I323436,I323404,);
nand I_18879 (I323835,I323796,I323705);
nand I_18880 (I323413,I323688,I323835);
not I_18881 (I323866,I323796);
nor I_18882 (I323883,I323866,I323606);
DFFARX1 I_18883 (I323883,I2859,I323436,I323425,);
nor I_18884 (I323914,I233239,I233239);
or I_18885 (I323416,I323663,I323914);
nor I_18886 (I323407,I323796,I323914);
or I_18887 (I323410,I323530,I323914);
DFFARX1 I_18888 (I323914,I2859,I323436,I323428,);
not I_18889 (I324014,I2866);
DFFARX1 I_18890 (I1532,I2859,I324014,I324040,);
not I_18891 (I324048,I324040);
nand I_18892 (I324065,I2580,I1852);
and I_18893 (I324082,I324065,I1652);
DFFARX1 I_18894 (I324082,I2859,I324014,I324108,);
not I_18895 (I324116,I1660);
DFFARX1 I_18896 (I2796,I2859,I324014,I324142,);
not I_18897 (I324150,I324142);
nor I_18898 (I324167,I324150,I324048);
and I_18899 (I324184,I324167,I1660);
nor I_18900 (I324201,I324150,I324116);
nor I_18901 (I323997,I324108,I324201);
DFFARX1 I_18902 (I2596,I2859,I324014,I324241,);
nor I_18903 (I324249,I324241,I324108);
not I_18904 (I324266,I324249);
not I_18905 (I324283,I324241);
nor I_18906 (I324300,I324283,I324184);
DFFARX1 I_18907 (I324300,I2859,I324014,I324000,);
nand I_18908 (I324331,I2396,I2156);
and I_18909 (I324348,I324331,I2124);
DFFARX1 I_18910 (I324348,I2859,I324014,I324374,);
nor I_18911 (I324382,I324374,I324241);
DFFARX1 I_18912 (I324382,I2859,I324014,I323982,);
nand I_18913 (I324413,I324374,I324283);
nand I_18914 (I323991,I324266,I324413);
not I_18915 (I324444,I324374);
nor I_18916 (I324461,I324444,I324184);
DFFARX1 I_18917 (I324461,I2859,I324014,I324003,);
nor I_18918 (I324492,I2076,I2156);
or I_18919 (I323994,I324241,I324492);
nor I_18920 (I323985,I324374,I324492);
or I_18921 (I323988,I324108,I324492);
DFFARX1 I_18922 (I324492,I2859,I324014,I324006,);
not I_18923 (I324592,I2866);
DFFARX1 I_18924 (I457008,I2859,I324592,I324618,);
not I_18925 (I324626,I324618);
nand I_18926 (I324643,I456990,I457002);
and I_18927 (I324660,I324643,I457005);
DFFARX1 I_18928 (I324660,I2859,I324592,I324686,);
not I_18929 (I324694,I456999);
DFFARX1 I_18930 (I456996,I2859,I324592,I324720,);
not I_18931 (I324728,I324720);
nor I_18932 (I324745,I324728,I324626);
and I_18933 (I324762,I324745,I456999);
nor I_18934 (I324779,I324728,I324694);
nor I_18935 (I324575,I324686,I324779);
DFFARX1 I_18936 (I457014,I2859,I324592,I324819,);
nor I_18937 (I324827,I324819,I324686);
not I_18938 (I324844,I324827);
not I_18939 (I324861,I324819);
nor I_18940 (I324878,I324861,I324762);
DFFARX1 I_18941 (I324878,I2859,I324592,I324578,);
nand I_18942 (I324909,I456993,I456993);
and I_18943 (I324926,I324909,I456990);
DFFARX1 I_18944 (I324926,I2859,I324592,I324952,);
nor I_18945 (I324960,I324952,I324819);
DFFARX1 I_18946 (I324960,I2859,I324592,I324560,);
nand I_18947 (I324991,I324952,I324861);
nand I_18948 (I324569,I324844,I324991);
not I_18949 (I325022,I324952);
nor I_18950 (I325039,I325022,I324762);
DFFARX1 I_18951 (I325039,I2859,I324592,I324581,);
nor I_18952 (I325070,I457011,I456993);
or I_18953 (I324572,I324819,I325070);
nor I_18954 (I324563,I324952,I325070);
or I_18955 (I324566,I324686,I325070);
DFFARX1 I_18956 (I325070,I2859,I324592,I324584,);
not I_18957 (I325170,I2866);
DFFARX1 I_18958 (I428691,I2859,I325170,I325196,);
not I_18959 (I325204,I325196);
nand I_18960 (I325221,I428688,I428706);
and I_18961 (I325238,I325221,I428703);
DFFARX1 I_18962 (I325238,I2859,I325170,I325264,);
not I_18963 (I325272,I428685);
DFFARX1 I_18964 (I428688,I2859,I325170,I325298,);
not I_18965 (I325306,I325298);
nor I_18966 (I325323,I325306,I325204);
and I_18967 (I325340,I325323,I428685);
nor I_18968 (I325357,I325306,I325272);
nor I_18969 (I325153,I325264,I325357);
DFFARX1 I_18970 (I428697,I2859,I325170,I325397,);
nor I_18971 (I325405,I325397,I325264);
not I_18972 (I325422,I325405);
not I_18973 (I325439,I325397);
nor I_18974 (I325456,I325439,I325340);
DFFARX1 I_18975 (I325456,I2859,I325170,I325156,);
nand I_18976 (I325487,I428700,I428685);
and I_18977 (I325504,I325487,I428691);
DFFARX1 I_18978 (I325504,I2859,I325170,I325530,);
nor I_18979 (I325538,I325530,I325397);
DFFARX1 I_18980 (I325538,I2859,I325170,I325138,);
nand I_18981 (I325569,I325530,I325439);
nand I_18982 (I325147,I325422,I325569);
not I_18983 (I325600,I325530);
nor I_18984 (I325617,I325600,I325340);
DFFARX1 I_18985 (I325617,I2859,I325170,I325159,);
nor I_18986 (I325648,I428694,I428685);
or I_18987 (I325150,I325397,I325648);
nor I_18988 (I325141,I325530,I325648);
or I_18989 (I325144,I325264,I325648);
DFFARX1 I_18990 (I325648,I2859,I325170,I325162,);
not I_18991 (I325748,I2866);
DFFARX1 I_18992 (I114005,I2859,I325748,I325774,);
not I_18993 (I325782,I325774);
nand I_18994 (I325799,I114008,I113984);
and I_18995 (I325816,I325799,I113981);
DFFARX1 I_18996 (I325816,I2859,I325748,I325842,);
not I_18997 (I325850,I113987);
DFFARX1 I_18998 (I113981,I2859,I325748,I325876,);
not I_18999 (I325884,I325876);
nor I_19000 (I325901,I325884,I325782);
and I_19001 (I325918,I325901,I113987);
nor I_19002 (I325935,I325884,I325850);
nor I_19003 (I325731,I325842,I325935);
DFFARX1 I_19004 (I113990,I2859,I325748,I325975,);
nor I_19005 (I325983,I325975,I325842);
not I_19006 (I326000,I325983);
not I_19007 (I326017,I325975);
nor I_19008 (I326034,I326017,I325918);
DFFARX1 I_19009 (I326034,I2859,I325748,I325734,);
nand I_19010 (I326065,I113993,I114002);
and I_19011 (I326082,I326065,I113999);
DFFARX1 I_19012 (I326082,I2859,I325748,I326108,);
nor I_19013 (I326116,I326108,I325975);
DFFARX1 I_19014 (I326116,I2859,I325748,I325716,);
nand I_19015 (I326147,I326108,I326017);
nand I_19016 (I325725,I326000,I326147);
not I_19017 (I326178,I326108);
nor I_19018 (I326195,I326178,I325918);
DFFARX1 I_19019 (I326195,I2859,I325748,I325737,);
nor I_19020 (I326226,I113996,I114002);
or I_19021 (I325728,I325975,I326226);
nor I_19022 (I325719,I326108,I326226);
or I_19023 (I325722,I325842,I326226);
DFFARX1 I_19024 (I326226,I2859,I325748,I325740,);
not I_19025 (I326326,I2866);
DFFARX1 I_19026 (I383523,I2859,I326326,I326352,);
not I_19027 (I326360,I326352);
nand I_19028 (I326377,I383499,I383514);
and I_19029 (I326394,I326377,I383526);
DFFARX1 I_19030 (I326394,I2859,I326326,I326420,);
not I_19031 (I326428,I383511);
DFFARX1 I_19032 (I383502,I2859,I326326,I326454,);
not I_19033 (I326462,I326454);
nor I_19034 (I326479,I326462,I326360);
and I_19035 (I326496,I326479,I383511);
nor I_19036 (I326513,I326462,I326428);
nor I_19037 (I326309,I326420,I326513);
DFFARX1 I_19038 (I383499,I2859,I326326,I326553,);
nor I_19039 (I326561,I326553,I326420);
not I_19040 (I326578,I326561);
not I_19041 (I326595,I326553);
nor I_19042 (I326612,I326595,I326496);
DFFARX1 I_19043 (I326612,I2859,I326326,I326312,);
nand I_19044 (I326643,I383517,I383508);
and I_19045 (I326660,I326643,I383520);
DFFARX1 I_19046 (I326660,I2859,I326326,I326686,);
nor I_19047 (I326694,I326686,I326553);
DFFARX1 I_19048 (I326694,I2859,I326326,I326294,);
nand I_19049 (I326725,I326686,I326595);
nand I_19050 (I326303,I326578,I326725);
not I_19051 (I326756,I326686);
nor I_19052 (I326773,I326756,I326496);
DFFARX1 I_19053 (I326773,I2859,I326326,I326315,);
nor I_19054 (I326804,I383505,I383508);
or I_19055 (I326306,I326553,I326804);
nor I_19056 (I326297,I326686,I326804);
or I_19057 (I326300,I326420,I326804);
DFFARX1 I_19058 (I326804,I2859,I326326,I326318,);
not I_19059 (I326904,I2866);
DFFARX1 I_19060 (I170532,I2859,I326904,I326930,);
not I_19061 (I326938,I326930);
nand I_19062 (I326955,I170523,I170541);
and I_19063 (I326972,I326955,I170544);
DFFARX1 I_19064 (I326972,I2859,I326904,I326998,);
not I_19065 (I327006,I170538);
DFFARX1 I_19066 (I170526,I2859,I326904,I327032,);
not I_19067 (I327040,I327032);
nor I_19068 (I327057,I327040,I326938);
and I_19069 (I327074,I327057,I170538);
nor I_19070 (I327091,I327040,I327006);
nor I_19071 (I326887,I326998,I327091);
DFFARX1 I_19072 (I170535,I2859,I326904,I327131,);
nor I_19073 (I327139,I327131,I326998);
not I_19074 (I327156,I327139);
not I_19075 (I327173,I327131);
nor I_19076 (I327190,I327173,I327074);
DFFARX1 I_19077 (I327190,I2859,I326904,I326890,);
nand I_19078 (I327221,I170550,I170547);
and I_19079 (I327238,I327221,I170529);
DFFARX1 I_19080 (I327238,I2859,I326904,I327264,);
nor I_19081 (I327272,I327264,I327131);
DFFARX1 I_19082 (I327272,I2859,I326904,I326872,);
nand I_19083 (I327303,I327264,I327173);
nand I_19084 (I326881,I327156,I327303);
not I_19085 (I327334,I327264);
nor I_19086 (I327351,I327334,I327074);
DFFARX1 I_19087 (I327351,I2859,I326904,I326893,);
nor I_19088 (I327382,I170523,I170547);
or I_19089 (I326884,I327131,I327382);
nor I_19090 (I326875,I327264,I327382);
or I_19091 (I326878,I326998,I327382);
DFFARX1 I_19092 (I327382,I2859,I326904,I326896,);
not I_19093 (I327482,I2866);
DFFARX1 I_19094 (I38385,I2859,I327482,I327508,);
not I_19095 (I327516,I327508);
nand I_19096 (I327533,I38394,I38403);
and I_19097 (I327550,I327533,I38382);
DFFARX1 I_19098 (I327550,I2859,I327482,I327576,);
not I_19099 (I327584,I38385);
DFFARX1 I_19100 (I38400,I2859,I327482,I327610,);
not I_19101 (I327618,I327610);
nor I_19102 (I327635,I327618,I327516);
and I_19103 (I327652,I327635,I38385);
nor I_19104 (I327669,I327618,I327584);
nor I_19105 (I327465,I327576,I327669);
DFFARX1 I_19106 (I38391,I2859,I327482,I327709,);
nor I_19107 (I327717,I327709,I327576);
not I_19108 (I327734,I327717);
not I_19109 (I327751,I327709);
nor I_19110 (I327768,I327751,I327652);
DFFARX1 I_19111 (I327768,I2859,I327482,I327468,);
nand I_19112 (I327799,I38406,I38382);
and I_19113 (I327816,I327799,I38388);
DFFARX1 I_19114 (I327816,I2859,I327482,I327842,);
nor I_19115 (I327850,I327842,I327709);
DFFARX1 I_19116 (I327850,I2859,I327482,I327450,);
nand I_19117 (I327881,I327842,I327751);
nand I_19118 (I327459,I327734,I327881);
not I_19119 (I327912,I327842);
nor I_19120 (I327929,I327912,I327652);
DFFARX1 I_19121 (I327929,I2859,I327482,I327471,);
nor I_19122 (I327960,I38397,I38382);
or I_19123 (I327462,I327709,I327960);
nor I_19124 (I327453,I327842,I327960);
or I_19125 (I327456,I327576,I327960);
DFFARX1 I_19126 (I327960,I2859,I327482,I327474,);
not I_19127 (I328060,I2866);
DFFARX1 I_19128 (I25737,I2859,I328060,I328086,);
not I_19129 (I328094,I328086);
nand I_19130 (I328111,I25746,I25755);
and I_19131 (I328128,I328111,I25734);
DFFARX1 I_19132 (I328128,I2859,I328060,I328154,);
not I_19133 (I328162,I25737);
DFFARX1 I_19134 (I25752,I2859,I328060,I328188,);
not I_19135 (I328196,I328188);
nor I_19136 (I328213,I328196,I328094);
and I_19137 (I328230,I328213,I25737);
nor I_19138 (I328247,I328196,I328162);
nor I_19139 (I328043,I328154,I328247);
DFFARX1 I_19140 (I25743,I2859,I328060,I328287,);
nor I_19141 (I328295,I328287,I328154);
not I_19142 (I328312,I328295);
not I_19143 (I328329,I328287);
nor I_19144 (I328346,I328329,I328230);
DFFARX1 I_19145 (I328346,I2859,I328060,I328046,);
nand I_19146 (I328377,I25758,I25734);
and I_19147 (I328394,I328377,I25740);
DFFARX1 I_19148 (I328394,I2859,I328060,I328420,);
nor I_19149 (I328428,I328420,I328287);
DFFARX1 I_19150 (I328428,I2859,I328060,I328028,);
nand I_19151 (I328459,I328420,I328329);
nand I_19152 (I328037,I328312,I328459);
not I_19153 (I328490,I328420);
nor I_19154 (I328507,I328490,I328230);
DFFARX1 I_19155 (I328507,I2859,I328060,I328049,);
nor I_19156 (I328538,I25749,I25734);
or I_19157 (I328040,I328287,I328538);
nor I_19158 (I328031,I328420,I328538);
or I_19159 (I328034,I328154,I328538);
DFFARX1 I_19160 (I328538,I2859,I328060,I328052,);
not I_19161 (I328638,I2866);
DFFARX1 I_19162 (I259246,I2859,I328638,I328664,);
not I_19163 (I328672,I328664);
nand I_19164 (I328689,I259255,I259264);
and I_19165 (I328706,I328689,I259270);
DFFARX1 I_19166 (I328706,I2859,I328638,I328732,);
not I_19167 (I328740,I259267);
DFFARX1 I_19168 (I259252,I2859,I328638,I328766,);
not I_19169 (I328774,I328766);
nor I_19170 (I328791,I328774,I328672);
and I_19171 (I328808,I328791,I259267);
nor I_19172 (I328825,I328774,I328740);
nor I_19173 (I328621,I328732,I328825);
DFFARX1 I_19174 (I259261,I2859,I328638,I328865,);
nor I_19175 (I328873,I328865,I328732);
not I_19176 (I328890,I328873);
not I_19177 (I328907,I328865);
nor I_19178 (I328924,I328907,I328808);
DFFARX1 I_19179 (I328924,I2859,I328638,I328624,);
nand I_19180 (I328955,I259258,I259249);
and I_19181 (I328972,I328955,I259246);
DFFARX1 I_19182 (I328972,I2859,I328638,I328998,);
nor I_19183 (I329006,I328998,I328865);
DFFARX1 I_19184 (I329006,I2859,I328638,I328606,);
nand I_19185 (I329037,I328998,I328907);
nand I_19186 (I328615,I328890,I329037);
not I_19187 (I329068,I328998);
nor I_19188 (I329085,I329068,I328808);
DFFARX1 I_19189 (I329085,I2859,I328638,I328627,);
nor I_19190 (I329116,I259249,I259249);
or I_19191 (I328618,I328865,I329116);
nor I_19192 (I328609,I328998,I329116);
or I_19193 (I328612,I328732,I329116);
DFFARX1 I_19194 (I329116,I2859,I328638,I328630,);
not I_19195 (I329216,I2866);
DFFARX1 I_19196 (I394505,I2859,I329216,I329242,);
not I_19197 (I329250,I329242);
nand I_19198 (I329267,I394481,I394496);
and I_19199 (I329284,I329267,I394508);
DFFARX1 I_19200 (I329284,I2859,I329216,I329310,);
not I_19201 (I329318,I394493);
DFFARX1 I_19202 (I394484,I2859,I329216,I329344,);
not I_19203 (I329352,I329344);
nor I_19204 (I329369,I329352,I329250);
and I_19205 (I329386,I329369,I394493);
nor I_19206 (I329403,I329352,I329318);
nor I_19207 (I329199,I329310,I329403);
DFFARX1 I_19208 (I394481,I2859,I329216,I329443,);
nor I_19209 (I329451,I329443,I329310);
not I_19210 (I329468,I329451);
not I_19211 (I329485,I329443);
nor I_19212 (I329502,I329485,I329386);
DFFARX1 I_19213 (I329502,I2859,I329216,I329202,);
nand I_19214 (I329533,I394499,I394490);
and I_19215 (I329550,I329533,I394502);
DFFARX1 I_19216 (I329550,I2859,I329216,I329576,);
nor I_19217 (I329584,I329576,I329443);
DFFARX1 I_19218 (I329584,I2859,I329216,I329184,);
nand I_19219 (I329615,I329576,I329485);
nand I_19220 (I329193,I329468,I329615);
not I_19221 (I329646,I329576);
nor I_19222 (I329663,I329646,I329386);
DFFARX1 I_19223 (I329663,I2859,I329216,I329205,);
nor I_19224 (I329694,I394487,I394490);
or I_19225 (I329196,I329443,I329694);
nor I_19226 (I329187,I329576,I329694);
or I_19227 (I329190,I329310,I329694);
DFFARX1 I_19228 (I329694,I2859,I329216,I329208,);
not I_19229 (I329794,I2866);
DFFARX1 I_19230 (I42074,I2859,I329794,I329820,);
not I_19231 (I329828,I329820);
nand I_19232 (I329845,I42083,I42092);
and I_19233 (I329862,I329845,I42071);
DFFARX1 I_19234 (I329862,I2859,I329794,I329888,);
not I_19235 (I329896,I42074);
DFFARX1 I_19236 (I42089,I2859,I329794,I329922,);
not I_19237 (I329930,I329922);
nor I_19238 (I329947,I329930,I329828);
and I_19239 (I329964,I329947,I42074);
nor I_19240 (I329981,I329930,I329896);
nor I_19241 (I329777,I329888,I329981);
DFFARX1 I_19242 (I42080,I2859,I329794,I330021,);
nor I_19243 (I330029,I330021,I329888);
not I_19244 (I330046,I330029);
not I_19245 (I330063,I330021);
nor I_19246 (I330080,I330063,I329964);
DFFARX1 I_19247 (I330080,I2859,I329794,I329780,);
nand I_19248 (I330111,I42095,I42071);
and I_19249 (I330128,I330111,I42077);
DFFARX1 I_19250 (I330128,I2859,I329794,I330154,);
nor I_19251 (I330162,I330154,I330021);
DFFARX1 I_19252 (I330162,I2859,I329794,I329762,);
nand I_19253 (I330193,I330154,I330063);
nand I_19254 (I329771,I330046,I330193);
not I_19255 (I330224,I330154);
nor I_19256 (I330241,I330224,I329964);
DFFARX1 I_19257 (I330241,I2859,I329794,I329783,);
nor I_19258 (I330272,I42086,I42071);
or I_19259 (I329774,I330021,I330272);
nor I_19260 (I329765,I330154,I330272);
or I_19261 (I329768,I329888,I330272);
DFFARX1 I_19262 (I330272,I2859,I329794,I329786,);
not I_19263 (I330372,I2866);
DFFARX1 I_19264 (I362179,I2859,I330372,I330398,);
not I_19265 (I330406,I330398);
nand I_19266 (I330423,I362167,I362185);
and I_19267 (I330440,I330423,I362182);
DFFARX1 I_19268 (I330440,I2859,I330372,I330466,);
not I_19269 (I330474,I362173);
DFFARX1 I_19270 (I362170,I2859,I330372,I330500,);
not I_19271 (I330508,I330500);
nor I_19272 (I330525,I330508,I330406);
and I_19273 (I330542,I330525,I362173);
nor I_19274 (I330559,I330508,I330474);
nor I_19275 (I330355,I330466,I330559);
DFFARX1 I_19276 (I362164,I2859,I330372,I330599,);
nor I_19277 (I330607,I330599,I330466);
not I_19278 (I330624,I330607);
not I_19279 (I330641,I330599);
nor I_19280 (I330658,I330641,I330542);
DFFARX1 I_19281 (I330658,I2859,I330372,I330358,);
nand I_19282 (I330689,I362164,I362167);
and I_19283 (I330706,I330689,I362170);
DFFARX1 I_19284 (I330706,I2859,I330372,I330732,);
nor I_19285 (I330740,I330732,I330599);
DFFARX1 I_19286 (I330740,I2859,I330372,I330340,);
nand I_19287 (I330771,I330732,I330641);
nand I_19288 (I330349,I330624,I330771);
not I_19289 (I330802,I330732);
nor I_19290 (I330819,I330802,I330542);
DFFARX1 I_19291 (I330819,I2859,I330372,I330361,);
nor I_19292 (I330850,I362176,I362167);
or I_19293 (I330352,I330599,I330850);
nor I_19294 (I330343,I330732,I330850);
or I_19295 (I330346,I330466,I330850);
DFFARX1 I_19296 (I330850,I2859,I330372,I330364,);
not I_19297 (I330950,I2866);
DFFARX1 I_19298 (I381585,I2859,I330950,I330976,);
not I_19299 (I330984,I330976);
nand I_19300 (I331001,I381561,I381576);
and I_19301 (I331018,I331001,I381588);
DFFARX1 I_19302 (I331018,I2859,I330950,I331044,);
not I_19303 (I331052,I381573);
DFFARX1 I_19304 (I381564,I2859,I330950,I331078,);
not I_19305 (I331086,I331078);
nor I_19306 (I331103,I331086,I330984);
and I_19307 (I331120,I331103,I381573);
nor I_19308 (I331137,I331086,I331052);
nor I_19309 (I330933,I331044,I331137);
DFFARX1 I_19310 (I381561,I2859,I330950,I331177,);
nor I_19311 (I331185,I331177,I331044);
not I_19312 (I331202,I331185);
not I_19313 (I331219,I331177);
nor I_19314 (I331236,I331219,I331120);
DFFARX1 I_19315 (I331236,I2859,I330950,I330936,);
nand I_19316 (I331267,I381579,I381570);
and I_19317 (I331284,I331267,I381582);
DFFARX1 I_19318 (I331284,I2859,I330950,I331310,);
nor I_19319 (I331318,I331310,I331177);
DFFARX1 I_19320 (I331318,I2859,I330950,I330918,);
nand I_19321 (I331349,I331310,I331219);
nand I_19322 (I330927,I331202,I331349);
not I_19323 (I331380,I331310);
nor I_19324 (I331397,I331380,I331120);
DFFARX1 I_19325 (I331397,I2859,I330950,I330939,);
nor I_19326 (I331428,I381567,I381570);
or I_19327 (I330930,I331177,I331428);
nor I_19328 (I330921,I331310,I331428);
or I_19329 (I330924,I331044,I331428);
DFFARX1 I_19330 (I331428,I2859,I330950,I330942,);
not I_19331 (I331528,I2866);
DFFARX1 I_19332 (I355855,I2859,I331528,I331554,);
not I_19333 (I331562,I331554);
nand I_19334 (I331579,I355843,I355861);
and I_19335 (I331596,I331579,I355858);
DFFARX1 I_19336 (I331596,I2859,I331528,I331622,);
not I_19337 (I331630,I355849);
DFFARX1 I_19338 (I355846,I2859,I331528,I331656,);
not I_19339 (I331664,I331656);
nor I_19340 (I331681,I331664,I331562);
and I_19341 (I331698,I331681,I355849);
nor I_19342 (I331715,I331664,I331630);
nor I_19343 (I331511,I331622,I331715);
DFFARX1 I_19344 (I355840,I2859,I331528,I331755,);
nor I_19345 (I331763,I331755,I331622);
not I_19346 (I331780,I331763);
not I_19347 (I331797,I331755);
nor I_19348 (I331814,I331797,I331698);
DFFARX1 I_19349 (I331814,I2859,I331528,I331514,);
nand I_19350 (I331845,I355840,I355843);
and I_19351 (I331862,I331845,I355846);
DFFARX1 I_19352 (I331862,I2859,I331528,I331888,);
nor I_19353 (I331896,I331888,I331755);
DFFARX1 I_19354 (I331896,I2859,I331528,I331496,);
nand I_19355 (I331927,I331888,I331797);
nand I_19356 (I331505,I331780,I331927);
not I_19357 (I331958,I331888);
nor I_19358 (I331975,I331958,I331698);
DFFARX1 I_19359 (I331975,I2859,I331528,I331517,);
nor I_19360 (I332006,I355852,I355843);
or I_19361 (I331508,I331755,I332006);
nor I_19362 (I331499,I331888,I332006);
or I_19363 (I331502,I331622,I332006);
DFFARX1 I_19364 (I332006,I2859,I331528,I331520,);
not I_19365 (I332106,I2866);
DFFARX1 I_19366 (I408071,I2859,I332106,I332132,);
not I_19367 (I332140,I332132);
nand I_19368 (I332157,I408047,I408062);
and I_19369 (I332174,I332157,I408074);
DFFARX1 I_19370 (I332174,I2859,I332106,I332200,);
not I_19371 (I332208,I408059);
DFFARX1 I_19372 (I408050,I2859,I332106,I332234,);
not I_19373 (I332242,I332234);
nor I_19374 (I332259,I332242,I332140);
and I_19375 (I332276,I332259,I408059);
nor I_19376 (I332293,I332242,I332208);
nor I_19377 (I332089,I332200,I332293);
DFFARX1 I_19378 (I408047,I2859,I332106,I332333,);
nor I_19379 (I332341,I332333,I332200);
not I_19380 (I332358,I332341);
not I_19381 (I332375,I332333);
nor I_19382 (I332392,I332375,I332276);
DFFARX1 I_19383 (I332392,I2859,I332106,I332092,);
nand I_19384 (I332423,I408065,I408056);
and I_19385 (I332440,I332423,I408068);
DFFARX1 I_19386 (I332440,I2859,I332106,I332466,);
nor I_19387 (I332474,I332466,I332333);
DFFARX1 I_19388 (I332474,I2859,I332106,I332074,);
nand I_19389 (I332505,I332466,I332375);
nand I_19390 (I332083,I332358,I332505);
not I_19391 (I332536,I332466);
nor I_19392 (I332553,I332536,I332276);
DFFARX1 I_19393 (I332553,I2859,I332106,I332095,);
nor I_19394 (I332584,I408053,I408056);
or I_19395 (I332086,I332333,I332584);
nor I_19396 (I332077,I332466,I332584);
or I_19397 (I332080,I332200,I332584);
DFFARX1 I_19398 (I332584,I2859,I332106,I332098,);
not I_19399 (I332681,I2866);
DFFARX1 I_19400 (I461632,I2859,I332681,I332707,);
not I_19401 (I332715,I332707);
nand I_19402 (I332732,I461614,I461614);
and I_19403 (I332749,I332732,I461620);
DFFARX1 I_19404 (I332749,I2859,I332681,I332775,);
DFFARX1 I_19405 (I332775,I2859,I332681,I332670,);
DFFARX1 I_19406 (I461617,I2859,I332681,I332806,);
nand I_19407 (I332814,I332806,I461626);
not I_19408 (I332831,I332814);
DFFARX1 I_19409 (I332831,I2859,I332681,I332857,);
not I_19410 (I332865,I332857);
nor I_19411 (I332673,I332715,I332865);
DFFARX1 I_19412 (I461638,I2859,I332681,I332905,);
nor I_19413 (I332664,I332905,I332775);
nor I_19414 (I332655,I332905,I332831);
nand I_19415 (I332941,I461629,I461623);
and I_19416 (I332958,I332941,I461617);
DFFARX1 I_19417 (I332958,I2859,I332681,I332984,);
not I_19418 (I332992,I332984);
nand I_19419 (I333009,I332992,I332905);
nand I_19420 (I332658,I332992,I332814);
nor I_19421 (I333040,I461635,I461623);
and I_19422 (I333057,I332905,I333040);
nor I_19423 (I333074,I332992,I333057);
DFFARX1 I_19424 (I333074,I2859,I332681,I332667,);
nor I_19425 (I333105,I332707,I333040);
DFFARX1 I_19426 (I333105,I2859,I332681,I332652,);
nor I_19427 (I333136,I332984,I333040);
not I_19428 (I333153,I333136);
nand I_19429 (I332661,I333153,I333009);
not I_19430 (I333208,I2866);
DFFARX1 I_19431 (I460476,I2859,I333208,I333234,);
not I_19432 (I333242,I333234);
nand I_19433 (I333259,I460458,I460458);
and I_19434 (I333276,I333259,I460464);
DFFARX1 I_19435 (I333276,I2859,I333208,I333302,);
DFFARX1 I_19436 (I333302,I2859,I333208,I333197,);
DFFARX1 I_19437 (I460461,I2859,I333208,I333333,);
nand I_19438 (I333341,I333333,I460470);
not I_19439 (I333358,I333341);
DFFARX1 I_19440 (I333358,I2859,I333208,I333384,);
not I_19441 (I333392,I333384);
nor I_19442 (I333200,I333242,I333392);
DFFARX1 I_19443 (I460482,I2859,I333208,I333432,);
nor I_19444 (I333191,I333432,I333302);
nor I_19445 (I333182,I333432,I333358);
nand I_19446 (I333468,I460473,I460467);
and I_19447 (I333485,I333468,I460461);
DFFARX1 I_19448 (I333485,I2859,I333208,I333511,);
not I_19449 (I333519,I333511);
nand I_19450 (I333536,I333519,I333432);
nand I_19451 (I333185,I333519,I333341);
nor I_19452 (I333567,I460479,I460467);
and I_19453 (I333584,I333432,I333567);
nor I_19454 (I333601,I333519,I333584);
DFFARX1 I_19455 (I333601,I2859,I333208,I333194,);
nor I_19456 (I333632,I333234,I333567);
DFFARX1 I_19457 (I333632,I2859,I333208,I333179,);
nor I_19458 (I333663,I333511,I333567);
not I_19459 (I333680,I333663);
nand I_19460 (I333188,I333680,I333536);
not I_19461 (I333735,I2866);
DFFARX1 I_19462 (I217874,I2859,I333735,I333761,);
not I_19463 (I333769,I333761);
nand I_19464 (I333786,I217892,I217883);
and I_19465 (I333803,I333786,I217886);
DFFARX1 I_19466 (I333803,I2859,I333735,I333829,);
DFFARX1 I_19467 (I333829,I2859,I333735,I333724,);
DFFARX1 I_19468 (I217880,I2859,I333735,I333860,);
nand I_19469 (I333868,I333860,I217871);
not I_19470 (I333885,I333868);
DFFARX1 I_19471 (I333885,I2859,I333735,I333911,);
not I_19472 (I333919,I333911);
nor I_19473 (I333727,I333769,I333919);
DFFARX1 I_19474 (I217877,I2859,I333735,I333959,);
nor I_19475 (I333718,I333959,I333829);
nor I_19476 (I333709,I333959,I333885);
nand I_19477 (I333995,I217871,I217868);
and I_19478 (I334012,I333995,I217889);
DFFARX1 I_19479 (I334012,I2859,I333735,I334038,);
not I_19480 (I334046,I334038);
nand I_19481 (I334063,I334046,I333959);
nand I_19482 (I333712,I334046,I333868);
nor I_19483 (I334094,I217868,I217868);
and I_19484 (I334111,I333959,I334094);
nor I_19485 (I334128,I334046,I334111);
DFFARX1 I_19486 (I334128,I2859,I333735,I333721,);
nor I_19487 (I334159,I333761,I334094);
DFFARX1 I_19488 (I334159,I2859,I333735,I333706,);
nor I_19489 (I334190,I334038,I334094);
not I_19490 (I334207,I334190);
nand I_19491 (I333715,I334207,I334063);
not I_19492 (I334262,I2866);
DFFARX1 I_19493 (I20473,I2859,I334262,I334288,);
not I_19494 (I334296,I334288);
nand I_19495 (I334313,I20485,I20488);
and I_19496 (I334330,I334313,I20464);
DFFARX1 I_19497 (I334330,I2859,I334262,I334356,);
DFFARX1 I_19498 (I334356,I2859,I334262,I334251,);
DFFARX1 I_19499 (I20482,I2859,I334262,I334387,);
nand I_19500 (I334395,I334387,I20470);
not I_19501 (I334412,I334395);
DFFARX1 I_19502 (I334412,I2859,I334262,I334438,);
not I_19503 (I334446,I334438);
nor I_19504 (I334254,I334296,I334446);
DFFARX1 I_19505 (I20467,I2859,I334262,I334486,);
nor I_19506 (I334245,I334486,I334356);
nor I_19507 (I334236,I334486,I334412);
nand I_19508 (I334522,I20476,I20467);
and I_19509 (I334539,I334522,I20464);
DFFARX1 I_19510 (I334539,I2859,I334262,I334565,);
not I_19511 (I334573,I334565);
nand I_19512 (I334590,I334573,I334486);
nand I_19513 (I334239,I334573,I334395);
nor I_19514 (I334621,I20479,I20467);
and I_19515 (I334638,I334486,I334621);
nor I_19516 (I334655,I334573,I334638);
DFFARX1 I_19517 (I334655,I2859,I334262,I334248,);
nor I_19518 (I334686,I334288,I334621);
DFFARX1 I_19519 (I334686,I2859,I334262,I334233,);
nor I_19520 (I334717,I334565,I334621);
not I_19521 (I334734,I334717);
nand I_19522 (I334242,I334734,I334590);
not I_19523 (I334789,I2866);
DFFARX1 I_19524 (I270228,I2859,I334789,I334815,);
not I_19525 (I334823,I334815);
nand I_19526 (I334840,I270231,I270228);
and I_19527 (I334857,I334840,I270240);
DFFARX1 I_19528 (I334857,I2859,I334789,I334883,);
DFFARX1 I_19529 (I334883,I2859,I334789,I334778,);
DFFARX1 I_19530 (I270237,I2859,I334789,I334914,);
nand I_19531 (I334922,I334914,I270243);
not I_19532 (I334939,I334922);
DFFARX1 I_19533 (I334939,I2859,I334789,I334965,);
not I_19534 (I334973,I334965);
nor I_19535 (I334781,I334823,I334973);
DFFARX1 I_19536 (I270252,I2859,I334789,I335013,);
nor I_19537 (I334772,I335013,I334883);
nor I_19538 (I334763,I335013,I334939);
nand I_19539 (I335049,I270246,I270234);
and I_19540 (I335066,I335049,I270231);
DFFARX1 I_19541 (I335066,I2859,I334789,I335092,);
not I_19542 (I335100,I335092);
nand I_19543 (I335117,I335100,I335013);
nand I_19544 (I334766,I335100,I334922);
nor I_19545 (I335148,I270249,I270234);
and I_19546 (I335165,I335013,I335148);
nor I_19547 (I335182,I335100,I335165);
DFFARX1 I_19548 (I335182,I2859,I334789,I334775,);
nor I_19549 (I335213,I334815,I335148);
DFFARX1 I_19550 (I335213,I2859,I334789,I334760,);
nor I_19551 (I335244,I335092,I335148);
not I_19552 (I335261,I335244);
nand I_19553 (I334769,I335261,I335117);
not I_19554 (I335316,I2866);
DFFARX1 I_19555 (I149826,I2859,I335316,I335342,);
not I_19556 (I335350,I335342);
nand I_19557 (I335367,I149817,I149817);
and I_19558 (I335384,I335367,I149835);
DFFARX1 I_19559 (I335384,I2859,I335316,I335410,);
DFFARX1 I_19560 (I335410,I2859,I335316,I335305,);
DFFARX1 I_19561 (I149838,I2859,I335316,I335441,);
nand I_19562 (I335449,I335441,I149820);
not I_19563 (I335466,I335449);
DFFARX1 I_19564 (I335466,I2859,I335316,I335492,);
not I_19565 (I335500,I335492);
nor I_19566 (I335308,I335350,I335500);
DFFARX1 I_19567 (I149832,I2859,I335316,I335540,);
nor I_19568 (I335299,I335540,I335410);
nor I_19569 (I335290,I335540,I335466);
nand I_19570 (I335576,I149844,I149823);
and I_19571 (I335593,I335576,I149829);
DFFARX1 I_19572 (I335593,I2859,I335316,I335619,);
not I_19573 (I335627,I335619);
nand I_19574 (I335644,I335627,I335540);
nand I_19575 (I335293,I335627,I335449);
nor I_19576 (I335675,I149841,I149823);
and I_19577 (I335692,I335540,I335675);
nor I_19578 (I335709,I335627,I335692);
DFFARX1 I_19579 (I335709,I2859,I335316,I335302,);
nor I_19580 (I335740,I335342,I335675);
DFFARX1 I_19581 (I335740,I2859,I335316,I335287,);
nor I_19582 (I335771,I335619,I335675);
not I_19583 (I335788,I335771);
nand I_19584 (I335296,I335788,I335644);
not I_19585 (I335843,I2866);
DFFARX1 I_19586 (I300284,I2859,I335843,I335869,);
not I_19587 (I335877,I335869);
nand I_19588 (I335894,I300287,I300284);
and I_19589 (I335911,I335894,I300296);
DFFARX1 I_19590 (I335911,I2859,I335843,I335937,);
DFFARX1 I_19591 (I335937,I2859,I335843,I335832,);
DFFARX1 I_19592 (I300293,I2859,I335843,I335968,);
nand I_19593 (I335976,I335968,I300299);
not I_19594 (I335993,I335976);
DFFARX1 I_19595 (I335993,I2859,I335843,I336019,);
not I_19596 (I336027,I336019);
nor I_19597 (I335835,I335877,I336027);
DFFARX1 I_19598 (I300308,I2859,I335843,I336067,);
nor I_19599 (I335826,I336067,I335937);
nor I_19600 (I335817,I336067,I335993);
nand I_19601 (I336103,I300302,I300290);
and I_19602 (I336120,I336103,I300287);
DFFARX1 I_19603 (I336120,I2859,I335843,I336146,);
not I_19604 (I336154,I336146);
nand I_19605 (I336171,I336154,I336067);
nand I_19606 (I335820,I336154,I335976);
nor I_19607 (I336202,I300305,I300290);
and I_19608 (I336219,I336067,I336202);
nor I_19609 (I336236,I336154,I336219);
DFFARX1 I_19610 (I336236,I2859,I335843,I335829,);
nor I_19611 (I336267,I335869,I336202);
DFFARX1 I_19612 (I336267,I2859,I335843,I335814,);
nor I_19613 (I336298,I336146,I336202);
not I_19614 (I336315,I336298);
nand I_19615 (I335823,I336315,I336171);
not I_19616 (I336370,I2866);
DFFARX1 I_19617 (I225014,I2859,I336370,I336396,);
not I_19618 (I336404,I336396);
nand I_19619 (I336421,I225032,I225023);
and I_19620 (I336438,I336421,I225026);
DFFARX1 I_19621 (I336438,I2859,I336370,I336464,);
DFFARX1 I_19622 (I336464,I2859,I336370,I336359,);
DFFARX1 I_19623 (I225020,I2859,I336370,I336495,);
nand I_19624 (I336503,I336495,I225011);
not I_19625 (I336520,I336503);
DFFARX1 I_19626 (I336520,I2859,I336370,I336546,);
not I_19627 (I336554,I336546);
nor I_19628 (I336362,I336404,I336554);
DFFARX1 I_19629 (I225017,I2859,I336370,I336594,);
nor I_19630 (I336353,I336594,I336464);
nor I_19631 (I336344,I336594,I336520);
nand I_19632 (I336630,I225011,I225008);
and I_19633 (I336647,I336630,I225029);
DFFARX1 I_19634 (I336647,I2859,I336370,I336673,);
not I_19635 (I336681,I336673);
nand I_19636 (I336698,I336681,I336594);
nand I_19637 (I336347,I336681,I336503);
nor I_19638 (I336729,I225008,I225008);
and I_19639 (I336746,I336594,I336729);
nor I_19640 (I336763,I336681,I336746);
DFFARX1 I_19641 (I336763,I2859,I336370,I336356,);
nor I_19642 (I336794,I336396,I336729);
DFFARX1 I_19643 (I336794,I2859,I336370,I336341,);
nor I_19644 (I336825,I336673,I336729);
not I_19645 (I336842,I336825);
nand I_19646 (I336350,I336842,I336698);
not I_19647 (I336897,I2866);
DFFARX1 I_19648 (I116625,I2859,I336897,I336923,);
not I_19649 (I336931,I336923);
nand I_19650 (I336948,I116616,I116616);
and I_19651 (I336965,I336948,I116634);
DFFARX1 I_19652 (I336965,I2859,I336897,I336991,);
DFFARX1 I_19653 (I336991,I2859,I336897,I336886,);
DFFARX1 I_19654 (I116637,I2859,I336897,I337022,);
nand I_19655 (I337030,I337022,I116619);
not I_19656 (I337047,I337030);
DFFARX1 I_19657 (I337047,I2859,I336897,I337073,);
not I_19658 (I337081,I337073);
nor I_19659 (I336889,I336931,I337081);
DFFARX1 I_19660 (I116631,I2859,I336897,I337121,);
nor I_19661 (I336880,I337121,I336991);
nor I_19662 (I336871,I337121,I337047);
nand I_19663 (I337157,I116643,I116622);
and I_19664 (I337174,I337157,I116628);
DFFARX1 I_19665 (I337174,I2859,I336897,I337200,);
not I_19666 (I337208,I337200);
nand I_19667 (I337225,I337208,I337121);
nand I_19668 (I336874,I337208,I337030);
nor I_19669 (I337256,I116640,I116622);
and I_19670 (I337273,I337121,I337256);
nor I_19671 (I337290,I337208,I337273);
DFFARX1 I_19672 (I337290,I2859,I336897,I336883,);
nor I_19673 (I337321,I336923,I337256);
DFFARX1 I_19674 (I337321,I2859,I336897,I336868,);
nor I_19675 (I337352,I337200,I337256);
not I_19676 (I337369,I337352);
nand I_19677 (I336877,I337369,I337225);
not I_19678 (I337424,I2866);
DFFARX1 I_19679 (I325716,I2859,I337424,I337450,);
not I_19680 (I337458,I337450);
nand I_19681 (I337475,I325719,I325716);
and I_19682 (I337492,I337475,I325728);
DFFARX1 I_19683 (I337492,I2859,I337424,I337518,);
DFFARX1 I_19684 (I337518,I2859,I337424,I337413,);
DFFARX1 I_19685 (I325725,I2859,I337424,I337549,);
nand I_19686 (I337557,I337549,I325731);
not I_19687 (I337574,I337557);
DFFARX1 I_19688 (I337574,I2859,I337424,I337600,);
not I_19689 (I337608,I337600);
nor I_19690 (I337416,I337458,I337608);
DFFARX1 I_19691 (I325740,I2859,I337424,I337648,);
nor I_19692 (I337407,I337648,I337518);
nor I_19693 (I337398,I337648,I337574);
nand I_19694 (I337684,I325734,I325722);
and I_19695 (I337701,I337684,I325719);
DFFARX1 I_19696 (I337701,I2859,I337424,I337727,);
not I_19697 (I337735,I337727);
nand I_19698 (I337752,I337735,I337648);
nand I_19699 (I337401,I337735,I337557);
nor I_19700 (I337783,I325737,I325722);
and I_19701 (I337800,I337648,I337783);
nor I_19702 (I337817,I337735,I337800);
DFFARX1 I_19703 (I337817,I2859,I337424,I337410,);
nor I_19704 (I337848,I337450,I337783);
DFFARX1 I_19705 (I337848,I2859,I337424,I337395,);
nor I_19706 (I337879,I337727,I337783);
not I_19707 (I337896,I337879);
nand I_19708 (I337404,I337896,I337752);
not I_19709 (I337951,I2866);
DFFARX1 I_19710 (I133489,I2859,I337951,I337977,);
not I_19711 (I337985,I337977);
nand I_19712 (I338002,I133480,I133480);
and I_19713 (I338019,I338002,I133498);
DFFARX1 I_19714 (I338019,I2859,I337951,I338045,);
DFFARX1 I_19715 (I338045,I2859,I337951,I337940,);
DFFARX1 I_19716 (I133501,I2859,I337951,I338076,);
nand I_19717 (I338084,I338076,I133483);
not I_19718 (I338101,I338084);
DFFARX1 I_19719 (I338101,I2859,I337951,I338127,);
not I_19720 (I338135,I338127);
nor I_19721 (I337943,I337985,I338135);
DFFARX1 I_19722 (I133495,I2859,I337951,I338175,);
nor I_19723 (I337934,I338175,I338045);
nor I_19724 (I337925,I338175,I338101);
nand I_19725 (I338211,I133507,I133486);
and I_19726 (I338228,I338211,I133492);
DFFARX1 I_19727 (I338228,I2859,I337951,I338254,);
not I_19728 (I338262,I338254);
nand I_19729 (I338279,I338262,I338175);
nand I_19730 (I337928,I338262,I338084);
nor I_19731 (I338310,I133504,I133486);
and I_19732 (I338327,I338175,I338310);
nor I_19733 (I338344,I338262,I338327);
DFFARX1 I_19734 (I338344,I2859,I337951,I337937,);
nor I_19735 (I338375,I337977,I338310);
DFFARX1 I_19736 (I338375,I2859,I337951,I337922,);
nor I_19737 (I338406,I338254,I338310);
not I_19738 (I338423,I338406);
nand I_19739 (I337931,I338423,I338279);
not I_19740 (I338478,I2866);
DFFARX1 I_19741 (I319936,I2859,I338478,I338504,);
not I_19742 (I338512,I338504);
nand I_19743 (I338529,I319939,I319936);
and I_19744 (I338546,I338529,I319948);
DFFARX1 I_19745 (I338546,I2859,I338478,I338572,);
DFFARX1 I_19746 (I338572,I2859,I338478,I338467,);
DFFARX1 I_19747 (I319945,I2859,I338478,I338603,);
nand I_19748 (I338611,I338603,I319951);
not I_19749 (I338628,I338611);
DFFARX1 I_19750 (I338628,I2859,I338478,I338654,);
not I_19751 (I338662,I338654);
nor I_19752 (I338470,I338512,I338662);
DFFARX1 I_19753 (I319960,I2859,I338478,I338702,);
nor I_19754 (I338461,I338702,I338572);
nor I_19755 (I338452,I338702,I338628);
nand I_19756 (I338738,I319954,I319942);
and I_19757 (I338755,I338738,I319939);
DFFARX1 I_19758 (I338755,I2859,I338478,I338781,);
not I_19759 (I338789,I338781);
nand I_19760 (I338806,I338789,I338702);
nand I_19761 (I338455,I338789,I338611);
nor I_19762 (I338837,I319957,I319942);
and I_19763 (I338854,I338702,I338837);
nor I_19764 (I338871,I338789,I338854);
DFFARX1 I_19765 (I338871,I2859,I338478,I338464,);
nor I_19766 (I338902,I338504,I338837);
DFFARX1 I_19767 (I338902,I2859,I338478,I338449,);
nor I_19768 (I338933,I338781,I338837);
not I_19769 (I338950,I338933);
nand I_19770 (I338458,I338950,I338806);
not I_19771 (I339005,I2866);
DFFARX1 I_19772 (I417094,I2859,I339005,I339031,);
not I_19773 (I339039,I339031);
nand I_19774 (I339056,I417109,I417091);
and I_19775 (I339073,I339056,I417091);
DFFARX1 I_19776 (I339073,I2859,I339005,I339099,);
DFFARX1 I_19777 (I339099,I2859,I339005,I338994,);
DFFARX1 I_19778 (I417100,I2859,I339005,I339130,);
nand I_19779 (I339138,I339130,I417118);
not I_19780 (I339155,I339138);
DFFARX1 I_19781 (I339155,I2859,I339005,I339181,);
not I_19782 (I339189,I339181);
nor I_19783 (I338997,I339039,I339189);
DFFARX1 I_19784 (I417115,I2859,I339005,I339229,);
nor I_19785 (I338988,I339229,I339099);
nor I_19786 (I338979,I339229,I339155);
nand I_19787 (I339265,I417112,I417103);
and I_19788 (I339282,I339265,I417097);
DFFARX1 I_19789 (I339282,I2859,I339005,I339308,);
not I_19790 (I339316,I339308);
nand I_19791 (I339333,I339316,I339229);
nand I_19792 (I338982,I339316,I339138);
nor I_19793 (I339364,I417106,I417103);
and I_19794 (I339381,I339229,I339364);
nor I_19795 (I339398,I339316,I339381);
DFFARX1 I_19796 (I339398,I2859,I339005,I338991,);
nor I_19797 (I339429,I339031,I339364);
DFFARX1 I_19798 (I339429,I2859,I339005,I338976,);
nor I_19799 (I339460,I339308,I339364);
not I_19800 (I339477,I339460);
nand I_19801 (I338985,I339477,I339333);
not I_19802 (I339532,I2866);
DFFARX1 I_19803 (I278898,I2859,I339532,I339558,);
not I_19804 (I339566,I339558);
nand I_19805 (I339583,I278901,I278898);
and I_19806 (I339600,I339583,I278910);
DFFARX1 I_19807 (I339600,I2859,I339532,I339626,);
DFFARX1 I_19808 (I339626,I2859,I339532,I339521,);
DFFARX1 I_19809 (I278907,I2859,I339532,I339657,);
nand I_19810 (I339665,I339657,I278913);
not I_19811 (I339682,I339665);
DFFARX1 I_19812 (I339682,I2859,I339532,I339708,);
not I_19813 (I339716,I339708);
nor I_19814 (I339524,I339566,I339716);
DFFARX1 I_19815 (I278922,I2859,I339532,I339756,);
nor I_19816 (I339515,I339756,I339626);
nor I_19817 (I339506,I339756,I339682);
nand I_19818 (I339792,I278916,I278904);
and I_19819 (I339809,I339792,I278901);
DFFARX1 I_19820 (I339809,I2859,I339532,I339835,);
not I_19821 (I339843,I339835);
nand I_19822 (I339860,I339843,I339756);
nand I_19823 (I339509,I339843,I339665);
nor I_19824 (I339891,I278919,I278904);
and I_19825 (I339908,I339756,I339891);
nor I_19826 (I339925,I339843,I339908);
DFFARX1 I_19827 (I339925,I2859,I339532,I339518,);
nor I_19828 (I339956,I339558,I339891);
DFFARX1 I_19829 (I339956,I2859,I339532,I339503,);
nor I_19830 (I339987,I339835,I339891);
not I_19831 (I340004,I339987);
nand I_19832 (I339512,I340004,I339860);
not I_19833 (I340059,I2866);
DFFARX1 I_19834 (I159839,I2859,I340059,I340085,);
not I_19835 (I340093,I340085);
nand I_19836 (I340110,I159830,I159830);
and I_19837 (I340127,I340110,I159848);
DFFARX1 I_19838 (I340127,I2859,I340059,I340153,);
DFFARX1 I_19839 (I340153,I2859,I340059,I340048,);
DFFARX1 I_19840 (I159851,I2859,I340059,I340184,);
nand I_19841 (I340192,I340184,I159833);
not I_19842 (I340209,I340192);
DFFARX1 I_19843 (I340209,I2859,I340059,I340235,);
not I_19844 (I340243,I340235);
nor I_19845 (I340051,I340093,I340243);
DFFARX1 I_19846 (I159845,I2859,I340059,I340283,);
nor I_19847 (I340042,I340283,I340153);
nor I_19848 (I340033,I340283,I340209);
nand I_19849 (I340319,I159857,I159836);
and I_19850 (I340336,I340319,I159842);
DFFARX1 I_19851 (I340336,I2859,I340059,I340362,);
not I_19852 (I340370,I340362);
nand I_19853 (I340387,I340370,I340283);
nand I_19854 (I340036,I340370,I340192);
nor I_19855 (I340418,I159854,I159836);
and I_19856 (I340435,I340283,I340418);
nor I_19857 (I340452,I340370,I340435);
DFFARX1 I_19858 (I340452,I2859,I340059,I340045,);
nor I_19859 (I340483,I340085,I340418);
DFFARX1 I_19860 (I340483,I2859,I340059,I340030,);
nor I_19861 (I340514,I340362,I340418);
not I_19862 (I340531,I340514);
nand I_19863 (I340039,I340531,I340387);
not I_19864 (I340586,I2866);
DFFARX1 I_19865 (I48419,I2859,I340586,I340612,);
not I_19866 (I340620,I340612);
nand I_19867 (I340637,I48395,I48404);
and I_19868 (I340654,I340637,I48398);
DFFARX1 I_19869 (I340654,I2859,I340586,I340680,);
DFFARX1 I_19870 (I340680,I2859,I340586,I340575,);
DFFARX1 I_19871 (I48416,I2859,I340586,I340711,);
nand I_19872 (I340719,I340711,I48407);
not I_19873 (I340736,I340719);
DFFARX1 I_19874 (I340736,I2859,I340586,I340762,);
not I_19875 (I340770,I340762);
nor I_19876 (I340578,I340620,I340770);
DFFARX1 I_19877 (I48401,I2859,I340586,I340810,);
nor I_19878 (I340569,I340810,I340680);
nor I_19879 (I340560,I340810,I340736);
nand I_19880 (I340846,I48413,I48410);
and I_19881 (I340863,I340846,I48398);
DFFARX1 I_19882 (I340863,I2859,I340586,I340889,);
not I_19883 (I340897,I340889);
nand I_19884 (I340914,I340897,I340810);
nand I_19885 (I340563,I340897,I340719);
nor I_19886 (I340945,I48395,I48410);
and I_19887 (I340962,I340810,I340945);
nor I_19888 (I340979,I340897,I340962);
DFFARX1 I_19889 (I340979,I2859,I340586,I340572,);
nor I_19890 (I341010,I340612,I340945);
DFFARX1 I_19891 (I341010,I2859,I340586,I340557,);
nor I_19892 (I341041,I340889,I340945);
not I_19893 (I341058,I341041);
nand I_19894 (I340566,I341058,I340914);
not I_19895 (I341113,I2866);
DFFARX1 I_19896 (I491688,I2859,I341113,I341139,);
not I_19897 (I341147,I341139);
nand I_19898 (I341164,I491670,I491670);
and I_19899 (I341181,I341164,I491676);
DFFARX1 I_19900 (I341181,I2859,I341113,I341207,);
DFFARX1 I_19901 (I341207,I2859,I341113,I341102,);
DFFARX1 I_19902 (I491673,I2859,I341113,I341238,);
nand I_19903 (I341246,I341238,I491682);
not I_19904 (I341263,I341246);
DFFARX1 I_19905 (I341263,I2859,I341113,I341289,);
not I_19906 (I341297,I341289);
nor I_19907 (I341105,I341147,I341297);
DFFARX1 I_19908 (I491694,I2859,I341113,I341337,);
nor I_19909 (I341096,I341337,I341207);
nor I_19910 (I341087,I341337,I341263);
nand I_19911 (I341373,I491685,I491679);
and I_19912 (I341390,I341373,I491673);
DFFARX1 I_19913 (I341390,I2859,I341113,I341416,);
not I_19914 (I341424,I341416);
nand I_19915 (I341441,I341424,I341337);
nand I_19916 (I341090,I341424,I341246);
nor I_19917 (I341472,I491691,I491679);
and I_19918 (I341489,I341337,I341472);
nor I_19919 (I341506,I341424,I341489);
DFFARX1 I_19920 (I341506,I2859,I341113,I341099,);
nor I_19921 (I341537,I341139,I341472);
DFFARX1 I_19922 (I341537,I2859,I341113,I341084,);
nor I_19923 (I341568,I341416,I341472);
not I_19924 (I341585,I341568);
nand I_19925 (I341093,I341585,I341441);
not I_19926 (I341640,I2866);
DFFARX1 I_19927 (I513510,I2859,I341640,I341666,);
not I_19928 (I341674,I341666);
nand I_19929 (I341691,I513516,I513498);
and I_19930 (I341708,I341691,I513507);
DFFARX1 I_19931 (I341708,I2859,I341640,I341734,);
DFFARX1 I_19932 (I341734,I2859,I341640,I341629,);
DFFARX1 I_19933 (I513513,I2859,I341640,I341765,);
nand I_19934 (I341773,I341765,I513501);
not I_19935 (I341790,I341773);
DFFARX1 I_19936 (I341790,I2859,I341640,I341816,);
not I_19937 (I341824,I341816);
nor I_19938 (I341632,I341674,I341824);
DFFARX1 I_19939 (I513519,I2859,I341640,I341864,);
nor I_19940 (I341623,I341864,I341734);
nor I_19941 (I341614,I341864,I341790);
nand I_19942 (I341900,I513498,I513504);
and I_19943 (I341917,I341900,I513522);
DFFARX1 I_19944 (I341917,I2859,I341640,I341943,);
not I_19945 (I341951,I341943);
nand I_19946 (I341968,I341951,I341864);
nand I_19947 (I341617,I341951,I341773);
nor I_19948 (I341999,I513501,I513504);
and I_19949 (I342016,I341864,I341999);
nor I_19950 (I342033,I341951,I342016);
DFFARX1 I_19951 (I342033,I2859,I341640,I341626,);
nor I_19952 (I342064,I341666,I341999);
DFFARX1 I_19953 (I342064,I2859,I341640,I341611,);
nor I_19954 (I342095,I341943,I341999);
not I_19955 (I342112,I342095);
nand I_19956 (I341620,I342112,I341968);
not I_19957 (I342167,I2866);
DFFARX1 I_19958 (I223229,I2859,I342167,I342193,);
not I_19959 (I342201,I342193);
nand I_19960 (I342218,I223247,I223238);
and I_19961 (I342235,I342218,I223241);
DFFARX1 I_19962 (I342235,I2859,I342167,I342261,);
DFFARX1 I_19963 (I342261,I2859,I342167,I342156,);
DFFARX1 I_19964 (I223235,I2859,I342167,I342292,);
nand I_19965 (I342300,I342292,I223226);
not I_19966 (I342317,I342300);
DFFARX1 I_19967 (I342317,I2859,I342167,I342343,);
not I_19968 (I342351,I342343);
nor I_19969 (I342159,I342201,I342351);
DFFARX1 I_19970 (I223232,I2859,I342167,I342391,);
nor I_19971 (I342150,I342391,I342261);
nor I_19972 (I342141,I342391,I342317);
nand I_19973 (I342427,I223226,I223223);
and I_19974 (I342444,I342427,I223244);
DFFARX1 I_19975 (I342444,I2859,I342167,I342470,);
not I_19976 (I342478,I342470);
nand I_19977 (I342495,I342478,I342391);
nand I_19978 (I342144,I342478,I342300);
nor I_19979 (I342526,I223223,I223223);
and I_19980 (I342543,I342391,I342526);
nor I_19981 (I342560,I342478,I342543);
DFFARX1 I_19982 (I342560,I2859,I342167,I342153,);
nor I_19983 (I342591,I342193,I342526);
DFFARX1 I_19984 (I342591,I2859,I342167,I342138,);
nor I_19985 (I342622,I342470,I342526);
not I_19986 (I342639,I342622);
nand I_19987 (I342147,I342639,I342495);
not I_19988 (I342694,I2866);
DFFARX1 I_19989 (I536692,I2859,I342694,I342720,);
not I_19990 (I342728,I342720);
nand I_19991 (I342745,I536686,I536704);
and I_19992 (I342762,I342745,I536689);
DFFARX1 I_19993 (I342762,I2859,I342694,I342788,);
DFFARX1 I_19994 (I342788,I2859,I342694,I342683,);
DFFARX1 I_19995 (I536710,I2859,I342694,I342819,);
nand I_19996 (I342827,I342819,I536695);
not I_19997 (I342844,I342827);
DFFARX1 I_19998 (I342844,I2859,I342694,I342870,);
not I_19999 (I342878,I342870);
nor I_20000 (I342686,I342728,I342878);
DFFARX1 I_20001 (I536707,I2859,I342694,I342918,);
nor I_20002 (I342677,I342918,I342788);
nor I_20003 (I342668,I342918,I342844);
nand I_20004 (I342954,I536698,I536713);
and I_20005 (I342971,I342954,I536701);
DFFARX1 I_20006 (I342971,I2859,I342694,I342997,);
not I_20007 (I343005,I342997);
nand I_20008 (I343022,I343005,I342918);
nand I_20009 (I342671,I343005,I342827);
nor I_20010 (I343053,I536686,I536713);
and I_20011 (I343070,I342918,I343053);
nor I_20012 (I343087,I343005,I343070);
DFFARX1 I_20013 (I343087,I2859,I342694,I342680,);
nor I_20014 (I343118,I342720,I343053);
DFFARX1 I_20015 (I343118,I2859,I342694,I342665,);
nor I_20016 (I343149,I342997,I343053);
not I_20017 (I343166,I343149);
nand I_20018 (I342674,I343166,I343022);
not I_20019 (I343221,I2866);
DFFARX1 I_20020 (I484174,I2859,I343221,I343247,);
not I_20021 (I343255,I343247);
nand I_20022 (I343272,I484156,I484156);
and I_20023 (I343289,I343272,I484162);
DFFARX1 I_20024 (I343289,I2859,I343221,I343315,);
DFFARX1 I_20025 (I343315,I2859,I343221,I343210,);
DFFARX1 I_20026 (I484159,I2859,I343221,I343346,);
nand I_20027 (I343354,I343346,I484168);
not I_20028 (I343371,I343354);
DFFARX1 I_20029 (I343371,I2859,I343221,I343397,);
not I_20030 (I343405,I343397);
nor I_20031 (I343213,I343255,I343405);
DFFARX1 I_20032 (I484180,I2859,I343221,I343445,);
nor I_20033 (I343204,I343445,I343315);
nor I_20034 (I343195,I343445,I343371);
nand I_20035 (I343481,I484171,I484165);
and I_20036 (I343498,I343481,I484159);
DFFARX1 I_20037 (I343498,I2859,I343221,I343524,);
not I_20038 (I343532,I343524);
nand I_20039 (I343549,I343532,I343445);
nand I_20040 (I343198,I343532,I343354);
nor I_20041 (I343580,I484177,I484165);
and I_20042 (I343597,I343445,I343580);
nor I_20043 (I343614,I343532,I343597);
DFFARX1 I_20044 (I343614,I2859,I343221,I343207,);
nor I_20045 (I343645,I343247,I343580);
DFFARX1 I_20046 (I343645,I2859,I343221,I343192,);
nor I_20047 (I343676,I343524,I343580);
not I_20048 (I343693,I343676);
nand I_20049 (I343201,I343693,I343549);
not I_20050 (I343748,I2866);
DFFARX1 I_20051 (I469724,I2859,I343748,I343774,);
not I_20052 (I343782,I343774);
nand I_20053 (I343799,I469706,I469706);
and I_20054 (I343816,I343799,I469712);
DFFARX1 I_20055 (I343816,I2859,I343748,I343842,);
DFFARX1 I_20056 (I343842,I2859,I343748,I343737,);
DFFARX1 I_20057 (I469709,I2859,I343748,I343873,);
nand I_20058 (I343881,I343873,I469718);
not I_20059 (I343898,I343881);
DFFARX1 I_20060 (I343898,I2859,I343748,I343924,);
not I_20061 (I343932,I343924);
nor I_20062 (I343740,I343782,I343932);
DFFARX1 I_20063 (I469730,I2859,I343748,I343972,);
nor I_20064 (I343731,I343972,I343842);
nor I_20065 (I343722,I343972,I343898);
nand I_20066 (I344008,I469721,I469715);
and I_20067 (I344025,I344008,I469709);
DFFARX1 I_20068 (I344025,I2859,I343748,I344051,);
not I_20069 (I344059,I344051);
nand I_20070 (I344076,I344059,I343972);
nand I_20071 (I343725,I344059,I343881);
nor I_20072 (I344107,I469727,I469715);
and I_20073 (I344124,I343972,I344107);
nor I_20074 (I344141,I344059,I344124);
DFFARX1 I_20075 (I344141,I2859,I343748,I343734,);
nor I_20076 (I344172,I343774,I344107);
DFFARX1 I_20077 (I344172,I2859,I343748,I343719,);
nor I_20078 (I344203,I344051,I344107);
not I_20079 (I344220,I344203);
nand I_20080 (I343728,I344220,I344076);
not I_20081 (I344275,I2866);
DFFARX1 I_20082 (I106612,I2859,I344275,I344301,);
not I_20083 (I344309,I344301);
nand I_20084 (I344326,I106603,I106603);
and I_20085 (I344343,I344326,I106621);
DFFARX1 I_20086 (I344343,I2859,I344275,I344369,);
DFFARX1 I_20087 (I344369,I2859,I344275,I344264,);
DFFARX1 I_20088 (I106624,I2859,I344275,I344400,);
nand I_20089 (I344408,I344400,I106606);
not I_20090 (I344425,I344408);
DFFARX1 I_20091 (I344425,I2859,I344275,I344451,);
not I_20092 (I344459,I344451);
nor I_20093 (I344267,I344309,I344459);
DFFARX1 I_20094 (I106618,I2859,I344275,I344499,);
nor I_20095 (I344258,I344499,I344369);
nor I_20096 (I344249,I344499,I344425);
nand I_20097 (I344535,I106630,I106609);
and I_20098 (I344552,I344535,I106615);
DFFARX1 I_20099 (I344552,I2859,I344275,I344578,);
not I_20100 (I344586,I344578);
nand I_20101 (I344603,I344586,I344499);
nand I_20102 (I344252,I344586,I344408);
nor I_20103 (I344634,I106627,I106609);
and I_20104 (I344651,I344499,I344634);
nor I_20105 (I344668,I344586,I344651);
DFFARX1 I_20106 (I344668,I2859,I344275,I344261,);
nor I_20107 (I344699,I344301,I344634);
DFFARX1 I_20108 (I344699,I2859,I344275,I344246,);
nor I_20109 (I344730,I344578,I344634);
not I_20110 (I344747,I344730);
nand I_20111 (I344255,I344747,I344603);
not I_20112 (I344802,I2866);
DFFARX1 I_20113 (I139286,I2859,I344802,I344828,);
not I_20114 (I344836,I344828);
nand I_20115 (I344853,I139277,I139277);
and I_20116 (I344870,I344853,I139295);
DFFARX1 I_20117 (I344870,I2859,I344802,I344896,);
DFFARX1 I_20118 (I344896,I2859,I344802,I344791,);
DFFARX1 I_20119 (I139298,I2859,I344802,I344927,);
nand I_20120 (I344935,I344927,I139280);
not I_20121 (I344952,I344935);
DFFARX1 I_20122 (I344952,I2859,I344802,I344978,);
not I_20123 (I344986,I344978);
nor I_20124 (I344794,I344836,I344986);
DFFARX1 I_20125 (I139292,I2859,I344802,I345026,);
nor I_20126 (I344785,I345026,I344896);
nor I_20127 (I344776,I345026,I344952);
nand I_20128 (I345062,I139304,I139283);
and I_20129 (I345079,I345062,I139289);
DFFARX1 I_20130 (I345079,I2859,I344802,I345105,);
not I_20131 (I345113,I345105);
nand I_20132 (I345130,I345113,I345026);
nand I_20133 (I344779,I345113,I344935);
nor I_20134 (I345161,I139301,I139283);
and I_20135 (I345178,I345026,I345161);
nor I_20136 (I345195,I345113,I345178);
DFFARX1 I_20137 (I345195,I2859,I344802,I344788,);
nor I_20138 (I345226,I344828,I345161);
DFFARX1 I_20139 (I345226,I2859,I344802,I344773,);
nor I_20140 (I345257,I345105,I345161);
not I_20141 (I345274,I345257);
nand I_20142 (I344782,I345274,I345130);
not I_20143 (I345329,I2866);
DFFARX1 I_20144 (I140340,I2859,I345329,I345355,);
not I_20145 (I345363,I345355);
nand I_20146 (I345380,I140331,I140331);
and I_20147 (I345397,I345380,I140349);
DFFARX1 I_20148 (I345397,I2859,I345329,I345423,);
DFFARX1 I_20149 (I345423,I2859,I345329,I345318,);
DFFARX1 I_20150 (I140352,I2859,I345329,I345454,);
nand I_20151 (I345462,I345454,I140334);
not I_20152 (I345479,I345462);
DFFARX1 I_20153 (I345479,I2859,I345329,I345505,);
not I_20154 (I345513,I345505);
nor I_20155 (I345321,I345363,I345513);
DFFARX1 I_20156 (I140346,I2859,I345329,I345553,);
nor I_20157 (I345312,I345553,I345423);
nor I_20158 (I345303,I345553,I345479);
nand I_20159 (I345589,I140358,I140337);
and I_20160 (I345606,I345589,I140343);
DFFARX1 I_20161 (I345606,I2859,I345329,I345632,);
not I_20162 (I345640,I345632);
nand I_20163 (I345657,I345640,I345553);
nand I_20164 (I345306,I345640,I345462);
nor I_20165 (I345688,I140355,I140337);
and I_20166 (I345705,I345553,I345688);
nor I_20167 (I345722,I345640,I345705);
DFFARX1 I_20168 (I345722,I2859,I345329,I345315,);
nor I_20169 (I345753,I345355,I345688);
DFFARX1 I_20170 (I345753,I2859,I345329,I345300,);
nor I_20171 (I345784,I345632,I345688);
not I_20172 (I345801,I345784);
nand I_20173 (I345309,I345801,I345657);
not I_20174 (I345856,I2866);
DFFARX1 I_20175 (I452384,I2859,I345856,I345882,);
not I_20176 (I345890,I345882);
nand I_20177 (I345907,I452366,I452366);
and I_20178 (I345924,I345907,I452372);
DFFARX1 I_20179 (I345924,I2859,I345856,I345950,);
DFFARX1 I_20180 (I345950,I2859,I345856,I345845,);
DFFARX1 I_20181 (I452369,I2859,I345856,I345981,);
nand I_20182 (I345989,I345981,I452378);
not I_20183 (I346006,I345989);
DFFARX1 I_20184 (I346006,I2859,I345856,I346032,);
not I_20185 (I346040,I346032);
nor I_20186 (I345848,I345890,I346040);
DFFARX1 I_20187 (I452390,I2859,I345856,I346080,);
nor I_20188 (I345839,I346080,I345950);
nor I_20189 (I345830,I346080,I346006);
nand I_20190 (I346116,I452381,I452375);
and I_20191 (I346133,I346116,I452369);
DFFARX1 I_20192 (I346133,I2859,I345856,I346159,);
not I_20193 (I346167,I346159);
nand I_20194 (I346184,I346167,I346080);
nand I_20195 (I345833,I346167,I345989);
nor I_20196 (I346215,I452387,I452375);
and I_20197 (I346232,I346080,I346215);
nor I_20198 (I346249,I346167,I346232);
DFFARX1 I_20199 (I346249,I2859,I345856,I345842,);
nor I_20200 (I346280,I345882,I346215);
DFFARX1 I_20201 (I346280,I2859,I345856,I345827,);
nor I_20202 (I346311,I346159,I346215);
not I_20203 (I346328,I346311);
nand I_20204 (I345836,I346328,I346184);
not I_20205 (I346383,I2866);
DFFARX1 I_20206 (I19419,I2859,I346383,I346409,);
not I_20207 (I346417,I346409);
nand I_20208 (I346434,I19431,I19434);
and I_20209 (I346451,I346434,I19410);
DFFARX1 I_20210 (I346451,I2859,I346383,I346477,);
DFFARX1 I_20211 (I346477,I2859,I346383,I346372,);
DFFARX1 I_20212 (I19428,I2859,I346383,I346508,);
nand I_20213 (I346516,I346508,I19416);
not I_20214 (I346533,I346516);
DFFARX1 I_20215 (I346533,I2859,I346383,I346559,);
not I_20216 (I346567,I346559);
nor I_20217 (I346375,I346417,I346567);
DFFARX1 I_20218 (I19413,I2859,I346383,I346607,);
nor I_20219 (I346366,I346607,I346477);
nor I_20220 (I346357,I346607,I346533);
nand I_20221 (I346643,I19422,I19413);
and I_20222 (I346660,I346643,I19410);
DFFARX1 I_20223 (I346660,I2859,I346383,I346686,);
not I_20224 (I346694,I346686);
nand I_20225 (I346711,I346694,I346607);
nand I_20226 (I346360,I346694,I346516);
nor I_20227 (I346742,I19425,I19413);
and I_20228 (I346759,I346607,I346742);
nor I_20229 (I346776,I346694,I346759);
DFFARX1 I_20230 (I346776,I2859,I346383,I346369,);
nor I_20231 (I346807,I346409,I346742);
DFFARX1 I_20232 (I346807,I2859,I346383,I346354,);
nor I_20233 (I346838,I346686,I346742);
not I_20234 (I346855,I346838);
nand I_20235 (I346363,I346855,I346711);
not I_20236 (I346910,I2866);
DFFARX1 I_20237 (I398360,I2859,I346910,I346936,);
not I_20238 (I346944,I346936);
nand I_20239 (I346961,I398375,I398357);
and I_20240 (I346978,I346961,I398357);
DFFARX1 I_20241 (I346978,I2859,I346910,I347004,);
DFFARX1 I_20242 (I347004,I2859,I346910,I346899,);
DFFARX1 I_20243 (I398366,I2859,I346910,I347035,);
nand I_20244 (I347043,I347035,I398384);
not I_20245 (I347060,I347043);
DFFARX1 I_20246 (I347060,I2859,I346910,I347086,);
not I_20247 (I347094,I347086);
nor I_20248 (I346902,I346944,I347094);
DFFARX1 I_20249 (I398381,I2859,I346910,I347134,);
nor I_20250 (I346893,I347134,I347004);
nor I_20251 (I346884,I347134,I347060);
nand I_20252 (I347170,I398378,I398369);
and I_20253 (I347187,I347170,I398363);
DFFARX1 I_20254 (I347187,I2859,I346910,I347213,);
not I_20255 (I347221,I347213);
nand I_20256 (I347238,I347221,I347134);
nand I_20257 (I346887,I347221,I347043);
nor I_20258 (I347269,I398372,I398369);
and I_20259 (I347286,I347134,I347269);
nor I_20260 (I347303,I347221,I347286);
DFFARX1 I_20261 (I347303,I2859,I346910,I346896,);
nor I_20262 (I347334,I346936,I347269);
DFFARX1 I_20263 (I347334,I2859,I346910,I346881,);
nor I_20264 (I347365,I347213,I347269);
not I_20265 (I347382,I347365);
nand I_20266 (I346890,I347382,I347238);
not I_20267 (I347437,I2866);
DFFARX1 I_20268 (I195553,I2859,I347437,I347463,);
not I_20269 (I347471,I347463);
nand I_20270 (I347488,I195550,I195559);
and I_20271 (I347505,I347488,I195568);
DFFARX1 I_20272 (I347505,I2859,I347437,I347531,);
DFFARX1 I_20273 (I347531,I2859,I347437,I347426,);
DFFARX1 I_20274 (I195571,I2859,I347437,I347562,);
nand I_20275 (I347570,I347562,I195574);
not I_20276 (I347587,I347570);
DFFARX1 I_20277 (I347587,I2859,I347437,I347613,);
not I_20278 (I347621,I347613);
nor I_20279 (I347429,I347471,I347621);
DFFARX1 I_20280 (I195547,I2859,I347437,I347661,);
nor I_20281 (I347420,I347661,I347531);
nor I_20282 (I347411,I347661,I347587);
nand I_20283 (I347697,I195562,I195565);
and I_20284 (I347714,I347697,I195556);
DFFARX1 I_20285 (I347714,I2859,I347437,I347740,);
not I_20286 (I347748,I347740);
nand I_20287 (I347765,I347748,I347661);
nand I_20288 (I347414,I347748,I347570);
nor I_20289 (I347796,I195547,I195565);
and I_20290 (I347813,I347661,I347796);
nor I_20291 (I347830,I347748,I347813);
DFFARX1 I_20292 (I347830,I2859,I347437,I347423,);
nor I_20293 (I347861,I347463,I347796);
DFFARX1 I_20294 (I347861,I2859,I347437,I347408,);
nor I_20295 (I347892,I347740,I347796);
not I_20296 (I347909,I347892);
nand I_20297 (I347417,I347909,I347765);
not I_20298 (I347964,I2866);
DFFARX1 I_20299 (I46838,I2859,I347964,I347990,);
not I_20300 (I347998,I347990);
nand I_20301 (I348015,I46814,I46823);
and I_20302 (I348032,I348015,I46817);
DFFARX1 I_20303 (I348032,I2859,I347964,I348058,);
DFFARX1 I_20304 (I348058,I2859,I347964,I347953,);
DFFARX1 I_20305 (I46835,I2859,I347964,I348089,);
nand I_20306 (I348097,I348089,I46826);
not I_20307 (I348114,I348097);
DFFARX1 I_20308 (I348114,I2859,I347964,I348140,);
not I_20309 (I348148,I348140);
nor I_20310 (I347956,I347998,I348148);
DFFARX1 I_20311 (I46820,I2859,I347964,I348188,);
nor I_20312 (I347947,I348188,I348058);
nor I_20313 (I347938,I348188,I348114);
nand I_20314 (I348224,I46832,I46829);
and I_20315 (I348241,I348224,I46817);
DFFARX1 I_20316 (I348241,I2859,I347964,I348267,);
not I_20317 (I348275,I348267);
nand I_20318 (I348292,I348275,I348188);
nand I_20319 (I347941,I348275,I348097);
nor I_20320 (I348323,I46814,I46829);
and I_20321 (I348340,I348188,I348323);
nor I_20322 (I348357,I348275,I348340);
DFFARX1 I_20323 (I348357,I2859,I347964,I347950,);
nor I_20324 (I348388,I347990,I348323);
DFFARX1 I_20325 (I348388,I2859,I347964,I347935,);
nor I_20326 (I348419,I348267,I348323);
not I_20327 (I348436,I348419);
nand I_20328 (I347944,I348436,I348292);
not I_20329 (I348491,I2866);
DFFARX1 I_20330 (I207521,I2859,I348491,I348517,);
not I_20331 (I348525,I348517);
nand I_20332 (I348542,I207518,I207527);
and I_20333 (I348559,I348542,I207536);
DFFARX1 I_20334 (I348559,I2859,I348491,I348585,);
DFFARX1 I_20335 (I348585,I2859,I348491,I348480,);
DFFARX1 I_20336 (I207539,I2859,I348491,I348616,);
nand I_20337 (I348624,I348616,I207542);
not I_20338 (I348641,I348624);
DFFARX1 I_20339 (I348641,I2859,I348491,I348667,);
not I_20340 (I348675,I348667);
nor I_20341 (I348483,I348525,I348675);
DFFARX1 I_20342 (I207515,I2859,I348491,I348715,);
nor I_20343 (I348474,I348715,I348585);
nor I_20344 (I348465,I348715,I348641);
nand I_20345 (I348751,I207530,I207533);
and I_20346 (I348768,I348751,I207524);
DFFARX1 I_20347 (I348768,I2859,I348491,I348794,);
not I_20348 (I348802,I348794);
nand I_20349 (I348819,I348802,I348715);
nand I_20350 (I348468,I348802,I348624);
nor I_20351 (I348850,I207515,I207533);
and I_20352 (I348867,I348715,I348850);
nor I_20353 (I348884,I348802,I348867);
DFFARX1 I_20354 (I348884,I2859,I348491,I348477,);
nor I_20355 (I348915,I348517,I348850);
DFFARX1 I_20356 (I348915,I2859,I348491,I348462,);
nor I_20357 (I348946,I348794,I348850);
not I_20358 (I348963,I348946);
nand I_20359 (I348471,I348963,I348819);
not I_20360 (I349018,I2866);
DFFARX1 I_20361 (I439914,I2859,I349018,I349044,);
not I_20362 (I349052,I349044);
nand I_20363 (I349069,I439923,I439911);
and I_20364 (I349086,I349069,I439908);
DFFARX1 I_20365 (I349086,I2859,I349018,I349112,);
DFFARX1 I_20366 (I349112,I2859,I349018,I349007,);
DFFARX1 I_20367 (I439908,I2859,I349018,I349143,);
nand I_20368 (I349151,I349143,I439905);
not I_20369 (I349168,I349151);
DFFARX1 I_20370 (I349168,I2859,I349018,I349194,);
not I_20371 (I349202,I349194);
nor I_20372 (I349010,I349052,I349202);
DFFARX1 I_20373 (I439911,I2859,I349018,I349242,);
nor I_20374 (I349001,I349242,I349112);
nor I_20375 (I348992,I349242,I349168);
nand I_20376 (I349278,I439926,I439917);
and I_20377 (I349295,I349278,I439920);
DFFARX1 I_20378 (I349295,I2859,I349018,I349321,);
not I_20379 (I349329,I349321);
nand I_20380 (I349346,I349329,I349242);
nand I_20381 (I348995,I349329,I349151);
nor I_20382 (I349377,I439905,I439917);
and I_20383 (I349394,I349242,I349377);
nor I_20384 (I349411,I349329,I349394);
DFFARX1 I_20385 (I349411,I2859,I349018,I349004,);
nor I_20386 (I349442,I349044,I349377);
DFFARX1 I_20387 (I349442,I2859,I349018,I348989,);
nor I_20388 (I349473,I349321,I349377);
not I_20389 (I349490,I349473);
nand I_20390 (I348998,I349490,I349346);
not I_20391 (I349545,I2866);
DFFARX1 I_20392 (I441597,I2859,I349545,I349571,);
not I_20393 (I349579,I349571);
nand I_20394 (I349596,I441606,I441594);
and I_20395 (I349613,I349596,I441591);
DFFARX1 I_20396 (I349613,I2859,I349545,I349639,);
DFFARX1 I_20397 (I349639,I2859,I349545,I349534,);
DFFARX1 I_20398 (I441591,I2859,I349545,I349670,);
nand I_20399 (I349678,I349670,I441588);
not I_20400 (I349695,I349678);
DFFARX1 I_20401 (I349695,I2859,I349545,I349721,);
not I_20402 (I349729,I349721);
nor I_20403 (I349537,I349579,I349729);
DFFARX1 I_20404 (I441594,I2859,I349545,I349769,);
nor I_20405 (I349528,I349769,I349639);
nor I_20406 (I349519,I349769,I349695);
nand I_20407 (I349805,I441609,I441600);
and I_20408 (I349822,I349805,I441603);
DFFARX1 I_20409 (I349822,I2859,I349545,I349848,);
not I_20410 (I349856,I349848);
nand I_20411 (I349873,I349856,I349769);
nand I_20412 (I349522,I349856,I349678);
nor I_20413 (I349904,I441588,I441600);
and I_20414 (I349921,I349769,I349904);
nor I_20415 (I349938,I349856,I349921);
DFFARX1 I_20416 (I349938,I2859,I349545,I349531,);
nor I_20417 (I349969,I349571,I349904);
DFFARX1 I_20418 (I349969,I2859,I349545,I349516,);
nor I_20419 (I350000,I349848,I349904);
not I_20420 (I350017,I350000);
nand I_20421 (I349525,I350017,I349873);
not I_20422 (I350072,I2866);
DFFARX1 I_20423 (I204257,I2859,I350072,I350098,);
not I_20424 (I350106,I350098);
nand I_20425 (I350123,I204254,I204263);
and I_20426 (I350140,I350123,I204272);
DFFARX1 I_20427 (I350140,I2859,I350072,I350166,);
DFFARX1 I_20428 (I350166,I2859,I350072,I350061,);
DFFARX1 I_20429 (I204275,I2859,I350072,I350197,);
nand I_20430 (I350205,I350197,I204278);
not I_20431 (I350222,I350205);
DFFARX1 I_20432 (I350222,I2859,I350072,I350248,);
not I_20433 (I350256,I350248);
nor I_20434 (I350064,I350106,I350256);
DFFARX1 I_20435 (I204251,I2859,I350072,I350296,);
nor I_20436 (I350055,I350296,I350166);
nor I_20437 (I350046,I350296,I350222);
nand I_20438 (I350332,I204266,I204269);
and I_20439 (I350349,I350332,I204260);
DFFARX1 I_20440 (I350349,I2859,I350072,I350375,);
not I_20441 (I350383,I350375);
nand I_20442 (I350400,I350383,I350296);
nand I_20443 (I350049,I350383,I350205);
nor I_20444 (I350431,I204251,I204269);
and I_20445 (I350448,I350296,I350431);
nor I_20446 (I350465,I350383,I350448);
DFFARX1 I_20447 (I350465,I2859,I350072,I350058,);
nor I_20448 (I350496,I350098,I350431);
DFFARX1 I_20449 (I350496,I2859,I350072,I350043,);
nor I_20450 (I350527,I350375,I350431);
not I_20451 (I350544,I350527);
nand I_20452 (I350052,I350544,I350400);
not I_20453 (I350599,I2866);
DFFARX1 I_20454 (I107139,I2859,I350599,I350625,);
not I_20455 (I350633,I350625);
nand I_20456 (I350650,I107130,I107130);
and I_20457 (I350667,I350650,I107148);
DFFARX1 I_20458 (I350667,I2859,I350599,I350693,);
DFFARX1 I_20459 (I350693,I2859,I350599,I350588,);
DFFARX1 I_20460 (I107151,I2859,I350599,I350724,);
nand I_20461 (I350732,I350724,I107133);
not I_20462 (I350749,I350732);
DFFARX1 I_20463 (I350749,I2859,I350599,I350775,);
not I_20464 (I350783,I350775);
nor I_20465 (I350591,I350633,I350783);
DFFARX1 I_20466 (I107145,I2859,I350599,I350823,);
nor I_20467 (I350582,I350823,I350693);
nor I_20468 (I350573,I350823,I350749);
nand I_20469 (I350859,I107157,I107136);
and I_20470 (I350876,I350859,I107142);
DFFARX1 I_20471 (I350876,I2859,I350599,I350902,);
not I_20472 (I350910,I350902);
nand I_20473 (I350927,I350910,I350823);
nand I_20474 (I350576,I350910,I350732);
nor I_20475 (I350958,I107154,I107136);
and I_20476 (I350975,I350823,I350958);
nor I_20477 (I350992,I350910,I350975);
DFFARX1 I_20478 (I350992,I2859,I350599,I350585,);
nor I_20479 (I351023,I350625,I350958);
DFFARX1 I_20480 (I351023,I2859,I350599,I350570,);
nor I_20481 (I351054,I350902,I350958);
not I_20482 (I351071,I351054);
nand I_20483 (I350579,I351071,I350927);
not I_20484 (I351126,I2866);
DFFARX1 I_20485 (I569290,I2859,I351126,I351152,);
not I_20486 (I351160,I351152);
nand I_20487 (I351177,I569287,I569296);
and I_20488 (I351194,I351177,I569275);
DFFARX1 I_20489 (I351194,I2859,I351126,I351220,);
DFFARX1 I_20490 (I351220,I2859,I351126,I351115,);
DFFARX1 I_20491 (I569278,I2859,I351126,I351251,);
nand I_20492 (I351259,I351251,I569293);
not I_20493 (I351276,I351259);
DFFARX1 I_20494 (I351276,I2859,I351126,I351302,);
not I_20495 (I351310,I351302);
nor I_20496 (I351118,I351160,I351310);
DFFARX1 I_20497 (I569299,I2859,I351126,I351350,);
nor I_20498 (I351109,I351350,I351220);
nor I_20499 (I351100,I351350,I351276);
nand I_20500 (I351386,I569281,I569302);
and I_20501 (I351403,I351386,I569284);
DFFARX1 I_20502 (I351403,I2859,I351126,I351429,);
not I_20503 (I351437,I351429);
nand I_20504 (I351454,I351437,I351350);
nand I_20505 (I351103,I351437,I351259);
nor I_20506 (I351485,I569275,I569302);
and I_20507 (I351502,I351350,I351485);
nor I_20508 (I351519,I351437,I351502);
DFFARX1 I_20509 (I351519,I2859,I351126,I351112,);
nor I_20510 (I351550,I351152,I351485);
DFFARX1 I_20511 (I351550,I2859,I351126,I351097,);
nor I_20512 (I351581,I351429,I351485);
not I_20513 (I351598,I351581);
nand I_20514 (I351106,I351598,I351454);
not I_20515 (I351653,I2866);
DFFARX1 I_20516 (I241343,I2859,I351653,I351679,);
not I_20517 (I351687,I351679);
nand I_20518 (I351704,I241328,I241349);
and I_20519 (I351721,I351704,I241337);
DFFARX1 I_20520 (I351721,I2859,I351653,I351747,);
DFFARX1 I_20521 (I351747,I2859,I351653,I351642,);
DFFARX1 I_20522 (I241331,I2859,I351653,I351778,);
nand I_20523 (I351786,I351778,I241340);
not I_20524 (I351803,I351786);
DFFARX1 I_20525 (I351803,I2859,I351653,I351829,);
not I_20526 (I351837,I351829);
nor I_20527 (I351645,I351687,I351837);
DFFARX1 I_20528 (I241346,I2859,I351653,I351877,);
nor I_20529 (I351636,I351877,I351747);
nor I_20530 (I351627,I351877,I351803);
nand I_20531 (I351913,I241328,I241331);
and I_20532 (I351930,I351913,I241352);
DFFARX1 I_20533 (I351930,I2859,I351653,I351956,);
not I_20534 (I351964,I351956);
nand I_20535 (I351981,I351964,I351877);
nand I_20536 (I351630,I351964,I351786);
nor I_20537 (I352012,I241334,I241331);
and I_20538 (I352029,I351877,I352012);
nor I_20539 (I352046,I351964,I352029);
DFFARX1 I_20540 (I352046,I2859,I351653,I351639,);
nor I_20541 (I352077,I351679,I352012);
DFFARX1 I_20542 (I352077,I2859,I351653,I351624,);
nor I_20543 (I352108,I351956,I352012);
not I_20544 (I352125,I352108);
nand I_20545 (I351633,I352125,I351981);
not I_20546 (I352180,I2866);
DFFARX1 I_20547 (I401590,I2859,I352180,I352206,);
not I_20548 (I352214,I352206);
nand I_20549 (I352231,I401605,I401587);
and I_20550 (I352248,I352231,I401587);
DFFARX1 I_20551 (I352248,I2859,I352180,I352274,);
DFFARX1 I_20552 (I352274,I2859,I352180,I352169,);
DFFARX1 I_20553 (I401596,I2859,I352180,I352305,);
nand I_20554 (I352313,I352305,I401614);
not I_20555 (I352330,I352313);
DFFARX1 I_20556 (I352330,I2859,I352180,I352356,);
not I_20557 (I352364,I352356);
nor I_20558 (I352172,I352214,I352364);
DFFARX1 I_20559 (I401611,I2859,I352180,I352404,);
nor I_20560 (I352163,I352404,I352274);
nor I_20561 (I352154,I352404,I352330);
nand I_20562 (I352440,I401608,I401599);
and I_20563 (I352457,I352440,I401593);
DFFARX1 I_20564 (I352457,I2859,I352180,I352483,);
not I_20565 (I352491,I352483);
nand I_20566 (I352508,I352491,I352404);
nand I_20567 (I352157,I352491,I352313);
nor I_20568 (I352539,I401602,I401599);
and I_20569 (I352556,I352404,I352539);
nor I_20570 (I352573,I352491,I352556);
DFFARX1 I_20571 (I352573,I2859,I352180,I352166,);
nor I_20572 (I352604,I352206,I352539);
DFFARX1 I_20573 (I352604,I2859,I352180,I352151,);
nor I_20574 (I352635,I352483,I352539);
not I_20575 (I352652,I352635);
nand I_20576 (I352160,I352652,I352508);
not I_20577 (I352707,I2866);
DFFARX1 I_20578 (I546680,I2859,I352707,I352733,);
not I_20579 (I352741,I352733);
nand I_20580 (I352758,I546677,I546686);
and I_20581 (I352775,I352758,I546665);
DFFARX1 I_20582 (I352775,I2859,I352707,I352801,);
DFFARX1 I_20583 (I352801,I2859,I352707,I352696,);
DFFARX1 I_20584 (I546668,I2859,I352707,I352832,);
nand I_20585 (I352840,I352832,I546683);
not I_20586 (I352857,I352840);
DFFARX1 I_20587 (I352857,I2859,I352707,I352883,);
not I_20588 (I352891,I352883);
nor I_20589 (I352699,I352741,I352891);
DFFARX1 I_20590 (I546689,I2859,I352707,I352931,);
nor I_20591 (I352690,I352931,I352801);
nor I_20592 (I352681,I352931,I352857);
nand I_20593 (I352967,I546671,I546692);
and I_20594 (I352984,I352967,I546674);
DFFARX1 I_20595 (I352984,I2859,I352707,I353010,);
not I_20596 (I353018,I353010);
nand I_20597 (I353035,I353018,I352931);
nand I_20598 (I352684,I353018,I352840);
nor I_20599 (I353066,I546665,I546692);
and I_20600 (I353083,I352931,I353066);
nor I_20601 (I353100,I353018,I353083);
DFFARX1 I_20602 (I353100,I2859,I352707,I352693,);
nor I_20603 (I353131,I352733,I353066);
DFFARX1 I_20604 (I353131,I2859,I352707,I352678,);
nor I_20605 (I353162,I353010,I353066);
not I_20606 (I353179,I353162);
nand I_20607 (I352687,I353179,I353035);
not I_20608 (I353234,I2866);
DFFARX1 I_20609 (I34717,I2859,I353234,I353260,);
not I_20610 (I353268,I353260);
nand I_20611 (I353285,I34693,I34702);
and I_20612 (I353302,I353285,I34696);
DFFARX1 I_20613 (I353302,I2859,I353234,I353328,);
DFFARX1 I_20614 (I353328,I2859,I353234,I353223,);
DFFARX1 I_20615 (I34714,I2859,I353234,I353359,);
nand I_20616 (I353367,I353359,I34705);
not I_20617 (I353384,I353367);
DFFARX1 I_20618 (I353384,I2859,I353234,I353410,);
not I_20619 (I353418,I353410);
nor I_20620 (I353226,I353268,I353418);
DFFARX1 I_20621 (I34699,I2859,I353234,I353458,);
nor I_20622 (I353217,I353458,I353328);
nor I_20623 (I353208,I353458,I353384);
nand I_20624 (I353494,I34711,I34708);
and I_20625 (I353511,I353494,I34696);
DFFARX1 I_20626 (I353511,I2859,I353234,I353537,);
not I_20627 (I353545,I353537);
nand I_20628 (I353562,I353545,I353458);
nand I_20629 (I353211,I353545,I353367);
nor I_20630 (I353593,I34693,I34708);
and I_20631 (I353610,I353458,I353593);
nor I_20632 (I353627,I353545,I353610);
DFFARX1 I_20633 (I353627,I2859,I353234,I353220,);
nor I_20634 (I353658,I353260,I353593);
DFFARX1 I_20635 (I353658,I2859,I353234,I353205,);
nor I_20636 (I353689,I353537,I353593);
not I_20637 (I353706,I353689);
nand I_20638 (I353214,I353706,I353562);
not I_20639 (I353761,I2866);
DFFARX1 I_20640 (I37352,I2859,I353761,I353787,);
not I_20641 (I353795,I353787);
nand I_20642 (I353812,I37328,I37337);
and I_20643 (I353829,I353812,I37331);
DFFARX1 I_20644 (I353829,I2859,I353761,I353855,);
DFFARX1 I_20645 (I353855,I2859,I353761,I353750,);
DFFARX1 I_20646 (I37349,I2859,I353761,I353886,);
nand I_20647 (I353894,I353886,I37340);
not I_20648 (I353911,I353894);
DFFARX1 I_20649 (I353911,I2859,I353761,I353937,);
not I_20650 (I353945,I353937);
nor I_20651 (I353753,I353795,I353945);
DFFARX1 I_20652 (I37334,I2859,I353761,I353985,);
nor I_20653 (I353744,I353985,I353855);
nor I_20654 (I353735,I353985,I353911);
nand I_20655 (I354021,I37346,I37343);
and I_20656 (I354038,I354021,I37331);
DFFARX1 I_20657 (I354038,I2859,I353761,I354064,);
not I_20658 (I354072,I354064);
nand I_20659 (I354089,I354072,I353985);
nand I_20660 (I353738,I354072,I353894);
nor I_20661 (I354120,I37328,I37343);
and I_20662 (I354137,I353985,I354120);
nor I_20663 (I354154,I354072,I354137);
DFFARX1 I_20664 (I354154,I2859,I353761,I353747,);
nor I_20665 (I354185,I353787,I354120);
DFFARX1 I_20666 (I354185,I2859,I353761,I353732,);
nor I_20667 (I354216,I354064,I354120);
not I_20668 (I354233,I354216);
nand I_20669 (I353741,I354233,I354089);
not I_20670 (I354288,I2866);
DFFARX1 I_20671 (I22069,I2859,I354288,I354314,);
not I_20672 (I354322,I354314);
nand I_20673 (I354339,I22045,I22054);
and I_20674 (I354356,I354339,I22048);
DFFARX1 I_20675 (I354356,I2859,I354288,I354382,);
DFFARX1 I_20676 (I354382,I2859,I354288,I354277,);
DFFARX1 I_20677 (I22066,I2859,I354288,I354413,);
nand I_20678 (I354421,I354413,I22057);
not I_20679 (I354438,I354421);
DFFARX1 I_20680 (I354438,I2859,I354288,I354464,);
not I_20681 (I354472,I354464);
nor I_20682 (I354280,I354322,I354472);
DFFARX1 I_20683 (I22051,I2859,I354288,I354512,);
nor I_20684 (I354271,I354512,I354382);
nor I_20685 (I354262,I354512,I354438);
nand I_20686 (I354548,I22063,I22060);
and I_20687 (I354565,I354548,I22048);
DFFARX1 I_20688 (I354565,I2859,I354288,I354591,);
not I_20689 (I354599,I354591);
nand I_20690 (I354616,I354599,I354512);
nand I_20691 (I354265,I354599,I354421);
nor I_20692 (I354647,I22045,I22060);
and I_20693 (I354664,I354512,I354647);
nor I_20694 (I354681,I354599,I354664);
DFFARX1 I_20695 (I354681,I2859,I354288,I354274,);
nor I_20696 (I354712,I354314,I354647);
DFFARX1 I_20697 (I354712,I2859,I354288,I354259,);
nor I_20698 (I354743,I354591,I354647);
not I_20699 (I354760,I354743);
nand I_20700 (I354268,I354760,I354616);
not I_20701 (I354815,I2866);
DFFARX1 I_20702 (I24177,I2859,I354815,I354841,);
not I_20703 (I354849,I354841);
nand I_20704 (I354866,I24153,I24162);
and I_20705 (I354883,I354866,I24156);
DFFARX1 I_20706 (I354883,I2859,I354815,I354909,);
DFFARX1 I_20707 (I354909,I2859,I354815,I354804,);
DFFARX1 I_20708 (I24174,I2859,I354815,I354940,);
nand I_20709 (I354948,I354940,I24165);
not I_20710 (I354965,I354948);
DFFARX1 I_20711 (I354965,I2859,I354815,I354991,);
not I_20712 (I354999,I354991);
nor I_20713 (I354807,I354849,I354999);
DFFARX1 I_20714 (I24159,I2859,I354815,I355039,);
nor I_20715 (I354798,I355039,I354909);
nor I_20716 (I354789,I355039,I354965);
nand I_20717 (I355075,I24171,I24168);
and I_20718 (I355092,I355075,I24156);
DFFARX1 I_20719 (I355092,I2859,I354815,I355118,);
not I_20720 (I355126,I355118);
nand I_20721 (I355143,I355126,I355039);
nand I_20722 (I354792,I355126,I354948);
nor I_20723 (I355174,I24153,I24168);
and I_20724 (I355191,I355039,I355174);
nor I_20725 (I355208,I355126,I355191);
DFFARX1 I_20726 (I355208,I2859,I354815,I354801,);
nor I_20727 (I355239,I354841,I355174);
DFFARX1 I_20728 (I355239,I2859,I354815,I354786,);
nor I_20729 (I355270,I355118,I355174);
not I_20730 (I355287,I355270);
nand I_20731 (I354795,I355287,I355143);
not I_20732 (I355342,I2866);
DFFARX1 I_20733 (I258683,I2859,I355342,I355368,);
not I_20734 (I355376,I355368);
nand I_20735 (I355393,I258668,I258689);
and I_20736 (I355410,I355393,I258677);
DFFARX1 I_20737 (I355410,I2859,I355342,I355436,);
DFFARX1 I_20738 (I355436,I2859,I355342,I355331,);
DFFARX1 I_20739 (I258671,I2859,I355342,I355467,);
nand I_20740 (I355475,I355467,I258680);
not I_20741 (I355492,I355475);
DFFARX1 I_20742 (I355492,I2859,I355342,I355518,);
not I_20743 (I355526,I355518);
nor I_20744 (I355334,I355376,I355526);
DFFARX1 I_20745 (I258686,I2859,I355342,I355566,);
nor I_20746 (I355325,I355566,I355436);
nor I_20747 (I355316,I355566,I355492);
nand I_20748 (I355602,I258668,I258671);
and I_20749 (I355619,I355602,I258692);
DFFARX1 I_20750 (I355619,I2859,I355342,I355645,);
not I_20751 (I355653,I355645);
nand I_20752 (I355670,I355653,I355566);
nand I_20753 (I355319,I355653,I355475);
nor I_20754 (I355701,I258674,I258671);
and I_20755 (I355718,I355566,I355701);
nor I_20756 (I355735,I355653,I355718);
DFFARX1 I_20757 (I355735,I2859,I355342,I355328,);
nor I_20758 (I355766,I355368,I355701);
DFFARX1 I_20759 (I355766,I2859,I355342,I355313,);
nor I_20760 (I355797,I355645,I355701);
not I_20761 (I355814,I355797);
nand I_20762 (I355322,I355814,I355670);
not I_20763 (I355869,I2866);
DFFARX1 I_20764 (I326294,I2859,I355869,I355895,);
not I_20765 (I355903,I355895);
nand I_20766 (I355920,I326297,I326294);
and I_20767 (I355937,I355920,I326306);
DFFARX1 I_20768 (I355937,I2859,I355869,I355963,);
DFFARX1 I_20769 (I355963,I2859,I355869,I355858,);
DFFARX1 I_20770 (I326303,I2859,I355869,I355994,);
nand I_20771 (I356002,I355994,I326309);
not I_20772 (I356019,I356002);
DFFARX1 I_20773 (I356019,I2859,I355869,I356045,);
not I_20774 (I356053,I356045);
nor I_20775 (I355861,I355903,I356053);
DFFARX1 I_20776 (I326318,I2859,I355869,I356093,);
nor I_20777 (I355852,I356093,I355963);
nor I_20778 (I355843,I356093,I356019);
nand I_20779 (I356129,I326312,I326300);
and I_20780 (I356146,I356129,I326297);
DFFARX1 I_20781 (I356146,I2859,I355869,I356172,);
not I_20782 (I356180,I356172);
nand I_20783 (I356197,I356180,I356093);
nand I_20784 (I355846,I356180,I356002);
nor I_20785 (I356228,I326315,I326300);
and I_20786 (I356245,I356093,I356228);
nor I_20787 (I356262,I356180,I356245);
DFFARX1 I_20788 (I356262,I2859,I355869,I355855,);
nor I_20789 (I356293,I355895,I356228);
DFFARX1 I_20790 (I356293,I2859,I355869,I355840,);
nor I_20791 (I356324,I356172,I356228);
not I_20792 (I356341,I356324);
nand I_20793 (I355849,I356341,I356197);
not I_20794 (I356396,I2866);
DFFARX1 I_20795 (I193921,I2859,I356396,I356422,);
not I_20796 (I356430,I356422);
nand I_20797 (I356447,I193918,I193927);
and I_20798 (I356464,I356447,I193936);
DFFARX1 I_20799 (I356464,I2859,I356396,I356490,);
DFFARX1 I_20800 (I356490,I2859,I356396,I356385,);
DFFARX1 I_20801 (I193939,I2859,I356396,I356521,);
nand I_20802 (I356529,I356521,I193942);
not I_20803 (I356546,I356529);
DFFARX1 I_20804 (I356546,I2859,I356396,I356572,);
not I_20805 (I356580,I356572);
nor I_20806 (I356388,I356430,I356580);
DFFARX1 I_20807 (I193915,I2859,I356396,I356620,);
nor I_20808 (I356379,I356620,I356490);
nor I_20809 (I356370,I356620,I356546);
nand I_20810 (I356656,I193930,I193933);
and I_20811 (I356673,I356656,I193924);
DFFARX1 I_20812 (I356673,I2859,I356396,I356699,);
not I_20813 (I356707,I356699);
nand I_20814 (I356724,I356707,I356620);
nand I_20815 (I356373,I356707,I356529);
nor I_20816 (I356755,I193915,I193933);
and I_20817 (I356772,I356620,I356755);
nor I_20818 (I356789,I356707,I356772);
DFFARX1 I_20819 (I356789,I2859,I356396,I356382,);
nor I_20820 (I356820,I356422,I356755);
DFFARX1 I_20821 (I356820,I2859,I356396,I356367,);
nor I_20822 (I356851,I356699,I356755);
not I_20823 (I356868,I356851);
nand I_20824 (I356376,I356868,I356724);
not I_20825 (I356923,I2866);
DFFARX1 I_20826 (I313578,I2859,I356923,I356949,);
not I_20827 (I356957,I356949);
nand I_20828 (I356974,I313581,I313578);
and I_20829 (I356991,I356974,I313590);
DFFARX1 I_20830 (I356991,I2859,I356923,I357017,);
DFFARX1 I_20831 (I357017,I2859,I356923,I356912,);
DFFARX1 I_20832 (I313587,I2859,I356923,I357048,);
nand I_20833 (I357056,I357048,I313593);
not I_20834 (I357073,I357056);
DFFARX1 I_20835 (I357073,I2859,I356923,I357099,);
not I_20836 (I357107,I357099);
nor I_20837 (I356915,I356957,I357107);
DFFARX1 I_20838 (I313602,I2859,I356923,I357147,);
nor I_20839 (I356906,I357147,I357017);
nor I_20840 (I356897,I357147,I357073);
nand I_20841 (I357183,I313596,I313584);
and I_20842 (I357200,I357183,I313581);
DFFARX1 I_20843 (I357200,I2859,I356923,I357226,);
not I_20844 (I357234,I357226);
nand I_20845 (I357251,I357234,I357147);
nand I_20846 (I356900,I357234,I357056);
nor I_20847 (I357282,I313599,I313584);
and I_20848 (I357299,I357147,I357282);
nor I_20849 (I357316,I357234,I357299);
DFFARX1 I_20850 (I357316,I2859,I356923,I356909,);
nor I_20851 (I357347,I356949,I357282);
DFFARX1 I_20852 (I357347,I2859,I356923,I356894,);
nor I_20853 (I357378,I357226,I357282);
not I_20854 (I357395,I357378);
nand I_20855 (I356903,I357395,I357251);
not I_20856 (I357450,I2866);
DFFARX1 I_20857 (I502630,I2859,I357450,I357476,);
not I_20858 (I357484,I357476);
nand I_20859 (I357501,I502636,I502618);
and I_20860 (I357518,I357501,I502627);
DFFARX1 I_20861 (I357518,I2859,I357450,I357544,);
DFFARX1 I_20862 (I357544,I2859,I357450,I357439,);
DFFARX1 I_20863 (I502633,I2859,I357450,I357575,);
nand I_20864 (I357583,I357575,I502621);
not I_20865 (I357600,I357583);
DFFARX1 I_20866 (I357600,I2859,I357450,I357626,);
not I_20867 (I357634,I357626);
nor I_20868 (I357442,I357484,I357634);
DFFARX1 I_20869 (I502639,I2859,I357450,I357674,);
nor I_20870 (I357433,I357674,I357544);
nor I_20871 (I357424,I357674,I357600);
nand I_20872 (I357710,I502618,I502624);
and I_20873 (I357727,I357710,I502642);
DFFARX1 I_20874 (I357727,I2859,I357450,I357753,);
not I_20875 (I357761,I357753);
nand I_20876 (I357778,I357761,I357674);
nand I_20877 (I357427,I357761,I357583);
nor I_20878 (I357809,I502621,I502624);
and I_20879 (I357826,I357674,I357809);
nor I_20880 (I357843,I357761,I357826);
DFFARX1 I_20881 (I357843,I2859,I357450,I357436,);
nor I_20882 (I357874,I357476,I357809);
DFFARX1 I_20883 (I357874,I2859,I357450,I357421,);
nor I_20884 (I357905,I357753,I357809);
not I_20885 (I357922,I357905);
nand I_20886 (I357430,I357922,I357778);
not I_20887 (I357977,I2866);
DFFARX1 I_20888 (I181953,I2859,I357977,I358003,);
not I_20889 (I358011,I358003);
nand I_20890 (I358028,I181950,I181959);
and I_20891 (I358045,I358028,I181968);
DFFARX1 I_20892 (I358045,I2859,I357977,I358071,);
DFFARX1 I_20893 (I358071,I2859,I357977,I357966,);
DFFARX1 I_20894 (I181971,I2859,I357977,I358102,);
nand I_20895 (I358110,I358102,I181974);
not I_20896 (I358127,I358110);
DFFARX1 I_20897 (I358127,I2859,I357977,I358153,);
not I_20898 (I358161,I358153);
nor I_20899 (I357969,I358011,I358161);
DFFARX1 I_20900 (I181947,I2859,I357977,I358201,);
nor I_20901 (I357960,I358201,I358071);
nor I_20902 (I357951,I358201,I358127);
nand I_20903 (I358237,I181962,I181965);
and I_20904 (I358254,I358237,I181956);
DFFARX1 I_20905 (I358254,I2859,I357977,I358280,);
not I_20906 (I358288,I358280);
nand I_20907 (I358305,I358288,I358201);
nand I_20908 (I357954,I358288,I358110);
nor I_20909 (I358336,I181947,I181965);
and I_20910 (I358353,I358201,I358336);
nor I_20911 (I358370,I358288,I358353);
DFFARX1 I_20912 (I358370,I2859,I357977,I357963,);
nor I_20913 (I358401,I358003,I358336);
DFFARX1 I_20914 (I358401,I2859,I357977,I357948,);
nor I_20915 (I358432,I358280,I358336);
not I_20916 (I358449,I358432);
nand I_20917 (I357957,I358449,I358305);
not I_20918 (I358504,I2866);
DFFARX1 I_20919 (I276586,I2859,I358504,I358530,);
not I_20920 (I358538,I358530);
nand I_20921 (I358555,I276589,I276586);
and I_20922 (I358572,I358555,I276598);
DFFARX1 I_20923 (I358572,I2859,I358504,I358598,);
DFFARX1 I_20924 (I358598,I2859,I358504,I358493,);
DFFARX1 I_20925 (I276595,I2859,I358504,I358629,);
nand I_20926 (I358637,I358629,I276601);
not I_20927 (I358654,I358637);
DFFARX1 I_20928 (I358654,I2859,I358504,I358680,);
not I_20929 (I358688,I358680);
nor I_20930 (I358496,I358538,I358688);
DFFARX1 I_20931 (I276610,I2859,I358504,I358728,);
nor I_20932 (I358487,I358728,I358598);
nor I_20933 (I358478,I358728,I358654);
nand I_20934 (I358764,I276604,I276592);
and I_20935 (I358781,I358764,I276589);
DFFARX1 I_20936 (I358781,I2859,I358504,I358807,);
not I_20937 (I358815,I358807);
nand I_20938 (I358832,I358815,I358728);
nand I_20939 (I358481,I358815,I358637);
nor I_20940 (I358863,I276607,I276592);
and I_20941 (I358880,I358728,I358863);
nor I_20942 (I358897,I358815,I358880);
DFFARX1 I_20943 (I358897,I2859,I358504,I358490,);
nor I_20944 (I358928,I358530,I358863);
DFFARX1 I_20945 (I358928,I2859,I358504,I358475,);
nor I_20946 (I358959,I358807,I358863);
not I_20947 (I358976,I358959);
nand I_20948 (I358484,I358976,I358832);
not I_20949 (I359031,I2866);
DFFARX1 I_20950 (I382210,I2859,I359031,I359057,);
not I_20951 (I359065,I359057);
nand I_20952 (I359082,I382225,I382207);
and I_20953 (I359099,I359082,I382207);
DFFARX1 I_20954 (I359099,I2859,I359031,I359125,);
DFFARX1 I_20955 (I359125,I2859,I359031,I359020,);
DFFARX1 I_20956 (I382216,I2859,I359031,I359156,);
nand I_20957 (I359164,I359156,I382234);
not I_20958 (I359181,I359164);
DFFARX1 I_20959 (I359181,I2859,I359031,I359207,);
not I_20960 (I359215,I359207);
nor I_20961 (I359023,I359065,I359215);
DFFARX1 I_20962 (I382231,I2859,I359031,I359255,);
nor I_20963 (I359014,I359255,I359125);
nor I_20964 (I359005,I359255,I359181);
nand I_20965 (I359291,I382228,I382219);
and I_20966 (I359308,I359291,I382213);
DFFARX1 I_20967 (I359308,I2859,I359031,I359334,);
not I_20968 (I359342,I359334);
nand I_20969 (I359359,I359342,I359255);
nand I_20970 (I359008,I359342,I359164);
nor I_20971 (I359390,I382222,I382219);
and I_20972 (I359407,I359255,I359390);
nor I_20973 (I359424,I359342,I359407);
DFFARX1 I_20974 (I359424,I2859,I359031,I359017,);
nor I_20975 (I359455,I359057,I359390);
DFFARX1 I_20976 (I359455,I2859,I359031,I359002,);
nor I_20977 (I359486,I359334,I359390);
not I_20978 (I359503,I359486);
nand I_20979 (I359011,I359503,I359359);
not I_20980 (I359558,I2866);
DFFARX1 I_20981 (I532692,I2859,I359558,I359584,);
not I_20982 (I359592,I359584);
nand I_20983 (I359609,I532674,I532677);
and I_20984 (I359626,I359609,I532689);
DFFARX1 I_20985 (I359626,I2859,I359558,I359652,);
DFFARX1 I_20986 (I359652,I2859,I359558,I359547,);
DFFARX1 I_20987 (I532698,I2859,I359558,I359683,);
nand I_20988 (I359691,I359683,I532683);
not I_20989 (I359708,I359691);
DFFARX1 I_20990 (I359708,I2859,I359558,I359734,);
not I_20991 (I359742,I359734);
nor I_20992 (I359550,I359592,I359742);
DFFARX1 I_20993 (I532695,I2859,I359558,I359782,);
nor I_20994 (I359541,I359782,I359652);
nor I_20995 (I359532,I359782,I359708);
nand I_20996 (I359818,I532686,I532680);
and I_20997 (I359835,I359818,I532674);
DFFARX1 I_20998 (I359835,I2859,I359558,I359861,);
not I_20999 (I359869,I359861);
nand I_21000 (I359886,I359869,I359782);
nand I_21001 (I359535,I359869,I359691);
nor I_21002 (I359917,I532677,I532680);
and I_21003 (I359934,I359782,I359917);
nor I_21004 (I359951,I359869,I359934);
DFFARX1 I_21005 (I359951,I2859,I359558,I359544,);
nor I_21006 (I359982,I359584,I359917);
DFFARX1 I_21007 (I359982,I2859,I359558,I359529,);
nor I_21008 (I360013,I359861,I359917);
not I_21009 (I360030,I360013);
nand I_21010 (I359538,I360030,I359886);
not I_21011 (I360085,I2866);
DFFARX1 I_21012 (I179777,I2859,I360085,I360111,);
not I_21013 (I360119,I360111);
nand I_21014 (I360136,I179774,I179783);
and I_21015 (I360153,I360136,I179792);
DFFARX1 I_21016 (I360153,I2859,I360085,I360179,);
DFFARX1 I_21017 (I360179,I2859,I360085,I360074,);
DFFARX1 I_21018 (I179795,I2859,I360085,I360210,);
nand I_21019 (I360218,I360210,I179798);
not I_21020 (I360235,I360218);
DFFARX1 I_21021 (I360235,I2859,I360085,I360261,);
not I_21022 (I360269,I360261);
nor I_21023 (I360077,I360119,I360269);
DFFARX1 I_21024 (I179771,I2859,I360085,I360309,);
nor I_21025 (I360068,I360309,I360179);
nor I_21026 (I360059,I360309,I360235);
nand I_21027 (I360345,I179786,I179789);
and I_21028 (I360362,I360345,I179780);
DFFARX1 I_21029 (I360362,I2859,I360085,I360388,);
not I_21030 (I360396,I360388);
nand I_21031 (I360413,I360396,I360309);
nand I_21032 (I360062,I360396,I360218);
nor I_21033 (I360444,I179771,I179789);
and I_21034 (I360461,I360309,I360444);
nor I_21035 (I360478,I360396,I360461);
DFFARX1 I_21036 (I360478,I2859,I360085,I360071,);
nor I_21037 (I360509,I360111,I360444);
DFFARX1 I_21038 (I360509,I2859,I360085,I360056,);
nor I_21039 (I360540,I360388,I360444);
not I_21040 (I360557,I360540);
nand I_21041 (I360065,I360557,I360413);
not I_21042 (I360612,I2866);
DFFARX1 I_21043 (I421616,I2859,I360612,I360638,);
not I_21044 (I360646,I360638);
nand I_21045 (I360663,I421631,I421613);
and I_21046 (I360680,I360663,I421613);
DFFARX1 I_21047 (I360680,I2859,I360612,I360706,);
DFFARX1 I_21048 (I360706,I2859,I360612,I360601,);
DFFARX1 I_21049 (I421622,I2859,I360612,I360737,);
nand I_21050 (I360745,I360737,I421640);
not I_21051 (I360762,I360745);
DFFARX1 I_21052 (I360762,I2859,I360612,I360788,);
not I_21053 (I360796,I360788);
nor I_21054 (I360604,I360646,I360796);
DFFARX1 I_21055 (I421637,I2859,I360612,I360836,);
nor I_21056 (I360595,I360836,I360706);
nor I_21057 (I360586,I360836,I360762);
nand I_21058 (I360872,I421634,I421625);
and I_21059 (I360889,I360872,I421619);
DFFARX1 I_21060 (I360889,I2859,I360612,I360915,);
not I_21061 (I360923,I360915);
nand I_21062 (I360940,I360923,I360836);
nand I_21063 (I360589,I360923,I360745);
nor I_21064 (I360971,I421628,I421625);
and I_21065 (I360988,I360836,I360971);
nor I_21066 (I361005,I360923,I360988);
DFFARX1 I_21067 (I361005,I2859,I360612,I360598,);
nor I_21068 (I361036,I360638,I360971);
DFFARX1 I_21069 (I361036,I2859,I360612,I360583,);
nor I_21070 (I361067,I360915,I360971);
not I_21071 (I361084,I361067);
nand I_21072 (I360592,I361084,I360940);
not I_21073 (I361139,I2866);
DFFARX1 I_21074 (I12041,I2859,I361139,I361165,);
not I_21075 (I361173,I361165);
nand I_21076 (I361190,I12053,I12056);
and I_21077 (I361207,I361190,I12032);
DFFARX1 I_21078 (I361207,I2859,I361139,I361233,);
DFFARX1 I_21079 (I361233,I2859,I361139,I361128,);
DFFARX1 I_21080 (I12050,I2859,I361139,I361264,);
nand I_21081 (I361272,I361264,I12038);
not I_21082 (I361289,I361272);
DFFARX1 I_21083 (I361289,I2859,I361139,I361315,);
not I_21084 (I361323,I361315);
nor I_21085 (I361131,I361173,I361323);
DFFARX1 I_21086 (I12035,I2859,I361139,I361363,);
nor I_21087 (I361122,I361363,I361233);
nor I_21088 (I361113,I361363,I361289);
nand I_21089 (I361399,I12044,I12035);
and I_21090 (I361416,I361399,I12032);
DFFARX1 I_21091 (I361416,I2859,I361139,I361442,);
not I_21092 (I361450,I361442);
nand I_21093 (I361467,I361450,I361363);
nand I_21094 (I361116,I361450,I361272);
nor I_21095 (I361498,I12047,I12035);
and I_21096 (I361515,I361363,I361498);
nor I_21097 (I361532,I361450,I361515);
DFFARX1 I_21098 (I361532,I2859,I361139,I361125,);
nor I_21099 (I361563,I361165,I361498);
DFFARX1 I_21100 (I361563,I2859,I361139,I361110,);
nor I_21101 (I361594,I361442,I361498);
not I_21102 (I361611,I361594);
nand I_21103 (I361119,I361611,I361467);
not I_21104 (I361666,I2866);
DFFARX1 I_21105 (I227989,I2859,I361666,I361692,);
not I_21106 (I361700,I361692);
nand I_21107 (I361717,I228007,I227998);
and I_21108 (I361734,I361717,I228001);
DFFARX1 I_21109 (I361734,I2859,I361666,I361760,);
DFFARX1 I_21110 (I361760,I2859,I361666,I361655,);
DFFARX1 I_21111 (I227995,I2859,I361666,I361791,);
nand I_21112 (I361799,I361791,I227986);
not I_21113 (I361816,I361799);
DFFARX1 I_21114 (I361816,I2859,I361666,I361842,);
not I_21115 (I361850,I361842);
nor I_21116 (I361658,I361700,I361850);
DFFARX1 I_21117 (I227992,I2859,I361666,I361890,);
nor I_21118 (I361649,I361890,I361760);
nor I_21119 (I361640,I361890,I361816);
nand I_21120 (I361926,I227986,I227983);
and I_21121 (I361943,I361926,I228004);
DFFARX1 I_21122 (I361943,I2859,I361666,I361969,);
not I_21123 (I361977,I361969);
nand I_21124 (I361994,I361977,I361890);
nand I_21125 (I361643,I361977,I361799);
nor I_21126 (I362025,I227983,I227983);
and I_21127 (I362042,I361890,I362025);
nor I_21128 (I362059,I361977,I362042);
DFFARX1 I_21129 (I362059,I2859,I361666,I361652,);
nor I_21130 (I362090,I361692,I362025);
DFFARX1 I_21131 (I362090,I2859,I361666,I361637,);
nor I_21132 (I362121,I361969,I362025);
not I_21133 (I362138,I362121);
nand I_21134 (I361646,I362138,I361994);
not I_21135 (I362193,I2866);
DFFARX1 I_21136 (I453540,I2859,I362193,I362219,);
not I_21137 (I362227,I362219);
nand I_21138 (I362244,I453522,I453522);
and I_21139 (I362261,I362244,I453528);
DFFARX1 I_21140 (I362261,I2859,I362193,I362287,);
DFFARX1 I_21141 (I362287,I2859,I362193,I362182,);
DFFARX1 I_21142 (I453525,I2859,I362193,I362318,);
nand I_21143 (I362326,I362318,I453534);
not I_21144 (I362343,I362326);
DFFARX1 I_21145 (I362343,I2859,I362193,I362369,);
not I_21146 (I362377,I362369);
nor I_21147 (I362185,I362227,I362377);
DFFARX1 I_21148 (I453546,I2859,I362193,I362417,);
nor I_21149 (I362176,I362417,I362287);
nor I_21150 (I362167,I362417,I362343);
nand I_21151 (I362453,I453537,I453531);
and I_21152 (I362470,I362453,I453525);
DFFARX1 I_21153 (I362470,I2859,I362193,I362496,);
not I_21154 (I362504,I362496);
nand I_21155 (I362521,I362504,I362417);
nand I_21156 (I362170,I362504,I362326);
nor I_21157 (I362552,I453543,I453531);
and I_21158 (I362569,I362417,I362552);
nor I_21159 (I362586,I362504,I362569);
DFFARX1 I_21160 (I362586,I2859,I362193,I362179,);
nor I_21161 (I362617,I362219,I362552);
DFFARX1 I_21162 (I362617,I2859,I362193,I362164,);
nor I_21163 (I362648,I362496,I362552);
not I_21164 (I362665,I362648);
nand I_21165 (I362173,I362665,I362521);
not I_21166 (I362720,I2866);
DFFARX1 I_21167 (I103634,I2859,I362720,I362746,);
not I_21168 (I362754,I362746);
nand I_21169 (I362771,I103631,I103649);
and I_21170 (I362788,I362771,I103640);
DFFARX1 I_21171 (I362788,I2859,I362720,I362814,);
DFFARX1 I_21172 (I362814,I2859,I362720,I362709,);
DFFARX1 I_21173 (I103646,I2859,I362720,I362845,);
nand I_21174 (I362853,I362845,I103643);
not I_21175 (I362870,I362853);
DFFARX1 I_21176 (I362870,I2859,I362720,I362896,);
not I_21177 (I362904,I362896);
nor I_21178 (I362712,I362754,I362904);
DFFARX1 I_21179 (I103637,I2859,I362720,I362944,);
nor I_21180 (I362703,I362944,I362814);
nor I_21181 (I362694,I362944,I362870);
nand I_21182 (I362980,I103628,I103652);
and I_21183 (I362997,I362980,I103631);
DFFARX1 I_21184 (I362997,I2859,I362720,I363023,);
not I_21185 (I363031,I363023);
nand I_21186 (I363048,I363031,I362944);
nand I_21187 (I362697,I363031,I362853);
nor I_21188 (I363079,I103628,I103652);
and I_21189 (I363096,I362944,I363079);
nor I_21190 (I363113,I363031,I363096);
DFFARX1 I_21191 (I363113,I2859,I362720,I362706,);
nor I_21192 (I363144,I362746,I363079);
DFFARX1 I_21193 (I363144,I2859,I362720,I362691,);
nor I_21194 (I363175,I363023,I363079);
not I_21195 (I363192,I363175);
nand I_21196 (I362700,I363192,I363048);
not I_21197 (I363247,I2866);
DFFARX1 I_21198 (I198817,I2859,I363247,I363273,);
not I_21199 (I363281,I363273);
nand I_21200 (I363298,I198814,I198823);
and I_21201 (I363315,I363298,I198832);
DFFARX1 I_21202 (I363315,I2859,I363247,I363341,);
DFFARX1 I_21203 (I363341,I2859,I363247,I363236,);
DFFARX1 I_21204 (I198835,I2859,I363247,I363372,);
nand I_21205 (I363380,I363372,I198838);
not I_21206 (I363397,I363380);
DFFARX1 I_21207 (I363397,I2859,I363247,I363423,);
not I_21208 (I363431,I363423);
nor I_21209 (I363239,I363281,I363431);
DFFARX1 I_21210 (I198811,I2859,I363247,I363471,);
nor I_21211 (I363230,I363471,I363341);
nor I_21212 (I363221,I363471,I363397);
nand I_21213 (I363507,I198826,I198829);
and I_21214 (I363524,I363507,I198820);
DFFARX1 I_21215 (I363524,I2859,I363247,I363550,);
not I_21216 (I363558,I363550);
nand I_21217 (I363575,I363558,I363471);
nand I_21218 (I363224,I363558,I363380);
nor I_21219 (I363606,I198811,I198829);
and I_21220 (I363623,I363471,I363606);
nor I_21221 (I363640,I363558,I363623);
DFFARX1 I_21222 (I363640,I2859,I363247,I363233,);
nor I_21223 (I363671,I363273,I363606);
DFFARX1 I_21224 (I363671,I2859,I363247,I363218,);
nor I_21225 (I363702,I363550,I363606);
not I_21226 (I363719,I363702);
nand I_21227 (I363227,I363719,I363575);
not I_21228 (I363774,I2866);
DFFARX1 I_21229 (I166177,I2859,I363774,I363800,);
not I_21230 (I363808,I363800);
nand I_21231 (I363825,I166174,I166183);
and I_21232 (I363842,I363825,I166192);
DFFARX1 I_21233 (I363842,I2859,I363774,I363868,);
DFFARX1 I_21234 (I363868,I2859,I363774,I363763,);
DFFARX1 I_21235 (I166195,I2859,I363774,I363899,);
nand I_21236 (I363907,I363899,I166198);
not I_21237 (I363924,I363907);
DFFARX1 I_21238 (I363924,I2859,I363774,I363950,);
not I_21239 (I363958,I363950);
nor I_21240 (I363766,I363808,I363958);
DFFARX1 I_21241 (I166171,I2859,I363774,I363998,);
nor I_21242 (I363757,I363998,I363868);
nor I_21243 (I363748,I363998,I363924);
nand I_21244 (I364034,I166186,I166189);
and I_21245 (I364051,I364034,I166180);
DFFARX1 I_21246 (I364051,I2859,I363774,I364077,);
not I_21247 (I364085,I364077);
nand I_21248 (I364102,I364085,I363998);
nand I_21249 (I363751,I364085,I363907);
nor I_21250 (I364133,I166171,I166189);
and I_21251 (I364150,I363998,I364133);
nor I_21252 (I364167,I364085,I364150);
DFFARX1 I_21253 (I364167,I2859,I363774,I363760,);
nor I_21254 (I364198,I363800,I364133);
DFFARX1 I_21255 (I364198,I2859,I363774,I363745,);
nor I_21256 (I364229,I364077,I364133);
not I_21257 (I364246,I364229);
nand I_21258 (I363754,I364246,I364102);
not I_21259 (I364301,I2866);
DFFARX1 I_21260 (I1692,I2859,I364301,I364327,);
not I_21261 (I364335,I364327);
nand I_21262 (I364352,I2852,I1708);
and I_21263 (I364369,I364352,I1876);
DFFARX1 I_21264 (I364369,I2859,I364301,I364395,);
DFFARX1 I_21265 (I364395,I2859,I364301,I364290,);
DFFARX1 I_21266 (I2812,I2859,I364301,I364426,);
nand I_21267 (I364434,I364426,I2756);
not I_21268 (I364451,I364434);
DFFARX1 I_21269 (I364451,I2859,I364301,I364477,);
not I_21270 (I364485,I364477);
nor I_21271 (I364293,I364335,I364485);
DFFARX1 I_21272 (I1420,I2859,I364301,I364525,);
nor I_21273 (I364284,I364525,I364395);
nor I_21274 (I364275,I364525,I364451);
nand I_21275 (I364561,I1956,I2532);
and I_21276 (I364578,I364561,I1452);
DFFARX1 I_21277 (I364578,I2859,I364301,I364604,);
not I_21278 (I364612,I364604);
nand I_21279 (I364629,I364612,I364525);
nand I_21280 (I364278,I364612,I364434);
nor I_21281 (I364660,I1428,I2532);
and I_21282 (I364677,I364525,I364660);
nor I_21283 (I364694,I364612,I364677);
DFFARX1 I_21284 (I364694,I2859,I364301,I364287,);
nor I_21285 (I364725,I364327,I364660);
DFFARX1 I_21286 (I364725,I2859,I364301,I364272,);
nor I_21287 (I364756,I364604,I364660);
not I_21288 (I364773,I364756);
nand I_21289 (I364281,I364773,I364629);
not I_21290 (I364828,I2866);
DFFARX1 I_21291 (I528068,I2859,I364828,I364854,);
not I_21292 (I364862,I364854);
nand I_21293 (I364879,I528050,I528053);
and I_21294 (I364896,I364879,I528065);
DFFARX1 I_21295 (I364896,I2859,I364828,I364922,);
DFFARX1 I_21296 (I364922,I2859,I364828,I364817,);
DFFARX1 I_21297 (I528074,I2859,I364828,I364953,);
nand I_21298 (I364961,I364953,I528059);
not I_21299 (I364978,I364961);
DFFARX1 I_21300 (I364978,I2859,I364828,I365004,);
not I_21301 (I365012,I365004);
nor I_21302 (I364820,I364862,I365012);
DFFARX1 I_21303 (I528071,I2859,I364828,I365052,);
nor I_21304 (I364811,I365052,I364922);
nor I_21305 (I364802,I365052,I364978);
nand I_21306 (I365088,I528062,I528056);
and I_21307 (I365105,I365088,I528050);
DFFARX1 I_21308 (I365105,I2859,I364828,I365131,);
not I_21309 (I365139,I365131);
nand I_21310 (I365156,I365139,I365052);
nand I_21311 (I364805,I365139,I364961);
nor I_21312 (I365187,I528053,I528056);
and I_21313 (I365204,I365052,I365187);
nor I_21314 (I365221,I365139,I365204);
DFFARX1 I_21315 (I365221,I2859,I364828,I364814,);
nor I_21316 (I365252,I364854,I365187);
DFFARX1 I_21317 (I365252,I2859,I364828,I364799,);
nor I_21318 (I365283,I365131,I365187);
not I_21319 (I365300,I365283);
nand I_21320 (I364808,I365300,I365156);
not I_21321 (I365355,I2866);
DFFARX1 I_21322 (I64364,I2859,I365355,I365381,);
not I_21323 (I365389,I365381);
nand I_21324 (I365406,I64361,I64379);
and I_21325 (I365423,I365406,I64370);
DFFARX1 I_21326 (I365423,I2859,I365355,I365449,);
DFFARX1 I_21327 (I365449,I2859,I365355,I365344,);
DFFARX1 I_21328 (I64376,I2859,I365355,I365480,);
nand I_21329 (I365488,I365480,I64373);
not I_21330 (I365505,I365488);
DFFARX1 I_21331 (I365505,I2859,I365355,I365531,);
not I_21332 (I365539,I365531);
nor I_21333 (I365347,I365389,I365539);
DFFARX1 I_21334 (I64367,I2859,I365355,I365579,);
nor I_21335 (I365338,I365579,I365449);
nor I_21336 (I365329,I365579,I365505);
nand I_21337 (I365615,I64358,I64382);
and I_21338 (I365632,I365615,I64361);
DFFARX1 I_21339 (I365632,I2859,I365355,I365658,);
not I_21340 (I365666,I365658);
nand I_21341 (I365683,I365666,I365579);
nand I_21342 (I365332,I365666,I365488);
nor I_21343 (I365714,I64358,I64382);
and I_21344 (I365731,I365579,I365714);
nor I_21345 (I365748,I365666,I365731);
DFFARX1 I_21346 (I365748,I2859,I365355,I365341,);
nor I_21347 (I365779,I365381,I365714);
DFFARX1 I_21348 (I365779,I2859,I365355,I365326,);
nor I_21349 (I365810,I365658,I365714);
not I_21350 (I365827,I365810);
nand I_21351 (I365335,I365827,I365683);
not I_21352 (I365882,I2866);
DFFARX1 I_21353 (I413218,I2859,I365882,I365908,);
not I_21354 (I365916,I365908);
nand I_21355 (I365933,I413233,I413215);
and I_21356 (I365950,I365933,I413215);
DFFARX1 I_21357 (I365950,I2859,I365882,I365976,);
DFFARX1 I_21358 (I365976,I2859,I365882,I365871,);
DFFARX1 I_21359 (I413224,I2859,I365882,I366007,);
nand I_21360 (I366015,I366007,I413242);
not I_21361 (I366032,I366015);
DFFARX1 I_21362 (I366032,I2859,I365882,I366058,);
not I_21363 (I366066,I366058);
nor I_21364 (I365874,I365916,I366066);
DFFARX1 I_21365 (I413239,I2859,I365882,I366106,);
nor I_21366 (I365865,I366106,I365976);
nor I_21367 (I365856,I366106,I366032);
nand I_21368 (I366142,I413236,I413227);
and I_21369 (I366159,I366142,I413221);
DFFARX1 I_21370 (I366159,I2859,I365882,I366185,);
not I_21371 (I366193,I366185);
nand I_21372 (I366210,I366193,I366106);
nand I_21373 (I365859,I366193,I366015);
nor I_21374 (I366241,I413230,I413227);
and I_21375 (I366258,I366106,I366241);
nor I_21376 (I366275,I366193,I366258);
DFFARX1 I_21377 (I366275,I2859,I365882,I365868,);
nor I_21378 (I366306,I365908,I366241);
DFFARX1 I_21379 (I366306,I2859,I365882,I365853,);
nor I_21380 (I366337,I366185,I366241);
not I_21381 (I366354,I366337);
nand I_21382 (I365862,I366354,I366210);
not I_21383 (I366409,I2866);
DFFARX1 I_21384 (I331496,I2859,I366409,I366435,);
not I_21385 (I366443,I366435);
nand I_21386 (I366460,I331499,I331496);
and I_21387 (I366477,I366460,I331508);
DFFARX1 I_21388 (I366477,I2859,I366409,I366503,);
DFFARX1 I_21389 (I366503,I2859,I366409,I366398,);
DFFARX1 I_21390 (I331505,I2859,I366409,I366534,);
nand I_21391 (I366542,I366534,I331511);
not I_21392 (I366559,I366542);
DFFARX1 I_21393 (I366559,I2859,I366409,I366585,);
not I_21394 (I366593,I366585);
nor I_21395 (I366401,I366443,I366593);
DFFARX1 I_21396 (I331520,I2859,I366409,I366633,);
nor I_21397 (I366392,I366633,I366503);
nor I_21398 (I366383,I366633,I366559);
nand I_21399 (I366669,I331514,I331502);
and I_21400 (I366686,I366669,I331499);
DFFARX1 I_21401 (I366686,I2859,I366409,I366712,);
not I_21402 (I366720,I366712);
nand I_21403 (I366737,I366720,I366633);
nand I_21404 (I366386,I366720,I366542);
nor I_21405 (I366768,I331517,I331502);
and I_21406 (I366785,I366633,I366768);
nor I_21407 (I366802,I366720,I366785);
DFFARX1 I_21408 (I366802,I2859,I366409,I366395,);
nor I_21409 (I366833,I366435,I366768);
DFFARX1 I_21410 (I366833,I2859,I366409,I366380,);
nor I_21411 (I366864,I366712,I366768);
not I_21412 (I366881,I366864);
nand I_21413 (I366389,I366881,I366737);
not I_21414 (I366936,I2866);
DFFARX1 I_21415 (I555010,I2859,I366936,I366962,);
not I_21416 (I366970,I366962);
nand I_21417 (I366987,I555007,I555016);
and I_21418 (I367004,I366987,I554995);
DFFARX1 I_21419 (I367004,I2859,I366936,I367030,);
DFFARX1 I_21420 (I367030,I2859,I366936,I366925,);
DFFARX1 I_21421 (I554998,I2859,I366936,I367061,);
nand I_21422 (I367069,I367061,I555013);
not I_21423 (I367086,I367069);
DFFARX1 I_21424 (I367086,I2859,I366936,I367112,);
not I_21425 (I367120,I367112);
nor I_21426 (I366928,I366970,I367120);
DFFARX1 I_21427 (I555019,I2859,I366936,I367160,);
nor I_21428 (I366919,I367160,I367030);
nor I_21429 (I366910,I367160,I367086);
nand I_21430 (I367196,I555001,I555022);
and I_21431 (I367213,I367196,I555004);
DFFARX1 I_21432 (I367213,I2859,I366936,I367239,);
not I_21433 (I367247,I367239);
nand I_21434 (I367264,I367247,I367160);
nand I_21435 (I366913,I367247,I367069);
nor I_21436 (I367295,I554995,I555022);
and I_21437 (I367312,I367160,I367295);
nor I_21438 (I367329,I367247,I367312);
DFFARX1 I_21439 (I367329,I2859,I366936,I366922,);
nor I_21440 (I367360,I366962,I367295);
DFFARX1 I_21441 (I367360,I2859,I366936,I366907,);
nor I_21442 (I367391,I367239,I367295);
not I_21443 (I367408,I367391);
nand I_21444 (I366916,I367408,I367264);
not I_21445 (I367463,I2866);
DFFARX1 I_21446 (I37879,I2859,I367463,I367489,);
not I_21447 (I367497,I367489);
nand I_21448 (I367514,I37855,I37864);
and I_21449 (I367531,I367514,I37858);
DFFARX1 I_21450 (I367531,I2859,I367463,I367557,);
DFFARX1 I_21451 (I367557,I2859,I367463,I367452,);
DFFARX1 I_21452 (I37876,I2859,I367463,I367588,);
nand I_21453 (I367596,I367588,I37867);
not I_21454 (I367613,I367596);
DFFARX1 I_21455 (I367613,I2859,I367463,I367639,);
not I_21456 (I367647,I367639);
nor I_21457 (I367455,I367497,I367647);
DFFARX1 I_21458 (I37861,I2859,I367463,I367687,);
nor I_21459 (I367446,I367687,I367557);
nor I_21460 (I367437,I367687,I367613);
nand I_21461 (I367723,I37873,I37870);
and I_21462 (I367740,I367723,I37858);
DFFARX1 I_21463 (I367740,I2859,I367463,I367766,);
not I_21464 (I367774,I367766);
nand I_21465 (I367791,I367774,I367687);
nand I_21466 (I367440,I367774,I367596);
nor I_21467 (I367822,I37855,I37870);
and I_21468 (I367839,I367687,I367822);
nor I_21469 (I367856,I367774,I367839);
DFFARX1 I_21470 (I367856,I2859,I367463,I367449,);
nor I_21471 (I367887,I367489,I367822);
DFFARX1 I_21472 (I367887,I2859,I367463,I367434,);
nor I_21473 (I367918,I367766,I367822);
not I_21474 (I367935,I367918);
nand I_21475 (I367443,I367935,I367791);
not I_21476 (I367990,I2866);
DFFARX1 I_21477 (I538945,I2859,I367990,I368016,);
not I_21478 (I368024,I368016);
nand I_21479 (I368041,I538942,I538951);
and I_21480 (I368058,I368041,I538930);
DFFARX1 I_21481 (I368058,I2859,I367990,I368084,);
DFFARX1 I_21482 (I368084,I2859,I367990,I367979,);
DFFARX1 I_21483 (I538933,I2859,I367990,I368115,);
nand I_21484 (I368123,I368115,I538948);
not I_21485 (I368140,I368123);
DFFARX1 I_21486 (I368140,I2859,I367990,I368166,);
not I_21487 (I368174,I368166);
nor I_21488 (I367982,I368024,I368174);
DFFARX1 I_21489 (I538954,I2859,I367990,I368214,);
nor I_21490 (I367973,I368214,I368084);
nor I_21491 (I367964,I368214,I368140);
nand I_21492 (I368250,I538936,I538957);
and I_21493 (I368267,I368250,I538939);
DFFARX1 I_21494 (I368267,I2859,I367990,I368293,);
not I_21495 (I368301,I368293);
nand I_21496 (I368318,I368301,I368214);
nand I_21497 (I367967,I368301,I368123);
nor I_21498 (I368349,I538930,I538957);
and I_21499 (I368366,I368214,I368349);
nor I_21500 (I368383,I368301,I368366);
DFFARX1 I_21501 (I368383,I2859,I367990,I367976,);
nor I_21502 (I368414,I368016,I368349);
DFFARX1 I_21503 (I368414,I2859,I367990,I367961,);
nor I_21504 (I368445,I368293,I368349);
not I_21505 (I368462,I368445);
nand I_21506 (I367970,I368462,I368318);
not I_21507 (I368517,I2866);
DFFARX1 I_21508 (I160366,I2859,I368517,I368543,);
not I_21509 (I368551,I368543);
nand I_21510 (I368568,I160357,I160357);
and I_21511 (I368585,I368568,I160375);
DFFARX1 I_21512 (I368585,I2859,I368517,I368611,);
DFFARX1 I_21513 (I368611,I2859,I368517,I368506,);
DFFARX1 I_21514 (I160378,I2859,I368517,I368642,);
nand I_21515 (I368650,I368642,I160360);
not I_21516 (I368667,I368650);
DFFARX1 I_21517 (I368667,I2859,I368517,I368693,);
not I_21518 (I368701,I368693);
nor I_21519 (I368509,I368551,I368701);
DFFARX1 I_21520 (I160372,I2859,I368517,I368741,);
nor I_21521 (I368500,I368741,I368611);
nor I_21522 (I368491,I368741,I368667);
nand I_21523 (I368777,I160384,I160363);
and I_21524 (I368794,I368777,I160369);
DFFARX1 I_21525 (I368794,I2859,I368517,I368820,);
not I_21526 (I368828,I368820);
nand I_21527 (I368845,I368828,I368741);
nand I_21528 (I368494,I368828,I368650);
nor I_21529 (I368876,I160381,I160363);
and I_21530 (I368893,I368741,I368876);
nor I_21531 (I368910,I368828,I368893);
DFFARX1 I_21532 (I368910,I2859,I368517,I368503,);
nor I_21533 (I368941,I368543,I368876);
DFFARX1 I_21534 (I368941,I2859,I368517,I368488,);
nor I_21535 (I368972,I368820,I368876);
not I_21536 (I368989,I368972);
nand I_21537 (I368497,I368989,I368845);
not I_21538 (I369044,I2866);
DFFARX1 I_21539 (I473770,I2859,I369044,I369070,);
not I_21540 (I369078,I369070);
nand I_21541 (I369095,I473752,I473752);
and I_21542 (I369112,I369095,I473758);
DFFARX1 I_21543 (I369112,I2859,I369044,I369138,);
DFFARX1 I_21544 (I369138,I2859,I369044,I369033,);
DFFARX1 I_21545 (I473755,I2859,I369044,I369169,);
nand I_21546 (I369177,I369169,I473764);
not I_21547 (I369194,I369177);
DFFARX1 I_21548 (I369194,I2859,I369044,I369220,);
not I_21549 (I369228,I369220);
nor I_21550 (I369036,I369078,I369228);
DFFARX1 I_21551 (I473776,I2859,I369044,I369268,);
nor I_21552 (I369027,I369268,I369138);
nor I_21553 (I369018,I369268,I369194);
nand I_21554 (I369304,I473767,I473761);
and I_21555 (I369321,I369304,I473755);
DFFARX1 I_21556 (I369321,I2859,I369044,I369347,);
not I_21557 (I369355,I369347);
nand I_21558 (I369372,I369355,I369268);
nand I_21559 (I369021,I369355,I369177);
nor I_21560 (I369403,I473773,I473761);
and I_21561 (I369420,I369268,I369403);
nor I_21562 (I369437,I369355,I369420);
DFFARX1 I_21563 (I369437,I2859,I369044,I369030,);
nor I_21564 (I369468,I369070,I369403);
DFFARX1 I_21565 (I369468,I2859,I369044,I369015,);
nor I_21566 (I369499,I369347,I369403);
not I_21567 (I369516,I369499);
nand I_21568 (I369024,I369516,I369372);
not I_21569 (I369571,I2866);
DFFARX1 I_21570 (I139813,I2859,I369571,I369597,);
not I_21571 (I369605,I369597);
nand I_21572 (I369622,I139804,I139804);
and I_21573 (I369639,I369622,I139822);
DFFARX1 I_21574 (I369639,I2859,I369571,I369665,);
DFFARX1 I_21575 (I369665,I2859,I369571,I369560,);
DFFARX1 I_21576 (I139825,I2859,I369571,I369696,);
nand I_21577 (I369704,I369696,I139807);
not I_21578 (I369721,I369704);
DFFARX1 I_21579 (I369721,I2859,I369571,I369747,);
not I_21580 (I369755,I369747);
nor I_21581 (I369563,I369605,I369755);
DFFARX1 I_21582 (I139819,I2859,I369571,I369795,);
nor I_21583 (I369554,I369795,I369665);
nor I_21584 (I369545,I369795,I369721);
nand I_21585 (I369831,I139831,I139810);
and I_21586 (I369848,I369831,I139816);
DFFARX1 I_21587 (I369848,I2859,I369571,I369874,);
not I_21588 (I369882,I369874);
nand I_21589 (I369899,I369882,I369795);
nand I_21590 (I369548,I369882,I369704);
nor I_21591 (I369930,I139828,I139810);
and I_21592 (I369947,I369795,I369930);
nor I_21593 (I369964,I369882,I369947);
DFFARX1 I_21594 (I369964,I2859,I369571,I369557,);
nor I_21595 (I369995,I369597,I369930);
DFFARX1 I_21596 (I369995,I2859,I369571,I369542,);
nor I_21597 (I370026,I369874,I369930);
not I_21598 (I370043,I370026);
nand I_21599 (I369551,I370043,I369899);
not I_21600 (I370098,I2866);
DFFARX1 I_21601 (I97089,I2859,I370098,I370124,);
not I_21602 (I370132,I370124);
nand I_21603 (I370149,I97086,I97104);
and I_21604 (I370166,I370149,I97095);
DFFARX1 I_21605 (I370166,I2859,I370098,I370192,);
DFFARX1 I_21606 (I370192,I2859,I370098,I370087,);
DFFARX1 I_21607 (I97101,I2859,I370098,I370223,);
nand I_21608 (I370231,I370223,I97098);
not I_21609 (I370248,I370231);
DFFARX1 I_21610 (I370248,I2859,I370098,I370274,);
not I_21611 (I370282,I370274);
nor I_21612 (I370090,I370132,I370282);
DFFARX1 I_21613 (I97092,I2859,I370098,I370322,);
nor I_21614 (I370081,I370322,I370192);
nor I_21615 (I370072,I370322,I370248);
nand I_21616 (I370358,I97083,I97107);
and I_21617 (I370375,I370358,I97086);
DFFARX1 I_21618 (I370375,I2859,I370098,I370401,);
not I_21619 (I370409,I370401);
nand I_21620 (I370426,I370409,I370322);
nand I_21621 (I370075,I370409,I370231);
nor I_21622 (I370457,I97083,I97107);
and I_21623 (I370474,I370322,I370457);
nor I_21624 (I370491,I370409,I370474);
DFFARX1 I_21625 (I370491,I2859,I370098,I370084,);
nor I_21626 (I370522,I370124,I370457);
DFFARX1 I_21627 (I370522,I2859,I370098,I370069,);
nor I_21628 (I370553,I370401,I370457);
not I_21629 (I370570,I370553);
nand I_21630 (I370078,I370570,I370426);
not I_21631 (I370625,I2866);
DFFARX1 I_21632 (I196641,I2859,I370625,I370651,);
not I_21633 (I370659,I370651);
nand I_21634 (I370676,I196638,I196647);
and I_21635 (I370693,I370676,I196656);
DFFARX1 I_21636 (I370693,I2859,I370625,I370719,);
DFFARX1 I_21637 (I370719,I2859,I370625,I370614,);
DFFARX1 I_21638 (I196659,I2859,I370625,I370750,);
nand I_21639 (I370758,I370750,I196662);
not I_21640 (I370775,I370758);
DFFARX1 I_21641 (I370775,I2859,I370625,I370801,);
not I_21642 (I370809,I370801);
nor I_21643 (I370617,I370659,I370809);
DFFARX1 I_21644 (I196635,I2859,I370625,I370849,);
nor I_21645 (I370608,I370849,I370719);
nor I_21646 (I370599,I370849,I370775);
nand I_21647 (I370885,I196650,I196653);
and I_21648 (I370902,I370885,I196644);
DFFARX1 I_21649 (I370902,I2859,I370625,I370928,);
not I_21650 (I370936,I370928);
nand I_21651 (I370953,I370936,I370849);
nand I_21652 (I370602,I370936,I370758);
nor I_21653 (I370984,I196635,I196653);
and I_21654 (I371001,I370849,I370984);
nor I_21655 (I371018,I370936,I371001);
DFFARX1 I_21656 (I371018,I2859,I370625,I370611,);
nor I_21657 (I371049,I370651,I370984);
DFFARX1 I_21658 (I371049,I2859,I370625,I370596,);
nor I_21659 (I371080,I370928,I370984);
not I_21660 (I371097,I371080);
nand I_21661 (I370605,I371097,I370953);
not I_21662 (I371152,I2866);
DFFARX1 I_21663 (I527490,I2859,I371152,I371178,);
not I_21664 (I371186,I371178);
nand I_21665 (I371203,I527472,I527475);
and I_21666 (I371220,I371203,I527487);
DFFARX1 I_21667 (I371220,I2859,I371152,I371246,);
DFFARX1 I_21668 (I371246,I2859,I371152,I371141,);
DFFARX1 I_21669 (I527496,I2859,I371152,I371277,);
nand I_21670 (I371285,I371277,I527481);
not I_21671 (I371302,I371285);
DFFARX1 I_21672 (I371302,I2859,I371152,I371328,);
not I_21673 (I371336,I371328);
nor I_21674 (I371144,I371186,I371336);
DFFARX1 I_21675 (I527493,I2859,I371152,I371376,);
nor I_21676 (I371135,I371376,I371246);
nor I_21677 (I371126,I371376,I371302);
nand I_21678 (I371412,I527484,I527478);
and I_21679 (I371429,I371412,I527472);
DFFARX1 I_21680 (I371429,I2859,I371152,I371455,);
not I_21681 (I371463,I371455);
nand I_21682 (I371480,I371463,I371376);
nand I_21683 (I371129,I371463,I371285);
nor I_21684 (I371511,I527475,I527478);
and I_21685 (I371528,I371376,I371511);
nor I_21686 (I371545,I371463,I371528);
DFFARX1 I_21687 (I371545,I2859,I371152,I371138,);
nor I_21688 (I371576,I371178,I371511);
DFFARX1 I_21689 (I371576,I2859,I371152,I371123,);
nor I_21690 (I371607,I371455,I371511);
not I_21691 (I371624,I371607);
nand I_21692 (I371132,I371624,I371480);
not I_21693 (I371679,I2866);
DFFARX1 I_21694 (I138232,I2859,I371679,I371705,);
not I_21695 (I371713,I371705);
nand I_21696 (I371730,I138223,I138223);
and I_21697 (I371747,I371730,I138241);
DFFARX1 I_21698 (I371747,I2859,I371679,I371773,);
DFFARX1 I_21699 (I371773,I2859,I371679,I371668,);
DFFARX1 I_21700 (I138244,I2859,I371679,I371804,);
nand I_21701 (I371812,I371804,I138226);
not I_21702 (I371829,I371812);
DFFARX1 I_21703 (I371829,I2859,I371679,I371855,);
not I_21704 (I371863,I371855);
nor I_21705 (I371671,I371713,I371863);
DFFARX1 I_21706 (I138238,I2859,I371679,I371903,);
nor I_21707 (I371662,I371903,I371773);
nor I_21708 (I371653,I371903,I371829);
nand I_21709 (I371939,I138250,I138229);
and I_21710 (I371956,I371939,I138235);
DFFARX1 I_21711 (I371956,I2859,I371679,I371982,);
not I_21712 (I371990,I371982);
nand I_21713 (I372007,I371990,I371903);
nand I_21714 (I371656,I371990,I371812);
nor I_21715 (I372038,I138247,I138229);
and I_21716 (I372055,I371903,I372038);
nor I_21717 (I372072,I371990,I372055);
DFFARX1 I_21718 (I372072,I2859,I371679,I371665,);
nor I_21719 (I372103,I371705,I372038);
DFFARX1 I_21720 (I372103,I2859,I371679,I371650,);
nor I_21721 (I372134,I371982,I372038);
not I_21722 (I372151,I372134);
nand I_21723 (I371659,I372151,I372007);
not I_21724 (I372206,I2866);
DFFARX1 I_21725 (I329184,I2859,I372206,I372232,);
not I_21726 (I372240,I372232);
nand I_21727 (I372257,I329187,I329184);
and I_21728 (I372274,I372257,I329196);
DFFARX1 I_21729 (I372274,I2859,I372206,I372300,);
DFFARX1 I_21730 (I372300,I2859,I372206,I372195,);
DFFARX1 I_21731 (I329193,I2859,I372206,I372331,);
nand I_21732 (I372339,I372331,I329199);
not I_21733 (I372356,I372339);
DFFARX1 I_21734 (I372356,I2859,I372206,I372382,);
not I_21735 (I372390,I372382);
nor I_21736 (I372198,I372240,I372390);
DFFARX1 I_21737 (I329208,I2859,I372206,I372430,);
nor I_21738 (I372189,I372430,I372300);
nor I_21739 (I372180,I372430,I372356);
nand I_21740 (I372466,I329202,I329190);
and I_21741 (I372483,I372466,I329187);
DFFARX1 I_21742 (I372483,I2859,I372206,I372509,);
not I_21743 (I372517,I372509);
nand I_21744 (I372534,I372517,I372430);
nand I_21745 (I372183,I372517,I372339);
nor I_21746 (I372565,I329205,I329190);
and I_21747 (I372582,I372430,I372565);
nor I_21748 (I372599,I372517,I372582);
DFFARX1 I_21749 (I372599,I2859,I372206,I372192,);
nor I_21750 (I372630,I372232,I372565);
DFFARX1 I_21751 (I372630,I2859,I372206,I372177,);
nor I_21752 (I372661,I372509,I372565);
not I_21753 (I372678,I372661);
nand I_21754 (I372186,I372678,I372534);
not I_21755 (I372733,I2866);
DFFARX1 I_21756 (I124003,I2859,I372733,I372759,);
not I_21757 (I372767,I372759);
nand I_21758 (I372784,I123994,I123994);
and I_21759 (I372801,I372784,I124012);
DFFARX1 I_21760 (I372801,I2859,I372733,I372827,);
DFFARX1 I_21761 (I372827,I2859,I372733,I372722,);
DFFARX1 I_21762 (I124015,I2859,I372733,I372858,);
nand I_21763 (I372866,I372858,I123997);
not I_21764 (I372883,I372866);
DFFARX1 I_21765 (I372883,I2859,I372733,I372909,);
not I_21766 (I372917,I372909);
nor I_21767 (I372725,I372767,I372917);
DFFARX1 I_21768 (I124009,I2859,I372733,I372957,);
nor I_21769 (I372716,I372957,I372827);
nor I_21770 (I372707,I372957,I372883);
nand I_21771 (I372993,I124021,I124000);
and I_21772 (I373010,I372993,I124006);
DFFARX1 I_21773 (I373010,I2859,I372733,I373036,);
not I_21774 (I373044,I373036);
nand I_21775 (I373061,I373044,I372957);
nand I_21776 (I372710,I373044,I372866);
nor I_21777 (I373092,I124018,I124000);
and I_21778 (I373109,I372957,I373092);
nor I_21779 (I373126,I373044,I373109);
DFFARX1 I_21780 (I373126,I2859,I372733,I372719,);
nor I_21781 (I373157,I372759,I373092);
DFFARX1 I_21782 (I373157,I2859,I372733,I372704,);
nor I_21783 (I373188,I373036,I373092);
not I_21784 (I373205,I373188);
nand I_21785 (I372713,I373205,I373061);
not I_21786 (I373260,I2866);
DFFARX1 I_21787 (I397714,I2859,I373260,I373286,);
not I_21788 (I373294,I373286);
nand I_21789 (I373311,I397729,I397711);
and I_21790 (I373328,I373311,I397711);
DFFARX1 I_21791 (I373328,I2859,I373260,I373354,);
DFFARX1 I_21792 (I373354,I2859,I373260,I373249,);
DFFARX1 I_21793 (I397720,I2859,I373260,I373385,);
nand I_21794 (I373393,I373385,I397738);
not I_21795 (I373410,I373393);
DFFARX1 I_21796 (I373410,I2859,I373260,I373436,);
not I_21797 (I373444,I373436);
nor I_21798 (I373252,I373294,I373444);
DFFARX1 I_21799 (I397735,I2859,I373260,I373484,);
nor I_21800 (I373243,I373484,I373354);
nor I_21801 (I373234,I373484,I373410);
nand I_21802 (I373520,I397732,I397723);
and I_21803 (I373537,I373520,I397717);
DFFARX1 I_21804 (I373537,I2859,I373260,I373563,);
not I_21805 (I373571,I373563);
nand I_21806 (I373588,I373571,I373484);
nand I_21807 (I373237,I373571,I373393);
nor I_21808 (I373619,I397726,I397723);
and I_21809 (I373636,I373484,I373619);
nor I_21810 (I373653,I373571,I373636);
DFFARX1 I_21811 (I373653,I2859,I373260,I373246,);
nor I_21812 (I373684,I373286,I373619);
DFFARX1 I_21813 (I373684,I2859,I373260,I373231,);
nor I_21814 (I373715,I373563,I373619);
not I_21815 (I373732,I373715);
nand I_21816 (I373240,I373732,I373588);
not I_21817 (I373787,I2866);
DFFARX1 I_21818 (I317624,I2859,I373787,I373813,);
not I_21819 (I373821,I373813);
nand I_21820 (I373838,I317627,I317624);
and I_21821 (I373855,I373838,I317636);
DFFARX1 I_21822 (I373855,I2859,I373787,I373881,);
DFFARX1 I_21823 (I373881,I2859,I373787,I373776,);
DFFARX1 I_21824 (I317633,I2859,I373787,I373912,);
nand I_21825 (I373920,I373912,I317639);
not I_21826 (I373937,I373920);
DFFARX1 I_21827 (I373937,I2859,I373787,I373963,);
not I_21828 (I373971,I373963);
nor I_21829 (I373779,I373821,I373971);
DFFARX1 I_21830 (I317648,I2859,I373787,I374011,);
nor I_21831 (I373770,I374011,I373881);
nor I_21832 (I373761,I374011,I373937);
nand I_21833 (I374047,I317642,I317630);
and I_21834 (I374064,I374047,I317627);
DFFARX1 I_21835 (I374064,I2859,I373787,I374090,);
not I_21836 (I374098,I374090);
nand I_21837 (I374115,I374098,I374011);
nand I_21838 (I373764,I374098,I373920);
nor I_21839 (I374146,I317645,I317630);
and I_21840 (I374163,I374011,I374146);
nor I_21841 (I374180,I374098,I374163);
DFFARX1 I_21842 (I374180,I2859,I373787,I373773,);
nor I_21843 (I374211,I373813,I374146);
DFFARX1 I_21844 (I374211,I2859,I373787,I373758,);
nor I_21845 (I374242,I374090,I374146);
not I_21846 (I374259,I374242);
nand I_21847 (I373767,I374259,I374115);
not I_21848 (I374314,I2866);
DFFARX1 I_21849 (I126111,I2859,I374314,I374340,);
not I_21850 (I374348,I374340);
nand I_21851 (I374365,I126102,I126102);
and I_21852 (I374382,I374365,I126120);
DFFARX1 I_21853 (I374382,I2859,I374314,I374408,);
DFFARX1 I_21854 (I374408,I2859,I374314,I374303,);
DFFARX1 I_21855 (I126123,I2859,I374314,I374439,);
nand I_21856 (I374447,I374439,I126105);
not I_21857 (I374464,I374447);
DFFARX1 I_21858 (I374464,I2859,I374314,I374490,);
not I_21859 (I374498,I374490);
nor I_21860 (I374306,I374348,I374498);
DFFARX1 I_21861 (I126117,I2859,I374314,I374538,);
nor I_21862 (I374297,I374538,I374408);
nor I_21863 (I374288,I374538,I374464);
nand I_21864 (I374574,I126129,I126108);
and I_21865 (I374591,I374574,I126114);
DFFARX1 I_21866 (I374591,I2859,I374314,I374617,);
not I_21867 (I374625,I374617);
nand I_21868 (I374642,I374625,I374538);
nand I_21869 (I374291,I374625,I374447);
nor I_21870 (I374673,I126126,I126108);
and I_21871 (I374690,I374538,I374673);
nor I_21872 (I374707,I374625,I374690);
DFFARX1 I_21873 (I374707,I2859,I374314,I374300,);
nor I_21874 (I374738,I374340,I374673);
DFFARX1 I_21875 (I374738,I2859,I374314,I374285,);
nor I_21876 (I374769,I374617,I374673);
not I_21877 (I374786,I374769);
nand I_21878 (I374294,I374786,I374642);
not I_21879 (I374841,I2866);
DFFARX1 I_21880 (I66149,I2859,I374841,I374867,);
not I_21881 (I374875,I374867);
nand I_21882 (I374892,I66146,I66164);
and I_21883 (I374909,I374892,I66155);
DFFARX1 I_21884 (I374909,I2859,I374841,I374935,);
DFFARX1 I_21885 (I374935,I2859,I374841,I374830,);
DFFARX1 I_21886 (I66161,I2859,I374841,I374966,);
nand I_21887 (I374974,I374966,I66158);
not I_21888 (I374991,I374974);
DFFARX1 I_21889 (I374991,I2859,I374841,I375017,);
not I_21890 (I375025,I375017);
nor I_21891 (I374833,I374875,I375025);
DFFARX1 I_21892 (I66152,I2859,I374841,I375065,);
nor I_21893 (I374824,I375065,I374935);
nor I_21894 (I374815,I375065,I374991);
nand I_21895 (I375101,I66143,I66167);
and I_21896 (I375118,I375101,I66146);
DFFARX1 I_21897 (I375118,I2859,I374841,I375144,);
not I_21898 (I375152,I375144);
nand I_21899 (I375169,I375152,I375065);
nand I_21900 (I374818,I375152,I374974);
nor I_21901 (I375200,I66143,I66167);
and I_21902 (I375217,I375065,I375200);
nor I_21903 (I375234,I375152,I375217);
DFFARX1 I_21904 (I375234,I2859,I374841,I374827,);
nor I_21905 (I375265,I374867,I375200);
DFFARX1 I_21906 (I375265,I2859,I374841,I374812,);
nor I_21907 (I375296,I375144,I375200);
not I_21908 (I375313,I375296);
nand I_21909 (I374821,I375313,I375169);
not I_21910 (I375368,I2866);
DFFARX1 I_21911 (I129800,I2859,I375368,I375394,);
not I_21912 (I375402,I375394);
nand I_21913 (I375419,I129791,I129791);
and I_21914 (I375436,I375419,I129809);
DFFARX1 I_21915 (I375436,I2859,I375368,I375462,);
DFFARX1 I_21916 (I375462,I2859,I375368,I375357,);
DFFARX1 I_21917 (I129812,I2859,I375368,I375493,);
nand I_21918 (I375501,I375493,I129794);
not I_21919 (I375518,I375501);
DFFARX1 I_21920 (I375518,I2859,I375368,I375544,);
not I_21921 (I375552,I375544);
nor I_21922 (I375360,I375402,I375552);
DFFARX1 I_21923 (I129806,I2859,I375368,I375592,);
nor I_21924 (I375351,I375592,I375462);
nor I_21925 (I375342,I375592,I375518);
nand I_21926 (I375628,I129818,I129797);
and I_21927 (I375645,I375628,I129803);
DFFARX1 I_21928 (I375645,I2859,I375368,I375671,);
not I_21929 (I375679,I375671);
nand I_21930 (I375696,I375679,I375592);
nand I_21931 (I375345,I375679,I375501);
nor I_21932 (I375727,I129815,I129797);
and I_21933 (I375744,I375592,I375727);
nor I_21934 (I375761,I375679,I375744);
DFFARX1 I_21935 (I375761,I2859,I375368,I375354,);
nor I_21936 (I375792,I375394,I375727);
DFFARX1 I_21937 (I375792,I2859,I375368,I375339,);
nor I_21938 (I375823,I375671,I375727);
not I_21939 (I375840,I375823);
nand I_21940 (I375348,I375840,I375696);
not I_21941 (I375895,I2866);
DFFARX1 I_21942 (I183585,I2859,I375895,I375921,);
not I_21943 (I375929,I375921);
nand I_21944 (I375946,I183582,I183591);
and I_21945 (I375963,I375946,I183600);
DFFARX1 I_21946 (I375963,I2859,I375895,I375989,);
DFFARX1 I_21947 (I375989,I2859,I375895,I375884,);
DFFARX1 I_21948 (I183603,I2859,I375895,I376020,);
nand I_21949 (I376028,I376020,I183606);
not I_21950 (I376045,I376028);
DFFARX1 I_21951 (I376045,I2859,I375895,I376071,);
not I_21952 (I376079,I376071);
nor I_21953 (I375887,I375929,I376079);
DFFARX1 I_21954 (I183579,I2859,I375895,I376119,);
nor I_21955 (I375878,I376119,I375989);
nor I_21956 (I375869,I376119,I376045);
nand I_21957 (I376155,I183594,I183597);
and I_21958 (I376172,I376155,I183588);
DFFARX1 I_21959 (I376172,I2859,I375895,I376198,);
not I_21960 (I376206,I376198);
nand I_21961 (I376223,I376206,I376119);
nand I_21962 (I375872,I376206,I376028);
nor I_21963 (I376254,I183579,I183597);
and I_21964 (I376271,I376119,I376254);
nor I_21965 (I376288,I376206,I376271);
DFFARX1 I_21966 (I376288,I2859,I375895,I375881,);
nor I_21967 (I376319,I375921,I376254);
DFFARX1 I_21968 (I376319,I2859,I375895,I375866,);
nor I_21969 (I376350,I376198,I376254);
not I_21970 (I376367,I376350);
nand I_21971 (I375875,I376367,I376223);
not I_21972 (I376428,I2866);
DFFARX1 I_21973 (I275436,I2859,I376428,I376454,);
DFFARX1 I_21974 (I275430,I2859,I376428,I376471,);
not I_21975 (I376479,I376471);
not I_21976 (I376496,I275445);
nor I_21977 (I376513,I376496,I275430);
not I_21978 (I376530,I275439);
nor I_21979 (I376547,I376513,I275448);
nor I_21980 (I376564,I376471,I376547);
DFFARX1 I_21981 (I376564,I2859,I376428,I376414,);
nor I_21982 (I376595,I275448,I275430);
nand I_21983 (I376612,I376595,I275445);
DFFARX1 I_21984 (I376612,I2859,I376428,I376417,);
nor I_21985 (I376643,I376530,I275448);
nand I_21986 (I376660,I376643,I275433);
nor I_21987 (I376677,I376454,I376660);
DFFARX1 I_21988 (I376677,I2859,I376428,I376393,);
not I_21989 (I376708,I376660);
nand I_21990 (I376405,I376471,I376708);
DFFARX1 I_21991 (I376660,I2859,I376428,I376748,);
not I_21992 (I376756,I376748);
not I_21993 (I376773,I275448);
not I_21994 (I376790,I275442);
nor I_21995 (I376807,I376790,I275439);
nor I_21996 (I376420,I376756,I376807);
nor I_21997 (I376838,I376790,I275451);
and I_21998 (I376855,I376838,I275454);
or I_21999 (I376872,I376855,I275433);
DFFARX1 I_22000 (I376872,I2859,I376428,I376898,);
nor I_22001 (I376408,I376898,I376454);
not I_22002 (I376920,I376898);
and I_22003 (I376937,I376920,I376454);
nor I_22004 (I376402,I376479,I376937);
nand I_22005 (I376968,I376920,I376530);
nor I_22006 (I376396,I376790,I376968);
nand I_22007 (I376399,I376920,I376708);
nand I_22008 (I377013,I376530,I275442);
nor I_22009 (I376411,I376773,I377013);
not I_22010 (I377074,I2866);
DFFARX1 I_22011 (I266766,I2859,I377074,I377100,);
DFFARX1 I_22012 (I266760,I2859,I377074,I377117,);
not I_22013 (I377125,I377117);
not I_22014 (I377142,I266775);
nor I_22015 (I377159,I377142,I266760);
not I_22016 (I377176,I266769);
nor I_22017 (I377193,I377159,I266778);
nor I_22018 (I377210,I377117,I377193);
DFFARX1 I_22019 (I377210,I2859,I377074,I377060,);
nor I_22020 (I377241,I266778,I266760);
nand I_22021 (I377258,I377241,I266775);
DFFARX1 I_22022 (I377258,I2859,I377074,I377063,);
nor I_22023 (I377289,I377176,I266778);
nand I_22024 (I377306,I377289,I266763);
nor I_22025 (I377323,I377100,I377306);
DFFARX1 I_22026 (I377323,I2859,I377074,I377039,);
not I_22027 (I377354,I377306);
nand I_22028 (I377051,I377117,I377354);
DFFARX1 I_22029 (I377306,I2859,I377074,I377394,);
not I_22030 (I377402,I377394);
not I_22031 (I377419,I266778);
not I_22032 (I377436,I266772);
nor I_22033 (I377453,I377436,I266769);
nor I_22034 (I377066,I377402,I377453);
nor I_22035 (I377484,I377436,I266781);
and I_22036 (I377501,I377484,I266784);
or I_22037 (I377518,I377501,I266763);
DFFARX1 I_22038 (I377518,I2859,I377074,I377544,);
nor I_22039 (I377054,I377544,I377100);
not I_22040 (I377566,I377544);
and I_22041 (I377583,I377566,I377100);
nor I_22042 (I377048,I377125,I377583);
nand I_22043 (I377614,I377566,I377176);
nor I_22044 (I377042,I377436,I377614);
nand I_22045 (I377045,I377566,I377354);
nand I_22046 (I377659,I377176,I266772);
nor I_22047 (I377057,I377419,I377659);
not I_22048 (I377720,I2866);
DFFARX1 I_22049 (I108711,I2859,I377720,I377746,);
DFFARX1 I_22050 (I108717,I2859,I377720,I377763,);
not I_22051 (I377771,I377763);
not I_22052 (I377788,I108738);
nor I_22053 (I377805,I377788,I108726);
not I_22054 (I377822,I108735);
nor I_22055 (I377839,I377805,I108720);
nor I_22056 (I377856,I377763,I377839);
DFFARX1 I_22057 (I377856,I2859,I377720,I377706,);
nor I_22058 (I377887,I108720,I108726);
nand I_22059 (I377904,I377887,I108738);
DFFARX1 I_22060 (I377904,I2859,I377720,I377709,);
nor I_22061 (I377935,I377822,I108720);
nand I_22062 (I377952,I377935,I108711);
nor I_22063 (I377969,I377746,I377952);
DFFARX1 I_22064 (I377969,I2859,I377720,I377685,);
not I_22065 (I378000,I377952);
nand I_22066 (I377697,I377763,I378000);
DFFARX1 I_22067 (I377952,I2859,I377720,I378040,);
not I_22068 (I378048,I378040);
not I_22069 (I378065,I108720);
not I_22070 (I378082,I108723);
nor I_22071 (I378099,I378082,I108735);
nor I_22072 (I377712,I378048,I378099);
nor I_22073 (I378130,I378082,I108732);
and I_22074 (I378147,I378130,I108714);
or I_22075 (I378164,I378147,I108729);
DFFARX1 I_22076 (I378164,I2859,I377720,I378190,);
nor I_22077 (I377700,I378190,I377746);
not I_22078 (I378212,I378190);
and I_22079 (I378229,I378212,I377746);
nor I_22080 (I377694,I377771,I378229);
nand I_22081 (I378260,I378212,I377822);
nor I_22082 (I377688,I378082,I378260);
nand I_22083 (I377691,I378212,I378000);
nand I_22084 (I378305,I377822,I108723);
nor I_22085 (I377703,I378065,I378305);
not I_22086 (I378366,I2866);
DFFARX1 I_22087 (I126629,I2859,I378366,I378392,);
DFFARX1 I_22088 (I126635,I2859,I378366,I378409,);
not I_22089 (I378417,I378409);
not I_22090 (I378434,I126656);
nor I_22091 (I378451,I378434,I126644);
not I_22092 (I378468,I126653);
nor I_22093 (I378485,I378451,I126638);
nor I_22094 (I378502,I378409,I378485);
DFFARX1 I_22095 (I378502,I2859,I378366,I378352,);
nor I_22096 (I378533,I126638,I126644);
nand I_22097 (I378550,I378533,I126656);
DFFARX1 I_22098 (I378550,I2859,I378366,I378355,);
nor I_22099 (I378581,I378468,I126638);
nand I_22100 (I378598,I378581,I126629);
nor I_22101 (I378615,I378392,I378598);
DFFARX1 I_22102 (I378615,I2859,I378366,I378331,);
not I_22103 (I378646,I378598);
nand I_22104 (I378343,I378409,I378646);
DFFARX1 I_22105 (I378598,I2859,I378366,I378686,);
not I_22106 (I378694,I378686);
not I_22107 (I378711,I126638);
not I_22108 (I378728,I126641);
nor I_22109 (I378745,I378728,I126653);
nor I_22110 (I378358,I378694,I378745);
nor I_22111 (I378776,I378728,I126650);
and I_22112 (I378793,I378776,I126632);
or I_22113 (I378810,I378793,I126647);
DFFARX1 I_22114 (I378810,I2859,I378366,I378836,);
nor I_22115 (I378346,I378836,I378392);
not I_22116 (I378858,I378836);
and I_22117 (I378875,I378858,I378392);
nor I_22118 (I378340,I378417,I378875);
nand I_22119 (I378906,I378858,I378468);
nor I_22120 (I378334,I378728,I378906);
nand I_22121 (I378337,I378858,I378646);
nand I_22122 (I378951,I378468,I126641);
nor I_22123 (I378349,I378711,I378951);
not I_22124 (I379012,I2866);
DFFARX1 I_22125 (I253469,I2859,I379012,I379038,);
DFFARX1 I_22126 (I253481,I2859,I379012,I379055,);
not I_22127 (I379063,I379055);
not I_22128 (I379080,I253490);
nor I_22129 (I379097,I379080,I253466);
not I_22130 (I379114,I253484);
nor I_22131 (I379131,I379097,I253478);
nor I_22132 (I379148,I379055,I379131);
DFFARX1 I_22133 (I379148,I2859,I379012,I378998,);
nor I_22134 (I379179,I253478,I253466);
nand I_22135 (I379196,I379179,I253490);
DFFARX1 I_22136 (I379196,I2859,I379012,I379001,);
nor I_22137 (I379227,I379114,I253478);
nand I_22138 (I379244,I379227,I253472);
nor I_22139 (I379261,I379038,I379244);
DFFARX1 I_22140 (I379261,I2859,I379012,I378977,);
not I_22141 (I379292,I379244);
nand I_22142 (I378989,I379055,I379292);
DFFARX1 I_22143 (I379244,I2859,I379012,I379332,);
not I_22144 (I379340,I379332);
not I_22145 (I379357,I253478);
not I_22146 (I379374,I253487);
nor I_22147 (I379391,I379374,I253484);
nor I_22148 (I379004,I379340,I379391);
nor I_22149 (I379422,I379374,I253469);
and I_22150 (I379439,I379422,I253466);
or I_22151 (I379456,I379439,I253475);
DFFARX1 I_22152 (I379456,I2859,I379012,I379482,);
nor I_22153 (I378992,I379482,I379038);
not I_22154 (I379504,I379482);
and I_22155 (I379521,I379504,I379038);
nor I_22156 (I378986,I379063,I379521);
nand I_22157 (I379552,I379504,I379114);
nor I_22158 (I378980,I379374,I379552);
nand I_22159 (I378983,I379504,I379292);
nand I_22160 (I379597,I379114,I253487);
nor I_22161 (I378995,I379357,I379597);
not I_22162 (I379658,I2866);
DFFARX1 I_22163 (I466256,I2859,I379658,I379684,);
DFFARX1 I_22164 (I466238,I2859,I379658,I379701,);
not I_22165 (I379709,I379701);
not I_22166 (I379726,I466247);
nor I_22167 (I379743,I379726,I466259);
not I_22168 (I379760,I466241);
nor I_22169 (I379777,I379743,I466250);
nor I_22170 (I379794,I379701,I379777);
DFFARX1 I_22171 (I379794,I2859,I379658,I379644,);
nor I_22172 (I379825,I466250,I466259);
nand I_22173 (I379842,I379825,I466247);
DFFARX1 I_22174 (I379842,I2859,I379658,I379647,);
nor I_22175 (I379873,I379760,I466250);
nand I_22176 (I379890,I379873,I466262);
nor I_22177 (I379907,I379684,I379890);
DFFARX1 I_22178 (I379907,I2859,I379658,I379623,);
not I_22179 (I379938,I379890);
nand I_22180 (I379635,I379701,I379938);
DFFARX1 I_22181 (I379890,I2859,I379658,I379978,);
not I_22182 (I379986,I379978);
not I_22183 (I380003,I466250);
not I_22184 (I380020,I466238);
nor I_22185 (I380037,I380020,I466241);
nor I_22186 (I379650,I379986,I380037);
nor I_22187 (I380068,I380020,I466244);
and I_22188 (I380085,I380068,I466253);
or I_22189 (I380102,I380085,I466241);
DFFARX1 I_22190 (I380102,I2859,I379658,I380128,);
nor I_22191 (I379638,I380128,I379684);
not I_22192 (I380150,I380128);
and I_22193 (I380167,I380150,I379684);
nor I_22194 (I379632,I379709,I380167);
nand I_22195 (I380198,I380150,I379760);
nor I_22196 (I379626,I380020,I380198);
nand I_22197 (I379629,I380150,I379938);
nand I_22198 (I380243,I379760,I466238);
nor I_22199 (I379641,I380003,I380243);
not I_22200 (I380304,I2866);
DFFARX1 I_22201 (I94709,I2859,I380304,I380330,);
DFFARX1 I_22202 (I94721,I2859,I380304,I380347,);
not I_22203 (I380355,I380347);
not I_22204 (I380372,I94727);
nor I_22205 (I380389,I380372,I94712);
not I_22206 (I380406,I94703);
nor I_22207 (I380423,I380389,I94724);
nor I_22208 (I380440,I380347,I380423);
DFFARX1 I_22209 (I380440,I2859,I380304,I380290,);
nor I_22210 (I380471,I94724,I94712);
nand I_22211 (I380488,I380471,I94727);
DFFARX1 I_22212 (I380488,I2859,I380304,I380293,);
nor I_22213 (I380519,I380406,I94724);
nand I_22214 (I380536,I380519,I94706);
nor I_22215 (I380553,I380330,I380536);
DFFARX1 I_22216 (I380553,I2859,I380304,I380269,);
not I_22217 (I380584,I380536);
nand I_22218 (I380281,I380347,I380584);
DFFARX1 I_22219 (I380536,I2859,I380304,I380624,);
not I_22220 (I380632,I380624);
not I_22221 (I380649,I94724);
not I_22222 (I380666,I94715);
nor I_22223 (I380683,I380666,I94703);
nor I_22224 (I380296,I380632,I380683);
nor I_22225 (I380714,I380666,I94718);
and I_22226 (I380731,I380714,I94706);
or I_22227 (I380748,I380731,I94703);
DFFARX1 I_22228 (I380748,I2859,I380304,I380774,);
nor I_22229 (I380284,I380774,I380330);
not I_22230 (I380796,I380774);
and I_22231 (I380813,I380796,I380330);
nor I_22232 (I380278,I380355,I380813);
nand I_22233 (I380844,I380796,I380406);
nor I_22234 (I380272,I380666,I380844);
nand I_22235 (I380275,I380796,I380584);
nand I_22236 (I380889,I380406,I94715);
nor I_22237 (I380287,I380649,I380889);
not I_22238 (I380950,I2866);
DFFARX1 I_22239 (I337401,I2859,I380950,I380976,);
DFFARX1 I_22240 (I337398,I2859,I380950,I380993,);
not I_22241 (I381001,I380993);
not I_22242 (I381018,I337398);
nor I_22243 (I381035,I381018,I337401);
not I_22244 (I381052,I337413);
nor I_22245 (I381069,I381035,I337407);
nor I_22246 (I381086,I380993,I381069);
DFFARX1 I_22247 (I381086,I2859,I380950,I380936,);
nor I_22248 (I381117,I337407,I337401);
nand I_22249 (I381134,I381117,I337398);
DFFARX1 I_22250 (I381134,I2859,I380950,I380939,);
nor I_22251 (I381165,I381052,I337407);
nand I_22252 (I381182,I381165,I337395);
nor I_22253 (I381199,I380976,I381182);
DFFARX1 I_22254 (I381199,I2859,I380950,I380915,);
not I_22255 (I381230,I381182);
nand I_22256 (I380927,I380993,I381230);
DFFARX1 I_22257 (I381182,I2859,I380950,I381270,);
not I_22258 (I381278,I381270);
not I_22259 (I381295,I337407);
not I_22260 (I381312,I337404);
nor I_22261 (I381329,I381312,I337413);
nor I_22262 (I380942,I381278,I381329);
nor I_22263 (I381360,I381312,I337410);
and I_22264 (I381377,I381360,I337416);
or I_22265 (I381394,I381377,I337395);
DFFARX1 I_22266 (I381394,I2859,I380950,I381420,);
nor I_22267 (I380930,I381420,I380976);
not I_22268 (I381442,I381420);
and I_22269 (I381459,I381442,I380976);
nor I_22270 (I380924,I381001,I381459);
nand I_22271 (I381490,I381442,I381052);
nor I_22272 (I380918,I381312,I381490);
nand I_22273 (I380921,I381442,I381230);
nand I_22274 (I381535,I381052,I337404);
nor I_22275 (I380933,I381295,I381535);
not I_22276 (I381596,I2866);
DFFARX1 I_22277 (I135588,I2859,I381596,I381622,);
DFFARX1 I_22278 (I135594,I2859,I381596,I381639,);
not I_22279 (I381647,I381639);
not I_22280 (I381664,I135615);
nor I_22281 (I381681,I381664,I135603);
not I_22282 (I381698,I135612);
nor I_22283 (I381715,I381681,I135597);
nor I_22284 (I381732,I381639,I381715);
DFFARX1 I_22285 (I381732,I2859,I381596,I381582,);
nor I_22286 (I381763,I135597,I135603);
nand I_22287 (I381780,I381763,I135615);
DFFARX1 I_22288 (I381780,I2859,I381596,I381585,);
nor I_22289 (I381811,I381698,I135597);
nand I_22290 (I381828,I381811,I135588);
nor I_22291 (I381845,I381622,I381828);
DFFARX1 I_22292 (I381845,I2859,I381596,I381561,);
not I_22293 (I381876,I381828);
nand I_22294 (I381573,I381639,I381876);
DFFARX1 I_22295 (I381828,I2859,I381596,I381916,);
not I_22296 (I381924,I381916);
not I_22297 (I381941,I135597);
not I_22298 (I381958,I135600);
nor I_22299 (I381975,I381958,I135612);
nor I_22300 (I381588,I381924,I381975);
nor I_22301 (I382006,I381958,I135609);
and I_22302 (I382023,I382006,I135591);
or I_22303 (I382040,I382023,I135606);
DFFARX1 I_22304 (I382040,I2859,I381596,I382066,);
nor I_22305 (I381576,I382066,I381622);
not I_22306 (I382088,I382066);
and I_22307 (I382105,I382088,I381622);
nor I_22308 (I381570,I381647,I382105);
nand I_22309 (I382136,I382088,I381698);
nor I_22310 (I381564,I381958,I382136);
nand I_22311 (I381567,I382088,I381876);
nand I_22312 (I382181,I381698,I135600);
nor I_22313 (I381579,I381941,I382181);
not I_22314 (I382242,I2866);
DFFARX1 I_22315 (I318786,I2859,I382242,I382268,);
DFFARX1 I_22316 (I318780,I2859,I382242,I382285,);
not I_22317 (I382293,I382285);
not I_22318 (I382310,I318795);
nor I_22319 (I382327,I382310,I318780);
not I_22320 (I382344,I318789);
nor I_22321 (I382361,I382327,I318798);
nor I_22322 (I382378,I382285,I382361);
DFFARX1 I_22323 (I382378,I2859,I382242,I382228,);
nor I_22324 (I382409,I318798,I318780);
nand I_22325 (I382426,I382409,I318795);
DFFARX1 I_22326 (I382426,I2859,I382242,I382231,);
nor I_22327 (I382457,I382344,I318798);
nand I_22328 (I382474,I382457,I318783);
nor I_22329 (I382491,I382268,I382474);
DFFARX1 I_22330 (I382491,I2859,I382242,I382207,);
not I_22331 (I382522,I382474);
nand I_22332 (I382219,I382285,I382522);
DFFARX1 I_22333 (I382474,I2859,I382242,I382562,);
not I_22334 (I382570,I382562);
not I_22335 (I382587,I318798);
not I_22336 (I382604,I318792);
nor I_22337 (I382621,I382604,I318789);
nor I_22338 (I382234,I382570,I382621);
nor I_22339 (I382652,I382604,I318801);
and I_22340 (I382669,I382652,I318804);
or I_22341 (I382686,I382669,I318783);
DFFARX1 I_22342 (I382686,I2859,I382242,I382712,);
nor I_22343 (I382222,I382712,I382268);
not I_22344 (I382734,I382712);
and I_22345 (I382751,I382734,I382268);
nor I_22346 (I382216,I382293,I382751);
nand I_22347 (I382782,I382734,I382344);
nor I_22348 (I382210,I382604,I382782);
nand I_22349 (I382213,I382734,I382522);
nand I_22350 (I382827,I382344,I318792);
nor I_22351 (I382225,I382587,I382827);
not I_22352 (I382888,I2866);
DFFARX1 I_22353 (I181409,I2859,I382888,I382914,);
DFFARX1 I_22354 (I181406,I2859,I382888,I382931,);
not I_22355 (I382939,I382931);
not I_22356 (I382956,I181421);
nor I_22357 (I382973,I382956,I181424);
not I_22358 (I382990,I181412);
nor I_22359 (I383007,I382973,I181418);
nor I_22360 (I383024,I382931,I383007);
DFFARX1 I_22361 (I383024,I2859,I382888,I382874,);
nor I_22362 (I383055,I181418,I181424);
nand I_22363 (I383072,I383055,I181421);
DFFARX1 I_22364 (I383072,I2859,I382888,I382877,);
nor I_22365 (I383103,I382990,I181418);
nand I_22366 (I383120,I383103,I181430);
nor I_22367 (I383137,I382914,I383120);
DFFARX1 I_22368 (I383137,I2859,I382888,I382853,);
not I_22369 (I383168,I383120);
nand I_22370 (I382865,I382931,I383168);
DFFARX1 I_22371 (I383120,I2859,I382888,I383208,);
not I_22372 (I383216,I383208);
not I_22373 (I383233,I181418);
not I_22374 (I383250,I181403);
nor I_22375 (I383267,I383250,I181412);
nor I_22376 (I382880,I383216,I383267);
nor I_22377 (I383298,I383250,I181415);
and I_22378 (I383315,I383298,I181403);
or I_22379 (I383332,I383315,I181427);
DFFARX1 I_22380 (I383332,I2859,I382888,I383358,);
nor I_22381 (I382868,I383358,I382914);
not I_22382 (I383380,I383358);
and I_22383 (I383397,I383380,I382914);
nor I_22384 (I382862,I382939,I383397);
nand I_22385 (I383428,I383380,I382990);
nor I_22386 (I382856,I383250,I383428);
nand I_22387 (I382859,I383380,I383168);
nand I_22388 (I383473,I382990,I181403);
nor I_22389 (I382871,I383233,I383473);
not I_22390 (I383534,I2866);
DFFARX1 I_22391 (I321676,I2859,I383534,I383560,);
DFFARX1 I_22392 (I321670,I2859,I383534,I383577,);
not I_22393 (I383585,I383577);
not I_22394 (I383602,I321685);
nor I_22395 (I383619,I383602,I321670);
not I_22396 (I383636,I321679);
nor I_22397 (I383653,I383619,I321688);
nor I_22398 (I383670,I383577,I383653);
DFFARX1 I_22399 (I383670,I2859,I383534,I383520,);
nor I_22400 (I383701,I321688,I321670);
nand I_22401 (I383718,I383701,I321685);
DFFARX1 I_22402 (I383718,I2859,I383534,I383523,);
nor I_22403 (I383749,I383636,I321688);
nand I_22404 (I383766,I383749,I321673);
nor I_22405 (I383783,I383560,I383766);
DFFARX1 I_22406 (I383783,I2859,I383534,I383499,);
not I_22407 (I383814,I383766);
nand I_22408 (I383511,I383577,I383814);
DFFARX1 I_22409 (I383766,I2859,I383534,I383854,);
not I_22410 (I383862,I383854);
not I_22411 (I383879,I321688);
not I_22412 (I383896,I321682);
nor I_22413 (I383913,I383896,I321679);
nor I_22414 (I383526,I383862,I383913);
nor I_22415 (I383944,I383896,I321691);
and I_22416 (I383961,I383944,I321694);
or I_22417 (I383978,I383961,I321673);
DFFARX1 I_22418 (I383978,I2859,I383534,I384004,);
nor I_22419 (I383514,I384004,I383560);
not I_22420 (I384026,I384004);
and I_22421 (I384043,I384026,I383560);
nor I_22422 (I383508,I383585,I384043);
nand I_22423 (I384074,I384026,I383636);
nor I_22424 (I383502,I383896,I384074);
nand I_22425 (I383505,I384026,I383814);
nand I_22426 (I384119,I383636,I321682);
nor I_22427 (I383517,I383879,I384119);
not I_22428 (I384180,I2866);
DFFARX1 I_22429 (I234973,I2859,I384180,I384206,);
DFFARX1 I_22430 (I234985,I2859,I384180,I384223,);
not I_22431 (I384231,I384223);
not I_22432 (I384248,I234994);
nor I_22433 (I384265,I384248,I234970);
not I_22434 (I384282,I234988);
nor I_22435 (I384299,I384265,I234982);
nor I_22436 (I384316,I384223,I384299);
DFFARX1 I_22437 (I384316,I2859,I384180,I384166,);
nor I_22438 (I384347,I234982,I234970);
nand I_22439 (I384364,I384347,I234994);
DFFARX1 I_22440 (I384364,I2859,I384180,I384169,);
nor I_22441 (I384395,I384282,I234982);
nand I_22442 (I384412,I384395,I234976);
nor I_22443 (I384429,I384206,I384412);
DFFARX1 I_22444 (I384429,I2859,I384180,I384145,);
not I_22445 (I384460,I384412);
nand I_22446 (I384157,I384223,I384460);
DFFARX1 I_22447 (I384412,I2859,I384180,I384500,);
not I_22448 (I384508,I384500);
not I_22449 (I384525,I234982);
not I_22450 (I384542,I234991);
nor I_22451 (I384559,I384542,I234988);
nor I_22452 (I384172,I384508,I384559);
nor I_22453 (I384590,I384542,I234973);
and I_22454 (I384607,I384590,I234970);
or I_22455 (I384624,I384607,I234979);
DFFARX1 I_22456 (I384624,I2859,I384180,I384650,);
nor I_22457 (I384160,I384650,I384206);
not I_22458 (I384672,I384650);
and I_22459 (I384689,I384672,I384206);
nor I_22460 (I384154,I384231,I384689);
nand I_22461 (I384720,I384672,I384282);
nor I_22462 (I384148,I384542,I384720);
nand I_22463 (I384151,I384672,I384460);
nand I_22464 (I384765,I384282,I234991);
nor I_22465 (I384163,I384525,I384765);
not I_22466 (I384826,I2866);
DFFARX1 I_22467 (I332080,I2859,I384826,I384852,);
DFFARX1 I_22468 (I332074,I2859,I384826,I384869,);
not I_22469 (I384877,I384869);
not I_22470 (I384894,I332089);
nor I_22471 (I384911,I384894,I332074);
not I_22472 (I384928,I332083);
nor I_22473 (I384945,I384911,I332092);
nor I_22474 (I384962,I384869,I384945);
DFFARX1 I_22475 (I384962,I2859,I384826,I384812,);
nor I_22476 (I384993,I332092,I332074);
nand I_22477 (I385010,I384993,I332089);
DFFARX1 I_22478 (I385010,I2859,I384826,I384815,);
nor I_22479 (I385041,I384928,I332092);
nand I_22480 (I385058,I385041,I332077);
nor I_22481 (I385075,I384852,I385058);
DFFARX1 I_22482 (I385075,I2859,I384826,I384791,);
not I_22483 (I385106,I385058);
nand I_22484 (I384803,I384869,I385106);
DFFARX1 I_22485 (I385058,I2859,I384826,I385146,);
not I_22486 (I385154,I385146);
not I_22487 (I385171,I332092);
not I_22488 (I385188,I332086);
nor I_22489 (I385205,I385188,I332083);
nor I_22490 (I384818,I385154,I385205);
nor I_22491 (I385236,I385188,I332095);
and I_22492 (I385253,I385236,I332098);
or I_22493 (I385270,I385253,I332077);
DFFARX1 I_22494 (I385270,I2859,I384826,I385296,);
nor I_22495 (I384806,I385296,I384852);
not I_22496 (I385318,I385296);
and I_22497 (I385335,I385318,I384852);
nor I_22498 (I384800,I384877,I385335);
nand I_22499 (I385366,I385318,I384928);
nor I_22500 (I384794,I385188,I385366);
nand I_22501 (I384797,I385318,I385106);
nand I_22502 (I385411,I384928,I332086);
nor I_22503 (I384809,I385171,I385411);
not I_22504 (I385472,I2866);
DFFARX1 I_22505 (I348468,I2859,I385472,I385498,);
DFFARX1 I_22506 (I348465,I2859,I385472,I385515,);
not I_22507 (I385523,I385515);
not I_22508 (I385540,I348465);
nor I_22509 (I385557,I385540,I348468);
not I_22510 (I385574,I348480);
nor I_22511 (I385591,I385557,I348474);
nor I_22512 (I385608,I385515,I385591);
DFFARX1 I_22513 (I385608,I2859,I385472,I385458,);
nor I_22514 (I385639,I348474,I348468);
nand I_22515 (I385656,I385639,I348465);
DFFARX1 I_22516 (I385656,I2859,I385472,I385461,);
nor I_22517 (I385687,I385574,I348474);
nand I_22518 (I385704,I385687,I348462);
nor I_22519 (I385721,I385498,I385704);
DFFARX1 I_22520 (I385721,I2859,I385472,I385437,);
not I_22521 (I385752,I385704);
nand I_22522 (I385449,I385515,I385752);
DFFARX1 I_22523 (I385704,I2859,I385472,I385792,);
not I_22524 (I385800,I385792);
not I_22525 (I385817,I348474);
not I_22526 (I385834,I348471);
nor I_22527 (I385851,I385834,I348480);
nor I_22528 (I385464,I385800,I385851);
nor I_22529 (I385882,I385834,I348477);
and I_22530 (I385899,I385882,I348483);
or I_22531 (I385916,I385899,I348462);
DFFARX1 I_22532 (I385916,I2859,I385472,I385942,);
nor I_22533 (I385452,I385942,I385498);
not I_22534 (I385964,I385942);
and I_22535 (I385981,I385964,I385498);
nor I_22536 (I385446,I385523,I385981);
nand I_22537 (I386012,I385964,I385574);
nor I_22538 (I385440,I385834,I386012);
nand I_22539 (I385443,I385964,I385752);
nand I_22540 (I386057,I385574,I348471);
nor I_22541 (I385455,I385817,I386057);
not I_22542 (I386118,I2866);
DFFARX1 I_22543 (I451228,I2859,I386118,I386144,);
DFFARX1 I_22544 (I451210,I2859,I386118,I386161,);
not I_22545 (I386169,I386161);
not I_22546 (I386186,I451219);
nor I_22547 (I386203,I386186,I451231);
not I_22548 (I386220,I451213);
nor I_22549 (I386237,I386203,I451222);
nor I_22550 (I386254,I386161,I386237);
DFFARX1 I_22551 (I386254,I2859,I386118,I386104,);
nor I_22552 (I386285,I451222,I451231);
nand I_22553 (I386302,I386285,I451219);
DFFARX1 I_22554 (I386302,I2859,I386118,I386107,);
nor I_22555 (I386333,I386220,I451222);
nand I_22556 (I386350,I386333,I451234);
nor I_22557 (I386367,I386144,I386350);
DFFARX1 I_22558 (I386367,I2859,I386118,I386083,);
not I_22559 (I386398,I386350);
nand I_22560 (I386095,I386161,I386398);
DFFARX1 I_22561 (I386350,I2859,I386118,I386438,);
not I_22562 (I386446,I386438);
not I_22563 (I386463,I451222);
not I_22564 (I386480,I451210);
nor I_22565 (I386497,I386480,I451213);
nor I_22566 (I386110,I386446,I386497);
nor I_22567 (I386528,I386480,I451216);
and I_22568 (I386545,I386528,I451225);
or I_22569 (I386562,I386545,I451213);
DFFARX1 I_22570 (I386562,I2859,I386118,I386588,);
nor I_22571 (I386098,I386588,I386144);
not I_22572 (I386610,I386588);
and I_22573 (I386627,I386610,I386144);
nor I_22574 (I386092,I386169,I386627);
nand I_22575 (I386658,I386610,I386220);
nor I_22576 (I386086,I386480,I386658);
nand I_22577 (I386089,I386610,I386398);
nand I_22578 (I386703,I386220,I451210);
nor I_22579 (I386101,I386463,I386703);
not I_22580 (I386764,I2866);
DFFARX1 I_22581 (I71504,I2859,I386764,I386790,);
DFFARX1 I_22582 (I71516,I2859,I386764,I386807,);
not I_22583 (I386815,I386807);
not I_22584 (I386832,I71522);
nor I_22585 (I386849,I386832,I71507);
not I_22586 (I386866,I71498);
nor I_22587 (I386883,I386849,I71519);
nor I_22588 (I386900,I386807,I386883);
DFFARX1 I_22589 (I386900,I2859,I386764,I386750,);
nor I_22590 (I386931,I71519,I71507);
nand I_22591 (I386948,I386931,I71522);
DFFARX1 I_22592 (I386948,I2859,I386764,I386753,);
nor I_22593 (I386979,I386866,I71519);
nand I_22594 (I386996,I386979,I71501);
nor I_22595 (I387013,I386790,I386996);
DFFARX1 I_22596 (I387013,I2859,I386764,I386729,);
not I_22597 (I387044,I386996);
nand I_22598 (I386741,I386807,I387044);
DFFARX1 I_22599 (I386996,I2859,I386764,I387084,);
not I_22600 (I387092,I387084);
not I_22601 (I387109,I71519);
not I_22602 (I387126,I71510);
nor I_22603 (I387143,I387126,I71498);
nor I_22604 (I386756,I387092,I387143);
nor I_22605 (I387174,I387126,I71513);
and I_22606 (I387191,I387174,I71501);
or I_22607 (I387208,I387191,I71498);
DFFARX1 I_22608 (I387208,I2859,I386764,I387234,);
nor I_22609 (I386744,I387234,I386790);
not I_22610 (I387256,I387234);
and I_22611 (I387273,I387256,I386790);
nor I_22612 (I386738,I386815,I387273);
nand I_22613 (I387304,I387256,I386866);
nor I_22614 (I386732,I387126,I387304);
nand I_22615 (I386735,I387256,I387044);
nand I_22616 (I387349,I386866,I71510);
nor I_22617 (I386747,I387109,I387349);
not I_22618 (I387410,I2866);
DFFARX1 I_22619 (I72099,I2859,I387410,I387436,);
DFFARX1 I_22620 (I72111,I2859,I387410,I387453,);
not I_22621 (I387461,I387453);
not I_22622 (I387478,I72117);
nor I_22623 (I387495,I387478,I72102);
not I_22624 (I387512,I72093);
nor I_22625 (I387529,I387495,I72114);
nor I_22626 (I387546,I387453,I387529);
DFFARX1 I_22627 (I387546,I2859,I387410,I387396,);
nor I_22628 (I387577,I72114,I72102);
nand I_22629 (I387594,I387577,I72117);
DFFARX1 I_22630 (I387594,I2859,I387410,I387399,);
nor I_22631 (I387625,I387512,I72114);
nand I_22632 (I387642,I387625,I72096);
nor I_22633 (I387659,I387436,I387642);
DFFARX1 I_22634 (I387659,I2859,I387410,I387375,);
not I_22635 (I387690,I387642);
nand I_22636 (I387387,I387453,I387690);
DFFARX1 I_22637 (I387642,I2859,I387410,I387730,);
not I_22638 (I387738,I387730);
not I_22639 (I387755,I72114);
not I_22640 (I387772,I72105);
nor I_22641 (I387789,I387772,I72093);
nor I_22642 (I387402,I387738,I387789);
nor I_22643 (I387820,I387772,I72108);
and I_22644 (I387837,I387820,I72096);
or I_22645 (I387854,I387837,I72093);
DFFARX1 I_22646 (I387854,I2859,I387410,I387880,);
nor I_22647 (I387390,I387880,I387436);
not I_22648 (I387902,I387880);
and I_22649 (I387919,I387902,I387436);
nor I_22650 (I387384,I387461,I387919);
nand I_22651 (I387950,I387902,I387512);
nor I_22652 (I387378,I387772,I387950);
nand I_22653 (I387381,I387902,I387690);
nand I_22654 (I387995,I387512,I72105);
nor I_22655 (I387393,I387755,I387995);
not I_22656 (I388056,I2866);
DFFARX1 I_22657 (I351103,I2859,I388056,I388082,);
DFFARX1 I_22658 (I351100,I2859,I388056,I388099,);
not I_22659 (I388107,I388099);
not I_22660 (I388124,I351100);
nor I_22661 (I388141,I388124,I351103);
not I_22662 (I388158,I351115);
nor I_22663 (I388175,I388141,I351109);
nor I_22664 (I388192,I388099,I388175);
DFFARX1 I_22665 (I388192,I2859,I388056,I388042,);
nor I_22666 (I388223,I351109,I351103);
nand I_22667 (I388240,I388223,I351100);
DFFARX1 I_22668 (I388240,I2859,I388056,I388045,);
nor I_22669 (I388271,I388158,I351109);
nand I_22670 (I388288,I388271,I351097);
nor I_22671 (I388305,I388082,I388288);
DFFARX1 I_22672 (I388305,I2859,I388056,I388021,);
not I_22673 (I388336,I388288);
nand I_22674 (I388033,I388099,I388336);
DFFARX1 I_22675 (I388288,I2859,I388056,I388376,);
not I_22676 (I388384,I388376);
not I_22677 (I388401,I351109);
not I_22678 (I388418,I351106);
nor I_22679 (I388435,I388418,I351115);
nor I_22680 (I388048,I388384,I388435);
nor I_22681 (I388466,I388418,I351112);
and I_22682 (I388483,I388466,I351118);
or I_22683 (I388500,I388483,I351097);
DFFARX1 I_22684 (I388500,I2859,I388056,I388526,);
nor I_22685 (I388036,I388526,I388082);
not I_22686 (I388548,I388526);
and I_22687 (I388565,I388548,I388082);
nor I_22688 (I388030,I388107,I388565);
nand I_22689 (I388596,I388548,I388158);
nor I_22690 (I388024,I388418,I388596);
nand I_22691 (I388027,I388548,I388336);
nand I_22692 (I388641,I388158,I351106);
nor I_22693 (I388039,I388401,I388641);
not I_22694 (I388702,I2866);
DFFARX1 I_22695 (I248267,I2859,I388702,I388728,);
DFFARX1 I_22696 (I248279,I2859,I388702,I388745,);
not I_22697 (I388753,I388745);
not I_22698 (I388770,I248288);
nor I_22699 (I388787,I388770,I248264);
not I_22700 (I388804,I248282);
nor I_22701 (I388821,I388787,I248276);
nor I_22702 (I388838,I388745,I388821);
DFFARX1 I_22703 (I388838,I2859,I388702,I388688,);
nor I_22704 (I388869,I248276,I248264);
nand I_22705 (I388886,I388869,I248288);
DFFARX1 I_22706 (I388886,I2859,I388702,I388691,);
nor I_22707 (I388917,I388804,I248276);
nand I_22708 (I388934,I388917,I248270);
nor I_22709 (I388951,I388728,I388934);
DFFARX1 I_22710 (I388951,I2859,I388702,I388667,);
not I_22711 (I388982,I388934);
nand I_22712 (I388679,I388745,I388982);
DFFARX1 I_22713 (I388934,I2859,I388702,I389022,);
not I_22714 (I389030,I389022);
not I_22715 (I389047,I248276);
not I_22716 (I389064,I248285);
nor I_22717 (I389081,I389064,I248282);
nor I_22718 (I388694,I389030,I389081);
nor I_22719 (I389112,I389064,I248267);
and I_22720 (I389129,I389112,I248264);
or I_22721 (I389146,I389129,I248273);
DFFARX1 I_22722 (I389146,I2859,I388702,I389172,);
nor I_22723 (I388682,I389172,I388728);
not I_22724 (I389194,I389172);
and I_22725 (I389211,I389194,I388728);
nor I_22726 (I388676,I388753,I389211);
nand I_22727 (I389242,I389194,I388804);
nor I_22728 (I388670,I389064,I389242);
nand I_22729 (I388673,I389194,I388982);
nand I_22730 (I389287,I388804,I248285);
nor I_22731 (I388685,I389047,I389287);
not I_22732 (I389348,I2866);
DFFARX1 I_22733 (I266188,I2859,I389348,I389374,);
DFFARX1 I_22734 (I266182,I2859,I389348,I389391,);
not I_22735 (I389399,I389391);
not I_22736 (I389416,I266197);
nor I_22737 (I389433,I389416,I266182);
not I_22738 (I389450,I266191);
nor I_22739 (I389467,I389433,I266200);
nor I_22740 (I389484,I389391,I389467);
DFFARX1 I_22741 (I389484,I2859,I389348,I389334,);
nor I_22742 (I389515,I266200,I266182);
nand I_22743 (I389532,I389515,I266197);
DFFARX1 I_22744 (I389532,I2859,I389348,I389337,);
nor I_22745 (I389563,I389450,I266200);
nand I_22746 (I389580,I389563,I266185);
nor I_22747 (I389597,I389374,I389580);
DFFARX1 I_22748 (I389597,I2859,I389348,I389313,);
not I_22749 (I389628,I389580);
nand I_22750 (I389325,I389391,I389628);
DFFARX1 I_22751 (I389580,I2859,I389348,I389668,);
not I_22752 (I389676,I389668);
not I_22753 (I389693,I266200);
not I_22754 (I389710,I266194);
nor I_22755 (I389727,I389710,I266191);
nor I_22756 (I389340,I389676,I389727);
nor I_22757 (I389758,I389710,I266203);
and I_22758 (I389775,I389758,I266206);
or I_22759 (I389792,I389775,I266185);
DFFARX1 I_22760 (I389792,I2859,I389348,I389818,);
nor I_22761 (I389328,I389818,I389374);
not I_22762 (I389840,I389818);
and I_22763 (I389857,I389840,I389374);
nor I_22764 (I389322,I389399,I389857);
nand I_22765 (I389888,I389840,I389450);
nor I_22766 (I389316,I389710,I389888);
nand I_22767 (I389319,I389840,I389628);
nand I_22768 (I389933,I389450,I266194);
nor I_22769 (I389331,I389693,I389933);
not I_22770 (I389994,I2866);
DFFARX1 I_22771 (I86379,I2859,I389994,I390020,);
DFFARX1 I_22772 (I86391,I2859,I389994,I390037,);
not I_22773 (I390045,I390037);
not I_22774 (I390062,I86397);
nor I_22775 (I390079,I390062,I86382);
not I_22776 (I390096,I86373);
nor I_22777 (I390113,I390079,I86394);
nor I_22778 (I390130,I390037,I390113);
DFFARX1 I_22779 (I390130,I2859,I389994,I389980,);
nor I_22780 (I390161,I86394,I86382);
nand I_22781 (I390178,I390161,I86397);
DFFARX1 I_22782 (I390178,I2859,I389994,I389983,);
nor I_22783 (I390209,I390096,I86394);
nand I_22784 (I390226,I390209,I86376);
nor I_22785 (I390243,I390020,I390226);
DFFARX1 I_22786 (I390243,I2859,I389994,I389959,);
not I_22787 (I390274,I390226);
nand I_22788 (I389971,I390037,I390274);
DFFARX1 I_22789 (I390226,I2859,I389994,I390314,);
not I_22790 (I390322,I390314);
not I_22791 (I390339,I86394);
not I_22792 (I390356,I86385);
nor I_22793 (I390373,I390356,I86373);
nor I_22794 (I389986,I390322,I390373);
nor I_22795 (I390404,I390356,I86388);
and I_22796 (I390421,I390404,I86376);
or I_22797 (I390438,I390421,I86373);
DFFARX1 I_22798 (I390438,I2859,I389994,I390464,);
nor I_22799 (I389974,I390464,I390020);
not I_22800 (I390486,I390464);
and I_22801 (I390503,I390486,I390020);
nor I_22802 (I389968,I390045,I390503);
nand I_22803 (I390534,I390486,I390096);
nor I_22804 (I389962,I390356,I390534);
nand I_22805 (I389965,I390486,I390274);
nand I_22806 (I390579,I390096,I86385);
nor I_22807 (I389977,I390339,I390579);
not I_22808 (I390640,I2866);
DFFARX1 I_22809 (I476082,I2859,I390640,I390666,);
DFFARX1 I_22810 (I476064,I2859,I390640,I390683,);
not I_22811 (I390691,I390683);
not I_22812 (I390708,I476073);
nor I_22813 (I390725,I390708,I476085);
not I_22814 (I390742,I476067);
nor I_22815 (I390759,I390725,I476076);
nor I_22816 (I390776,I390683,I390759);
DFFARX1 I_22817 (I390776,I2859,I390640,I390626,);
nor I_22818 (I390807,I476076,I476085);
nand I_22819 (I390824,I390807,I476073);
DFFARX1 I_22820 (I390824,I2859,I390640,I390629,);
nor I_22821 (I390855,I390742,I476076);
nand I_22822 (I390872,I390855,I476088);
nor I_22823 (I390889,I390666,I390872);
DFFARX1 I_22824 (I390889,I2859,I390640,I390605,);
not I_22825 (I390920,I390872);
nand I_22826 (I390617,I390683,I390920);
DFFARX1 I_22827 (I390872,I2859,I390640,I390960,);
not I_22828 (I390968,I390960);
not I_22829 (I390985,I476076);
not I_22830 (I391002,I476064);
nor I_22831 (I391019,I391002,I476067);
nor I_22832 (I390632,I390968,I391019);
nor I_22833 (I391050,I391002,I476070);
and I_22834 (I391067,I391050,I476079);
or I_22835 (I391084,I391067,I476067);
DFFARX1 I_22836 (I391084,I2859,I390640,I391110,);
nor I_22837 (I390620,I391110,I390666);
not I_22838 (I391132,I391110);
and I_22839 (I391149,I391132,I390666);
nor I_22840 (I390614,I390691,I391149);
nand I_22841 (I391180,I391132,I390742);
nor I_22842 (I390608,I391002,I391180);
nand I_22843 (I390611,I391132,I390920);
nand I_22844 (I391225,I390742,I476064);
nor I_22845 (I390623,I390985,I391225);
not I_22846 (I391286,I2866);
DFFARX1 I_22847 (I251735,I2859,I391286,I391312,);
DFFARX1 I_22848 (I251747,I2859,I391286,I391329,);
not I_22849 (I391337,I391329);
not I_22850 (I391354,I251756);
nor I_22851 (I391371,I391354,I251732);
not I_22852 (I391388,I251750);
nor I_22853 (I391405,I391371,I251744);
nor I_22854 (I391422,I391329,I391405);
DFFARX1 I_22855 (I391422,I2859,I391286,I391272,);
nor I_22856 (I391453,I251744,I251732);
nand I_22857 (I391470,I391453,I251756);
DFFARX1 I_22858 (I391470,I2859,I391286,I391275,);
nor I_22859 (I391501,I391388,I251744);
nand I_22860 (I391518,I391501,I251738);
nor I_22861 (I391535,I391312,I391518);
DFFARX1 I_22862 (I391535,I2859,I391286,I391251,);
not I_22863 (I391566,I391518);
nand I_22864 (I391263,I391329,I391566);
DFFARX1 I_22865 (I391518,I2859,I391286,I391606,);
not I_22866 (I391614,I391606);
not I_22867 (I391631,I251744);
not I_22868 (I391648,I251753);
nor I_22869 (I391665,I391648,I251750);
nor I_22870 (I391278,I391614,I391665);
nor I_22871 (I391696,I391648,I251735);
and I_22872 (I391713,I391696,I251732);
or I_22873 (I391730,I391713,I251741);
DFFARX1 I_22874 (I391730,I2859,I391286,I391756,);
nor I_22875 (I391266,I391756,I391312);
not I_22876 (I391778,I391756);
and I_22877 (I391795,I391778,I391312);
nor I_22878 (I391260,I391337,I391795);
nand I_22879 (I391826,I391778,I391388);
nor I_22880 (I391254,I391648,I391826);
nand I_22881 (I391257,I391778,I391566);
nand I_22882 (I391871,I391388,I251753);
nor I_22883 (I391269,I391631,I391871);
not I_22884 (I391932,I2866);
DFFARX1 I_22885 (I110819,I2859,I391932,I391958,);
DFFARX1 I_22886 (I110825,I2859,I391932,I391975,);
not I_22887 (I391983,I391975);
not I_22888 (I392000,I110846);
nor I_22889 (I392017,I392000,I110834);
not I_22890 (I392034,I110843);
nor I_22891 (I392051,I392017,I110828);
nor I_22892 (I392068,I391975,I392051);
DFFARX1 I_22893 (I392068,I2859,I391932,I391918,);
nor I_22894 (I392099,I110828,I110834);
nand I_22895 (I392116,I392099,I110846);
DFFARX1 I_22896 (I392116,I2859,I391932,I391921,);
nor I_22897 (I392147,I392034,I110828);
nand I_22898 (I392164,I392147,I110819);
nor I_22899 (I392181,I391958,I392164);
DFFARX1 I_22900 (I392181,I2859,I391932,I391897,);
not I_22901 (I392212,I392164);
nand I_22902 (I391909,I391975,I392212);
DFFARX1 I_22903 (I392164,I2859,I391932,I392252,);
not I_22904 (I392260,I392252);
not I_22905 (I392277,I110828);
not I_22906 (I392294,I110831);
nor I_22907 (I392311,I392294,I110843);
nor I_22908 (I391924,I392260,I392311);
nor I_22909 (I392342,I392294,I110840);
and I_22910 (I392359,I392342,I110822);
or I_22911 (I392376,I392359,I110837);
DFFARX1 I_22912 (I392376,I2859,I391932,I392402,);
nor I_22913 (I391912,I392402,I391958);
not I_22914 (I392424,I392402);
and I_22915 (I392441,I392424,I391958);
nor I_22916 (I391906,I391983,I392441);
nand I_22917 (I392472,I392424,I392034);
nor I_22918 (I391900,I392294,I392472);
nand I_22919 (I391903,I392424,I392212);
nand I_22920 (I392517,I392034,I110831);
nor I_22921 (I391915,I392277,I392517);
not I_22922 (I392578,I2866);
DFFARX1 I_22923 (I6762,I2859,I392578,I392604,);
DFFARX1 I_22924 (I6768,I2859,I392578,I392621,);
not I_22925 (I392629,I392621);
not I_22926 (I392646,I6762);
nor I_22927 (I392663,I392646,I6774);
not I_22928 (I392680,I6786);
nor I_22929 (I392697,I392663,I6780);
nor I_22930 (I392714,I392621,I392697);
DFFARX1 I_22931 (I392714,I2859,I392578,I392564,);
nor I_22932 (I392745,I6780,I6774);
nand I_22933 (I392762,I392745,I6762);
DFFARX1 I_22934 (I392762,I2859,I392578,I392567,);
nor I_22935 (I392793,I392680,I6780);
nand I_22936 (I392810,I392793,I6765);
nor I_22937 (I392827,I392604,I392810);
DFFARX1 I_22938 (I392827,I2859,I392578,I392543,);
not I_22939 (I392858,I392810);
nand I_22940 (I392555,I392621,I392858);
DFFARX1 I_22941 (I392810,I2859,I392578,I392898,);
not I_22942 (I392906,I392898);
not I_22943 (I392923,I6780);
not I_22944 (I392940,I6765);
nor I_22945 (I392957,I392940,I6786);
nor I_22946 (I392570,I392906,I392957);
nor I_22947 (I392988,I392940,I6783);
and I_22948 (I393005,I392988,I6777);
or I_22949 (I393022,I393005,I6771);
DFFARX1 I_22950 (I393022,I2859,I392578,I393048,);
nor I_22951 (I392558,I393048,I392604);
not I_22952 (I393070,I393048);
and I_22953 (I393087,I393070,I392604);
nor I_22954 (I392552,I392629,I393087);
nand I_22955 (I393118,I393070,I392680);
nor I_22956 (I392546,I392940,I393118);
nand I_22957 (I392549,I393070,I392858);
nand I_22958 (I393163,I392680,I6765);
nor I_22959 (I392561,I392923,I393163);
not I_22960 (I393224,I2866);
DFFARX1 I_22961 (I89354,I2859,I393224,I393250,);
DFFARX1 I_22962 (I89366,I2859,I393224,I393267,);
not I_22963 (I393275,I393267);
not I_22964 (I393292,I89372);
nor I_22965 (I393309,I393292,I89357);
not I_22966 (I393326,I89348);
nor I_22967 (I393343,I393309,I89369);
nor I_22968 (I393360,I393267,I393343);
DFFARX1 I_22969 (I393360,I2859,I393224,I393210,);
nor I_22970 (I393391,I89369,I89357);
nand I_22971 (I393408,I393391,I89372);
DFFARX1 I_22972 (I393408,I2859,I393224,I393213,);
nor I_22973 (I393439,I393326,I89369);
nand I_22974 (I393456,I393439,I89351);
nor I_22975 (I393473,I393250,I393456);
DFFARX1 I_22976 (I393473,I2859,I393224,I393189,);
not I_22977 (I393504,I393456);
nand I_22978 (I393201,I393267,I393504);
DFFARX1 I_22979 (I393456,I2859,I393224,I393544,);
not I_22980 (I393552,I393544);
not I_22981 (I393569,I89369);
not I_22982 (I393586,I89360);
nor I_22983 (I393603,I393586,I89348);
nor I_22984 (I393216,I393552,I393603);
nor I_22985 (I393634,I393586,I89363);
and I_22986 (I393651,I393634,I89351);
or I_22987 (I393668,I393651,I89348);
DFFARX1 I_22988 (I393668,I2859,I393224,I393694,);
nor I_22989 (I393204,I393694,I393250);
not I_22990 (I393716,I393694);
and I_22991 (I393733,I393716,I393250);
nor I_22992 (I393198,I393275,I393733);
nand I_22993 (I393764,I393716,I393326);
nor I_22994 (I393192,I393586,I393764);
nand I_22995 (I393195,I393716,I393504);
nand I_22996 (I393809,I393326,I89360);
nor I_22997 (I393207,I393569,I393809);
not I_22998 (I393870,I2866);
DFFARX1 I_22999 (I200449,I2859,I393870,I393896,);
DFFARX1 I_23000 (I200446,I2859,I393870,I393913,);
not I_23001 (I393921,I393913);
not I_23002 (I393938,I200461);
nor I_23003 (I393955,I393938,I200464);
not I_23004 (I393972,I200452);
nor I_23005 (I393989,I393955,I200458);
nor I_23006 (I394006,I393913,I393989);
DFFARX1 I_23007 (I394006,I2859,I393870,I393856,);
nor I_23008 (I394037,I200458,I200464);
nand I_23009 (I394054,I394037,I200461);
DFFARX1 I_23010 (I394054,I2859,I393870,I393859,);
nor I_23011 (I394085,I393972,I200458);
nand I_23012 (I394102,I394085,I200470);
nor I_23013 (I394119,I393896,I394102);
DFFARX1 I_23014 (I394119,I2859,I393870,I393835,);
not I_23015 (I394150,I394102);
nand I_23016 (I393847,I393913,I394150);
DFFARX1 I_23017 (I394102,I2859,I393870,I394190,);
not I_23018 (I394198,I394190);
not I_23019 (I394215,I200458);
not I_23020 (I394232,I200443);
nor I_23021 (I394249,I394232,I200452);
nor I_23022 (I393862,I394198,I394249);
nor I_23023 (I394280,I394232,I200455);
and I_23024 (I394297,I394280,I200443);
or I_23025 (I394314,I394297,I200467);
DFFARX1 I_23026 (I394314,I2859,I393870,I394340,);
nor I_23027 (I393850,I394340,I393896);
not I_23028 (I394362,I394340);
and I_23029 (I394379,I394362,I393896);
nor I_23030 (I393844,I393921,I394379);
nand I_23031 (I394410,I394362,I393972);
nor I_23032 (I393838,I394232,I394410);
nand I_23033 (I393841,I394362,I394150);
nand I_23034 (I394455,I393972,I200443);
nor I_23035 (I393853,I394215,I394455);
not I_23036 (I394516,I2866);
DFFARX1 I_23037 (I483596,I2859,I394516,I394542,);
DFFARX1 I_23038 (I483578,I2859,I394516,I394559,);
not I_23039 (I394567,I394559);
not I_23040 (I394584,I483587);
nor I_23041 (I394601,I394584,I483599);
not I_23042 (I394618,I483581);
nor I_23043 (I394635,I394601,I483590);
nor I_23044 (I394652,I394559,I394635);
DFFARX1 I_23045 (I394652,I2859,I394516,I394502,);
nor I_23046 (I394683,I483590,I483599);
nand I_23047 (I394700,I394683,I483587);
DFFARX1 I_23048 (I394700,I2859,I394516,I394505,);
nor I_23049 (I394731,I394618,I483590);
nand I_23050 (I394748,I394731,I483602);
nor I_23051 (I394765,I394542,I394748);
DFFARX1 I_23052 (I394765,I2859,I394516,I394481,);
not I_23053 (I394796,I394748);
nand I_23054 (I394493,I394559,I394796);
DFFARX1 I_23055 (I394748,I2859,I394516,I394836,);
not I_23056 (I394844,I394836);
not I_23057 (I394861,I483590);
not I_23058 (I394878,I483578);
nor I_23059 (I394895,I394878,I483581);
nor I_23060 (I394508,I394844,I394895);
nor I_23061 (I394926,I394878,I483584);
and I_23062 (I394943,I394926,I483593);
or I_23063 (I394960,I394943,I483581);
DFFARX1 I_23064 (I394960,I2859,I394516,I394986,);
nor I_23065 (I394496,I394986,I394542);
not I_23066 (I395008,I394986);
and I_23067 (I395025,I395008,I394542);
nor I_23068 (I394490,I394567,I395025);
nand I_23069 (I395056,I395008,I394618);
nor I_23070 (I394484,I394878,I395056);
nand I_23071 (I394487,I395008,I394796);
nand I_23072 (I395101,I394618,I483578);
nor I_23073 (I394499,I394861,I395101);
not I_23074 (I395162,I2866);
DFFARX1 I_23075 (I254625,I2859,I395162,I395188,);
DFFARX1 I_23076 (I254637,I2859,I395162,I395205,);
not I_23077 (I395213,I395205);
not I_23078 (I395230,I254646);
nor I_23079 (I395247,I395230,I254622);
not I_23080 (I395264,I254640);
nor I_23081 (I395281,I395247,I254634);
nor I_23082 (I395298,I395205,I395281);
DFFARX1 I_23083 (I395298,I2859,I395162,I395148,);
nor I_23084 (I395329,I254634,I254622);
nand I_23085 (I395346,I395329,I254646);
DFFARX1 I_23086 (I395346,I2859,I395162,I395151,);
nor I_23087 (I395377,I395264,I254634);
nand I_23088 (I395394,I395377,I254628);
nor I_23089 (I395411,I395188,I395394);
DFFARX1 I_23090 (I395411,I2859,I395162,I395127,);
not I_23091 (I395442,I395394);
nand I_23092 (I395139,I395205,I395442);
DFFARX1 I_23093 (I395394,I2859,I395162,I395482,);
not I_23094 (I395490,I395482);
not I_23095 (I395507,I254634);
not I_23096 (I395524,I254643);
nor I_23097 (I395541,I395524,I254640);
nor I_23098 (I395154,I395490,I395541);
nor I_23099 (I395572,I395524,I254625);
and I_23100 (I395589,I395572,I254622);
or I_23101 (I395606,I395589,I254631);
DFFARX1 I_23102 (I395606,I2859,I395162,I395632,);
nor I_23103 (I395142,I395632,I395188);
not I_23104 (I395654,I395632);
and I_23105 (I395671,I395654,I395188);
nor I_23106 (I395136,I395213,I395671);
nand I_23107 (I395702,I395654,I395264);
nor I_23108 (I395130,I395524,I395702);
nand I_23109 (I395133,I395654,I395442);
nand I_23110 (I395747,I395264,I254643);
nor I_23111 (I395145,I395507,I395747);
not I_23112 (I395808,I2866);
DFFARX1 I_23113 (I273124,I2859,I395808,I395834,);
DFFARX1 I_23114 (I273118,I2859,I395808,I395851,);
not I_23115 (I395859,I395851);
not I_23116 (I395876,I273133);
nor I_23117 (I395893,I395876,I273118);
not I_23118 (I395910,I273127);
nor I_23119 (I395927,I395893,I273136);
nor I_23120 (I395944,I395851,I395927);
DFFARX1 I_23121 (I395944,I2859,I395808,I395794,);
nor I_23122 (I395975,I273136,I273118);
nand I_23123 (I395992,I395975,I273133);
DFFARX1 I_23124 (I395992,I2859,I395808,I395797,);
nor I_23125 (I396023,I395910,I273136);
nand I_23126 (I396040,I396023,I273121);
nor I_23127 (I396057,I395834,I396040);
DFFARX1 I_23128 (I396057,I2859,I395808,I395773,);
not I_23129 (I396088,I396040);
nand I_23130 (I395785,I395851,I396088);
DFFARX1 I_23131 (I396040,I2859,I395808,I396128,);
not I_23132 (I396136,I396128);
not I_23133 (I396153,I273136);
not I_23134 (I396170,I273130);
nor I_23135 (I396187,I396170,I273127);
nor I_23136 (I395800,I396136,I396187);
nor I_23137 (I396218,I396170,I273139);
and I_23138 (I396235,I396218,I273142);
or I_23139 (I396252,I396235,I273121);
DFFARX1 I_23140 (I396252,I2859,I395808,I396278,);
nor I_23141 (I395788,I396278,I395834);
not I_23142 (I396300,I396278);
and I_23143 (I396317,I396300,I395834);
nor I_23144 (I395782,I395859,I396317);
nand I_23145 (I396348,I396300,I395910);
nor I_23146 (I395776,I396170,I396348);
nand I_23147 (I395779,I396300,I396088);
nand I_23148 (I396393,I395910,I273130);
nor I_23149 (I395791,I396153,I396393);
not I_23150 (I396454,I2866);
DFFARX1 I_23151 (I186849,I2859,I396454,I396480,);
DFFARX1 I_23152 (I186846,I2859,I396454,I396497,);
not I_23153 (I396505,I396497);
not I_23154 (I396522,I186861);
nor I_23155 (I396539,I396522,I186864);
not I_23156 (I396556,I186852);
nor I_23157 (I396573,I396539,I186858);
nor I_23158 (I396590,I396497,I396573);
DFFARX1 I_23159 (I396590,I2859,I396454,I396440,);
nor I_23160 (I396621,I186858,I186864);
nand I_23161 (I396638,I396621,I186861);
DFFARX1 I_23162 (I396638,I2859,I396454,I396443,);
nor I_23163 (I396669,I396556,I186858);
nand I_23164 (I396686,I396669,I186870);
nor I_23165 (I396703,I396480,I396686);
DFFARX1 I_23166 (I396703,I2859,I396454,I396419,);
not I_23167 (I396734,I396686);
nand I_23168 (I396431,I396497,I396734);
DFFARX1 I_23169 (I396686,I2859,I396454,I396774,);
not I_23170 (I396782,I396774);
not I_23171 (I396799,I186858);
not I_23172 (I396816,I186843);
nor I_23173 (I396833,I396816,I186852);
nor I_23174 (I396446,I396782,I396833);
nor I_23175 (I396864,I396816,I186855);
and I_23176 (I396881,I396864,I186843);
or I_23177 (I396898,I396881,I186867);
DFFARX1 I_23178 (I396898,I2859,I396454,I396924,);
nor I_23179 (I396434,I396924,I396480);
not I_23180 (I396946,I396924);
and I_23181 (I396963,I396946,I396480);
nor I_23182 (I396428,I396505,I396963);
nand I_23183 (I396994,I396946,I396556);
nor I_23184 (I396422,I396816,I396994);
nand I_23185 (I396425,I396946,I396734);
nand I_23186 (I397039,I396556,I186843);
nor I_23187 (I396437,I396799,I397039);
not I_23188 (I397100,I2866);
DFFARX1 I_23189 (I173249,I2859,I397100,I397126,);
DFFARX1 I_23190 (I173246,I2859,I397100,I397143,);
not I_23191 (I397151,I397143);
not I_23192 (I397168,I173261);
nor I_23193 (I397185,I397168,I173264);
not I_23194 (I397202,I173252);
nor I_23195 (I397219,I397185,I173258);
nor I_23196 (I397236,I397143,I397219);
DFFARX1 I_23197 (I397236,I2859,I397100,I397086,);
nor I_23198 (I397267,I173258,I173264);
nand I_23199 (I397284,I397267,I173261);
DFFARX1 I_23200 (I397284,I2859,I397100,I397089,);
nor I_23201 (I397315,I397202,I173258);
nand I_23202 (I397332,I397315,I173270);
nor I_23203 (I397349,I397126,I397332);
DFFARX1 I_23204 (I397349,I2859,I397100,I397065,);
not I_23205 (I397380,I397332);
nand I_23206 (I397077,I397143,I397380);
DFFARX1 I_23207 (I397332,I2859,I397100,I397420,);
not I_23208 (I397428,I397420);
not I_23209 (I397445,I173258);
not I_23210 (I397462,I173243);
nor I_23211 (I397479,I397462,I173252);
nor I_23212 (I397092,I397428,I397479);
nor I_23213 (I397510,I397462,I173255);
and I_23214 (I397527,I397510,I173243);
or I_23215 (I397544,I397527,I173267);
DFFARX1 I_23216 (I397544,I2859,I397100,I397570,);
nor I_23217 (I397080,I397570,I397126);
not I_23218 (I397592,I397570);
and I_23219 (I397609,I397592,I397126);
nor I_23220 (I397074,I397151,I397609);
nand I_23221 (I397640,I397592,I397202);
nor I_23222 (I397068,I397462,I397640);
nand I_23223 (I397071,I397592,I397380);
nand I_23224 (I397685,I397202,I173243);
nor I_23225 (I397083,I397445,I397685);
not I_23226 (I397746,I2866);
DFFARX1 I_23227 (I500936,I2859,I397746,I397772,);
DFFARX1 I_23228 (I500918,I2859,I397746,I397789,);
not I_23229 (I397797,I397789);
not I_23230 (I397814,I500927);
nor I_23231 (I397831,I397814,I500939);
not I_23232 (I397848,I500921);
nor I_23233 (I397865,I397831,I500930);
nor I_23234 (I397882,I397789,I397865);
DFFARX1 I_23235 (I397882,I2859,I397746,I397732,);
nor I_23236 (I397913,I500930,I500939);
nand I_23237 (I397930,I397913,I500927);
DFFARX1 I_23238 (I397930,I2859,I397746,I397735,);
nor I_23239 (I397961,I397848,I500930);
nand I_23240 (I397978,I397961,I500942);
nor I_23241 (I397995,I397772,I397978);
DFFARX1 I_23242 (I397995,I2859,I397746,I397711,);
not I_23243 (I398026,I397978);
nand I_23244 (I397723,I397789,I398026);
DFFARX1 I_23245 (I397978,I2859,I397746,I398066,);
not I_23246 (I398074,I398066);
not I_23247 (I398091,I500930);
not I_23248 (I398108,I500918);
nor I_23249 (I398125,I398108,I500921);
nor I_23250 (I397738,I398074,I398125);
nor I_23251 (I398156,I398108,I500924);
and I_23252 (I398173,I398156,I500933);
or I_23253 (I398190,I398173,I500921);
DFFARX1 I_23254 (I398190,I2859,I397746,I398216,);
nor I_23255 (I397726,I398216,I397772);
not I_23256 (I398238,I398216);
and I_23257 (I398255,I398238,I397772);
nor I_23258 (I397720,I397797,I398255);
nand I_23259 (I398286,I398238,I397848);
nor I_23260 (I397714,I398108,I398286);
nand I_23261 (I397717,I398238,I398026);
nand I_23262 (I398331,I397848,I500918);
nor I_23263 (I397729,I398091,I398331);
not I_23264 (I398392,I2866);
DFFARX1 I_23265 (I451806,I2859,I398392,I398418,);
DFFARX1 I_23266 (I451788,I2859,I398392,I398435,);
not I_23267 (I398443,I398435);
not I_23268 (I398460,I451797);
nor I_23269 (I398477,I398460,I451809);
not I_23270 (I398494,I451791);
nor I_23271 (I398511,I398477,I451800);
nor I_23272 (I398528,I398435,I398511);
DFFARX1 I_23273 (I398528,I2859,I398392,I398378,);
nor I_23274 (I398559,I451800,I451809);
nand I_23275 (I398576,I398559,I451797);
DFFARX1 I_23276 (I398576,I2859,I398392,I398381,);
nor I_23277 (I398607,I398494,I451800);
nand I_23278 (I398624,I398607,I451812);
nor I_23279 (I398641,I398418,I398624);
DFFARX1 I_23280 (I398641,I2859,I398392,I398357,);
not I_23281 (I398672,I398624);
nand I_23282 (I398369,I398435,I398672);
DFFARX1 I_23283 (I398624,I2859,I398392,I398712,);
not I_23284 (I398720,I398712);
not I_23285 (I398737,I451800);
not I_23286 (I398754,I451788);
nor I_23287 (I398771,I398754,I451791);
nor I_23288 (I398384,I398720,I398771);
nor I_23289 (I398802,I398754,I451794);
and I_23290 (I398819,I398802,I451803);
or I_23291 (I398836,I398819,I451791);
DFFARX1 I_23292 (I398836,I2859,I398392,I398862,);
nor I_23293 (I398372,I398862,I398418);
not I_23294 (I398884,I398862);
and I_23295 (I398901,I398884,I398418);
nor I_23296 (I398366,I398443,I398901);
nand I_23297 (I398932,I398884,I398494);
nor I_23298 (I398360,I398754,I398932);
nand I_23299 (I398363,I398884,I398672);
nand I_23300 (I398977,I398494,I451788);
nor I_23301 (I398375,I398737,I398977);
not I_23302 (I399038,I2866);
DFFARX1 I_23303 (I333185,I2859,I399038,I399064,);
DFFARX1 I_23304 (I333182,I2859,I399038,I399081,);
not I_23305 (I399089,I399081);
not I_23306 (I399106,I333182);
nor I_23307 (I399123,I399106,I333185);
not I_23308 (I399140,I333197);
nor I_23309 (I399157,I399123,I333191);
nor I_23310 (I399174,I399081,I399157);
DFFARX1 I_23311 (I399174,I2859,I399038,I399024,);
nor I_23312 (I399205,I333191,I333185);
nand I_23313 (I399222,I399205,I333182);
DFFARX1 I_23314 (I399222,I2859,I399038,I399027,);
nor I_23315 (I399253,I399140,I333191);
nand I_23316 (I399270,I399253,I333179);
nor I_23317 (I399287,I399064,I399270);
DFFARX1 I_23318 (I399287,I2859,I399038,I399003,);
not I_23319 (I399318,I399270);
nand I_23320 (I399015,I399081,I399318);
DFFARX1 I_23321 (I399270,I2859,I399038,I399358,);
not I_23322 (I399366,I399358);
not I_23323 (I399383,I333191);
not I_23324 (I399400,I333188);
nor I_23325 (I399417,I399400,I333197);
nor I_23326 (I399030,I399366,I399417);
nor I_23327 (I399448,I399400,I333194);
and I_23328 (I399465,I399448,I333200);
or I_23329 (I399482,I399465,I333179);
DFFARX1 I_23330 (I399482,I2859,I399038,I399508,);
nor I_23331 (I399018,I399508,I399064);
not I_23332 (I399530,I399508);
and I_23333 (I399547,I399530,I399064);
nor I_23334 (I399012,I399089,I399547);
nand I_23335 (I399578,I399530,I399140);
nor I_23336 (I399006,I399400,I399578);
nand I_23337 (I399009,I399530,I399318);
nand I_23338 (I399623,I399140,I333188);
nor I_23339 (I399021,I399383,I399623);
not I_23340 (I399684,I2866);
DFFARX1 I_23341 (I216086,I2859,I399684,I399710,);
DFFARX1 I_23342 (I216098,I2859,I399684,I399727,);
not I_23343 (I399735,I399727);
not I_23344 (I399752,I216083);
nor I_23345 (I399769,I399752,I216101);
not I_23346 (I399786,I216107);
nor I_23347 (I399803,I399769,I216089);
nor I_23348 (I399820,I399727,I399803);
DFFARX1 I_23349 (I399820,I2859,I399684,I399670,);
nor I_23350 (I399851,I216089,I216101);
nand I_23351 (I399868,I399851,I216083);
DFFARX1 I_23352 (I399868,I2859,I399684,I399673,);
nor I_23353 (I399899,I399786,I216089);
nand I_23354 (I399916,I399899,I216092);
nor I_23355 (I399933,I399710,I399916);
DFFARX1 I_23356 (I399933,I2859,I399684,I399649,);
not I_23357 (I399964,I399916);
nand I_23358 (I399661,I399727,I399964);
DFFARX1 I_23359 (I399916,I2859,I399684,I400004,);
not I_23360 (I400012,I400004);
not I_23361 (I400029,I216089);
not I_23362 (I400046,I216095);
nor I_23363 (I400063,I400046,I216107);
nor I_23364 (I399676,I400012,I400063);
nor I_23365 (I400094,I400046,I216104);
and I_23366 (I400111,I400094,I216083);
or I_23367 (I400128,I400111,I216086);
DFFARX1 I_23368 (I400128,I2859,I399684,I400154,);
nor I_23369 (I399664,I400154,I399710);
not I_23370 (I400176,I400154);
and I_23371 (I400193,I400176,I399710);
nor I_23372 (I399658,I399735,I400193);
nand I_23373 (I400224,I400176,I399786);
nor I_23374 (I399652,I400046,I400224);
nand I_23375 (I399655,I400176,I399964);
nand I_23376 (I400269,I399786,I216095);
nor I_23377 (I399667,I400029,I400269);
not I_23378 (I400330,I2866);
DFFARX1 I_23379 (I113454,I2859,I400330,I400356,);
DFFARX1 I_23380 (I113460,I2859,I400330,I400373,);
not I_23381 (I400381,I400373);
not I_23382 (I400398,I113481);
nor I_23383 (I400415,I400398,I113469);
not I_23384 (I400432,I113478);
nor I_23385 (I400449,I400415,I113463);
nor I_23386 (I400466,I400373,I400449);
DFFARX1 I_23387 (I400466,I2859,I400330,I400316,);
nor I_23388 (I400497,I113463,I113469);
nand I_23389 (I400514,I400497,I113481);
DFFARX1 I_23390 (I400514,I2859,I400330,I400319,);
nor I_23391 (I400545,I400432,I113463);
nand I_23392 (I400562,I400545,I113454);
nor I_23393 (I400579,I400356,I400562);
DFFARX1 I_23394 (I400579,I2859,I400330,I400295,);
not I_23395 (I400610,I400562);
nand I_23396 (I400307,I400373,I400610);
DFFARX1 I_23397 (I400562,I2859,I400330,I400650,);
not I_23398 (I400658,I400650);
not I_23399 (I400675,I113463);
not I_23400 (I400692,I113466);
nor I_23401 (I400709,I400692,I113478);
nor I_23402 (I400322,I400658,I400709);
nor I_23403 (I400740,I400692,I113475);
and I_23404 (I400757,I400740,I113457);
or I_23405 (I400774,I400757,I113472);
DFFARX1 I_23406 (I400774,I2859,I400330,I400800,);
nor I_23407 (I400310,I400800,I400356);
not I_23408 (I400822,I400800);
and I_23409 (I400839,I400822,I400356);
nor I_23410 (I400304,I400381,I400839);
nand I_23411 (I400870,I400822,I400432);
nor I_23412 (I400298,I400692,I400870);
nand I_23413 (I400301,I400822,I400610);
nand I_23414 (I400915,I400432,I113466);
nor I_23415 (I400313,I400675,I400915);
not I_23416 (I400976,I2866);
DFFARX1 I_23417 (I285262,I2859,I400976,I401002,);
DFFARX1 I_23418 (I285256,I2859,I400976,I401019,);
not I_23419 (I401027,I401019);
not I_23420 (I401044,I285271);
nor I_23421 (I401061,I401044,I285256);
not I_23422 (I401078,I285265);
nor I_23423 (I401095,I401061,I285274);
nor I_23424 (I401112,I401019,I401095);
DFFARX1 I_23425 (I401112,I2859,I400976,I400962,);
nor I_23426 (I401143,I285274,I285256);
nand I_23427 (I401160,I401143,I285271);
DFFARX1 I_23428 (I401160,I2859,I400976,I400965,);
nor I_23429 (I401191,I401078,I285274);
nand I_23430 (I401208,I401191,I285259);
nor I_23431 (I401225,I401002,I401208);
DFFARX1 I_23432 (I401225,I2859,I400976,I400941,);
not I_23433 (I401256,I401208);
nand I_23434 (I400953,I401019,I401256);
DFFARX1 I_23435 (I401208,I2859,I400976,I401296,);
not I_23436 (I401304,I401296);
not I_23437 (I401321,I285274);
not I_23438 (I401338,I285268);
nor I_23439 (I401355,I401338,I285265);
nor I_23440 (I400968,I401304,I401355);
nor I_23441 (I401386,I401338,I285277);
and I_23442 (I401403,I401386,I285280);
or I_23443 (I401420,I401403,I285259);
DFFARX1 I_23444 (I401420,I2859,I400976,I401446,);
nor I_23445 (I400956,I401446,I401002);
not I_23446 (I401468,I401446);
and I_23447 (I401485,I401468,I401002);
nor I_23448 (I400950,I401027,I401485);
nand I_23449 (I401516,I401468,I401078);
nor I_23450 (I400944,I401338,I401516);
nand I_23451 (I400947,I401468,I401256);
nand I_23452 (I401561,I401078,I285268);
nor I_23453 (I400959,I401321,I401561);
not I_23454 (I401622,I2866);
DFFARX1 I_23455 (I187937,I2859,I401622,I401648,);
DFFARX1 I_23456 (I187934,I2859,I401622,I401665,);
not I_23457 (I401673,I401665);
not I_23458 (I401690,I187949);
nor I_23459 (I401707,I401690,I187952);
not I_23460 (I401724,I187940);
nor I_23461 (I401741,I401707,I187946);
nor I_23462 (I401758,I401665,I401741);
DFFARX1 I_23463 (I401758,I2859,I401622,I401608,);
nor I_23464 (I401789,I187946,I187952);
nand I_23465 (I401806,I401789,I187949);
DFFARX1 I_23466 (I401806,I2859,I401622,I401611,);
nor I_23467 (I401837,I401724,I187946);
nand I_23468 (I401854,I401837,I187958);
nor I_23469 (I401871,I401648,I401854);
DFFARX1 I_23470 (I401871,I2859,I401622,I401587,);
not I_23471 (I401902,I401854);
nand I_23472 (I401599,I401665,I401902);
DFFARX1 I_23473 (I401854,I2859,I401622,I401942,);
not I_23474 (I401950,I401942);
not I_23475 (I401967,I187946);
not I_23476 (I401984,I187931);
nor I_23477 (I402001,I401984,I187940);
nor I_23478 (I401614,I401950,I402001);
nor I_23479 (I402032,I401984,I187943);
and I_23480 (I402049,I402032,I187931);
or I_23481 (I402066,I402049,I187955);
DFFARX1 I_23482 (I402066,I2859,I401622,I402092,);
nor I_23483 (I401602,I402092,I401648);
not I_23484 (I402114,I402092);
and I_23485 (I402131,I402114,I401648);
nor I_23486 (I401596,I401673,I402131);
nand I_23487 (I402162,I402114,I401724);
nor I_23488 (I401590,I401984,I402162);
nand I_23489 (I401593,I402114,I401902);
nand I_23490 (I402207,I401724,I187931);
nor I_23491 (I401605,I401967,I402207);
not I_23492 (I402268,I2866);
DFFARX1 I_23493 (I547260,I2859,I402268,I402294,);
DFFARX1 I_23494 (I547284,I2859,I402268,I402311,);
not I_23495 (I402319,I402311);
not I_23496 (I402336,I547266);
nor I_23497 (I402353,I402336,I547275);
not I_23498 (I402370,I547260);
nor I_23499 (I402387,I402353,I547281);
nor I_23500 (I402404,I402311,I402387);
DFFARX1 I_23501 (I402404,I2859,I402268,I402254,);
nor I_23502 (I402435,I547281,I547275);
nand I_23503 (I402452,I402435,I547266);
DFFARX1 I_23504 (I402452,I2859,I402268,I402257,);
nor I_23505 (I402483,I402370,I547281);
nand I_23506 (I402500,I402483,I547278);
nor I_23507 (I402517,I402294,I402500);
DFFARX1 I_23508 (I402517,I2859,I402268,I402233,);
not I_23509 (I402548,I402500);
nand I_23510 (I402245,I402311,I402548);
DFFARX1 I_23511 (I402500,I2859,I402268,I402588,);
not I_23512 (I402596,I402588);
not I_23513 (I402613,I547281);
not I_23514 (I402630,I547272);
nor I_23515 (I402647,I402630,I547260);
nor I_23516 (I402260,I402596,I402647);
nor I_23517 (I402678,I402630,I547263);
and I_23518 (I402695,I402678,I547287);
or I_23519 (I402712,I402695,I547269);
DFFARX1 I_23520 (I402712,I2859,I402268,I402738,);
nor I_23521 (I402248,I402738,I402294);
not I_23522 (I402760,I402738);
and I_23523 (I402777,I402760,I402294);
nor I_23524 (I402242,I402319,I402777);
nand I_23525 (I402808,I402760,I402370);
nor I_23526 (I402236,I402630,I402808);
nand I_23527 (I402239,I402760,I402548);
nand I_23528 (I402853,I402370,I547272);
nor I_23529 (I402251,I402613,I402853);
not I_23530 (I402914,I2866);
DFFARX1 I_23531 (I438783,I2859,I402914,I402940,);
DFFARX1 I_23532 (I438786,I2859,I402914,I402957,);
not I_23533 (I402965,I402957);
not I_23534 (I402982,I438783);
nor I_23535 (I402999,I402982,I438795);
not I_23536 (I403016,I438804);
nor I_23537 (I403033,I402999,I438792);
nor I_23538 (I403050,I402957,I403033);
DFFARX1 I_23539 (I403050,I2859,I402914,I402900,);
nor I_23540 (I403081,I438792,I438795);
nand I_23541 (I403098,I403081,I438783);
DFFARX1 I_23542 (I403098,I2859,I402914,I402903,);
nor I_23543 (I403129,I403016,I438792);
nand I_23544 (I403146,I403129,I438798);
nor I_23545 (I403163,I402940,I403146);
DFFARX1 I_23546 (I403163,I2859,I402914,I402879,);
not I_23547 (I403194,I403146);
nand I_23548 (I402891,I402957,I403194);
DFFARX1 I_23549 (I403146,I2859,I402914,I403234,);
not I_23550 (I403242,I403234);
not I_23551 (I403259,I438792);
not I_23552 (I403276,I438789);
nor I_23553 (I403293,I403276,I438804);
nor I_23554 (I402906,I403242,I403293);
nor I_23555 (I403324,I403276,I438801);
and I_23556 (I403341,I403324,I438789);
or I_23557 (I403358,I403341,I438786);
DFFARX1 I_23558 (I403358,I2859,I402914,I403384,);
nor I_23559 (I402894,I403384,I402940);
not I_23560 (I403406,I403384);
and I_23561 (I403423,I403406,I402940);
nor I_23562 (I402888,I402965,I403423);
nand I_23563 (I403454,I403406,I403016);
nor I_23564 (I402882,I403276,I403454);
nand I_23565 (I402885,I403406,I403194);
nand I_23566 (I403499,I403016,I438789);
nor I_23567 (I402897,I403259,I403499);
not I_23568 (I403560,I2866);
DFFARX1 I_23569 (I517868,I2859,I403560,I403586,);
DFFARX1 I_23570 (I517874,I2859,I403560,I403603,);
not I_23571 (I403611,I403603);
not I_23572 (I403628,I517871);
nor I_23573 (I403645,I403628,I517850);
not I_23574 (I403662,I517853);
nor I_23575 (I403679,I403645,I517859);
nor I_23576 (I403696,I403603,I403679);
DFFARX1 I_23577 (I403696,I2859,I403560,I403546,);
nor I_23578 (I403727,I517859,I517850);
nand I_23579 (I403744,I403727,I517871);
DFFARX1 I_23580 (I403744,I2859,I403560,I403549,);
nor I_23581 (I403775,I403662,I517859);
nand I_23582 (I403792,I403775,I517853);
nor I_23583 (I403809,I403586,I403792);
DFFARX1 I_23584 (I403809,I2859,I403560,I403525,);
not I_23585 (I403840,I403792);
nand I_23586 (I403537,I403603,I403840);
DFFARX1 I_23587 (I403792,I2859,I403560,I403880,);
not I_23588 (I403888,I403880);
not I_23589 (I403905,I517859);
not I_23590 (I403922,I517862);
nor I_23591 (I403939,I403922,I517853);
nor I_23592 (I403552,I403888,I403939);
nor I_23593 (I403970,I403922,I517850);
and I_23594 (I403987,I403970,I517856);
or I_23595 (I404004,I403987,I517865);
DFFARX1 I_23596 (I404004,I2859,I403560,I404030,);
nor I_23597 (I403540,I404030,I403586);
not I_23598 (I404052,I404030);
and I_23599 (I404069,I404052,I403586);
nor I_23600 (I403534,I403611,I404069);
nand I_23601 (I404100,I404052,I403662);
nor I_23602 (I403528,I403922,I404100);
nand I_23603 (I403531,I404052,I403840);
nand I_23604 (I404145,I403662,I517862);
nor I_23605 (I403543,I403905,I404145);
not I_23606 (I404206,I2866);
DFFARX1 I_23607 (I86974,I2859,I404206,I404232,);
DFFARX1 I_23608 (I86986,I2859,I404206,I404249,);
not I_23609 (I404257,I404249);
not I_23610 (I404274,I86992);
nor I_23611 (I404291,I404274,I86977);
not I_23612 (I404308,I86968);
nor I_23613 (I404325,I404291,I86989);
nor I_23614 (I404342,I404249,I404325);
DFFARX1 I_23615 (I404342,I2859,I404206,I404192,);
nor I_23616 (I404373,I86989,I86977);
nand I_23617 (I404390,I404373,I86992);
DFFARX1 I_23618 (I404390,I2859,I404206,I404195,);
nor I_23619 (I404421,I404308,I86989);
nand I_23620 (I404438,I404421,I86971);
nor I_23621 (I404455,I404232,I404438);
DFFARX1 I_23622 (I404455,I2859,I404206,I404171,);
not I_23623 (I404486,I404438);
nand I_23624 (I404183,I404249,I404486);
DFFARX1 I_23625 (I404438,I2859,I404206,I404526,);
not I_23626 (I404534,I404526);
not I_23627 (I404551,I86989);
not I_23628 (I404568,I86980);
nor I_23629 (I404585,I404568,I86968);
nor I_23630 (I404198,I404534,I404585);
nor I_23631 (I404616,I404568,I86983);
and I_23632 (I404633,I404616,I86971);
or I_23633 (I404650,I404633,I86968);
DFFARX1 I_23634 (I404650,I2859,I404206,I404676,);
nor I_23635 (I404186,I404676,I404232);
not I_23636 (I404698,I404676);
and I_23637 (I404715,I404698,I404232);
nor I_23638 (I404180,I404257,I404715);
nand I_23639 (I404746,I404698,I404308);
nor I_23640 (I404174,I404568,I404746);
nand I_23641 (I404177,I404698,I404486);
nand I_23642 (I404791,I404308,I86980);
nor I_23643 (I404189,I404551,I404791);
not I_23644 (I404852,I2866);
DFFARX1 I_23645 (I344779,I2859,I404852,I404878,);
DFFARX1 I_23646 (I344776,I2859,I404852,I404895,);
not I_23647 (I404903,I404895);
not I_23648 (I404920,I344776);
nor I_23649 (I404937,I404920,I344779);
not I_23650 (I404954,I344791);
nor I_23651 (I404971,I404937,I344785);
nor I_23652 (I404988,I404895,I404971);
DFFARX1 I_23653 (I404988,I2859,I404852,I404838,);
nor I_23654 (I405019,I344785,I344779);
nand I_23655 (I405036,I405019,I344776);
DFFARX1 I_23656 (I405036,I2859,I404852,I404841,);
nor I_23657 (I405067,I404954,I344785);
nand I_23658 (I405084,I405067,I344773);
nor I_23659 (I405101,I404878,I405084);
DFFARX1 I_23660 (I405101,I2859,I404852,I404817,);
not I_23661 (I405132,I405084);
nand I_23662 (I404829,I404895,I405132);
DFFARX1 I_23663 (I405084,I2859,I404852,I405172,);
not I_23664 (I405180,I405172);
not I_23665 (I405197,I344785);
not I_23666 (I405214,I344782);
nor I_23667 (I405231,I405214,I344791);
nor I_23668 (I404844,I405180,I405231);
nor I_23669 (I405262,I405214,I344788);
and I_23670 (I405279,I405262,I344794);
or I_23671 (I405296,I405279,I344773);
DFFARX1 I_23672 (I405296,I2859,I404852,I405322,);
nor I_23673 (I404832,I405322,I404878);
not I_23674 (I405344,I405322);
and I_23675 (I405361,I405344,I404878);
nor I_23676 (I404826,I404903,I405361);
nand I_23677 (I405392,I405344,I404954);
nor I_23678 (I404820,I405214,I405392);
nand I_23679 (I404823,I405344,I405132);
nand I_23680 (I405437,I404954,I344782);
nor I_23681 (I404835,I405197,I405437);
not I_23682 (I405498,I2866);
DFFARX1 I_23683 (I223821,I2859,I405498,I405524,);
DFFARX1 I_23684 (I223833,I2859,I405498,I405541,);
not I_23685 (I405549,I405541);
not I_23686 (I405566,I223818);
nor I_23687 (I405583,I405566,I223836);
not I_23688 (I405600,I223842);
nor I_23689 (I405617,I405583,I223824);
nor I_23690 (I405634,I405541,I405617);
DFFARX1 I_23691 (I405634,I2859,I405498,I405484,);
nor I_23692 (I405665,I223824,I223836);
nand I_23693 (I405682,I405665,I223818);
DFFARX1 I_23694 (I405682,I2859,I405498,I405487,);
nor I_23695 (I405713,I405600,I223824);
nand I_23696 (I405730,I405713,I223827);
nor I_23697 (I405747,I405524,I405730);
DFFARX1 I_23698 (I405747,I2859,I405498,I405463,);
not I_23699 (I405778,I405730);
nand I_23700 (I405475,I405541,I405778);
DFFARX1 I_23701 (I405730,I2859,I405498,I405818,);
not I_23702 (I405826,I405818);
not I_23703 (I405843,I223824);
not I_23704 (I405860,I223830);
nor I_23705 (I405877,I405860,I223842);
nor I_23706 (I405490,I405826,I405877);
nor I_23707 (I405908,I405860,I223839);
and I_23708 (I405925,I405908,I223818);
or I_23709 (I405942,I405925,I223821);
DFFARX1 I_23710 (I405942,I2859,I405498,I405968,);
nor I_23711 (I405478,I405968,I405524);
not I_23712 (I405990,I405968);
and I_23713 (I406007,I405990,I405524);
nor I_23714 (I405472,I405549,I406007);
nand I_23715 (I406038,I405990,I405600);
nor I_23716 (I405466,I405860,I406038);
nand I_23717 (I405469,I405990,I405778);
nand I_23718 (I406083,I405600,I223830);
nor I_23719 (I405481,I405843,I406083);
not I_23720 (I406144,I2866);
DFFARX1 I_23721 (I328612,I2859,I406144,I406170,);
DFFARX1 I_23722 (I328606,I2859,I406144,I406187,);
not I_23723 (I406195,I406187);
not I_23724 (I406212,I328621);
nor I_23725 (I406229,I406212,I328606);
not I_23726 (I406246,I328615);
nor I_23727 (I406263,I406229,I328624);
nor I_23728 (I406280,I406187,I406263);
DFFARX1 I_23729 (I406280,I2859,I406144,I406130,);
nor I_23730 (I406311,I328624,I328606);
nand I_23731 (I406328,I406311,I328621);
DFFARX1 I_23732 (I406328,I2859,I406144,I406133,);
nor I_23733 (I406359,I406246,I328624);
nand I_23734 (I406376,I406359,I328609);
nor I_23735 (I406393,I406170,I406376);
DFFARX1 I_23736 (I406393,I2859,I406144,I406109,);
not I_23737 (I406424,I406376);
nand I_23738 (I406121,I406187,I406424);
DFFARX1 I_23739 (I406376,I2859,I406144,I406464,);
not I_23740 (I406472,I406464);
not I_23741 (I406489,I328624);
not I_23742 (I406506,I328618);
nor I_23743 (I406523,I406506,I328615);
nor I_23744 (I406136,I406472,I406523);
nor I_23745 (I406554,I406506,I328627);
and I_23746 (I406571,I406554,I328630);
or I_23747 (I406588,I406571,I328609);
DFFARX1 I_23748 (I406588,I2859,I406144,I406614,);
nor I_23749 (I406124,I406614,I406170);
not I_23750 (I406636,I406614);
and I_23751 (I406653,I406636,I406170);
nor I_23752 (I406118,I406195,I406653);
nand I_23753 (I406684,I406636,I406246);
nor I_23754 (I406112,I406506,I406684);
nand I_23755 (I406115,I406636,I406424);
nand I_23756 (I406729,I406246,I328618);
nor I_23757 (I406127,I406489,I406729);
not I_23758 (I406790,I2866);
DFFARX1 I_23759 (I98279,I2859,I406790,I406816,);
DFFARX1 I_23760 (I98291,I2859,I406790,I406833,);
not I_23761 (I406841,I406833);
not I_23762 (I406858,I98297);
nor I_23763 (I406875,I406858,I98282);
not I_23764 (I406892,I98273);
nor I_23765 (I406909,I406875,I98294);
nor I_23766 (I406926,I406833,I406909);
DFFARX1 I_23767 (I406926,I2859,I406790,I406776,);
nor I_23768 (I406957,I98294,I98282);
nand I_23769 (I406974,I406957,I98297);
DFFARX1 I_23770 (I406974,I2859,I406790,I406779,);
nor I_23771 (I407005,I406892,I98294);
nand I_23772 (I407022,I407005,I98276);
nor I_23773 (I407039,I406816,I407022);
DFFARX1 I_23774 (I407039,I2859,I406790,I406755,);
not I_23775 (I407070,I407022);
nand I_23776 (I406767,I406833,I407070);
DFFARX1 I_23777 (I407022,I2859,I406790,I407110,);
not I_23778 (I407118,I407110);
not I_23779 (I407135,I98294);
not I_23780 (I407152,I98285);
nor I_23781 (I407169,I407152,I98273);
nor I_23782 (I406782,I407118,I407169);
nor I_23783 (I407200,I407152,I98288);
and I_23784 (I407217,I407200,I98276);
or I_23785 (I407234,I407217,I98273);
DFFARX1 I_23786 (I407234,I2859,I406790,I407260,);
nor I_23787 (I406770,I407260,I406816);
not I_23788 (I407282,I407260);
and I_23789 (I407299,I407282,I406816);
nor I_23790 (I406764,I406841,I407299);
nand I_23791 (I407330,I407282,I406892);
nor I_23792 (I406758,I407152,I407330);
nand I_23793 (I406761,I407282,I407070);
nand I_23794 (I407375,I406892,I98285);
nor I_23795 (I406773,I407135,I407375);
not I_23796 (I407436,I2866);
DFFARX1 I_23797 (I226796,I2859,I407436,I407462,);
DFFARX1 I_23798 (I226808,I2859,I407436,I407479,);
not I_23799 (I407487,I407479);
not I_23800 (I407504,I226793);
nor I_23801 (I407521,I407504,I226811);
not I_23802 (I407538,I226817);
nor I_23803 (I407555,I407521,I226799);
nor I_23804 (I407572,I407479,I407555);
DFFARX1 I_23805 (I407572,I2859,I407436,I407422,);
nor I_23806 (I407603,I226799,I226811);
nand I_23807 (I407620,I407603,I226793);
DFFARX1 I_23808 (I407620,I2859,I407436,I407425,);
nor I_23809 (I407651,I407538,I226799);
nand I_23810 (I407668,I407651,I226802);
nor I_23811 (I407685,I407462,I407668);
DFFARX1 I_23812 (I407685,I2859,I407436,I407401,);
not I_23813 (I407716,I407668);
nand I_23814 (I407413,I407479,I407716);
DFFARX1 I_23815 (I407668,I2859,I407436,I407756,);
not I_23816 (I407764,I407756);
not I_23817 (I407781,I226799);
not I_23818 (I407798,I226805);
nor I_23819 (I407815,I407798,I226817);
nor I_23820 (I407428,I407764,I407815);
nor I_23821 (I407846,I407798,I226814);
and I_23822 (I407863,I407846,I226793);
or I_23823 (I407880,I407863,I226796);
DFFARX1 I_23824 (I407880,I2859,I407436,I407906,);
nor I_23825 (I407416,I407906,I407462);
not I_23826 (I407928,I407906);
and I_23827 (I407945,I407928,I407462);
nor I_23828 (I407410,I407487,I407945);
nand I_23829 (I407976,I407928,I407538);
nor I_23830 (I407404,I407798,I407976);
nand I_23831 (I407407,I407928,I407716);
nand I_23832 (I408021,I407538,I226805);
nor I_23833 (I407419,I407781,I408021);
not I_23834 (I408082,I2866);
DFFARX1 I_23835 (I447759,I2859,I408082,I408108,);
DFFARX1 I_23836 (I447762,I2859,I408082,I408125,);
not I_23837 (I408133,I408125);
not I_23838 (I408150,I447759);
nor I_23839 (I408167,I408150,I447771);
not I_23840 (I408184,I447780);
nor I_23841 (I408201,I408167,I447768);
nor I_23842 (I408218,I408125,I408201);
DFFARX1 I_23843 (I408218,I2859,I408082,I408068,);
nor I_23844 (I408249,I447768,I447771);
nand I_23845 (I408266,I408249,I447759);
DFFARX1 I_23846 (I408266,I2859,I408082,I408071,);
nor I_23847 (I408297,I408184,I447768);
nand I_23848 (I408314,I408297,I447774);
nor I_23849 (I408331,I408108,I408314);
DFFARX1 I_23850 (I408331,I2859,I408082,I408047,);
not I_23851 (I408362,I408314);
nand I_23852 (I408059,I408125,I408362);
DFFARX1 I_23853 (I408314,I2859,I408082,I408402,);
not I_23854 (I408410,I408402);
not I_23855 (I408427,I447768);
not I_23856 (I408444,I447765);
nor I_23857 (I408461,I408444,I447780);
nor I_23858 (I408074,I408410,I408461);
nor I_23859 (I408492,I408444,I447777);
and I_23860 (I408509,I408492,I447765);
or I_23861 (I408526,I408509,I447762);
DFFARX1 I_23862 (I408526,I2859,I408082,I408552,);
nor I_23863 (I408062,I408552,I408108);
not I_23864 (I408574,I408552);
and I_23865 (I408591,I408574,I408108);
nor I_23866 (I408056,I408133,I408591);
nand I_23867 (I408622,I408574,I408184);
nor I_23868 (I408050,I408444,I408622);
nand I_23869 (I408053,I408574,I408362);
nand I_23870 (I408667,I408184,I447765);
nor I_23871 (I408065,I408427,I408667);
not I_23872 (I408728,I2866);
DFFARX1 I_23873 (I540715,I2859,I408728,I408754,);
DFFARX1 I_23874 (I540739,I2859,I408728,I408771,);
not I_23875 (I408779,I408771);
not I_23876 (I408796,I540721);
nor I_23877 (I408813,I408796,I540730);
not I_23878 (I408830,I540715);
nor I_23879 (I408847,I408813,I540736);
nor I_23880 (I408864,I408771,I408847);
DFFARX1 I_23881 (I408864,I2859,I408728,I408714,);
nor I_23882 (I408895,I540736,I540730);
nand I_23883 (I408912,I408895,I540721);
DFFARX1 I_23884 (I408912,I2859,I408728,I408717,);
nor I_23885 (I408943,I408830,I540736);
nand I_23886 (I408960,I408943,I540733);
nor I_23887 (I408977,I408754,I408960);
DFFARX1 I_23888 (I408977,I2859,I408728,I408693,);
not I_23889 (I409008,I408960);
nand I_23890 (I408705,I408771,I409008);
DFFARX1 I_23891 (I408960,I2859,I408728,I409048,);
not I_23892 (I409056,I409048);
not I_23893 (I409073,I540736);
not I_23894 (I409090,I540727);
nor I_23895 (I409107,I409090,I540715);
nor I_23896 (I408720,I409056,I409107);
nor I_23897 (I409138,I409090,I540718);
and I_23898 (I409155,I409138,I540742);
or I_23899 (I409172,I409155,I540724);
DFFARX1 I_23900 (I409172,I2859,I408728,I409198,);
nor I_23901 (I408708,I409198,I408754);
not I_23902 (I409220,I409198);
and I_23903 (I409237,I409220,I408754);
nor I_23904 (I408702,I408779,I409237);
nand I_23905 (I409268,I409220,I408830);
nor I_23906 (I408696,I409090,I409268);
nand I_23907 (I408699,I409220,I409008);
nand I_23908 (I409313,I408830,I540727);
nor I_23909 (I408711,I409073,I409313);
not I_23910 (I409374,I2866);
DFFARX1 I_23911 (I208065,I2859,I409374,I409400,);
DFFARX1 I_23912 (I208062,I2859,I409374,I409417,);
not I_23913 (I409425,I409417);
not I_23914 (I409442,I208077);
nor I_23915 (I409459,I409442,I208080);
not I_23916 (I409476,I208068);
nor I_23917 (I409493,I409459,I208074);
nor I_23918 (I409510,I409417,I409493);
DFFARX1 I_23919 (I409510,I2859,I409374,I409360,);
nor I_23920 (I409541,I208074,I208080);
nand I_23921 (I409558,I409541,I208077);
DFFARX1 I_23922 (I409558,I2859,I409374,I409363,);
nor I_23923 (I409589,I409476,I208074);
nand I_23924 (I409606,I409589,I208086);
nor I_23925 (I409623,I409400,I409606);
DFFARX1 I_23926 (I409623,I2859,I409374,I409339,);
not I_23927 (I409654,I409606);
nand I_23928 (I409351,I409417,I409654);
DFFARX1 I_23929 (I409606,I2859,I409374,I409694,);
not I_23930 (I409702,I409694);
not I_23931 (I409719,I208074);
not I_23932 (I409736,I208059);
nor I_23933 (I409753,I409736,I208068);
nor I_23934 (I409366,I409702,I409753);
nor I_23935 (I409784,I409736,I208071);
and I_23936 (I409801,I409784,I208059);
or I_23937 (I409818,I409801,I208083);
DFFARX1 I_23938 (I409818,I2859,I409374,I409844,);
nor I_23939 (I409354,I409844,I409400);
not I_23940 (I409866,I409844);
and I_23941 (I409883,I409866,I409400);
nor I_23942 (I409348,I409425,I409883);
nand I_23943 (I409914,I409866,I409476);
nor I_23944 (I409342,I409736,I409914);
nand I_23945 (I409345,I409866,I409654);
nand I_23946 (I409959,I409476,I208059);
nor I_23947 (I409357,I409719,I409959);
not I_23948 (I410020,I2866);
DFFARX1 I_23949 (I456430,I2859,I410020,I410046,);
DFFARX1 I_23950 (I456412,I2859,I410020,I410063,);
not I_23951 (I410071,I410063);
not I_23952 (I410088,I456421);
nor I_23953 (I410105,I410088,I456433);
not I_23954 (I410122,I456415);
nor I_23955 (I410139,I410105,I456424);
nor I_23956 (I410156,I410063,I410139);
DFFARX1 I_23957 (I410156,I2859,I410020,I410006,);
nor I_23958 (I410187,I456424,I456433);
nand I_23959 (I410204,I410187,I456421);
DFFARX1 I_23960 (I410204,I2859,I410020,I410009,);
nor I_23961 (I410235,I410122,I456424);
nand I_23962 (I410252,I410235,I456436);
nor I_23963 (I410269,I410046,I410252);
DFFARX1 I_23964 (I410269,I2859,I410020,I409985,);
not I_23965 (I410300,I410252);
nand I_23966 (I409997,I410063,I410300);
DFFARX1 I_23967 (I410252,I2859,I410020,I410340,);
not I_23968 (I410348,I410340);
not I_23969 (I410365,I456424);
not I_23970 (I410382,I456412);
nor I_23971 (I410399,I410382,I456415);
nor I_23972 (I410012,I410348,I410399);
nor I_23973 (I410430,I410382,I456418);
and I_23974 (I410447,I410430,I456427);
or I_23975 (I410464,I410447,I456415);
DFFARX1 I_23976 (I410464,I2859,I410020,I410490,);
nor I_23977 (I410000,I410490,I410046);
not I_23978 (I410512,I410490);
and I_23979 (I410529,I410512,I410046);
nor I_23980 (I409994,I410071,I410529);
nand I_23981 (I410560,I410512,I410122);
nor I_23982 (I409988,I410382,I410560);
nand I_23983 (I409991,I410512,I410300);
nand I_23984 (I410605,I410122,I456412);
nor I_23985 (I410003,I410365,I410605);
not I_23986 (I410666,I2866);
DFFARX1 I_23987 (I44706,I2859,I410666,I410692,);
DFFARX1 I_23988 (I44712,I2859,I410666,I410709,);
not I_23989 (I410717,I410709);
not I_23990 (I410734,I44730);
nor I_23991 (I410751,I410734,I44709);
not I_23992 (I410768,I44715);
nor I_23993 (I410785,I410751,I44721);
nor I_23994 (I410802,I410709,I410785);
DFFARX1 I_23995 (I410802,I2859,I410666,I410652,);
nor I_23996 (I410833,I44721,I44709);
nand I_23997 (I410850,I410833,I44730);
DFFARX1 I_23998 (I410850,I2859,I410666,I410655,);
nor I_23999 (I410881,I410768,I44721);
nand I_24000 (I410898,I410881,I44727);
nor I_24001 (I410915,I410692,I410898);
DFFARX1 I_24002 (I410915,I2859,I410666,I410631,);
not I_24003 (I410946,I410898);
nand I_24004 (I410643,I410709,I410946);
DFFARX1 I_24005 (I410898,I2859,I410666,I410986,);
not I_24006 (I410994,I410986);
not I_24007 (I411011,I44721);
not I_24008 (I411028,I44709);
nor I_24009 (I411045,I411028,I44715);
nor I_24010 (I410658,I410994,I411045);
nor I_24011 (I411076,I411028,I44718);
and I_24012 (I411093,I411076,I44706);
or I_24013 (I411110,I411093,I44724);
DFFARX1 I_24014 (I411110,I2859,I410666,I411136,);
nor I_24015 (I410646,I411136,I410692);
not I_24016 (I411158,I411136);
and I_24017 (I411175,I411158,I410692);
nor I_24018 (I410640,I410717,I411175);
nand I_24019 (I411206,I411158,I410768);
nor I_24020 (I410634,I411028,I411206);
nand I_24021 (I410637,I411158,I410946);
nand I_24022 (I411251,I410768,I44709);
nor I_24023 (I410649,I411011,I411251);
not I_24024 (I411312,I2866);
DFFARX1 I_24025 (I195009,I2859,I411312,I411338,);
DFFARX1 I_24026 (I195006,I2859,I411312,I411355,);
not I_24027 (I411363,I411355);
not I_24028 (I411380,I195021);
nor I_24029 (I411397,I411380,I195024);
not I_24030 (I411414,I195012);
nor I_24031 (I411431,I411397,I195018);
nor I_24032 (I411448,I411355,I411431);
DFFARX1 I_24033 (I411448,I2859,I411312,I411298,);
nor I_24034 (I411479,I195018,I195024);
nand I_24035 (I411496,I411479,I195021);
DFFARX1 I_24036 (I411496,I2859,I411312,I411301,);
nor I_24037 (I411527,I411414,I195018);
nand I_24038 (I411544,I411527,I195030);
nor I_24039 (I411561,I411338,I411544);
DFFARX1 I_24040 (I411561,I2859,I411312,I411277,);
not I_24041 (I411592,I411544);
nand I_24042 (I411289,I411355,I411592);
DFFARX1 I_24043 (I411544,I2859,I411312,I411632,);
not I_24044 (I411640,I411632);
not I_24045 (I411657,I195018);
not I_24046 (I411674,I195003);
nor I_24047 (I411691,I411674,I195012);
nor I_24048 (I411304,I411640,I411691);
nor I_24049 (I411722,I411674,I195015);
and I_24050 (I411739,I411722,I195003);
or I_24051 (I411756,I411739,I195027);
DFFARX1 I_24052 (I411756,I2859,I411312,I411782,);
nor I_24053 (I411292,I411782,I411338);
not I_24054 (I411804,I411782);
and I_24055 (I411821,I411804,I411338);
nor I_24056 (I411286,I411363,I411821);
nand I_24057 (I411852,I411804,I411414);
nor I_24058 (I411280,I411674,I411852);
nand I_24059 (I411283,I411804,I411592);
nand I_24060 (I411897,I411414,I195003);
nor I_24061 (I411295,I411657,I411897);
not I_24062 (I411958,I2866);
DFFARX1 I_24063 (I174881,I2859,I411958,I411984,);
DFFARX1 I_24064 (I174878,I2859,I411958,I412001,);
not I_24065 (I412009,I412001);
not I_24066 (I412026,I174893);
nor I_24067 (I412043,I412026,I174896);
not I_24068 (I412060,I174884);
nor I_24069 (I412077,I412043,I174890);
nor I_24070 (I412094,I412001,I412077);
DFFARX1 I_24071 (I412094,I2859,I411958,I411944,);
nor I_24072 (I412125,I174890,I174896);
nand I_24073 (I412142,I412125,I174893);
DFFARX1 I_24074 (I412142,I2859,I411958,I411947,);
nor I_24075 (I412173,I412060,I174890);
nand I_24076 (I412190,I412173,I174902);
nor I_24077 (I412207,I411984,I412190);
DFFARX1 I_24078 (I412207,I2859,I411958,I411923,);
not I_24079 (I412238,I412190);
nand I_24080 (I411935,I412001,I412238);
DFFARX1 I_24081 (I412190,I2859,I411958,I412278,);
not I_24082 (I412286,I412278);
not I_24083 (I412303,I174890);
not I_24084 (I412320,I174875);
nor I_24085 (I412337,I412320,I174884);
nor I_24086 (I411950,I412286,I412337);
nor I_24087 (I412368,I412320,I174887);
and I_24088 (I412385,I412368,I174875);
or I_24089 (I412402,I412385,I174899);
DFFARX1 I_24090 (I412402,I2859,I411958,I412428,);
nor I_24091 (I411938,I412428,I411984);
not I_24092 (I412450,I412428);
and I_24093 (I412467,I412450,I411984);
nor I_24094 (I411932,I412009,I412467);
nand I_24095 (I412498,I412450,I412060);
nor I_24096 (I411926,I412320,I412498);
nand I_24097 (I411929,I412450,I412238);
nand I_24098 (I412543,I412060,I174875);
nor I_24099 (I411941,I412303,I412543);
not I_24100 (I412604,I2866);
DFFARX1 I_24101 (I142966,I2859,I412604,I412630,);
DFFARX1 I_24102 (I142972,I2859,I412604,I412647,);
not I_24103 (I412655,I412647);
not I_24104 (I412672,I142993);
nor I_24105 (I412689,I412672,I142981);
not I_24106 (I412706,I142990);
nor I_24107 (I412723,I412689,I142975);
nor I_24108 (I412740,I412647,I412723);
DFFARX1 I_24109 (I412740,I2859,I412604,I412590,);
nor I_24110 (I412771,I142975,I142981);
nand I_24111 (I412788,I412771,I142993);
DFFARX1 I_24112 (I412788,I2859,I412604,I412593,);
nor I_24113 (I412819,I412706,I142975);
nand I_24114 (I412836,I412819,I142966);
nor I_24115 (I412853,I412630,I412836);
DFFARX1 I_24116 (I412853,I2859,I412604,I412569,);
not I_24117 (I412884,I412836);
nand I_24118 (I412581,I412647,I412884);
DFFARX1 I_24119 (I412836,I2859,I412604,I412924,);
not I_24120 (I412932,I412924);
not I_24121 (I412949,I142975);
not I_24122 (I412966,I142978);
nor I_24123 (I412983,I412966,I142990);
nor I_24124 (I412596,I412932,I412983);
nor I_24125 (I413014,I412966,I142987);
and I_24126 (I413031,I413014,I142969);
or I_24127 (I413048,I413031,I142984);
DFFARX1 I_24128 (I413048,I2859,I412604,I413074,);
nor I_24129 (I412584,I413074,I412630);
not I_24130 (I413096,I413074);
and I_24131 (I413113,I413096,I412630);
nor I_24132 (I412578,I412655,I413113);
nand I_24133 (I413144,I413096,I412706);
nor I_24134 (I412572,I412966,I413144);
nand I_24135 (I412575,I413096,I412884);
nand I_24136 (I413189,I412706,I142978);
nor I_24137 (I412587,I412949,I413189);
not I_24138 (I413250,I2866);
DFFARX1 I_24139 (I566300,I2859,I413250,I413276,);
DFFARX1 I_24140 (I566324,I2859,I413250,I413293,);
not I_24141 (I413301,I413293);
not I_24142 (I413318,I566306);
nor I_24143 (I413335,I413318,I566315);
not I_24144 (I413352,I566300);
nor I_24145 (I413369,I413335,I566321);
nor I_24146 (I413386,I413293,I413369);
DFFARX1 I_24147 (I413386,I2859,I413250,I413236,);
nor I_24148 (I413417,I566321,I566315);
nand I_24149 (I413434,I413417,I566306);
DFFARX1 I_24150 (I413434,I2859,I413250,I413239,);
nor I_24151 (I413465,I413352,I566321);
nand I_24152 (I413482,I413465,I566318);
nor I_24153 (I413499,I413276,I413482);
DFFARX1 I_24154 (I413499,I2859,I413250,I413215,);
not I_24155 (I413530,I413482);
nand I_24156 (I413227,I413293,I413530);
DFFARX1 I_24157 (I413482,I2859,I413250,I413570,);
not I_24158 (I413578,I413570);
not I_24159 (I413595,I566321);
not I_24160 (I413612,I566312);
nor I_24161 (I413629,I413612,I566300);
nor I_24162 (I413242,I413578,I413629);
nor I_24163 (I413660,I413612,I566303);
and I_24164 (I413677,I413660,I566327);
or I_24165 (I413694,I413677,I566309);
DFFARX1 I_24166 (I413694,I2859,I413250,I413720,);
nor I_24167 (I413230,I413720,I413276);
not I_24168 (I413742,I413720);
and I_24169 (I413759,I413742,I413276);
nor I_24170 (I413224,I413301,I413759);
nand I_24171 (I413790,I413742,I413352);
nor I_24172 (I413218,I413612,I413790);
nand I_24173 (I413221,I413742,I413530);
nand I_24174 (I413835,I413352,I566312);
nor I_24175 (I413233,I413595,I413835);
not I_24176 (I413896,I2866);
DFFARX1 I_24177 (I316474,I2859,I413896,I413922,);
DFFARX1 I_24178 (I316468,I2859,I413896,I413939,);
not I_24179 (I413947,I413939);
not I_24180 (I413964,I316483);
nor I_24181 (I413981,I413964,I316468);
not I_24182 (I413998,I316477);
nor I_24183 (I414015,I413981,I316486);
nor I_24184 (I414032,I413939,I414015);
DFFARX1 I_24185 (I414032,I2859,I413896,I413882,);
nor I_24186 (I414063,I316486,I316468);
nand I_24187 (I414080,I414063,I316483);
DFFARX1 I_24188 (I414080,I2859,I413896,I413885,);
nor I_24189 (I414111,I413998,I316486);
nand I_24190 (I414128,I414111,I316471);
nor I_24191 (I414145,I413922,I414128);
DFFARX1 I_24192 (I414145,I2859,I413896,I413861,);
not I_24193 (I414176,I414128);
nand I_24194 (I413873,I413939,I414176);
DFFARX1 I_24195 (I414128,I2859,I413896,I414216,);
not I_24196 (I414224,I414216);
not I_24197 (I414241,I316486);
not I_24198 (I414258,I316480);
nor I_24199 (I414275,I414258,I316477);
nor I_24200 (I413888,I414224,I414275);
nor I_24201 (I414306,I414258,I316489);
and I_24202 (I414323,I414306,I316492);
or I_24203 (I414340,I414323,I316471);
DFFARX1 I_24204 (I414340,I2859,I413896,I414366,);
nor I_24205 (I413876,I414366,I413922);
not I_24206 (I414388,I414366);
and I_24207 (I414405,I414388,I413922);
nor I_24208 (I413870,I413947,I414405);
nand I_24209 (I414436,I414388,I413998);
nor I_24210 (I413864,I414258,I414436);
nand I_24211 (I413867,I414388,I414176);
nand I_24212 (I414481,I413998,I316480);
nor I_24213 (I413879,I414241,I414481);
not I_24214 (I414542,I2866);
DFFARX1 I_24215 (I219656,I2859,I414542,I414568,);
DFFARX1 I_24216 (I219668,I2859,I414542,I414585,);
not I_24217 (I414593,I414585);
not I_24218 (I414610,I219653);
nor I_24219 (I414627,I414610,I219671);
not I_24220 (I414644,I219677);
nor I_24221 (I414661,I414627,I219659);
nor I_24222 (I414678,I414585,I414661);
DFFARX1 I_24223 (I414678,I2859,I414542,I414528,);
nor I_24224 (I414709,I219659,I219671);
nand I_24225 (I414726,I414709,I219653);
DFFARX1 I_24226 (I414726,I2859,I414542,I414531,);
nor I_24227 (I414757,I414644,I219659);
nand I_24228 (I414774,I414757,I219662);
nor I_24229 (I414791,I414568,I414774);
DFFARX1 I_24230 (I414791,I2859,I414542,I414507,);
not I_24231 (I414822,I414774);
nand I_24232 (I414519,I414585,I414822);
DFFARX1 I_24233 (I414774,I2859,I414542,I414862,);
not I_24234 (I414870,I414862);
not I_24235 (I414887,I219659);
not I_24236 (I414904,I219665);
nor I_24237 (I414921,I414904,I219677);
nor I_24238 (I414534,I414870,I414921);
nor I_24239 (I414952,I414904,I219674);
and I_24240 (I414969,I414952,I219653);
or I_24241 (I414986,I414969,I219656);
DFFARX1 I_24242 (I414986,I2859,I414542,I415012,);
nor I_24243 (I414522,I415012,I414568);
not I_24244 (I415034,I415012);
and I_24245 (I415051,I415034,I414568);
nor I_24246 (I414516,I414593,I415051);
nand I_24247 (I415082,I415034,I414644);
nor I_24248 (I414510,I414904,I415082);
nand I_24249 (I414513,I415034,I414822);
nand I_24250 (I415127,I414644,I219665);
nor I_24251 (I414525,I414887,I415127);
not I_24252 (I415188,I2866);
DFFARX1 I_24253 (I197729,I2859,I415188,I415214,);
DFFARX1 I_24254 (I197726,I2859,I415188,I415231,);
not I_24255 (I415239,I415231);
not I_24256 (I415256,I197741);
nor I_24257 (I415273,I415256,I197744);
not I_24258 (I415290,I197732);
nor I_24259 (I415307,I415273,I197738);
nor I_24260 (I415324,I415231,I415307);
DFFARX1 I_24261 (I415324,I2859,I415188,I415174,);
nor I_24262 (I415355,I197738,I197744);
nand I_24263 (I415372,I415355,I197741);
DFFARX1 I_24264 (I415372,I2859,I415188,I415177,);
nor I_24265 (I415403,I415290,I197738);
nand I_24266 (I415420,I415403,I197750);
nor I_24267 (I415437,I415214,I415420);
DFFARX1 I_24268 (I415437,I2859,I415188,I415153,);
not I_24269 (I415468,I415420);
nand I_24270 (I415165,I415231,I415468);
DFFARX1 I_24271 (I415420,I2859,I415188,I415508,);
not I_24272 (I415516,I415508);
not I_24273 (I415533,I197738);
not I_24274 (I415550,I197723);
nor I_24275 (I415567,I415550,I197732);
nor I_24276 (I415180,I415516,I415567);
nor I_24277 (I415598,I415550,I197735);
and I_24278 (I415615,I415598,I197723);
or I_24279 (I415632,I415615,I197747);
DFFARX1 I_24280 (I415632,I2859,I415188,I415658,);
nor I_24281 (I415168,I415658,I415214);
not I_24282 (I415680,I415658);
and I_24283 (I415697,I415680,I415214);
nor I_24284 (I415162,I415239,I415697);
nand I_24285 (I415728,I415680,I415290);
nor I_24286 (I415156,I415550,I415728);
nand I_24287 (I415159,I415680,I415468);
nand I_24288 (I415773,I415290,I197723);
nor I_24289 (I415171,I415533,I415773);
not I_24290 (I415834,I2866);
DFFARX1 I_24291 (I373237,I2859,I415834,I415860,);
DFFARX1 I_24292 (I373234,I2859,I415834,I415877,);
not I_24293 (I415885,I415877);
not I_24294 (I415902,I373234);
nor I_24295 (I415919,I415902,I373237);
not I_24296 (I415936,I373249);
nor I_24297 (I415953,I415919,I373243);
nor I_24298 (I415970,I415877,I415953);
DFFARX1 I_24299 (I415970,I2859,I415834,I415820,);
nor I_24300 (I416001,I373243,I373237);
nand I_24301 (I416018,I416001,I373234);
DFFARX1 I_24302 (I416018,I2859,I415834,I415823,);
nor I_24303 (I416049,I415936,I373243);
nand I_24304 (I416066,I416049,I373231);
nor I_24305 (I416083,I415860,I416066);
DFFARX1 I_24306 (I416083,I2859,I415834,I415799,);
not I_24307 (I416114,I416066);
nand I_24308 (I415811,I415877,I416114);
DFFARX1 I_24309 (I416066,I2859,I415834,I416154,);
not I_24310 (I416162,I416154);
not I_24311 (I416179,I373243);
not I_24312 (I416196,I373240);
nor I_24313 (I416213,I416196,I373249);
nor I_24314 (I415826,I416162,I416213);
nor I_24315 (I416244,I416196,I373246);
and I_24316 (I416261,I416244,I373252);
or I_24317 (I416278,I416261,I373231);
DFFARX1 I_24318 (I416278,I2859,I415834,I416304,);
nor I_24319 (I415814,I416304,I415860);
not I_24320 (I416326,I416304);
and I_24321 (I416343,I416326,I415860);
nor I_24322 (I415808,I415885,I416343);
nand I_24323 (I416374,I416326,I415936);
nor I_24324 (I415802,I416196,I416374);
nand I_24325 (I415805,I416326,I416114);
nand I_24326 (I416419,I415936,I373240);
nor I_24327 (I415817,I416179,I416419);
not I_24328 (I416480,I2866);
DFFARX1 I_24329 (I565705,I2859,I416480,I416506,);
DFFARX1 I_24330 (I565729,I2859,I416480,I416523,);
not I_24331 (I416531,I416523);
not I_24332 (I416548,I565711);
nor I_24333 (I416565,I416548,I565720);
not I_24334 (I416582,I565705);
nor I_24335 (I416599,I416565,I565726);
nor I_24336 (I416616,I416523,I416599);
DFFARX1 I_24337 (I416616,I2859,I416480,I416466,);
nor I_24338 (I416647,I565726,I565720);
nand I_24339 (I416664,I416647,I565711);
DFFARX1 I_24340 (I416664,I2859,I416480,I416469,);
nor I_24341 (I416695,I416582,I565726);
nand I_24342 (I416712,I416695,I565723);
nor I_24343 (I416729,I416506,I416712);
DFFARX1 I_24344 (I416729,I2859,I416480,I416445,);
not I_24345 (I416760,I416712);
nand I_24346 (I416457,I416523,I416760);
DFFARX1 I_24347 (I416712,I2859,I416480,I416800,);
not I_24348 (I416808,I416800);
not I_24349 (I416825,I565726);
not I_24350 (I416842,I565717);
nor I_24351 (I416859,I416842,I565705);
nor I_24352 (I416472,I416808,I416859);
nor I_24353 (I416890,I416842,I565708);
and I_24354 (I416907,I416890,I565732);
or I_24355 (I416924,I416907,I565714);
DFFARX1 I_24356 (I416924,I2859,I416480,I416950,);
nor I_24357 (I416460,I416950,I416506);
not I_24358 (I416972,I416950);
and I_24359 (I416989,I416972,I416506);
nor I_24360 (I416454,I416531,I416989);
nand I_24361 (I417020,I416972,I416582);
nor I_24362 (I416448,I416842,I417020);
nand I_24363 (I416451,I416972,I416760);
nand I_24364 (I417065,I416582,I565717);
nor I_24365 (I416463,I416825,I417065);
not I_24366 (I417126,I2866);
DFFARX1 I_24367 (I477238,I2859,I417126,I417152,);
DFFARX1 I_24368 (I477220,I2859,I417126,I417169,);
not I_24369 (I417177,I417169);
not I_24370 (I417194,I477229);
nor I_24371 (I417211,I417194,I477241);
not I_24372 (I417228,I477223);
nor I_24373 (I417245,I417211,I477232);
nor I_24374 (I417262,I417169,I417245);
DFFARX1 I_24375 (I417262,I2859,I417126,I417112,);
nor I_24376 (I417293,I477232,I477241);
nand I_24377 (I417310,I417293,I477229);
DFFARX1 I_24378 (I417310,I2859,I417126,I417115,);
nor I_24379 (I417341,I417228,I477232);
nand I_24380 (I417358,I417341,I477244);
nor I_24381 (I417375,I417152,I417358);
DFFARX1 I_24382 (I417375,I2859,I417126,I417091,);
not I_24383 (I417406,I417358);
nand I_24384 (I417103,I417169,I417406);
DFFARX1 I_24385 (I417358,I2859,I417126,I417446,);
not I_24386 (I417454,I417446);
not I_24387 (I417471,I477232);
not I_24388 (I417488,I477220);
nor I_24389 (I417505,I417488,I477223);
nor I_24390 (I417118,I417454,I417505);
nor I_24391 (I417536,I417488,I477226);
and I_24392 (I417553,I417536,I477235);
or I_24393 (I417570,I417553,I477223);
DFFARX1 I_24394 (I417570,I2859,I417126,I417596,);
nor I_24395 (I417106,I417596,I417152);
not I_24396 (I417618,I417596);
and I_24397 (I417635,I417618,I417152);
nor I_24398 (I417100,I417177,I417635);
nand I_24399 (I417666,I417618,I417228);
nor I_24400 (I417094,I417488,I417666);
nand I_24401 (I417097,I417618,I417406);
nand I_24402 (I417711,I417228,I477220);
nor I_24403 (I417109,I417471,I417711);
not I_24404 (I417772,I2866);
DFFARX1 I_24405 (I492266,I2859,I417772,I417798,);
DFFARX1 I_24406 (I492248,I2859,I417772,I417815,);
not I_24407 (I417823,I417815);
not I_24408 (I417840,I492257);
nor I_24409 (I417857,I417840,I492269);
not I_24410 (I417874,I492251);
nor I_24411 (I417891,I417857,I492260);
nor I_24412 (I417908,I417815,I417891);
DFFARX1 I_24413 (I417908,I2859,I417772,I417758,);
nor I_24414 (I417939,I492260,I492269);
nand I_24415 (I417956,I417939,I492257);
DFFARX1 I_24416 (I417956,I2859,I417772,I417761,);
nor I_24417 (I417987,I417874,I492260);
nand I_24418 (I418004,I417987,I492272);
nor I_24419 (I418021,I417798,I418004);
DFFARX1 I_24420 (I418021,I2859,I417772,I417737,);
not I_24421 (I418052,I418004);
nand I_24422 (I417749,I417815,I418052);
DFFARX1 I_24423 (I418004,I2859,I417772,I418092,);
not I_24424 (I418100,I418092);
not I_24425 (I418117,I492260);
not I_24426 (I418134,I492248);
nor I_24427 (I418151,I418134,I492251);
nor I_24428 (I417764,I418100,I418151);
nor I_24429 (I418182,I418134,I492254);
and I_24430 (I418199,I418182,I492263);
or I_24431 (I418216,I418199,I492251);
DFFARX1 I_24432 (I418216,I2859,I417772,I418242,);
nor I_24433 (I417752,I418242,I417798);
not I_24434 (I418264,I418242);
and I_24435 (I418281,I418264,I417798);
nor I_24436 (I417746,I417823,I418281);
nand I_24437 (I418312,I418264,I417874);
nor I_24438 (I417740,I418134,I418312);
nand I_24439 (I417743,I418264,I418052);
nand I_24440 (I418357,I417874,I492248);
nor I_24441 (I417755,I418117,I418357);
not I_24442 (I418418,I2866);
DFFARX1 I_24443 (I347941,I2859,I418418,I418444,);
DFFARX1 I_24444 (I347938,I2859,I418418,I418461,);
not I_24445 (I418469,I418461);
not I_24446 (I418486,I347938);
nor I_24447 (I418503,I418486,I347941);
not I_24448 (I418520,I347953);
nor I_24449 (I418537,I418503,I347947);
nor I_24450 (I418554,I418461,I418537);
DFFARX1 I_24451 (I418554,I2859,I418418,I418404,);
nor I_24452 (I418585,I347947,I347941);
nand I_24453 (I418602,I418585,I347938);
DFFARX1 I_24454 (I418602,I2859,I418418,I418407,);
nor I_24455 (I418633,I418520,I347947);
nand I_24456 (I418650,I418633,I347935);
nor I_24457 (I418667,I418444,I418650);
DFFARX1 I_24458 (I418667,I2859,I418418,I418383,);
not I_24459 (I418698,I418650);
nand I_24460 (I418395,I418461,I418698);
DFFARX1 I_24461 (I418650,I2859,I418418,I418738,);
not I_24462 (I418746,I418738);
not I_24463 (I418763,I347947);
not I_24464 (I418780,I347944);
nor I_24465 (I418797,I418780,I347953);
nor I_24466 (I418410,I418746,I418797);
nor I_24467 (I418828,I418780,I347950);
and I_24468 (I418845,I418828,I347956);
or I_24469 (I418862,I418845,I347935);
DFFARX1 I_24470 (I418862,I2859,I418418,I418888,);
nor I_24471 (I418398,I418888,I418444);
not I_24472 (I418910,I418888);
and I_24473 (I418927,I418910,I418444);
nor I_24474 (I418392,I418469,I418927);
nand I_24475 (I418958,I418910,I418520);
nor I_24476 (I418386,I418780,I418958);
nand I_24477 (I418389,I418910,I418698);
nand I_24478 (I419003,I418520,I347944);
nor I_24479 (I418401,I418763,I419003);
not I_24480 (I419064,I2866);
DFFARX1 I_24481 (I330924,I2859,I419064,I419090,);
DFFARX1 I_24482 (I330918,I2859,I419064,I419107,);
not I_24483 (I419115,I419107);
not I_24484 (I419132,I330933);
nor I_24485 (I419149,I419132,I330918);
not I_24486 (I419166,I330927);
nor I_24487 (I419183,I419149,I330936);
nor I_24488 (I419200,I419107,I419183);
DFFARX1 I_24489 (I419200,I2859,I419064,I419050,);
nor I_24490 (I419231,I330936,I330918);
nand I_24491 (I419248,I419231,I330933);
DFFARX1 I_24492 (I419248,I2859,I419064,I419053,);
nor I_24493 (I419279,I419166,I330936);
nand I_24494 (I419296,I419279,I330921);
nor I_24495 (I419313,I419090,I419296);
DFFARX1 I_24496 (I419313,I2859,I419064,I419029,);
not I_24497 (I419344,I419296);
nand I_24498 (I419041,I419107,I419344);
DFFARX1 I_24499 (I419296,I2859,I419064,I419384,);
not I_24500 (I419392,I419384);
not I_24501 (I419409,I330936);
not I_24502 (I419426,I330930);
nor I_24503 (I419443,I419426,I330927);
nor I_24504 (I419056,I419392,I419443);
nor I_24505 (I419474,I419426,I330939);
and I_24506 (I419491,I419474,I330942);
or I_24507 (I419508,I419491,I330921);
DFFARX1 I_24508 (I419508,I2859,I419064,I419534,);
nor I_24509 (I419044,I419534,I419090);
not I_24510 (I419556,I419534);
and I_24511 (I419573,I419556,I419090);
nor I_24512 (I419038,I419115,I419573);
nand I_24513 (I419604,I419556,I419166);
nor I_24514 (I419032,I419426,I419604);
nand I_24515 (I419035,I419556,I419344);
nand I_24516 (I419649,I419166,I330930);
nor I_24517 (I419047,I419409,I419649);
not I_24518 (I419710,I2866);
DFFARX1 I_24519 (I255203,I2859,I419710,I419736,);
DFFARX1 I_24520 (I255215,I2859,I419710,I419753,);
not I_24521 (I419761,I419753);
not I_24522 (I419778,I255224);
nor I_24523 (I419795,I419778,I255200);
not I_24524 (I419812,I255218);
nor I_24525 (I419829,I419795,I255212);
nor I_24526 (I419846,I419753,I419829);
DFFARX1 I_24527 (I419846,I2859,I419710,I419696,);
nor I_24528 (I419877,I255212,I255200);
nand I_24529 (I419894,I419877,I255224);
DFFARX1 I_24530 (I419894,I2859,I419710,I419699,);
nor I_24531 (I419925,I419812,I255212);
nand I_24532 (I419942,I419925,I255206);
nor I_24533 (I419959,I419736,I419942);
DFFARX1 I_24534 (I419959,I2859,I419710,I419675,);
not I_24535 (I419990,I419942);
nand I_24536 (I419687,I419753,I419990);
DFFARX1 I_24537 (I419942,I2859,I419710,I420030,);
not I_24538 (I420038,I420030);
not I_24539 (I420055,I255212);
not I_24540 (I420072,I255221);
nor I_24541 (I420089,I420072,I255218);
nor I_24542 (I419702,I420038,I420089);
nor I_24543 (I420120,I420072,I255203);
and I_24544 (I420137,I420120,I255200);
or I_24545 (I420154,I420137,I255209);
DFFARX1 I_24546 (I420154,I2859,I419710,I420180,);
nor I_24547 (I419690,I420180,I419736);
not I_24548 (I420202,I420180);
and I_24549 (I420219,I420202,I419736);
nor I_24550 (I419684,I419761,I420219);
nand I_24551 (I420250,I420202,I419812);
nor I_24552 (I419678,I420072,I420250);
nand I_24553 (I419681,I420202,I419990);
nand I_24554 (I420295,I419812,I255221);
nor I_24555 (I419693,I420055,I420295);
not I_24556 (I420356,I2866);
DFFARX1 I_24557 (I272546,I2859,I420356,I420382,);
DFFARX1 I_24558 (I272540,I2859,I420356,I420399,);
not I_24559 (I420407,I420399);
not I_24560 (I420424,I272555);
nor I_24561 (I420441,I420424,I272540);
not I_24562 (I420458,I272549);
nor I_24563 (I420475,I420441,I272558);
nor I_24564 (I420492,I420399,I420475);
DFFARX1 I_24565 (I420492,I2859,I420356,I420342,);
nor I_24566 (I420523,I272558,I272540);
nand I_24567 (I420540,I420523,I272555);
DFFARX1 I_24568 (I420540,I2859,I420356,I420345,);
nor I_24569 (I420571,I420458,I272558);
nand I_24570 (I420588,I420571,I272543);
nor I_24571 (I420605,I420382,I420588);
DFFARX1 I_24572 (I420605,I2859,I420356,I420321,);
not I_24573 (I420636,I420588);
nand I_24574 (I420333,I420399,I420636);
DFFARX1 I_24575 (I420588,I2859,I420356,I420676,);
not I_24576 (I420684,I420676);
not I_24577 (I420701,I272558);
not I_24578 (I420718,I272552);
nor I_24579 (I420735,I420718,I272549);
nor I_24580 (I420348,I420684,I420735);
nor I_24581 (I420766,I420718,I272561);
and I_24582 (I420783,I420766,I272564);
or I_24583 (I420800,I420783,I272543);
DFFARX1 I_24584 (I420800,I2859,I420356,I420826,);
nor I_24585 (I420336,I420826,I420382);
not I_24586 (I420848,I420826);
and I_24587 (I420865,I420848,I420382);
nor I_24588 (I420330,I420407,I420865);
nand I_24589 (I420896,I420848,I420458);
nor I_24590 (I420324,I420718,I420896);
nand I_24591 (I420327,I420848,I420636);
nand I_24592 (I420941,I420458,I272552);
nor I_24593 (I420339,I420701,I420941);
not I_24594 (I421002,I2866);
DFFARX1 I_24595 (I304336,I2859,I421002,I421028,);
DFFARX1 I_24596 (I304330,I2859,I421002,I421045,);
not I_24597 (I421053,I421045);
not I_24598 (I421070,I304345);
nor I_24599 (I421087,I421070,I304330);
not I_24600 (I421104,I304339);
nor I_24601 (I421121,I421087,I304348);
nor I_24602 (I421138,I421045,I421121);
DFFARX1 I_24603 (I421138,I2859,I421002,I420988,);
nor I_24604 (I421169,I304348,I304330);
nand I_24605 (I421186,I421169,I304345);
DFFARX1 I_24606 (I421186,I2859,I421002,I420991,);
nor I_24607 (I421217,I421104,I304348);
nand I_24608 (I421234,I421217,I304333);
nor I_24609 (I421251,I421028,I421234);
DFFARX1 I_24610 (I421251,I2859,I421002,I420967,);
not I_24611 (I421282,I421234);
nand I_24612 (I420979,I421045,I421282);
DFFARX1 I_24613 (I421234,I2859,I421002,I421322,);
not I_24614 (I421330,I421322);
not I_24615 (I421347,I304348);
not I_24616 (I421364,I304342);
nor I_24617 (I421381,I421364,I304339);
nor I_24618 (I420994,I421330,I421381);
nor I_24619 (I421412,I421364,I304351);
and I_24620 (I421429,I421412,I304354);
or I_24621 (I421446,I421429,I304333);
DFFARX1 I_24622 (I421446,I2859,I421002,I421472,);
nor I_24623 (I420982,I421472,I421028);
not I_24624 (I421494,I421472);
and I_24625 (I421511,I421494,I421028);
nor I_24626 (I420976,I421053,I421511);
nand I_24627 (I421542,I421494,I421104);
nor I_24628 (I420970,I421364,I421542);
nand I_24629 (I420973,I421494,I421282);
nand I_24630 (I421587,I421104,I304342);
nor I_24631 (I420985,I421347,I421587);
not I_24632 (I421648,I2866);
DFFARX1 I_24633 (I312428,I2859,I421648,I421674,);
DFFARX1 I_24634 (I312422,I2859,I421648,I421691,);
not I_24635 (I421699,I421691);
not I_24636 (I421716,I312437);
nor I_24637 (I421733,I421716,I312422);
not I_24638 (I421750,I312431);
nor I_24639 (I421767,I421733,I312440);
nor I_24640 (I421784,I421691,I421767);
DFFARX1 I_24641 (I421784,I2859,I421648,I421634,);
nor I_24642 (I421815,I312440,I312422);
nand I_24643 (I421832,I421815,I312437);
DFFARX1 I_24644 (I421832,I2859,I421648,I421637,);
nor I_24645 (I421863,I421750,I312440);
nand I_24646 (I421880,I421863,I312425);
nor I_24647 (I421897,I421674,I421880);
DFFARX1 I_24648 (I421897,I2859,I421648,I421613,);
not I_24649 (I421928,I421880);
nand I_24650 (I421625,I421691,I421928);
DFFARX1 I_24651 (I421880,I2859,I421648,I421968,);
not I_24652 (I421976,I421968);
not I_24653 (I421993,I312440);
not I_24654 (I422010,I312434);
nor I_24655 (I422027,I422010,I312431);
nor I_24656 (I421640,I421976,I422027);
nor I_24657 (I422058,I422010,I312443);
and I_24658 (I422075,I422058,I312446);
or I_24659 (I422092,I422075,I312425);
DFFARX1 I_24660 (I422092,I2859,I421648,I422118,);
nor I_24661 (I421628,I422118,I421674);
not I_24662 (I422140,I422118);
and I_24663 (I422157,I422140,I421674);
nor I_24664 (I421622,I421699,I422157);
nand I_24665 (I422188,I422140,I421750);
nor I_24666 (I421616,I422010,I422188);
nand I_24667 (I421619,I422140,I421928);
nand I_24668 (I422233,I421750,I312434);
nor I_24669 (I421631,I421993,I422233);
not I_24670 (I422294,I2866);
DFFARX1 I_24671 (I425319,I2859,I422294,I422320,);
DFFARX1 I_24672 (I425322,I2859,I422294,I422337,);
not I_24673 (I422345,I422337);
not I_24674 (I422362,I425319);
nor I_24675 (I422379,I422362,I425331);
not I_24676 (I422396,I425340);
nor I_24677 (I422413,I422379,I425328);
nor I_24678 (I422430,I422337,I422413);
DFFARX1 I_24679 (I422430,I2859,I422294,I422280,);
nor I_24680 (I422461,I425328,I425331);
nand I_24681 (I422478,I422461,I425319);
DFFARX1 I_24682 (I422478,I2859,I422294,I422283,);
nor I_24683 (I422509,I422396,I425328);
nand I_24684 (I422526,I422509,I425334);
nor I_24685 (I422543,I422320,I422526);
DFFARX1 I_24686 (I422543,I2859,I422294,I422259,);
not I_24687 (I422574,I422526);
nand I_24688 (I422271,I422337,I422574);
DFFARX1 I_24689 (I422526,I2859,I422294,I422614,);
not I_24690 (I422622,I422614);
not I_24691 (I422639,I425328);
not I_24692 (I422656,I425325);
nor I_24693 (I422673,I422656,I425340);
nor I_24694 (I422286,I422622,I422673);
nor I_24695 (I422704,I422656,I425337);
and I_24696 (I422721,I422704,I425325);
or I_24697 (I422738,I422721,I425322);
DFFARX1 I_24698 (I422738,I2859,I422294,I422764,);
nor I_24699 (I422274,I422764,I422320);
not I_24700 (I422786,I422764);
and I_24701 (I422803,I422786,I422320);
nor I_24702 (I422268,I422345,I422803);
nand I_24703 (I422834,I422786,I422396);
nor I_24704 (I422262,I422656,I422834);
nand I_24705 (I422265,I422786,I422574);
nand I_24706 (I422879,I422396,I425325);
nor I_24707 (I422277,I422639,I422879);
not I_24708 (I422940,I2866);
DFFARX1 I_24709 (I479550,I2859,I422940,I422966,);
DFFARX1 I_24710 (I479532,I2859,I422940,I422983,);
not I_24711 (I422991,I422983);
not I_24712 (I423008,I479541);
nor I_24713 (I423025,I423008,I479553);
not I_24714 (I423042,I479535);
nor I_24715 (I423059,I423025,I479544);
nor I_24716 (I423076,I422983,I423059);
DFFARX1 I_24717 (I423076,I2859,I422940,I422926,);
nor I_24718 (I423107,I479544,I479553);
nand I_24719 (I423124,I423107,I479541);
DFFARX1 I_24720 (I423124,I2859,I422940,I422929,);
nor I_24721 (I423155,I423042,I479544);
nand I_24722 (I423172,I423155,I479556);
nor I_24723 (I423189,I422966,I423172);
DFFARX1 I_24724 (I423189,I2859,I422940,I422905,);
not I_24725 (I423220,I423172);
nand I_24726 (I422917,I422983,I423220);
DFFARX1 I_24727 (I423172,I2859,I422940,I423260,);
not I_24728 (I423268,I423260);
not I_24729 (I423285,I479544);
not I_24730 (I423302,I479532);
nor I_24731 (I423319,I423302,I479535);
nor I_24732 (I422932,I423268,I423319);
nor I_24733 (I423350,I423302,I479538);
and I_24734 (I423367,I423350,I479547);
or I_24735 (I423384,I423367,I479535);
DFFARX1 I_24736 (I423384,I2859,I422940,I423410,);
nor I_24737 (I422920,I423410,I422966);
not I_24738 (I423432,I423410);
and I_24739 (I423449,I423432,I422966);
nor I_24740 (I422914,I422991,I423449);
nand I_24741 (I423480,I423432,I423042);
nor I_24742 (I422908,I423302,I423480);
nand I_24743 (I422911,I423432,I423220);
nand I_24744 (I423525,I423042,I479532);
nor I_24745 (I422923,I423285,I423525);
not I_24746 (I423586,I2866);
DFFARX1 I_24747 (I361116,I2859,I423586,I423612,);
DFFARX1 I_24748 (I361113,I2859,I423586,I423629,);
not I_24749 (I423637,I423629);
not I_24750 (I423654,I361113);
nor I_24751 (I423671,I423654,I361116);
not I_24752 (I423688,I361128);
nor I_24753 (I423705,I423671,I361122);
nor I_24754 (I423722,I423629,I423705);
DFFARX1 I_24755 (I423722,I2859,I423586,I423572,);
nor I_24756 (I423753,I361122,I361116);
nand I_24757 (I423770,I423753,I361113);
DFFARX1 I_24758 (I423770,I2859,I423586,I423575,);
nor I_24759 (I423801,I423688,I361122);
nand I_24760 (I423818,I423801,I361110);
nor I_24761 (I423835,I423612,I423818);
DFFARX1 I_24762 (I423835,I2859,I423586,I423551,);
not I_24763 (I423866,I423818);
nand I_24764 (I423563,I423629,I423866);
DFFARX1 I_24765 (I423818,I2859,I423586,I423906,);
not I_24766 (I423914,I423906);
not I_24767 (I423931,I361122);
not I_24768 (I423948,I361119);
nor I_24769 (I423965,I423948,I361128);
nor I_24770 (I423578,I423914,I423965);
nor I_24771 (I423996,I423948,I361125);
and I_24772 (I424013,I423996,I361131);
or I_24773 (I424030,I424013,I361110);
DFFARX1 I_24774 (I424030,I2859,I423586,I424056,);
nor I_24775 (I423566,I424056,I423612);
not I_24776 (I424078,I424056);
and I_24777 (I424095,I424078,I423612);
nor I_24778 (I423560,I423637,I424095);
nand I_24779 (I424126,I424078,I423688);
nor I_24780 (I423554,I423948,I424126);
nand I_24781 (I423557,I424078,I423866);
nand I_24782 (I424171,I423688,I361119);
nor I_24783 (I423569,I423931,I424171);
not I_24784 (I424226,I2866);
DFFARX1 I_24785 (I409339,I2859,I424226,I424252,);
DFFARX1 I_24786 (I424252,I2859,I424226,I424269,);
not I_24787 (I424218,I424269);
not I_24788 (I424291,I424252);
DFFARX1 I_24789 (I409366,I2859,I424226,I424317,);
nand I_24790 (I424325,I424317,I409357);
not I_24791 (I424342,I409357);
not I_24792 (I424359,I409339);
nand I_24793 (I424376,I409351,I409354);
and I_24794 (I424393,I409351,I409354);
not I_24795 (I424410,I409363);
nand I_24796 (I424427,I424410,I424359);
nor I_24797 (I424200,I424427,I424325);
nor I_24798 (I424458,I424342,I424427);
nand I_24799 (I424203,I424393,I424458);
not I_24800 (I424489,I409348);
nor I_24801 (I424506,I424489,I409351);
nor I_24802 (I424523,I424506,I409363);
nor I_24803 (I424540,I424291,I424523);
DFFARX1 I_24804 (I424540,I2859,I424226,I424212,);
not I_24805 (I424571,I424506);
DFFARX1 I_24806 (I424571,I2859,I424226,I424215,);
and I_24807 (I424209,I424317,I424506);
nor I_24808 (I424616,I424489,I409342);
and I_24809 (I424633,I424616,I409345);
or I_24810 (I424650,I424633,I409360);
DFFARX1 I_24811 (I424650,I2859,I424226,I424676,);
nor I_24812 (I424684,I424676,I424410);
DFFARX1 I_24813 (I424684,I2859,I424226,I424197,);
nand I_24814 (I424715,I424676,I424317);
nand I_24815 (I424732,I424410,I424715);
nor I_24816 (I424206,I424732,I424376);
not I_24817 (I424787,I2866);
DFFARX1 I_24818 (I529787,I2859,I424787,I424813,);
DFFARX1 I_24819 (I424813,I2859,I424787,I424830,);
not I_24820 (I424779,I424830);
not I_24821 (I424852,I424813);
DFFARX1 I_24822 (I529784,I2859,I424787,I424878,);
nand I_24823 (I424886,I424878,I529790);
not I_24824 (I424903,I529790);
not I_24825 (I424920,I529799);
nand I_24826 (I424937,I529793,I529787);
and I_24827 (I424954,I529793,I529787);
not I_24828 (I424971,I529805);
nand I_24829 (I424988,I424971,I424920);
nor I_24830 (I424761,I424988,I424886);
nor I_24831 (I425019,I424903,I424988);
nand I_24832 (I424764,I424954,I425019);
not I_24833 (I425050,I529802);
nor I_24834 (I425067,I425050,I529793);
nor I_24835 (I425084,I425067,I529805);
nor I_24836 (I425101,I424852,I425084);
DFFARX1 I_24837 (I425101,I2859,I424787,I424773,);
not I_24838 (I425132,I425067);
DFFARX1 I_24839 (I425132,I2859,I424787,I424776,);
and I_24840 (I424770,I424878,I425067);
nor I_24841 (I425177,I425050,I529796);
and I_24842 (I425194,I425177,I529808);
or I_24843 (I425211,I425194,I529784);
DFFARX1 I_24844 (I425211,I2859,I424787,I425237,);
nor I_24845 (I425245,I425237,I424971);
DFFARX1 I_24846 (I425245,I2859,I424787,I424758,);
nand I_24847 (I425276,I425237,I424878);
nand I_24848 (I425293,I424971,I425276);
nor I_24849 (I424767,I425293,I424937);
not I_24850 (I425348,I2866);
DFFARX1 I_24851 (I559770,I2859,I425348,I425374,);
DFFARX1 I_24852 (I425374,I2859,I425348,I425391,);
not I_24853 (I425340,I425391);
not I_24854 (I425413,I425374);
DFFARX1 I_24855 (I559764,I2859,I425348,I425439,);
nand I_24856 (I425447,I425439,I559755);
not I_24857 (I425464,I559755);
not I_24858 (I425481,I559782);
nand I_24859 (I425498,I559767,I559776);
and I_24860 (I425515,I559767,I559776);
not I_24861 (I425532,I559761);
nand I_24862 (I425549,I425532,I425481);
nor I_24863 (I425322,I425549,I425447);
nor I_24864 (I425580,I425464,I425549);
nand I_24865 (I425325,I425515,I425580);
not I_24866 (I425611,I559779);
nor I_24867 (I425628,I425611,I559767);
nor I_24868 (I425645,I425628,I559761);
nor I_24869 (I425662,I425413,I425645);
DFFARX1 I_24870 (I425662,I2859,I425348,I425334,);
not I_24871 (I425693,I425628);
DFFARX1 I_24872 (I425693,I2859,I425348,I425337,);
and I_24873 (I425331,I425439,I425628);
nor I_24874 (I425738,I425611,I559773);
and I_24875 (I425755,I425738,I559755);
or I_24876 (I425772,I425755,I559758);
DFFARX1 I_24877 (I425772,I2859,I425348,I425798,);
nor I_24878 (I425806,I425798,I425532);
DFFARX1 I_24879 (I425806,I2859,I425348,I425319,);
nand I_24880 (I425837,I425798,I425439);
nand I_24881 (I425854,I425532,I425837);
nor I_24882 (I425328,I425854,I425498);
not I_24883 (I425909,I2866);
DFFARX1 I_24884 (I63766,I2859,I425909,I425935,);
DFFARX1 I_24885 (I425935,I2859,I425909,I425952,);
not I_24886 (I425901,I425952);
not I_24887 (I425974,I425935);
DFFARX1 I_24888 (I63781,I2859,I425909,I426000,);
nand I_24889 (I426008,I426000,I63763);
not I_24890 (I426025,I63763);
not I_24891 (I426042,I63772);
nand I_24892 (I426059,I63778,I63769);
and I_24893 (I426076,I63778,I63769);
not I_24894 (I426093,I63766);
nand I_24895 (I426110,I426093,I426042);
nor I_24896 (I425883,I426110,I426008);
nor I_24897 (I426141,I426025,I426110);
nand I_24898 (I425886,I426076,I426141);
not I_24899 (I426172,I63763);
nor I_24900 (I426189,I426172,I63778);
nor I_24901 (I426206,I426189,I63766);
nor I_24902 (I426223,I425974,I426206);
DFFARX1 I_24903 (I426223,I2859,I425909,I425895,);
not I_24904 (I426254,I426189);
DFFARX1 I_24905 (I426254,I2859,I425909,I425898,);
and I_24906 (I425892,I426000,I426189);
nor I_24907 (I426299,I426172,I63787);
and I_24908 (I426316,I426299,I63784);
or I_24909 (I426333,I426316,I63775);
DFFARX1 I_24910 (I426333,I2859,I425909,I426359,);
nor I_24911 (I426367,I426359,I426093);
DFFARX1 I_24912 (I426367,I2859,I425909,I425880,);
nand I_24913 (I426398,I426359,I426000);
nand I_24914 (I426415,I426093,I426398);
nor I_24915 (I425889,I426415,I426059);
not I_24916 (I426470,I2866);
DFFARX1 I_24917 (I277167,I2859,I426470,I426496,);
DFFARX1 I_24918 (I426496,I2859,I426470,I426513,);
not I_24919 (I426462,I426513);
not I_24920 (I426535,I426496);
DFFARX1 I_24921 (I277179,I2859,I426470,I426561,);
nand I_24922 (I426569,I426561,I277188);
not I_24923 (I426586,I277188);
not I_24924 (I426603,I277170);
nand I_24925 (I426620,I277173,I277164);
and I_24926 (I426637,I277173,I277164);
not I_24927 (I426654,I277182);
nand I_24928 (I426671,I426654,I426603);
nor I_24929 (I426444,I426671,I426569);
nor I_24930 (I426702,I426586,I426671);
nand I_24931 (I426447,I426637,I426702);
not I_24932 (I426733,I277185);
nor I_24933 (I426750,I426733,I277173);
nor I_24934 (I426767,I426750,I277182);
nor I_24935 (I426784,I426535,I426767);
DFFARX1 I_24936 (I426784,I2859,I426470,I426456,);
not I_24937 (I426815,I426750);
DFFARX1 I_24938 (I426815,I2859,I426470,I426459,);
and I_24939 (I426453,I426561,I426750);
nor I_24940 (I426860,I426733,I277164);
and I_24941 (I426877,I426860,I277176);
or I_24942 (I426894,I426877,I277167);
DFFARX1 I_24943 (I426894,I2859,I426470,I426920,);
nor I_24944 (I426928,I426920,I426654);
DFFARX1 I_24945 (I426928,I2859,I426470,I426441,);
nand I_24946 (I426959,I426920,I426561);
nand I_24947 (I426976,I426654,I426959);
nor I_24948 (I426450,I426976,I426620);
not I_24949 (I427031,I2866);
DFFARX1 I_24950 (I377039,I2859,I427031,I427057,);
DFFARX1 I_24951 (I427057,I2859,I427031,I427074,);
not I_24952 (I427023,I427074);
not I_24953 (I427096,I427057);
DFFARX1 I_24954 (I377066,I2859,I427031,I427122,);
nand I_24955 (I427130,I427122,I377057);
not I_24956 (I427147,I377057);
not I_24957 (I427164,I377039);
nand I_24958 (I427181,I377051,I377054);
and I_24959 (I427198,I377051,I377054);
not I_24960 (I427215,I377063);
nand I_24961 (I427232,I427215,I427164);
nor I_24962 (I427005,I427232,I427130);
nor I_24963 (I427263,I427147,I427232);
nand I_24964 (I427008,I427198,I427263);
not I_24965 (I427294,I377048);
nor I_24966 (I427311,I427294,I377051);
nor I_24967 (I427328,I427311,I377063);
nor I_24968 (I427345,I427096,I427328);
DFFARX1 I_24969 (I427345,I2859,I427031,I427017,);
not I_24970 (I427376,I427311);
DFFARX1 I_24971 (I427376,I2859,I427031,I427020,);
and I_24972 (I427014,I427122,I427311);
nor I_24973 (I427421,I427294,I377042);
and I_24974 (I427438,I427421,I377045);
or I_24975 (I427455,I427438,I377060);
DFFARX1 I_24976 (I427455,I2859,I427031,I427481,);
nor I_24977 (I427489,I427481,I427215);
DFFARX1 I_24978 (I427489,I2859,I427031,I427002,);
nand I_24979 (I427520,I427481,I427122);
nand I_24980 (I427537,I427215,I427520);
nor I_24981 (I427011,I427537,I427181);
not I_24982 (I427592,I2866);
DFFARX1 I_24983 (I284681,I2859,I427592,I427618,);
DFFARX1 I_24984 (I427618,I2859,I427592,I427635,);
not I_24985 (I427584,I427635);
not I_24986 (I427657,I427618);
DFFARX1 I_24987 (I284693,I2859,I427592,I427683,);
nand I_24988 (I427691,I427683,I284702);
not I_24989 (I427708,I284702);
not I_24990 (I427725,I284684);
nand I_24991 (I427742,I284687,I284678);
and I_24992 (I427759,I284687,I284678);
not I_24993 (I427776,I284696);
nand I_24994 (I427793,I427776,I427725);
nor I_24995 (I427566,I427793,I427691);
nor I_24996 (I427824,I427708,I427793);
nand I_24997 (I427569,I427759,I427824);
not I_24998 (I427855,I284699);
nor I_24999 (I427872,I427855,I284687);
nor I_25000 (I427889,I427872,I284696);
nor I_25001 (I427906,I427657,I427889);
DFFARX1 I_25002 (I427906,I2859,I427592,I427578,);
not I_25003 (I427937,I427872);
DFFARX1 I_25004 (I427937,I2859,I427592,I427581,);
and I_25005 (I427575,I427683,I427872);
nor I_25006 (I427982,I427855,I284678);
and I_25007 (I427999,I427982,I284690);
or I_25008 (I428016,I427999,I284681);
DFFARX1 I_25009 (I428016,I2859,I427592,I428042,);
nor I_25010 (I428050,I428042,I427776);
DFFARX1 I_25011 (I428050,I2859,I427592,I427563,);
nand I_25012 (I428081,I428042,I427683);
nand I_25013 (I428098,I427776,I428081);
nor I_25014 (I427572,I428098,I427742);
not I_25015 (I428153,I2866);
DFFARX1 I_25016 (I103036,I2859,I428153,I428179,);
DFFARX1 I_25017 (I428179,I2859,I428153,I428196,);
not I_25018 (I428145,I428196);
not I_25019 (I428218,I428179);
DFFARX1 I_25020 (I103051,I2859,I428153,I428244,);
nand I_25021 (I428252,I428244,I103033);
not I_25022 (I428269,I103033);
not I_25023 (I428286,I103042);
nand I_25024 (I428303,I103048,I103039);
and I_25025 (I428320,I103048,I103039);
not I_25026 (I428337,I103036);
nand I_25027 (I428354,I428337,I428286);
nor I_25028 (I428127,I428354,I428252);
nor I_25029 (I428385,I428269,I428354);
nand I_25030 (I428130,I428320,I428385);
not I_25031 (I428416,I103033);
nor I_25032 (I428433,I428416,I103048);
nor I_25033 (I428450,I428433,I103036);
nor I_25034 (I428467,I428218,I428450);
DFFARX1 I_25035 (I428467,I2859,I428153,I428139,);
not I_25036 (I428498,I428433);
DFFARX1 I_25037 (I428498,I2859,I428153,I428142,);
and I_25038 (I428136,I428244,I428433);
nor I_25039 (I428543,I428416,I103057);
and I_25040 (I428560,I428543,I103054);
or I_25041 (I428577,I428560,I103045);
DFFARX1 I_25042 (I428577,I2859,I428153,I428603,);
nor I_25043 (I428611,I428603,I428337);
DFFARX1 I_25044 (I428611,I2859,I428153,I428124,);
nand I_25045 (I428642,I428603,I428244);
nand I_25046 (I428659,I428337,I428642);
nor I_25047 (I428133,I428659,I428303);
not I_25048 (I428714,I2866);
DFFARX1 I_25049 (I125069,I2859,I428714,I428740,);
DFFARX1 I_25050 (I428740,I2859,I428714,I428757,);
not I_25051 (I428706,I428757);
not I_25052 (I428779,I428740);
DFFARX1 I_25053 (I125066,I2859,I428714,I428805,);
nand I_25054 (I428813,I428805,I125060);
not I_25055 (I428830,I125060);
not I_25056 (I428847,I125057);
nand I_25057 (I428864,I125051,I125048);
and I_25058 (I428881,I125051,I125048);
not I_25059 (I428898,I125063);
nand I_25060 (I428915,I428898,I428847);
nor I_25061 (I428688,I428915,I428813);
nor I_25062 (I428946,I428830,I428915);
nand I_25063 (I428691,I428881,I428946);
not I_25064 (I428977,I125075);
nor I_25065 (I428994,I428977,I125051);
nor I_25066 (I429011,I428994,I125063);
nor I_25067 (I429028,I428779,I429011);
DFFARX1 I_25068 (I429028,I2859,I428714,I428700,);
not I_25069 (I429059,I428994);
DFFARX1 I_25070 (I429059,I2859,I428714,I428703,);
and I_25071 (I428697,I428805,I428994);
nor I_25072 (I429104,I428977,I125072);
and I_25073 (I429121,I429104,I125048);
or I_25074 (I429138,I429121,I125054);
DFFARX1 I_25075 (I429138,I2859,I428714,I429164,);
nor I_25076 (I429172,I429164,I428898);
DFFARX1 I_25077 (I429172,I2859,I428714,I428685,);
nand I_25078 (I429203,I429164,I428805);
nand I_25079 (I429220,I428898,I429203);
nor I_25080 (I428694,I429220,I428864);
not I_25081 (I429275,I2866);
DFFARX1 I_25082 (I559175,I2859,I429275,I429301,);
DFFARX1 I_25083 (I429301,I2859,I429275,I429318,);
not I_25084 (I429267,I429318);
not I_25085 (I429340,I429301);
DFFARX1 I_25086 (I559169,I2859,I429275,I429366,);
nand I_25087 (I429374,I429366,I559160);
not I_25088 (I429391,I559160);
not I_25089 (I429408,I559187);
nand I_25090 (I429425,I559172,I559181);
and I_25091 (I429442,I559172,I559181);
not I_25092 (I429459,I559166);
nand I_25093 (I429476,I429459,I429408);
nor I_25094 (I429249,I429476,I429374);
nor I_25095 (I429507,I429391,I429476);
nand I_25096 (I429252,I429442,I429507);
not I_25097 (I429538,I559184);
nor I_25098 (I429555,I429538,I559172);
nor I_25099 (I429572,I429555,I559166);
nor I_25100 (I429589,I429340,I429572);
DFFARX1 I_25101 (I429589,I2859,I429275,I429261,);
not I_25102 (I429620,I429555);
DFFARX1 I_25103 (I429620,I2859,I429275,I429264,);
and I_25104 (I429258,I429366,I429555);
nor I_25105 (I429665,I429538,I559178);
and I_25106 (I429682,I429665,I559160);
or I_25107 (I429699,I429682,I559163);
DFFARX1 I_25108 (I429699,I2859,I429275,I429725,);
nor I_25109 (I429733,I429725,I429459);
DFFARX1 I_25110 (I429733,I2859,I429275,I429246,);
nand I_25111 (I429764,I429725,I429366);
nand I_25112 (I429781,I429459,I429764);
nor I_25113 (I429255,I429781,I429425);
not I_25114 (I429836,I2866);
DFFARX1 I_25115 (I30489,I2859,I429836,I429862,);
DFFARX1 I_25116 (I429862,I2859,I429836,I429879,);
not I_25117 (I429828,I429879);
not I_25118 (I429901,I429862);
DFFARX1 I_25119 (I30477,I2859,I429836,I429927,);
nand I_25120 (I429935,I429927,I30492);
not I_25121 (I429952,I30492);
not I_25122 (I429969,I30480);
nand I_25123 (I429986,I30501,I30495);
and I_25124 (I430003,I30501,I30495);
not I_25125 (I430020,I30483);
nand I_25126 (I430037,I430020,I429969);
nor I_25127 (I429810,I430037,I429935);
nor I_25128 (I430068,I429952,I430037);
nand I_25129 (I429813,I430003,I430068);
not I_25130 (I430099,I30486);
nor I_25131 (I430116,I430099,I30501);
nor I_25132 (I430133,I430116,I30483);
nor I_25133 (I430150,I429901,I430133);
DFFARX1 I_25134 (I430150,I2859,I429836,I429822,);
not I_25135 (I430181,I430116);
DFFARX1 I_25136 (I430181,I2859,I429836,I429825,);
and I_25137 (I429819,I429927,I430116);
nor I_25138 (I430226,I430099,I30480);
and I_25139 (I430243,I430226,I30477);
or I_25140 (I430260,I430243,I30498);
DFFARX1 I_25141 (I430260,I2859,I429836,I430286,);
nor I_25142 (I430294,I430286,I430020);
DFFARX1 I_25143 (I430294,I2859,I429836,I429807,);
nand I_25144 (I430325,I430286,I429927);
nand I_25145 (I430342,I430020,I430325);
nor I_25146 (I429816,I430342,I429986);
not I_25147 (I430397,I2866);
DFFARX1 I_25148 (I204819,I2859,I430397,I430423,);
DFFARX1 I_25149 (I430423,I2859,I430397,I430440,);
not I_25150 (I430389,I430440);
not I_25151 (I430462,I430423);
DFFARX1 I_25152 (I204807,I2859,I430397,I430488,);
nand I_25153 (I430496,I430488,I204813);
not I_25154 (I430513,I204813);
not I_25155 (I430530,I204810);
nand I_25156 (I430547,I204798,I204795);
and I_25157 (I430564,I204798,I204795);
not I_25158 (I430581,I204822);
nand I_25159 (I430598,I430581,I430530);
nor I_25160 (I430371,I430598,I430496);
nor I_25161 (I430629,I430513,I430598);
nand I_25162 (I430374,I430564,I430629);
not I_25163 (I430660,I204795);
nor I_25164 (I430677,I430660,I204798);
nor I_25165 (I430694,I430677,I204822);
nor I_25166 (I430711,I430462,I430694);
DFFARX1 I_25167 (I430711,I2859,I430397,I430383,);
not I_25168 (I430742,I430677);
DFFARX1 I_25169 (I430742,I2859,I430397,I430386,);
and I_25170 (I430380,I430488,I430677);
nor I_25171 (I430787,I430660,I204804);
and I_25172 (I430804,I430787,I204801);
or I_25173 (I430821,I430804,I204816);
DFFARX1 I_25174 (I430821,I2859,I430397,I430847,);
nor I_25175 (I430855,I430847,I430581);
DFFARX1 I_25176 (I430855,I2859,I430397,I430368,);
nand I_25177 (I430886,I430847,I430488);
nand I_25178 (I430903,I430581,I430886);
nor I_25179 (I430377,I430903,I430547);
not I_25180 (I430958,I2866);
DFFARX1 I_25181 (I560960,I2859,I430958,I430984,);
DFFARX1 I_25182 (I430984,I2859,I430958,I431001,);
not I_25183 (I430950,I431001);
not I_25184 (I431023,I430984);
DFFARX1 I_25185 (I560954,I2859,I430958,I431049,);
nand I_25186 (I431057,I431049,I560945);
not I_25187 (I431074,I560945);
not I_25188 (I431091,I560972);
nand I_25189 (I431108,I560957,I560966);
and I_25190 (I431125,I560957,I560966);
not I_25191 (I431142,I560951);
nand I_25192 (I431159,I431142,I431091);
nor I_25193 (I430932,I431159,I431057);
nor I_25194 (I431190,I431074,I431159);
nand I_25195 (I430935,I431125,I431190);
not I_25196 (I431221,I560969);
nor I_25197 (I431238,I431221,I560957);
nor I_25198 (I431255,I431238,I560951);
nor I_25199 (I431272,I431023,I431255);
DFFARX1 I_25200 (I431272,I2859,I430958,I430944,);
not I_25201 (I431303,I431238);
DFFARX1 I_25202 (I431303,I2859,I430958,I430947,);
and I_25203 (I430941,I431049,I431238);
nor I_25204 (I431348,I431221,I560963);
and I_25205 (I431365,I431348,I560945);
or I_25206 (I431382,I431365,I560948);
DFFARX1 I_25207 (I431382,I2859,I430958,I431408,);
nor I_25208 (I431416,I431408,I431142);
DFFARX1 I_25209 (I431416,I2859,I430958,I430929,);
nand I_25210 (I431447,I431408,I431049);
nand I_25211 (I431464,I431142,I431447);
nor I_25212 (I430938,I431464,I431108);
not I_25213 (I431519,I2866);
DFFARX1 I_25214 (I305489,I2859,I431519,I431545,);
DFFARX1 I_25215 (I431545,I2859,I431519,I431562,);
not I_25216 (I431511,I431562);
not I_25217 (I431584,I431545);
DFFARX1 I_25218 (I305501,I2859,I431519,I431610,);
nand I_25219 (I431618,I431610,I305510);
not I_25220 (I431635,I305510);
not I_25221 (I431652,I305492);
nand I_25222 (I431669,I305495,I305486);
and I_25223 (I431686,I305495,I305486);
not I_25224 (I431703,I305504);
nand I_25225 (I431720,I431703,I431652);
nor I_25226 (I431493,I431720,I431618);
nor I_25227 (I431751,I431635,I431720);
nand I_25228 (I431496,I431686,I431751);
not I_25229 (I431782,I305507);
nor I_25230 (I431799,I431782,I305495);
nor I_25231 (I431816,I431799,I305504);
nor I_25232 (I431833,I431584,I431816);
DFFARX1 I_25233 (I431833,I2859,I431519,I431505,);
not I_25234 (I431864,I431799);
DFFARX1 I_25235 (I431864,I2859,I431519,I431508,);
and I_25236 (I431502,I431610,I431799);
nor I_25237 (I431909,I431782,I305486);
and I_25238 (I431926,I431909,I305498);
or I_25239 (I431943,I431926,I305489);
DFFARX1 I_25240 (I431943,I2859,I431519,I431969,);
nor I_25241 (I431977,I431969,I431703);
DFFARX1 I_25242 (I431977,I2859,I431519,I431490,);
nand I_25243 (I432008,I431969,I431610);
nand I_25244 (I432025,I431703,I432008);
nor I_25245 (I431499,I432025,I431669);
not I_25246 (I432080,I2866);
DFFARX1 I_25247 (I249998,I2859,I432080,I432106,);
DFFARX1 I_25248 (I432106,I2859,I432080,I432123,);
not I_25249 (I432072,I432123);
not I_25250 (I432145,I432106);
DFFARX1 I_25251 (I250013,I2859,I432080,I432171,);
nand I_25252 (I432179,I432171,I250004);
not I_25253 (I432196,I250004);
not I_25254 (I432213,I250010);
nand I_25255 (I432230,I250007,I250016);
and I_25256 (I432247,I250007,I250016);
not I_25257 (I432264,I250001);
nand I_25258 (I432281,I432264,I432213);
nor I_25259 (I432054,I432281,I432179);
nor I_25260 (I432312,I432196,I432281);
nand I_25261 (I432057,I432247,I432312);
not I_25262 (I432343,I249998);
nor I_25263 (I432360,I432343,I250007);
nor I_25264 (I432377,I432360,I250001);
nor I_25265 (I432394,I432145,I432377);
DFFARX1 I_25266 (I432394,I2859,I432080,I432066,);
not I_25267 (I432425,I432360);
DFFARX1 I_25268 (I432425,I2859,I432080,I432069,);
and I_25269 (I432063,I432171,I432360);
nor I_25270 (I432470,I432343,I250022);
and I_25271 (I432487,I432470,I250001);
or I_25272 (I432504,I432487,I250019);
DFFARX1 I_25273 (I432504,I2859,I432080,I432530,);
nor I_25274 (I432538,I432530,I432264);
DFFARX1 I_25275 (I432538,I2859,I432080,I432051,);
nand I_25276 (I432569,I432530,I432171);
nand I_25277 (I432586,I432264,I432569);
nor I_25278 (I432060,I432586,I432230);
not I_25279 (I432641,I2866);
DFFARX1 I_25280 (I417737,I2859,I432641,I432667,);
DFFARX1 I_25281 (I432667,I2859,I432641,I432684,);
not I_25282 (I432633,I432684);
not I_25283 (I432706,I432667);
DFFARX1 I_25284 (I417764,I2859,I432641,I432732,);
nand I_25285 (I432740,I432732,I417755);
not I_25286 (I432757,I417755);
not I_25287 (I432774,I417737);
nand I_25288 (I432791,I417749,I417752);
and I_25289 (I432808,I417749,I417752);
not I_25290 (I432825,I417761);
nand I_25291 (I432842,I432825,I432774);
nor I_25292 (I432615,I432842,I432740);
nor I_25293 (I432873,I432757,I432842);
nand I_25294 (I432618,I432808,I432873);
not I_25295 (I432904,I417746);
nor I_25296 (I432921,I432904,I417749);
nor I_25297 (I432938,I432921,I417761);
nor I_25298 (I432955,I432706,I432938);
DFFARX1 I_25299 (I432955,I2859,I432641,I432627,);
not I_25300 (I432986,I432921);
DFFARX1 I_25301 (I432986,I2859,I432641,I432630,);
and I_25302 (I432624,I432732,I432921);
nor I_25303 (I433031,I432904,I417740);
and I_25304 (I433048,I433031,I417743);
or I_25305 (I433065,I433048,I417758);
DFFARX1 I_25306 (I433065,I2859,I432641,I433091,);
nor I_25307 (I433099,I433091,I432825);
DFFARX1 I_25308 (I433099,I2859,I432641,I432612,);
nand I_25309 (I433130,I433091,I432732);
nand I_25310 (I433147,I432825,I433130);
nor I_25311 (I432621,I433147,I432791);
not I_25312 (I433202,I2866);
DFFARX1 I_25313 (I512960,I2859,I433202,I433228,);
DFFARX1 I_25314 (I433228,I2859,I433202,I433245,);
not I_25315 (I433194,I433245);
not I_25316 (I433267,I433228);
DFFARX1 I_25317 (I512966,I2859,I433202,I433293,);
nand I_25318 (I433301,I433293,I512975);
not I_25319 (I433318,I512975);
not I_25320 (I433335,I512954);
nand I_25321 (I433352,I512957,I512957);
and I_25322 (I433369,I512957,I512957);
not I_25323 (I433386,I512969);
nand I_25324 (I433403,I433386,I433335);
nor I_25325 (I433176,I433403,I433301);
nor I_25326 (I433434,I433318,I433403);
nand I_25327 (I433179,I433369,I433434);
not I_25328 (I433465,I512963);
nor I_25329 (I433482,I433465,I512957);
nor I_25330 (I433499,I433482,I512969);
nor I_25331 (I433516,I433267,I433499);
DFFARX1 I_25332 (I433516,I2859,I433202,I433188,);
not I_25333 (I433547,I433482);
DFFARX1 I_25334 (I433547,I2859,I433202,I433191,);
and I_25335 (I433185,I433293,I433482);
nor I_25336 (I433592,I433465,I512978);
and I_25337 (I433609,I433592,I512954);
or I_25338 (I433626,I433609,I512972);
DFFARX1 I_25339 (I433626,I2859,I433202,I433652,);
nor I_25340 (I433660,I433652,I433386);
DFFARX1 I_25341 (I433660,I2859,I433202,I433173,);
nand I_25342 (I433691,I433652,I433293);
nand I_25343 (I433708,I433386,I433691);
nor I_25344 (I433182,I433708,I433352);
not I_25345 (I433763,I2866);
DFFARX1 I_25346 (I463941,I2859,I433763,I433789,);
DFFARX1 I_25347 (I433789,I2859,I433763,I433806,);
not I_25348 (I433755,I433806);
not I_25349 (I433828,I433789);
DFFARX1 I_25350 (I463932,I2859,I433763,I433854,);
nand I_25351 (I433862,I433854,I463929);
not I_25352 (I433879,I463929);
not I_25353 (I433896,I463938);
nand I_25354 (I433913,I463947,I463929);
and I_25355 (I433930,I463947,I463929);
not I_25356 (I433947,I463926);
nand I_25357 (I433964,I433947,I433896);
nor I_25358 (I433737,I433964,I433862);
nor I_25359 (I433995,I433879,I433964);
nand I_25360 (I433740,I433930,I433995);
not I_25361 (I434026,I463935);
nor I_25362 (I434043,I434026,I463947);
nor I_25363 (I434060,I434043,I463926);
nor I_25364 (I434077,I433828,I434060);
DFFARX1 I_25365 (I434077,I2859,I433763,I433749,);
not I_25366 (I434108,I434043);
DFFARX1 I_25367 (I434108,I2859,I433763,I433752,);
and I_25368 (I433746,I433854,I434043);
nor I_25369 (I434153,I434026,I463950);
and I_25370 (I434170,I434153,I463926);
or I_25371 (I434187,I434170,I463944);
DFFARX1 I_25372 (I434187,I2859,I433763,I434213,);
nor I_25373 (I434221,I434213,I433947);
DFFARX1 I_25374 (I434221,I2859,I433763,I433734,);
nand I_25375 (I434252,I434213,I433854);
nand I_25376 (I434269,I433947,I434252);
nor I_25377 (I433743,I434269,I433913);
not I_25378 (I434324,I2866);
DFFARX1 I_25379 (I496887,I2859,I434324,I434350,);
DFFARX1 I_25380 (I434350,I2859,I434324,I434367,);
not I_25381 (I434316,I434367);
not I_25382 (I434389,I434350);
DFFARX1 I_25383 (I496878,I2859,I434324,I434415,);
nand I_25384 (I434423,I434415,I496875);
not I_25385 (I434440,I496875);
not I_25386 (I434457,I496884);
nand I_25387 (I434474,I496893,I496875);
and I_25388 (I434491,I496893,I496875);
not I_25389 (I434508,I496872);
nand I_25390 (I434525,I434508,I434457);
nor I_25391 (I434298,I434525,I434423);
nor I_25392 (I434556,I434440,I434525);
nand I_25393 (I434301,I434491,I434556);
not I_25394 (I434587,I496881);
nor I_25395 (I434604,I434587,I496893);
nor I_25396 (I434621,I434604,I496872);
nor I_25397 (I434638,I434389,I434621);
DFFARX1 I_25398 (I434638,I2859,I434324,I434310,);
not I_25399 (I434669,I434604);
DFFARX1 I_25400 (I434669,I2859,I434324,I434313,);
and I_25401 (I434307,I434415,I434604);
nor I_25402 (I434714,I434587,I496896);
and I_25403 (I434731,I434714,I496872);
or I_25404 (I434748,I434731,I496890);
DFFARX1 I_25405 (I434748,I2859,I434324,I434774,);
nor I_25406 (I434782,I434774,I434508);
DFFARX1 I_25407 (I434782,I2859,I434324,I434295,);
nand I_25408 (I434813,I434774,I434415);
nand I_25409 (I434830,I434508,I434813);
nor I_25410 (I434304,I434830,I434474);
not I_25411 (I434885,I2866);
DFFARX1 I_25412 (I525741,I2859,I434885,I434911,);
DFFARX1 I_25413 (I434911,I2859,I434885,I434928,);
not I_25414 (I434877,I434928);
not I_25415 (I434950,I434911);
DFFARX1 I_25416 (I525738,I2859,I434885,I434976,);
nand I_25417 (I434984,I434976,I525744);
not I_25418 (I435001,I525744);
not I_25419 (I435018,I525753);
nand I_25420 (I435035,I525747,I525741);
and I_25421 (I435052,I525747,I525741);
not I_25422 (I435069,I525759);
nand I_25423 (I435086,I435069,I435018);
nor I_25424 (I434859,I435086,I434984);
nor I_25425 (I435117,I435001,I435086);
nand I_25426 (I434862,I435052,I435117);
not I_25427 (I435148,I525756);
nor I_25428 (I435165,I435148,I525747);
nor I_25429 (I435182,I435165,I525759);
nor I_25430 (I435199,I434950,I435182);
DFFARX1 I_25431 (I435199,I2859,I434885,I434871,);
not I_25432 (I435230,I435165);
DFFARX1 I_25433 (I435230,I2859,I434885,I434874,);
and I_25434 (I434868,I434976,I435165);
nor I_25435 (I435275,I435148,I525750);
and I_25436 (I435292,I435275,I525762);
or I_25437 (I435309,I435292,I525738);
DFFARX1 I_25438 (I435309,I2859,I434885,I435335,);
nor I_25439 (I435343,I435335,I435069);
DFFARX1 I_25440 (I435343,I2859,I434885,I434856,);
nand I_25441 (I435374,I435335,I434976);
nand I_25442 (I435391,I435069,I435374);
nor I_25443 (I434865,I435391,I435035);
not I_25444 (I435446,I2866);
DFFARX1 I_25445 (I473189,I2859,I435446,I435472,);
DFFARX1 I_25446 (I435472,I2859,I435446,I435489,);
not I_25447 (I435438,I435489);
not I_25448 (I435511,I435472);
DFFARX1 I_25449 (I473180,I2859,I435446,I435537,);
nand I_25450 (I435545,I435537,I473177);
not I_25451 (I435562,I473177);
not I_25452 (I435579,I473186);
nand I_25453 (I435596,I473195,I473177);
and I_25454 (I435613,I473195,I473177);
not I_25455 (I435630,I473174);
nand I_25456 (I435647,I435630,I435579);
nor I_25457 (I435420,I435647,I435545);
nor I_25458 (I435678,I435562,I435647);
nand I_25459 (I435423,I435613,I435678);
not I_25460 (I435709,I473183);
nor I_25461 (I435726,I435709,I473195);
nor I_25462 (I435743,I435726,I473174);
nor I_25463 (I435760,I435511,I435743);
DFFARX1 I_25464 (I435760,I2859,I435446,I435432,);
not I_25465 (I435791,I435726);
DFFARX1 I_25466 (I435791,I2859,I435446,I435435,);
and I_25467 (I435429,I435537,I435726);
nor I_25468 (I435836,I435709,I473198);
and I_25469 (I435853,I435836,I473174);
or I_25470 (I435870,I435853,I473192);
DFFARX1 I_25471 (I435870,I2859,I435446,I435896,);
nor I_25472 (I435904,I435896,I435630);
DFFARX1 I_25473 (I435904,I2859,I435446,I435417,);
nand I_25474 (I435935,I435896,I435537);
nand I_25475 (I435952,I435630,I435935);
nor I_25476 (I435426,I435952,I435596);
not I_25477 (I436007,I2866);
DFFARX1 I_25478 (I137190,I2859,I436007,I436033,);
DFFARX1 I_25479 (I436033,I2859,I436007,I436050,);
not I_25480 (I435999,I436050);
not I_25481 (I436072,I436033);
DFFARX1 I_25482 (I137187,I2859,I436007,I436098,);
nand I_25483 (I436106,I436098,I137181);
not I_25484 (I436123,I137181);
not I_25485 (I436140,I137178);
nand I_25486 (I436157,I137172,I137169);
and I_25487 (I436174,I137172,I137169);
not I_25488 (I436191,I137184);
nand I_25489 (I436208,I436191,I436140);
nor I_25490 (I435981,I436208,I436106);
nor I_25491 (I436239,I436123,I436208);
nand I_25492 (I435984,I436174,I436239);
not I_25493 (I436270,I137196);
nor I_25494 (I436287,I436270,I137172);
nor I_25495 (I436304,I436287,I137184);
nor I_25496 (I436321,I436072,I436304);
DFFARX1 I_25497 (I436321,I2859,I436007,I435993,);
not I_25498 (I436352,I436287);
DFFARX1 I_25499 (I436352,I2859,I436007,I435996,);
and I_25500 (I435990,I436098,I436287);
nor I_25501 (I436397,I436270,I137193);
and I_25502 (I436414,I436397,I137169);
or I_25503 (I436431,I436414,I137175);
DFFARX1 I_25504 (I436431,I2859,I436007,I436457,);
nor I_25505 (I436465,I436457,I436191);
DFFARX1 I_25506 (I436465,I2859,I436007,I435978,);
nand I_25507 (I436496,I436457,I436098);
nand I_25508 (I436513,I436191,I436496);
nor I_25509 (I435987,I436513,I436157);
not I_25510 (I436568,I2866);
DFFARX1 I_25511 (I51569,I2859,I436568,I436594,);
DFFARX1 I_25512 (I436594,I2859,I436568,I436611,);
not I_25513 (I436560,I436611);
not I_25514 (I436633,I436594);
DFFARX1 I_25515 (I51557,I2859,I436568,I436659,);
nand I_25516 (I436667,I436659,I51572);
not I_25517 (I436684,I51572);
not I_25518 (I436701,I51560);
nand I_25519 (I436718,I51581,I51575);
and I_25520 (I436735,I51581,I51575);
not I_25521 (I436752,I51563);
nand I_25522 (I436769,I436752,I436701);
nor I_25523 (I436542,I436769,I436667);
nor I_25524 (I436800,I436684,I436769);
nand I_25525 (I436545,I436735,I436800);
not I_25526 (I436831,I51566);
nor I_25527 (I436848,I436831,I51581);
nor I_25528 (I436865,I436848,I51563);
nor I_25529 (I436882,I436633,I436865);
DFFARX1 I_25530 (I436882,I2859,I436568,I436554,);
not I_25531 (I436913,I436848);
DFFARX1 I_25532 (I436913,I2859,I436568,I436557,);
and I_25533 (I436551,I436659,I436848);
nor I_25534 (I436958,I436831,I51560);
and I_25535 (I436975,I436958,I51557);
or I_25536 (I436992,I436975,I51578);
DFFARX1 I_25537 (I436992,I2859,I436568,I437018,);
nor I_25538 (I437026,I437018,I436752);
DFFARX1 I_25539 (I437026,I2859,I436568,I436539,);
nand I_25540 (I437057,I437018,I436659);
nand I_25541 (I437074,I436752,I437057);
nor I_25542 (I436548,I437074,I436718);
not I_25543 (I437129,I2866);
DFFARX1 I_25544 (I493419,I2859,I437129,I437155,);
DFFARX1 I_25545 (I437155,I2859,I437129,I437172,);
not I_25546 (I437121,I437172);
not I_25547 (I437194,I437155);
DFFARX1 I_25548 (I493410,I2859,I437129,I437220,);
nand I_25549 (I437228,I437220,I493407);
not I_25550 (I437245,I493407);
not I_25551 (I437262,I493416);
nand I_25552 (I437279,I493425,I493407);
and I_25553 (I437296,I493425,I493407);
not I_25554 (I437313,I493404);
nand I_25555 (I437330,I437313,I437262);
nor I_25556 (I437103,I437330,I437228);
nor I_25557 (I437361,I437245,I437330);
nand I_25558 (I437106,I437296,I437361);
not I_25559 (I437392,I493413);
nor I_25560 (I437409,I437392,I493425);
nor I_25561 (I437426,I437409,I493404);
nor I_25562 (I437443,I437194,I437426);
DFFARX1 I_25563 (I437443,I2859,I437129,I437115,);
not I_25564 (I437474,I437409);
DFFARX1 I_25565 (I437474,I2859,I437129,I437118,);
and I_25566 (I437112,I437220,I437409);
nor I_25567 (I437519,I437392,I493428);
and I_25568 (I437536,I437519,I493404);
or I_25569 (I437553,I437536,I493422);
DFFARX1 I_25570 (I437553,I2859,I437129,I437579,);
nor I_25571 (I437587,I437579,I437313);
DFFARX1 I_25572 (I437587,I2859,I437129,I437100,);
nand I_25573 (I437618,I437579,I437220);
nand I_25574 (I437635,I437313,I437618);
nor I_25575 (I437109,I437635,I437279);
not I_25576 (I437690,I2866);
DFFARX1 I_25577 (I388667,I2859,I437690,I437716,);
DFFARX1 I_25578 (I437716,I2859,I437690,I437733,);
not I_25579 (I437682,I437733);
not I_25580 (I437755,I437716);
DFFARX1 I_25581 (I388694,I2859,I437690,I437781,);
nand I_25582 (I437789,I437781,I388685);
not I_25583 (I437806,I388685);
not I_25584 (I437823,I388667);
nand I_25585 (I437840,I388679,I388682);
and I_25586 (I437857,I388679,I388682);
not I_25587 (I437874,I388691);
nand I_25588 (I437891,I437874,I437823);
nor I_25589 (I437664,I437891,I437789);
nor I_25590 (I437922,I437806,I437891);
nand I_25591 (I437667,I437857,I437922);
not I_25592 (I437953,I388676);
nor I_25593 (I437970,I437953,I388679);
nor I_25594 (I437987,I437970,I388691);
nor I_25595 (I438004,I437755,I437987);
DFFARX1 I_25596 (I438004,I2859,I437690,I437676,);
not I_25597 (I438035,I437970);
DFFARX1 I_25598 (I438035,I2859,I437690,I437679,);
and I_25599 (I437673,I437781,I437970);
nor I_25600 (I438080,I437953,I388670);
and I_25601 (I438097,I438080,I388673);
or I_25602 (I438114,I438097,I388688);
DFFARX1 I_25603 (I438114,I2859,I437690,I438140,);
nor I_25604 (I438148,I438140,I437874);
DFFARX1 I_25605 (I438148,I2859,I437690,I437661,);
nand I_25606 (I438179,I438140,I437781);
nand I_25607 (I438196,I437874,I438179);
nor I_25608 (I437670,I438196,I437840);
not I_25609 (I438251,I2866);
DFFARX1 I_25610 (I462785,I2859,I438251,I438277,);
DFFARX1 I_25611 (I438277,I2859,I438251,I438294,);
not I_25612 (I438243,I438294);
not I_25613 (I438316,I438277);
DFFARX1 I_25614 (I462776,I2859,I438251,I438342,);
nand I_25615 (I438350,I438342,I462773);
not I_25616 (I438367,I462773);
not I_25617 (I438384,I462782);
nand I_25618 (I438401,I462791,I462773);
and I_25619 (I438418,I462791,I462773);
not I_25620 (I438435,I462770);
nand I_25621 (I438452,I438435,I438384);
nor I_25622 (I438225,I438452,I438350);
nor I_25623 (I438483,I438367,I438452);
nand I_25624 (I438228,I438418,I438483);
not I_25625 (I438514,I462779);
nor I_25626 (I438531,I438514,I462791);
nor I_25627 (I438548,I438531,I462770);
nor I_25628 (I438565,I438316,I438548);
DFFARX1 I_25629 (I438565,I2859,I438251,I438237,);
not I_25630 (I438596,I438531);
DFFARX1 I_25631 (I438596,I2859,I438251,I438240,);
and I_25632 (I438234,I438342,I438531);
nor I_25633 (I438641,I438514,I462794);
and I_25634 (I438658,I438641,I462770);
or I_25635 (I438675,I438658,I462788);
DFFARX1 I_25636 (I438675,I2859,I438251,I438701,);
nor I_25637 (I438709,I438701,I438435);
DFFARX1 I_25638 (I438709,I2859,I438251,I438222,);
nand I_25639 (I438740,I438701,I438342);
nand I_25640 (I438757,I438435,I438740);
nor I_25641 (I438231,I438757,I438401);
not I_25642 (I438812,I2866);
DFFARX1 I_25643 (I267919,I2859,I438812,I438838,);
DFFARX1 I_25644 (I438838,I2859,I438812,I438855,);
not I_25645 (I438804,I438855);
not I_25646 (I438877,I438838);
DFFARX1 I_25647 (I267931,I2859,I438812,I438903,);
nand I_25648 (I438911,I438903,I267940);
not I_25649 (I438928,I267940);
not I_25650 (I438945,I267922);
nand I_25651 (I438962,I267925,I267916);
and I_25652 (I438979,I267925,I267916);
not I_25653 (I438996,I267934);
nand I_25654 (I439013,I438996,I438945);
nor I_25655 (I438786,I439013,I438911);
nor I_25656 (I439044,I438928,I439013);
nand I_25657 (I438789,I438979,I439044);
not I_25658 (I439075,I267937);
nor I_25659 (I439092,I439075,I267925);
nor I_25660 (I439109,I439092,I267934);
nor I_25661 (I439126,I438877,I439109);
DFFARX1 I_25662 (I439126,I2859,I438812,I438798,);
not I_25663 (I439157,I439092);
DFFARX1 I_25664 (I439157,I2859,I438812,I438801,);
and I_25665 (I438795,I438903,I439092);
nor I_25666 (I439202,I439075,I267916);
and I_25667 (I439219,I439202,I267928);
or I_25668 (I439236,I439219,I267919);
DFFARX1 I_25669 (I439236,I2859,I438812,I439262,);
nor I_25670 (I439270,I439262,I438996);
DFFARX1 I_25671 (I439270,I2859,I438812,I438783,);
nand I_25672 (I439301,I439262,I438903);
nand I_25673 (I439318,I438996,I439301);
nor I_25674 (I438792,I439318,I438962);
not I_25675 (I439373,I2866);
DFFARX1 I_25676 (I21530,I2859,I439373,I439399,);
DFFARX1 I_25677 (I439399,I2859,I439373,I439416,);
not I_25678 (I439365,I439416);
not I_25679 (I439438,I439399);
DFFARX1 I_25680 (I21518,I2859,I439373,I439464,);
nand I_25681 (I439472,I439464,I21533);
not I_25682 (I439489,I21533);
not I_25683 (I439506,I21521);
nand I_25684 (I439523,I21542,I21536);
and I_25685 (I439540,I21542,I21536);
not I_25686 (I439557,I21524);
nand I_25687 (I439574,I439557,I439506);
nor I_25688 (I439347,I439574,I439472);
nor I_25689 (I439605,I439489,I439574);
nand I_25690 (I439350,I439540,I439605);
not I_25691 (I439636,I21527);
nor I_25692 (I439653,I439636,I21542);
nor I_25693 (I439670,I439653,I21524);
nor I_25694 (I439687,I439438,I439670);
DFFARX1 I_25695 (I439687,I2859,I439373,I439359,);
not I_25696 (I439718,I439653);
DFFARX1 I_25697 (I439718,I2859,I439373,I439362,);
and I_25698 (I439356,I439464,I439653);
nor I_25699 (I439763,I439636,I21521);
and I_25700 (I439780,I439763,I21518);
or I_25701 (I439797,I439780,I21539);
DFFARX1 I_25702 (I439797,I2859,I439373,I439823,);
nor I_25703 (I439831,I439823,I439557);
DFFARX1 I_25704 (I439831,I2859,I439373,I439344,);
nand I_25705 (I439862,I439823,I439464);
nand I_25706 (I439879,I439557,I439862);
nor I_25707 (I439353,I439879,I439523);
not I_25708 (I439934,I2866);
DFFARX1 I_25709 (I296241,I2859,I439934,I439960,);
DFFARX1 I_25710 (I439960,I2859,I439934,I439977,);
not I_25711 (I439926,I439977);
not I_25712 (I439999,I439960);
DFFARX1 I_25713 (I296253,I2859,I439934,I440025,);
nand I_25714 (I440033,I440025,I296262);
not I_25715 (I440050,I296262);
not I_25716 (I440067,I296244);
nand I_25717 (I440084,I296247,I296238);
and I_25718 (I440101,I296247,I296238);
not I_25719 (I440118,I296256);
nand I_25720 (I440135,I440118,I440067);
nor I_25721 (I439908,I440135,I440033);
nor I_25722 (I440166,I440050,I440135);
nand I_25723 (I439911,I440101,I440166);
not I_25724 (I440197,I296259);
nor I_25725 (I440214,I440197,I296247);
nor I_25726 (I440231,I440214,I296256);
nor I_25727 (I440248,I439999,I440231);
DFFARX1 I_25728 (I440248,I2859,I439934,I439920,);
not I_25729 (I440279,I440214);
DFFARX1 I_25730 (I440279,I2859,I439934,I439923,);
and I_25731 (I439917,I440025,I440214);
nor I_25732 (I440324,I440197,I296238);
and I_25733 (I440341,I440324,I296250);
or I_25734 (I440358,I440341,I296241);
DFFARX1 I_25735 (I440358,I2859,I439934,I440384,);
nor I_25736 (I440392,I440384,I440118);
DFFARX1 I_25737 (I440392,I2859,I439934,I439905,);
nand I_25738 (I440423,I440384,I440025);
nand I_25739 (I440440,I440118,I440423);
nor I_25740 (I439914,I440440,I440084);
not I_25741 (I440495,I2866);
DFFARX1 I_25742 (I129285,I2859,I440495,I440521,);
DFFARX1 I_25743 (I440521,I2859,I440495,I440538,);
not I_25744 (I440487,I440538);
not I_25745 (I440560,I440521);
DFFARX1 I_25746 (I129282,I2859,I440495,I440586,);
nand I_25747 (I440594,I440586,I129276);
not I_25748 (I440611,I129276);
not I_25749 (I440628,I129273);
nand I_25750 (I440645,I129267,I129264);
and I_25751 (I440662,I129267,I129264);
not I_25752 (I440679,I129279);
nand I_25753 (I440696,I440679,I440628);
nor I_25754 (I440469,I440696,I440594);
nor I_25755 (I440727,I440611,I440696);
nand I_25756 (I440472,I440662,I440727);
not I_25757 (I440758,I129291);
nor I_25758 (I440775,I440758,I129267);
nor I_25759 (I440792,I440775,I129279);
nor I_25760 (I440809,I440560,I440792);
DFFARX1 I_25761 (I440809,I2859,I440495,I440481,);
not I_25762 (I440840,I440775);
DFFARX1 I_25763 (I440840,I2859,I440495,I440484,);
and I_25764 (I440478,I440586,I440775);
nor I_25765 (I440885,I440758,I129288);
and I_25766 (I440902,I440885,I129264);
or I_25767 (I440919,I440902,I129270);
DFFARX1 I_25768 (I440919,I2859,I440495,I440945,);
nor I_25769 (I440953,I440945,I440679);
DFFARX1 I_25770 (I440953,I2859,I440495,I440466,);
nand I_25771 (I440984,I440945,I440586);
nand I_25772 (I441001,I440679,I440984);
nor I_25773 (I440475,I441001,I440645);
not I_25774 (I441056,I2866);
DFFARX1 I_25775 (I227406,I2859,I441056,I441082,);
DFFARX1 I_25776 (I441082,I2859,I441056,I441099,);
not I_25777 (I441048,I441099);
not I_25778 (I441121,I441082);
DFFARX1 I_25779 (I227403,I2859,I441056,I441147,);
nand I_25780 (I441155,I441147,I227397);
not I_25781 (I441172,I227397);
not I_25782 (I441189,I227409);
nand I_25783 (I441206,I227412,I227391);
and I_25784 (I441223,I227412,I227391);
not I_25785 (I441240,I227388);
nand I_25786 (I441257,I441240,I441189);
nor I_25787 (I441030,I441257,I441155);
nor I_25788 (I441288,I441172,I441257);
nand I_25789 (I441033,I441223,I441288);
not I_25790 (I441319,I227394);
nor I_25791 (I441336,I441319,I227412);
nor I_25792 (I441353,I441336,I227388);
nor I_25793 (I441370,I441121,I441353);
DFFARX1 I_25794 (I441370,I2859,I441056,I441042,);
not I_25795 (I441401,I441336);
DFFARX1 I_25796 (I441401,I2859,I441056,I441045,);
and I_25797 (I441039,I441147,I441336);
nor I_25798 (I441446,I441319,I227388);
and I_25799 (I441463,I441446,I227400);
or I_25800 (I441480,I441463,I227391);
DFFARX1 I_25801 (I441480,I2859,I441056,I441506,);
nor I_25802 (I441514,I441506,I441240);
DFFARX1 I_25803 (I441514,I2859,I441056,I441027,);
nand I_25804 (I441545,I441506,I441147);
nand I_25805 (I441562,I441240,I441545);
nor I_25806 (I441036,I441562,I441206);
not I_25807 (I441617,I2866);
DFFARX1 I_25808 (I169459,I2859,I441617,I441643,);
DFFARX1 I_25809 (I441643,I2859,I441617,I441660,);
not I_25810 (I441609,I441660);
not I_25811 (I441682,I441643);
DFFARX1 I_25812 (I169447,I2859,I441617,I441708,);
nand I_25813 (I441716,I441708,I169453);
not I_25814 (I441733,I169453);
not I_25815 (I441750,I169450);
nand I_25816 (I441767,I169438,I169435);
and I_25817 (I441784,I169438,I169435);
not I_25818 (I441801,I169462);
nand I_25819 (I441818,I441801,I441750);
nor I_25820 (I441591,I441818,I441716);
nor I_25821 (I441849,I441733,I441818);
nand I_25822 (I441594,I441784,I441849);
not I_25823 (I441880,I169435);
nor I_25824 (I441897,I441880,I169438);
nor I_25825 (I441914,I441897,I169462);
nor I_25826 (I441931,I441682,I441914);
DFFARX1 I_25827 (I441931,I2859,I441617,I441603,);
not I_25828 (I441962,I441897);
DFFARX1 I_25829 (I441962,I2859,I441617,I441606,);
and I_25830 (I441600,I441708,I441897);
nor I_25831 (I442007,I441880,I169444);
and I_25832 (I442024,I442007,I169441);
or I_25833 (I442041,I442024,I169456);
DFFARX1 I_25834 (I442041,I2859,I441617,I442067,);
nor I_25835 (I442075,I442067,I441801);
DFFARX1 I_25836 (I442075,I2859,I441617,I441588,);
nand I_25837 (I442106,I442067,I441708);
nand I_25838 (I442123,I441801,I442106);
nor I_25839 (I441597,I442123,I441767);
not I_25840 (I442178,I2866);
DFFARX1 I_25841 (I524585,I2859,I442178,I442204,);
DFFARX1 I_25842 (I442204,I2859,I442178,I442221,);
not I_25843 (I442170,I442221);
not I_25844 (I442243,I442204);
DFFARX1 I_25845 (I524582,I2859,I442178,I442269,);
nand I_25846 (I442277,I442269,I524588);
not I_25847 (I442294,I524588);
not I_25848 (I442311,I524597);
nand I_25849 (I442328,I524591,I524585);
and I_25850 (I442345,I524591,I524585);
not I_25851 (I442362,I524603);
nand I_25852 (I442379,I442362,I442311);
nor I_25853 (I442152,I442379,I442277);
nor I_25854 (I442410,I442294,I442379);
nand I_25855 (I442155,I442345,I442410);
not I_25856 (I442441,I524600);
nor I_25857 (I442458,I442441,I524591);
nor I_25858 (I442475,I442458,I524603);
nor I_25859 (I442492,I442243,I442475);
DFFARX1 I_25860 (I442492,I2859,I442178,I442164,);
not I_25861 (I442523,I442458);
DFFARX1 I_25862 (I442523,I2859,I442178,I442167,);
and I_25863 (I442161,I442269,I442458);
nor I_25864 (I442568,I442441,I524594);
and I_25865 (I442585,I442568,I524606);
or I_25866 (I442602,I442585,I524582);
DFFARX1 I_25867 (I442602,I2859,I442178,I442628,);
nor I_25868 (I442636,I442628,I442362);
DFFARX1 I_25869 (I442636,I2859,I442178,I442149,);
nand I_25870 (I442667,I442628,I442269);
nand I_25871 (I442684,I442362,I442667);
nor I_25872 (I442158,I442684,I442328);
not I_25873 (I442739,I2866);
DFFARX1 I_25874 (I308379,I2859,I442739,I442765,);
DFFARX1 I_25875 (I442765,I2859,I442739,I442782,);
not I_25876 (I442731,I442782);
not I_25877 (I442804,I442765);
DFFARX1 I_25878 (I308391,I2859,I442739,I442830,);
nand I_25879 (I442838,I442830,I308400);
not I_25880 (I442855,I308400);
not I_25881 (I442872,I308382);
nand I_25882 (I442889,I308385,I308376);
and I_25883 (I442906,I308385,I308376);
not I_25884 (I442923,I308394);
nand I_25885 (I442940,I442923,I442872);
nor I_25886 (I442713,I442940,I442838);
nor I_25887 (I442971,I442855,I442940);
nand I_25888 (I442716,I442906,I442971);
not I_25889 (I443002,I308397);
nor I_25890 (I443019,I443002,I308385);
nor I_25891 (I443036,I443019,I308394);
nor I_25892 (I443053,I442804,I443036);
DFFARX1 I_25893 (I443053,I2859,I442739,I442725,);
not I_25894 (I443084,I443019);
DFFARX1 I_25895 (I443084,I2859,I442739,I442728,);
and I_25896 (I442722,I442830,I443019);
nor I_25897 (I443129,I443002,I308376);
and I_25898 (I443146,I443129,I308388);
or I_25899 (I443163,I443146,I308379);
DFFARX1 I_25900 (I443163,I2859,I442739,I443189,);
nor I_25901 (I443197,I443189,I442923);
DFFARX1 I_25902 (I443197,I2859,I442739,I442710,);
nand I_25903 (I443228,I443189,I442830);
nand I_25904 (I443245,I442923,I443228);
nor I_25905 (I442719,I443245,I442889);
not I_25906 (I443300,I2866);
DFFARX1 I_25907 (I335823,I2859,I443300,I443326,);
DFFARX1 I_25908 (I443326,I2859,I443300,I443343,);
not I_25909 (I443292,I443343);
not I_25910 (I443365,I443326);
DFFARX1 I_25911 (I335820,I2859,I443300,I443391,);
nand I_25912 (I443399,I443391,I335835);
not I_25913 (I443416,I335835);
not I_25914 (I443433,I335832);
nand I_25915 (I443450,I335829,I335817);
and I_25916 (I443467,I335829,I335817);
not I_25917 (I443484,I335814);
nand I_25918 (I443501,I443484,I443433);
nor I_25919 (I443274,I443501,I443399);
nor I_25920 (I443532,I443416,I443501);
nand I_25921 (I443277,I443467,I443532);
not I_25922 (I443563,I335820);
nor I_25923 (I443580,I443563,I335829);
nor I_25924 (I443597,I443580,I335814);
nor I_25925 (I443614,I443365,I443597);
DFFARX1 I_25926 (I443614,I2859,I443300,I443286,);
not I_25927 (I443645,I443580);
DFFARX1 I_25928 (I443645,I2859,I443300,I443289,);
and I_25929 (I443283,I443391,I443580);
nor I_25930 (I443690,I443563,I335826);
and I_25931 (I443707,I443690,I335814);
or I_25932 (I443724,I443707,I335817);
DFFARX1 I_25933 (I443724,I2859,I443300,I443750,);
nor I_25934 (I443758,I443750,I443484);
DFFARX1 I_25935 (I443758,I2859,I443300,I443271,);
nand I_25936 (I443789,I443750,I443391);
nand I_25937 (I443806,I443484,I443789);
nor I_25938 (I443280,I443806,I443450);
not I_25939 (I443861,I2866);
DFFARX1 I_25940 (I177075,I2859,I443861,I443887,);
DFFARX1 I_25941 (I443887,I2859,I443861,I443904,);
not I_25942 (I443853,I443904);
not I_25943 (I443926,I443887);
DFFARX1 I_25944 (I177063,I2859,I443861,I443952,);
nand I_25945 (I443960,I443952,I177069);
not I_25946 (I443977,I177069);
not I_25947 (I443994,I177066);
nand I_25948 (I444011,I177054,I177051);
and I_25949 (I444028,I177054,I177051);
not I_25950 (I444045,I177078);
nand I_25951 (I444062,I444045,I443994);
nor I_25952 (I443835,I444062,I443960);
nor I_25953 (I444093,I443977,I444062);
nand I_25954 (I443838,I444028,I444093);
not I_25955 (I444124,I177051);
nor I_25956 (I444141,I444124,I177054);
nor I_25957 (I444158,I444141,I177078);
nor I_25958 (I444175,I443926,I444158);
DFFARX1 I_25959 (I444175,I2859,I443861,I443847,);
not I_25960 (I444206,I444141);
DFFARX1 I_25961 (I444206,I2859,I443861,I443850,);
and I_25962 (I443844,I443952,I444141);
nor I_25963 (I444251,I444124,I177060);
and I_25964 (I444268,I444251,I177057);
or I_25965 (I444285,I444268,I177072);
DFFARX1 I_25966 (I444285,I2859,I443861,I444311,);
nor I_25967 (I444319,I444311,I444045);
DFFARX1 I_25968 (I444319,I2859,I443861,I443832,);
nand I_25969 (I444350,I444311,I443952);
nand I_25970 (I444367,I444045,I444350);
nor I_25971 (I443841,I444367,I444011);
not I_25972 (I444422,I2866);
DFFARX1 I_25973 (I65551,I2859,I444422,I444448,);
DFFARX1 I_25974 (I444448,I2859,I444422,I444465,);
not I_25975 (I444414,I444465);
not I_25976 (I444487,I444448);
DFFARX1 I_25977 (I65566,I2859,I444422,I444513,);
nand I_25978 (I444521,I444513,I65548);
not I_25979 (I444538,I65548);
not I_25980 (I444555,I65557);
nand I_25981 (I444572,I65563,I65554);
and I_25982 (I444589,I65563,I65554);
not I_25983 (I444606,I65551);
nand I_25984 (I444623,I444606,I444555);
nor I_25985 (I444396,I444623,I444521);
nor I_25986 (I444654,I444538,I444623);
nand I_25987 (I444399,I444589,I444654);
not I_25988 (I444685,I65548);
nor I_25989 (I444702,I444685,I65563);
nor I_25990 (I444719,I444702,I65551);
nor I_25991 (I444736,I444487,I444719);
DFFARX1 I_25992 (I444736,I2859,I444422,I444408,);
not I_25993 (I444767,I444702);
DFFARX1 I_25994 (I444767,I2859,I444422,I444411,);
and I_25995 (I444405,I444513,I444702);
nor I_25996 (I444812,I444685,I65572);
and I_25997 (I444829,I444812,I65569);
or I_25998 (I444846,I444829,I65560);
DFFARX1 I_25999 (I444846,I2859,I444422,I444872,);
nor I_26000 (I444880,I444872,I444606);
DFFARX1 I_26001 (I444880,I2859,I444422,I444393,);
nand I_26002 (I444911,I444872,I444513);
nand I_26003 (I444928,I444606,I444911);
nor I_26004 (I444402,I444928,I444572);
not I_26005 (I444983,I2866);
DFFARX1 I_26006 (I553225,I2859,I444983,I445009,);
DFFARX1 I_26007 (I445009,I2859,I444983,I445026,);
not I_26008 (I444975,I445026);
not I_26009 (I445048,I445009);
DFFARX1 I_26010 (I553219,I2859,I444983,I445074,);
nand I_26011 (I445082,I445074,I553210);
not I_26012 (I445099,I553210);
not I_26013 (I445116,I553237);
nand I_26014 (I445133,I553222,I553231);
and I_26015 (I445150,I553222,I553231);
not I_26016 (I445167,I553216);
nand I_26017 (I445184,I445167,I445116);
nor I_26018 (I444957,I445184,I445082);
nor I_26019 (I445215,I445099,I445184);
nand I_26020 (I444960,I445150,I445215);
not I_26021 (I445246,I553234);
nor I_26022 (I445263,I445246,I553222);
nor I_26023 (I445280,I445263,I553216);
nor I_26024 (I445297,I445048,I445280);
DFFARX1 I_26025 (I445297,I2859,I444983,I444969,);
not I_26026 (I445328,I445263);
DFFARX1 I_26027 (I445328,I2859,I444983,I444972,);
and I_26028 (I444966,I445074,I445263);
nor I_26029 (I445373,I445246,I553228);
and I_26030 (I445390,I445373,I553210);
or I_26031 (I445407,I445390,I553213);
DFFARX1 I_26032 (I445407,I2859,I444983,I445433,);
nor I_26033 (I445441,I445433,I445167);
DFFARX1 I_26034 (I445441,I2859,I444983,I444954,);
nand I_26035 (I445472,I445433,I445074);
nand I_26036 (I445489,I445167,I445472);
nor I_26037 (I444963,I445489,I445133);
not I_26038 (I445544,I2866);
DFFARX1 I_26039 (I109259,I2859,I445544,I445570,);
DFFARX1 I_26040 (I445570,I2859,I445544,I445587,);
not I_26041 (I445536,I445587);
not I_26042 (I445609,I445570);
DFFARX1 I_26043 (I109256,I2859,I445544,I445635,);
nand I_26044 (I445643,I445635,I109250);
not I_26045 (I445660,I109250);
not I_26046 (I445677,I109247);
nand I_26047 (I445694,I109241,I109238);
and I_26048 (I445711,I109241,I109238);
not I_26049 (I445728,I109253);
nand I_26050 (I445745,I445728,I445677);
nor I_26051 (I445518,I445745,I445643);
nor I_26052 (I445776,I445660,I445745);
nand I_26053 (I445521,I445711,I445776);
not I_26054 (I445807,I109265);
nor I_26055 (I445824,I445807,I109241);
nor I_26056 (I445841,I445824,I109253);
nor I_26057 (I445858,I445609,I445841);
DFFARX1 I_26058 (I445858,I2859,I445544,I445530,);
not I_26059 (I445889,I445824);
DFFARX1 I_26060 (I445889,I2859,I445544,I445533,);
and I_26061 (I445527,I445635,I445824);
nor I_26062 (I445934,I445807,I109262);
and I_26063 (I445951,I445934,I109238);
or I_26064 (I445968,I445951,I109244);
DFFARX1 I_26065 (I445968,I2859,I445544,I445994,);
nor I_26066 (I446002,I445994,I445728);
DFFARX1 I_26067 (I446002,I2859,I445544,I445515,);
nand I_26068 (I446033,I445994,I445635);
nand I_26069 (I446050,I445728,I446033);
nor I_26070 (I445524,I446050,I445694);
not I_26071 (I446105,I2866);
DFFARX1 I_26072 (I541920,I2859,I446105,I446131,);
DFFARX1 I_26073 (I446131,I2859,I446105,I446148,);
not I_26074 (I446097,I446148);
not I_26075 (I446170,I446131);
DFFARX1 I_26076 (I541914,I2859,I446105,I446196,);
nand I_26077 (I446204,I446196,I541905);
not I_26078 (I446221,I541905);
not I_26079 (I446238,I541932);
nand I_26080 (I446255,I541917,I541926);
and I_26081 (I446272,I541917,I541926);
not I_26082 (I446289,I541911);
nand I_26083 (I446306,I446289,I446238);
nor I_26084 (I446079,I446306,I446204);
nor I_26085 (I446337,I446221,I446306);
nand I_26086 (I446082,I446272,I446337);
not I_26087 (I446368,I541929);
nor I_26088 (I446385,I446368,I541917);
nor I_26089 (I446402,I446385,I541911);
nor I_26090 (I446419,I446170,I446402);
DFFARX1 I_26091 (I446419,I2859,I446105,I446091,);
not I_26092 (I446450,I446385);
DFFARX1 I_26093 (I446450,I2859,I446105,I446094,);
and I_26094 (I446088,I446196,I446385);
nor I_26095 (I446495,I446368,I541923);
and I_26096 (I446512,I446495,I541905);
or I_26097 (I446529,I446512,I541908);
DFFARX1 I_26098 (I446529,I2859,I446105,I446555,);
nor I_26099 (I446563,I446555,I446289);
DFFARX1 I_26100 (I446563,I2859,I446105,I446076,);
nand I_26101 (I446594,I446555,I446196);
nand I_26102 (I446611,I446289,I446594);
nor I_26103 (I446085,I446611,I446255);
not I_26104 (I446666,I2866);
DFFARX1 I_26105 (I21003,I2859,I446666,I446692,);
DFFARX1 I_26106 (I446692,I2859,I446666,I446709,);
not I_26107 (I446658,I446709);
not I_26108 (I446731,I446692);
DFFARX1 I_26109 (I20991,I2859,I446666,I446757,);
nand I_26110 (I446765,I446757,I21006);
not I_26111 (I446782,I21006);
not I_26112 (I446799,I20994);
nand I_26113 (I446816,I21015,I21009);
and I_26114 (I446833,I21015,I21009);
not I_26115 (I446850,I20997);
nand I_26116 (I446867,I446850,I446799);
nor I_26117 (I446640,I446867,I446765);
nor I_26118 (I446898,I446782,I446867);
nand I_26119 (I446643,I446833,I446898);
not I_26120 (I446929,I21000);
nor I_26121 (I446946,I446929,I21015);
nor I_26122 (I446963,I446946,I20997);
nor I_26123 (I446980,I446731,I446963);
DFFARX1 I_26124 (I446980,I2859,I446666,I446652,);
not I_26125 (I447011,I446946);
DFFARX1 I_26126 (I447011,I2859,I446666,I446655,);
and I_26127 (I446649,I446757,I446946);
nor I_26128 (I447056,I446929,I20994);
and I_26129 (I447073,I447056,I20991);
or I_26130 (I447090,I447073,I21012);
DFFARX1 I_26131 (I447090,I2859,I446666,I447116,);
nor I_26132 (I447124,I447116,I446850);
DFFARX1 I_26133 (I447124,I2859,I446666,I446637,);
nand I_26134 (I447155,I447116,I446757);
nand I_26135 (I447172,I446850,I447155);
nor I_26136 (I446646,I447172,I446816);
not I_26137 (I447227,I2866);
DFFARX1 I_26138 (I546085,I2859,I447227,I447253,);
DFFARX1 I_26139 (I447253,I2859,I447227,I447270,);
not I_26140 (I447219,I447270);
not I_26141 (I447292,I447253);
DFFARX1 I_26142 (I546079,I2859,I447227,I447318,);
nand I_26143 (I447326,I447318,I546070);
not I_26144 (I447343,I546070);
not I_26145 (I447360,I546097);
nand I_26146 (I447377,I546082,I546091);
and I_26147 (I447394,I546082,I546091);
not I_26148 (I447411,I546076);
nand I_26149 (I447428,I447411,I447360);
nor I_26150 (I447201,I447428,I447326);
nor I_26151 (I447459,I447343,I447428);
nand I_26152 (I447204,I447394,I447459);
not I_26153 (I447490,I546094);
nor I_26154 (I447507,I447490,I546082);
nor I_26155 (I447524,I447507,I546076);
nor I_26156 (I447541,I447292,I447524);
DFFARX1 I_26157 (I447541,I2859,I447227,I447213,);
not I_26158 (I447572,I447507);
DFFARX1 I_26159 (I447572,I2859,I447227,I447216,);
and I_26160 (I447210,I447318,I447507);
nor I_26161 (I447617,I447490,I546088);
and I_26162 (I447634,I447617,I546070);
or I_26163 (I447651,I447634,I546073);
DFFARX1 I_26164 (I447651,I2859,I447227,I447677,);
nor I_26165 (I447685,I447677,I447411);
DFFARX1 I_26166 (I447685,I2859,I447227,I447198,);
nand I_26167 (I447716,I447677,I447318);
nand I_26168 (I447733,I447411,I447716);
nor I_26169 (I447207,I447733,I447377);
not I_26170 (I447788,I2866);
DFFARX1 I_26171 (I396419,I2859,I447788,I447814,);
DFFARX1 I_26172 (I447814,I2859,I447788,I447831,);
not I_26173 (I447780,I447831);
not I_26174 (I447853,I447814);
DFFARX1 I_26175 (I396446,I2859,I447788,I447879,);
nand I_26176 (I447887,I447879,I396437);
not I_26177 (I447904,I396437);
not I_26178 (I447921,I396419);
nand I_26179 (I447938,I396431,I396434);
and I_26180 (I447955,I396431,I396434);
not I_26181 (I447972,I396443);
nand I_26182 (I447989,I447972,I447921);
nor I_26183 (I447762,I447989,I447887);
nor I_26184 (I448020,I447904,I447989);
nand I_26185 (I447765,I447955,I448020);
not I_26186 (I448051,I396428);
nor I_26187 (I448068,I448051,I396431);
nor I_26188 (I448085,I448068,I396443);
nor I_26189 (I448102,I447853,I448085);
DFFARX1 I_26190 (I448102,I2859,I447788,I447774,);
not I_26191 (I448133,I448068);
DFFARX1 I_26192 (I448133,I2859,I447788,I447777,);
and I_26193 (I447771,I447879,I448068);
nor I_26194 (I448178,I448051,I396422);
and I_26195 (I448195,I448178,I396425);
or I_26196 (I448212,I448195,I396440);
DFFARX1 I_26197 (I448212,I2859,I447788,I448238,);
nor I_26198 (I448246,I448238,I447972);
DFFARX1 I_26199 (I448246,I2859,I447788,I447759,);
nand I_26200 (I448277,I448238,I447879);
nand I_26201 (I448294,I447972,I448277);
nor I_26202 (I447768,I448294,I447938);
not I_26203 (I448352,I2866);
DFFARX1 I_26204 (I2380,I2859,I448352,I448378,);
and I_26205 (I448386,I448378,I1604);
DFFARX1 I_26206 (I448386,I2859,I448352,I448335,);
DFFARX1 I_26207 (I2100,I2859,I448352,I448426,);
not I_26208 (I448434,I1612);
not I_26209 (I448451,I2196);
nand I_26210 (I448468,I448451,I448434);
nor I_26211 (I448323,I448426,I448468);
DFFARX1 I_26212 (I448468,I2859,I448352,I448508,);
not I_26213 (I448344,I448508);
not I_26214 (I448530,I2844);
nand I_26215 (I448547,I448451,I448530);
DFFARX1 I_26216 (I448547,I2859,I448352,I448573,);
not I_26217 (I448581,I448573);
not I_26218 (I448598,I1900);
nand I_26219 (I448615,I448598,I1716);
and I_26220 (I448632,I448434,I448615);
nor I_26221 (I448649,I448547,I448632);
DFFARX1 I_26222 (I448649,I2859,I448352,I448320,);
DFFARX1 I_26223 (I448632,I2859,I448352,I448341,);
nor I_26224 (I448694,I1900,I1588);
nor I_26225 (I448332,I448547,I448694);
or I_26226 (I448725,I1900,I1588);
nor I_26227 (I448742,I2708,I2052);
DFFARX1 I_26228 (I448742,I2859,I448352,I448768,);
not I_26229 (I448776,I448768);
nor I_26230 (I448338,I448776,I448581);
nand I_26231 (I448807,I448776,I448426);
not I_26232 (I448824,I2708);
nand I_26233 (I448841,I448824,I448530);
nand I_26234 (I448858,I448776,I448841);
nand I_26235 (I448329,I448858,I448807);
nand I_26236 (I448326,I448841,I448725);
not I_26237 (I448930,I2866);
DFFARX1 I_26238 (I209147,I2859,I448930,I448956,);
and I_26239 (I448964,I448956,I209162);
DFFARX1 I_26240 (I448964,I2859,I448930,I448913,);
DFFARX1 I_26241 (I209165,I2859,I448930,I449004,);
not I_26242 (I449012,I209159);
not I_26243 (I449029,I209174);
nand I_26244 (I449046,I449029,I449012);
nor I_26245 (I448901,I449004,I449046);
DFFARX1 I_26246 (I449046,I2859,I448930,I449086,);
not I_26247 (I448922,I449086);
not I_26248 (I449108,I209150);
nand I_26249 (I449125,I449029,I449108);
DFFARX1 I_26250 (I449125,I2859,I448930,I449151,);
not I_26251 (I449159,I449151);
not I_26252 (I449176,I209153);
nand I_26253 (I449193,I449176,I209147);
and I_26254 (I449210,I449012,I449193);
nor I_26255 (I449227,I449125,I449210);
DFFARX1 I_26256 (I449227,I2859,I448930,I448898,);
DFFARX1 I_26257 (I449210,I2859,I448930,I448919,);
nor I_26258 (I449272,I209153,I209156);
nor I_26259 (I448910,I449125,I449272);
or I_26260 (I449303,I209153,I209156);
nor I_26261 (I449320,I209171,I209168);
DFFARX1 I_26262 (I449320,I2859,I448930,I449346,);
not I_26263 (I449354,I449346);
nor I_26264 (I448916,I449354,I449159);
nand I_26265 (I449385,I449354,I449004);
not I_26266 (I449402,I209171);
nand I_26267 (I449419,I449402,I449108);
nand I_26268 (I449436,I449354,I449419);
nand I_26269 (I448907,I449436,I449385);
nand I_26270 (I448904,I449419,I449303);
not I_26271 (I449508,I2866);
DFFARX1 I_26272 (I419681,I2859,I449508,I449534,);
and I_26273 (I449542,I449534,I419675);
DFFARX1 I_26274 (I449542,I2859,I449508,I449491,);
DFFARX1 I_26275 (I419693,I2859,I449508,I449582,);
not I_26276 (I449590,I419684);
not I_26277 (I449607,I419696);
nand I_26278 (I449624,I449607,I449590);
nor I_26279 (I449479,I449582,I449624);
DFFARX1 I_26280 (I449624,I2859,I449508,I449664,);
not I_26281 (I449500,I449664);
not I_26282 (I449686,I419702);
nand I_26283 (I449703,I449607,I449686);
DFFARX1 I_26284 (I449703,I2859,I449508,I449729,);
not I_26285 (I449737,I449729);
not I_26286 (I449754,I419678);
nand I_26287 (I449771,I449754,I419699);
and I_26288 (I449788,I449590,I449771);
nor I_26289 (I449805,I449703,I449788);
DFFARX1 I_26290 (I449805,I2859,I449508,I449476,);
DFFARX1 I_26291 (I449788,I2859,I449508,I449497,);
nor I_26292 (I449850,I419678,I419690);
nor I_26293 (I449488,I449703,I449850);
or I_26294 (I449881,I419678,I419690);
nor I_26295 (I449898,I419675,I419687);
DFFARX1 I_26296 (I449898,I2859,I449508,I449924,);
not I_26297 (I449932,I449924);
nor I_26298 (I449494,I449932,I449737);
nand I_26299 (I449963,I449932,I449582);
not I_26300 (I449980,I419675);
nand I_26301 (I449997,I449980,I449686);
nand I_26302 (I450014,I449932,I449997);
nand I_26303 (I449485,I450014,I449963);
nand I_26304 (I449482,I449997,I449881);
not I_26305 (I450086,I2866);
DFFARX1 I_26306 (I308969,I2859,I450086,I450112,);
and I_26307 (I450120,I450112,I308957);
DFFARX1 I_26308 (I450120,I2859,I450086,I450069,);
DFFARX1 I_26309 (I308960,I2859,I450086,I450160,);
not I_26310 (I450168,I308954);
not I_26311 (I450185,I308978);
nand I_26312 (I450202,I450185,I450168);
nor I_26313 (I450057,I450160,I450202);
DFFARX1 I_26314 (I450202,I2859,I450086,I450242,);
not I_26315 (I450078,I450242);
not I_26316 (I450264,I308966);
nand I_26317 (I450281,I450185,I450264);
DFFARX1 I_26318 (I450281,I2859,I450086,I450307,);
not I_26319 (I450315,I450307);
not I_26320 (I450332,I308975);
nand I_26321 (I450349,I450332,I308972);
and I_26322 (I450366,I450168,I450349);
nor I_26323 (I450383,I450281,I450366);
DFFARX1 I_26324 (I450383,I2859,I450086,I450054,);
DFFARX1 I_26325 (I450366,I2859,I450086,I450075,);
nor I_26326 (I450428,I308975,I308963);
nor I_26327 (I450066,I450281,I450428);
or I_26328 (I450459,I308975,I308963);
nor I_26329 (I450476,I308954,I308957);
DFFARX1 I_26330 (I450476,I2859,I450086,I450502,);
not I_26331 (I450510,I450502);
nor I_26332 (I450072,I450510,I450315);
nand I_26333 (I450541,I450510,I450160);
not I_26334 (I450558,I308954);
nand I_26335 (I450575,I450558,I450264);
nand I_26336 (I450592,I450510,I450575);
nand I_26337 (I450063,I450592,I450541);
nand I_26338 (I450060,I450575,I450459);
not I_26339 (I450664,I2866);
DFFARX1 I_26340 (I399655,I2859,I450664,I450690,);
and I_26341 (I450698,I450690,I399649);
DFFARX1 I_26342 (I450698,I2859,I450664,I450647,);
DFFARX1 I_26343 (I399667,I2859,I450664,I450738,);
not I_26344 (I450746,I399658);
not I_26345 (I450763,I399670);
nand I_26346 (I450780,I450763,I450746);
nor I_26347 (I450635,I450738,I450780);
DFFARX1 I_26348 (I450780,I2859,I450664,I450820,);
not I_26349 (I450656,I450820);
not I_26350 (I450842,I399676);
nand I_26351 (I450859,I450763,I450842);
DFFARX1 I_26352 (I450859,I2859,I450664,I450885,);
not I_26353 (I450893,I450885);
not I_26354 (I450910,I399652);
nand I_26355 (I450927,I450910,I399673);
and I_26356 (I450944,I450746,I450927);
nor I_26357 (I450961,I450859,I450944);
DFFARX1 I_26358 (I450961,I2859,I450664,I450632,);
DFFARX1 I_26359 (I450944,I2859,I450664,I450653,);
nor I_26360 (I451006,I399652,I399664);
nor I_26361 (I450644,I450859,I451006);
or I_26362 (I451037,I399652,I399664);
nor I_26363 (I451054,I399649,I399661);
DFFARX1 I_26364 (I451054,I2859,I450664,I451080,);
not I_26365 (I451088,I451080);
nor I_26366 (I450650,I451088,I450893);
nand I_26367 (I451119,I451088,I450738);
not I_26368 (I451136,I399649);
nand I_26369 (I451153,I451136,I450842);
nand I_26370 (I451170,I451088,I451153);
nand I_26371 (I450641,I451170,I451119);
nand I_26372 (I450638,I451153,I451037);
not I_26373 (I451242,I2866);
DFFARX1 I_26374 (I118751,I2859,I451242,I451268,);
and I_26375 (I451276,I451268,I118736);
DFFARX1 I_26376 (I451276,I2859,I451242,I451225,);
DFFARX1 I_26377 (I118742,I2859,I451242,I451316,);
not I_26378 (I451324,I118724);
not I_26379 (I451341,I118745);
nand I_26380 (I451358,I451341,I451324);
nor I_26381 (I451213,I451316,I451358);
DFFARX1 I_26382 (I451358,I2859,I451242,I451398,);
not I_26383 (I451234,I451398);
not I_26384 (I451420,I118748);
nand I_26385 (I451437,I451341,I451420);
DFFARX1 I_26386 (I451437,I2859,I451242,I451463,);
not I_26387 (I451471,I451463);
not I_26388 (I451488,I118739);
nand I_26389 (I451505,I451488,I118727);
and I_26390 (I451522,I451324,I451505);
nor I_26391 (I451539,I451437,I451522);
DFFARX1 I_26392 (I451539,I2859,I451242,I451210,);
DFFARX1 I_26393 (I451522,I2859,I451242,I451231,);
nor I_26394 (I451584,I118739,I118733);
nor I_26395 (I451222,I451437,I451584);
or I_26396 (I451615,I118739,I118733);
nor I_26397 (I451632,I118730,I118724);
DFFARX1 I_26398 (I451632,I2859,I451242,I451658,);
not I_26399 (I451666,I451658);
nor I_26400 (I451228,I451666,I451471);
nand I_26401 (I451697,I451666,I451316);
not I_26402 (I451714,I118730);
nand I_26403 (I451731,I451714,I451420);
nand I_26404 (I451748,I451666,I451731);
nand I_26405 (I451219,I451748,I451697);
nand I_26406 (I451216,I451731,I451615);
not I_26407 (I451820,I2866);
DFFARX1 I_26408 (I259839,I2859,I451820,I451846,);
and I_26409 (I451854,I451846,I259827);
DFFARX1 I_26410 (I451854,I2859,I451820,I451803,);
DFFARX1 I_26411 (I259842,I2859,I451820,I451894,);
not I_26412 (I451902,I259833);
not I_26413 (I451919,I259824);
nand I_26414 (I451936,I451919,I451902);
nor I_26415 (I451791,I451894,I451936);
DFFARX1 I_26416 (I451936,I2859,I451820,I451976,);
not I_26417 (I451812,I451976);
not I_26418 (I451998,I259830);
nand I_26419 (I452015,I451919,I451998);
DFFARX1 I_26420 (I452015,I2859,I451820,I452041,);
not I_26421 (I452049,I452041);
not I_26422 (I452066,I259845);
nand I_26423 (I452083,I452066,I259848);
and I_26424 (I452100,I451902,I452083);
nor I_26425 (I452117,I452015,I452100);
DFFARX1 I_26426 (I452117,I2859,I451820,I451788,);
DFFARX1 I_26427 (I452100,I2859,I451820,I451809,);
nor I_26428 (I452162,I259845,I259824);
nor I_26429 (I451800,I452015,I452162);
or I_26430 (I452193,I259845,I259824);
nor I_26431 (I452210,I259836,I259827);
DFFARX1 I_26432 (I452210,I2859,I451820,I452236,);
not I_26433 (I452244,I452236);
nor I_26434 (I451806,I452244,I452049);
nand I_26435 (I452275,I452244,I451894);
not I_26436 (I452292,I259836);
nand I_26437 (I452309,I452292,I451998);
nand I_26438 (I452326,I452244,I452309);
nand I_26439 (I451797,I452326,I452275);
nand I_26440 (I451794,I452309,I452193);
not I_26441 (I452398,I2866);
DFFARX1 I_26442 (I1676,I2859,I452398,I452424,);
and I_26443 (I452432,I452424,I1932);
DFFARX1 I_26444 (I452432,I2859,I452398,I452381,);
DFFARX1 I_26445 (I1948,I2859,I452398,I452472,);
not I_26446 (I452480,I2524);
not I_26447 (I452497,I1772);
nand I_26448 (I452514,I452497,I452480);
nor I_26449 (I452369,I452472,I452514);
DFFARX1 I_26450 (I452514,I2859,I452398,I452554,);
not I_26451 (I452390,I452554);
not I_26452 (I452576,I2684);
nand I_26453 (I452593,I452497,I452576);
DFFARX1 I_26454 (I452593,I2859,I452398,I452619,);
not I_26455 (I452627,I452619);
not I_26456 (I452644,I2692);
nand I_26457 (I452661,I452644,I2012);
and I_26458 (I452678,I452480,I452661);
nor I_26459 (I452695,I452593,I452678);
DFFARX1 I_26460 (I452695,I2859,I452398,I452366,);
DFFARX1 I_26461 (I452678,I2859,I452398,I452387,);
nor I_26462 (I452740,I2692,I2244);
nor I_26463 (I452378,I452593,I452740);
or I_26464 (I452771,I2692,I2244);
nor I_26465 (I452788,I2436,I2516);
DFFARX1 I_26466 (I452788,I2859,I452398,I452814,);
not I_26467 (I452822,I452814);
nor I_26468 (I452384,I452822,I452627);
nand I_26469 (I452853,I452822,I452472);
not I_26470 (I452870,I2436);
nand I_26471 (I452887,I452870,I452576);
nand I_26472 (I452904,I452822,I452887);
nand I_26473 (I452375,I452904,I452853);
nand I_26474 (I452372,I452887,I452771);
not I_26475 (I452976,I2866);
DFFARX1 I_26476 (I348992,I2859,I452976,I453002,);
and I_26477 (I453010,I453002,I348998);
DFFARX1 I_26478 (I453010,I2859,I452976,I452959,);
DFFARX1 I_26479 (I349004,I2859,I452976,I453050,);
not I_26480 (I453058,I348989);
not I_26481 (I453075,I348989);
nand I_26482 (I453092,I453075,I453058);
nor I_26483 (I452947,I453050,I453092);
DFFARX1 I_26484 (I453092,I2859,I452976,I453132,);
not I_26485 (I452968,I453132);
not I_26486 (I453154,I349007);
nand I_26487 (I453171,I453075,I453154);
DFFARX1 I_26488 (I453171,I2859,I452976,I453197,);
not I_26489 (I453205,I453197);
not I_26490 (I453222,I349001);
nand I_26491 (I453239,I453222,I348992);
and I_26492 (I453256,I453058,I453239);
nor I_26493 (I453273,I453171,I453256);
DFFARX1 I_26494 (I453273,I2859,I452976,I452944,);
DFFARX1 I_26495 (I453256,I2859,I452976,I452965,);
nor I_26496 (I453318,I349001,I349010);
nor I_26497 (I452956,I453171,I453318);
or I_26498 (I453349,I349001,I349010);
nor I_26499 (I453366,I348995,I348995);
DFFARX1 I_26500 (I453366,I2859,I452976,I453392,);
not I_26501 (I453400,I453392);
nor I_26502 (I452962,I453400,I453205);
nand I_26503 (I453431,I453400,I453050);
not I_26504 (I453448,I348995);
nand I_26505 (I453465,I453448,I453154);
nand I_26506 (I453482,I453400,I453465);
nand I_26507 (I452953,I453482,I453431);
nand I_26508 (I452950,I453465,I453349);
not I_26509 (I453554,I2866);
DFFARX1 I_26510 (I141412,I2859,I453554,I453580,);
and I_26511 (I453588,I453580,I141397);
DFFARX1 I_26512 (I453588,I2859,I453554,I453537,);
DFFARX1 I_26513 (I141403,I2859,I453554,I453628,);
not I_26514 (I453636,I141385);
not I_26515 (I453653,I141406);
nand I_26516 (I453670,I453653,I453636);
nor I_26517 (I453525,I453628,I453670);
DFFARX1 I_26518 (I453670,I2859,I453554,I453710,);
not I_26519 (I453546,I453710);
not I_26520 (I453732,I141409);
nand I_26521 (I453749,I453653,I453732);
DFFARX1 I_26522 (I453749,I2859,I453554,I453775,);
not I_26523 (I453783,I453775);
not I_26524 (I453800,I141400);
nand I_26525 (I453817,I453800,I141388);
and I_26526 (I453834,I453636,I453817);
nor I_26527 (I453851,I453749,I453834);
DFFARX1 I_26528 (I453851,I2859,I453554,I453522,);
DFFARX1 I_26529 (I453834,I2859,I453554,I453543,);
nor I_26530 (I453896,I141400,I141394);
nor I_26531 (I453534,I453749,I453896);
or I_26532 (I453927,I141400,I141394);
nor I_26533 (I453944,I141391,I141385);
DFFARX1 I_26534 (I453944,I2859,I453554,I453970,);
not I_26535 (I453978,I453970);
nor I_26536 (I453540,I453978,I453783);
nand I_26537 (I454009,I453978,I453628);
not I_26538 (I454026,I141391);
nand I_26539 (I454043,I454026,I453732);
nand I_26540 (I454060,I453978,I454043);
nand I_26541 (I453531,I454060,I454009);
nand I_26542 (I453528,I454043,I453927);
not I_26543 (I454132,I2866);
DFFARX1 I_26544 (I57905,I2859,I454132,I454158,);
and I_26545 (I454166,I454158,I57881);
DFFARX1 I_26546 (I454166,I2859,I454132,I454115,);
DFFARX1 I_26547 (I57899,I2859,I454132,I454206,);
not I_26548 (I454214,I57887);
not I_26549 (I454231,I57884);
nand I_26550 (I454248,I454231,I454214);
nor I_26551 (I454103,I454206,I454248);
DFFARX1 I_26552 (I454248,I2859,I454132,I454288,);
not I_26553 (I454124,I454288);
not I_26554 (I454310,I57893);
nand I_26555 (I454327,I454231,I454310);
DFFARX1 I_26556 (I454327,I2859,I454132,I454353,);
not I_26557 (I454361,I454353);
not I_26558 (I454378,I57884);
nand I_26559 (I454395,I454378,I57902);
and I_26560 (I454412,I454214,I454395);
nor I_26561 (I454429,I454327,I454412);
DFFARX1 I_26562 (I454429,I2859,I454132,I454100,);
DFFARX1 I_26563 (I454412,I2859,I454132,I454121,);
nor I_26564 (I454474,I57884,I57896);
nor I_26565 (I454112,I454327,I454474);
or I_26566 (I454505,I57884,I57896);
nor I_26567 (I454522,I57890,I57881);
DFFARX1 I_26568 (I454522,I2859,I454132,I454548,);
not I_26569 (I454556,I454548);
nor I_26570 (I454118,I454556,I454361);
nand I_26571 (I454587,I454556,I454206);
not I_26572 (I454604,I57890);
nand I_26573 (I454621,I454604,I454310);
nand I_26574 (I454638,I454556,I454621);
nand I_26575 (I454109,I454638,I454587);
nand I_26576 (I454106,I454621,I454505);
not I_26577 (I454710,I2866);
DFFARX1 I_26578 (I552642,I2859,I454710,I454736,);
and I_26579 (I454744,I454736,I552624);
DFFARX1 I_26580 (I454744,I2859,I454710,I454693,);
DFFARX1 I_26581 (I552615,I2859,I454710,I454784,);
not I_26582 (I454792,I552630);
not I_26583 (I454809,I552618);
nand I_26584 (I454826,I454809,I454792);
nor I_26585 (I454681,I454784,I454826);
DFFARX1 I_26586 (I454826,I2859,I454710,I454866,);
not I_26587 (I454702,I454866);
not I_26588 (I454888,I552627);
nand I_26589 (I454905,I454809,I454888);
DFFARX1 I_26590 (I454905,I2859,I454710,I454931,);
not I_26591 (I454939,I454931);
not I_26592 (I454956,I552636);
nand I_26593 (I454973,I454956,I552615);
and I_26594 (I454990,I454792,I454973);
nor I_26595 (I455007,I454905,I454990);
DFFARX1 I_26596 (I455007,I2859,I454710,I454678,);
DFFARX1 I_26597 (I454990,I2859,I454710,I454699,);
nor I_26598 (I455052,I552636,I552639);
nor I_26599 (I454690,I454905,I455052);
or I_26600 (I455083,I552636,I552639);
nor I_26601 (I455100,I552633,I552621);
DFFARX1 I_26602 (I455100,I2859,I454710,I455126,);
not I_26603 (I455134,I455126);
nor I_26604 (I454696,I455134,I454939);
nand I_26605 (I455165,I455134,I454784);
not I_26606 (I455182,I552633);
nand I_26607 (I455199,I455182,I454888);
nand I_26608 (I455216,I455134,I455199);
nand I_26609 (I454687,I455216,I455165);
nand I_26610 (I454684,I455199,I455083);
not I_26611 (I455288,I2866);
DFFARX1 I_26612 (I104223,I2859,I455288,I455314,);
and I_26613 (I455322,I455314,I104226);
DFFARX1 I_26614 (I455322,I2859,I455288,I455271,);
DFFARX1 I_26615 (I104226,I2859,I455288,I455362,);
not I_26616 (I455370,I104241);
not I_26617 (I455387,I104247);
nand I_26618 (I455404,I455387,I455370);
nor I_26619 (I455259,I455362,I455404);
DFFARX1 I_26620 (I455404,I2859,I455288,I455444,);
not I_26621 (I455280,I455444);
not I_26622 (I455466,I104235);
nand I_26623 (I455483,I455387,I455466);
DFFARX1 I_26624 (I455483,I2859,I455288,I455509,);
not I_26625 (I455517,I455509);
not I_26626 (I455534,I104232);
nand I_26627 (I455551,I455534,I104229);
and I_26628 (I455568,I455370,I455551);
nor I_26629 (I455585,I455483,I455568);
DFFARX1 I_26630 (I455585,I2859,I455288,I455256,);
DFFARX1 I_26631 (I455568,I2859,I455288,I455277,);
nor I_26632 (I455630,I104232,I104223);
nor I_26633 (I455268,I455483,I455630);
or I_26634 (I455661,I104232,I104223);
nor I_26635 (I455678,I104238,I104244);
DFFARX1 I_26636 (I455678,I2859,I455288,I455704,);
not I_26637 (I455712,I455704);
nor I_26638 (I455274,I455712,I455517);
nand I_26639 (I455743,I455712,I455362);
not I_26640 (I455760,I104238);
nand I_26641 (I455777,I455760,I455466);
nand I_26642 (I455794,I455712,I455777);
nand I_26643 (I455265,I455794,I455743);
nand I_26644 (I455262,I455777,I455661);
not I_26645 (I455866,I2866);
DFFARX1 I_26646 (I3479,I2859,I455866,I455892,);
and I_26647 (I455900,I455892,I3485);
DFFARX1 I_26648 (I455900,I2859,I455866,I455849,);
DFFARX1 I_26649 (I3464,I2859,I455866,I455940,);
not I_26650 (I455948,I3470);
not I_26651 (I455965,I3476);
nand I_26652 (I455982,I455965,I455948);
nor I_26653 (I455837,I455940,I455982);
DFFARX1 I_26654 (I455982,I2859,I455866,I456022,);
not I_26655 (I455858,I456022);
not I_26656 (I456044,I3467);
nand I_26657 (I456061,I455965,I456044);
DFFARX1 I_26658 (I456061,I2859,I455866,I456087,);
not I_26659 (I456095,I456087);
not I_26660 (I456112,I3482);
nand I_26661 (I456129,I456112,I3467);
and I_26662 (I456146,I455948,I456129);
nor I_26663 (I456163,I456061,I456146);
DFFARX1 I_26664 (I456163,I2859,I455866,I455834,);
DFFARX1 I_26665 (I456146,I2859,I455866,I455855,);
nor I_26666 (I456208,I3482,I3470);
nor I_26667 (I455846,I456061,I456208);
or I_26668 (I456239,I3482,I3470);
nor I_26669 (I456256,I3473,I3464);
DFFARX1 I_26670 (I456256,I2859,I455866,I456282,);
not I_26671 (I456290,I456282);
nor I_26672 (I455852,I456290,I456095);
nand I_26673 (I456321,I456290,I455940);
not I_26674 (I456338,I3473);
nand I_26675 (I456355,I456338,I456044);
nand I_26676 (I456372,I456290,I456355);
nand I_26677 (I455843,I456372,I456321);
nand I_26678 (I455840,I456355,I456239);
not I_26679 (I456444,I2866);
DFFARX1 I_26680 (I303189,I2859,I456444,I456470,);
and I_26681 (I456478,I456470,I303177);
DFFARX1 I_26682 (I456478,I2859,I456444,I456427,);
DFFARX1 I_26683 (I303180,I2859,I456444,I456518,);
not I_26684 (I456526,I303174);
not I_26685 (I456543,I303198);
nand I_26686 (I456560,I456543,I456526);
nor I_26687 (I456415,I456518,I456560);
DFFARX1 I_26688 (I456560,I2859,I456444,I456600,);
not I_26689 (I456436,I456600);
not I_26690 (I456622,I303186);
nand I_26691 (I456639,I456543,I456622);
DFFARX1 I_26692 (I456639,I2859,I456444,I456665,);
not I_26693 (I456673,I456665);
not I_26694 (I456690,I303195);
nand I_26695 (I456707,I456690,I303192);
and I_26696 (I456724,I456526,I456707);
nor I_26697 (I456741,I456639,I456724);
DFFARX1 I_26698 (I456741,I2859,I456444,I456412,);
DFFARX1 I_26699 (I456724,I2859,I456444,I456433,);
nor I_26700 (I456786,I303195,I303183);
nor I_26701 (I456424,I456639,I456786);
or I_26702 (I456817,I303195,I303183);
nor I_26703 (I456834,I303174,I303177);
DFFARX1 I_26704 (I456834,I2859,I456444,I456860,);
not I_26705 (I456868,I456860);
nor I_26706 (I456430,I456868,I456673);
nand I_26707 (I456899,I456868,I456518);
not I_26708 (I456916,I303174);
nand I_26709 (I456933,I456916,I456622);
nand I_26710 (I456950,I456868,I456933);
nand I_26711 (I456421,I456950,I456899);
nand I_26712 (I456418,I456933,I456817);
not I_26713 (I457022,I2866);
DFFARX1 I_26714 (I120859,I2859,I457022,I457048,);
and I_26715 (I457056,I457048,I120844);
DFFARX1 I_26716 (I457056,I2859,I457022,I457005,);
DFFARX1 I_26717 (I120850,I2859,I457022,I457096,);
not I_26718 (I457104,I120832);
not I_26719 (I457121,I120853);
nand I_26720 (I457138,I457121,I457104);
nor I_26721 (I456993,I457096,I457138);
DFFARX1 I_26722 (I457138,I2859,I457022,I457178,);
not I_26723 (I457014,I457178);
not I_26724 (I457200,I120856);
nand I_26725 (I457217,I457121,I457200);
DFFARX1 I_26726 (I457217,I2859,I457022,I457243,);
not I_26727 (I457251,I457243);
not I_26728 (I457268,I120847);
nand I_26729 (I457285,I457268,I120835);
and I_26730 (I457302,I457104,I457285);
nor I_26731 (I457319,I457217,I457302);
DFFARX1 I_26732 (I457319,I2859,I457022,I456990,);
DFFARX1 I_26733 (I457302,I2859,I457022,I457011,);
nor I_26734 (I457364,I120847,I120841);
nor I_26735 (I457002,I457217,I457364);
or I_26736 (I457395,I120847,I120841);
nor I_26737 (I457412,I120838,I120832);
DFFARX1 I_26738 (I457412,I2859,I457022,I457438,);
not I_26739 (I457446,I457438);
nor I_26740 (I457008,I457446,I457251);
nand I_26741 (I457477,I457446,I457096);
not I_26742 (I457494,I120838);
nand I_26743 (I457511,I457494,I457200);
nand I_26744 (I457528,I457446,I457511);
nand I_26745 (I456999,I457528,I457477);
nand I_26746 (I456996,I457511,I457395);
not I_26747 (I457600,I2866);
DFFARX1 I_26748 (I78043,I2859,I457600,I457626,);
and I_26749 (I457634,I457626,I78046);
DFFARX1 I_26750 (I457634,I2859,I457600,I457583,);
DFFARX1 I_26751 (I78046,I2859,I457600,I457674,);
not I_26752 (I457682,I78061);
not I_26753 (I457699,I78067);
nand I_26754 (I457716,I457699,I457682);
nor I_26755 (I457571,I457674,I457716);
DFFARX1 I_26756 (I457716,I2859,I457600,I457756,);
not I_26757 (I457592,I457756);
not I_26758 (I457778,I78055);
nand I_26759 (I457795,I457699,I457778);
DFFARX1 I_26760 (I457795,I2859,I457600,I457821,);
not I_26761 (I457829,I457821);
not I_26762 (I457846,I78052);
nand I_26763 (I457863,I457846,I78049);
and I_26764 (I457880,I457682,I457863);
nor I_26765 (I457897,I457795,I457880);
DFFARX1 I_26766 (I457897,I2859,I457600,I457568,);
DFFARX1 I_26767 (I457880,I2859,I457600,I457589,);
nor I_26768 (I457942,I78052,I78043);
nor I_26769 (I457580,I457795,I457942);
or I_26770 (I457973,I78052,I78043);
nor I_26771 (I457990,I78058,I78064);
DFFARX1 I_26772 (I457990,I2859,I457600,I458016,);
not I_26773 (I458024,I458016);
nor I_26774 (I457586,I458024,I457829);
nand I_26775 (I458055,I458024,I457674);
not I_26776 (I458072,I78058);
nand I_26777 (I458089,I458072,I457778);
nand I_26778 (I458106,I458024,I458089);
nand I_26779 (I457577,I458106,I458055);
nand I_26780 (I457574,I458089,I457973);
not I_26781 (I458178,I2866);
DFFARX1 I_26782 (I556807,I2859,I458178,I458204,);
and I_26783 (I458212,I458204,I556789);
DFFARX1 I_26784 (I458212,I2859,I458178,I458161,);
DFFARX1 I_26785 (I556780,I2859,I458178,I458252,);
not I_26786 (I458260,I556795);
not I_26787 (I458277,I556783);
nand I_26788 (I458294,I458277,I458260);
nor I_26789 (I458149,I458252,I458294);
DFFARX1 I_26790 (I458294,I2859,I458178,I458334,);
not I_26791 (I458170,I458334);
not I_26792 (I458356,I556792);
nand I_26793 (I458373,I458277,I458356);
DFFARX1 I_26794 (I458373,I2859,I458178,I458399,);
not I_26795 (I458407,I458399);
not I_26796 (I458424,I556801);
nand I_26797 (I458441,I458424,I556780);
and I_26798 (I458458,I458260,I458441);
nor I_26799 (I458475,I458373,I458458);
DFFARX1 I_26800 (I458475,I2859,I458178,I458146,);
DFFARX1 I_26801 (I458458,I2859,I458178,I458167,);
nor I_26802 (I458520,I556801,I556804);
nor I_26803 (I458158,I458373,I458520);
or I_26804 (I458551,I556801,I556804);
nor I_26805 (I458568,I556798,I556786);
DFFARX1 I_26806 (I458568,I2859,I458178,I458594,);
not I_26807 (I458602,I458594);
nor I_26808 (I458164,I458602,I458407);
nand I_26809 (I458633,I458602,I458252);
not I_26810 (I458650,I556798);
nand I_26811 (I458667,I458650,I458356);
nand I_26812 (I458684,I458602,I458667);
nand I_26813 (I458155,I458684,I458633);
nand I_26814 (I458152,I458667,I458551);
not I_26815 (I458756,I2866);
DFFARX1 I_26816 (I1516,I2859,I458756,I458782,);
and I_26817 (I458790,I458782,I1988);
DFFARX1 I_26818 (I458790,I2859,I458756,I458739,);
DFFARX1 I_26819 (I2412,I2859,I458756,I458830,);
not I_26820 (I458838,I1380);
not I_26821 (I458855,I2644);
nand I_26822 (I458872,I458855,I458838);
nor I_26823 (I458727,I458830,I458872);
DFFARX1 I_26824 (I458872,I2859,I458756,I458912,);
not I_26825 (I458748,I458912);
not I_26826 (I458934,I1700);
nand I_26827 (I458951,I458855,I458934);
DFFARX1 I_26828 (I458951,I2859,I458756,I458977,);
not I_26829 (I458985,I458977);
not I_26830 (I459002,I2276);
nand I_26831 (I459019,I459002,I2004);
and I_26832 (I459036,I458838,I459019);
nor I_26833 (I459053,I458951,I459036);
DFFARX1 I_26834 (I459053,I2859,I458756,I458724,);
DFFARX1 I_26835 (I459036,I2859,I458756,I458745,);
nor I_26836 (I459098,I2276,I1396);
nor I_26837 (I458736,I458951,I459098);
or I_26838 (I459129,I2276,I1396);
nor I_26839 (I459146,I1684,I1924);
DFFARX1 I_26840 (I459146,I2859,I458756,I459172,);
not I_26841 (I459180,I459172);
nor I_26842 (I458742,I459180,I458985);
nand I_26843 (I459211,I459180,I458830);
not I_26844 (I459228,I1684);
nand I_26845 (I459245,I459228,I458934);
nand I_26846 (I459262,I459180,I459245);
nand I_26847 (I458733,I459262,I459211);
nand I_26848 (I458730,I459245,I459129);
not I_26849 (I459334,I2866);
DFFARX1 I_26850 (I363221,I2859,I459334,I459360,);
and I_26851 (I459368,I459360,I363227);
DFFARX1 I_26852 (I459368,I2859,I459334,I459317,);
DFFARX1 I_26853 (I363233,I2859,I459334,I459408,);
not I_26854 (I459416,I363218);
not I_26855 (I459433,I363218);
nand I_26856 (I459450,I459433,I459416);
nor I_26857 (I459305,I459408,I459450);
DFFARX1 I_26858 (I459450,I2859,I459334,I459490,);
not I_26859 (I459326,I459490);
not I_26860 (I459512,I363236);
nand I_26861 (I459529,I459433,I459512);
DFFARX1 I_26862 (I459529,I2859,I459334,I459555,);
not I_26863 (I459563,I459555);
not I_26864 (I459580,I363230);
nand I_26865 (I459597,I459580,I363221);
and I_26866 (I459614,I459416,I459597);
nor I_26867 (I459631,I459529,I459614);
DFFARX1 I_26868 (I459631,I2859,I459334,I459302,);
DFFARX1 I_26869 (I459614,I2859,I459334,I459323,);
nor I_26870 (I459676,I363230,I363239);
nor I_26871 (I459314,I459529,I459676);
or I_26872 (I459707,I363230,I363239);
nor I_26873 (I459724,I363224,I363224);
DFFARX1 I_26874 (I459724,I2859,I459334,I459750,);
not I_26875 (I459758,I459750);
nor I_26876 (I459320,I459758,I459563);
nand I_26877 (I459789,I459758,I459408);
not I_26878 (I459806,I363224);
nand I_26879 (I459823,I459806,I459512);
nand I_26880 (I459840,I459758,I459823);
nand I_26881 (I459311,I459840,I459789);
nand I_26882 (I459308,I459823,I459707);
not I_26883 (I459912,I2866);
DFFARX1 I_26884 (I297409,I2859,I459912,I459938,);
and I_26885 (I459946,I459938,I297397);
DFFARX1 I_26886 (I459946,I2859,I459912,I459895,);
DFFARX1 I_26887 (I297400,I2859,I459912,I459986,);
not I_26888 (I459994,I297394);
not I_26889 (I460011,I297418);
nand I_26890 (I460028,I460011,I459994);
nor I_26891 (I459883,I459986,I460028);
DFFARX1 I_26892 (I460028,I2859,I459912,I460068,);
not I_26893 (I459904,I460068);
not I_26894 (I460090,I297406);
nand I_26895 (I460107,I460011,I460090);
DFFARX1 I_26896 (I460107,I2859,I459912,I460133,);
not I_26897 (I460141,I460133);
not I_26898 (I460158,I297415);
nand I_26899 (I460175,I460158,I297412);
and I_26900 (I460192,I459994,I460175);
nor I_26901 (I460209,I460107,I460192);
DFFARX1 I_26902 (I460209,I2859,I459912,I459880,);
DFFARX1 I_26903 (I460192,I2859,I459912,I459901,);
nor I_26904 (I460254,I297415,I297403);
nor I_26905 (I459892,I460107,I460254);
or I_26906 (I460285,I297415,I297403);
nor I_26907 (I460302,I297394,I297397);
DFFARX1 I_26908 (I460302,I2859,I459912,I460328,);
not I_26909 (I460336,I460328);
nor I_26910 (I459898,I460336,I460141);
nand I_26911 (I460367,I460336,I459986);
not I_26912 (I460384,I297394);
nand I_26913 (I460401,I460384,I460090);
nand I_26914 (I460418,I460336,I460401);
nand I_26915 (I459889,I460418,I460367);
nand I_26916 (I459886,I460401,I460285);
not I_26917 (I460490,I2866);
DFFARX1 I_26918 (I371653,I2859,I460490,I460516,);
and I_26919 (I460524,I460516,I371659);
DFFARX1 I_26920 (I460524,I2859,I460490,I460473,);
DFFARX1 I_26921 (I371665,I2859,I460490,I460564,);
not I_26922 (I460572,I371650);
not I_26923 (I460589,I371650);
nand I_26924 (I460606,I460589,I460572);
nor I_26925 (I460461,I460564,I460606);
DFFARX1 I_26926 (I460606,I2859,I460490,I460646,);
not I_26927 (I460482,I460646);
not I_26928 (I460668,I371668);
nand I_26929 (I460685,I460589,I460668);
DFFARX1 I_26930 (I460685,I2859,I460490,I460711,);
not I_26931 (I460719,I460711);
not I_26932 (I460736,I371662);
nand I_26933 (I460753,I460736,I371653);
and I_26934 (I460770,I460572,I460753);
nor I_26935 (I460787,I460685,I460770);
DFFARX1 I_26936 (I460787,I2859,I460490,I460458,);
DFFARX1 I_26937 (I460770,I2859,I460490,I460479,);
nor I_26938 (I460832,I371662,I371671);
nor I_26939 (I460470,I460685,I460832);
or I_26940 (I460863,I371662,I371671);
nor I_26941 (I460880,I371656,I371656);
DFFARX1 I_26942 (I460880,I2859,I460490,I460906,);
not I_26943 (I460914,I460906);
nor I_26944 (I460476,I460914,I460719);
nand I_26945 (I460945,I460914,I460564);
not I_26946 (I460962,I371656);
nand I_26947 (I460979,I460962,I460668);
nand I_26948 (I460996,I460914,I460979);
nand I_26949 (I460467,I460996,I460945);
nand I_26950 (I460464,I460979,I460863);
not I_26951 (I461068,I2866);
DFFARX1 I_26952 (I264463,I2859,I461068,I461094,);
and I_26953 (I461102,I461094,I264451);
DFFARX1 I_26954 (I461102,I2859,I461068,I461051,);
DFFARX1 I_26955 (I264466,I2859,I461068,I461142,);
not I_26956 (I461150,I264457);
not I_26957 (I461167,I264448);
nand I_26958 (I461184,I461167,I461150);
nor I_26959 (I461039,I461142,I461184);
DFFARX1 I_26960 (I461184,I2859,I461068,I461224,);
not I_26961 (I461060,I461224);
not I_26962 (I461246,I264454);
nand I_26963 (I461263,I461167,I461246);
DFFARX1 I_26964 (I461263,I2859,I461068,I461289,);
not I_26965 (I461297,I461289);
not I_26966 (I461314,I264469);
nand I_26967 (I461331,I461314,I264472);
and I_26968 (I461348,I461150,I461331);
nor I_26969 (I461365,I461263,I461348);
DFFARX1 I_26970 (I461365,I2859,I461068,I461036,);
DFFARX1 I_26971 (I461348,I2859,I461068,I461057,);
nor I_26972 (I461410,I264469,I264448);
nor I_26973 (I461048,I461263,I461410);
or I_26974 (I461441,I264469,I264448);
nor I_26975 (I461458,I264460,I264451);
DFFARX1 I_26976 (I461458,I2859,I461068,I461484,);
not I_26977 (I461492,I461484);
nor I_26978 (I461054,I461492,I461297);
nand I_26979 (I461523,I461492,I461142);
not I_26980 (I461540,I264460);
nand I_26981 (I461557,I461540,I461246);
nand I_26982 (I461574,I461492,I461557);
nand I_26983 (I461045,I461574,I461523);
nand I_26984 (I461042,I461557,I461441);
not I_26985 (I461646,I2866);
DFFARX1 I_26986 (I85183,I2859,I461646,I461672,);
and I_26987 (I461680,I461672,I85186);
DFFARX1 I_26988 (I461680,I2859,I461646,I461629,);
DFFARX1 I_26989 (I85186,I2859,I461646,I461720,);
not I_26990 (I461728,I85201);
not I_26991 (I461745,I85207);
nand I_26992 (I461762,I461745,I461728);
nor I_26993 (I461617,I461720,I461762);
DFFARX1 I_26994 (I461762,I2859,I461646,I461802,);
not I_26995 (I461638,I461802);
not I_26996 (I461824,I85195);
nand I_26997 (I461841,I461745,I461824);
DFFARX1 I_26998 (I461841,I2859,I461646,I461867,);
not I_26999 (I461875,I461867);
not I_27000 (I461892,I85192);
nand I_27001 (I461909,I461892,I85189);
and I_27002 (I461926,I461728,I461909);
nor I_27003 (I461943,I461841,I461926);
DFFARX1 I_27004 (I461943,I2859,I461646,I461614,);
DFFARX1 I_27005 (I461926,I2859,I461646,I461635,);
nor I_27006 (I461988,I85192,I85183);
nor I_27007 (I461626,I461841,I461988);
or I_27008 (I462019,I85192,I85183);
nor I_27009 (I462036,I85198,I85204);
DFFARX1 I_27010 (I462036,I2859,I461646,I462062,);
not I_27011 (I462070,I462062);
nor I_27012 (I461632,I462070,I461875);
nand I_27013 (I462101,I462070,I461720);
not I_27014 (I462118,I85198);
nand I_27015 (I462135,I462118,I461824);
nand I_27016 (I462152,I462070,I462135);
nand I_27017 (I461623,I462152,I462101);
nand I_27018 (I461620,I462135,I462019);
not I_27019 (I462224,I2866);
DFFARX1 I_27020 (I356897,I2859,I462224,I462250,);
and I_27021 (I462258,I462250,I356903);
DFFARX1 I_27022 (I462258,I2859,I462224,I462207,);
DFFARX1 I_27023 (I356909,I2859,I462224,I462298,);
not I_27024 (I462306,I356894);
not I_27025 (I462323,I356894);
nand I_27026 (I462340,I462323,I462306);
nor I_27027 (I462195,I462298,I462340);
DFFARX1 I_27028 (I462340,I2859,I462224,I462380,);
not I_27029 (I462216,I462380);
not I_27030 (I462402,I356912);
nand I_27031 (I462419,I462323,I462402);
DFFARX1 I_27032 (I462419,I2859,I462224,I462445,);
not I_27033 (I462453,I462445);
not I_27034 (I462470,I356906);
nand I_27035 (I462487,I462470,I356897);
and I_27036 (I462504,I462306,I462487);
nor I_27037 (I462521,I462419,I462504);
DFFARX1 I_27038 (I462521,I2859,I462224,I462192,);
DFFARX1 I_27039 (I462504,I2859,I462224,I462213,);
nor I_27040 (I462566,I356906,I356915);
nor I_27041 (I462204,I462419,I462566);
or I_27042 (I462597,I356906,I356915);
nor I_27043 (I462614,I356900,I356900);
DFFARX1 I_27044 (I462614,I2859,I462224,I462640,);
not I_27045 (I462648,I462640);
nor I_27046 (I462210,I462648,I462453);
nand I_27047 (I462679,I462648,I462298);
not I_27048 (I462696,I356900);
nand I_27049 (I462713,I462696,I462402);
nand I_27050 (I462730,I462648,I462713);
nand I_27051 (I462201,I462730,I462679);
nand I_27052 (I462198,I462713,I462597);
not I_27053 (I462802,I2866);
DFFARX1 I_27054 (I519503,I2859,I462802,I462828,);
and I_27055 (I462836,I462828,I519497);
DFFARX1 I_27056 (I462836,I2859,I462802,I462785,);
DFFARX1 I_27057 (I519482,I2859,I462802,I462876,);
not I_27058 (I462884,I519488);
not I_27059 (I462901,I519500);
nand I_27060 (I462918,I462901,I462884);
nor I_27061 (I462773,I462876,I462918);
DFFARX1 I_27062 (I462918,I2859,I462802,I462958,);
not I_27063 (I462794,I462958);
not I_27064 (I462980,I519482);
nand I_27065 (I462997,I462901,I462980);
DFFARX1 I_27066 (I462997,I2859,I462802,I463023,);
not I_27067 (I463031,I463023);
not I_27068 (I463048,I519506);
nand I_27069 (I463065,I463048,I519494);
and I_27070 (I463082,I462884,I463065);
nor I_27071 (I463099,I462997,I463082);
DFFARX1 I_27072 (I463099,I2859,I462802,I462770,);
DFFARX1 I_27073 (I463082,I2859,I462802,I462791,);
nor I_27074 (I463144,I519506,I519485);
nor I_27075 (I462782,I462997,I463144);
or I_27076 (I463175,I519506,I519485);
nor I_27077 (I463192,I519491,I519485);
DFFARX1 I_27078 (I463192,I2859,I462802,I463218,);
not I_27079 (I463226,I463218);
nor I_27080 (I462788,I463226,I463031);
nand I_27081 (I463257,I463226,I462876);
not I_27082 (I463274,I519491);
nand I_27083 (I463291,I463274,I462980);
nand I_27084 (I463308,I463226,I463291);
nand I_27085 (I462779,I463308,I463257);
nand I_27086 (I462776,I463291,I463175);
not I_27087 (I463380,I2866);
DFFARX1 I_27088 (I446640,I2859,I463380,I463406,);
and I_27089 (I463414,I463406,I446637);
DFFARX1 I_27090 (I463414,I2859,I463380,I463363,);
DFFARX1 I_27091 (I446643,I2859,I463380,I463454,);
not I_27092 (I463462,I446646);
not I_27093 (I463479,I446640);
nand I_27094 (I463496,I463479,I463462);
nor I_27095 (I463351,I463454,I463496);
DFFARX1 I_27096 (I463496,I2859,I463380,I463536,);
not I_27097 (I463372,I463536);
not I_27098 (I463558,I446655);
nand I_27099 (I463575,I463479,I463558);
DFFARX1 I_27100 (I463575,I2859,I463380,I463601,);
not I_27101 (I463609,I463601);
not I_27102 (I463626,I446652);
nand I_27103 (I463643,I463626,I446658);
and I_27104 (I463660,I463462,I463643);
nor I_27105 (I463677,I463575,I463660);
DFFARX1 I_27106 (I463677,I2859,I463380,I463348,);
DFFARX1 I_27107 (I463660,I2859,I463380,I463369,);
nor I_27108 (I463722,I446652,I446637);
nor I_27109 (I463360,I463575,I463722);
or I_27110 (I463753,I446652,I446637);
nor I_27111 (I463770,I446649,I446643);
DFFARX1 I_27112 (I463770,I2859,I463380,I463796,);
not I_27113 (I463804,I463796);
nor I_27114 (I463366,I463804,I463609);
nand I_27115 (I463835,I463804,I463454);
not I_27116 (I463852,I446649);
nand I_27117 (I463869,I463852,I463558);
nand I_27118 (I463886,I463804,I463869);
nand I_27119 (I463357,I463886,I463835);
nand I_27120 (I463354,I463869,I463753);
not I_27121 (I463958,I2866);
DFFARX1 I_27122 (I155641,I2859,I463958,I463984,);
and I_27123 (I463992,I463984,I155626);
DFFARX1 I_27124 (I463992,I2859,I463958,I463941,);
DFFARX1 I_27125 (I155632,I2859,I463958,I464032,);
not I_27126 (I464040,I155614);
not I_27127 (I464057,I155635);
nand I_27128 (I464074,I464057,I464040);
nor I_27129 (I463929,I464032,I464074);
DFFARX1 I_27130 (I464074,I2859,I463958,I464114,);
not I_27131 (I463950,I464114);
not I_27132 (I464136,I155638);
nand I_27133 (I464153,I464057,I464136);
DFFARX1 I_27134 (I464153,I2859,I463958,I464179,);
not I_27135 (I464187,I464179);
not I_27136 (I464204,I155629);
nand I_27137 (I464221,I464204,I155617);
and I_27138 (I464238,I464040,I464221);
nor I_27139 (I464255,I464153,I464238);
DFFARX1 I_27140 (I464255,I2859,I463958,I463926,);
DFFARX1 I_27141 (I464238,I2859,I463958,I463947,);
nor I_27142 (I464300,I155629,I155623);
nor I_27143 (I463938,I464153,I464300);
or I_27144 (I464331,I155629,I155623);
nor I_27145 (I464348,I155620,I155614);
DFFARX1 I_27146 (I464348,I2859,I463958,I464374,);
not I_27147 (I464382,I464374);
nor I_27148 (I463944,I464382,I464187);
nand I_27149 (I464413,I464382,I464032);
not I_27150 (I464430,I155620);
nand I_27151 (I464447,I464430,I464136);
nand I_27152 (I464464,I464382,I464447);
nand I_27153 (I463935,I464464,I464413);
nand I_27154 (I463932,I464447,I464331);
not I_27155 (I464536,I2866);
DFFARX1 I_27156 (I121913,I2859,I464536,I464562,);
and I_27157 (I464570,I464562,I121898);
DFFARX1 I_27158 (I464570,I2859,I464536,I464519,);
DFFARX1 I_27159 (I121904,I2859,I464536,I464610,);
not I_27160 (I464618,I121886);
not I_27161 (I464635,I121907);
nand I_27162 (I464652,I464635,I464618);
nor I_27163 (I464507,I464610,I464652);
DFFARX1 I_27164 (I464652,I2859,I464536,I464692,);
not I_27165 (I464528,I464692);
not I_27166 (I464714,I121910);
nand I_27167 (I464731,I464635,I464714);
DFFARX1 I_27168 (I464731,I2859,I464536,I464757,);
not I_27169 (I464765,I464757);
not I_27170 (I464782,I121901);
nand I_27171 (I464799,I464782,I121889);
and I_27172 (I464816,I464618,I464799);
nor I_27173 (I464833,I464731,I464816);
DFFARX1 I_27174 (I464833,I2859,I464536,I464504,);
DFFARX1 I_27175 (I464816,I2859,I464536,I464525,);
nor I_27176 (I464878,I121901,I121895);
nor I_27177 (I464516,I464731,I464878);
or I_27178 (I464909,I121901,I121895);
nor I_27179 (I464926,I121892,I121886);
DFFARX1 I_27180 (I464926,I2859,I464536,I464952,);
not I_27181 (I464960,I464952);
nor I_27182 (I464522,I464960,I464765);
nand I_27183 (I464991,I464960,I464610);
not I_27184 (I465008,I121892);
nand I_27185 (I465025,I465008,I464714);
nand I_27186 (I465042,I464960,I465025);
nand I_27187 (I464513,I465042,I464991);
nand I_27188 (I464510,I465025,I464909);
not I_27189 (I465114,I2866);
DFFARX1 I_27190 (I177595,I2859,I465114,I465140,);
and I_27191 (I465148,I465140,I177610);
DFFARX1 I_27192 (I465148,I2859,I465114,I465097,);
DFFARX1 I_27193 (I177613,I2859,I465114,I465188,);
not I_27194 (I465196,I177607);
not I_27195 (I465213,I177622);
nand I_27196 (I465230,I465213,I465196);
nor I_27197 (I465085,I465188,I465230);
DFFARX1 I_27198 (I465230,I2859,I465114,I465270,);
not I_27199 (I465106,I465270);
not I_27200 (I465292,I177598);
nand I_27201 (I465309,I465213,I465292);
DFFARX1 I_27202 (I465309,I2859,I465114,I465335,);
not I_27203 (I465343,I465335);
not I_27204 (I465360,I177601);
nand I_27205 (I465377,I465360,I177595);
and I_27206 (I465394,I465196,I465377);
nor I_27207 (I465411,I465309,I465394);
DFFARX1 I_27208 (I465411,I2859,I465114,I465082,);
DFFARX1 I_27209 (I465394,I2859,I465114,I465103,);
nor I_27210 (I465456,I177601,I177604);
nor I_27211 (I465094,I465309,I465456);
or I_27212 (I465487,I177601,I177604);
nor I_27213 (I465504,I177619,I177616);
DFFARX1 I_27214 (I465504,I2859,I465114,I465530,);
not I_27215 (I465538,I465530);
nor I_27216 (I465100,I465538,I465343);
nand I_27217 (I465569,I465538,I465188);
not I_27218 (I465586,I177619);
nand I_27219 (I465603,I465586,I465292);
nand I_27220 (I465620,I465538,I465603);
nand I_27221 (I465091,I465620,I465569);
nand I_27222 (I465088,I465603,I465487);
not I_27223 (I465692,I2866);
DFFARX1 I_27224 (I161965,I2859,I465692,I465718,);
and I_27225 (I465726,I465718,I161950);
DFFARX1 I_27226 (I465726,I2859,I465692,I465675,);
DFFARX1 I_27227 (I161956,I2859,I465692,I465766,);
not I_27228 (I465774,I161938);
not I_27229 (I465791,I161959);
nand I_27230 (I465808,I465791,I465774);
nor I_27231 (I465663,I465766,I465808);
DFFARX1 I_27232 (I465808,I2859,I465692,I465848,);
not I_27233 (I465684,I465848);
not I_27234 (I465870,I161962);
nand I_27235 (I465887,I465791,I465870);
DFFARX1 I_27236 (I465887,I2859,I465692,I465913,);
not I_27237 (I465921,I465913);
not I_27238 (I465938,I161953);
nand I_27239 (I465955,I465938,I161941);
and I_27240 (I465972,I465774,I465955);
nor I_27241 (I465989,I465887,I465972);
DFFARX1 I_27242 (I465989,I2859,I465692,I465660,);
DFFARX1 I_27243 (I465972,I2859,I465692,I465681,);
nor I_27244 (I466034,I161953,I161947);
nor I_27245 (I465672,I465887,I466034);
or I_27246 (I466065,I161953,I161947);
nor I_27247 (I466082,I161944,I161938);
DFFARX1 I_27248 (I466082,I2859,I465692,I466108,);
not I_27249 (I466116,I466108);
nor I_27250 (I465678,I466116,I465921);
nand I_27251 (I466147,I466116,I465766);
not I_27252 (I466164,I161944);
nand I_27253 (I466181,I466164,I465870);
nand I_27254 (I466198,I466116,I466181);
nand I_27255 (I465669,I466198,I466147);
nand I_27256 (I465666,I466181,I466065);
not I_27257 (I466270,I2866);
DFFARX1 I_27258 (I549072,I2859,I466270,I466296,);
and I_27259 (I466304,I466296,I549054);
DFFARX1 I_27260 (I466304,I2859,I466270,I466253,);
DFFARX1 I_27261 (I549045,I2859,I466270,I466344,);
not I_27262 (I466352,I549060);
not I_27263 (I466369,I549048);
nand I_27264 (I466386,I466369,I466352);
nor I_27265 (I466241,I466344,I466386);
DFFARX1 I_27266 (I466386,I2859,I466270,I466426,);
not I_27267 (I466262,I466426);
not I_27268 (I466448,I549057);
nand I_27269 (I466465,I466369,I466448);
DFFARX1 I_27270 (I466465,I2859,I466270,I466491,);
not I_27271 (I466499,I466491);
not I_27272 (I466516,I549066);
nand I_27273 (I466533,I466516,I549045);
and I_27274 (I466550,I466352,I466533);
nor I_27275 (I466567,I466465,I466550);
DFFARX1 I_27276 (I466567,I2859,I466270,I466238,);
DFFARX1 I_27277 (I466550,I2859,I466270,I466259,);
nor I_27278 (I466612,I549066,I549069);
nor I_27279 (I466250,I466465,I466612);
or I_27280 (I466643,I549066,I549069);
nor I_27281 (I466660,I549063,I549051);
DFFARX1 I_27282 (I466660,I2859,I466270,I466686,);
not I_27283 (I466694,I466686);
nor I_27284 (I466256,I466694,I466499);
nand I_27285 (I466725,I466694,I466344);
not I_27286 (I466742,I549063);
nand I_27287 (I466759,I466742,I466448);
nand I_27288 (I466776,I466694,I466759);
nand I_27289 (I466247,I466776,I466725);
nand I_27290 (I466244,I466759,I466643);
not I_27291 (I466848,I2866);
DFFARX1 I_27292 (I38933,I2859,I466848,I466874,);
and I_27293 (I466882,I466874,I38909);
DFFARX1 I_27294 (I466882,I2859,I466848,I466831,);
DFFARX1 I_27295 (I38927,I2859,I466848,I466922,);
not I_27296 (I466930,I38915);
not I_27297 (I466947,I38912);
nand I_27298 (I466964,I466947,I466930);
nor I_27299 (I466819,I466922,I466964);
DFFARX1 I_27300 (I466964,I2859,I466848,I467004,);
not I_27301 (I466840,I467004);
not I_27302 (I467026,I38921);
nand I_27303 (I467043,I466947,I467026);
DFFARX1 I_27304 (I467043,I2859,I466848,I467069,);
not I_27305 (I467077,I467069);
not I_27306 (I467094,I38912);
nand I_27307 (I467111,I467094,I38930);
and I_27308 (I467128,I466930,I467111);
nor I_27309 (I467145,I467043,I467128);
DFFARX1 I_27310 (I467145,I2859,I466848,I466816,);
DFFARX1 I_27311 (I467128,I2859,I466848,I466837,);
nor I_27312 (I467190,I38912,I38924);
nor I_27313 (I466828,I467043,I467190);
or I_27314 (I467221,I38912,I38924);
nor I_27315 (I467238,I38918,I38909);
DFFARX1 I_27316 (I467238,I2859,I466848,I467264,);
not I_27317 (I467272,I467264);
nor I_27318 (I466834,I467272,I467077);
nand I_27319 (I467303,I467272,I466922);
not I_27320 (I467320,I38918);
nand I_27321 (I467337,I467320,I467026);
nand I_27322 (I467354,I467272,I467337);
nand I_27323 (I466825,I467354,I467303);
nand I_27324 (I466822,I467337,I467221);
not I_27325 (I467426,I2866);
DFFARX1 I_27326 (I518959,I2859,I467426,I467452,);
and I_27327 (I467460,I467452,I518953);
DFFARX1 I_27328 (I467460,I2859,I467426,I467409,);
DFFARX1 I_27329 (I518938,I2859,I467426,I467500,);
not I_27330 (I467508,I518944);
not I_27331 (I467525,I518956);
nand I_27332 (I467542,I467525,I467508);
nor I_27333 (I467397,I467500,I467542);
DFFARX1 I_27334 (I467542,I2859,I467426,I467582,);
not I_27335 (I467418,I467582);
not I_27336 (I467604,I518938);
nand I_27337 (I467621,I467525,I467604);
DFFARX1 I_27338 (I467621,I2859,I467426,I467647,);
not I_27339 (I467655,I467647);
not I_27340 (I467672,I518962);
nand I_27341 (I467689,I467672,I518950);
and I_27342 (I467706,I467508,I467689);
nor I_27343 (I467723,I467621,I467706);
DFFARX1 I_27344 (I467723,I2859,I467426,I467394,);
DFFARX1 I_27345 (I467706,I2859,I467426,I467415,);
nor I_27346 (I467768,I518962,I518941);
nor I_27347 (I467406,I467621,I467768);
or I_27348 (I467799,I518962,I518941);
nor I_27349 (I467816,I518947,I518941);
DFFARX1 I_27350 (I467816,I2859,I467426,I467842,);
not I_27351 (I467850,I467842);
nor I_27352 (I467412,I467850,I467655);
nand I_27353 (I467881,I467850,I467500);
not I_27354 (I467898,I518947);
nand I_27355 (I467915,I467898,I467604);
nand I_27356 (I467932,I467850,I467915);
nand I_27357 (I467403,I467932,I467881);
nand I_27358 (I467400,I467915,I467799);
not I_27359 (I468004,I2866);
DFFARX1 I_27360 (I344249,I2859,I468004,I468030,);
and I_27361 (I468038,I468030,I344255);
DFFARX1 I_27362 (I468038,I2859,I468004,I467987,);
DFFARX1 I_27363 (I344261,I2859,I468004,I468078,);
not I_27364 (I468086,I344246);
not I_27365 (I468103,I344246);
nand I_27366 (I468120,I468103,I468086);
nor I_27367 (I467975,I468078,I468120);
DFFARX1 I_27368 (I468120,I2859,I468004,I468160,);
not I_27369 (I467996,I468160);
not I_27370 (I468182,I344264);
nand I_27371 (I468199,I468103,I468182);
DFFARX1 I_27372 (I468199,I2859,I468004,I468225,);
not I_27373 (I468233,I468225);
not I_27374 (I468250,I344258);
nand I_27375 (I468267,I468250,I344249);
and I_27376 (I468284,I468086,I468267);
nor I_27377 (I468301,I468199,I468284);
DFFARX1 I_27378 (I468301,I2859,I468004,I467972,);
DFFARX1 I_27379 (I468284,I2859,I468004,I467993,);
nor I_27380 (I468346,I344258,I344267);
nor I_27381 (I467984,I468199,I468346);
or I_27382 (I468377,I344258,I344267);
nor I_27383 (I468394,I344252,I344252);
DFFARX1 I_27384 (I468394,I2859,I468004,I468420,);
not I_27385 (I468428,I468420);
nor I_27386 (I467990,I468428,I468233);
nand I_27387 (I468459,I468428,I468078);
not I_27388 (I468476,I344252);
nand I_27389 (I468493,I468476,I468182);
nand I_27390 (I468510,I468428,I468493);
nand I_27391 (I467981,I468510,I468459);
nand I_27392 (I467978,I468493,I468377);
not I_27393 (I468582,I2866);
DFFARX1 I_27394 (I74473,I2859,I468582,I468608,);
and I_27395 (I468616,I468608,I74476);
DFFARX1 I_27396 (I468616,I2859,I468582,I468565,);
DFFARX1 I_27397 (I74476,I2859,I468582,I468656,);
not I_27398 (I468664,I74491);
not I_27399 (I468681,I74497);
nand I_27400 (I468698,I468681,I468664);
nor I_27401 (I468553,I468656,I468698);
DFFARX1 I_27402 (I468698,I2859,I468582,I468738,);
not I_27403 (I468574,I468738);
not I_27404 (I468760,I74485);
nand I_27405 (I468777,I468681,I468760);
DFFARX1 I_27406 (I468777,I2859,I468582,I468803,);
not I_27407 (I468811,I468803);
not I_27408 (I468828,I74482);
nand I_27409 (I468845,I468828,I74479);
and I_27410 (I468862,I468664,I468845);
nor I_27411 (I468879,I468777,I468862);
DFFARX1 I_27412 (I468879,I2859,I468582,I468550,);
DFFARX1 I_27413 (I468862,I2859,I468582,I468571,);
nor I_27414 (I468924,I74482,I74473);
nor I_27415 (I468562,I468777,I468924);
or I_27416 (I468955,I74482,I74473);
nor I_27417 (I468972,I74488,I74494);
DFFARX1 I_27418 (I468972,I2859,I468582,I468998,);
not I_27419 (I469006,I468998);
nor I_27420 (I468568,I469006,I468811);
nand I_27421 (I469037,I469006,I468656);
not I_27422 (I469054,I74488);
nand I_27423 (I469071,I469054,I468760);
nand I_27424 (I469088,I469006,I469071);
nand I_27425 (I468559,I469088,I469037);
nand I_27426 (I468556,I469071,I468955);
not I_27427 (I469160,I2866);
DFFARX1 I_27428 (I210779,I2859,I469160,I469186,);
and I_27429 (I469194,I469186,I210794);
DFFARX1 I_27430 (I469194,I2859,I469160,I469143,);
DFFARX1 I_27431 (I210797,I2859,I469160,I469234,);
not I_27432 (I469242,I210791);
not I_27433 (I469259,I210806);
nand I_27434 (I469276,I469259,I469242);
nor I_27435 (I469131,I469234,I469276);
DFFARX1 I_27436 (I469276,I2859,I469160,I469316,);
not I_27437 (I469152,I469316);
not I_27438 (I469338,I210782);
nand I_27439 (I469355,I469259,I469338);
DFFARX1 I_27440 (I469355,I2859,I469160,I469381,);
not I_27441 (I469389,I469381);
not I_27442 (I469406,I210785);
nand I_27443 (I469423,I469406,I210779);
and I_27444 (I469440,I469242,I469423);
nor I_27445 (I469457,I469355,I469440);
DFFARX1 I_27446 (I469457,I2859,I469160,I469128,);
DFFARX1 I_27447 (I469440,I2859,I469160,I469149,);
nor I_27448 (I469502,I210785,I210788);
nor I_27449 (I469140,I469355,I469502);
or I_27450 (I469533,I210785,I210788);
nor I_27451 (I469550,I210803,I210800);
DFFARX1 I_27452 (I469550,I2859,I469160,I469576,);
not I_27453 (I469584,I469576);
nor I_27454 (I469146,I469584,I469389);
nand I_27455 (I469615,I469584,I469234);
not I_27456 (I469632,I210803);
nand I_27457 (I469649,I469632,I469338);
nand I_27458 (I469666,I469584,I469649);
nand I_27459 (I469137,I469666,I469615);
nand I_27460 (I469134,I469649,I469533);
not I_27461 (I469738,I2866);
DFFARX1 I_27462 (I282959,I2859,I469738,I469764,);
and I_27463 (I469772,I469764,I282947);
DFFARX1 I_27464 (I469772,I2859,I469738,I469721,);
DFFARX1 I_27465 (I282950,I2859,I469738,I469812,);
not I_27466 (I469820,I282944);
not I_27467 (I469837,I282968);
nand I_27468 (I469854,I469837,I469820);
nor I_27469 (I469709,I469812,I469854);
DFFARX1 I_27470 (I469854,I2859,I469738,I469894,);
not I_27471 (I469730,I469894);
not I_27472 (I469916,I282956);
nand I_27473 (I469933,I469837,I469916);
DFFARX1 I_27474 (I469933,I2859,I469738,I469959,);
not I_27475 (I469967,I469959);
not I_27476 (I469984,I282965);
nand I_27477 (I470001,I469984,I282962);
and I_27478 (I470018,I469820,I470001);
nor I_27479 (I470035,I469933,I470018);
DFFARX1 I_27480 (I470035,I2859,I469738,I469706,);
DFFARX1 I_27481 (I470018,I2859,I469738,I469727,);
nor I_27482 (I470080,I282965,I282953);
nor I_27483 (I469718,I469933,I470080);
or I_27484 (I470111,I282965,I282953);
nor I_27485 (I470128,I282944,I282947);
DFFARX1 I_27486 (I470128,I2859,I469738,I470154,);
not I_27487 (I470162,I470154);
nor I_27488 (I469724,I470162,I469967);
nand I_27489 (I470193,I470162,I469812);
not I_27490 (I470210,I282944);
nand I_27491 (I470227,I470210,I469916);
nand I_27492 (I470244,I470162,I470227);
nand I_27493 (I469715,I470244,I470193);
nand I_27494 (I469712,I470227,I470111);
not I_27495 (I470316,I2866);
DFFARX1 I_27496 (I171067,I2859,I470316,I470342,);
and I_27497 (I470350,I470342,I171082);
DFFARX1 I_27498 (I470350,I2859,I470316,I470299,);
DFFARX1 I_27499 (I171085,I2859,I470316,I470390,);
not I_27500 (I470398,I171079);
not I_27501 (I470415,I171094);
nand I_27502 (I470432,I470415,I470398);
nor I_27503 (I470287,I470390,I470432);
DFFARX1 I_27504 (I470432,I2859,I470316,I470472,);
not I_27505 (I470308,I470472);
not I_27506 (I470494,I171070);
nand I_27507 (I470511,I470415,I470494);
DFFARX1 I_27508 (I470511,I2859,I470316,I470537,);
not I_27509 (I470545,I470537);
not I_27510 (I470562,I171073);
nand I_27511 (I470579,I470562,I171067);
and I_27512 (I470596,I470398,I470579);
nor I_27513 (I470613,I470511,I470596);
DFFARX1 I_27514 (I470613,I2859,I470316,I470284,);
DFFARX1 I_27515 (I470596,I2859,I470316,I470305,);
nor I_27516 (I470658,I171073,I171076);
nor I_27517 (I470296,I470511,I470658);
or I_27518 (I470689,I171073,I171076);
nor I_27519 (I470706,I171091,I171088);
DFFARX1 I_27520 (I470706,I2859,I470316,I470732,);
not I_27521 (I470740,I470732);
nor I_27522 (I470302,I470740,I470545);
nand I_27523 (I470771,I470740,I470390);
not I_27524 (I470788,I171091);
nand I_27525 (I470805,I470788,I470494);
nand I_27526 (I470822,I470740,I470805);
nand I_27527 (I470293,I470822,I470771);
nand I_27528 (I470290,I470805,I470689);
not I_27529 (I470894,I2866);
DFFARX1 I_27530 (I545502,I2859,I470894,I470920,);
and I_27531 (I470928,I470920,I545484);
DFFARX1 I_27532 (I470928,I2859,I470894,I470877,);
DFFARX1 I_27533 (I545475,I2859,I470894,I470968,);
not I_27534 (I470976,I545490);
not I_27535 (I470993,I545478);
nand I_27536 (I471010,I470993,I470976);
nor I_27537 (I470865,I470968,I471010);
DFFARX1 I_27538 (I471010,I2859,I470894,I471050,);
not I_27539 (I470886,I471050);
not I_27540 (I471072,I545487);
nand I_27541 (I471089,I470993,I471072);
DFFARX1 I_27542 (I471089,I2859,I470894,I471115,);
not I_27543 (I471123,I471115);
not I_27544 (I471140,I545496);
nand I_27545 (I471157,I471140,I545475);
and I_27546 (I471174,I470976,I471157);
nor I_27547 (I471191,I471089,I471174);
DFFARX1 I_27548 (I471191,I2859,I470894,I470862,);
DFFARX1 I_27549 (I471174,I2859,I470894,I470883,);
nor I_27550 (I471236,I545496,I545499);
nor I_27551 (I470874,I471089,I471236);
or I_27552 (I471267,I545496,I545499);
nor I_27553 (I471284,I545493,I545481);
DFFARX1 I_27554 (I471284,I2859,I470894,I471310,);
not I_27555 (I471318,I471310);
nor I_27556 (I470880,I471318,I471123);
nand I_27557 (I471349,I471318,I470968);
not I_27558 (I471366,I545493);
nand I_27559 (I471383,I471366,I471072);
nand I_27560 (I471400,I471318,I471383);
nand I_27561 (I470871,I471400,I471349);
nand I_27562 (I470868,I471383,I471267);
not I_27563 (I471472,I2866);
DFFARX1 I_27564 (I166715,I2859,I471472,I471498,);
and I_27565 (I471506,I471498,I166730);
DFFARX1 I_27566 (I471506,I2859,I471472,I471455,);
DFFARX1 I_27567 (I166733,I2859,I471472,I471546,);
not I_27568 (I471554,I166727);
not I_27569 (I471571,I166742);
nand I_27570 (I471588,I471571,I471554);
nor I_27571 (I471443,I471546,I471588);
DFFARX1 I_27572 (I471588,I2859,I471472,I471628,);
not I_27573 (I471464,I471628);
not I_27574 (I471650,I166718);
nand I_27575 (I471667,I471571,I471650);
DFFARX1 I_27576 (I471667,I2859,I471472,I471693,);
not I_27577 (I471701,I471693);
not I_27578 (I471718,I166721);
nand I_27579 (I471735,I471718,I166715);
and I_27580 (I471752,I471554,I471735);
nor I_27581 (I471769,I471667,I471752);
DFFARX1 I_27582 (I471769,I2859,I471472,I471440,);
DFFARX1 I_27583 (I471752,I2859,I471472,I471461,);
nor I_27584 (I471814,I166721,I166724);
nor I_27585 (I471452,I471667,I471814);
or I_27586 (I471845,I166721,I166724);
nor I_27587 (I471862,I166739,I166736);
DFFARX1 I_27588 (I471862,I2859,I471472,I471888,);
not I_27589 (I471896,I471888);
nor I_27590 (I471458,I471896,I471701);
nand I_27591 (I471927,I471896,I471546);
not I_27592 (I471944,I166739);
nand I_27593 (I471961,I471944,I471650);
nand I_27594 (I471978,I471896,I471961);
nand I_27595 (I471449,I471978,I471927);
nand I_27596 (I471446,I471961,I471845);
not I_27597 (I472050,I2866);
DFFARX1 I_27598 (I23123,I2859,I472050,I472076,);
and I_27599 (I472084,I472076,I23099);
DFFARX1 I_27600 (I472084,I2859,I472050,I472033,);
DFFARX1 I_27601 (I23117,I2859,I472050,I472124,);
not I_27602 (I472132,I23105);
not I_27603 (I472149,I23102);
nand I_27604 (I472166,I472149,I472132);
nor I_27605 (I472021,I472124,I472166);
DFFARX1 I_27606 (I472166,I2859,I472050,I472206,);
not I_27607 (I472042,I472206);
not I_27608 (I472228,I23111);
nand I_27609 (I472245,I472149,I472228);
DFFARX1 I_27610 (I472245,I2859,I472050,I472271,);
not I_27611 (I472279,I472271);
not I_27612 (I472296,I23102);
nand I_27613 (I472313,I472296,I23120);
and I_27614 (I472330,I472132,I472313);
nor I_27615 (I472347,I472245,I472330);
DFFARX1 I_27616 (I472347,I2859,I472050,I472018,);
DFFARX1 I_27617 (I472330,I2859,I472050,I472039,);
nor I_27618 (I472392,I23102,I23114);
nor I_27619 (I472030,I472245,I472392);
or I_27620 (I472423,I23102,I23114);
nor I_27621 (I472440,I23108,I23099);
DFFARX1 I_27622 (I472440,I2859,I472050,I472466,);
not I_27623 (I472474,I472466);
nor I_27624 (I472036,I472474,I472279);
nand I_27625 (I472505,I472474,I472124);
not I_27626 (I472522,I23108);
nand I_27627 (I472539,I472522,I472228);
nand I_27628 (I472556,I472474,I472539);
nand I_27629 (I472027,I472556,I472505);
nand I_27630 (I472024,I472539,I472423);
not I_27631 (I472628,I2866);
DFFARX1 I_27632 (I1828,I2859,I472628,I472654,);
and I_27633 (I472662,I472654,I2228);
DFFARX1 I_27634 (I472662,I2859,I472628,I472611,);
DFFARX1 I_27635 (I1796,I2859,I472628,I472702,);
not I_27636 (I472710,I2084);
not I_27637 (I472727,I2564);
nand I_27638 (I472744,I472727,I472710);
nor I_27639 (I472599,I472702,I472744);
DFFARX1 I_27640 (I472744,I2859,I472628,I472784,);
not I_27641 (I472620,I472784);
not I_27642 (I472806,I2316);
nand I_27643 (I472823,I472727,I472806);
DFFARX1 I_27644 (I472823,I2859,I472628,I472849,);
not I_27645 (I472857,I472849);
not I_27646 (I472874,I2652);
nand I_27647 (I472891,I472874,I1748);
and I_27648 (I472908,I472710,I472891);
nor I_27649 (I472925,I472823,I472908);
DFFARX1 I_27650 (I472925,I2859,I472628,I472596,);
DFFARX1 I_27651 (I472908,I2859,I472628,I472617,);
nor I_27652 (I472970,I2652,I2180);
nor I_27653 (I472608,I472823,I472970);
or I_27654 (I473001,I2652,I2180);
nor I_27655 (I473018,I1548,I2764);
DFFARX1 I_27656 (I473018,I2859,I472628,I473044,);
not I_27657 (I473052,I473044);
nor I_27658 (I472614,I473052,I472857);
nand I_27659 (I473083,I473052,I472702);
not I_27660 (I473100,I1548);
nand I_27661 (I473117,I473100,I472806);
nand I_27662 (I473134,I473052,I473117);
nand I_27663 (I472605,I473134,I473083);
nand I_27664 (I472602,I473117,I473001);
not I_27665 (I473206,I2866);
DFFARX1 I_27666 (I289317,I2859,I473206,I473232,);
and I_27667 (I473240,I473232,I289305);
DFFARX1 I_27668 (I473240,I2859,I473206,I473189,);
DFFARX1 I_27669 (I289308,I2859,I473206,I473280,);
not I_27670 (I473288,I289302);
not I_27671 (I473305,I289326);
nand I_27672 (I473322,I473305,I473288);
nor I_27673 (I473177,I473280,I473322);
DFFARX1 I_27674 (I473322,I2859,I473206,I473362,);
not I_27675 (I473198,I473362);
not I_27676 (I473384,I289314);
nand I_27677 (I473401,I473305,I473384);
DFFARX1 I_27678 (I473401,I2859,I473206,I473427,);
not I_27679 (I473435,I473427);
not I_27680 (I473452,I289323);
nand I_27681 (I473469,I473452,I289320);
and I_27682 (I473486,I473288,I473469);
nor I_27683 (I473503,I473401,I473486);
DFFARX1 I_27684 (I473503,I2859,I473206,I473174,);
DFFARX1 I_27685 (I473486,I2859,I473206,I473195,);
nor I_27686 (I473548,I289323,I289311);
nor I_27687 (I473186,I473401,I473548);
or I_27688 (I473579,I289323,I289311);
nor I_27689 (I473596,I289302,I289305);
DFFARX1 I_27690 (I473596,I2859,I473206,I473622,);
not I_27691 (I473630,I473622);
nor I_27692 (I473192,I473630,I473435);
nand I_27693 (I473661,I473630,I473280);
not I_27694 (I473678,I289302);
nand I_27695 (I473695,I473678,I473384);
nand I_27696 (I473712,I473630,I473695);
nand I_27697 (I473183,I473712,I473661);
nand I_27698 (I473180,I473695,I473579);
not I_27699 (I473784,I2866);
DFFARX1 I_27700 (I431493,I2859,I473784,I473810,);
and I_27701 (I473818,I473810,I431490);
DFFARX1 I_27702 (I473818,I2859,I473784,I473767,);
DFFARX1 I_27703 (I431496,I2859,I473784,I473858,);
not I_27704 (I473866,I431499);
not I_27705 (I473883,I431493);
nand I_27706 (I473900,I473883,I473866);
nor I_27707 (I473755,I473858,I473900);
DFFARX1 I_27708 (I473900,I2859,I473784,I473940,);
not I_27709 (I473776,I473940);
not I_27710 (I473962,I431508);
nand I_27711 (I473979,I473883,I473962);
DFFARX1 I_27712 (I473979,I2859,I473784,I474005,);
not I_27713 (I474013,I474005);
not I_27714 (I474030,I431505);
nand I_27715 (I474047,I474030,I431511);
and I_27716 (I474064,I473866,I474047);
nor I_27717 (I474081,I473979,I474064);
DFFARX1 I_27718 (I474081,I2859,I473784,I473752,);
DFFARX1 I_27719 (I474064,I2859,I473784,I473773,);
nor I_27720 (I474126,I431505,I431490);
nor I_27721 (I473764,I473979,I474126);
or I_27722 (I474157,I431505,I431490);
nor I_27723 (I474174,I431502,I431496);
DFFARX1 I_27724 (I474174,I2859,I473784,I474200,);
not I_27725 (I474208,I474200);
nor I_27726 (I473770,I474208,I474013);
nand I_27727 (I474239,I474208,I473858);
not I_27728 (I474256,I431502);
nand I_27729 (I474273,I474256,I473962);
nand I_27730 (I474290,I474208,I474273);
nand I_27731 (I473761,I474290,I474239);
nand I_27732 (I473758,I474273,I474157);
not I_27733 (I474362,I2866);
DFFARX1 I_27734 (I270821,I2859,I474362,I474388,);
and I_27735 (I474396,I474388,I270809);
DFFARX1 I_27736 (I474396,I2859,I474362,I474345,);
DFFARX1 I_27737 (I270812,I2859,I474362,I474436,);
not I_27738 (I474444,I270806);
not I_27739 (I474461,I270830);
nand I_27740 (I474478,I474461,I474444);
nor I_27741 (I474333,I474436,I474478);
DFFARX1 I_27742 (I474478,I2859,I474362,I474518,);
not I_27743 (I474354,I474518);
not I_27744 (I474540,I270818);
nand I_27745 (I474557,I474461,I474540);
DFFARX1 I_27746 (I474557,I2859,I474362,I474583,);
not I_27747 (I474591,I474583);
not I_27748 (I474608,I270827);
nand I_27749 (I474625,I474608,I270824);
and I_27750 (I474642,I474444,I474625);
nor I_27751 (I474659,I474557,I474642);
DFFARX1 I_27752 (I474659,I2859,I474362,I474330,);
DFFARX1 I_27753 (I474642,I2859,I474362,I474351,);
nor I_27754 (I474704,I270827,I270815);
nor I_27755 (I474342,I474557,I474704);
or I_27756 (I474735,I270827,I270815);
nor I_27757 (I474752,I270806,I270809);
DFFARX1 I_27758 (I474752,I2859,I474362,I474778,);
not I_27759 (I474786,I474778);
nor I_27760 (I474348,I474786,I474591);
nand I_27761 (I474817,I474786,I474436);
not I_27762 (I474834,I270806);
nand I_27763 (I474851,I474834,I474540);
nand I_27764 (I474868,I474786,I474851);
nand I_27765 (I474339,I474868,I474817);
nand I_27766 (I474336,I474851,I474735);
not I_27767 (I474940,I2866);
DFFARX1 I_27768 (I68523,I2859,I474940,I474966,);
and I_27769 (I474974,I474966,I68526);
DFFARX1 I_27770 (I474974,I2859,I474940,I474923,);
DFFARX1 I_27771 (I68526,I2859,I474940,I475014,);
not I_27772 (I475022,I68541);
not I_27773 (I475039,I68547);
nand I_27774 (I475056,I475039,I475022);
nor I_27775 (I474911,I475014,I475056);
DFFARX1 I_27776 (I475056,I2859,I474940,I475096,);
not I_27777 (I474932,I475096);
not I_27778 (I475118,I68535);
nand I_27779 (I475135,I475039,I475118);
DFFARX1 I_27780 (I475135,I2859,I474940,I475161,);
not I_27781 (I475169,I475161);
not I_27782 (I475186,I68532);
nand I_27783 (I475203,I475186,I68529);
and I_27784 (I475220,I475022,I475203);
nor I_27785 (I475237,I475135,I475220);
DFFARX1 I_27786 (I475237,I2859,I474940,I474908,);
DFFARX1 I_27787 (I475220,I2859,I474940,I474929,);
nor I_27788 (I475282,I68532,I68523);
nor I_27789 (I474920,I475135,I475282);
or I_27790 (I475313,I68532,I68523);
nor I_27791 (I475330,I68538,I68544);
DFFARX1 I_27792 (I475330,I2859,I474940,I475356,);
not I_27793 (I475364,I475356);
nor I_27794 (I474926,I475364,I475169);
nand I_27795 (I475395,I475364,I475014);
not I_27796 (I475412,I68538);
nand I_27797 (I475429,I475412,I475118);
nand I_27798 (I475446,I475364,I475429);
nand I_27799 (I474917,I475446,I475395);
nand I_27800 (I474914,I475429,I475313);
not I_27801 (I475518,I2866);
DFFARX1 I_27802 (I131399,I2859,I475518,I475544,);
and I_27803 (I475552,I475544,I131384);
DFFARX1 I_27804 (I475552,I2859,I475518,I475501,);
DFFARX1 I_27805 (I131390,I2859,I475518,I475592,);
not I_27806 (I475600,I131372);
not I_27807 (I475617,I131393);
nand I_27808 (I475634,I475617,I475600);
nor I_27809 (I475489,I475592,I475634);
DFFARX1 I_27810 (I475634,I2859,I475518,I475674,);
not I_27811 (I475510,I475674);
not I_27812 (I475696,I131396);
nand I_27813 (I475713,I475617,I475696);
DFFARX1 I_27814 (I475713,I2859,I475518,I475739,);
not I_27815 (I475747,I475739);
not I_27816 (I475764,I131387);
nand I_27817 (I475781,I475764,I131375);
and I_27818 (I475798,I475600,I475781);
nor I_27819 (I475815,I475713,I475798);
DFFARX1 I_27820 (I475815,I2859,I475518,I475486,);
DFFARX1 I_27821 (I475798,I2859,I475518,I475507,);
nor I_27822 (I475860,I131387,I131381);
nor I_27823 (I475498,I475713,I475860);
or I_27824 (I475891,I131387,I131381);
nor I_27825 (I475908,I131378,I131372);
DFFARX1 I_27826 (I475908,I2859,I475518,I475934,);
not I_27827 (I475942,I475934);
nor I_27828 (I475504,I475942,I475747);
nand I_27829 (I475973,I475942,I475592);
not I_27830 (I475990,I131378);
nand I_27831 (I476007,I475990,I475696);
nand I_27832 (I476024,I475942,I476007);
nand I_27833 (I475495,I476024,I475973);
nand I_27834 (I475492,I476007,I475891);
not I_27835 (I476096,I2866);
DFFARX1 I_27836 (I63168,I2859,I476096,I476122,);
and I_27837 (I476130,I476122,I63171);
DFFARX1 I_27838 (I476130,I2859,I476096,I476079,);
DFFARX1 I_27839 (I63171,I2859,I476096,I476170,);
not I_27840 (I476178,I63186);
not I_27841 (I476195,I63192);
nand I_27842 (I476212,I476195,I476178);
nor I_27843 (I476067,I476170,I476212);
DFFARX1 I_27844 (I476212,I2859,I476096,I476252,);
not I_27845 (I476088,I476252);
not I_27846 (I476274,I63180);
nand I_27847 (I476291,I476195,I476274);
DFFARX1 I_27848 (I476291,I2859,I476096,I476317,);
not I_27849 (I476325,I476317);
not I_27850 (I476342,I63177);
nand I_27851 (I476359,I476342,I63174);
and I_27852 (I476376,I476178,I476359);
nor I_27853 (I476393,I476291,I476376);
DFFARX1 I_27854 (I476393,I2859,I476096,I476064,);
DFFARX1 I_27855 (I476376,I2859,I476096,I476085,);
nor I_27856 (I476438,I63177,I63168);
nor I_27857 (I476076,I476291,I476438);
or I_27858 (I476469,I63177,I63168);
nor I_27859 (I476486,I63183,I63189);
DFFARX1 I_27860 (I476486,I2859,I476096,I476512,);
not I_27861 (I476520,I476512);
nor I_27862 (I476082,I476520,I476325);
nand I_27863 (I476551,I476520,I476170);
not I_27864 (I476568,I63183);
nand I_27865 (I476585,I476568,I476274);
nand I_27866 (I476602,I476520,I476585);
nand I_27867 (I476073,I476602,I476551);
nand I_27868 (I476070,I476585,I476469);
not I_27869 (I476674,I2866);
DFFARX1 I_27870 (I290473,I2859,I476674,I476700,);
and I_27871 (I476708,I476700,I290461);
DFFARX1 I_27872 (I476708,I2859,I476674,I476657,);
DFFARX1 I_27873 (I290464,I2859,I476674,I476748,);
not I_27874 (I476756,I290458);
not I_27875 (I476773,I290482);
nand I_27876 (I476790,I476773,I476756);
nor I_27877 (I476645,I476748,I476790);
DFFARX1 I_27878 (I476790,I2859,I476674,I476830,);
not I_27879 (I476666,I476830);
not I_27880 (I476852,I290470);
nand I_27881 (I476869,I476773,I476852);
DFFARX1 I_27882 (I476869,I2859,I476674,I476895,);
not I_27883 (I476903,I476895);
not I_27884 (I476920,I290479);
nand I_27885 (I476937,I476920,I290476);
and I_27886 (I476954,I476756,I476937);
nor I_27887 (I476971,I476869,I476954);
DFFARX1 I_27888 (I476971,I2859,I476674,I476642,);
DFFARX1 I_27889 (I476954,I2859,I476674,I476663,);
nor I_27890 (I477016,I290479,I290467);
nor I_27891 (I476654,I476869,I477016);
or I_27892 (I477047,I290479,I290467);
nor I_27893 (I477064,I290458,I290461);
DFFARX1 I_27894 (I477064,I2859,I476674,I477090,);
not I_27895 (I477098,I477090);
nor I_27896 (I476660,I477098,I476903);
nand I_27897 (I477129,I477098,I476748);
not I_27898 (I477146,I290458);
nand I_27899 (I477163,I477146,I476852);
nand I_27900 (I477180,I477098,I477163);
nand I_27901 (I476651,I477180,I477129);
nand I_27902 (I476648,I477163,I477047);
not I_27903 (I477252,I2866);
DFFARX1 I_27904 (I346357,I2859,I477252,I477278,);
and I_27905 (I477286,I477278,I346363);
DFFARX1 I_27906 (I477286,I2859,I477252,I477235,);
DFFARX1 I_27907 (I346369,I2859,I477252,I477326,);
not I_27908 (I477334,I346354);
not I_27909 (I477351,I346354);
nand I_27910 (I477368,I477351,I477334);
nor I_27911 (I477223,I477326,I477368);
DFFARX1 I_27912 (I477368,I2859,I477252,I477408,);
not I_27913 (I477244,I477408);
not I_27914 (I477430,I346372);
nand I_27915 (I477447,I477351,I477430);
DFFARX1 I_27916 (I477447,I2859,I477252,I477473,);
not I_27917 (I477481,I477473);
not I_27918 (I477498,I346366);
nand I_27919 (I477515,I477498,I346357);
and I_27920 (I477532,I477334,I477515);
nor I_27921 (I477549,I477447,I477532);
DFFARX1 I_27922 (I477549,I2859,I477252,I477220,);
DFFARX1 I_27923 (I477532,I2859,I477252,I477241,);
nor I_27924 (I477594,I346366,I346375);
nor I_27925 (I477232,I477447,I477594);
or I_27926 (I477625,I346366,I346375);
nor I_27927 (I477642,I346360,I346360);
DFFARX1 I_27928 (I477642,I2859,I477252,I477668,);
not I_27929 (I477676,I477668);
nor I_27930 (I477238,I477676,I477481);
nand I_27931 (I477707,I477676,I477326);
not I_27932 (I477724,I346360);
nand I_27933 (I477741,I477724,I477430);
nand I_27934 (I477758,I477676,I477741);
nand I_27935 (I477229,I477758,I477707);
nand I_27936 (I477226,I477741,I477625);
not I_27937 (I477830,I2866);
DFFARX1 I_27938 (I330355,I2859,I477830,I477856,);
and I_27939 (I477864,I477856,I330343);
DFFARX1 I_27940 (I477864,I2859,I477830,I477813,);
DFFARX1 I_27941 (I330346,I2859,I477830,I477904,);
not I_27942 (I477912,I330340);
not I_27943 (I477929,I330364);
nand I_27944 (I477946,I477929,I477912);
nor I_27945 (I477801,I477904,I477946);
DFFARX1 I_27946 (I477946,I2859,I477830,I477986,);
not I_27947 (I477822,I477986);
not I_27948 (I478008,I330352);
nand I_27949 (I478025,I477929,I478008);
DFFARX1 I_27950 (I478025,I2859,I477830,I478051,);
not I_27951 (I478059,I478051);
not I_27952 (I478076,I330361);
nand I_27953 (I478093,I478076,I330358);
and I_27954 (I478110,I477912,I478093);
nor I_27955 (I478127,I478025,I478110);
DFFARX1 I_27956 (I478127,I2859,I477830,I477798,);
DFFARX1 I_27957 (I478110,I2859,I477830,I477819,);
nor I_27958 (I478172,I330361,I330349);
nor I_27959 (I477810,I478025,I478172);
or I_27960 (I478203,I330361,I330349);
nor I_27961 (I478220,I330340,I330343);
DFFARX1 I_27962 (I478220,I2859,I477830,I478246,);
not I_27963 (I478254,I478246);
nor I_27964 (I477816,I478254,I478059);
nand I_27965 (I478285,I478254,I477904);
not I_27966 (I478302,I330340);
nand I_27967 (I478319,I478302,I478008);
nand I_27968 (I478336,I478254,I478319);
nand I_27969 (I477807,I478336,I478285);
nand I_27970 (I477804,I478319,I478203);
not I_27971 (I478408,I2866);
DFFARX1 I_27972 (I324575,I2859,I478408,I478434,);
and I_27973 (I478442,I478434,I324563);
DFFARX1 I_27974 (I478442,I2859,I478408,I478391,);
DFFARX1 I_27975 (I324566,I2859,I478408,I478482,);
not I_27976 (I478490,I324560);
not I_27977 (I478507,I324584);
nand I_27978 (I478524,I478507,I478490);
nor I_27979 (I478379,I478482,I478524);
DFFARX1 I_27980 (I478524,I2859,I478408,I478564,);
not I_27981 (I478400,I478564);
not I_27982 (I478586,I324572);
nand I_27983 (I478603,I478507,I478586);
DFFARX1 I_27984 (I478603,I2859,I478408,I478629,);
not I_27985 (I478637,I478629);
not I_27986 (I478654,I324581);
nand I_27987 (I478671,I478654,I324578);
and I_27988 (I478688,I478490,I478671);
nor I_27989 (I478705,I478603,I478688);
DFFARX1 I_27990 (I478705,I2859,I478408,I478376,);
DFFARX1 I_27991 (I478688,I2859,I478408,I478397,);
nor I_27992 (I478750,I324581,I324569);
nor I_27993 (I478388,I478603,I478750);
or I_27994 (I478781,I324581,I324569);
nor I_27995 (I478798,I324560,I324563);
DFFARX1 I_27996 (I478798,I2859,I478408,I478824,);
not I_27997 (I478832,I478824);
nor I_27998 (I478394,I478832,I478637);
nand I_27999 (I478863,I478832,I478482);
not I_28000 (I478880,I324560);
nand I_28001 (I478897,I478880,I478586);
nand I_28002 (I478914,I478832,I478897);
nand I_28003 (I478385,I478914,I478863);
nand I_28004 (I478382,I478897,I478781);
not I_28005 (I478986,I2866);
DFFARX1 I_28006 (I273711,I2859,I478986,I479012,);
and I_28007 (I479020,I479012,I273699);
DFFARX1 I_28008 (I479020,I2859,I478986,I478969,);
DFFARX1 I_28009 (I273702,I2859,I478986,I479060,);
not I_28010 (I479068,I273696);
not I_28011 (I479085,I273720);
nand I_28012 (I479102,I479085,I479068);
nor I_28013 (I478957,I479060,I479102);
DFFARX1 I_28014 (I479102,I2859,I478986,I479142,);
not I_28015 (I478978,I479142);
not I_28016 (I479164,I273708);
nand I_28017 (I479181,I479085,I479164);
DFFARX1 I_28018 (I479181,I2859,I478986,I479207,);
not I_28019 (I479215,I479207);
not I_28020 (I479232,I273717);
nand I_28021 (I479249,I479232,I273714);
and I_28022 (I479266,I479068,I479249);
nor I_28023 (I479283,I479181,I479266);
DFFARX1 I_28024 (I479283,I2859,I478986,I478954,);
DFFARX1 I_28025 (I479266,I2859,I478986,I478975,);
nor I_28026 (I479328,I273717,I273705);
nor I_28027 (I478966,I479181,I479328);
or I_28028 (I479359,I273717,I273705);
nor I_28029 (I479376,I273696,I273699);
DFFARX1 I_28030 (I479376,I2859,I478986,I479402,);
not I_28031 (I479410,I479402);
nor I_28032 (I478972,I479410,I479215);
nand I_28033 (I479441,I479410,I479060);
not I_28034 (I479458,I273696);
nand I_28035 (I479475,I479458,I479164);
nand I_28036 (I479492,I479410,I479475);
nand I_28037 (I478963,I479492,I479441);
nand I_28038 (I478960,I479475,I479359);
not I_28039 (I479564,I2866);
DFFARX1 I_28040 (I311281,I2859,I479564,I479590,);
and I_28041 (I479598,I479590,I311269);
DFFARX1 I_28042 (I479598,I2859,I479564,I479547,);
DFFARX1 I_28043 (I311272,I2859,I479564,I479638,);
not I_28044 (I479646,I311266);
not I_28045 (I479663,I311290);
nand I_28046 (I479680,I479663,I479646);
nor I_28047 (I479535,I479638,I479680);
DFFARX1 I_28048 (I479680,I2859,I479564,I479720,);
not I_28049 (I479556,I479720);
not I_28050 (I479742,I311278);
nand I_28051 (I479759,I479663,I479742);
DFFARX1 I_28052 (I479759,I2859,I479564,I479785,);
not I_28053 (I479793,I479785);
not I_28054 (I479810,I311287);
nand I_28055 (I479827,I479810,I311284);
and I_28056 (I479844,I479646,I479827);
nor I_28057 (I479861,I479759,I479844);
DFFARX1 I_28058 (I479861,I2859,I479564,I479532,);
DFFARX1 I_28059 (I479844,I2859,I479564,I479553,);
nor I_28060 (I479906,I311287,I311275);
nor I_28061 (I479544,I479759,I479906);
or I_28062 (I479937,I311287,I311275);
nor I_28063 (I479954,I311266,I311269);
DFFARX1 I_28064 (I479954,I2859,I479564,I479980,);
not I_28065 (I479988,I479980);
nor I_28066 (I479550,I479988,I479793);
nand I_28067 (I480019,I479988,I479638);
not I_28068 (I480036,I311266);
nand I_28069 (I480053,I480036,I479742);
nand I_28070 (I480070,I479988,I480053);
nand I_28071 (I479541,I480070,I480019);
nand I_28072 (I479538,I480053,I479937);
not I_28073 (I480142,I2866);
DFFARX1 I_28074 (I168347,I2859,I480142,I480168,);
and I_28075 (I480176,I480168,I168362);
DFFARX1 I_28076 (I480176,I2859,I480142,I480125,);
DFFARX1 I_28077 (I168365,I2859,I480142,I480216,);
not I_28078 (I480224,I168359);
not I_28079 (I480241,I168374);
nand I_28080 (I480258,I480241,I480224);
nor I_28081 (I480113,I480216,I480258);
DFFARX1 I_28082 (I480258,I2859,I480142,I480298,);
not I_28083 (I480134,I480298);
not I_28084 (I480320,I168350);
nand I_28085 (I480337,I480241,I480320);
DFFARX1 I_28086 (I480337,I2859,I480142,I480363,);
not I_28087 (I480371,I480363);
not I_28088 (I480388,I168353);
nand I_28089 (I480405,I480388,I168347);
and I_28090 (I480422,I480224,I480405);
nor I_28091 (I480439,I480337,I480422);
DFFARX1 I_28092 (I480439,I2859,I480142,I480110,);
DFFARX1 I_28093 (I480422,I2859,I480142,I480131,);
nor I_28094 (I480484,I168353,I168356);
nor I_28095 (I480122,I480337,I480484);
or I_28096 (I480515,I168353,I168356);
nor I_28097 (I480532,I168371,I168368);
DFFARX1 I_28098 (I480532,I2859,I480142,I480558,);
not I_28099 (I480566,I480558);
nor I_28100 (I480128,I480566,I480371);
nand I_28101 (I480597,I480566,I480216);
not I_28102 (I480614,I168371);
nand I_28103 (I480631,I480614,I480320);
nand I_28104 (I480648,I480566,I480631);
nand I_28105 (I480119,I480648,I480597);
nand I_28106 (I480116,I480631,I480515);
not I_28107 (I480720,I2866);
DFFARX1 I_28108 (I140885,I2859,I480720,I480746,);
and I_28109 (I480754,I480746,I140870);
DFFARX1 I_28110 (I480754,I2859,I480720,I480703,);
DFFARX1 I_28111 (I140876,I2859,I480720,I480794,);
not I_28112 (I480802,I140858);
not I_28113 (I480819,I140879);
nand I_28114 (I480836,I480819,I480802);
nor I_28115 (I480691,I480794,I480836);
DFFARX1 I_28116 (I480836,I2859,I480720,I480876,);
not I_28117 (I480712,I480876);
not I_28118 (I480898,I140882);
nand I_28119 (I480915,I480819,I480898);
DFFARX1 I_28120 (I480915,I2859,I480720,I480941,);
not I_28121 (I480949,I480941);
not I_28122 (I480966,I140873);
nand I_28123 (I480983,I480966,I140861);
and I_28124 (I481000,I480802,I480983);
nor I_28125 (I481017,I480915,I481000);
DFFARX1 I_28126 (I481017,I2859,I480720,I480688,);
DFFARX1 I_28127 (I481000,I2859,I480720,I480709,);
nor I_28128 (I481062,I140873,I140867);
nor I_28129 (I480700,I480915,I481062);
or I_28130 (I481093,I140873,I140867);
nor I_28131 (I481110,I140864,I140858);
DFFARX1 I_28132 (I481110,I2859,I480720,I481136,);
not I_28133 (I481144,I481136);
nor I_28134 (I480706,I481144,I480949);
nand I_28135 (I481175,I481144,I480794);
not I_28136 (I481192,I140864);
nand I_28137 (I481209,I481192,I480898);
nand I_28138 (I481226,I481144,I481209);
nand I_28139 (I480697,I481226,I481175);
nand I_28140 (I480694,I481209,I481093);
not I_28141 (I481298,I2866);
DFFARX1 I_28142 (I416451,I2859,I481298,I481324,);
and I_28143 (I481332,I481324,I416445);
DFFARX1 I_28144 (I481332,I2859,I481298,I481281,);
DFFARX1 I_28145 (I416463,I2859,I481298,I481372,);
not I_28146 (I481380,I416454);
not I_28147 (I481397,I416466);
nand I_28148 (I481414,I481397,I481380);
nor I_28149 (I481269,I481372,I481414);
DFFARX1 I_28150 (I481414,I2859,I481298,I481454,);
not I_28151 (I481290,I481454);
not I_28152 (I481476,I416472);
nand I_28153 (I481493,I481397,I481476);
DFFARX1 I_28154 (I481493,I2859,I481298,I481519,);
not I_28155 (I481527,I481519);
not I_28156 (I481544,I416448);
nand I_28157 (I481561,I481544,I416469);
and I_28158 (I481578,I481380,I481561);
nor I_28159 (I481595,I481493,I481578);
DFFARX1 I_28160 (I481595,I2859,I481298,I481266,);
DFFARX1 I_28161 (I481578,I2859,I481298,I481287,);
nor I_28162 (I481640,I416448,I416460);
nor I_28163 (I481278,I481493,I481640);
or I_28164 (I481671,I416448,I416460);
nor I_28165 (I481688,I416445,I416457);
DFFARX1 I_28166 (I481688,I2859,I481298,I481714,);
not I_28167 (I481722,I481714);
nor I_28168 (I481284,I481722,I481527);
nand I_28169 (I481753,I481722,I481372);
not I_28170 (I481770,I416445);
nand I_28171 (I481787,I481770,I481476);
nand I_28172 (I481804,I481722,I481787);
nand I_28173 (I481275,I481804,I481753);
nand I_28174 (I481272,I481787,I481671);
not I_28175 (I481876,I2866);
DFFARX1 I_28176 (I438225,I2859,I481876,I481902,);
and I_28177 (I481910,I481902,I438222);
DFFARX1 I_28178 (I481910,I2859,I481876,I481859,);
DFFARX1 I_28179 (I438228,I2859,I481876,I481950,);
not I_28180 (I481958,I438231);
not I_28181 (I481975,I438225);
nand I_28182 (I481992,I481975,I481958);
nor I_28183 (I481847,I481950,I481992);
DFFARX1 I_28184 (I481992,I2859,I481876,I482032,);
not I_28185 (I481868,I482032);
not I_28186 (I482054,I438240);
nand I_28187 (I482071,I481975,I482054);
DFFARX1 I_28188 (I482071,I2859,I481876,I482097,);
not I_28189 (I482105,I482097);
not I_28190 (I482122,I438237);
nand I_28191 (I482139,I482122,I438243);
and I_28192 (I482156,I481958,I482139);
nor I_28193 (I482173,I482071,I482156);
DFFARX1 I_28194 (I482173,I2859,I481876,I481844,);
DFFARX1 I_28195 (I482156,I2859,I481876,I481865,);
nor I_28196 (I482218,I438237,I438222);
nor I_28197 (I481856,I482071,I482218);
or I_28198 (I482249,I438237,I438222);
nor I_28199 (I482266,I438234,I438228);
DFFARX1 I_28200 (I482266,I2859,I481876,I482292,);
not I_28201 (I482300,I482292);
nor I_28202 (I481862,I482300,I482105);
nand I_28203 (I482331,I482300,I481950);
not I_28204 (I482348,I438234);
nand I_28205 (I482365,I482348,I482054);
nand I_28206 (I482382,I482300,I482365);
nand I_28207 (I481853,I482382,I482331);
nand I_28208 (I481850,I482365,I482249);
not I_28209 (I482454,I2866);
DFFARX1 I_28210 (I386735,I2859,I482454,I482480,);
and I_28211 (I482488,I482480,I386729);
DFFARX1 I_28212 (I482488,I2859,I482454,I482437,);
DFFARX1 I_28213 (I386747,I2859,I482454,I482528,);
not I_28214 (I482536,I386738);
not I_28215 (I482553,I386750);
nand I_28216 (I482570,I482553,I482536);
nor I_28217 (I482425,I482528,I482570);
DFFARX1 I_28218 (I482570,I2859,I482454,I482610,);
not I_28219 (I482446,I482610);
not I_28220 (I482632,I386756);
nand I_28221 (I482649,I482553,I482632);
DFFARX1 I_28222 (I482649,I2859,I482454,I482675,);
not I_28223 (I482683,I482675);
not I_28224 (I482700,I386732);
nand I_28225 (I482717,I482700,I386753);
and I_28226 (I482734,I482536,I482717);
nor I_28227 (I482751,I482649,I482734);
DFFARX1 I_28228 (I482751,I2859,I482454,I482422,);
DFFARX1 I_28229 (I482734,I2859,I482454,I482443,);
nor I_28230 (I482796,I386732,I386744);
nor I_28231 (I482434,I482649,I482796);
or I_28232 (I482827,I386732,I386744);
nor I_28233 (I482844,I386729,I386741);
DFFARX1 I_28234 (I482844,I2859,I482454,I482870,);
not I_28235 (I482878,I482870);
nor I_28236 (I482440,I482878,I482683);
nand I_28237 (I482909,I482878,I482528);
not I_28238 (I482926,I386729);
nand I_28239 (I482943,I482926,I482632);
nand I_28240 (I482960,I482878,I482943);
nand I_28241 (I482431,I482960,I482909);
nand I_28242 (I482428,I482943,I482827);
not I_28243 (I483032,I2866);
DFFARX1 I_28244 (I540147,I2859,I483032,I483058,);
and I_28245 (I483066,I483058,I540129);
DFFARX1 I_28246 (I483066,I2859,I483032,I483015,);
DFFARX1 I_28247 (I540120,I2859,I483032,I483106,);
not I_28248 (I483114,I540135);
not I_28249 (I483131,I540123);
nand I_28250 (I483148,I483131,I483114);
nor I_28251 (I483003,I483106,I483148);
DFFARX1 I_28252 (I483148,I2859,I483032,I483188,);
not I_28253 (I483024,I483188);
not I_28254 (I483210,I540132);
nand I_28255 (I483227,I483131,I483210);
DFFARX1 I_28256 (I483227,I2859,I483032,I483253,);
not I_28257 (I483261,I483253);
not I_28258 (I483278,I540141);
nand I_28259 (I483295,I483278,I540120);
and I_28260 (I483312,I483114,I483295);
nor I_28261 (I483329,I483227,I483312);
DFFARX1 I_28262 (I483329,I2859,I483032,I483000,);
DFFARX1 I_28263 (I483312,I2859,I483032,I483021,);
nor I_28264 (I483374,I540141,I540144);
nor I_28265 (I483012,I483227,I483374);
or I_28266 (I483405,I540141,I540144);
nor I_28267 (I483422,I540138,I540126);
DFFARX1 I_28268 (I483422,I2859,I483032,I483448,);
not I_28269 (I483456,I483448);
nor I_28270 (I483018,I483456,I483261);
nand I_28271 (I483487,I483456,I483106);
not I_28272 (I483504,I540138);
nand I_28273 (I483521,I483504,I483210);
nand I_28274 (I483538,I483456,I483521);
nand I_28275 (I483009,I483538,I483487);
nand I_28276 (I483006,I483521,I483405);
not I_28277 (I483610,I2866);
DFFARX1 I_28278 (I382859,I2859,I483610,I483636,);
and I_28279 (I483644,I483636,I382853);
DFFARX1 I_28280 (I483644,I2859,I483610,I483593,);
DFFARX1 I_28281 (I382871,I2859,I483610,I483684,);
not I_28282 (I483692,I382862);
not I_28283 (I483709,I382874);
nand I_28284 (I483726,I483709,I483692);
nor I_28285 (I483581,I483684,I483726);
DFFARX1 I_28286 (I483726,I2859,I483610,I483766,);
not I_28287 (I483602,I483766);
not I_28288 (I483788,I382880);
nand I_28289 (I483805,I483709,I483788);
DFFARX1 I_28290 (I483805,I2859,I483610,I483831,);
not I_28291 (I483839,I483831);
not I_28292 (I483856,I382856);
nand I_28293 (I483873,I483856,I382877);
and I_28294 (I483890,I483692,I483873);
nor I_28295 (I483907,I483805,I483890);
DFFARX1 I_28296 (I483907,I2859,I483610,I483578,);
DFFARX1 I_28297 (I483890,I2859,I483610,I483599,);
nor I_28298 (I483952,I382856,I382868);
nor I_28299 (I483590,I483805,I483952);
or I_28300 (I483983,I382856,I382868);
nor I_28301 (I484000,I382853,I382865);
DFFARX1 I_28302 (I484000,I2859,I483610,I484026,);
not I_28303 (I484034,I484026);
nor I_28304 (I483596,I484034,I483839);
nand I_28305 (I484065,I484034,I483684);
not I_28306 (I484082,I382853);
nand I_28307 (I484099,I484082,I483788);
nand I_28308 (I484116,I484034,I484099);
nand I_28309 (I483587,I484116,I484065);
nand I_28310 (I483584,I484099,I483983);
not I_28311 (I484188,I2866);
DFFARX1 I_28312 (I303767,I2859,I484188,I484214,);
and I_28313 (I484222,I484214,I303755);
DFFARX1 I_28314 (I484222,I2859,I484188,I484171,);
DFFARX1 I_28315 (I303758,I2859,I484188,I484262,);
not I_28316 (I484270,I303752);
not I_28317 (I484287,I303776);
nand I_28318 (I484304,I484287,I484270);
nor I_28319 (I484159,I484262,I484304);
DFFARX1 I_28320 (I484304,I2859,I484188,I484344,);
not I_28321 (I484180,I484344);
not I_28322 (I484366,I303764);
nand I_28323 (I484383,I484287,I484366);
DFFARX1 I_28324 (I484383,I2859,I484188,I484409,);
not I_28325 (I484417,I484409);
not I_28326 (I484434,I303773);
nand I_28327 (I484451,I484434,I303770);
and I_28328 (I484468,I484270,I484451);
nor I_28329 (I484485,I484383,I484468);
DFFARX1 I_28330 (I484485,I2859,I484188,I484156,);
DFFARX1 I_28331 (I484468,I2859,I484188,I484177,);
nor I_28332 (I484530,I303773,I303761);
nor I_28333 (I484168,I484383,I484530);
or I_28334 (I484561,I303773,I303761);
nor I_28335 (I484578,I303752,I303755);
DFFARX1 I_28336 (I484578,I2859,I484188,I484604,);
not I_28337 (I484612,I484604);
nor I_28338 (I484174,I484612,I484417);
nand I_28339 (I484643,I484612,I484262);
not I_28340 (I484660,I303752);
nand I_28341 (I484677,I484660,I484366);
nand I_28342 (I484694,I484612,I484677);
nand I_28343 (I484165,I484694,I484643);
nand I_28344 (I484162,I484677,I484561);
not I_28345 (I484766,I2866);
DFFARX1 I_28346 (I189019,I2859,I484766,I484792,);
and I_28347 (I484800,I484792,I189034);
DFFARX1 I_28348 (I484800,I2859,I484766,I484749,);
DFFARX1 I_28349 (I189037,I2859,I484766,I484840,);
not I_28350 (I484848,I189031);
not I_28351 (I484865,I189046);
nand I_28352 (I484882,I484865,I484848);
nor I_28353 (I484737,I484840,I484882);
DFFARX1 I_28354 (I484882,I2859,I484766,I484922,);
not I_28355 (I484758,I484922);
not I_28356 (I484944,I189022);
nand I_28357 (I484961,I484865,I484944);
DFFARX1 I_28358 (I484961,I2859,I484766,I484987,);
not I_28359 (I484995,I484987);
not I_28360 (I485012,I189025);
nand I_28361 (I485029,I485012,I189019);
and I_28362 (I485046,I484848,I485029);
nor I_28363 (I485063,I484961,I485046);
DFFARX1 I_28364 (I485063,I2859,I484766,I484734,);
DFFARX1 I_28365 (I485046,I2859,I484766,I484755,);
nor I_28366 (I485108,I189025,I189028);
nor I_28367 (I484746,I484961,I485108);
or I_28368 (I485139,I189025,I189028);
nor I_28369 (I485156,I189043,I189040);
DFFARX1 I_28370 (I485156,I2859,I484766,I485182,);
not I_28371 (I485190,I485182);
nor I_28372 (I484752,I485190,I484995);
nand I_28373 (I485221,I485190,I484840);
not I_28374 (I485238,I189043);
nand I_28375 (I485255,I485238,I484944);
nand I_28376 (I485272,I485190,I485255);
nand I_28377 (I484743,I485272,I485221);
nand I_28378 (I484740,I485255,I485139);
not I_28379 (I485344,I2866);
DFFARX1 I_28380 (I422911,I2859,I485344,I485370,);
and I_28381 (I485378,I485370,I422905);
DFFARX1 I_28382 (I485378,I2859,I485344,I485327,);
DFFARX1 I_28383 (I422923,I2859,I485344,I485418,);
not I_28384 (I485426,I422914);
not I_28385 (I485443,I422926);
nand I_28386 (I485460,I485443,I485426);
nor I_28387 (I485315,I485418,I485460);
DFFARX1 I_28388 (I485460,I2859,I485344,I485500,);
not I_28389 (I485336,I485500);
not I_28390 (I485522,I422932);
nand I_28391 (I485539,I485443,I485522);
DFFARX1 I_28392 (I485539,I2859,I485344,I485565,);
not I_28393 (I485573,I485565);
not I_28394 (I485590,I422908);
nand I_28395 (I485607,I485590,I422929);
and I_28396 (I485624,I485426,I485607);
nor I_28397 (I485641,I485539,I485624);
DFFARX1 I_28398 (I485641,I2859,I485344,I485312,);
DFFARX1 I_28399 (I485624,I2859,I485344,I485333,);
nor I_28400 (I485686,I422908,I422920);
nor I_28401 (I485324,I485539,I485686);
or I_28402 (I485717,I422908,I422920);
nor I_28403 (I485734,I422905,I422917);
DFFARX1 I_28404 (I485734,I2859,I485344,I485760,);
not I_28405 (I485768,I485760);
nor I_28406 (I485330,I485768,I485573);
nand I_28407 (I485799,I485768,I485418);
not I_28408 (I485816,I422905);
nand I_28409 (I485833,I485816,I485522);
nand I_28410 (I485850,I485768,I485833);
nand I_28411 (I485321,I485850,I485799);
nand I_28412 (I485318,I485833,I485717);
not I_28413 (I485922,I2866);
DFFARX1 I_28414 (I4654,I2859,I485922,I485948,);
and I_28415 (I485956,I485948,I4657);
DFFARX1 I_28416 (I485956,I2859,I485922,I485905,);
DFFARX1 I_28417 (I4657,I2859,I485922,I485996,);
not I_28418 (I486004,I4660);
not I_28419 (I486021,I4675);
nand I_28420 (I486038,I486021,I486004);
nor I_28421 (I485893,I485996,I486038);
DFFARX1 I_28422 (I486038,I2859,I485922,I486078,);
not I_28423 (I485914,I486078);
not I_28424 (I486100,I4669);
nand I_28425 (I486117,I486021,I486100);
DFFARX1 I_28426 (I486117,I2859,I485922,I486143,);
not I_28427 (I486151,I486143);
not I_28428 (I486168,I4672);
nand I_28429 (I486185,I486168,I4654);
and I_28430 (I486202,I486004,I486185);
nor I_28431 (I486219,I486117,I486202);
DFFARX1 I_28432 (I486219,I2859,I485922,I485890,);
DFFARX1 I_28433 (I486202,I2859,I485922,I485911,);
nor I_28434 (I486264,I4672,I4666);
nor I_28435 (I485902,I486117,I486264);
or I_28436 (I486295,I4672,I4666);
nor I_28437 (I486312,I4663,I4678);
DFFARX1 I_28438 (I486312,I2859,I485922,I486338,);
not I_28439 (I486346,I486338);
nor I_28440 (I485908,I486346,I486151);
nand I_28441 (I486377,I486346,I485996);
not I_28442 (I486394,I4663);
nand I_28443 (I486411,I486394,I486100);
nand I_28444 (I486428,I486346,I486411);
nand I_28445 (I485899,I486428,I486377);
nand I_28446 (I485896,I486411,I486295);
not I_28447 (I486500,I2866);
DFFARX1 I_28448 (I293941,I2859,I486500,I486526,);
and I_28449 (I486534,I486526,I293929);
DFFARX1 I_28450 (I486534,I2859,I486500,I486483,);
DFFARX1 I_28451 (I293932,I2859,I486500,I486574,);
not I_28452 (I486582,I293926);
not I_28453 (I486599,I293950);
nand I_28454 (I486616,I486599,I486582);
nor I_28455 (I486471,I486574,I486616);
DFFARX1 I_28456 (I486616,I2859,I486500,I486656,);
not I_28457 (I486492,I486656);
not I_28458 (I486678,I293938);
nand I_28459 (I486695,I486599,I486678);
DFFARX1 I_28460 (I486695,I2859,I486500,I486721,);
not I_28461 (I486729,I486721);
not I_28462 (I486746,I293947);
nand I_28463 (I486763,I486746,I293944);
and I_28464 (I486780,I486582,I486763);
nor I_28465 (I486797,I486695,I486780);
DFFARX1 I_28466 (I486797,I2859,I486500,I486468,);
DFFARX1 I_28467 (I486780,I2859,I486500,I486489,);
nor I_28468 (I486842,I293947,I293935);
nor I_28469 (I486480,I486695,I486842);
or I_28470 (I486873,I293947,I293935);
nor I_28471 (I486890,I293926,I293929);
DFFARX1 I_28472 (I486890,I2859,I486500,I486916,);
not I_28473 (I486924,I486916);
nor I_28474 (I486486,I486924,I486729);
nand I_28475 (I486955,I486924,I486574);
not I_28476 (I486972,I293926);
nand I_28477 (I486989,I486972,I486678);
nand I_28478 (I487006,I486924,I486989);
nand I_28479 (I486477,I487006,I486955);
nand I_28480 (I486474,I486989,I486873);
not I_28481 (I487078,I2866);
DFFARX1 I_28482 (I10451,I2859,I487078,I487104,);
and I_28483 (I487112,I487104,I10454);
DFFARX1 I_28484 (I487112,I2859,I487078,I487061,);
DFFARX1 I_28485 (I10454,I2859,I487078,I487152,);
not I_28486 (I487160,I10457);
not I_28487 (I487177,I10472);
nand I_28488 (I487194,I487177,I487160);
nor I_28489 (I487049,I487152,I487194);
DFFARX1 I_28490 (I487194,I2859,I487078,I487234,);
not I_28491 (I487070,I487234);
not I_28492 (I487256,I10466);
nand I_28493 (I487273,I487177,I487256);
DFFARX1 I_28494 (I487273,I2859,I487078,I487299,);
not I_28495 (I487307,I487299);
not I_28496 (I487324,I10469);
nand I_28497 (I487341,I487324,I10451);
and I_28498 (I487358,I487160,I487341);
nor I_28499 (I487375,I487273,I487358);
DFFARX1 I_28500 (I487375,I2859,I487078,I487046,);
DFFARX1 I_28501 (I487358,I2859,I487078,I487067,);
nor I_28502 (I487420,I10469,I10463);
nor I_28503 (I487058,I487273,I487420);
or I_28504 (I487451,I10469,I10463);
nor I_28505 (I487468,I10460,I10475);
DFFARX1 I_28506 (I487468,I2859,I487078,I487494,);
not I_28507 (I487502,I487494);
nor I_28508 (I487064,I487502,I487307);
nand I_28509 (I487533,I487502,I487152);
not I_28510 (I487550,I10460);
nand I_28511 (I487567,I487550,I487256);
nand I_28512 (I487584,I487502,I487567);
nand I_28513 (I487055,I487584,I487533);
nand I_28514 (I487052,I487567,I487451);
not I_28515 (I487656,I2866);
DFFARX1 I_28516 (I205339,I2859,I487656,I487682,);
and I_28517 (I487690,I487682,I205354);
DFFARX1 I_28518 (I487690,I2859,I487656,I487639,);
DFFARX1 I_28519 (I205357,I2859,I487656,I487730,);
not I_28520 (I487738,I205351);
not I_28521 (I487755,I205366);
nand I_28522 (I487772,I487755,I487738);
nor I_28523 (I487627,I487730,I487772);
DFFARX1 I_28524 (I487772,I2859,I487656,I487812,);
not I_28525 (I487648,I487812);
not I_28526 (I487834,I205342);
nand I_28527 (I487851,I487755,I487834);
DFFARX1 I_28528 (I487851,I2859,I487656,I487877,);
not I_28529 (I487885,I487877);
not I_28530 (I487902,I205345);
nand I_28531 (I487919,I487902,I205339);
and I_28532 (I487936,I487738,I487919);
nor I_28533 (I487953,I487851,I487936);
DFFARX1 I_28534 (I487953,I2859,I487656,I487624,);
DFFARX1 I_28535 (I487936,I2859,I487656,I487645,);
nor I_28536 (I487998,I205345,I205348);
nor I_28537 (I487636,I487851,I487998);
or I_28538 (I488029,I205345,I205348);
nor I_28539 (I488046,I205363,I205360);
DFFARX1 I_28540 (I488046,I2859,I487656,I488072,);
not I_28541 (I488080,I488072);
nor I_28542 (I487642,I488080,I487885);
nand I_28543 (I488111,I488080,I487730);
not I_28544 (I488128,I205363);
nand I_28545 (I488145,I488128,I487834);
nand I_28546 (I488162,I488080,I488145);
nand I_28547 (I487633,I488162,I488111);
nand I_28548 (I487630,I488145,I488029);
not I_28549 (I488234,I2866);
DFFARX1 I_28550 (I137723,I2859,I488234,I488260,);
and I_28551 (I488268,I488260,I137708);
DFFARX1 I_28552 (I488268,I2859,I488234,I488217,);
DFFARX1 I_28553 (I137714,I2859,I488234,I488308,);
not I_28554 (I488316,I137696);
not I_28555 (I488333,I137717);
nand I_28556 (I488350,I488333,I488316);
nor I_28557 (I488205,I488308,I488350);
DFFARX1 I_28558 (I488350,I2859,I488234,I488390,);
not I_28559 (I488226,I488390);
not I_28560 (I488412,I137720);
nand I_28561 (I488429,I488333,I488412);
DFFARX1 I_28562 (I488429,I2859,I488234,I488455,);
not I_28563 (I488463,I488455);
not I_28564 (I488480,I137711);
nand I_28565 (I488497,I488480,I137699);
and I_28566 (I488514,I488316,I488497);
nor I_28567 (I488531,I488429,I488514);
DFFARX1 I_28568 (I488531,I2859,I488234,I488202,);
DFFARX1 I_28569 (I488514,I2859,I488234,I488223,);
nor I_28570 (I488576,I137711,I137705);
nor I_28571 (I488214,I488429,I488576);
or I_28572 (I488607,I137711,I137705);
nor I_28573 (I488624,I137702,I137696);
DFFARX1 I_28574 (I488624,I2859,I488234,I488650,);
not I_28575 (I488658,I488650);
nor I_28576 (I488220,I488658,I488463);
nand I_28577 (I488689,I488658,I488308);
not I_28578 (I488706,I137702);
nand I_28579 (I488723,I488706,I488412);
nand I_28580 (I488740,I488658,I488723);
nand I_28581 (I488211,I488740,I488689);
nand I_28582 (I488208,I488723,I488607);
not I_28583 (I488812,I2866);
DFFARX1 I_28584 (I44203,I2859,I488812,I488838,);
and I_28585 (I488846,I488838,I44179);
DFFARX1 I_28586 (I488846,I2859,I488812,I488795,);
DFFARX1 I_28587 (I44197,I2859,I488812,I488886,);
not I_28588 (I488894,I44185);
not I_28589 (I488911,I44182);
nand I_28590 (I488928,I488911,I488894);
nor I_28591 (I488783,I488886,I488928);
DFFARX1 I_28592 (I488928,I2859,I488812,I488968,);
not I_28593 (I488804,I488968);
not I_28594 (I488990,I44191);
nand I_28595 (I489007,I488911,I488990);
DFFARX1 I_28596 (I489007,I2859,I488812,I489033,);
not I_28597 (I489041,I489033);
not I_28598 (I489058,I44182);
nand I_28599 (I489075,I489058,I44200);
and I_28600 (I489092,I488894,I489075);
nor I_28601 (I489109,I489007,I489092);
DFFARX1 I_28602 (I489109,I2859,I488812,I488780,);
DFFARX1 I_28603 (I489092,I2859,I488812,I488801,);
nor I_28604 (I489154,I44182,I44194);
nor I_28605 (I488792,I489007,I489154);
or I_28606 (I489185,I44182,I44194);
nor I_28607 (I489202,I44188,I44179);
DFFARX1 I_28608 (I489202,I2859,I488812,I489228,);
not I_28609 (I489236,I489228);
nor I_28610 (I488798,I489236,I489041);
nand I_28611 (I489267,I489236,I488886);
not I_28612 (I489284,I44188);
nand I_28613 (I489301,I489284,I488990);
nand I_28614 (I489318,I489236,I489301);
nand I_28615 (I488789,I489318,I489267);
nand I_28616 (I488786,I489301,I489185);
not I_28617 (I489390,I2866);
DFFARX1 I_28618 (I320529,I2859,I489390,I489416,);
and I_28619 (I489424,I489416,I320517);
DFFARX1 I_28620 (I489424,I2859,I489390,I489373,);
DFFARX1 I_28621 (I320520,I2859,I489390,I489464,);
not I_28622 (I489472,I320514);
not I_28623 (I489489,I320538);
nand I_28624 (I489506,I489489,I489472);
nor I_28625 (I489361,I489464,I489506);
DFFARX1 I_28626 (I489506,I2859,I489390,I489546,);
not I_28627 (I489382,I489546);
not I_28628 (I489568,I320526);
nand I_28629 (I489585,I489489,I489568);
DFFARX1 I_28630 (I489585,I2859,I489390,I489611,);
not I_28631 (I489619,I489611);
not I_28632 (I489636,I320535);
nand I_28633 (I489653,I489636,I320532);
and I_28634 (I489670,I489472,I489653);
nor I_28635 (I489687,I489585,I489670);
DFFARX1 I_28636 (I489687,I2859,I489390,I489358,);
DFFARX1 I_28637 (I489670,I2859,I489390,I489379,);
nor I_28638 (I489732,I320535,I320523);
nor I_28639 (I489370,I489585,I489732);
or I_28640 (I489763,I320535,I320523);
nor I_28641 (I489780,I320514,I320517);
DFFARX1 I_28642 (I489780,I2859,I489390,I489806,);
not I_28643 (I489814,I489806);
nor I_28644 (I489376,I489814,I489619);
nand I_28645 (I489845,I489814,I489464);
not I_28646 (I489862,I320514);
nand I_28647 (I489879,I489862,I489568);
nand I_28648 (I489896,I489814,I489879);
nand I_28649 (I489367,I489896,I489845);
nand I_28650 (I489364,I489879,I489763);
not I_28651 (I489968,I2866);
DFFARX1 I_28652 (I35771,I2859,I489968,I489994,);
and I_28653 (I490002,I489994,I35747);
DFFARX1 I_28654 (I490002,I2859,I489968,I489951,);
DFFARX1 I_28655 (I35765,I2859,I489968,I490042,);
not I_28656 (I490050,I35753);
not I_28657 (I490067,I35750);
nand I_28658 (I490084,I490067,I490050);
nor I_28659 (I489939,I490042,I490084);
DFFARX1 I_28660 (I490084,I2859,I489968,I490124,);
not I_28661 (I489960,I490124);
not I_28662 (I490146,I35759);
nand I_28663 (I490163,I490067,I490146);
DFFARX1 I_28664 (I490163,I2859,I489968,I490189,);
not I_28665 (I490197,I490189);
not I_28666 (I490214,I35750);
nand I_28667 (I490231,I490214,I35768);
and I_28668 (I490248,I490050,I490231);
nor I_28669 (I490265,I490163,I490248);
DFFARX1 I_28670 (I490265,I2859,I489968,I489936,);
DFFARX1 I_28671 (I490248,I2859,I489968,I489957,);
nor I_28672 (I490310,I35750,I35762);
nor I_28673 (I489948,I490163,I490310);
or I_28674 (I490341,I35750,I35762);
nor I_28675 (I490358,I35756,I35747);
DFFARX1 I_28676 (I490358,I2859,I489968,I490384,);
not I_28677 (I490392,I490384);
nor I_28678 (I489954,I490392,I490197);
nand I_28679 (I490423,I490392,I490042);
not I_28680 (I490440,I35756);
nand I_28681 (I490457,I490440,I490146);
nand I_28682 (I490474,I490392,I490457);
nand I_28683 (I489945,I490474,I490423);
nand I_28684 (I489942,I490457,I490341);
not I_28685 (I490546,I2866);
DFFARX1 I_28686 (I45784,I2859,I490546,I490572,);
and I_28687 (I490580,I490572,I45760);
DFFARX1 I_28688 (I490580,I2859,I490546,I490529,);
DFFARX1 I_28689 (I45778,I2859,I490546,I490620,);
not I_28690 (I490628,I45766);
not I_28691 (I490645,I45763);
nand I_28692 (I490662,I490645,I490628);
nor I_28693 (I490517,I490620,I490662);
DFFARX1 I_28694 (I490662,I2859,I490546,I490702,);
not I_28695 (I490538,I490702);
not I_28696 (I490724,I45772);
nand I_28697 (I490741,I490645,I490724);
DFFARX1 I_28698 (I490741,I2859,I490546,I490767,);
not I_28699 (I490775,I490767);
not I_28700 (I490792,I45763);
nand I_28701 (I490809,I490792,I45781);
and I_28702 (I490826,I490628,I490809);
nor I_28703 (I490843,I490741,I490826);
DFFARX1 I_28704 (I490843,I2859,I490546,I490514,);
DFFARX1 I_28705 (I490826,I2859,I490546,I490535,);
nor I_28706 (I490888,I45763,I45775);
nor I_28707 (I490526,I490741,I490888);
or I_28708 (I490919,I45763,I45775);
nor I_28709 (I490936,I45769,I45760);
DFFARX1 I_28710 (I490936,I2859,I490546,I490962,);
not I_28711 (I490970,I490962);
nor I_28712 (I490532,I490970,I490775);
nand I_28713 (I491001,I490970,I490620);
not I_28714 (I491018,I45769);
nand I_28715 (I491035,I491018,I490724);
nand I_28716 (I491052,I490970,I491035);
nand I_28717 (I490523,I491052,I491001);
nand I_28718 (I490520,I491035,I490919);
not I_28719 (I491124,I2866);
DFFARX1 I_28720 (I526918,I2859,I491124,I491150,);
and I_28721 (I491158,I491150,I526900);
DFFARX1 I_28722 (I491158,I2859,I491124,I491107,);
DFFARX1 I_28723 (I526909,I2859,I491124,I491198,);
not I_28724 (I491206,I526894);
not I_28725 (I491223,I526906);
nand I_28726 (I491240,I491223,I491206);
nor I_28727 (I491095,I491198,I491240);
DFFARX1 I_28728 (I491240,I2859,I491124,I491280,);
not I_28729 (I491116,I491280);
not I_28730 (I491302,I526897);
nand I_28731 (I491319,I491223,I491302);
DFFARX1 I_28732 (I491319,I2859,I491124,I491345,);
not I_28733 (I491353,I491345);
not I_28734 (I491370,I526894);
nand I_28735 (I491387,I491370,I526897);
and I_28736 (I491404,I491206,I491387);
nor I_28737 (I491421,I491319,I491404);
DFFARX1 I_28738 (I491421,I2859,I491124,I491092,);
DFFARX1 I_28739 (I491404,I2859,I491124,I491113,);
nor I_28740 (I491466,I526894,I526915);
nor I_28741 (I491104,I491319,I491466);
or I_28742 (I491497,I526894,I526915);
nor I_28743 (I491514,I526903,I526912);
DFFARX1 I_28744 (I491514,I2859,I491124,I491540,);
not I_28745 (I491548,I491540);
nor I_28746 (I491110,I491548,I491353);
nand I_28747 (I491579,I491548,I491198);
not I_28748 (I491596,I526903);
nand I_28749 (I491613,I491596,I491302);
nand I_28750 (I491630,I491548,I491613);
nand I_28751 (I491101,I491630,I491579);
nand I_28752 (I491098,I491613,I491497);
not I_28753 (I491702,I2866);
DFFARX1 I_28754 (I353208,I2859,I491702,I491728,);
and I_28755 (I491736,I491728,I353214);
DFFARX1 I_28756 (I491736,I2859,I491702,I491685,);
DFFARX1 I_28757 (I353220,I2859,I491702,I491776,);
not I_28758 (I491784,I353205);
not I_28759 (I491801,I353205);
nand I_28760 (I491818,I491801,I491784);
nor I_28761 (I491673,I491776,I491818);
DFFARX1 I_28762 (I491818,I2859,I491702,I491858,);
not I_28763 (I491694,I491858);
not I_28764 (I491880,I353223);
nand I_28765 (I491897,I491801,I491880);
DFFARX1 I_28766 (I491897,I2859,I491702,I491923,);
not I_28767 (I491931,I491923);
not I_28768 (I491948,I353217);
nand I_28769 (I491965,I491948,I353208);
and I_28770 (I491982,I491784,I491965);
nor I_28771 (I491999,I491897,I491982);
DFFARX1 I_28772 (I491999,I2859,I491702,I491670,);
DFFARX1 I_28773 (I491982,I2859,I491702,I491691,);
nor I_28774 (I492044,I353217,I353226);
nor I_28775 (I491682,I491897,I492044);
or I_28776 (I492075,I353217,I353226);
nor I_28777 (I492092,I353211,I353211);
DFFARX1 I_28778 (I492092,I2859,I491702,I492118,);
not I_28779 (I492126,I492118);
nor I_28780 (I491688,I492126,I491931);
nand I_28781 (I492157,I492126,I491776);
not I_28782 (I492174,I353211);
nand I_28783 (I492191,I492174,I491880);
nand I_28784 (I492208,I492126,I492191);
nand I_28785 (I491679,I492208,I492157);
nand I_28786 (I491676,I492191,I492075);
not I_28787 (I492280,I2866);
DFFARX1 I_28788 (I311859,I2859,I492280,I492306,);
and I_28789 (I492314,I492306,I311847);
DFFARX1 I_28790 (I492314,I2859,I492280,I492263,);
DFFARX1 I_28791 (I311850,I2859,I492280,I492354,);
not I_28792 (I492362,I311844);
not I_28793 (I492379,I311868);
nand I_28794 (I492396,I492379,I492362);
nor I_28795 (I492251,I492354,I492396);
DFFARX1 I_28796 (I492396,I2859,I492280,I492436,);
not I_28797 (I492272,I492436);
not I_28798 (I492458,I311856);
nand I_28799 (I492475,I492379,I492458);
DFFARX1 I_28800 (I492475,I2859,I492280,I492501,);
not I_28801 (I492509,I492501);
not I_28802 (I492526,I311865);
nand I_28803 (I492543,I492526,I311862);
and I_28804 (I492560,I492362,I492543);
nor I_28805 (I492577,I492475,I492560);
DFFARX1 I_28806 (I492577,I2859,I492280,I492248,);
DFFARX1 I_28807 (I492560,I2859,I492280,I492269,);
nor I_28808 (I492622,I311865,I311853);
nor I_28809 (I492260,I492475,I492622);
or I_28810 (I492653,I311865,I311853);
nor I_28811 (I492670,I311844,I311847);
DFFARX1 I_28812 (I492670,I2859,I492280,I492696,);
not I_28813 (I492704,I492696);
nor I_28814 (I492266,I492704,I492509);
nand I_28815 (I492735,I492704,I492354);
not I_28816 (I492752,I311844);
nand I_28817 (I492769,I492752,I492458);
nand I_28818 (I492786,I492704,I492769);
nand I_28819 (I492257,I492786,I492735);
nand I_28820 (I492254,I492769,I492653);
not I_28821 (I492858,I2866);
DFFARX1 I_28822 (I194459,I2859,I492858,I492884,);
and I_28823 (I492892,I492884,I194474);
DFFARX1 I_28824 (I492892,I2859,I492858,I492841,);
DFFARX1 I_28825 (I194477,I2859,I492858,I492932,);
not I_28826 (I492940,I194471);
not I_28827 (I492957,I194486);
nand I_28828 (I492974,I492957,I492940);
nor I_28829 (I492829,I492932,I492974);
DFFARX1 I_28830 (I492974,I2859,I492858,I493014,);
not I_28831 (I492850,I493014);
not I_28832 (I493036,I194462);
nand I_28833 (I493053,I492957,I493036);
DFFARX1 I_28834 (I493053,I2859,I492858,I493079,);
not I_28835 (I493087,I493079);
not I_28836 (I493104,I194465);
nand I_28837 (I493121,I493104,I194459);
and I_28838 (I493138,I492940,I493121);
nor I_28839 (I493155,I493053,I493138);
DFFARX1 I_28840 (I493155,I2859,I492858,I492826,);
DFFARX1 I_28841 (I493138,I2859,I492858,I492847,);
nor I_28842 (I493200,I194465,I194468);
nor I_28843 (I492838,I493053,I493200);
or I_28844 (I493231,I194465,I194468);
nor I_28845 (I493248,I194483,I194480);
DFFARX1 I_28846 (I493248,I2859,I492858,I493274,);
not I_28847 (I493282,I493274);
nor I_28848 (I492844,I493282,I493087);
nand I_28849 (I493313,I493282,I492932);
not I_28850 (I493330,I194483);
nand I_28851 (I493347,I493330,I493036);
nand I_28852 (I493364,I493282,I493347);
nand I_28853 (I492835,I493364,I493313);
nand I_28854 (I492832,I493347,I493231);
not I_28855 (I493436,I2866);
DFFARX1 I_28856 (I424761,I2859,I493436,I493462,);
and I_28857 (I493470,I493462,I424758);
DFFARX1 I_28858 (I493470,I2859,I493436,I493419,);
DFFARX1 I_28859 (I424764,I2859,I493436,I493510,);
not I_28860 (I493518,I424767);
not I_28861 (I493535,I424761);
nand I_28862 (I493552,I493535,I493518);
nor I_28863 (I493407,I493510,I493552);
DFFARX1 I_28864 (I493552,I2859,I493436,I493592,);
not I_28865 (I493428,I493592);
not I_28866 (I493614,I424776);
nand I_28867 (I493631,I493535,I493614);
DFFARX1 I_28868 (I493631,I2859,I493436,I493657,);
not I_28869 (I493665,I493657);
not I_28870 (I493682,I424773);
nand I_28871 (I493699,I493682,I424779);
and I_28872 (I493716,I493518,I493699);
nor I_28873 (I493733,I493631,I493716);
DFFARX1 I_28874 (I493733,I2859,I493436,I493404,);
DFFARX1 I_28875 (I493716,I2859,I493436,I493425,);
nor I_28876 (I493778,I424773,I424758);
nor I_28877 (I493416,I493631,I493778);
or I_28878 (I493809,I424773,I424758);
nor I_28879 (I493826,I424770,I424764);
DFFARX1 I_28880 (I493826,I2859,I493436,I493852,);
not I_28881 (I493860,I493852);
nor I_28882 (I493422,I493860,I493665);
nand I_28883 (I493891,I493860,I493510);
not I_28884 (I493908,I424770);
nand I_28885 (I493925,I493908,I493614);
nand I_28886 (I493942,I493860,I493925);
nand I_28887 (I493413,I493942,I493891);
nand I_28888 (I493410,I493925,I493809);
not I_28889 (I494014,I2866);
DFFARX1 I_28890 (I50000,I2859,I494014,I494040,);
and I_28891 (I494048,I494040,I49976);
DFFARX1 I_28892 (I494048,I2859,I494014,I493997,);
DFFARX1 I_28893 (I49994,I2859,I494014,I494088,);
not I_28894 (I494096,I49982);
not I_28895 (I494113,I49979);
nand I_28896 (I494130,I494113,I494096);
nor I_28897 (I493985,I494088,I494130);
DFFARX1 I_28898 (I494130,I2859,I494014,I494170,);
not I_28899 (I494006,I494170);
not I_28900 (I494192,I49988);
nand I_28901 (I494209,I494113,I494192);
DFFARX1 I_28902 (I494209,I2859,I494014,I494235,);
not I_28903 (I494243,I494235);
not I_28904 (I494260,I49979);
nand I_28905 (I494277,I494260,I49997);
and I_28906 (I494294,I494096,I494277);
nor I_28907 (I494311,I494209,I494294);
DFFARX1 I_28908 (I494311,I2859,I494014,I493982,);
DFFARX1 I_28909 (I494294,I2859,I494014,I494003,);
nor I_28910 (I494356,I49979,I49991);
nor I_28911 (I493994,I494209,I494356);
or I_28912 (I494387,I49979,I49991);
nor I_28913 (I494404,I49985,I49976);
DFFARX1 I_28914 (I494404,I2859,I494014,I494430,);
not I_28915 (I494438,I494430);
nor I_28916 (I494000,I494438,I494243);
nand I_28917 (I494469,I494438,I494088);
not I_28918 (I494486,I49985);
nand I_28919 (I494503,I494486,I494192);
nand I_28920 (I494520,I494438,I494503);
nand I_28921 (I493991,I494520,I494469);
nand I_28922 (I493988,I494503,I494387);
not I_28923 (I494592,I2866);
DFFARX1 I_28924 (I307235,I2859,I494592,I494618,);
and I_28925 (I494626,I494618,I307223);
DFFARX1 I_28926 (I494626,I2859,I494592,I494575,);
DFFARX1 I_28927 (I307226,I2859,I494592,I494666,);
not I_28928 (I494674,I307220);
not I_28929 (I494691,I307244);
nand I_28930 (I494708,I494691,I494674);
nor I_28931 (I494563,I494666,I494708);
DFFARX1 I_28932 (I494708,I2859,I494592,I494748,);
not I_28933 (I494584,I494748);
not I_28934 (I494770,I307232);
nand I_28935 (I494787,I494691,I494770);
DFFARX1 I_28936 (I494787,I2859,I494592,I494813,);
not I_28937 (I494821,I494813);
not I_28938 (I494838,I307241);
nand I_28939 (I494855,I494838,I307238);
and I_28940 (I494872,I494674,I494855);
nor I_28941 (I494889,I494787,I494872);
DFFARX1 I_28942 (I494889,I2859,I494592,I494560,);
DFFARX1 I_28943 (I494872,I2859,I494592,I494581,);
nor I_28944 (I494934,I307241,I307229);
nor I_28945 (I494572,I494787,I494934);
or I_28946 (I494965,I307241,I307229);
nor I_28947 (I494982,I307220,I307223);
DFFARX1 I_28948 (I494982,I2859,I494592,I495008,);
not I_28949 (I495016,I495008);
nor I_28950 (I494578,I495016,I494821);
nand I_28951 (I495047,I495016,I494666);
not I_28952 (I495064,I307220);
nand I_28953 (I495081,I495064,I494770);
nand I_28954 (I495098,I495016,I495081);
nand I_28955 (I494569,I495098,I495047);
nand I_28956 (I494566,I495081,I494965);
not I_28957 (I495170,I2866);
DFFARX1 I_28958 (I147209,I2859,I495170,I495196,);
and I_28959 (I495204,I495196,I147194);
DFFARX1 I_28960 (I495204,I2859,I495170,I495153,);
DFFARX1 I_28961 (I147200,I2859,I495170,I495244,);
not I_28962 (I495252,I147182);
not I_28963 (I495269,I147203);
nand I_28964 (I495286,I495269,I495252);
nor I_28965 (I495141,I495244,I495286);
DFFARX1 I_28966 (I495286,I2859,I495170,I495326,);
not I_28967 (I495162,I495326);
not I_28968 (I495348,I147206);
nand I_28969 (I495365,I495269,I495348);
DFFARX1 I_28970 (I495365,I2859,I495170,I495391,);
not I_28971 (I495399,I495391);
not I_28972 (I495416,I147197);
nand I_28973 (I495433,I495416,I147185);
and I_28974 (I495450,I495252,I495433);
nor I_28975 (I495467,I495365,I495450);
DFFARX1 I_28976 (I495467,I2859,I495170,I495138,);
DFFARX1 I_28977 (I495450,I2859,I495170,I495159,);
nor I_28978 (I495512,I147197,I147191);
nor I_28979 (I495150,I495365,I495512);
or I_28980 (I495543,I147197,I147191);
nor I_28981 (I495560,I147188,I147182);
DFFARX1 I_28982 (I495560,I2859,I495170,I495586,);
not I_28983 (I495594,I495586);
nor I_28984 (I495156,I495594,I495399);
nand I_28985 (I495625,I495594,I495244);
not I_28986 (I495642,I147188);
nand I_28987 (I495659,I495642,I495348);
nand I_28988 (I495676,I495594,I495659);
nand I_28989 (I495147,I495676,I495625);
nand I_28990 (I495144,I495659,I495543);
not I_28991 (I495748,I2866);
DFFARX1 I_28992 (I256371,I2859,I495748,I495774,);
and I_28993 (I495782,I495774,I256359);
DFFARX1 I_28994 (I495782,I2859,I495748,I495731,);
DFFARX1 I_28995 (I256374,I2859,I495748,I495822,);
not I_28996 (I495830,I256365);
not I_28997 (I495847,I256356);
nand I_28998 (I495864,I495847,I495830);
nor I_28999 (I495719,I495822,I495864);
DFFARX1 I_29000 (I495864,I2859,I495748,I495904,);
not I_29001 (I495740,I495904);
not I_29002 (I495926,I256362);
nand I_29003 (I495943,I495847,I495926);
DFFARX1 I_29004 (I495943,I2859,I495748,I495969,);
not I_29005 (I495977,I495969);
not I_29006 (I495994,I256377);
nand I_29007 (I496011,I495994,I256380);
and I_29008 (I496028,I495830,I496011);
nor I_29009 (I496045,I495943,I496028);
DFFARX1 I_29010 (I496045,I2859,I495748,I495716,);
DFFARX1 I_29011 (I496028,I2859,I495748,I495737,);
nor I_29012 (I496090,I256377,I256356);
nor I_29013 (I495728,I495943,I496090);
or I_29014 (I496121,I256377,I256356);
nor I_29015 (I496138,I256368,I256359);
DFFARX1 I_29016 (I496138,I2859,I495748,I496164,);
not I_29017 (I496172,I496164);
nor I_29018 (I495734,I496172,I495977);
nand I_29019 (I496203,I496172,I495822);
not I_29020 (I496220,I256368);
nand I_29021 (I496237,I496220,I495926);
nand I_29022 (I496254,I496172,I496237);
nand I_29023 (I495725,I496254,I496203);
nand I_29024 (I495722,I496237,I496121);
not I_29025 (I496326,I2866);
DFFARX1 I_29026 (I132453,I2859,I496326,I496352,);
and I_29027 (I496360,I496352,I132438);
DFFARX1 I_29028 (I496360,I2859,I496326,I496309,);
DFFARX1 I_29029 (I132444,I2859,I496326,I496400,);
not I_29030 (I496408,I132426);
not I_29031 (I496425,I132447);
nand I_29032 (I496442,I496425,I496408);
nor I_29033 (I496297,I496400,I496442);
DFFARX1 I_29034 (I496442,I2859,I496326,I496482,);
not I_29035 (I496318,I496482);
not I_29036 (I496504,I132450);
nand I_29037 (I496521,I496425,I496504);
DFFARX1 I_29038 (I496521,I2859,I496326,I496547,);
not I_29039 (I496555,I496547);
not I_29040 (I496572,I132441);
nand I_29041 (I496589,I496572,I132429);
and I_29042 (I496606,I496408,I496589);
nor I_29043 (I496623,I496521,I496606);
DFFARX1 I_29044 (I496623,I2859,I496326,I496294,);
DFFARX1 I_29045 (I496606,I2859,I496326,I496315,);
nor I_29046 (I496668,I132441,I132435);
nor I_29047 (I496306,I496521,I496668);
or I_29048 (I496699,I132441,I132435);
nor I_29049 (I496716,I132432,I132426);
DFFARX1 I_29050 (I496716,I2859,I496326,I496742,);
not I_29051 (I496750,I496742);
nor I_29052 (I496312,I496750,I496555);
nand I_29053 (I496781,I496750,I496400);
not I_29054 (I496798,I132432);
nand I_29055 (I496815,I496798,I496504);
nand I_29056 (I496832,I496750,I496815);
nand I_29057 (I496303,I496832,I496781);
nand I_29058 (I496300,I496815,I496699);
not I_29059 (I496904,I2866);
DFFARX1 I_29060 (I2188,I2859,I496904,I496930,);
and I_29061 (I496938,I496930,I2340);
DFFARX1 I_29062 (I496938,I2859,I496904,I496887,);
DFFARX1 I_29063 (I2420,I2859,I496904,I496978,);
not I_29064 (I496986,I2540);
not I_29065 (I497003,I2740);
nand I_29066 (I497020,I497003,I496986);
nor I_29067 (I496875,I496978,I497020);
DFFARX1 I_29068 (I497020,I2859,I496904,I497060,);
not I_29069 (I496896,I497060);
not I_29070 (I497082,I1740);
nand I_29071 (I497099,I497003,I497082);
DFFARX1 I_29072 (I497099,I2859,I496904,I497125,);
not I_29073 (I497133,I497125);
not I_29074 (I497150,I2476);
nand I_29075 (I497167,I497150,I1668);
and I_29076 (I497184,I496986,I497167);
nor I_29077 (I497201,I497099,I497184);
DFFARX1 I_29078 (I497201,I2859,I496904,I496872,);
DFFARX1 I_29079 (I497184,I2859,I496904,I496893,);
nor I_29080 (I497246,I2476,I2660);
nor I_29081 (I496884,I497099,I497246);
or I_29082 (I497277,I2476,I2660);
nor I_29083 (I497294,I1620,I2628);
DFFARX1 I_29084 (I497294,I2859,I496904,I497320,);
not I_29085 (I497328,I497320);
nor I_29086 (I496890,I497328,I497133);
nand I_29087 (I497359,I497328,I496978);
not I_29088 (I497376,I1620);
nand I_29089 (I497393,I497376,I497082);
nand I_29090 (I497410,I497328,I497393);
nand I_29091 (I496881,I497410,I497359);
nand I_29092 (I496878,I497393,I497277);
not I_29093 (I497482,I2866);
DFFARX1 I_29094 (I389319,I2859,I497482,I497508,);
and I_29095 (I497516,I497508,I389313);
DFFARX1 I_29096 (I497516,I2859,I497482,I497465,);
DFFARX1 I_29097 (I389331,I2859,I497482,I497556,);
not I_29098 (I497564,I389322);
not I_29099 (I497581,I389334);
nand I_29100 (I497598,I497581,I497564);
nor I_29101 (I497453,I497556,I497598);
DFFARX1 I_29102 (I497598,I2859,I497482,I497638,);
not I_29103 (I497474,I497638);
not I_29104 (I497660,I389340);
nand I_29105 (I497677,I497581,I497660);
DFFARX1 I_29106 (I497677,I2859,I497482,I497703,);
not I_29107 (I497711,I497703);
not I_29108 (I497728,I389316);
nand I_29109 (I497745,I497728,I389337);
and I_29110 (I497762,I497564,I497745);
nor I_29111 (I497779,I497677,I497762);
DFFARX1 I_29112 (I497779,I2859,I497482,I497450,);
DFFARX1 I_29113 (I497762,I2859,I497482,I497471,);
nor I_29114 (I497824,I389316,I389328);
nor I_29115 (I497462,I497677,I497824);
or I_29116 (I497855,I389316,I389328);
nor I_29117 (I497872,I389313,I389325);
DFFARX1 I_29118 (I497872,I2859,I497482,I497898,);
not I_29119 (I497906,I497898);
nor I_29120 (I497468,I497906,I497711);
nand I_29121 (I497937,I497906,I497556);
not I_29122 (I497954,I389313);
nand I_29123 (I497971,I497954,I497660);
nand I_29124 (I497988,I497906,I497971);
nand I_29125 (I497459,I497988,I497937);
nand I_29126 (I497456,I497971,I497855);
not I_29127 (I498060,I2866);
DFFARX1 I_29128 (I246545,I2859,I498060,I498086,);
and I_29129 (I498094,I498086,I246533);
DFFARX1 I_29130 (I498094,I2859,I498060,I498043,);
DFFARX1 I_29131 (I246548,I2859,I498060,I498134,);
not I_29132 (I498142,I246539);
not I_29133 (I498159,I246530);
nand I_29134 (I498176,I498159,I498142);
nor I_29135 (I498031,I498134,I498176);
DFFARX1 I_29136 (I498176,I2859,I498060,I498216,);
not I_29137 (I498052,I498216);
not I_29138 (I498238,I246536);
nand I_29139 (I498255,I498159,I498238);
DFFARX1 I_29140 (I498255,I2859,I498060,I498281,);
not I_29141 (I498289,I498281);
not I_29142 (I498306,I246551);
nand I_29143 (I498323,I498306,I246554);
and I_29144 (I498340,I498142,I498323);
nor I_29145 (I498357,I498255,I498340);
DFFARX1 I_29146 (I498357,I2859,I498060,I498028,);
DFFARX1 I_29147 (I498340,I2859,I498060,I498049,);
nor I_29148 (I498402,I246551,I246530);
nor I_29149 (I498040,I498255,I498402);
or I_29150 (I498433,I246551,I246530);
nor I_29151 (I498450,I246542,I246533);
DFFARX1 I_29152 (I498450,I2859,I498060,I498476,);
not I_29153 (I498484,I498476);
nor I_29154 (I498046,I498484,I498289);
nand I_29155 (I498515,I498484,I498134);
not I_29156 (I498532,I246542);
nand I_29157 (I498549,I498532,I498238);
nand I_29158 (I498566,I498484,I498549);
nand I_29159 (I498037,I498566,I498515);
nand I_29160 (I498034,I498549,I498433);
not I_29161 (I498638,I2866);
DFFARX1 I_29162 (I2460,I2859,I498638,I498664,);
and I_29163 (I498672,I498664,I1556);
DFFARX1 I_29164 (I498672,I2859,I498638,I498621,);
DFFARX1 I_29165 (I1636,I2859,I498638,I498712,);
not I_29166 (I498720,I2492);
not I_29167 (I498737,I1892);
nand I_29168 (I498754,I498737,I498720);
nor I_29169 (I498609,I498712,I498754);
DFFARX1 I_29170 (I498754,I2859,I498638,I498794,);
not I_29171 (I498630,I498794);
not I_29172 (I498816,I1844);
nand I_29173 (I498833,I498737,I498816);
DFFARX1 I_29174 (I498833,I2859,I498638,I498859,);
not I_29175 (I498867,I498859);
not I_29176 (I498884,I2748);
nand I_29177 (I498901,I498884,I1372);
and I_29178 (I498918,I498720,I498901);
nor I_29179 (I498935,I498833,I498918);
DFFARX1 I_29180 (I498935,I2859,I498638,I498606,);
DFFARX1 I_29181 (I498918,I2859,I498638,I498627,);
nor I_29182 (I498980,I2748,I2308);
nor I_29183 (I498618,I498833,I498980);
or I_29184 (I499011,I2748,I2308);
nor I_29185 (I499028,I2508,I1404);
DFFARX1 I_29186 (I499028,I2859,I498638,I499054,);
not I_29187 (I499062,I499054);
nor I_29188 (I498624,I499062,I498867);
nand I_29189 (I499093,I499062,I498712);
not I_29190 (I499110,I2508);
nand I_29191 (I499127,I499110,I498816);
nand I_29192 (I499144,I499062,I499127);
nand I_29193 (I498615,I499144,I499093);
nand I_29194 (I498612,I499127,I499011);
not I_29195 (I499216,I2866);
DFFARX1 I_29196 (I286427,I2859,I499216,I499242,);
and I_29197 (I499250,I499242,I286415);
DFFARX1 I_29198 (I499250,I2859,I499216,I499199,);
DFFARX1 I_29199 (I286418,I2859,I499216,I499290,);
not I_29200 (I499298,I286412);
not I_29201 (I499315,I286436);
nand I_29202 (I499332,I499315,I499298);
nor I_29203 (I499187,I499290,I499332);
DFFARX1 I_29204 (I499332,I2859,I499216,I499372,);
not I_29205 (I499208,I499372);
not I_29206 (I499394,I286424);
nand I_29207 (I499411,I499315,I499394);
DFFARX1 I_29208 (I499411,I2859,I499216,I499437,);
not I_29209 (I499445,I499437);
not I_29210 (I499462,I286433);
nand I_29211 (I499479,I499462,I286430);
and I_29212 (I499496,I499298,I499479);
nor I_29213 (I499513,I499411,I499496);
DFFARX1 I_29214 (I499513,I2859,I499216,I499184,);
DFFARX1 I_29215 (I499496,I2859,I499216,I499205,);
nor I_29216 (I499558,I286433,I286421);
nor I_29217 (I499196,I499411,I499558);
or I_29218 (I499589,I286433,I286421);
nor I_29219 (I499606,I286412,I286415);
DFFARX1 I_29220 (I499606,I2859,I499216,I499632,);
not I_29221 (I499640,I499632);
nor I_29222 (I499202,I499640,I499445);
nand I_29223 (I499671,I499640,I499290);
not I_29224 (I499688,I286412);
nand I_29225 (I499705,I499688,I499394);
nand I_29226 (I499722,I499640,I499705);
nand I_29227 (I499193,I499722,I499671);
nand I_29228 (I499190,I499705,I499589);
not I_29229 (I499794,I2866);
DFFARX1 I_29230 (I61978,I2859,I499794,I499820,);
and I_29231 (I499828,I499820,I62002);
DFFARX1 I_29232 (I499828,I2859,I499794,I499777,);
DFFARX1 I_29233 (I61978,I2859,I499794,I499868,);
not I_29234 (I499876,I61996);
not I_29235 (I499893,I61981);
nand I_29236 (I499910,I499893,I499876);
nor I_29237 (I499765,I499868,I499910);
DFFARX1 I_29238 (I499910,I2859,I499794,I499950,);
not I_29239 (I499786,I499950);
not I_29240 (I499972,I61990);
nand I_29241 (I499989,I499893,I499972);
DFFARX1 I_29242 (I499989,I2859,I499794,I500015,);
not I_29243 (I500023,I500015);
not I_29244 (I500040,I61987);
nand I_29245 (I500057,I500040,I61984);
and I_29246 (I500074,I499876,I500057);
nor I_29247 (I500091,I499989,I500074);
DFFARX1 I_29248 (I500091,I2859,I499794,I499762,);
DFFARX1 I_29249 (I500074,I2859,I499794,I499783,);
nor I_29250 (I500136,I61987,I61993);
nor I_29251 (I499774,I499989,I500136);
or I_29252 (I500167,I61987,I61993);
nor I_29253 (I500184,I61999,I62005);
DFFARX1 I_29254 (I500184,I2859,I499794,I500210,);
not I_29255 (I500218,I500210);
nor I_29256 (I499780,I500218,I500023);
nand I_29257 (I500249,I500218,I499868);
not I_29258 (I500266,I61999);
nand I_29259 (I500283,I500266,I499972);
nand I_29260 (I500300,I500218,I500283);
nand I_29261 (I499771,I500300,I500249);
nand I_29262 (I499768,I500283,I500167);
not I_29263 (I500372,I2866);
DFFARX1 I_29264 (I380921,I2859,I500372,I500398,);
and I_29265 (I500406,I500398,I380915);
DFFARX1 I_29266 (I500406,I2859,I500372,I500355,);
DFFARX1 I_29267 (I380933,I2859,I500372,I500446,);
not I_29268 (I500454,I380924);
not I_29269 (I500471,I380936);
nand I_29270 (I500488,I500471,I500454);
nor I_29271 (I500343,I500446,I500488);
DFFARX1 I_29272 (I500488,I2859,I500372,I500528,);
not I_29273 (I500364,I500528);
not I_29274 (I500550,I380942);
nand I_29275 (I500567,I500471,I500550);
DFFARX1 I_29276 (I500567,I2859,I500372,I500593,);
not I_29277 (I500601,I500593);
not I_29278 (I500618,I380918);
nand I_29279 (I500635,I500618,I380939);
and I_29280 (I500652,I500454,I500635);
nor I_29281 (I500669,I500567,I500652);
DFFARX1 I_29282 (I500669,I2859,I500372,I500340,);
DFFARX1 I_29283 (I500652,I2859,I500372,I500361,);
nor I_29284 (I500714,I380918,I380930);
nor I_29285 (I500352,I500567,I500714);
or I_29286 (I500745,I380918,I380930);
nor I_29287 (I500762,I380915,I380927);
DFFARX1 I_29288 (I500762,I2859,I500372,I500788,);
not I_29289 (I500796,I500788);
nor I_29290 (I500358,I500796,I500601);
nand I_29291 (I500827,I500796,I500446);
not I_29292 (I500844,I380915);
nand I_29293 (I500861,I500844,I500550);
nand I_29294 (I500878,I500796,I500861);
nand I_29295 (I500349,I500878,I500827);
nand I_29296 (I500346,I500861,I500745);
not I_29297 (I500950,I2866);
DFFARX1 I_29298 (I70308,I2859,I500950,I500976,);
and I_29299 (I500984,I500976,I70311);
DFFARX1 I_29300 (I500984,I2859,I500950,I500933,);
DFFARX1 I_29301 (I70311,I2859,I500950,I501024,);
not I_29302 (I501032,I70326);
not I_29303 (I501049,I70332);
nand I_29304 (I501066,I501049,I501032);
nor I_29305 (I500921,I501024,I501066);
DFFARX1 I_29306 (I501066,I2859,I500950,I501106,);
not I_29307 (I500942,I501106);
not I_29308 (I501128,I70320);
nand I_29309 (I501145,I501049,I501128);
DFFARX1 I_29310 (I501145,I2859,I500950,I501171,);
not I_29311 (I501179,I501171);
not I_29312 (I501196,I70317);
nand I_29313 (I501213,I501196,I70314);
and I_29314 (I501230,I501032,I501213);
nor I_29315 (I501247,I501145,I501230);
DFFARX1 I_29316 (I501247,I2859,I500950,I500918,);
DFFARX1 I_29317 (I501230,I2859,I500950,I500939,);
nor I_29318 (I501292,I70317,I70308);
nor I_29319 (I500930,I501145,I501292);
or I_29320 (I501323,I70317,I70308);
nor I_29321 (I501340,I70323,I70329);
DFFARX1 I_29322 (I501340,I2859,I500950,I501366,);
not I_29323 (I501374,I501366);
nor I_29324 (I500936,I501374,I501179);
nand I_29325 (I501405,I501374,I501024);
not I_29326 (I501422,I70323);
nand I_29327 (I501439,I501422,I501128);
nand I_29328 (I501456,I501374,I501439);
nand I_29329 (I500927,I501456,I501405);
nand I_29330 (I500924,I501439,I501323);
not I_29331 (I501528,I2866);
DFFARX1 I_29332 (I8870,I2859,I501528,I501554,);
and I_29333 (I501562,I501554,I8873);
DFFARX1 I_29334 (I501562,I2859,I501528,I501511,);
DFFARX1 I_29335 (I8873,I2859,I501528,I501602,);
not I_29336 (I501610,I8876);
not I_29337 (I501627,I8891);
nand I_29338 (I501644,I501627,I501610);
nor I_29339 (I501499,I501602,I501644);
DFFARX1 I_29340 (I501644,I2859,I501528,I501684,);
not I_29341 (I501520,I501684);
not I_29342 (I501706,I8885);
nand I_29343 (I501723,I501627,I501706);
DFFARX1 I_29344 (I501723,I2859,I501528,I501749,);
not I_29345 (I501757,I501749);
not I_29346 (I501774,I8888);
nand I_29347 (I501791,I501774,I8870);
and I_29348 (I501808,I501610,I501791);
nor I_29349 (I501825,I501723,I501808);
DFFARX1 I_29350 (I501825,I2859,I501528,I501496,);
DFFARX1 I_29351 (I501808,I2859,I501528,I501517,);
nor I_29352 (I501870,I8888,I8882);
nor I_29353 (I501508,I501723,I501870);
or I_29354 (I501901,I8888,I8882);
nor I_29355 (I501918,I8879,I8894);
DFFARX1 I_29356 (I501918,I2859,I501528,I501944,);
not I_29357 (I501952,I501944);
nor I_29358 (I501514,I501952,I501757);
nand I_29359 (I501983,I501952,I501602);
not I_29360 (I502000,I8879);
nand I_29361 (I502017,I502000,I501706);
nand I_29362 (I502034,I501952,I502017);
nand I_29363 (I501505,I502034,I501983);
nand I_29364 (I501502,I502017,I501901);
not I_29365 (I502106,I2866);
DFFARX1 I_29366 (I465684,I2859,I502106,I502132,);
nand I_29367 (I502140,I502132,I465663);
DFFARX1 I_29368 (I465660,I2859,I502106,I502166,);
DFFARX1 I_29369 (I502166,I2859,I502106,I502183,);
not I_29370 (I502098,I502183);
not I_29371 (I502205,I465672);
nor I_29372 (I502222,I465672,I465681);
not I_29373 (I502239,I465669);
nand I_29374 (I502256,I502205,I502239);
nor I_29375 (I502273,I465669,I465672);
and I_29376 (I502077,I502273,I502140);
not I_29377 (I502304,I465678);
nand I_29378 (I502321,I502304,I465675);
nor I_29379 (I502338,I465678,I465660);
not I_29380 (I502355,I502338);
nand I_29381 (I502080,I502222,I502355);
DFFARX1 I_29382 (I502338,I2859,I502106,I502095,);
nor I_29383 (I502400,I465663,I465669);
nor I_29384 (I502417,I502400,I465681);
and I_29385 (I502434,I502417,I502321);
DFFARX1 I_29386 (I502434,I2859,I502106,I502092,);
nor I_29387 (I502089,I502400,I502256);
or I_29388 (I502086,I502338,I502400);
nor I_29389 (I502493,I465663,I465666);
DFFARX1 I_29390 (I502493,I2859,I502106,I502519,);
not I_29391 (I502527,I502519);
nand I_29392 (I502544,I502527,I502205);
nor I_29393 (I502561,I502544,I465681);
DFFARX1 I_29394 (I502561,I2859,I502106,I502074,);
nor I_29395 (I502592,I502527,I502256);
nor I_29396 (I502083,I502400,I502592);
not I_29397 (I502650,I2866);
DFFARX1 I_29398 (I132965,I2859,I502650,I502676,);
nand I_29399 (I502684,I502676,I132968);
DFFARX1 I_29400 (I132962,I2859,I502650,I502710,);
DFFARX1 I_29401 (I502710,I2859,I502650,I502727,);
not I_29402 (I502642,I502727);
not I_29403 (I502749,I132971);
nor I_29404 (I502766,I132971,I132956);
not I_29405 (I502783,I132980);
nand I_29406 (I502800,I502749,I502783);
nor I_29407 (I502817,I132980,I132971);
and I_29408 (I502621,I502817,I502684);
not I_29409 (I502848,I132959);
nand I_29410 (I502865,I502848,I132977);
nor I_29411 (I502882,I132959,I132953);
not I_29412 (I502899,I502882);
nand I_29413 (I502624,I502766,I502899);
DFFARX1 I_29414 (I502882,I2859,I502650,I502639,);
nor I_29415 (I502944,I132974,I132980);
nor I_29416 (I502961,I502944,I132956);
and I_29417 (I502978,I502961,I502865);
DFFARX1 I_29418 (I502978,I2859,I502650,I502636,);
nor I_29419 (I502633,I502944,I502800);
or I_29420 (I502630,I502882,I502944);
nor I_29421 (I503037,I132974,I132953);
DFFARX1 I_29422 (I503037,I2859,I502650,I503063,);
not I_29423 (I503071,I503063);
nand I_29424 (I503088,I503071,I502749);
nor I_29425 (I503105,I503088,I132956);
DFFARX1 I_29426 (I503105,I2859,I502650,I502618,);
nor I_29427 (I503136,I503071,I502800);
nor I_29428 (I502627,I502944,I503136);
not I_29429 (I503194,I2866);
DFFARX1 I_29430 (I494584,I2859,I503194,I503220,);
nand I_29431 (I503228,I503220,I494563);
DFFARX1 I_29432 (I494560,I2859,I503194,I503254,);
DFFARX1 I_29433 (I503254,I2859,I503194,I503271,);
not I_29434 (I503186,I503271);
not I_29435 (I503293,I494572);
nor I_29436 (I503310,I494572,I494581);
not I_29437 (I503327,I494569);
nand I_29438 (I503344,I503293,I503327);
nor I_29439 (I503361,I494569,I494572);
and I_29440 (I503165,I503361,I503228);
not I_29441 (I503392,I494578);
nand I_29442 (I503409,I503392,I494575);
nor I_29443 (I503426,I494578,I494560);
not I_29444 (I503443,I503426);
nand I_29445 (I503168,I503310,I503443);
DFFARX1 I_29446 (I503426,I2859,I503194,I503183,);
nor I_29447 (I503488,I494563,I494569);
nor I_29448 (I503505,I503488,I494581);
and I_29449 (I503522,I503505,I503409);
DFFARX1 I_29450 (I503522,I2859,I503194,I503180,);
nor I_29451 (I503177,I503488,I503344);
or I_29452 (I503174,I503426,I503488);
nor I_29453 (I503581,I494563,I494566);
DFFARX1 I_29454 (I503581,I2859,I503194,I503607,);
not I_29455 (I503615,I503607);
nand I_29456 (I503632,I503615,I503293);
nor I_29457 (I503649,I503632,I494581);
DFFARX1 I_29458 (I503649,I2859,I503194,I503162,);
nor I_29459 (I503680,I503615,I503344);
nor I_29460 (I503171,I503488,I503680);
not I_29461 (I503738,I2866);
DFFARX1 I_29462 (I471464,I2859,I503738,I503764,);
nand I_29463 (I503772,I503764,I471443);
DFFARX1 I_29464 (I471440,I2859,I503738,I503798,);
DFFARX1 I_29465 (I503798,I2859,I503738,I503815,);
not I_29466 (I503730,I503815);
not I_29467 (I503837,I471452);
nor I_29468 (I503854,I471452,I471461);
not I_29469 (I503871,I471449);
nand I_29470 (I503888,I503837,I503871);
nor I_29471 (I503905,I471449,I471452);
and I_29472 (I503709,I503905,I503772);
not I_29473 (I503936,I471458);
nand I_29474 (I503953,I503936,I471455);
nor I_29475 (I503970,I471458,I471440);
not I_29476 (I503987,I503970);
nand I_29477 (I503712,I503854,I503987);
DFFARX1 I_29478 (I503970,I2859,I503738,I503727,);
nor I_29479 (I504032,I471443,I471449);
nor I_29480 (I504049,I504032,I471461);
and I_29481 (I504066,I504049,I503953);
DFFARX1 I_29482 (I504066,I2859,I503738,I503724,);
nor I_29483 (I503721,I504032,I503888);
or I_29484 (I503718,I503970,I504032);
nor I_29485 (I504125,I471443,I471446);
DFFARX1 I_29486 (I504125,I2859,I503738,I504151,);
not I_29487 (I504159,I504151);
nand I_29488 (I504176,I504159,I503837);
nor I_29489 (I504193,I504176,I471461);
DFFARX1 I_29490 (I504193,I2859,I503738,I503706,);
nor I_29491 (I504224,I504159,I503888);
nor I_29492 (I503715,I504032,I504224);
not I_29493 (I504282,I2866);
DFFARX1 I_29494 (I379623,I2859,I504282,I504308,);
nand I_29495 (I504316,I504308,I379623);
DFFARX1 I_29496 (I379635,I2859,I504282,I504342,);
DFFARX1 I_29497 (I504342,I2859,I504282,I504359,);
not I_29498 (I504274,I504359);
not I_29499 (I504381,I379629);
nor I_29500 (I504398,I379629,I379650);
not I_29501 (I504415,I379638);
nand I_29502 (I504432,I504381,I504415);
nor I_29503 (I504449,I379638,I379629);
and I_29504 (I504253,I504449,I504316);
not I_29505 (I504480,I379632);
nand I_29506 (I504497,I504480,I379647);
nor I_29507 (I504514,I379632,I379641);
not I_29508 (I504531,I504514);
nand I_29509 (I504256,I504398,I504531);
DFFARX1 I_29510 (I504514,I2859,I504282,I504271,);
nor I_29511 (I504576,I379644,I379638);
nor I_29512 (I504593,I504576,I379650);
and I_29513 (I504610,I504593,I504497);
DFFARX1 I_29514 (I504610,I2859,I504282,I504268,);
nor I_29515 (I504265,I504576,I504432);
or I_29516 (I504262,I504514,I504576);
nor I_29517 (I504669,I379644,I379626);
DFFARX1 I_29518 (I504669,I2859,I504282,I504695,);
not I_29519 (I504703,I504695);
nand I_29520 (I504720,I504703,I504381);
nor I_29521 (I504737,I504720,I379650);
DFFARX1 I_29522 (I504737,I2859,I504282,I504250,);
nor I_29523 (I504768,I504703,I504432);
nor I_29524 (I504259,I504576,I504768);
not I_29525 (I504826,I2866);
DFFARX1 I_29526 (I377685,I2859,I504826,I504852,);
nand I_29527 (I504860,I504852,I377685);
DFFARX1 I_29528 (I377697,I2859,I504826,I504886,);
DFFARX1 I_29529 (I504886,I2859,I504826,I504903,);
not I_29530 (I504818,I504903);
not I_29531 (I504925,I377691);
nor I_29532 (I504942,I377691,I377712);
not I_29533 (I504959,I377700);
nand I_29534 (I504976,I504925,I504959);
nor I_29535 (I504993,I377700,I377691);
and I_29536 (I504797,I504993,I504860);
not I_29537 (I505024,I377694);
nand I_29538 (I505041,I505024,I377709);
nor I_29539 (I505058,I377694,I377703);
not I_29540 (I505075,I505058);
nand I_29541 (I504800,I504942,I505075);
DFFARX1 I_29542 (I505058,I2859,I504826,I504815,);
nor I_29543 (I505120,I377706,I377700);
nor I_29544 (I505137,I505120,I377712);
and I_29545 (I505154,I505137,I505041);
DFFARX1 I_29546 (I505154,I2859,I504826,I504812,);
nor I_29547 (I504809,I505120,I504976);
or I_29548 (I504806,I505058,I505120);
nor I_29549 (I505213,I377706,I377688);
DFFARX1 I_29550 (I505213,I2859,I504826,I505239,);
not I_29551 (I505247,I505239);
nand I_29552 (I505264,I505247,I504925);
nor I_29553 (I505281,I505264,I377712);
DFFARX1 I_29554 (I505281,I2859,I504826,I504794,);
nor I_29555 (I505312,I505247,I504976);
nor I_29556 (I504803,I505120,I505312);
not I_29557 (I505370,I2866);
DFFARX1 I_29558 (I276011,I2859,I505370,I505396,);
nand I_29559 (I505404,I505396,I276026);
DFFARX1 I_29560 (I276020,I2859,I505370,I505430,);
DFFARX1 I_29561 (I505430,I2859,I505370,I505447,);
not I_29562 (I505362,I505447);
not I_29563 (I505469,I276023);
nor I_29564 (I505486,I276023,I276029);
not I_29565 (I505503,I276011);
nand I_29566 (I505520,I505469,I505503);
nor I_29567 (I505537,I276011,I276023);
and I_29568 (I505341,I505537,I505404);
not I_29569 (I505568,I276008);
nand I_29570 (I505585,I505568,I276014);
nor I_29571 (I505602,I276008,I276008);
not I_29572 (I505619,I505602);
nand I_29573 (I505344,I505486,I505619);
DFFARX1 I_29574 (I505602,I2859,I505370,I505359,);
nor I_29575 (I505664,I276017,I276011);
nor I_29576 (I505681,I505664,I276029);
and I_29577 (I505698,I505681,I505585);
DFFARX1 I_29578 (I505698,I2859,I505370,I505356,);
nor I_29579 (I505353,I505664,I505520);
or I_29580 (I505350,I505602,I505664);
nor I_29581 (I505757,I276017,I276032);
DFFARX1 I_29582 (I505757,I2859,I505370,I505783,);
not I_29583 (I505791,I505783);
nand I_29584 (I505808,I505791,I505469);
nor I_29585 (I505825,I505808,I276029);
DFFARX1 I_29586 (I505825,I2859,I505370,I505338,);
nor I_29587 (I505856,I505791,I505520);
nor I_29588 (I505347,I505664,I505856);
not I_29589 (I505914,I2866);
DFFARX1 I_29590 (I85787,I2859,I505914,I505940,);
nand I_29591 (I505948,I505940,I85802);
DFFARX1 I_29592 (I85799,I2859,I505914,I505974,);
DFFARX1 I_29593 (I505974,I2859,I505914,I505991,);
not I_29594 (I505906,I505991);
not I_29595 (I506013,I85778);
nor I_29596 (I506030,I85778,I85784);
not I_29597 (I506047,I85790);
nand I_29598 (I506064,I506013,I506047);
nor I_29599 (I506081,I85790,I85778);
and I_29600 (I505885,I506081,I505948);
not I_29601 (I506112,I85796);
nand I_29602 (I506129,I506112,I85778);
nor I_29603 (I506146,I85796,I85781);
not I_29604 (I506163,I506146);
nand I_29605 (I505888,I506030,I506163);
DFFARX1 I_29606 (I506146,I2859,I505914,I505903,);
nor I_29607 (I506208,I85781,I85790);
nor I_29608 (I506225,I506208,I85784);
and I_29609 (I506242,I506225,I506129);
DFFARX1 I_29610 (I506242,I2859,I505914,I505900,);
nor I_29611 (I505897,I506208,I506064);
or I_29612 (I505894,I506146,I506208);
nor I_29613 (I506301,I85781,I85793);
DFFARX1 I_29614 (I506301,I2859,I505914,I506327,);
not I_29615 (I506335,I506327);
nand I_29616 (I506352,I506335,I506013);
nor I_29617 (I506369,I506352,I85784);
DFFARX1 I_29618 (I506369,I2859,I505914,I505882,);
nor I_29619 (I506400,I506335,I506064);
nor I_29620 (I505891,I506208,I506400);
not I_29621 (I506458,I2866);
DFFARX1 I_29622 (I51051,I2859,I506458,I506484,);
nand I_29623 (I506492,I506484,I51033);
DFFARX1 I_29624 (I51030,I2859,I506458,I506518,);
DFFARX1 I_29625 (I506518,I2859,I506458,I506535,);
not I_29626 (I506450,I506535);
not I_29627 (I506557,I51048);
nor I_29628 (I506574,I51048,I51042);
not I_29629 (I506591,I51030);
nand I_29630 (I506608,I506557,I506591);
nor I_29631 (I506625,I51030,I51048);
and I_29632 (I506429,I506625,I506492);
not I_29633 (I506656,I51039);
nand I_29634 (I506673,I506656,I51045);
nor I_29635 (I506690,I51039,I51033);
not I_29636 (I506707,I506690);
nand I_29637 (I506432,I506574,I506707);
DFFARX1 I_29638 (I506690,I2859,I506458,I506447,);
nor I_29639 (I506752,I51036,I51030);
nor I_29640 (I506769,I506752,I51042);
and I_29641 (I506786,I506769,I506673);
DFFARX1 I_29642 (I506786,I2859,I506458,I506444,);
nor I_29643 (I506441,I506752,I506608);
or I_29644 (I506438,I506690,I506752);
nor I_29645 (I506845,I51036,I51054);
DFFARX1 I_29646 (I506845,I2859,I506458,I506871,);
not I_29647 (I506879,I506871);
nand I_29648 (I506896,I506879,I506557);
nor I_29649 (I506913,I506896,I51042);
DFFARX1 I_29650 (I506913,I2859,I506458,I506426,);
nor I_29651 (I506944,I506879,I506608);
nor I_29652 (I506435,I506752,I506944);
not I_29653 (I507002,I2866);
DFFARX1 I_29654 (I429825,I2859,I507002,I507028,);
nand I_29655 (I507036,I507028,I429813);
DFFARX1 I_29656 (I429807,I2859,I507002,I507062,);
DFFARX1 I_29657 (I507062,I2859,I507002,I507079,);
not I_29658 (I506994,I507079);
not I_29659 (I507101,I429807);
nor I_29660 (I507118,I429807,I429819);
not I_29661 (I507135,I429816);
nand I_29662 (I507152,I507101,I507135);
nor I_29663 (I507169,I429816,I429807);
and I_29664 (I506973,I507169,I507036);
not I_29665 (I507200,I429810);
nand I_29666 (I507217,I507200,I429822);
nor I_29667 (I507234,I429810,I429828);
not I_29668 (I507251,I507234);
nand I_29669 (I506976,I507118,I507251);
DFFARX1 I_29670 (I507234,I2859,I507002,I506991,);
nor I_29671 (I507296,I429813,I429816);
nor I_29672 (I507313,I507296,I429819);
and I_29673 (I507330,I507313,I507217);
DFFARX1 I_29674 (I507330,I2859,I507002,I506988,);
nor I_29675 (I506985,I507296,I507152);
or I_29676 (I506982,I507234,I507296);
nor I_29677 (I507389,I429813,I429810);
DFFARX1 I_29678 (I507389,I2859,I507002,I507415,);
not I_29679 (I507423,I507415);
nand I_29680 (I507440,I507423,I507101);
nor I_29681 (I507457,I507440,I429819);
DFFARX1 I_29682 (I507457,I2859,I507002,I506970,);
nor I_29683 (I507488,I507423,I507152);
nor I_29684 (I506979,I507296,I507488);
not I_29685 (I507546,I2866);
DFFARX1 I_29686 (I80432,I2859,I507546,I507572,);
nand I_29687 (I507580,I507572,I80447);
DFFARX1 I_29688 (I80444,I2859,I507546,I507606,);
DFFARX1 I_29689 (I507606,I2859,I507546,I507623,);
not I_29690 (I507538,I507623);
not I_29691 (I507645,I80423);
nor I_29692 (I507662,I80423,I80429);
not I_29693 (I507679,I80435);
nand I_29694 (I507696,I507645,I507679);
nor I_29695 (I507713,I80435,I80423);
and I_29696 (I507517,I507713,I507580);
not I_29697 (I507744,I80441);
nand I_29698 (I507761,I507744,I80423);
nor I_29699 (I507778,I80441,I80426);
not I_29700 (I507795,I507778);
nand I_29701 (I507520,I507662,I507795);
DFFARX1 I_29702 (I507778,I2859,I507546,I507535,);
nor I_29703 (I507840,I80426,I80435);
nor I_29704 (I507857,I507840,I80429);
and I_29705 (I507874,I507857,I507761);
DFFARX1 I_29706 (I507874,I2859,I507546,I507532,);
nor I_29707 (I507529,I507840,I507696);
or I_29708 (I507526,I507778,I507840);
nor I_29709 (I507933,I80426,I80438);
DFFARX1 I_29710 (I507933,I2859,I507546,I507959,);
not I_29711 (I507967,I507959);
nand I_29712 (I507984,I507967,I507645);
nor I_29713 (I508001,I507984,I80429);
DFFARX1 I_29714 (I508001,I2859,I507546,I507514,);
nor I_29715 (I508032,I507967,I507696);
nor I_29716 (I507523,I507840,I508032);
not I_29717 (I508090,I2866);
DFFARX1 I_29718 (I542527,I2859,I508090,I508116,);
nand I_29719 (I508124,I508116,I542512);
DFFARX1 I_29720 (I542506,I2859,I508090,I508150,);
DFFARX1 I_29721 (I508150,I2859,I508090,I508167,);
not I_29722 (I508082,I508167);
not I_29723 (I508189,I542500);
nor I_29724 (I508206,I542500,I542521);
not I_29725 (I508223,I542509);
nand I_29726 (I508240,I508189,I508223);
nor I_29727 (I508257,I542509,I542500);
and I_29728 (I508061,I508257,I508124);
not I_29729 (I508288,I542518);
nand I_29730 (I508305,I508288,I542524);
nor I_29731 (I508322,I542518,I542515);
not I_29732 (I508339,I508322);
nand I_29733 (I508064,I508206,I508339);
DFFARX1 I_29734 (I508322,I2859,I508090,I508079,);
nor I_29735 (I508384,I542503,I542509);
nor I_29736 (I508401,I508384,I542521);
and I_29737 (I508418,I508401,I508305);
DFFARX1 I_29738 (I508418,I2859,I508090,I508076,);
nor I_29739 (I508073,I508384,I508240);
or I_29740 (I508070,I508322,I508384);
nor I_29741 (I508477,I542503,I542500);
DFFARX1 I_29742 (I508477,I2859,I508090,I508503,);
not I_29743 (I508511,I508503);
nand I_29744 (I508528,I508511,I508189);
nor I_29745 (I508545,I508528,I542521);
DFFARX1 I_29746 (I508545,I2859,I508090,I508058,);
nor I_29747 (I508576,I508511,I508240);
nor I_29748 (I508067,I508384,I508576);
not I_29749 (I508634,I2866);
DFFARX1 I_29750 (I480712,I2859,I508634,I508660,);
nand I_29751 (I508668,I508660,I480691);
DFFARX1 I_29752 (I480688,I2859,I508634,I508694,);
DFFARX1 I_29753 (I508694,I2859,I508634,I508711,);
not I_29754 (I508626,I508711);
not I_29755 (I508733,I480700);
nor I_29756 (I508750,I480700,I480709);
not I_29757 (I508767,I480697);
nand I_29758 (I508784,I508733,I508767);
nor I_29759 (I508801,I480697,I480700);
and I_29760 (I508605,I508801,I508668);
not I_29761 (I508832,I480706);
nand I_29762 (I508849,I508832,I480703);
nor I_29763 (I508866,I480706,I480688);
not I_29764 (I508883,I508866);
nand I_29765 (I508608,I508750,I508883);
DFFARX1 I_29766 (I508866,I2859,I508634,I508623,);
nor I_29767 (I508928,I480691,I480697);
nor I_29768 (I508945,I508928,I480709);
and I_29769 (I508962,I508945,I508849);
DFFARX1 I_29770 (I508962,I2859,I508634,I508620,);
nor I_29771 (I508617,I508928,I508784);
or I_29772 (I508614,I508866,I508928);
nor I_29773 (I509021,I480691,I480694);
DFFARX1 I_29774 (I509021,I2859,I508634,I509047,);
not I_29775 (I509055,I509047);
nand I_29776 (I509072,I509055,I508733);
nor I_29777 (I509089,I509072,I480709);
DFFARX1 I_29778 (I509089,I2859,I508634,I508602,);
nor I_29779 (I509120,I509055,I508784);
nor I_29780 (I508611,I508928,I509120);
not I_29781 (I509178,I2866);
DFFARX1 I_29782 (I39457,I2859,I509178,I509204,);
nand I_29783 (I509212,I509204,I39439);
DFFARX1 I_29784 (I39436,I2859,I509178,I509238,);
DFFARX1 I_29785 (I509238,I2859,I509178,I509255,);
not I_29786 (I509170,I509255);
not I_29787 (I509277,I39454);
nor I_29788 (I509294,I39454,I39448);
not I_29789 (I509311,I39436);
nand I_29790 (I509328,I509277,I509311);
nor I_29791 (I509345,I39436,I39454);
and I_29792 (I509149,I509345,I509212);
not I_29793 (I509376,I39445);
nand I_29794 (I509393,I509376,I39451);
nor I_29795 (I509410,I39445,I39439);
not I_29796 (I509427,I509410);
nand I_29797 (I509152,I509294,I509427);
DFFARX1 I_29798 (I509410,I2859,I509178,I509167,);
nor I_29799 (I509472,I39442,I39436);
nor I_29800 (I509489,I509472,I39448);
and I_29801 (I509506,I509489,I509393);
DFFARX1 I_29802 (I509506,I2859,I509178,I509164,);
nor I_29803 (I509161,I509472,I509328);
or I_29804 (I509158,I509410,I509472);
nor I_29805 (I509565,I39442,I39460);
DFFARX1 I_29806 (I509565,I2859,I509178,I509591,);
not I_29807 (I509599,I509591);
nand I_29808 (I509616,I509599,I509277);
nor I_29809 (I509633,I509616,I39448);
DFFARX1 I_29810 (I509633,I2859,I509178,I509146,);
nor I_29811 (I509664,I509599,I509328);
nor I_29812 (I509155,I509472,I509664);
not I_29813 (I509722,I2866);
DFFARX1 I_29814 (I560377,I2859,I509722,I509748,);
nand I_29815 (I509756,I509748,I560362);
DFFARX1 I_29816 (I560356,I2859,I509722,I509782,);
DFFARX1 I_29817 (I509782,I2859,I509722,I509799,);
not I_29818 (I509714,I509799);
not I_29819 (I509821,I560350);
nor I_29820 (I509838,I560350,I560371);
not I_29821 (I509855,I560359);
nand I_29822 (I509872,I509821,I509855);
nor I_29823 (I509889,I560359,I560350);
and I_29824 (I509693,I509889,I509756);
not I_29825 (I509920,I560368);
nand I_29826 (I509937,I509920,I560374);
nor I_29827 (I509954,I560368,I560365);
not I_29828 (I509971,I509954);
nand I_29829 (I509696,I509838,I509971);
DFFARX1 I_29830 (I509954,I2859,I509722,I509711,);
nor I_29831 (I510016,I560353,I560359);
nor I_29832 (I510033,I510016,I560371);
and I_29833 (I510050,I510033,I509937);
DFFARX1 I_29834 (I510050,I2859,I509722,I509708,);
nor I_29835 (I509705,I510016,I509872);
or I_29836 (I509702,I509954,I510016);
nor I_29837 (I510109,I560353,I560350);
DFFARX1 I_29838 (I510109,I2859,I509722,I510135,);
not I_29839 (I510143,I510135);
nand I_29840 (I510160,I510143,I509821);
nor I_29841 (I510177,I510160,I560371);
DFFARX1 I_29842 (I510177,I2859,I509722,I509690,);
nor I_29843 (I510208,I510143,I509872);
nor I_29844 (I509699,I510016,I510208);
not I_29845 (I510266,I2866);
DFFARX1 I_29846 (I427581,I2859,I510266,I510292,);
nand I_29847 (I510300,I510292,I427569);
DFFARX1 I_29848 (I427563,I2859,I510266,I510326,);
DFFARX1 I_29849 (I510326,I2859,I510266,I510343,);
not I_29850 (I510258,I510343);
not I_29851 (I510365,I427563);
nor I_29852 (I510382,I427563,I427575);
not I_29853 (I510399,I427572);
nand I_29854 (I510416,I510365,I510399);
nor I_29855 (I510433,I427572,I427563);
and I_29856 (I510237,I510433,I510300);
not I_29857 (I510464,I427566);
nand I_29858 (I510481,I510464,I427578);
nor I_29859 (I510498,I427566,I427584);
not I_29860 (I510515,I510498);
nand I_29861 (I510240,I510382,I510515);
DFFARX1 I_29862 (I510498,I2859,I510266,I510255,);
nor I_29863 (I510560,I427569,I427572);
nor I_29864 (I510577,I510560,I427575);
and I_29865 (I510594,I510577,I510481);
DFFARX1 I_29866 (I510594,I2859,I510266,I510252,);
nor I_29867 (I510249,I510560,I510416);
or I_29868 (I510246,I510498,I510560);
nor I_29869 (I510653,I427569,I427566);
DFFARX1 I_29870 (I510653,I2859,I510266,I510679,);
not I_29871 (I510687,I510679);
nand I_29872 (I510704,I510687,I510365);
nor I_29873 (I510721,I510704,I427575);
DFFARX1 I_29874 (I510721,I2859,I510266,I510234,);
nor I_29875 (I510752,I510687,I510416);
nor I_29876 (I510243,I510560,I510752);
not I_29877 (I510810,I2866);
DFFARX1 I_29878 (I185779,I2859,I510810,I510836,);
nand I_29879 (I510844,I510836,I185776);
DFFARX1 I_29880 (I185755,I2859,I510810,I510870,);
DFFARX1 I_29881 (I510870,I2859,I510810,I510887,);
not I_29882 (I510802,I510887);
not I_29883 (I510909,I185770);
nor I_29884 (I510926,I185770,I185773);
not I_29885 (I510943,I185764);
nand I_29886 (I510960,I510909,I510943);
nor I_29887 (I510977,I185764,I185770);
and I_29888 (I510781,I510977,I510844);
not I_29889 (I511008,I185761);
nand I_29890 (I511025,I511008,I185782);
nor I_29891 (I511042,I185761,I185758);
not I_29892 (I511059,I511042);
nand I_29893 (I510784,I510926,I511059);
DFFARX1 I_29894 (I511042,I2859,I510810,I510799,);
nor I_29895 (I511104,I185767,I185764);
nor I_29896 (I511121,I511104,I185773);
and I_29897 (I511138,I511121,I511025);
DFFARX1 I_29898 (I511138,I2859,I510810,I510796,);
nor I_29899 (I510793,I511104,I510960);
or I_29900 (I510790,I511042,I511104);
nor I_29901 (I511197,I185767,I185755);
DFFARX1 I_29902 (I511197,I2859,I510810,I511223,);
not I_29903 (I511231,I511223);
nand I_29904 (I511248,I511231,I510909);
nor I_29905 (I511265,I511248,I185773);
DFFARX1 I_29906 (I511265,I2859,I510810,I510778,);
nor I_29907 (I511296,I511231,I510960);
nor I_29908 (I510787,I511104,I511296);
not I_29909 (I511354,I2866);
DFFARX1 I_29910 (I448344,I2859,I511354,I511380,);
nand I_29911 (I511388,I511380,I448323);
DFFARX1 I_29912 (I448320,I2859,I511354,I511414,);
DFFARX1 I_29913 (I511414,I2859,I511354,I511431,);
not I_29914 (I511346,I511431);
not I_29915 (I511453,I448332);
nor I_29916 (I511470,I448332,I448341);
not I_29917 (I511487,I448329);
nand I_29918 (I511504,I511453,I511487);
nor I_29919 (I511521,I448329,I448332);
and I_29920 (I511325,I511521,I511388);
not I_29921 (I511552,I448338);
nand I_29922 (I511569,I511552,I448335);
nor I_29923 (I511586,I448338,I448320);
not I_29924 (I511603,I511586);
nand I_29925 (I511328,I511470,I511603);
DFFARX1 I_29926 (I511586,I2859,I511354,I511343,);
nor I_29927 (I511648,I448323,I448329);
nor I_29928 (I511665,I511648,I448341);
and I_29929 (I511682,I511665,I511569);
DFFARX1 I_29930 (I511682,I2859,I511354,I511340,);
nor I_29931 (I511337,I511648,I511504);
or I_29932 (I511334,I511586,I511648);
nor I_29933 (I511741,I448323,I448326);
DFFARX1 I_29934 (I511741,I2859,I511354,I511767,);
not I_29935 (I511775,I511767);
nand I_29936 (I511792,I511775,I511453);
nor I_29937 (I511809,I511792,I448341);
DFFARX1 I_29938 (I511809,I2859,I511354,I511322,);
nor I_29939 (I511840,I511775,I511504);
nor I_29940 (I511331,I511648,I511840);
not I_29941 (I511898,I2866);
DFFARX1 I_29942 (I498052,I2859,I511898,I511924,);
nand I_29943 (I511932,I511924,I498031);
DFFARX1 I_29944 (I498028,I2859,I511898,I511958,);
DFFARX1 I_29945 (I511958,I2859,I511898,I511975,);
not I_29946 (I511890,I511975);
not I_29947 (I511997,I498040);
nor I_29948 (I512014,I498040,I498049);
not I_29949 (I512031,I498037);
nand I_29950 (I512048,I511997,I512031);
nor I_29951 (I512065,I498037,I498040);
and I_29952 (I511869,I512065,I511932);
not I_29953 (I512096,I498046);
nand I_29954 (I512113,I512096,I498043);
nor I_29955 (I512130,I498046,I498028);
not I_29956 (I512147,I512130);
nand I_29957 (I511872,I512014,I512147);
DFFARX1 I_29958 (I512130,I2859,I511898,I511887,);
nor I_29959 (I512192,I498031,I498037);
nor I_29960 (I512209,I512192,I498049);
and I_29961 (I512226,I512209,I512113);
DFFARX1 I_29962 (I512226,I2859,I511898,I511884,);
nor I_29963 (I511881,I512192,I512048);
or I_29964 (I511878,I512130,I512192);
nor I_29965 (I512285,I498031,I498034);
DFFARX1 I_29966 (I512285,I2859,I511898,I512311,);
not I_29967 (I512319,I512311);
nand I_29968 (I512336,I512319,I511997);
nor I_29969 (I512353,I512336,I498049);
DFFARX1 I_29970 (I512353,I2859,I511898,I511866,);
nor I_29971 (I512384,I512319,I512048);
nor I_29972 (I511875,I512192,I512384);
not I_29973 (I512442,I2866);
DFFARX1 I_29974 (I9933,I2859,I512442,I512468,);
nand I_29975 (I512476,I512468,I9927);
DFFARX1 I_29976 (I9948,I2859,I512442,I512502,);
DFFARX1 I_29977 (I512502,I2859,I512442,I512519,);
not I_29978 (I512434,I512519);
not I_29979 (I512541,I9936);
nor I_29980 (I512558,I9936,I9945);
not I_29981 (I512575,I9924);
nand I_29982 (I512592,I512541,I512575);
nor I_29983 (I512609,I9924,I9936);
and I_29984 (I512413,I512609,I512476);
not I_29985 (I512640,I9942);
nand I_29986 (I512657,I512640,I9930);
nor I_29987 (I512674,I9942,I9924);
not I_29988 (I512691,I512674);
nand I_29989 (I512416,I512558,I512691);
DFFARX1 I_29990 (I512674,I2859,I512442,I512431,);
nor I_29991 (I512736,I9927,I9924);
nor I_29992 (I512753,I512736,I9945);
and I_29993 (I512770,I512753,I512657);
DFFARX1 I_29994 (I512770,I2859,I512442,I512428,);
nor I_29995 (I512425,I512736,I512592);
or I_29996 (I512422,I512674,I512736);
nor I_29997 (I512829,I9927,I9939);
DFFARX1 I_29998 (I512829,I2859,I512442,I512855,);
not I_29999 (I512863,I512855);
nand I_30000 (I512880,I512863,I512541);
nor I_30001 (I512897,I512880,I9945);
DFFARX1 I_30002 (I512897,I2859,I512442,I512410,);
nor I_30003 (I512928,I512863,I512592);
nor I_30004 (I512419,I512736,I512928);
not I_30005 (I512986,I2866);
DFFARX1 I_30006 (I217273,I2859,I512986,I513012,);
nand I_30007 (I513020,I513012,I217297);
DFFARX1 I_30008 (I217276,I2859,I512986,I513046,);
DFFARX1 I_30009 (I513046,I2859,I512986,I513063,);
not I_30010 (I512978,I513063);
not I_30011 (I513085,I217279);
nor I_30012 (I513102,I217279,I217294);
not I_30013 (I513119,I217285);
nand I_30014 (I513136,I513085,I513119);
nor I_30015 (I513153,I217285,I217279);
and I_30016 (I512957,I513153,I513020);
not I_30017 (I513184,I217282);
nand I_30018 (I513201,I513184,I217276);
nor I_30019 (I513218,I217282,I217291);
not I_30020 (I513235,I513218);
nand I_30021 (I512960,I513102,I513235);
DFFARX1 I_30022 (I513218,I2859,I512986,I512975,);
nor I_30023 (I513280,I217288,I217285);
nor I_30024 (I513297,I513280,I217294);
and I_30025 (I513314,I513297,I513201);
DFFARX1 I_30026 (I513314,I2859,I512986,I512972,);
nor I_30027 (I512969,I513280,I513136);
or I_30028 (I512966,I513218,I513280);
nor I_30029 (I513373,I217288,I217273);
DFFARX1 I_30030 (I513373,I2859,I512986,I513399,);
not I_30031 (I513407,I513399);
nand I_30032 (I513424,I513407,I513085);
nor I_30033 (I513441,I513424,I217294);
DFFARX1 I_30034 (I513441,I2859,I512986,I512954,);
nor I_30035 (I513472,I513407,I513136);
nor I_30036 (I512963,I513280,I513472);
not I_30037 (I513530,I2866);
DFFARX1 I_30038 (I521701,I2859,I513530,I513556,);
nand I_30039 (I513564,I513556,I521710);
DFFARX1 I_30040 (I521713,I2859,I513530,I513590,);
DFFARX1 I_30041 (I513590,I2859,I513530,I513607,);
not I_30042 (I513522,I513607);
not I_30043 (I513629,I521707);
nor I_30044 (I513646,I521707,I521704);
not I_30045 (I513663,I521698);
nand I_30046 (I513680,I513629,I513663);
nor I_30047 (I513697,I521698,I521707);
and I_30048 (I513501,I513697,I513564);
not I_30049 (I513728,I521695);
nand I_30050 (I513745,I513728,I521692);
nor I_30051 (I513762,I521695,I521692);
not I_30052 (I513779,I513762);
nand I_30053 (I513504,I513646,I513779);
DFFARX1 I_30054 (I513762,I2859,I513530,I513519,);
nor I_30055 (I513824,I521695,I521698);
nor I_30056 (I513841,I513824,I521704);
and I_30057 (I513858,I513841,I513745);
DFFARX1 I_30058 (I513858,I2859,I513530,I513516,);
nor I_30059 (I513513,I513824,I513680);
or I_30060 (I513510,I513762,I513824);
nor I_30061 (I513917,I521695,I521716);
DFFARX1 I_30062 (I513917,I2859,I513530,I513943,);
not I_30063 (I513951,I513943);
nand I_30064 (I513968,I513951,I513629);
nor I_30065 (I513985,I513968,I521704);
DFFARX1 I_30066 (I513985,I2859,I513530,I513498,);
nor I_30067 (I514016,I513951,I513680);
nor I_30068 (I513507,I513824,I514016);
not I_30069 (I514074,I2866);
DFFARX1 I_30070 (I232679,I2859,I514074,I514100,);
nand I_30071 (I514108,I514100,I232667);
DFFARX1 I_30072 (I232673,I2859,I514074,I514134,);
DFFARX1 I_30073 (I514134,I2859,I514074,I514151,);
not I_30074 (I514066,I514151);
not I_30075 (I514173,I232658);
nor I_30076 (I514190,I232658,I232670);
not I_30077 (I514207,I232661);
nand I_30078 (I514224,I514173,I514207);
nor I_30079 (I514241,I232661,I232658);
and I_30080 (I514045,I514241,I514108);
not I_30081 (I514272,I232676);
nand I_30082 (I514289,I514272,I232658);
nor I_30083 (I514306,I232676,I232682);
not I_30084 (I514323,I514306);
nand I_30085 (I514048,I514190,I514323);
DFFARX1 I_30086 (I514306,I2859,I514074,I514063,);
nor I_30087 (I514368,I232664,I232661);
nor I_30088 (I514385,I514368,I232670);
and I_30089 (I514402,I514385,I514289);
DFFARX1 I_30090 (I514402,I2859,I514074,I514060,);
nor I_30091 (I514057,I514368,I514224);
or I_30092 (I514054,I514306,I514368);
nor I_30093 (I514461,I232664,I232661);
DFFARX1 I_30094 (I514461,I2859,I514074,I514487,);
not I_30095 (I514495,I514487);
nand I_30096 (I514512,I514495,I514173);
nor I_30097 (I514529,I514512,I232670);
DFFARX1 I_30098 (I514529,I2859,I514074,I514042,);
nor I_30099 (I514560,I514495,I514224);
nor I_30100 (I514051,I514368,I514560);
not I_30101 (I514618,I2866);
DFFARX1 I_30102 (I24701,I2859,I514618,I514644,);
nand I_30103 (I514652,I514644,I24683);
DFFARX1 I_30104 (I24680,I2859,I514618,I514678,);
DFFARX1 I_30105 (I514678,I2859,I514618,I514695,);
not I_30106 (I514610,I514695);
not I_30107 (I514717,I24698);
nor I_30108 (I514734,I24698,I24692);
not I_30109 (I514751,I24680);
nand I_30110 (I514768,I514717,I514751);
nor I_30111 (I514785,I24680,I24698);
and I_30112 (I514589,I514785,I514652);
not I_30113 (I514816,I24689);
nand I_30114 (I514833,I514816,I24695);
nor I_30115 (I514850,I24689,I24683);
not I_30116 (I514867,I514850);
nand I_30117 (I514592,I514734,I514867);
DFFARX1 I_30118 (I514850,I2859,I514618,I514607,);
nor I_30119 (I514912,I24686,I24680);
nor I_30120 (I514929,I514912,I24692);
and I_30121 (I514946,I514929,I514833);
DFFARX1 I_30122 (I514946,I2859,I514618,I514604,);
nor I_30123 (I514601,I514912,I514768);
or I_30124 (I514598,I514850,I514912);
nor I_30125 (I515005,I24686,I24704);
DFFARX1 I_30126 (I515005,I2859,I514618,I515031,);
not I_30127 (I515039,I515031);
nand I_30128 (I515056,I515039,I514717);
nor I_30129 (I515073,I515056,I24692);
DFFARX1 I_30130 (I515073,I2859,I514618,I514586,);
nor I_30131 (I515104,I515039,I514768);
nor I_30132 (I514595,I514912,I515104);
not I_30133 (I515162,I2866);
DFFARX1 I_30134 (I389959,I2859,I515162,I515188,);
nand I_30135 (I515196,I515188,I389959);
DFFARX1 I_30136 (I389971,I2859,I515162,I515222,);
DFFARX1 I_30137 (I515222,I2859,I515162,I515239,);
not I_30138 (I515154,I515239);
not I_30139 (I515261,I389965);
nor I_30140 (I515278,I389965,I389986);
not I_30141 (I515295,I389974);
nand I_30142 (I515312,I515261,I515295);
nor I_30143 (I515329,I389974,I389965);
and I_30144 (I515133,I515329,I515196);
not I_30145 (I515360,I389968);
nand I_30146 (I515377,I515360,I389983);
nor I_30147 (I515394,I389968,I389977);
not I_30148 (I515411,I515394);
nand I_30149 (I515136,I515278,I515411);
DFFARX1 I_30150 (I515394,I2859,I515162,I515151,);
nor I_30151 (I515456,I389980,I389974);
nor I_30152 (I515473,I515456,I389986);
and I_30153 (I515490,I515473,I515377);
DFFARX1 I_30154 (I515490,I2859,I515162,I515148,);
nor I_30155 (I515145,I515456,I515312);
or I_30156 (I515142,I515394,I515456);
nor I_30157 (I515549,I389980,I389962);
DFFARX1 I_30158 (I515549,I2859,I515162,I515575,);
not I_30159 (I515583,I515575);
nand I_30160 (I515600,I515583,I515261);
nor I_30161 (I515617,I515600,I389986);
DFFARX1 I_30162 (I515617,I2859,I515162,I515130,);
nor I_30163 (I515648,I515583,I515312);
nor I_30164 (I515139,I515456,I515648);
not I_30165 (I515706,I2866);
DFFARX1 I_30166 (I9406,I2859,I515706,I515732,);
nand I_30167 (I515740,I515732,I9400);
DFFARX1 I_30168 (I9421,I2859,I515706,I515766,);
DFFARX1 I_30169 (I515766,I2859,I515706,I515783,);
not I_30170 (I515698,I515783);
not I_30171 (I515805,I9409);
nor I_30172 (I515822,I9409,I9418);
not I_30173 (I515839,I9397);
nand I_30174 (I515856,I515805,I515839);
nor I_30175 (I515873,I9397,I9409);
and I_30176 (I515677,I515873,I515740);
not I_30177 (I515904,I9415);
nand I_30178 (I515921,I515904,I9403);
nor I_30179 (I515938,I9415,I9397);
not I_30180 (I515955,I515938);
nand I_30181 (I515680,I515822,I515955);
DFFARX1 I_30182 (I515938,I2859,I515706,I515695,);
nor I_30183 (I516000,I9400,I9397);
nor I_30184 (I516017,I516000,I9418);
and I_30185 (I516034,I516017,I515921);
DFFARX1 I_30186 (I516034,I2859,I515706,I515692,);
nor I_30187 (I515689,I516000,I515856);
or I_30188 (I515686,I515938,I516000);
nor I_30189 (I516093,I9400,I9412);
DFFARX1 I_30190 (I516093,I2859,I515706,I516119,);
not I_30191 (I516127,I516119);
nand I_30192 (I516144,I516127,I515805);
nor I_30193 (I516161,I516144,I9418);
DFFARX1 I_30194 (I516161,I2859,I515706,I515674,);
nor I_30195 (I516192,I516127,I515856);
nor I_30196 (I515683,I516000,I516192);
not I_30197 (I516250,I2866);
DFFARX1 I_30198 (I282369,I2859,I516250,I516276,);
nand I_30199 (I516284,I516276,I282384);
DFFARX1 I_30200 (I282378,I2859,I516250,I516310,);
DFFARX1 I_30201 (I516310,I2859,I516250,I516327,);
not I_30202 (I516242,I516327);
not I_30203 (I516349,I282381);
nor I_30204 (I516366,I282381,I282387);
not I_30205 (I516383,I282369);
nand I_30206 (I516400,I516349,I516383);
nor I_30207 (I516417,I282369,I282381);
and I_30208 (I516221,I516417,I516284);
not I_30209 (I516448,I282366);
nand I_30210 (I516465,I516448,I282372);
nor I_30211 (I516482,I282366,I282366);
not I_30212 (I516499,I516482);
nand I_30213 (I516224,I516366,I516499);
DFFARX1 I_30214 (I516482,I2859,I516250,I516239,);
nor I_30215 (I516544,I282375,I282369);
nor I_30216 (I516561,I516544,I282387);
and I_30217 (I516578,I516561,I516465);
DFFARX1 I_30218 (I516578,I2859,I516250,I516236,);
nor I_30219 (I516233,I516544,I516400);
or I_30220 (I516230,I516482,I516544);
nor I_30221 (I516637,I282375,I282390);
DFFARX1 I_30222 (I516637,I2859,I516250,I516663,);
not I_30223 (I516671,I516663);
nand I_30224 (I516688,I516671,I516349);
nor I_30225 (I516705,I516688,I282387);
DFFARX1 I_30226 (I516705,I2859,I516250,I516218,);
nor I_30227 (I516736,I516671,I516400);
nor I_30228 (I516227,I516544,I516736);
not I_30229 (I516794,I2866);
DFFARX1 I_30230 (I25228,I2859,I516794,I516820,);
nand I_30231 (I516828,I516820,I25210);
DFFARX1 I_30232 (I25207,I2859,I516794,I516854,);
DFFARX1 I_30233 (I516854,I2859,I516794,I516871,);
not I_30234 (I516786,I516871);
not I_30235 (I516893,I25225);
nor I_30236 (I516910,I25225,I25219);
not I_30237 (I516927,I25207);
nand I_30238 (I516944,I516893,I516927);
nor I_30239 (I516961,I25207,I25225);
and I_30240 (I516765,I516961,I516828);
not I_30241 (I516992,I25216);
nand I_30242 (I517009,I516992,I25222);
nor I_30243 (I517026,I25216,I25210);
not I_30244 (I517043,I517026);
nand I_30245 (I516768,I516910,I517043);
DFFARX1 I_30246 (I517026,I2859,I516794,I516783,);
nor I_30247 (I517088,I25213,I25207);
nor I_30248 (I517105,I517088,I25219);
and I_30249 (I517122,I517105,I517009);
DFFARX1 I_30250 (I517122,I2859,I516794,I516780,);
nor I_30251 (I516777,I517088,I516944);
or I_30252 (I516774,I517026,I517088);
nor I_30253 (I517181,I25213,I25231);
DFFARX1 I_30254 (I517181,I2859,I516794,I517207,);
not I_30255 (I517215,I517207);
nand I_30256 (I517232,I517215,I516893);
nor I_30257 (I517249,I517232,I25219);
DFFARX1 I_30258 (I517249,I2859,I516794,I516762,);
nor I_30259 (I517280,I517215,I516944);
nor I_30260 (I516771,I517088,I517280);
not I_30261 (I517338,I2866);
DFFARX1 I_30262 (I66747,I2859,I517338,I517364,);
nand I_30263 (I517372,I517364,I66762);
DFFARX1 I_30264 (I66759,I2859,I517338,I517398,);
DFFARX1 I_30265 (I517398,I2859,I517338,I517415,);
not I_30266 (I517330,I517415);
not I_30267 (I517437,I66738);
nor I_30268 (I517454,I66738,I66744);
not I_30269 (I517471,I66750);
nand I_30270 (I517488,I517437,I517471);
nor I_30271 (I517505,I66750,I66738);
and I_30272 (I517309,I517505,I517372);
not I_30273 (I517536,I66756);
nand I_30274 (I517553,I517536,I66738);
nor I_30275 (I517570,I66756,I66741);
not I_30276 (I517587,I517570);
nand I_30277 (I517312,I517454,I517587);
DFFARX1 I_30278 (I517570,I2859,I517338,I517327,);
nor I_30279 (I517632,I66741,I66750);
nor I_30280 (I517649,I517632,I66744);
and I_30281 (I517666,I517649,I517553);
DFFARX1 I_30282 (I517666,I2859,I517338,I517324,);
nor I_30283 (I517321,I517632,I517488);
or I_30284 (I517318,I517570,I517632);
nor I_30285 (I517725,I66741,I66753);
DFFARX1 I_30286 (I517725,I2859,I517338,I517751,);
not I_30287 (I517759,I517751);
nand I_30288 (I517776,I517759,I517437);
nor I_30289 (I517793,I517776,I66744);
DFFARX1 I_30290 (I517793,I2859,I517338,I517306,);
nor I_30291 (I517824,I517759,I517488);
nor I_30292 (I517315,I517632,I517824);
not I_30293 (I517882,I2866);
DFFARX1 I_30294 (I171635,I2859,I517882,I517908,);
nand I_30295 (I517916,I517908,I171632);
DFFARX1 I_30296 (I171611,I2859,I517882,I517942,);
DFFARX1 I_30297 (I517942,I2859,I517882,I517959,);
not I_30298 (I517874,I517959);
not I_30299 (I517981,I171626);
nor I_30300 (I517998,I171626,I171629);
not I_30301 (I518015,I171620);
nand I_30302 (I518032,I517981,I518015);
nor I_30303 (I518049,I171620,I171626);
and I_30304 (I517853,I518049,I517916);
not I_30305 (I518080,I171617);
nand I_30306 (I518097,I518080,I171638);
nor I_30307 (I518114,I171617,I171614);
not I_30308 (I518131,I518114);
nand I_30309 (I517856,I517998,I518131);
DFFARX1 I_30310 (I518114,I2859,I517882,I517871,);
nor I_30311 (I518176,I171623,I171620);
nor I_30312 (I518193,I518176,I171629);
and I_30313 (I518210,I518193,I518097);
DFFARX1 I_30314 (I518210,I2859,I517882,I517868,);
nor I_30315 (I517865,I518176,I518032);
or I_30316 (I517862,I518114,I518176);
nor I_30317 (I518269,I171623,I171611);
DFFARX1 I_30318 (I518269,I2859,I517882,I518295,);
not I_30319 (I518303,I518295);
nand I_30320 (I518320,I518303,I517981);
nor I_30321 (I518337,I518320,I171629);
DFFARX1 I_30322 (I518337,I2859,I517882,I517850,);
nor I_30323 (I518368,I518303,I518032);
nor I_30324 (I517859,I518176,I518368);
not I_30325 (I518426,I2866);
DFFARX1 I_30326 (I358481,I2859,I518426,I518452,);
nand I_30327 (I518460,I518452,I358475);
DFFARX1 I_30328 (I358478,I2859,I518426,I518486,);
DFFARX1 I_30329 (I518486,I2859,I518426,I518503,);
not I_30330 (I518418,I518503);
not I_30331 (I518525,I358484);
nor I_30332 (I518542,I358484,I358478);
not I_30333 (I518559,I358487);
nand I_30334 (I518576,I518525,I518559);
nor I_30335 (I518593,I358487,I358484);
and I_30336 (I518397,I518593,I518460);
not I_30337 (I518624,I358496);
nand I_30338 (I518641,I518624,I358490);
nor I_30339 (I518658,I358496,I358493);
not I_30340 (I518675,I518658);
nand I_30341 (I518400,I518542,I518675);
DFFARX1 I_30342 (I518658,I2859,I518426,I518415,);
nor I_30343 (I518720,I358475,I358487);
nor I_30344 (I518737,I518720,I358478);
and I_30345 (I518754,I518737,I518641);
DFFARX1 I_30346 (I518754,I2859,I518426,I518412,);
nor I_30347 (I518409,I518720,I518576);
or I_30348 (I518406,I518658,I518720);
nor I_30349 (I518813,I358475,I358481);
DFFARX1 I_30350 (I518813,I2859,I518426,I518839,);
not I_30351 (I518847,I518839);
nand I_30352 (I518864,I518847,I518525);
nor I_30353 (I518881,I518864,I358478);
DFFARX1 I_30354 (I518881,I2859,I518426,I518394,);
nor I_30355 (I518912,I518847,I518576);
nor I_30356 (I518403,I518720,I518912);
not I_30357 (I518970,I2866);
DFFARX1 I_30358 (I554427,I2859,I518970,I518996,);
nand I_30359 (I519004,I518996,I554412);
DFFARX1 I_30360 (I554406,I2859,I518970,I519030,);
DFFARX1 I_30361 (I519030,I2859,I518970,I519047,);
not I_30362 (I518962,I519047);
not I_30363 (I519069,I554400);
nor I_30364 (I519086,I554400,I554421);
not I_30365 (I519103,I554409);
nand I_30366 (I519120,I519069,I519103);
nor I_30367 (I519137,I554409,I554400);
and I_30368 (I518941,I519137,I519004);
not I_30369 (I519168,I554418);
nand I_30370 (I519185,I519168,I554424);
nor I_30371 (I519202,I554418,I554415);
not I_30372 (I519219,I519202);
nand I_30373 (I518944,I519086,I519219);
DFFARX1 I_30374 (I519202,I2859,I518970,I518959,);
nor I_30375 (I519264,I554403,I554409);
nor I_30376 (I519281,I519264,I554421);
and I_30377 (I519298,I519281,I519185);
DFFARX1 I_30378 (I519298,I2859,I518970,I518956,);
nor I_30379 (I518953,I519264,I519120);
or I_30380 (I518950,I519202,I519264);
nor I_30381 (I519357,I554403,I554400);
DFFARX1 I_30382 (I519357,I2859,I518970,I519383,);
not I_30383 (I519391,I519383);
nand I_30384 (I519408,I519391,I519069);
nor I_30385 (I519425,I519408,I554421);
DFFARX1 I_30386 (I519425,I2859,I518970,I518938,);
nor I_30387 (I519456,I519391,I519120);
nor I_30388 (I518947,I519264,I519456);
not I_30389 (I519514,I2866);
DFFARX1 I_30390 (I119790,I2859,I519514,I519540,);
nand I_30391 (I519548,I519540,I119793);
DFFARX1 I_30392 (I119787,I2859,I519514,I519574,);
DFFARX1 I_30393 (I519574,I2859,I519514,I519591,);
not I_30394 (I519506,I519591);
not I_30395 (I519613,I119796);
nor I_30396 (I519630,I119796,I119781);
not I_30397 (I519647,I119805);
nand I_30398 (I519664,I519613,I519647);
nor I_30399 (I519681,I119805,I119796);
and I_30400 (I519485,I519681,I519548);
not I_30401 (I519712,I119784);
nand I_30402 (I519729,I519712,I119802);
nor I_30403 (I519746,I119784,I119778);
not I_30404 (I519763,I519746);
nand I_30405 (I519488,I519630,I519763);
DFFARX1 I_30406 (I519746,I2859,I519514,I519503,);
nor I_30407 (I519808,I119799,I119805);
nor I_30408 (I519825,I519808,I119781);
and I_30409 (I519842,I519825,I519729);
DFFARX1 I_30410 (I519842,I2859,I519514,I519500,);
nor I_30411 (I519497,I519808,I519664);
or I_30412 (I519494,I519746,I519808);
nor I_30413 (I519901,I119799,I119778);
DFFARX1 I_30414 (I519901,I2859,I519514,I519927,);
not I_30415 (I519935,I519927);
nand I_30416 (I519952,I519935,I519613);
nor I_30417 (I519969,I519952,I119781);
DFFARX1 I_30418 (I519969,I2859,I519514,I519482,);
nor I_30419 (I520000,I519935,I519664);
nor I_30420 (I519491,I519808,I520000);
not I_30421 (I520058,I2866);
DFFARX1 I_30422 (I239615,I2859,I520058,I520084,);
nand I_30423 (I520092,I520084,I239603);
DFFARX1 I_30424 (I239609,I2859,I520058,I520118,);
DFFARX1 I_30425 (I520118,I2859,I520058,I520135,);
not I_30426 (I520050,I520135);
not I_30427 (I520157,I239594);
nor I_30428 (I520174,I239594,I239606);
not I_30429 (I520191,I239597);
nand I_30430 (I520208,I520157,I520191);
nor I_30431 (I520225,I239597,I239594);
and I_30432 (I520029,I520225,I520092);
not I_30433 (I520256,I239612);
nand I_30434 (I520273,I520256,I239594);
nor I_30435 (I520290,I239612,I239618);
not I_30436 (I520307,I520290);
nand I_30437 (I520032,I520174,I520307);
DFFARX1 I_30438 (I520290,I2859,I520058,I520047,);
nor I_30439 (I520352,I239600,I239597);
nor I_30440 (I520369,I520352,I239606);
and I_30441 (I520386,I520369,I520273);
DFFARX1 I_30442 (I520386,I2859,I520058,I520044,);
nor I_30443 (I520041,I520352,I520208);
or I_30444 (I520038,I520290,I520352);
nor I_30445 (I520445,I239600,I239597);
DFFARX1 I_30446 (I520445,I2859,I520058,I520471,);
not I_30447 (I520479,I520471);
nand I_30448 (I520496,I520479,I520157);
nor I_30449 (I520513,I520496,I239606);
DFFARX1 I_30450 (I520513,I2859,I520058,I520026,);
nor I_30451 (I520544,I520479,I520208);
nor I_30452 (I520035,I520352,I520544);
not I_30453 (I520602,I2866);
DFFARX1 I_30454 (I375872,I2859,I520602,I520628,);
nand I_30455 (I520636,I520628,I375866);
DFFARX1 I_30456 (I375869,I2859,I520602,I520662,);
DFFARX1 I_30457 (I520662,I2859,I520602,I520679,);
not I_30458 (I520594,I520679);
not I_30459 (I520701,I375875);
nor I_30460 (I520718,I375875,I375869);
not I_30461 (I520735,I375878);
nand I_30462 (I520752,I520701,I520735);
nor I_30463 (I520769,I375878,I375875);
and I_30464 (I520573,I520769,I520636);
not I_30465 (I520800,I375887);
nand I_30466 (I520817,I520800,I375881);
nor I_30467 (I520834,I375887,I375884);
not I_30468 (I520851,I520834);
nand I_30469 (I520576,I520718,I520851);
DFFARX1 I_30470 (I520834,I2859,I520602,I520591,);
nor I_30471 (I520896,I375866,I375878);
nor I_30472 (I520913,I520896,I375869);
and I_30473 (I520930,I520913,I520817);
DFFARX1 I_30474 (I520930,I2859,I520602,I520588,);
nor I_30475 (I520585,I520896,I520752);
or I_30476 (I520582,I520834,I520896);
nor I_30477 (I520989,I375866,I375872);
DFFARX1 I_30478 (I520989,I2859,I520602,I521015,);
not I_30479 (I521023,I521015);
nand I_30480 (I521040,I521023,I520701);
nor I_30481 (I521057,I521040,I375869);
DFFARX1 I_30482 (I521057,I2859,I520602,I520570,);
nor I_30483 (I521088,I521023,I520752);
nor I_30484 (I520579,I520896,I521088);
not I_30485 (I521146,I2866);
DFFARX1 I_30486 (I550854,I2859,I521146,I521172,);
nand I_30487 (I521180,I521172,I550845);
not I_30488 (I521197,I521180);
DFFARX1 I_30489 (I550830,I2859,I521146,I521223,);
not I_30490 (I521231,I521223);
not I_30491 (I521248,I550833);
or I_30492 (I521265,I550842,I550833);
nor I_30493 (I521282,I550842,I550833);
or I_30494 (I521299,I550839,I550842);
DFFARX1 I_30495 (I521299,I2859,I521146,I521138,);
not I_30496 (I521330,I550851);
nand I_30497 (I521347,I521330,I550830);
nand I_30498 (I521364,I521248,I521347);
and I_30499 (I521117,I521231,I521364);
nor I_30500 (I521395,I550851,I550836);
and I_30501 (I521412,I521231,I521395);
nor I_30502 (I521123,I521197,I521412);
DFFARX1 I_30503 (I521395,I2859,I521146,I521452,);
not I_30504 (I521460,I521452);
nor I_30505 (I521132,I521231,I521460);
or I_30506 (I521491,I521299,I550857);
nor I_30507 (I521508,I550857,I550839);
nand I_30508 (I521525,I521364,I521508);
nand I_30509 (I521542,I521491,I521525);
DFFARX1 I_30510 (I521542,I2859,I521146,I521135,);
nor I_30511 (I521573,I521508,I521265);
DFFARX1 I_30512 (I521573,I2859,I521146,I521114,);
nor I_30513 (I521604,I550857,I550848);
DFFARX1 I_30514 (I521604,I2859,I521146,I521630,);
DFFARX1 I_30515 (I521630,I2859,I521146,I521129,);
not I_30516 (I521652,I521630);
nand I_30517 (I521126,I521652,I521180);
nand I_30518 (I521120,I521652,I521282);
not I_30519 (I521724,I2866);
DFFARX1 I_30520 (I158255,I2859,I521724,I521750,);
nand I_30521 (I521758,I521750,I158276);
not I_30522 (I521775,I521758);
DFFARX1 I_30523 (I158270,I2859,I521724,I521801,);
not I_30524 (I521809,I521801);
not I_30525 (I521826,I158258);
or I_30526 (I521843,I158273,I158258);
nor I_30527 (I521860,I158273,I158258);
or I_30528 (I521877,I158264,I158273);
DFFARX1 I_30529 (I521877,I2859,I521724,I521716,);
not I_30530 (I521908,I158252);
nand I_30531 (I521925,I521908,I158249);
nand I_30532 (I521942,I521826,I521925);
and I_30533 (I521695,I521809,I521942);
nor I_30534 (I521973,I158252,I158261);
and I_30535 (I521990,I521809,I521973);
nor I_30536 (I521701,I521775,I521990);
DFFARX1 I_30537 (I521973,I2859,I521724,I522030,);
not I_30538 (I522038,I522030);
nor I_30539 (I521710,I521809,I522038);
or I_30540 (I522069,I521877,I158267);
nor I_30541 (I522086,I158267,I158264);
nand I_30542 (I522103,I521942,I522086);
nand I_30543 (I522120,I522069,I522103);
DFFARX1 I_30544 (I522120,I2859,I521724,I521713,);
nor I_30545 (I522151,I522086,I521843);
DFFARX1 I_30546 (I522151,I2859,I521724,I521692,);
nor I_30547 (I522182,I158267,I158249);
DFFARX1 I_30548 (I522182,I2859,I521724,I522208,);
DFFARX1 I_30549 (I522208,I2859,I521724,I521707,);
not I_30550 (I522230,I522208);
nand I_30551 (I521704,I522230,I521758);
nand I_30552 (I521698,I522230,I521860);
not I_30553 (I522302,I2866);
DFFARX1 I_30554 (I128216,I2859,I522302,I522328,);
nand I_30555 (I522336,I522328,I128237);
not I_30556 (I522353,I522336);
DFFARX1 I_30557 (I128231,I2859,I522302,I522379,);
not I_30558 (I522387,I522379);
not I_30559 (I522404,I128219);
or I_30560 (I522421,I128234,I128219);
nor I_30561 (I522438,I128234,I128219);
or I_30562 (I522455,I128225,I128234);
DFFARX1 I_30563 (I522455,I2859,I522302,I522294,);
not I_30564 (I522486,I128213);
nand I_30565 (I522503,I522486,I128210);
nand I_30566 (I522520,I522404,I522503);
and I_30567 (I522273,I522387,I522520);
nor I_30568 (I522551,I128213,I128222);
and I_30569 (I522568,I522387,I522551);
nor I_30570 (I522279,I522353,I522568);
DFFARX1 I_30571 (I522551,I2859,I522302,I522608,);
not I_30572 (I522616,I522608);
nor I_30573 (I522288,I522387,I522616);
or I_30574 (I522647,I522455,I128228);
nor I_30575 (I522664,I128228,I128225);
nand I_30576 (I522681,I522520,I522664);
nand I_30577 (I522698,I522647,I522681);
DFFARX1 I_30578 (I522698,I2859,I522302,I522291,);
nor I_30579 (I522729,I522664,I522421);
DFFARX1 I_30580 (I522729,I2859,I522302,I522270,);
nor I_30581 (I522760,I128228,I128210);
DFFARX1 I_30582 (I522760,I2859,I522302,I522786,);
DFFARX1 I_30583 (I522786,I2859,I522302,I522285,);
not I_30584 (I522808,I522786);
nand I_30585 (I522282,I522808,I522336);
nand I_30586 (I522276,I522808,I522438);
not I_30587 (I522880,I2866);
DFFARX1 I_30588 (I369018,I2859,I522880,I522906,);
nand I_30589 (I522914,I522906,I369018);
not I_30590 (I522931,I522914);
DFFARX1 I_30591 (I369024,I2859,I522880,I522957,);
not I_30592 (I522965,I522957);
not I_30593 (I522982,I369036);
or I_30594 (I522999,I369021,I369036);
nor I_30595 (I523016,I369021,I369036);
or I_30596 (I523033,I369015,I369021);
DFFARX1 I_30597 (I523033,I2859,I522880,I522872,);
not I_30598 (I523064,I369033);
nand I_30599 (I523081,I523064,I369027);
nand I_30600 (I523098,I522982,I523081);
and I_30601 (I522851,I522965,I523098);
nor I_30602 (I523129,I369033,I369015);
and I_30603 (I523146,I522965,I523129);
nor I_30604 (I522857,I522931,I523146);
DFFARX1 I_30605 (I523129,I2859,I522880,I523186,);
not I_30606 (I523194,I523186);
nor I_30607 (I522866,I522965,I523194);
or I_30608 (I523225,I523033,I369030);
nor I_30609 (I523242,I369030,I369015);
nand I_30610 (I523259,I523098,I523242);
nand I_30611 (I523276,I523225,I523259);
DFFARX1 I_30612 (I523276,I2859,I522880,I522869,);
nor I_30613 (I523307,I523242,I522999);
DFFARX1 I_30614 (I523307,I2859,I522880,I522848,);
nor I_30615 (I523338,I369030,I369021);
DFFARX1 I_30616 (I523338,I2859,I522880,I523364,);
DFFARX1 I_30617 (I523364,I2859,I522880,I522863,);
not I_30618 (I523386,I523364);
nand I_30619 (I522860,I523386,I522914);
nand I_30620 (I522854,I523386,I523016);
not I_30621 (I523458,I2866);
DFFARX1 I_30622 (I342668,I2859,I523458,I523484,);
nand I_30623 (I523492,I523484,I342668);
not I_30624 (I523509,I523492);
DFFARX1 I_30625 (I342674,I2859,I523458,I523535,);
not I_30626 (I523543,I523535);
not I_30627 (I523560,I342686);
or I_30628 (I523577,I342671,I342686);
nor I_30629 (I523594,I342671,I342686);
or I_30630 (I523611,I342665,I342671);
DFFARX1 I_30631 (I523611,I2859,I523458,I523450,);
not I_30632 (I523642,I342683);
nand I_30633 (I523659,I523642,I342677);
nand I_30634 (I523676,I523560,I523659);
and I_30635 (I523429,I523543,I523676);
nor I_30636 (I523707,I342683,I342665);
and I_30637 (I523724,I523543,I523707);
nor I_30638 (I523435,I523509,I523724);
DFFARX1 I_30639 (I523707,I2859,I523458,I523764,);
not I_30640 (I523772,I523764);
nor I_30641 (I523444,I523543,I523772);
or I_30642 (I523803,I523611,I342680);
nor I_30643 (I523820,I342680,I342665);
nand I_30644 (I523837,I523676,I523820);
nand I_30645 (I523854,I523803,I523837);
DFFARX1 I_30646 (I523854,I2859,I523458,I523447,);
nor I_30647 (I523885,I523820,I523577);
DFFARX1 I_30648 (I523885,I2859,I523458,I523426,);
nor I_30649 (I523916,I342680,I342671);
DFFARX1 I_30650 (I523916,I2859,I523458,I523942,);
DFFARX1 I_30651 (I523942,I2859,I523458,I523441,);
not I_30652 (I523964,I523942);
nand I_30653 (I523438,I523964,I523492);
nand I_30654 (I523432,I523964,I523594);
not I_30655 (I524036,I2866);
DFFARX1 I_30656 (I449494,I2859,I524036,I524062,);
nand I_30657 (I524070,I524062,I449479);
not I_30658 (I524087,I524070);
DFFARX1 I_30659 (I449482,I2859,I524036,I524113,);
not I_30660 (I524121,I524113);
not I_30661 (I524138,I449497);
or I_30662 (I524155,I449500,I449497);
nor I_30663 (I524172,I449500,I449497);
or I_30664 (I524189,I449476,I449500);
DFFARX1 I_30665 (I524189,I2859,I524036,I524028,);
not I_30666 (I524220,I449488);
nand I_30667 (I524237,I524220,I449491);
nand I_30668 (I524254,I524138,I524237);
and I_30669 (I524007,I524121,I524254);
nor I_30670 (I524285,I449488,I449485);
and I_30671 (I524302,I524121,I524285);
nor I_30672 (I524013,I524087,I524302);
DFFARX1 I_30673 (I524285,I2859,I524036,I524342,);
not I_30674 (I524350,I524342);
nor I_30675 (I524022,I524121,I524350);
or I_30676 (I524381,I524189,I449476);
nor I_30677 (I524398,I449476,I449476);
nand I_30678 (I524415,I524254,I524398);
nand I_30679 (I524432,I524381,I524415);
DFFARX1 I_30680 (I524432,I2859,I524036,I524025,);
nor I_30681 (I524463,I524398,I524155);
DFFARX1 I_30682 (I524463,I2859,I524036,I524004,);
nor I_30683 (I524494,I449476,I449479);
DFFARX1 I_30684 (I524494,I2859,I524036,I524520,);
DFFARX1 I_30685 (I524520,I2859,I524036,I524019,);
not I_30686 (I524542,I524520);
nand I_30687 (I524016,I524542,I524070);
nand I_30688 (I524010,I524542,I524172);
not I_30689 (I524614,I2866);
DFFARX1 I_30690 (I442719,I2859,I524614,I524640,);
nand I_30691 (I524648,I524640,I442716);
not I_30692 (I524665,I524648);
DFFARX1 I_30693 (I442716,I2859,I524614,I524691,);
not I_30694 (I524699,I524691);
not I_30695 (I524716,I442713);
or I_30696 (I524733,I442722,I442713);
nor I_30697 (I524750,I442722,I442713);
or I_30698 (I524767,I442725,I442722);
DFFARX1 I_30699 (I524767,I2859,I524614,I524606,);
not I_30700 (I524798,I442713);
nand I_30701 (I524815,I524798,I442710);
nand I_30702 (I524832,I524716,I524815);
and I_30703 (I524585,I524699,I524832);
nor I_30704 (I524863,I442713,I442728);
and I_30705 (I524880,I524699,I524863);
nor I_30706 (I524591,I524665,I524880);
DFFARX1 I_30707 (I524863,I2859,I524614,I524920,);
not I_30708 (I524928,I524920);
nor I_30709 (I524600,I524699,I524928);
or I_30710 (I524959,I524767,I442731);
nor I_30711 (I524976,I442731,I442725);
nand I_30712 (I524993,I524832,I524976);
nand I_30713 (I525010,I524959,I524993);
DFFARX1 I_30714 (I525010,I2859,I524614,I524603,);
nor I_30715 (I525041,I524976,I524733);
DFFARX1 I_30716 (I525041,I2859,I524614,I524582,);
nor I_30717 (I525072,I442731,I442710);
DFFARX1 I_30718 (I525072,I2859,I524614,I525098,);
DFFARX1 I_30719 (I525098,I2859,I524614,I524597,);
not I_30720 (I525120,I525098);
nand I_30721 (I524594,I525120,I524648);
nand I_30722 (I524588,I525120,I524750);
not I_30723 (I525192,I2866);
DFFARX1 I_30724 (I457586,I2859,I525192,I525218,);
nand I_30725 (I525226,I525218,I457571);
not I_30726 (I525243,I525226);
DFFARX1 I_30727 (I457574,I2859,I525192,I525269,);
not I_30728 (I525277,I525269);
not I_30729 (I525294,I457589);
or I_30730 (I525311,I457592,I457589);
nor I_30731 (I525328,I457592,I457589);
or I_30732 (I525345,I457568,I457592);
DFFARX1 I_30733 (I525345,I2859,I525192,I525184,);
not I_30734 (I525376,I457580);
nand I_30735 (I525393,I525376,I457583);
nand I_30736 (I525410,I525294,I525393);
and I_30737 (I525163,I525277,I525410);
nor I_30738 (I525441,I457580,I457577);
and I_30739 (I525458,I525277,I525441);
nor I_30740 (I525169,I525243,I525458);
DFFARX1 I_30741 (I525441,I2859,I525192,I525498,);
not I_30742 (I525506,I525498);
nor I_30743 (I525178,I525277,I525506);
or I_30744 (I525537,I525345,I457568);
nor I_30745 (I525554,I457568,I457568);
nand I_30746 (I525571,I525410,I525554);
nand I_30747 (I525588,I525537,I525571);
DFFARX1 I_30748 (I525588,I2859,I525192,I525181,);
nor I_30749 (I525619,I525554,I525311);
DFFARX1 I_30750 (I525619,I2859,I525192,I525160,);
nor I_30751 (I525650,I457568,I457571);
DFFARX1 I_30752 (I525650,I2859,I525192,I525676,);
DFFARX1 I_30753 (I525676,I2859,I525192,I525175,);
not I_30754 (I525698,I525676);
nand I_30755 (I525172,I525698,I525226);
nand I_30756 (I525166,I525698,I525328);
not I_30757 (I525770,I2866);
DFFARX1 I_30758 (I199358,I2859,I525770,I525796,);
nand I_30759 (I525804,I525796,I199367);
not I_30760 (I525821,I525804);
DFFARX1 I_30761 (I199355,I2859,I525770,I525847,);
not I_30762 (I525855,I525847);
not I_30763 (I525872,I199361);
or I_30764 (I525889,I199355,I199361);
nor I_30765 (I525906,I199355,I199361);
or I_30766 (I525923,I199370,I199355);
DFFARX1 I_30767 (I525923,I2859,I525770,I525762,);
not I_30768 (I525954,I199364);
nand I_30769 (I525971,I525954,I199379);
nand I_30770 (I525988,I525872,I525971);
and I_30771 (I525741,I525855,I525988);
nor I_30772 (I526019,I199364,I199382);
and I_30773 (I526036,I525855,I526019);
nor I_30774 (I525747,I525821,I526036);
DFFARX1 I_30775 (I526019,I2859,I525770,I526076,);
not I_30776 (I526084,I526076);
nor I_30777 (I525756,I525855,I526084);
or I_30778 (I526115,I525923,I199373);
nor I_30779 (I526132,I199373,I199370);
nand I_30780 (I526149,I525988,I526132);
nand I_30781 (I526166,I526115,I526149);
DFFARX1 I_30782 (I526166,I2859,I525770,I525759,);
nor I_30783 (I526197,I526132,I525889);
DFFARX1 I_30784 (I526197,I2859,I525770,I525738,);
nor I_30785 (I526228,I199373,I199376);
DFFARX1 I_30786 (I526228,I2859,I525770,I526254,);
DFFARX1 I_30787 (I526254,I2859,I525770,I525753,);
not I_30788 (I526276,I526254);
nand I_30789 (I525750,I526276,I525804);
nand I_30790 (I525744,I526276,I525906);
not I_30791 (I526348,I2866);
DFFARX1 I_30792 (I551449,I2859,I526348,I526374,);
nand I_30793 (I526382,I526374,I551440);
not I_30794 (I526399,I526382);
DFFARX1 I_30795 (I551425,I2859,I526348,I526425,);
not I_30796 (I526433,I526425);
not I_30797 (I526450,I551428);
or I_30798 (I526467,I551437,I551428);
nor I_30799 (I526484,I551437,I551428);
or I_30800 (I526501,I551434,I551437);
DFFARX1 I_30801 (I526501,I2859,I526348,I526340,);
not I_30802 (I526532,I551446);
nand I_30803 (I526549,I526532,I551425);
nand I_30804 (I526566,I526450,I526549);
and I_30805 (I526319,I526433,I526566);
nor I_30806 (I526597,I551446,I551431);
and I_30807 (I526614,I526433,I526597);
nor I_30808 (I526325,I526399,I526614);
DFFARX1 I_30809 (I526597,I2859,I526348,I526654,);
not I_30810 (I526662,I526654);
nor I_30811 (I526334,I526433,I526662);
or I_30812 (I526693,I526501,I551452);
nor I_30813 (I526710,I551452,I551434);
nand I_30814 (I526727,I526566,I526710);
nand I_30815 (I526744,I526693,I526727);
DFFARX1 I_30816 (I526744,I2859,I526348,I526337,);
nor I_30817 (I526775,I526710,I526467);
DFFARX1 I_30818 (I526775,I2859,I526348,I526316,);
nor I_30819 (I526806,I551452,I551443);
DFFARX1 I_30820 (I526806,I2859,I526348,I526832,);
DFFARX1 I_30821 (I526832,I2859,I526348,I526331,);
not I_30822 (I526854,I526832);
nand I_30823 (I526328,I526854,I526382);
nand I_30824 (I526322,I526854,I526484);
not I_30825 (I526926,I2866);
DFFARX1 I_30826 (I134540,I2859,I526926,I526952,);
nand I_30827 (I526960,I526952,I134561);
not I_30828 (I526977,I526960);
DFFARX1 I_30829 (I134555,I2859,I526926,I527003,);
not I_30830 (I527011,I527003);
not I_30831 (I527028,I134543);
or I_30832 (I527045,I134558,I134543);
nor I_30833 (I527062,I134558,I134543);
or I_30834 (I527079,I134549,I134558);
DFFARX1 I_30835 (I527079,I2859,I526926,I526918,);
not I_30836 (I527110,I134537);
nand I_30837 (I527127,I527110,I134534);
nand I_30838 (I527144,I527028,I527127);
and I_30839 (I526897,I527011,I527144);
nor I_30840 (I527175,I134537,I134546);
and I_30841 (I527192,I527011,I527175);
nor I_30842 (I526903,I526977,I527192);
DFFARX1 I_30843 (I527175,I2859,I526926,I527232,);
not I_30844 (I527240,I527232);
nor I_30845 (I526912,I527011,I527240);
or I_30846 (I527271,I527079,I134552);
nor I_30847 (I527288,I134552,I134549);
nand I_30848 (I527305,I527144,I527288);
nand I_30849 (I527322,I527271,I527305);
DFFARX1 I_30850 (I527322,I2859,I526926,I526915,);
nor I_30851 (I527353,I527288,I527045);
DFFARX1 I_30852 (I527353,I2859,I526926,I526894,);
nor I_30853 (I527384,I134552,I134534);
DFFARX1 I_30854 (I527384,I2859,I526926,I527410,);
DFFARX1 I_30855 (I527410,I2859,I526926,I526909,);
not I_30856 (I527432,I527410);
nand I_30857 (I526906,I527432,I526960);
nand I_30858 (I526900,I527432,I527062);
not I_30859 (I527504,I2866);
DFFARX1 I_30860 (I209694,I2859,I527504,I527530,);
nand I_30861 (I527538,I527530,I209703);
not I_30862 (I527555,I527538);
DFFARX1 I_30863 (I209691,I2859,I527504,I527581,);
not I_30864 (I527589,I527581);
not I_30865 (I527606,I209697);
or I_30866 (I527623,I209691,I209697);
nor I_30867 (I527640,I209691,I209697);
or I_30868 (I527657,I209706,I209691);
DFFARX1 I_30869 (I527657,I2859,I527504,I527496,);
not I_30870 (I527688,I209700);
nand I_30871 (I527705,I527688,I209715);
nand I_30872 (I527722,I527606,I527705);
and I_30873 (I527475,I527589,I527722);
nor I_30874 (I527753,I209700,I209718);
and I_30875 (I527770,I527589,I527753);
nor I_30876 (I527481,I527555,I527770);
DFFARX1 I_30877 (I527753,I2859,I527504,I527810,);
not I_30878 (I527818,I527810);
nor I_30879 (I527490,I527589,I527818);
or I_30880 (I527849,I527657,I209709);
nor I_30881 (I527866,I209709,I209706);
nand I_30882 (I527883,I527722,I527866);
nand I_30883 (I527900,I527849,I527883);
DFFARX1 I_30884 (I527900,I2859,I527504,I527493,);
nor I_30885 (I527931,I527866,I527623);
DFFARX1 I_30886 (I527931,I2859,I527504,I527472,);
nor I_30887 (I527962,I209709,I209712);
DFFARX1 I_30888 (I527962,I2859,I527504,I527988,);
DFFARX1 I_30889 (I527988,I2859,I527504,I527487,);
not I_30890 (I528010,I527988);
nand I_30891 (I527484,I528010,I527538);
nand I_30892 (I527478,I528010,I527640);
not I_30893 (I528082,I2866);
DFFARX1 I_30894 (I470880,I2859,I528082,I528108,);
nand I_30895 (I528116,I528108,I470865);
not I_30896 (I528133,I528116);
DFFARX1 I_30897 (I470868,I2859,I528082,I528159,);
not I_30898 (I528167,I528159);
not I_30899 (I528184,I470883);
or I_30900 (I528201,I470886,I470883);
nor I_30901 (I528218,I470886,I470883);
or I_30902 (I528235,I470862,I470886);
DFFARX1 I_30903 (I528235,I2859,I528082,I528074,);
not I_30904 (I528266,I470874);
nand I_30905 (I528283,I528266,I470877);
nand I_30906 (I528300,I528184,I528283);
and I_30907 (I528053,I528167,I528300);
nor I_30908 (I528331,I470874,I470871);
and I_30909 (I528348,I528167,I528331);
nor I_30910 (I528059,I528133,I528348);
DFFARX1 I_30911 (I528331,I2859,I528082,I528388,);
not I_30912 (I528396,I528388);
nor I_30913 (I528068,I528167,I528396);
or I_30914 (I528427,I528235,I470862);
nor I_30915 (I528444,I470862,I470862);
nand I_30916 (I528461,I528300,I528444);
nand I_30917 (I528478,I528427,I528461);
DFFARX1 I_30918 (I528478,I2859,I528082,I528071,);
nor I_30919 (I528509,I528444,I528201);
DFFARX1 I_30920 (I528509,I2859,I528082,I528050,);
nor I_30921 (I528540,I470862,I470865);
DFFARX1 I_30922 (I528540,I2859,I528082,I528566,);
DFFARX1 I_30923 (I528566,I2859,I528082,I528065,);
not I_30924 (I528588,I528566);
nand I_30925 (I528062,I528588,I528116);
nand I_30926 (I528056,I528588,I528218);
not I_30927 (I528660,I2866);
DFFARX1 I_30928 (I310110,I2859,I528660,I528686,);
nand I_30929 (I528694,I528686,I310113);
not I_30930 (I528711,I528694);
DFFARX1 I_30931 (I310125,I2859,I528660,I528737,);
not I_30932 (I528745,I528737);
not I_30933 (I528762,I310110);
or I_30934 (I528779,I310119,I310110);
nor I_30935 (I528796,I310119,I310110);
or I_30936 (I528813,I310128,I310119);
DFFARX1 I_30937 (I528813,I2859,I528660,I528652,);
not I_30938 (I528844,I310131);
nand I_30939 (I528861,I528844,I310113);
nand I_30940 (I528878,I528762,I528861);
and I_30941 (I528631,I528745,I528878);
nor I_30942 (I528909,I310131,I310116);
and I_30943 (I528926,I528745,I528909);
nor I_30944 (I528637,I528711,I528926);
DFFARX1 I_30945 (I528909,I2859,I528660,I528966,);
not I_30946 (I528974,I528966);
nor I_30947 (I528646,I528745,I528974);
or I_30948 (I529005,I528813,I310122);
nor I_30949 (I529022,I310122,I310128);
nand I_30950 (I529039,I528878,I529022);
nand I_30951 (I529056,I529005,I529039);
DFFARX1 I_30952 (I529056,I2859,I528660,I528649,);
nor I_30953 (I529087,I529022,I528779);
DFFARX1 I_30954 (I529087,I2859,I528660,I528628,);
nor I_30955 (I529118,I310122,I310134);
DFFARX1 I_30956 (I529118,I2859,I528660,I529144,);
DFFARX1 I_30957 (I529144,I2859,I528660,I528643,);
not I_30958 (I529166,I529144);
nand I_30959 (I528640,I529166,I528694);
nand I_30960 (I528634,I529166,I528796);
not I_30961 (I529238,I2866);
DFFARX1 I_30962 (I59018,I2859,I529238,I529264,);
nand I_30963 (I529272,I529264,I59027);
not I_30964 (I529289,I529272);
DFFARX1 I_30965 (I59009,I2859,I529238,I529315,);
not I_30966 (I529323,I529315);
not I_30967 (I529340,I59015);
or I_30968 (I529357,I59024,I59015);
nor I_30969 (I529374,I59024,I59015);
or I_30970 (I529391,I59012,I59024);
DFFARX1 I_30971 (I529391,I2859,I529238,I529230,);
not I_30972 (I529422,I59030);
nand I_30973 (I529439,I529422,I59003);
nand I_30974 (I529456,I529340,I529439);
and I_30975 (I529209,I529323,I529456);
nor I_30976 (I529487,I59030,I59006);
and I_30977 (I529504,I529323,I529487);
nor I_30978 (I529215,I529289,I529504);
DFFARX1 I_30979 (I529487,I2859,I529238,I529544,);
not I_30980 (I529552,I529544);
nor I_30981 (I529224,I529323,I529552);
or I_30982 (I529583,I529391,I59021);
nor I_30983 (I529600,I59021,I59012);
nand I_30984 (I529617,I529456,I529600);
nand I_30985 (I529634,I529583,I529617);
DFFARX1 I_30986 (I529634,I2859,I529238,I529227,);
nor I_30987 (I529665,I529600,I529357);
DFFARX1 I_30988 (I529665,I2859,I529238,I529206,);
nor I_30989 (I529696,I59021,I59003);
DFFARX1 I_30990 (I529696,I2859,I529238,I529722,);
DFFARX1 I_30991 (I529722,I2859,I529238,I529221,);
not I_30992 (I529744,I529722);
nand I_30993 (I529218,I529744,I529272);
nand I_30994 (I529212,I529744,I529374);
not I_30995 (I529816,I2866);
DFFARX1 I_30996 (I337925,I2859,I529816,I529842,);
nand I_30997 (I529850,I529842,I337925);
not I_30998 (I529867,I529850);
DFFARX1 I_30999 (I337931,I2859,I529816,I529893,);
not I_31000 (I529901,I529893);
not I_31001 (I529918,I337943);
or I_31002 (I529935,I337928,I337943);
nor I_31003 (I529952,I337928,I337943);
or I_31004 (I529969,I337922,I337928);
DFFARX1 I_31005 (I529969,I2859,I529816,I529808,);
not I_31006 (I530000,I337940);
nand I_31007 (I530017,I530000,I337934);
nand I_31008 (I530034,I529918,I530017);
and I_31009 (I529787,I529901,I530034);
nor I_31010 (I530065,I337940,I337922);
and I_31011 (I530082,I529901,I530065);
nor I_31012 (I529793,I529867,I530082);
DFFARX1 I_31013 (I530065,I2859,I529816,I530122,);
not I_31014 (I530130,I530122);
nor I_31015 (I529802,I529901,I530130);
or I_31016 (I530161,I529969,I337937);
nor I_31017 (I530178,I337937,I337922);
nand I_31018 (I530195,I530034,I530178);
nand I_31019 (I530212,I530161,I530195);
DFFARX1 I_31020 (I530212,I2859,I529816,I529805,);
nor I_31021 (I530243,I530178,I529935);
DFFARX1 I_31022 (I530243,I2859,I529816,I529784,);
nor I_31023 (I530274,I337937,I337928);
DFFARX1 I_31024 (I530274,I2859,I529816,I530300,);
DFFARX1 I_31025 (I530300,I2859,I529816,I529799,);
not I_31026 (I530322,I530300);
nand I_31027 (I529796,I530322,I529850);
nand I_31028 (I529790,I530322,I529952);
not I_31029 (I530394,I2866);
DFFARX1 I_31030 (I31543,I2859,I530394,I530420,);
nand I_31031 (I530428,I530420,I31534);
not I_31032 (I530445,I530428);
DFFARX1 I_31033 (I31531,I2859,I530394,I530471,);
not I_31034 (I530479,I530471);
not I_31035 (I530496,I31540);
or I_31036 (I530513,I31531,I31540);
nor I_31037 (I530530,I31531,I31540);
or I_31038 (I530547,I31537,I31531);
DFFARX1 I_31039 (I530547,I2859,I530394,I530386,);
not I_31040 (I530578,I31546);
nand I_31041 (I530595,I530578,I31555);
nand I_31042 (I530612,I530496,I530595);
and I_31043 (I530365,I530479,I530612);
nor I_31044 (I530643,I31546,I31549);
and I_31045 (I530660,I530479,I530643);
nor I_31046 (I530371,I530445,I530660);
DFFARX1 I_31047 (I530643,I2859,I530394,I530700,);
not I_31048 (I530708,I530700);
nor I_31049 (I530380,I530479,I530708);
or I_31050 (I530739,I530547,I31534);
nor I_31051 (I530756,I31534,I31537);
nand I_31052 (I530773,I530612,I530756);
nand I_31053 (I530790,I530739,I530773);
DFFARX1 I_31054 (I530790,I2859,I530394,I530383,);
nor I_31055 (I530821,I530756,I530513);
DFFARX1 I_31056 (I530821,I2859,I530394,I530362,);
nor I_31057 (I530852,I31534,I31552);
DFFARX1 I_31058 (I530852,I2859,I530394,I530878,);
DFFARX1 I_31059 (I530878,I2859,I530394,I530377,);
not I_31060 (I530900,I530878);
nand I_31061 (I530374,I530900,I530428);
nand I_31062 (I530368,I530900,I530530);
not I_31063 (I530972,I2866);
DFFARX1 I_31064 (I428133,I2859,I530972,I530998,);
nand I_31065 (I531006,I530998,I428130);
not I_31066 (I531023,I531006);
DFFARX1 I_31067 (I428130,I2859,I530972,I531049,);
not I_31068 (I531057,I531049);
not I_31069 (I531074,I428127);
or I_31070 (I531091,I428136,I428127);
nor I_31071 (I531108,I428136,I428127);
or I_31072 (I531125,I428139,I428136);
DFFARX1 I_31073 (I531125,I2859,I530972,I530964,);
not I_31074 (I531156,I428127);
nand I_31075 (I531173,I531156,I428124);
nand I_31076 (I531190,I531074,I531173);
and I_31077 (I530943,I531057,I531190);
nor I_31078 (I531221,I428127,I428142);
and I_31079 (I531238,I531057,I531221);
nor I_31080 (I530949,I531023,I531238);
DFFARX1 I_31081 (I531221,I2859,I530972,I531278,);
not I_31082 (I531286,I531278);
nor I_31083 (I530958,I531057,I531286);
or I_31084 (I531317,I531125,I428145);
nor I_31085 (I531334,I428145,I428139);
nand I_31086 (I531351,I531190,I531334);
nand I_31087 (I531368,I531317,I531351);
DFFARX1 I_31088 (I531368,I2859,I530972,I530961,);
nor I_31089 (I531399,I531334,I531091);
DFFARX1 I_31090 (I531399,I2859,I530972,I530940,);
nor I_31091 (I531430,I428145,I428124);
DFFARX1 I_31092 (I531430,I2859,I530972,I531456,);
DFFARX1 I_31093 (I531456,I2859,I530972,I530955,);
not I_31094 (I531478,I531456);
nand I_31095 (I530952,I531478,I531006);
nand I_31096 (I530946,I531478,I531108);
not I_31097 (I531550,I2866);
DFFARX1 I_31098 (I148242,I2859,I531550,I531576,);
nand I_31099 (I531584,I531576,I148263);
not I_31100 (I531601,I531584);
DFFARX1 I_31101 (I148257,I2859,I531550,I531627,);
not I_31102 (I531635,I531627);
not I_31103 (I531652,I148245);
or I_31104 (I531669,I148260,I148245);
nor I_31105 (I531686,I148260,I148245);
or I_31106 (I531703,I148251,I148260);
DFFARX1 I_31107 (I531703,I2859,I531550,I531542,);
not I_31108 (I531734,I148239);
nand I_31109 (I531751,I531734,I148236);
nand I_31110 (I531768,I531652,I531751);
and I_31111 (I531521,I531635,I531768);
nor I_31112 (I531799,I148239,I148248);
and I_31113 (I531816,I531635,I531799);
nor I_31114 (I531527,I531601,I531816);
DFFARX1 I_31115 (I531799,I2859,I531550,I531856,);
not I_31116 (I531864,I531856);
nor I_31117 (I531536,I531635,I531864);
or I_31118 (I531895,I531703,I148254);
nor I_31119 (I531912,I148254,I148251);
nand I_31120 (I531929,I531768,I531912);
nand I_31121 (I531946,I531895,I531929);
DFFARX1 I_31122 (I531946,I2859,I531550,I531539,);
nor I_31123 (I531977,I531912,I531669);
DFFARX1 I_31124 (I531977,I2859,I531550,I531518,);
nor I_31125 (I532008,I148254,I148236);
DFFARX1 I_31126 (I532008,I2859,I531550,I532034,);
DFFARX1 I_31127 (I532034,I2859,I531550,I531533,);
not I_31128 (I532056,I532034);
nand I_31129 (I531530,I532056,I531584);
nand I_31130 (I531524,I532056,I531686);
not I_31131 (I532128,I2866);
DFFARX1 I_31132 (I537826,I2859,I532128,I532154,);
nand I_31133 (I532162,I532154,I537820);
not I_31134 (I532179,I532162);
DFFARX1 I_31135 (I537835,I2859,I532128,I532205,);
not I_31136 (I532213,I532205);
not I_31137 (I532230,I537811);
or I_31138 (I532247,I537808,I537811);
nor I_31139 (I532264,I537808,I537811);
or I_31140 (I532281,I537814,I537808);
DFFARX1 I_31141 (I532281,I2859,I532128,I532120,);
not I_31142 (I532312,I537808);
nand I_31143 (I532329,I532312,I537823);
nand I_31144 (I532346,I532230,I532329);
and I_31145 (I532099,I532213,I532346);
nor I_31146 (I532377,I537808,I537817);
and I_31147 (I532394,I532213,I532377);
nor I_31148 (I532105,I532179,I532394);
DFFARX1 I_31149 (I532377,I2859,I532128,I532434,);
not I_31150 (I532442,I532434);
nor I_31151 (I532114,I532213,I532442);
or I_31152 (I532473,I532281,I537832);
nor I_31153 (I532490,I537832,I537814);
nand I_31154 (I532507,I532346,I532490);
nand I_31155 (I532524,I532473,I532507);
DFFARX1 I_31156 (I532524,I2859,I532128,I532117,);
nor I_31157 (I532555,I532490,I532247);
DFFARX1 I_31158 (I532555,I2859,I532128,I532096,);
nor I_31159 (I532586,I537832,I537829);
DFFARX1 I_31160 (I532586,I2859,I532128,I532612,);
DFFARX1 I_31161 (I532612,I2859,I532128,I532111,);
not I_31162 (I532634,I532612);
nand I_31163 (I532108,I532634,I532162);
nand I_31164 (I532102,I532634,I532264);
not I_31165 (I532706,I2866);
DFFARX1 I_31166 (I508617,I2859,I532706,I532732,);
nand I_31167 (I532740,I532732,I508626);
not I_31168 (I532757,I532740);
DFFARX1 I_31169 (I508602,I2859,I532706,I532783,);
not I_31170 (I532791,I532783);
not I_31171 (I532808,I508605);
or I_31172 (I532825,I508602,I508605);
nor I_31173 (I532842,I508602,I508605);
or I_31174 (I532859,I508620,I508602);
DFFARX1 I_31175 (I532859,I2859,I532706,I532698,);
not I_31176 (I532890,I508608);
nand I_31177 (I532907,I532890,I508623);
nand I_31178 (I532924,I532808,I532907);
and I_31179 (I532677,I532791,I532924);
nor I_31180 (I532955,I508608,I508611);
and I_31181 (I532972,I532791,I532955);
nor I_31182 (I532683,I532757,I532972);
DFFARX1 I_31183 (I532955,I2859,I532706,I533012,);
not I_31184 (I533020,I533012);
nor I_31185 (I532692,I532791,I533020);
or I_31186 (I533051,I532859,I508614);
nor I_31187 (I533068,I508614,I508620);
nand I_31188 (I533085,I532924,I533068);
nand I_31189 (I533102,I533051,I533085);
DFFARX1 I_31190 (I533102,I2859,I532706,I532695,);
nor I_31191 (I533133,I533068,I532825);
DFFARX1 I_31192 (I533133,I2859,I532706,I532674,);
nor I_31193 (I533164,I508614,I508605);
DFFARX1 I_31194 (I533164,I2859,I532706,I533190,);
DFFARX1 I_31195 (I533190,I2859,I532706,I532689,);
not I_31196 (I533212,I533190);
nand I_31197 (I532686,I533212,I532740);
nand I_31198 (I532680,I533212,I532842);
not I_31199 (I533284,I2866);
DFFARX1 I_31200 (I343195,I2859,I533284,I533310,);
nand I_31201 (I533318,I533310,I343195);
not I_31202 (I533335,I533318);
DFFARX1 I_31203 (I343201,I2859,I533284,I533361,);
not I_31204 (I533369,I533361);
not I_31205 (I533386,I343213);
or I_31206 (I533403,I343198,I343213);
nor I_31207 (I533420,I343198,I343213);
or I_31208 (I533437,I343192,I343198);
DFFARX1 I_31209 (I533437,I2859,I533284,I533276,);
not I_31210 (I533468,I343210);
nand I_31211 (I533485,I533468,I343204);
nand I_31212 (I533502,I533386,I533485);
and I_31213 (I533255,I533369,I533502);
nor I_31214 (I533533,I343210,I343192);
and I_31215 (I533550,I533369,I533533);
nor I_31216 (I533261,I533335,I533550);
DFFARX1 I_31217 (I533533,I2859,I533284,I533590,);
not I_31218 (I533598,I533590);
nor I_31219 (I533270,I533369,I533598);
or I_31220 (I533629,I533437,I343207);
nor I_31221 (I533646,I343207,I343192);
nand I_31222 (I533663,I533502,I533646);
nand I_31223 (I533680,I533629,I533663);
DFFARX1 I_31224 (I533680,I2859,I533284,I533273,);
nor I_31225 (I533711,I533646,I533403);
DFFARX1 I_31226 (I533711,I2859,I533284,I533252,);
nor I_31227 (I533742,I343207,I343198);
DFFARX1 I_31228 (I533742,I2859,I533284,I533768,);
DFFARX1 I_31229 (I533768,I2859,I533284,I533267,);
not I_31230 (I533790,I533768);
nand I_31231 (I533264,I533790,I533318);
nand I_31232 (I533258,I533790,I533420);
not I_31233 (I533862,I2866);
DFFARX1 I_31234 (I326872,I2859,I533862,I533888,);
nand I_31235 (I533896,I533888,I326875);
not I_31236 (I533913,I533896);
DFFARX1 I_31237 (I326887,I2859,I533862,I533939,);
not I_31238 (I533947,I533939);
not I_31239 (I533964,I326872);
or I_31240 (I533981,I326881,I326872);
nor I_31241 (I533998,I326881,I326872);
or I_31242 (I534015,I326890,I326881);
DFFARX1 I_31243 (I534015,I2859,I533862,I533854,);
not I_31244 (I534046,I326893);
nand I_31245 (I534063,I534046,I326875);
nand I_31246 (I534080,I533964,I534063);
and I_31247 (I533833,I533947,I534080);
nor I_31248 (I534111,I326893,I326878);
and I_31249 (I534128,I533947,I534111);
nor I_31250 (I533839,I533913,I534128);
DFFARX1 I_31251 (I534111,I2859,I533862,I534168,);
not I_31252 (I534176,I534168);
nor I_31253 (I533848,I533947,I534176);
or I_31254 (I534207,I534015,I326884);
nor I_31255 (I534224,I326884,I326890);
nand I_31256 (I534241,I534080,I534224);
nand I_31257 (I534258,I534207,I534241);
DFFARX1 I_31258 (I534258,I2859,I533862,I533851,);
nor I_31259 (I534289,I534224,I533981);
DFFARX1 I_31260 (I534289,I2859,I533862,I533830,);
nor I_31261 (I534320,I326884,I326896);
DFFARX1 I_31262 (I534320,I2859,I533862,I534346,);
DFFARX1 I_31263 (I534346,I2859,I533862,I533845,);
not I_31264 (I534368,I534346);
nand I_31265 (I533842,I534368,I533896);
nand I_31266 (I533836,I534368,I533998);
not I_31267 (I534440,I2866);
DFFARX1 I_31268 (I476660,I2859,I534440,I534466,);
nand I_31269 (I534474,I534466,I476645);
not I_31270 (I534491,I534474);
DFFARX1 I_31271 (I476648,I2859,I534440,I534517,);
not I_31272 (I534525,I534517);
not I_31273 (I534542,I476663);
or I_31274 (I534559,I476666,I476663);
nor I_31275 (I534576,I476666,I476663);
or I_31276 (I534593,I476642,I476666);
DFFARX1 I_31277 (I534593,I2859,I534440,I534432,);
not I_31278 (I534624,I476654);
nand I_31279 (I534641,I534624,I476657);
nand I_31280 (I534658,I534542,I534641);
and I_31281 (I534411,I534525,I534658);
nor I_31282 (I534689,I476654,I476651);
and I_31283 (I534706,I534525,I534689);
nor I_31284 (I534417,I534491,I534706);
DFFARX1 I_31285 (I534689,I2859,I534440,I534746,);
not I_31286 (I534754,I534746);
nor I_31287 (I534426,I534525,I534754);
or I_31288 (I534785,I534593,I476642);
nor I_31289 (I534802,I476642,I476642);
nand I_31290 (I534819,I534658,I534802);
nand I_31291 (I534836,I534785,I534819);
DFFARX1 I_31292 (I534836,I2859,I534440,I534429,);
nor I_31293 (I534867,I534802,I534559);
DFFARX1 I_31294 (I534867,I2859,I534440,I534408,);
nor I_31295 (I534898,I476642,I476645);
DFFARX1 I_31296 (I534898,I2859,I534440,I534924,);
DFFARX1 I_31297 (I534924,I2859,I534440,I534423,);
not I_31298 (I534946,I534924);
nand I_31299 (I534420,I534946,I534474);
nand I_31300 (I534414,I534946,I534576);
not I_31301 (I535018,I2866);
DFFARX1 I_31302 (I41029,I2859,I535018,I535044,);
nand I_31303 (I535052,I535044,I41020);
not I_31304 (I535069,I535052);
DFFARX1 I_31305 (I41017,I2859,I535018,I535095,);
not I_31306 (I535103,I535095);
not I_31307 (I535120,I41026);
or I_31308 (I535137,I41017,I41026);
nor I_31309 (I535154,I41017,I41026);
or I_31310 (I535171,I41023,I41017);
DFFARX1 I_31311 (I535171,I2859,I535018,I535010,);
not I_31312 (I535202,I41032);
nand I_31313 (I535219,I535202,I41041);
nand I_31314 (I535236,I535120,I535219);
and I_31315 (I534989,I535103,I535236);
nor I_31316 (I535267,I41032,I41035);
and I_31317 (I535284,I535103,I535267);
nor I_31318 (I534995,I535069,I535284);
DFFARX1 I_31319 (I535267,I2859,I535018,I535324,);
not I_31320 (I535332,I535324);
nor I_31321 (I535004,I535103,I535332);
or I_31322 (I535363,I535171,I41020);
nor I_31323 (I535380,I41020,I41023);
nand I_31324 (I535397,I535236,I535380);
nand I_31325 (I535414,I535363,I535397);
DFFARX1 I_31326 (I535414,I2859,I535018,I535007,);
nor I_31327 (I535445,I535380,I535137);
DFFARX1 I_31328 (I535445,I2859,I535018,I534986,);
nor I_31329 (I535476,I41020,I41038);
DFFARX1 I_31330 (I535476,I2859,I535018,I535502,);
DFFARX1 I_31331 (I535502,I2859,I535018,I535001,);
not I_31332 (I535524,I535502);
nand I_31333 (I534998,I535524,I535052);
nand I_31334 (I534992,I535524,I535154);
not I_31335 (I535599,I2866);
DFFARX1 I_31336 (I327468,I2859,I535599,I535625,);
nand I_31337 (I535633,I535625,I327453);
not I_31338 (I535650,I535633);
DFFARX1 I_31339 (I327471,I2859,I535599,I535676,);
not I_31340 (I535684,I535676);
nor I_31341 (I535701,I327450,I327465);
not I_31342 (I535718,I535701);
DFFARX1 I_31343 (I535718,I2859,I535599,I535585,);
or I_31344 (I535749,I327462,I327450);
DFFARX1 I_31345 (I535749,I2859,I535599,I535588,);
not I_31346 (I535780,I327450);
nor I_31347 (I535797,I535780,I327459);
nor I_31348 (I535814,I535797,I327465);
nor I_31349 (I535831,I327459,I327453);
nor I_31350 (I535848,I535684,I535831);
nor I_31351 (I535573,I535650,I535848);
not I_31352 (I535879,I535831);
nand I_31353 (I535576,I535879,I535633);
nand I_31354 (I535570,I535879,I535701);
nor I_31355 (I535567,I535831,I535814);
nor I_31356 (I535938,I327456,I327462);
not I_31357 (I535955,I535938);
DFFARX1 I_31358 (I535938,I2859,I535599,I535981,);
not I_31359 (I535591,I535981);
nor I_31360 (I536003,I327456,I327474);
DFFARX1 I_31361 (I536003,I2859,I535599,I536029,);
and I_31362 (I536037,I536029,I327450);
nor I_31363 (I536054,I536037,I535955);
DFFARX1 I_31364 (I536054,I2859,I535599,I535582,);
nor I_31365 (I536085,I536029,I535814);
DFFARX1 I_31366 (I536085,I2859,I535599,I535564,);
nor I_31367 (I535579,I536029,I535718);
not I_31368 (I536160,I2866);
DFFARX1 I_31369 (I154054,I2859,I536160,I536186,);
nand I_31370 (I536194,I536186,I154033);
not I_31371 (I536211,I536194);
DFFARX1 I_31372 (I154042,I2859,I536160,I536237,);
not I_31373 (I536245,I536237);
nor I_31374 (I536262,I154036,I154048);
not I_31375 (I536279,I536262);
DFFARX1 I_31376 (I536279,I2859,I536160,I536146,);
or I_31377 (I536310,I154039,I154036);
DFFARX1 I_31378 (I536310,I2859,I536160,I536149,);
not I_31379 (I536341,I154060);
nor I_31380 (I536358,I536341,I154045);
nor I_31381 (I536375,I536358,I154048);
nor I_31382 (I536392,I154045,I154033);
nor I_31383 (I536409,I536245,I536392);
nor I_31384 (I536134,I536211,I536409);
not I_31385 (I536440,I536392);
nand I_31386 (I536137,I536440,I536194);
nand I_31387 (I536131,I536440,I536262);
nor I_31388 (I536128,I536392,I536375);
nor I_31389 (I536499,I154051,I154039);
not I_31390 (I536516,I536499);
DFFARX1 I_31391 (I536499,I2859,I536160,I536542,);
not I_31392 (I536152,I536542);
nor I_31393 (I536564,I154051,I154057);
DFFARX1 I_31394 (I536564,I2859,I536160,I536590,);
and I_31395 (I536598,I536590,I154036);
nor I_31396 (I536615,I536598,I536516);
DFFARX1 I_31397 (I536615,I2859,I536160,I536143,);
nor I_31398 (I536646,I536590,I536375);
DFFARX1 I_31399 (I536646,I2859,I536160,I536125,);
nor I_31400 (I536140,I536590,I536279);
not I_31401 (I536721,I2866);
DFFARX1 I_31402 (I426453,I2859,I536721,I536747,);
nand I_31403 (I536755,I536747,I426456);
not I_31404 (I536772,I536755);
DFFARX1 I_31405 (I426444,I2859,I536721,I536798,);
not I_31406 (I536806,I536798);
nor I_31407 (I536823,I426462,I426459);
not I_31408 (I536840,I536823);
DFFARX1 I_31409 (I536840,I2859,I536721,I536707,);
or I_31410 (I536871,I426441,I426462);
DFFARX1 I_31411 (I536871,I2859,I536721,I536710,);
not I_31412 (I536902,I426441);
nor I_31413 (I536919,I536902,I426444);
nor I_31414 (I536936,I536919,I426459);
nor I_31415 (I536953,I426444,I426447);
nor I_31416 (I536970,I536806,I536953);
nor I_31417 (I536695,I536772,I536970);
not I_31418 (I537001,I536953);
nand I_31419 (I536698,I537001,I536755);
nand I_31420 (I536692,I537001,I536823);
nor I_31421 (I536689,I536953,I536936);
nor I_31422 (I537060,I426450,I426441);
not I_31423 (I537077,I537060);
DFFARX1 I_31424 (I537060,I2859,I536721,I537103,);
not I_31425 (I536713,I537103);
nor I_31426 (I537125,I426450,I426447);
DFFARX1 I_31427 (I537125,I2859,I536721,I537151,);
and I_31428 (I537159,I537151,I426462);
nor I_31429 (I537176,I537159,I537077);
DFFARX1 I_31430 (I537176,I2859,I536721,I536704,);
nor I_31431 (I537207,I537151,I536936);
DFFARX1 I_31432 (I537207,I2859,I536721,I536686,);
nor I_31433 (I536701,I537151,I536840);
not I_31434 (I537282,I2866);
DFFARX1 I_31435 (I2875,I2859,I537282,I537308,);
nand I_31436 (I537316,I537308,I2872);
not I_31437 (I537333,I537316);
DFFARX1 I_31438 (I2872,I2859,I537282,I537359,);
not I_31439 (I537367,I537359);
nor I_31440 (I537384,I2890,I2884);
not I_31441 (I537401,I537384);
DFFARX1 I_31442 (I537401,I2859,I537282,I537268,);
or I_31443 (I537432,I2887,I2890);
DFFARX1 I_31444 (I537432,I2859,I537282,I537271,);
not I_31445 (I537463,I2875);
nor I_31446 (I537480,I537463,I2869);
nor I_31447 (I537497,I537480,I2884);
nor I_31448 (I537514,I2869,I2881);
nor I_31449 (I537531,I537367,I537514);
nor I_31450 (I537256,I537333,I537531);
not I_31451 (I537562,I537514);
nand I_31452 (I537259,I537562,I537316);
nand I_31453 (I537253,I537562,I537384);
nor I_31454 (I537250,I537514,I537497);
nor I_31455 (I537621,I2878,I2887);
not I_31456 (I537638,I537621);
DFFARX1 I_31457 (I537621,I2859,I537282,I537664,);
not I_31458 (I537274,I537664);
nor I_31459 (I537686,I2878,I2869);
DFFARX1 I_31460 (I537686,I2859,I537282,I537712,);
and I_31461 (I537720,I537712,I2890);
nor I_31462 (I537737,I537720,I537638);
DFFARX1 I_31463 (I537737,I2859,I537282,I537265,);
nor I_31464 (I537768,I537712,I537497);
DFFARX1 I_31465 (I537768,I2859,I537282,I537247,);
nor I_31466 (I537262,I537712,I537401);
not I_31467 (I537843,I2866);
DFFARX1 I_31468 (I352681,I2859,I537843,I537869,);
nand I_31469 (I537877,I537869,I352699);
not I_31470 (I537894,I537877);
DFFARX1 I_31471 (I352678,I2859,I537843,I537920,);
not I_31472 (I537928,I537920);
nor I_31473 (I537945,I352693,I352687);
not I_31474 (I537962,I537945);
DFFARX1 I_31475 (I537962,I2859,I537843,I537829,);
or I_31476 (I537993,I352684,I352693);
DFFARX1 I_31477 (I537993,I2859,I537843,I537832,);
not I_31478 (I538024,I352684);
nor I_31479 (I538041,I538024,I352690);
nor I_31480 (I538058,I538041,I352687);
nor I_31481 (I538075,I352690,I352678);
nor I_31482 (I538092,I537928,I538075);
nor I_31483 (I537817,I537894,I538092);
not I_31484 (I538123,I538075);
nand I_31485 (I537820,I538123,I537877);
nand I_31486 (I537814,I538123,I537945);
nor I_31487 (I537811,I538075,I538058);
nor I_31488 (I538182,I352681,I352684);
not I_31489 (I538199,I538182);
DFFARX1 I_31490 (I538182,I2859,I537843,I538225,);
not I_31491 (I537835,I538225);
nor I_31492 (I538247,I352681,I352696);
DFFARX1 I_31493 (I538247,I2859,I537843,I538273,);
and I_31494 (I538281,I538273,I352693);
nor I_31495 (I538298,I538281,I538199);
DFFARX1 I_31496 (I538298,I2859,I537843,I537826,);
nor I_31497 (I538329,I538273,I538058);
DFFARX1 I_31498 (I538329,I2859,I537843,I537808,);
nor I_31499 (I537823,I538273,I537962);
not I_31500 (I538404,I2866);
DFFARX1 I_31501 (I472021,I2859,I538404,I538430,);
nand I_31502 (I538438,I538430,I472018);
not I_31503 (I538455,I538438);
DFFARX1 I_31504 (I472021,I2859,I538404,I538481,);
not I_31505 (I538489,I538481);
nor I_31506 (I538506,I472039,I472033);
not I_31507 (I538523,I538506);
DFFARX1 I_31508 (I538523,I2859,I538404,I538390,);
or I_31509 (I538554,I472042,I472039);
DFFARX1 I_31510 (I538554,I2859,I538404,I538393,);
not I_31511 (I538585,I472030);
nor I_31512 (I538602,I538585,I472027);
nor I_31513 (I538619,I538602,I472033);
nor I_31514 (I538636,I472027,I472018);
nor I_31515 (I538653,I538489,I538636);
nor I_31516 (I538378,I538455,I538653);
not I_31517 (I538684,I538636);
nand I_31518 (I538381,I538684,I538438);
nand I_31519 (I538375,I538684,I538506);
nor I_31520 (I538372,I538636,I538619);
nor I_31521 (I538743,I472024,I472042);
not I_31522 (I538760,I538743);
DFFARX1 I_31523 (I538743,I2859,I538404,I538786,);
not I_31524 (I538396,I538786);
nor I_31525 (I538808,I472024,I472036);
DFFARX1 I_31526 (I538808,I2859,I538404,I538834,);
and I_31527 (I538842,I538834,I472039);
nor I_31528 (I538859,I538842,I538760);
DFFARX1 I_31529 (I538859,I2859,I538404,I538387,);
nor I_31530 (I538890,I538834,I538619);
DFFARX1 I_31531 (I538890,I2859,I538404,I538369,);
nor I_31532 (I538384,I538834,I538523);
not I_31533 (I538965,I2866);
DFFARX1 I_31534 (I336877,I2859,I538965,I538991,);
DFFARX1 I_31535 (I336874,I2859,I538965,I539008,);
not I_31536 (I539016,I539008);
nor I_31537 (I538933,I538991,I539016);
DFFARX1 I_31538 (I539016,I2859,I538965,I538948,);
nor I_31539 (I539061,I336889,I336871);
and I_31540 (I539078,I539061,I336868);
nor I_31541 (I539095,I539078,I336889);
not I_31542 (I539112,I336889);
and I_31543 (I539129,I539112,I336874);
nand I_31544 (I539146,I539129,I336886);
nor I_31545 (I539163,I539112,I539146);
DFFARX1 I_31546 (I539163,I2859,I538965,I538930,);
not I_31547 (I539194,I539146);
nand I_31548 (I539211,I539016,I539194);
nand I_31549 (I538942,I539078,I539194);
DFFARX1 I_31550 (I539112,I2859,I538965,I538957,);
not I_31551 (I539256,I336880);
nor I_31552 (I539273,I539256,I336874);
nor I_31553 (I539290,I539273,I539095);
DFFARX1 I_31554 (I539290,I2859,I538965,I538954,);
not I_31555 (I539321,I539273);
DFFARX1 I_31556 (I539321,I2859,I538965,I539347,);
not I_31557 (I539355,I539347);
nor I_31558 (I538951,I539355,I539273);
nor I_31559 (I539386,I539256,I336868);
and I_31560 (I539403,I539386,I336883);
or I_31561 (I539420,I539403,I336871);
DFFARX1 I_31562 (I539420,I2859,I538965,I539446,);
not I_31563 (I539454,I539446);
nand I_31564 (I539471,I539454,I539194);
not I_31565 (I538945,I539471);
nand I_31566 (I538939,I539471,I539211);
nand I_31567 (I538936,I539454,I539078);
not I_31568 (I539560,I2866);
DFFARX1 I_31569 (I196091,I2859,I539560,I539586,);
DFFARX1 I_31570 (I196097,I2859,I539560,I539603,);
not I_31571 (I539611,I539603);
nor I_31572 (I539528,I539586,I539611);
DFFARX1 I_31573 (I539611,I2859,I539560,I539543,);
nor I_31574 (I539656,I196106,I196091);
and I_31575 (I539673,I539656,I196118);
nor I_31576 (I539690,I539673,I196106);
not I_31577 (I539707,I196106);
and I_31578 (I539724,I539707,I196094);
nand I_31579 (I539741,I539724,I196115);
nor I_31580 (I539758,I539707,I539741);
DFFARX1 I_31581 (I539758,I2859,I539560,I539525,);
not I_31582 (I539789,I539741);
nand I_31583 (I539806,I539611,I539789);
nand I_31584 (I539537,I539673,I539789);
DFFARX1 I_31585 (I539707,I2859,I539560,I539552,);
not I_31586 (I539851,I196103);
nor I_31587 (I539868,I539851,I196094);
nor I_31588 (I539885,I539868,I539690);
DFFARX1 I_31589 (I539885,I2859,I539560,I539549,);
not I_31590 (I539916,I539868);
DFFARX1 I_31591 (I539916,I2859,I539560,I539942,);
not I_31592 (I539950,I539942);
nor I_31593 (I539546,I539950,I539868);
nor I_31594 (I539981,I539851,I196100);
and I_31595 (I539998,I539981,I196112);
or I_31596 (I540015,I539998,I196109);
DFFARX1 I_31597 (I540015,I2859,I539560,I540041,);
not I_31598 (I540049,I540041);
nand I_31599 (I540066,I540049,I539789);
not I_31600 (I539540,I540066);
nand I_31601 (I539534,I540066,I539806);
nand I_31602 (I539531,I540049,I539673);
not I_31603 (I540155,I2866);
DFFARX1 I_31604 (I123488,I2859,I540155,I540181,);
DFFARX1 I_31605 (I123482,I2859,I540155,I540198,);
not I_31606 (I540206,I540198);
nor I_31607 (I540123,I540181,I540206);
DFFARX1 I_31608 (I540206,I2859,I540155,I540138,);
nor I_31609 (I540251,I123470,I123491);
and I_31610 (I540268,I540251,I123485);
nor I_31611 (I540285,I540268,I123470);
not I_31612 (I540302,I123470);
and I_31613 (I540319,I540302,I123467);
nand I_31614 (I540336,I540319,I123479);
nor I_31615 (I540353,I540302,I540336);
DFFARX1 I_31616 (I540353,I2859,I540155,I540120,);
not I_31617 (I540384,I540336);
nand I_31618 (I540401,I540206,I540384);
nand I_31619 (I540132,I540268,I540384);
DFFARX1 I_31620 (I540302,I2859,I540155,I540147,);
not I_31621 (I540446,I123494);
nor I_31622 (I540463,I540446,I123467);
nor I_31623 (I540480,I540463,I540285);
DFFARX1 I_31624 (I540480,I2859,I540155,I540144,);
not I_31625 (I540511,I540463);
DFFARX1 I_31626 (I540511,I2859,I540155,I540537,);
not I_31627 (I540545,I540537);
nor I_31628 (I540141,I540545,I540463);
nor I_31629 (I540576,I540446,I123476);
and I_31630 (I540593,I540576,I123473);
or I_31631 (I540610,I540593,I123467);
DFFARX1 I_31632 (I540610,I2859,I540155,I540636,);
not I_31633 (I540644,I540636);
nand I_31634 (I540661,I540644,I540384);
not I_31635 (I540135,I540661);
nand I_31636 (I540129,I540661,I540401);
nand I_31637 (I540126,I540644,I540268);
not I_31638 (I540750,I2866);
DFFARX1 I_31639 (I368497,I2859,I540750,I540776,);
DFFARX1 I_31640 (I368494,I2859,I540750,I540793,);
not I_31641 (I540801,I540793);
nor I_31642 (I540718,I540776,I540801);
DFFARX1 I_31643 (I540801,I2859,I540750,I540733,);
nor I_31644 (I540846,I368509,I368491);
and I_31645 (I540863,I540846,I368488);
nor I_31646 (I540880,I540863,I368509);
not I_31647 (I540897,I368509);
and I_31648 (I540914,I540897,I368494);
nand I_31649 (I540931,I540914,I368506);
nor I_31650 (I540948,I540897,I540931);
DFFARX1 I_31651 (I540948,I2859,I540750,I540715,);
not I_31652 (I540979,I540931);
nand I_31653 (I540996,I540801,I540979);
nand I_31654 (I540727,I540863,I540979);
DFFARX1 I_31655 (I540897,I2859,I540750,I540742,);
not I_31656 (I541041,I368500);
nor I_31657 (I541058,I541041,I368494);
nor I_31658 (I541075,I541058,I540880);
DFFARX1 I_31659 (I541075,I2859,I540750,I540739,);
not I_31660 (I541106,I541058);
DFFARX1 I_31661 (I541106,I2859,I540750,I541132,);
not I_31662 (I541140,I541132);
nor I_31663 (I540736,I541140,I541058);
nor I_31664 (I541171,I541041,I368488);
and I_31665 (I541188,I541171,I368503);
or I_31666 (I541205,I541188,I368491);
DFFARX1 I_31667 (I541205,I2859,I540750,I541231,);
not I_31668 (I541239,I541231);
nand I_31669 (I541256,I541239,I540979);
not I_31670 (I540730,I541256);
nand I_31671 (I540724,I541256,I540996);
nand I_31672 (I540721,I541239,I540863);
not I_31673 (I541345,I2866);
DFFARX1 I_31674 (I385443,I2859,I541345,I541371,);
DFFARX1 I_31675 (I385461,I2859,I541345,I541388,);
not I_31676 (I541396,I541388);
nor I_31677 (I541313,I541371,I541396);
DFFARX1 I_31678 (I541396,I2859,I541345,I541328,);
nor I_31679 (I541441,I385440,I385452);
and I_31680 (I541458,I541441,I385437);
nor I_31681 (I541475,I541458,I385440);
not I_31682 (I541492,I385440);
and I_31683 (I541509,I541492,I385446);
nand I_31684 (I541526,I541509,I385458);
nor I_31685 (I541543,I541492,I541526);
DFFARX1 I_31686 (I541543,I2859,I541345,I541310,);
not I_31687 (I541574,I541526);
nand I_31688 (I541591,I541396,I541574);
nand I_31689 (I541322,I541458,I541574);
DFFARX1 I_31690 (I541492,I2859,I541345,I541337,);
not I_31691 (I541636,I385449);
nor I_31692 (I541653,I541636,I385446);
nor I_31693 (I541670,I541653,I541475);
DFFARX1 I_31694 (I541670,I2859,I541345,I541334,);
not I_31695 (I541701,I541653);
DFFARX1 I_31696 (I541701,I2859,I541345,I541727,);
not I_31697 (I541735,I541727);
nor I_31698 (I541331,I541735,I541653);
nor I_31699 (I541766,I541636,I385437);
and I_31700 (I541783,I541766,I385464);
or I_31701 (I541800,I541783,I385455);
DFFARX1 I_31702 (I541800,I2859,I541345,I541826,);
not I_31703 (I541834,I541826);
nand I_31704 (I541851,I541834,I541574);
not I_31705 (I541325,I541851);
nand I_31706 (I541319,I541851,I541591);
nand I_31707 (I541316,I541834,I541458);
not I_31708 (I541940,I2866);
DFFARX1 I_31709 (I267359,I2859,I541940,I541966,);
DFFARX1 I_31710 (I267341,I2859,I541940,I541983,);
not I_31711 (I541991,I541983);
nor I_31712 (I541908,I541966,I541991);
DFFARX1 I_31713 (I541991,I2859,I541940,I541923,);
nor I_31714 (I542036,I267347,I267350);
and I_31715 (I542053,I542036,I267338);
nor I_31716 (I542070,I542053,I267347);
not I_31717 (I542087,I267347);
and I_31718 (I542104,I542087,I267356);
nand I_31719 (I542121,I542104,I267344);
nor I_31720 (I542138,I542087,I542121);
DFFARX1 I_31721 (I542138,I2859,I541940,I541905,);
not I_31722 (I542169,I542121);
nand I_31723 (I542186,I541991,I542169);
nand I_31724 (I541917,I542053,I542169);
DFFARX1 I_31725 (I542087,I2859,I541940,I541932,);
not I_31726 (I542231,I267341);
nor I_31727 (I542248,I542231,I267356);
nor I_31728 (I542265,I542248,I542070);
DFFARX1 I_31729 (I542265,I2859,I541940,I541929,);
not I_31730 (I542296,I542248);
DFFARX1 I_31731 (I542296,I2859,I541940,I542322,);
not I_31732 (I542330,I542322);
nor I_31733 (I541926,I542330,I542248);
nor I_31734 (I542361,I542231,I267353);
and I_31735 (I542378,I542361,I267362);
or I_31736 (I542395,I542378,I267338);
DFFARX1 I_31737 (I542395,I2859,I541940,I542421,);
not I_31738 (I542429,I542421);
nand I_31739 (I542446,I542429,I542169);
not I_31740 (I541920,I542446);
nand I_31741 (I541914,I542446,I542186);
nand I_31742 (I541911,I542429,I542053);
not I_31743 (I542535,I2866);
DFFARX1 I_31744 (I334769,I2859,I542535,I542561,);
DFFARX1 I_31745 (I334766,I2859,I542535,I542578,);
not I_31746 (I542586,I542578);
nor I_31747 (I542503,I542561,I542586);
DFFARX1 I_31748 (I542586,I2859,I542535,I542518,);
nor I_31749 (I542631,I334781,I334763);
and I_31750 (I542648,I542631,I334760);
nor I_31751 (I542665,I542648,I334781);
not I_31752 (I542682,I334781);
and I_31753 (I542699,I542682,I334766);
nand I_31754 (I542716,I542699,I334778);
nor I_31755 (I542733,I542682,I542716);
DFFARX1 I_31756 (I542733,I2859,I542535,I542500,);
not I_31757 (I542764,I542716);
nand I_31758 (I542781,I542586,I542764);
nand I_31759 (I542512,I542648,I542764);
DFFARX1 I_31760 (I542682,I2859,I542535,I542527,);
not I_31761 (I542826,I334772);
nor I_31762 (I542843,I542826,I334766);
nor I_31763 (I542860,I542843,I542665);
DFFARX1 I_31764 (I542860,I2859,I542535,I542524,);
not I_31765 (I542891,I542843);
DFFARX1 I_31766 (I542891,I2859,I542535,I542917,);
not I_31767 (I542925,I542917);
nor I_31768 (I542521,I542925,I542843);
nor I_31769 (I542956,I542826,I334760);
and I_31770 (I542973,I542956,I334775);
or I_31771 (I542990,I542973,I334763);
DFFARX1 I_31772 (I542990,I2859,I542535,I543016,);
not I_31773 (I543024,I543016);
nand I_31774 (I543041,I543024,I542764);
not I_31775 (I542515,I543041);
nand I_31776 (I542509,I543041,I542781);
nand I_31777 (I542506,I543024,I542648);
not I_31778 (I543130,I2866);
DFFARX1 I_31779 (I321113,I2859,I543130,I543156,);
DFFARX1 I_31780 (I321095,I2859,I543130,I543173,);
not I_31781 (I543181,I543173);
nor I_31782 (I543098,I543156,I543181);
DFFARX1 I_31783 (I543181,I2859,I543130,I543113,);
nor I_31784 (I543226,I321101,I321104);
and I_31785 (I543243,I543226,I321092);
nor I_31786 (I543260,I543243,I321101);
not I_31787 (I543277,I321101);
and I_31788 (I543294,I543277,I321110);
nand I_31789 (I543311,I543294,I321098);
nor I_31790 (I543328,I543277,I543311);
DFFARX1 I_31791 (I543328,I2859,I543130,I543095,);
not I_31792 (I543359,I543311);
nand I_31793 (I543376,I543181,I543359);
nand I_31794 (I543107,I543243,I543359);
DFFARX1 I_31795 (I543277,I2859,I543130,I543122,);
not I_31796 (I543421,I321095);
nor I_31797 (I543438,I543421,I321110);
nor I_31798 (I543455,I543438,I543260);
DFFARX1 I_31799 (I543455,I2859,I543130,I543119,);
not I_31800 (I543486,I543438);
DFFARX1 I_31801 (I543486,I2859,I543130,I543512,);
not I_31802 (I543520,I543512);
nor I_31803 (I543116,I543520,I543438);
nor I_31804 (I543551,I543421,I321107);
and I_31805 (I543568,I543551,I321116);
or I_31806 (I543585,I543568,I321092);
DFFARX1 I_31807 (I543585,I2859,I543130,I543611,);
not I_31808 (I543619,I543611);
nand I_31809 (I543636,I543619,I543359);
not I_31810 (I543110,I543636);
nand I_31811 (I543104,I543636,I543376);
nand I_31812 (I543101,I543619,I543243);
not I_31813 (I543725,I2866);
DFFARX1 I_31814 (I288745,I2859,I543725,I543751,);
DFFARX1 I_31815 (I288727,I2859,I543725,I543768,);
not I_31816 (I543776,I543768);
nor I_31817 (I543693,I543751,I543776);
DFFARX1 I_31818 (I543776,I2859,I543725,I543708,);
nor I_31819 (I543821,I288733,I288736);
and I_31820 (I543838,I543821,I288724);
nor I_31821 (I543855,I543838,I288733);
not I_31822 (I543872,I288733);
and I_31823 (I543889,I543872,I288742);
nand I_31824 (I543906,I543889,I288730);
nor I_31825 (I543923,I543872,I543906);
DFFARX1 I_31826 (I543923,I2859,I543725,I543690,);
not I_31827 (I543954,I543906);
nand I_31828 (I543971,I543776,I543954);
nand I_31829 (I543702,I543838,I543954);
DFFARX1 I_31830 (I543872,I2859,I543725,I543717,);
not I_31831 (I544016,I288727);
nor I_31832 (I544033,I544016,I288742);
nor I_31833 (I544050,I544033,I543855);
DFFARX1 I_31834 (I544050,I2859,I543725,I543714,);
not I_31835 (I544081,I544033);
DFFARX1 I_31836 (I544081,I2859,I543725,I544107,);
not I_31837 (I544115,I544107);
nor I_31838 (I543711,I544115,I544033);
nor I_31839 (I544146,I544016,I288739);
and I_31840 (I544163,I544146,I288748);
or I_31841 (I544180,I544163,I288724);
DFFARX1 I_31842 (I544180,I2859,I543725,I544206,);
not I_31843 (I544214,I544206);
nand I_31844 (I544231,I544214,I543954);
not I_31845 (I543705,I544231);
nand I_31846 (I543699,I544231,I543971);
nand I_31847 (I543696,I544214,I543838);
not I_31848 (I544320,I2866);
DFFARX1 I_31849 (I47889,I2859,I544320,I544346,);
DFFARX1 I_31850 (I47877,I2859,I544320,I544363,);
not I_31851 (I544371,I544363);
nor I_31852 (I544288,I544346,I544371);
DFFARX1 I_31853 (I544371,I2859,I544320,I544303,);
nor I_31854 (I544416,I47868,I47892);
and I_31855 (I544433,I544416,I47871);
nor I_31856 (I544450,I544433,I47868);
not I_31857 (I544467,I47868);
and I_31858 (I544484,I544467,I47874);
nand I_31859 (I544501,I544484,I47886);
nor I_31860 (I544518,I544467,I544501);
DFFARX1 I_31861 (I544518,I2859,I544320,I544285,);
not I_31862 (I544549,I544501);
nand I_31863 (I544566,I544371,I544549);
nand I_31864 (I544297,I544433,I544549);
DFFARX1 I_31865 (I544467,I2859,I544320,I544312,);
not I_31866 (I544611,I47868);
nor I_31867 (I544628,I544611,I47874);
nor I_31868 (I544645,I544628,I544450);
DFFARX1 I_31869 (I544645,I2859,I544320,I544309,);
not I_31870 (I544676,I544628);
DFFARX1 I_31871 (I544676,I2859,I544320,I544702,);
not I_31872 (I544710,I544702);
nor I_31873 (I544306,I544710,I544628);
nor I_31874 (I544741,I544611,I47871);
and I_31875 (I544758,I544741,I47880);
or I_31876 (I544775,I544758,I47883);
DFFARX1 I_31877 (I544775,I2859,I544320,I544801,);
not I_31878 (I544809,I544801);
nand I_31879 (I544826,I544809,I544549);
not I_31880 (I544300,I544826);
nand I_31881 (I544294,I544826,I544566);
nand I_31882 (I544291,I544809,I544433);
not I_31883 (I544915,I2866);
DFFARX1 I_31884 (I33660,I2859,I544915,I544941,);
DFFARX1 I_31885 (I33648,I2859,I544915,I544958,);
not I_31886 (I544966,I544958);
nor I_31887 (I544883,I544941,I544966);
DFFARX1 I_31888 (I544966,I2859,I544915,I544898,);
nor I_31889 (I545011,I33639,I33663);
and I_31890 (I545028,I545011,I33642);
nor I_31891 (I545045,I545028,I33639);
not I_31892 (I545062,I33639);
and I_31893 (I545079,I545062,I33645);
nand I_31894 (I545096,I545079,I33657);
nor I_31895 (I545113,I545062,I545096);
DFFARX1 I_31896 (I545113,I2859,I544915,I544880,);
not I_31897 (I545144,I545096);
nand I_31898 (I545161,I544966,I545144);
nand I_31899 (I544892,I545028,I545144);
DFFARX1 I_31900 (I545062,I2859,I544915,I544907,);
not I_31901 (I545206,I33639);
nor I_31902 (I545223,I545206,I33645);
nor I_31903 (I545240,I545223,I545045);
DFFARX1 I_31904 (I545240,I2859,I544915,I544904,);
not I_31905 (I545271,I545223);
DFFARX1 I_31906 (I545271,I2859,I544915,I545297,);
not I_31907 (I545305,I545297);
nor I_31908 (I544901,I545305,I545223);
nor I_31909 (I545336,I545206,I33642);
and I_31910 (I545353,I545336,I33651);
or I_31911 (I545370,I545353,I33654);
DFFARX1 I_31912 (I545370,I2859,I544915,I545396,);
not I_31913 (I545404,I545396);
nand I_31914 (I545421,I545404,I545144);
not I_31915 (I544895,I545421);
nand I_31916 (I544889,I545421,I545161);
nand I_31917 (I544886,I545404,I545028);
not I_31918 (I545510,I2866);
DFFARX1 I_31919 (I210235,I2859,I545510,I545536,);
DFFARX1 I_31920 (I210241,I2859,I545510,I545553,);
not I_31921 (I545561,I545553);
nor I_31922 (I545478,I545536,I545561);
DFFARX1 I_31923 (I545561,I2859,I545510,I545493,);
nor I_31924 (I545606,I210250,I210235);
and I_31925 (I545623,I545606,I210262);
nor I_31926 (I545640,I545623,I210250);
not I_31927 (I545657,I210250);
and I_31928 (I545674,I545657,I210238);
nand I_31929 (I545691,I545674,I210259);
nor I_31930 (I545708,I545657,I545691);
DFFARX1 I_31931 (I545708,I2859,I545510,I545475,);
not I_31932 (I545739,I545691);
nand I_31933 (I545756,I545561,I545739);
nand I_31934 (I545487,I545623,I545739);
DFFARX1 I_31935 (I545657,I2859,I545510,I545502,);
not I_31936 (I545801,I210247);
nor I_31937 (I545818,I545801,I210238);
nor I_31938 (I545835,I545818,I545640);
DFFARX1 I_31939 (I545835,I2859,I545510,I545499,);
not I_31940 (I545866,I545818);
DFFARX1 I_31941 (I545866,I2859,I545510,I545892,);
not I_31942 (I545900,I545892);
nor I_31943 (I545496,I545900,I545818);
nor I_31944 (I545931,I545801,I210244);
and I_31945 (I545948,I545931,I210256);
or I_31946 (I545965,I545948,I210253);
DFFARX1 I_31947 (I545965,I2859,I545510,I545991,);
not I_31948 (I545999,I545991);
nand I_31949 (I546016,I545999,I545739);
not I_31950 (I545490,I546016);
nand I_31951 (I545484,I546016,I545756);
nand I_31952 (I545481,I545999,I545623);
not I_31953 (I546105,I2866);
DFFARX1 I_31954 (I413867,I2859,I546105,I546131,);
DFFARX1 I_31955 (I413885,I2859,I546105,I546148,);
not I_31956 (I546156,I546148);
nor I_31957 (I546073,I546131,I546156);
DFFARX1 I_31958 (I546156,I2859,I546105,I546088,);
nor I_31959 (I546201,I413864,I413876);
and I_31960 (I546218,I546201,I413861);
nor I_31961 (I546235,I546218,I413864);
not I_31962 (I546252,I413864);
and I_31963 (I546269,I546252,I413870);
nand I_31964 (I546286,I546269,I413882);
nor I_31965 (I546303,I546252,I546286);
DFFARX1 I_31966 (I546303,I2859,I546105,I546070,);
not I_31967 (I546334,I546286);
nand I_31968 (I546351,I546156,I546334);
nand I_31969 (I546082,I546218,I546334);
DFFARX1 I_31970 (I546252,I2859,I546105,I546097,);
not I_31971 (I546396,I413873);
nor I_31972 (I546413,I546396,I413870);
nor I_31973 (I546430,I546413,I546235);
DFFARX1 I_31974 (I546430,I2859,I546105,I546094,);
not I_31975 (I546461,I546413);
DFFARX1 I_31976 (I546461,I2859,I546105,I546487,);
not I_31977 (I546495,I546487);
nor I_31978 (I546091,I546495,I546413);
nor I_31979 (I546526,I546396,I413861);
and I_31980 (I546543,I546526,I413888);
or I_31981 (I546560,I546543,I413879);
DFFARX1 I_31982 (I546560,I2859,I546105,I546586,);
not I_31983 (I546594,I546586);
nand I_31984 (I546611,I546594,I546334);
not I_31985 (I546085,I546611);
nand I_31986 (I546079,I546611,I546351);
nand I_31987 (I546076,I546594,I546218);
not I_31988 (I546700,I2866);
DFFARX1 I_31989 (I244239,I2859,I546700,I546726,);
DFFARX1 I_31990 (I244233,I2859,I546700,I546743,);
not I_31991 (I546751,I546743);
nor I_31992 (I546668,I546726,I546751);
DFFARX1 I_31993 (I546751,I2859,I546700,I546683,);
nor I_31994 (I546796,I244230,I244221);
and I_31995 (I546813,I546796,I244218);
nor I_31996 (I546830,I546813,I244230);
not I_31997 (I546847,I244230);
and I_31998 (I546864,I546847,I244224);
nand I_31999 (I546881,I546864,I244236);
nor I_32000 (I546898,I546847,I546881);
DFFARX1 I_32001 (I546898,I2859,I546700,I546665,);
not I_32002 (I546929,I546881);
nand I_32003 (I546946,I546751,I546929);
nand I_32004 (I546677,I546813,I546929);
DFFARX1 I_32005 (I546847,I2859,I546700,I546692,);
not I_32006 (I546991,I244242);
nor I_32007 (I547008,I546991,I244224);
nor I_32008 (I547025,I547008,I546830);
DFFARX1 I_32009 (I547025,I2859,I546700,I546689,);
not I_32010 (I547056,I547008);
DFFARX1 I_32011 (I547056,I2859,I546700,I547082,);
not I_32012 (I547090,I547082);
nor I_32013 (I546686,I547090,I547008);
nor I_32014 (I547121,I546991,I244221);
and I_32015 (I547138,I547121,I244227);
or I_32016 (I547155,I547138,I244218);
DFFARX1 I_32017 (I547155,I2859,I546700,I547181,);
not I_32018 (I547189,I547181);
nand I_32019 (I547206,I547189,I546929);
not I_32020 (I546680,I547206);
nand I_32021 (I546674,I547206,I546946);
nand I_32022 (I546671,I547189,I546813);
not I_32023 (I547295,I2866);
DFFARX1 I_32024 (I237881,I2859,I547295,I547321,);
DFFARX1 I_32025 (I237875,I2859,I547295,I547338,);
not I_32026 (I547346,I547338);
nor I_32027 (I547263,I547321,I547346);
DFFARX1 I_32028 (I547346,I2859,I547295,I547278,);
nor I_32029 (I547391,I237872,I237863);
and I_32030 (I547408,I547391,I237860);
nor I_32031 (I547425,I547408,I237872);
not I_32032 (I547442,I237872);
and I_32033 (I547459,I547442,I237866);
nand I_32034 (I547476,I547459,I237878);
nor I_32035 (I547493,I547442,I547476);
DFFARX1 I_32036 (I547493,I2859,I547295,I547260,);
not I_32037 (I547524,I547476);
nand I_32038 (I547541,I547346,I547524);
nand I_32039 (I547272,I547408,I547524);
DFFARX1 I_32040 (I547442,I2859,I547295,I547287,);
not I_32041 (I547586,I237884);
nor I_32042 (I547603,I547586,I237866);
nor I_32043 (I547620,I547603,I547425);
DFFARX1 I_32044 (I547620,I2859,I547295,I547284,);
not I_32045 (I547651,I547603);
DFFARX1 I_32046 (I547651,I2859,I547295,I547677,);
not I_32047 (I547685,I547677);
nor I_32048 (I547281,I547685,I547603);
nor I_32049 (I547716,I547586,I237863);
and I_32050 (I547733,I547716,I237869);
or I_32051 (I547750,I547733,I237860);
DFFARX1 I_32052 (I547750,I2859,I547295,I547776,);
not I_32053 (I547784,I547776);
nand I_32054 (I547801,I547784,I547524);
not I_32055 (I547275,I547801);
nand I_32056 (I547269,I547801,I547541);
nand I_32057 (I547266,I547784,I547408);
not I_32058 (I547890,I2866);
DFFARX1 I_32059 (I514586,I2859,I547890,I547916,);
DFFARX1 I_32060 (I514589,I2859,I547890,I547933,);
not I_32061 (I547941,I547933);
nor I_32062 (I547858,I547916,I547941);
DFFARX1 I_32063 (I547941,I2859,I547890,I547873,);
nor I_32064 (I547986,I514589,I514604);
and I_32065 (I548003,I547986,I514598);
nor I_32066 (I548020,I548003,I514589);
not I_32067 (I548037,I514589);
and I_32068 (I548054,I548037,I514607);
nand I_32069 (I548071,I548054,I514595);
nor I_32070 (I548088,I548037,I548071);
DFFARX1 I_32071 (I548088,I2859,I547890,I547855,);
not I_32072 (I548119,I548071);
nand I_32073 (I548136,I547941,I548119);
nand I_32074 (I547867,I548003,I548119);
DFFARX1 I_32075 (I548037,I2859,I547890,I547882,);
not I_32076 (I548181,I514601);
nor I_32077 (I548198,I548181,I514607);
nor I_32078 (I548215,I548198,I548020);
DFFARX1 I_32079 (I548215,I2859,I547890,I547879,);
not I_32080 (I548246,I548198);
DFFARX1 I_32081 (I548246,I2859,I547890,I548272,);
not I_32082 (I548280,I548272);
nor I_32083 (I547876,I548280,I548198);
nor I_32084 (I548311,I548181,I514586);
and I_32085 (I548328,I548311,I514610);
or I_32086 (I548345,I548328,I514592);
DFFARX1 I_32087 (I548345,I2859,I547890,I548371,);
not I_32088 (I548379,I548371);
nand I_32089 (I548396,I548379,I548119);
not I_32090 (I547870,I548396);
nand I_32091 (I547864,I548396,I548136);
nand I_32092 (I547861,I548379,I548003);
not I_32093 (I548485,I2866);
DFFARX1 I_32094 (I32606,I2859,I548485,I548511,);
DFFARX1 I_32095 (I32594,I2859,I548485,I548528,);
not I_32096 (I548536,I548528);
nor I_32097 (I548453,I548511,I548536);
DFFARX1 I_32098 (I548536,I2859,I548485,I548468,);
nor I_32099 (I548581,I32585,I32609);
and I_32100 (I548598,I548581,I32588);
nor I_32101 (I548615,I548598,I32585);
not I_32102 (I548632,I32585);
and I_32103 (I548649,I548632,I32591);
nand I_32104 (I548666,I548649,I32603);
nor I_32105 (I548683,I548632,I548666);
DFFARX1 I_32106 (I548683,I2859,I548485,I548450,);
not I_32107 (I548714,I548666);
nand I_32108 (I548731,I548536,I548714);
nand I_32109 (I548462,I548598,I548714);
DFFARX1 I_32110 (I548632,I2859,I548485,I548477,);
not I_32111 (I548776,I32585);
nor I_32112 (I548793,I548776,I32591);
nor I_32113 (I548810,I548793,I548615);
DFFARX1 I_32114 (I548810,I2859,I548485,I548474,);
not I_32115 (I548841,I548793);
DFFARX1 I_32116 (I548841,I2859,I548485,I548867,);
not I_32117 (I548875,I548867);
nor I_32118 (I548471,I548875,I548793);
nor I_32119 (I548906,I548776,I32588);
and I_32120 (I548923,I548906,I32597);
or I_32121 (I548940,I548923,I32600);
DFFARX1 I_32122 (I548940,I2859,I548485,I548966,);
not I_32123 (I548974,I548966);
nand I_32124 (I548991,I548974,I548714);
not I_32125 (I548465,I548991);
nand I_32126 (I548459,I548991,I548731);
nand I_32127 (I548456,I548974,I548598);
not I_32128 (I549080,I2866);
DFFARX1 I_32129 (I406761,I2859,I549080,I549106,);
DFFARX1 I_32130 (I406779,I2859,I549080,I549123,);
not I_32131 (I549131,I549123);
nor I_32132 (I549048,I549106,I549131);
DFFARX1 I_32133 (I549131,I2859,I549080,I549063,);
nor I_32134 (I549176,I406758,I406770);
and I_32135 (I549193,I549176,I406755);
nor I_32136 (I549210,I549193,I406758);
not I_32137 (I549227,I406758);
and I_32138 (I549244,I549227,I406764);
nand I_32139 (I549261,I549244,I406776);
nor I_32140 (I549278,I549227,I549261);
DFFARX1 I_32141 (I549278,I2859,I549080,I549045,);
not I_32142 (I549309,I549261);
nand I_32143 (I549326,I549131,I549309);
nand I_32144 (I549057,I549193,I549309);
DFFARX1 I_32145 (I549227,I2859,I549080,I549072,);
not I_32146 (I549371,I406767);
nor I_32147 (I549388,I549371,I406764);
nor I_32148 (I549405,I549388,I549210);
DFFARX1 I_32149 (I549405,I2859,I549080,I549069,);
not I_32150 (I549436,I549388);
DFFARX1 I_32151 (I549436,I2859,I549080,I549462,);
not I_32152 (I549470,I549462);
nor I_32153 (I549066,I549470,I549388);
nor I_32154 (I549501,I549371,I406755);
and I_32155 (I549518,I549501,I406782);
or I_32156 (I549535,I549518,I406773);
DFFARX1 I_32157 (I549535,I2859,I549080,I549561,);
not I_32158 (I549569,I549561);
nand I_32159 (I549586,I549569,I549309);
not I_32160 (I549060,I549586);
nand I_32161 (I549054,I549586,I549326);
nand I_32162 (I549051,I549569,I549193);
not I_32163 (I549675,I2866);
DFFARX1 I_32164 (I17847,I2859,I549675,I549701,);
DFFARX1 I_32165 (I17829,I2859,I549675,I549718,);
not I_32166 (I549726,I549718);
nor I_32167 (I549643,I549701,I549726);
DFFARX1 I_32168 (I549726,I2859,I549675,I549658,);
nor I_32169 (I549771,I17829,I17844);
and I_32170 (I549788,I549771,I17838);
nor I_32171 (I549805,I549788,I17829);
not I_32172 (I549822,I17829);
and I_32173 (I549839,I549822,I17832);
nand I_32174 (I549856,I549839,I17835);
nor I_32175 (I549873,I549822,I549856);
DFFARX1 I_32176 (I549873,I2859,I549675,I549640,);
not I_32177 (I549904,I549856);
nand I_32178 (I549921,I549726,I549904);
nand I_32179 (I549652,I549788,I549904);
DFFARX1 I_32180 (I549822,I2859,I549675,I549667,);
not I_32181 (I549966,I17841);
nor I_32182 (I549983,I549966,I17832);
nor I_32183 (I550000,I549983,I549805);
DFFARX1 I_32184 (I550000,I2859,I549675,I549664,);
not I_32185 (I550031,I549983);
DFFARX1 I_32186 (I550031,I2859,I549675,I550057,);
not I_32187 (I550065,I550057);
nor I_32188 (I549661,I550065,I549983);
nor I_32189 (I550096,I549966,I17853);
and I_32190 (I550113,I550096,I17850);
or I_32191 (I550130,I550113,I17832);
DFFARX1 I_32192 (I550130,I2859,I549675,I550156,);
not I_32193 (I550164,I550156);
nand I_32194 (I550181,I550164,I549904);
not I_32195 (I549655,I550181);
nand I_32196 (I549649,I550181,I549921);
nand I_32197 (I549646,I550164,I549788);
not I_32198 (I550270,I2866);
DFFARX1 I_32199 (I119272,I2859,I550270,I550296,);
DFFARX1 I_32200 (I119266,I2859,I550270,I550313,);
not I_32201 (I550321,I550313);
nor I_32202 (I550238,I550296,I550321);
DFFARX1 I_32203 (I550321,I2859,I550270,I550253,);
nor I_32204 (I550366,I119254,I119275);
and I_32205 (I550383,I550366,I119269);
nor I_32206 (I550400,I550383,I119254);
not I_32207 (I550417,I119254);
and I_32208 (I550434,I550417,I119251);
nand I_32209 (I550451,I550434,I119263);
nor I_32210 (I550468,I550417,I550451);
DFFARX1 I_32211 (I550468,I2859,I550270,I550235,);
not I_32212 (I550499,I550451);
nand I_32213 (I550516,I550321,I550499);
nand I_32214 (I550247,I550383,I550499);
DFFARX1 I_32215 (I550417,I2859,I550270,I550262,);
not I_32216 (I550561,I119278);
nor I_32217 (I550578,I550561,I119251);
nor I_32218 (I550595,I550578,I550400);
DFFARX1 I_32219 (I550595,I2859,I550270,I550259,);
not I_32220 (I550626,I550578);
DFFARX1 I_32221 (I550626,I2859,I550270,I550652,);
not I_32222 (I550660,I550652);
nor I_32223 (I550256,I550660,I550578);
nor I_32224 (I550691,I550561,I119260);
and I_32225 (I550708,I550691,I119257);
or I_32226 (I550725,I550708,I119251);
DFFARX1 I_32227 (I550725,I2859,I550270,I550751,);
not I_32228 (I550759,I550751);
nand I_32229 (I550776,I550759,I550499);
not I_32230 (I550250,I550776);
nand I_32231 (I550244,I550776,I550516);
nand I_32232 (I550241,I550759,I550383);
not I_32233 (I550865,I2866);
DFFARX1 I_32234 (I509690,I2859,I550865,I550891,);
DFFARX1 I_32235 (I509693,I2859,I550865,I550908,);
not I_32236 (I550916,I550908);
nor I_32237 (I550833,I550891,I550916);
DFFARX1 I_32238 (I550916,I2859,I550865,I550848,);
nor I_32239 (I550961,I509693,I509708);
and I_32240 (I550978,I550961,I509702);
nor I_32241 (I550995,I550978,I509693);
not I_32242 (I551012,I509693);
and I_32243 (I551029,I551012,I509711);
nand I_32244 (I551046,I551029,I509699);
nor I_32245 (I551063,I551012,I551046);
DFFARX1 I_32246 (I551063,I2859,I550865,I550830,);
not I_32247 (I551094,I551046);
nand I_32248 (I551111,I550916,I551094);
nand I_32249 (I550842,I550978,I551094);
DFFARX1 I_32250 (I551012,I2859,I550865,I550857,);
not I_32251 (I551156,I509705);
nor I_32252 (I551173,I551156,I509711);
nor I_32253 (I551190,I551173,I550995);
DFFARX1 I_32254 (I551190,I2859,I550865,I550854,);
not I_32255 (I551221,I551173);
DFFARX1 I_32256 (I551221,I2859,I550865,I551247,);
not I_32257 (I551255,I551247);
nor I_32258 (I550851,I551255,I551173);
nor I_32259 (I551286,I551156,I509690);
and I_32260 (I551303,I551286,I509714);
or I_32261 (I551320,I551303,I509696);
DFFARX1 I_32262 (I551320,I2859,I550865,I551346,);
not I_32263 (I551354,I551346);
nand I_32264 (I551371,I551354,I551094);
not I_32265 (I550845,I551371);
nand I_32266 (I550839,I551371,I551111);
nand I_32267 (I550836,I551354,I550978);
not I_32268 (I551460,I2866);
DFFARX1 I_32269 (I36822,I2859,I551460,I551486,);
DFFARX1 I_32270 (I36810,I2859,I551460,I551503,);
not I_32271 (I551511,I551503);
nor I_32272 (I551428,I551486,I551511);
DFFARX1 I_32273 (I551511,I2859,I551460,I551443,);
nor I_32274 (I551556,I36801,I36825);
and I_32275 (I551573,I551556,I36804);
nor I_32276 (I551590,I551573,I36801);
not I_32277 (I551607,I36801);
and I_32278 (I551624,I551607,I36807);
nand I_32279 (I551641,I551624,I36819);
nor I_32280 (I551658,I551607,I551641);
DFFARX1 I_32281 (I551658,I2859,I551460,I551425,);
not I_32282 (I551689,I551641);
nand I_32283 (I551706,I551511,I551689);
nand I_32284 (I551437,I551573,I551689);
DFFARX1 I_32285 (I551607,I2859,I551460,I551452,);
not I_32286 (I551751,I36801);
nor I_32287 (I551768,I551751,I36807);
nor I_32288 (I551785,I551768,I551590);
DFFARX1 I_32289 (I551785,I2859,I551460,I551449,);
not I_32290 (I551816,I551768);
DFFARX1 I_32291 (I551816,I2859,I551460,I551842,);
not I_32292 (I551850,I551842);
nor I_32293 (I551446,I551850,I551768);
nor I_32294 (I551881,I551751,I36804);
and I_32295 (I551898,I551881,I36813);
or I_32296 (I551915,I551898,I36816);
DFFARX1 I_32297 (I551915,I2859,I551460,I551941,);
not I_32298 (I551949,I551941);
nand I_32299 (I551966,I551949,I551689);
not I_32300 (I551440,I551966);
nand I_32301 (I551434,I551966,I551706);
nand I_32302 (I551431,I551949,I551573);
not I_32303 (I552055,I2866);
DFFARX1 I_32304 (I203163,I2859,I552055,I552081,);
DFFARX1 I_32305 (I203169,I2859,I552055,I552098,);
not I_32306 (I552106,I552098);
nor I_32307 (I552023,I552081,I552106);
DFFARX1 I_32308 (I552106,I2859,I552055,I552038,);
nor I_32309 (I552151,I203178,I203163);
and I_32310 (I552168,I552151,I203190);
nor I_32311 (I552185,I552168,I203178);
not I_32312 (I552202,I203178);
and I_32313 (I552219,I552202,I203166);
nand I_32314 (I552236,I552219,I203187);
nor I_32315 (I552253,I552202,I552236);
DFFARX1 I_32316 (I552253,I2859,I552055,I552020,);
not I_32317 (I552284,I552236);
nand I_32318 (I552301,I552106,I552284);
nand I_32319 (I552032,I552168,I552284);
DFFARX1 I_32320 (I552202,I2859,I552055,I552047,);
not I_32321 (I552346,I203175);
nor I_32322 (I552363,I552346,I203166);
nor I_32323 (I552380,I552363,I552185);
DFFARX1 I_32324 (I552380,I2859,I552055,I552044,);
not I_32325 (I552411,I552363);
DFFARX1 I_32326 (I552411,I2859,I552055,I552437,);
not I_32327 (I552445,I552437);
nor I_32328 (I552041,I552445,I552363);
nor I_32329 (I552476,I552346,I203172);
and I_32330 (I552493,I552476,I203184);
or I_32331 (I552510,I552493,I203181);
DFFARX1 I_32332 (I552510,I2859,I552055,I552536,);
not I_32333 (I552544,I552536);
nand I_32334 (I552561,I552544,I552284);
not I_32335 (I552035,I552561);
nand I_32336 (I552029,I552561,I552301);
nand I_32337 (I552026,I552544,I552168);
not I_32338 (I552650,I2866);
DFFARX1 I_32339 (I292213,I2859,I552650,I552676,);
DFFARX1 I_32340 (I292195,I2859,I552650,I552693,);
not I_32341 (I552701,I552693);
nor I_32342 (I552618,I552676,I552701);
DFFARX1 I_32343 (I552701,I2859,I552650,I552633,);
nor I_32344 (I552746,I292201,I292204);
and I_32345 (I552763,I552746,I292192);
nor I_32346 (I552780,I552763,I292201);
not I_32347 (I552797,I292201);
and I_32348 (I552814,I552797,I292210);
nand I_32349 (I552831,I552814,I292198);
nor I_32350 (I552848,I552797,I552831);
DFFARX1 I_32351 (I552848,I2859,I552650,I552615,);
not I_32352 (I552879,I552831);
nand I_32353 (I552896,I552701,I552879);
nand I_32354 (I552627,I552763,I552879);
DFFARX1 I_32355 (I552797,I2859,I552650,I552642,);
not I_32356 (I552941,I292195);
nor I_32357 (I552958,I552941,I292210);
nor I_32358 (I552975,I552958,I552780);
DFFARX1 I_32359 (I552975,I2859,I552650,I552639,);
not I_32360 (I553006,I552958);
DFFARX1 I_32361 (I553006,I2859,I552650,I553032,);
not I_32362 (I553040,I553032);
nor I_32363 (I552636,I553040,I552958);
nor I_32364 (I553071,I552941,I292207);
and I_32365 (I553088,I553071,I292216);
or I_32366 (I553105,I553088,I292192);
DFFARX1 I_32367 (I553105,I2859,I552650,I553131,);
not I_32368 (I553139,I553131);
nand I_32369 (I553156,I553139,I552879);
not I_32370 (I552630,I553156);
nand I_32371 (I552624,I553156,I552896);
nand I_32372 (I552621,I553139,I552763);
not I_32373 (I553245,I2866);
DFFARX1 I_32374 (I520026,I2859,I553245,I553271,);
DFFARX1 I_32375 (I520029,I2859,I553245,I553288,);
not I_32376 (I553296,I553288);
nor I_32377 (I553213,I553271,I553296);
DFFARX1 I_32378 (I553296,I2859,I553245,I553228,);
nor I_32379 (I553341,I520029,I520044);
and I_32380 (I553358,I553341,I520038);
nor I_32381 (I553375,I553358,I520029);
not I_32382 (I553392,I520029);
and I_32383 (I553409,I553392,I520047);
nand I_32384 (I553426,I553409,I520035);
nor I_32385 (I553443,I553392,I553426);
DFFARX1 I_32386 (I553443,I2859,I553245,I553210,);
not I_32387 (I553474,I553426);
nand I_32388 (I553491,I553296,I553474);
nand I_32389 (I553222,I553358,I553474);
DFFARX1 I_32390 (I553392,I2859,I553245,I553237,);
not I_32391 (I553536,I520041);
nor I_32392 (I553553,I553536,I520047);
nor I_32393 (I553570,I553553,I553375);
DFFARX1 I_32394 (I553570,I2859,I553245,I553234,);
not I_32395 (I553601,I553553);
DFFARX1 I_32396 (I553601,I2859,I553245,I553627,);
not I_32397 (I553635,I553627);
nor I_32398 (I553231,I553635,I553553);
nor I_32399 (I553666,I553536,I520026);
and I_32400 (I553683,I553666,I520050);
or I_32401 (I553700,I553683,I520032);
DFFARX1 I_32402 (I553700,I2859,I553245,I553726,);
not I_32403 (I553734,I553726);
nand I_32404 (I553751,I553734,I553474);
not I_32405 (I553225,I553751);
nand I_32406 (I553219,I553751,I553491);
nand I_32407 (I553216,I553734,I553358);
not I_32408 (I553840,I2866);
DFFARX1 I_32409 (I127177,I2859,I553840,I553866,);
DFFARX1 I_32410 (I127171,I2859,I553840,I553883,);
not I_32411 (I553891,I553883);
nor I_32412 (I553808,I553866,I553891);
DFFARX1 I_32413 (I553891,I2859,I553840,I553823,);
nor I_32414 (I553936,I127159,I127180);
and I_32415 (I553953,I553936,I127174);
nor I_32416 (I553970,I553953,I127159);
not I_32417 (I553987,I127159);
and I_32418 (I554004,I553987,I127156);
nand I_32419 (I554021,I554004,I127168);
nor I_32420 (I554038,I553987,I554021);
DFFARX1 I_32421 (I554038,I2859,I553840,I553805,);
not I_32422 (I554069,I554021);
nand I_32423 (I554086,I553891,I554069);
nand I_32424 (I553817,I553953,I554069);
DFFARX1 I_32425 (I553987,I2859,I553840,I553832,);
not I_32426 (I554131,I127183);
nor I_32427 (I554148,I554131,I127156);
nor I_32428 (I554165,I554148,I553970);
DFFARX1 I_32429 (I554165,I2859,I553840,I553829,);
not I_32430 (I554196,I554148);
DFFARX1 I_32431 (I554196,I2859,I553840,I554222,);
not I_32432 (I554230,I554222);
nor I_32433 (I553826,I554230,I554148);
nor I_32434 (I554261,I554131,I127165);
and I_32435 (I554278,I554261,I127162);
or I_32436 (I554295,I554278,I127156);
DFFARX1 I_32437 (I554295,I2859,I553840,I554321,);
not I_32438 (I554329,I554321);
nand I_32439 (I554346,I554329,I554069);
not I_32440 (I553820,I554346);
nand I_32441 (I553814,I554346,I554086);
nand I_32442 (I553811,I554329,I553953);
not I_32443 (I554435,I2866);
DFFARX1 I_32444 (I167259,I2859,I554435,I554461,);
DFFARX1 I_32445 (I167265,I2859,I554435,I554478,);
not I_32446 (I554486,I554478);
nor I_32447 (I554403,I554461,I554486);
DFFARX1 I_32448 (I554486,I2859,I554435,I554418,);
nor I_32449 (I554531,I167274,I167259);
and I_32450 (I554548,I554531,I167286);
nor I_32451 (I554565,I554548,I167274);
not I_32452 (I554582,I167274);
and I_32453 (I554599,I554582,I167262);
nand I_32454 (I554616,I554599,I167283);
nor I_32455 (I554633,I554582,I554616);
DFFARX1 I_32456 (I554633,I2859,I554435,I554400,);
not I_32457 (I554664,I554616);
nand I_32458 (I554681,I554486,I554664);
nand I_32459 (I554412,I554548,I554664);
DFFARX1 I_32460 (I554582,I2859,I554435,I554427,);
not I_32461 (I554726,I167271);
nor I_32462 (I554743,I554726,I167262);
nor I_32463 (I554760,I554743,I554565);
DFFARX1 I_32464 (I554760,I2859,I554435,I554424,);
not I_32465 (I554791,I554743);
DFFARX1 I_32466 (I554791,I2859,I554435,I554817,);
not I_32467 (I554825,I554817);
nor I_32468 (I554421,I554825,I554743);
nor I_32469 (I554856,I554726,I167268);
and I_32470 (I554873,I554856,I167280);
or I_32471 (I554890,I554873,I167277);
DFFARX1 I_32472 (I554890,I2859,I554435,I554916,);
not I_32473 (I554924,I554916);
nand I_32474 (I554941,I554924,I554664);
not I_32475 (I554415,I554941);
nand I_32476 (I554409,I554941,I554681);
nand I_32477 (I554406,I554924,I554548);
not I_32478 (I555030,I2866);
DFFARX1 I_32479 (I83993,I2859,I555030,I555056,);
DFFARX1 I_32480 (I83996,I2859,I555030,I555073,);
not I_32481 (I555081,I555073);
nor I_32482 (I554998,I555056,I555081);
DFFARX1 I_32483 (I555081,I2859,I555030,I555013,);
nor I_32484 (I555126,I84002,I83996);
and I_32485 (I555143,I555126,I83999);
nor I_32486 (I555160,I555143,I84002);
not I_32487 (I555177,I84002);
and I_32488 (I555194,I555177,I83993);
nand I_32489 (I555211,I555194,I84011);
nor I_32490 (I555228,I555177,I555211);
DFFARX1 I_32491 (I555228,I2859,I555030,I554995,);
not I_32492 (I555259,I555211);
nand I_32493 (I555276,I555081,I555259);
nand I_32494 (I555007,I555143,I555259);
DFFARX1 I_32495 (I555177,I2859,I555030,I555022,);
not I_32496 (I555321,I84005);
nor I_32497 (I555338,I555321,I83993);
nor I_32498 (I555355,I555338,I555160);
DFFARX1 I_32499 (I555355,I2859,I555030,I555019,);
not I_32500 (I555386,I555338);
DFFARX1 I_32501 (I555386,I2859,I555030,I555412,);
not I_32502 (I555420,I555412);
nor I_32503 (I555016,I555420,I555338);
nor I_32504 (I555451,I555321,I84008);
and I_32505 (I555468,I555451,I84014);
or I_32506 (I555485,I555468,I84017);
DFFARX1 I_32507 (I555485,I2859,I555030,I555511,);
not I_32508 (I555519,I555511);
nand I_32509 (I555536,I555519,I555259);
not I_32510 (I555010,I555536);
nand I_32511 (I555004,I555536,I555276);
nand I_32512 (I555001,I555519,I555143);
not I_32513 (I555625,I2866);
DFFARX1 I_32514 (I411929,I2859,I555625,I555651,);
DFFARX1 I_32515 (I411947,I2859,I555625,I555668,);
not I_32516 (I555676,I555668);
nor I_32517 (I555593,I555651,I555676);
DFFARX1 I_32518 (I555676,I2859,I555625,I555608,);
nor I_32519 (I555721,I411926,I411938);
and I_32520 (I555738,I555721,I411923);
nor I_32521 (I555755,I555738,I411926);
not I_32522 (I555772,I411926);
and I_32523 (I555789,I555772,I411932);
nand I_32524 (I555806,I555789,I411944);
nor I_32525 (I555823,I555772,I555806);
DFFARX1 I_32526 (I555823,I2859,I555625,I555590,);
not I_32527 (I555854,I555806);
nand I_32528 (I555871,I555676,I555854);
nand I_32529 (I555602,I555738,I555854);
DFFARX1 I_32530 (I555772,I2859,I555625,I555617,);
not I_32531 (I555916,I411935);
nor I_32532 (I555933,I555916,I411932);
nor I_32533 (I555950,I555933,I555755);
DFFARX1 I_32534 (I555950,I2859,I555625,I555614,);
not I_32535 (I555981,I555933);
DFFARX1 I_32536 (I555981,I2859,I555625,I556007,);
not I_32537 (I556015,I556007);
nor I_32538 (I555611,I556015,I555933);
nor I_32539 (I556046,I555916,I411923);
and I_32540 (I556063,I556046,I411950);
or I_32541 (I556080,I556063,I411941);
DFFARX1 I_32542 (I556080,I2859,I555625,I556106,);
not I_32543 (I556114,I556106);
nand I_32544 (I556131,I556114,I555854);
not I_32545 (I555605,I556131);
nand I_32546 (I555599,I556131,I555871);
nand I_32547 (I555596,I556114,I555738);
not I_32548 (I556220,I2866);
DFFARX1 I_32549 (I141933,I2859,I556220,I556246,);
DFFARX1 I_32550 (I141927,I2859,I556220,I556263,);
not I_32551 (I556271,I556263);
nor I_32552 (I556188,I556246,I556271);
DFFARX1 I_32553 (I556271,I2859,I556220,I556203,);
nor I_32554 (I556316,I141915,I141936);
and I_32555 (I556333,I556316,I141930);
nor I_32556 (I556350,I556333,I141915);
not I_32557 (I556367,I141915);
and I_32558 (I556384,I556367,I141912);
nand I_32559 (I556401,I556384,I141924);
nor I_32560 (I556418,I556367,I556401);
DFFARX1 I_32561 (I556418,I2859,I556220,I556185,);
not I_32562 (I556449,I556401);
nand I_32563 (I556466,I556271,I556449);
nand I_32564 (I556197,I556333,I556449);
DFFARX1 I_32565 (I556367,I2859,I556220,I556212,);
not I_32566 (I556511,I141939);
nor I_32567 (I556528,I556511,I141912);
nor I_32568 (I556545,I556528,I556350);
DFFARX1 I_32569 (I556545,I2859,I556220,I556209,);
not I_32570 (I556576,I556528);
DFFARX1 I_32571 (I556576,I2859,I556220,I556602,);
not I_32572 (I556610,I556602);
nor I_32573 (I556206,I556610,I556528);
nor I_32574 (I556641,I556511,I141921);
and I_32575 (I556658,I556641,I141918);
or I_32576 (I556675,I556658,I141912);
DFFARX1 I_32577 (I556675,I2859,I556220,I556701,);
not I_32578 (I556709,I556701);
nand I_32579 (I556726,I556709,I556449);
not I_32580 (I556200,I556726);
nand I_32581 (I556194,I556726,I556466);
nand I_32582 (I556191,I556709,I556333);
not I_32583 (I556815,I2866);
DFFARX1 I_32584 (I478379,I2859,I556815,I556841,);
DFFARX1 I_32585 (I478391,I2859,I556815,I556858,);
not I_32586 (I556866,I556858);
nor I_32587 (I556783,I556841,I556866);
DFFARX1 I_32588 (I556866,I2859,I556815,I556798,);
nor I_32589 (I556911,I478388,I478382);
and I_32590 (I556928,I556911,I478376);
nor I_32591 (I556945,I556928,I478388);
not I_32592 (I556962,I478388);
and I_32593 (I556979,I556962,I478385);
nand I_32594 (I556996,I556979,I478376);
nor I_32595 (I557013,I556962,I556996);
DFFARX1 I_32596 (I557013,I2859,I556815,I556780,);
not I_32597 (I557044,I556996);
nand I_32598 (I557061,I556866,I557044);
nand I_32599 (I556792,I556928,I557044);
DFFARX1 I_32600 (I556962,I2859,I556815,I556807,);
not I_32601 (I557106,I478400);
nor I_32602 (I557123,I557106,I478385);
nor I_32603 (I557140,I557123,I556945);
DFFARX1 I_32604 (I557140,I2859,I556815,I556804,);
not I_32605 (I557171,I557123);
DFFARX1 I_32606 (I557171,I2859,I556815,I557197,);
not I_32607 (I557205,I557197);
nor I_32608 (I556801,I557205,I557123);
nor I_32609 (I557236,I557106,I478394);
and I_32610 (I557253,I557236,I478397);
or I_32611 (I557270,I557253,I478379);
DFFARX1 I_32612 (I557270,I2859,I556815,I557296,);
not I_32613 (I557304,I557296);
nand I_32614 (I557321,I557304,I557044);
not I_32615 (I556795,I557321);
nand I_32616 (I556789,I557321,I557061);
nand I_32617 (I556786,I557304,I556928);
not I_32618 (I557410,I2866);
DFFARX1 I_32619 (I131920,I2859,I557410,I557436,);
DFFARX1 I_32620 (I131914,I2859,I557410,I557453,);
not I_32621 (I557461,I557453);
nor I_32622 (I557378,I557436,I557461);
DFFARX1 I_32623 (I557461,I2859,I557410,I557393,);
nor I_32624 (I557506,I131902,I131923);
and I_32625 (I557523,I557506,I131917);
nor I_32626 (I557540,I557523,I131902);
not I_32627 (I557557,I131902);
and I_32628 (I557574,I557557,I131899);
nand I_32629 (I557591,I557574,I131911);
nor I_32630 (I557608,I557557,I557591);
DFFARX1 I_32631 (I557608,I2859,I557410,I557375,);
not I_32632 (I557639,I557591);
nand I_32633 (I557656,I557461,I557639);
nand I_32634 (I557387,I557523,I557639);
DFFARX1 I_32635 (I557557,I2859,I557410,I557402,);
not I_32636 (I557701,I131926);
nor I_32637 (I557718,I557701,I131899);
nor I_32638 (I557735,I557718,I557540);
DFFARX1 I_32639 (I557735,I2859,I557410,I557399,);
not I_32640 (I557766,I557718);
DFFARX1 I_32641 (I557766,I2859,I557410,I557792,);
not I_32642 (I557800,I557792);
nor I_32643 (I557396,I557800,I557718);
nor I_32644 (I557831,I557701,I131908);
and I_32645 (I557848,I557831,I131905);
or I_32646 (I557865,I557848,I131899);
DFFARX1 I_32647 (I557865,I2859,I557410,I557891,);
not I_32648 (I557899,I557891);
nand I_32649 (I557916,I557899,I557639);
not I_32650 (I557390,I557916);
nand I_32651 (I557384,I557916,I557656);
nand I_32652 (I557381,I557899,I557523);
not I_32653 (I558005,I2866);
DFFARX1 I_32654 (I274295,I2859,I558005,I558031,);
DFFARX1 I_32655 (I274277,I2859,I558005,I558048,);
not I_32656 (I558056,I558048);
nor I_32657 (I557973,I558031,I558056);
DFFARX1 I_32658 (I558056,I2859,I558005,I557988,);
nor I_32659 (I558101,I274283,I274286);
and I_32660 (I558118,I558101,I274274);
nor I_32661 (I558135,I558118,I274283);
not I_32662 (I558152,I274283);
and I_32663 (I558169,I558152,I274292);
nand I_32664 (I558186,I558169,I274280);
nor I_32665 (I558203,I558152,I558186);
DFFARX1 I_32666 (I558203,I2859,I558005,I557970,);
not I_32667 (I558234,I558186);
nand I_32668 (I558251,I558056,I558234);
nand I_32669 (I557982,I558118,I558234);
DFFARX1 I_32670 (I558152,I2859,I558005,I557997,);
not I_32671 (I558296,I274277);
nor I_32672 (I558313,I558296,I274292);
nor I_32673 (I558330,I558313,I558135);
DFFARX1 I_32674 (I558330,I2859,I558005,I557994,);
not I_32675 (I558361,I558313);
DFFARX1 I_32676 (I558361,I2859,I558005,I558387,);
not I_32677 (I558395,I558387);
nor I_32678 (I557991,I558395,I558313);
nor I_32679 (I558426,I558296,I274289);
and I_32680 (I558443,I558426,I274298);
or I_32681 (I558460,I558443,I274274);
DFFARX1 I_32682 (I558460,I2859,I558005,I558486,);
not I_32683 (I558494,I558486);
nand I_32684 (I558511,I558494,I558234);
not I_32685 (I557985,I558511);
nand I_32686 (I557979,I558511,I558251);
nand I_32687 (I557976,I558494,I558118);
not I_32688 (I558600,I2866);
DFFARX1 I_32689 (I390611,I2859,I558600,I558626,);
DFFARX1 I_32690 (I390629,I2859,I558600,I558643,);
not I_32691 (I558651,I558643);
nor I_32692 (I558568,I558626,I558651);
DFFARX1 I_32693 (I558651,I2859,I558600,I558583,);
nor I_32694 (I558696,I390608,I390620);
and I_32695 (I558713,I558696,I390605);
nor I_32696 (I558730,I558713,I390608);
not I_32697 (I558747,I390608);
and I_32698 (I558764,I558747,I390614);
nand I_32699 (I558781,I558764,I390626);
nor I_32700 (I558798,I558747,I558781);
DFFARX1 I_32701 (I558798,I2859,I558600,I558565,);
not I_32702 (I558829,I558781);
nand I_32703 (I558846,I558651,I558829);
nand I_32704 (I558577,I558713,I558829);
DFFARX1 I_32705 (I558747,I2859,I558600,I558592,);
not I_32706 (I558891,I390617);
nor I_32707 (I558908,I558891,I390614);
nor I_32708 (I558925,I558908,I558730);
DFFARX1 I_32709 (I558925,I2859,I558600,I558589,);
not I_32710 (I558956,I558908);
DFFARX1 I_32711 (I558956,I2859,I558600,I558982,);
not I_32712 (I558990,I558982);
nor I_32713 (I558586,I558990,I558908);
nor I_32714 (I559021,I558891,I390605);
and I_32715 (I559038,I559021,I390632);
or I_32716 (I559055,I559038,I390623);
DFFARX1 I_32717 (I559055,I2859,I558600,I559081,);
not I_32718 (I559089,I559081);
nand I_32719 (I559106,I559089,I558829);
not I_32720 (I558580,I559106);
nand I_32721 (I558574,I559106,I558846);
nand I_32722 (I558571,I559089,I558713);
not I_32723 (I559195,I2866);
DFFARX1 I_32724 (I472599,I2859,I559195,I559221,);
DFFARX1 I_32725 (I472611,I2859,I559195,I559238,);
not I_32726 (I559246,I559238);
nor I_32727 (I559163,I559221,I559246);
DFFARX1 I_32728 (I559246,I2859,I559195,I559178,);
nor I_32729 (I559291,I472608,I472602);
and I_32730 (I559308,I559291,I472596);
nor I_32731 (I559325,I559308,I472608);
not I_32732 (I559342,I472608);
and I_32733 (I559359,I559342,I472605);
nand I_32734 (I559376,I559359,I472596);
nor I_32735 (I559393,I559342,I559376);
DFFARX1 I_32736 (I559393,I2859,I559195,I559160,);
not I_32737 (I559424,I559376);
nand I_32738 (I559441,I559246,I559424);
nand I_32739 (I559172,I559308,I559424);
DFFARX1 I_32740 (I559342,I2859,I559195,I559187,);
not I_32741 (I559486,I472620);
nor I_32742 (I559503,I559486,I472605);
nor I_32743 (I559520,I559503,I559325);
DFFARX1 I_32744 (I559520,I2859,I559195,I559184,);
not I_32745 (I559551,I559503);
DFFARX1 I_32746 (I559551,I2859,I559195,I559577,);
not I_32747 (I559585,I559577);
nor I_32748 (I559181,I559585,I559503);
nor I_32749 (I559616,I559486,I472614);
and I_32750 (I559633,I559616,I472617);
or I_32751 (I559650,I559633,I472599);
DFFARX1 I_32752 (I559650,I2859,I559195,I559676,);
not I_32753 (I559684,I559676);
nand I_32754 (I559701,I559684,I559424);
not I_32755 (I559175,I559701);
nand I_32756 (I559169,I559701,I559441);
nand I_32757 (I559166,I559684,I559308);
not I_32758 (I559790,I2866);
DFFARX1 I_32759 (I28917,I2859,I559790,I559816,);
DFFARX1 I_32760 (I28905,I2859,I559790,I559833,);
not I_32761 (I559841,I559833);
nor I_32762 (I559758,I559816,I559841);
DFFARX1 I_32763 (I559841,I2859,I559790,I559773,);
nor I_32764 (I559886,I28896,I28920);
and I_32765 (I559903,I559886,I28899);
nor I_32766 (I559920,I559903,I28896);
not I_32767 (I559937,I28896);
and I_32768 (I559954,I559937,I28902);
nand I_32769 (I559971,I559954,I28914);
nor I_32770 (I559988,I559937,I559971);
DFFARX1 I_32771 (I559988,I2859,I559790,I559755,);
not I_32772 (I560019,I559971);
nand I_32773 (I560036,I559841,I560019);
nand I_32774 (I559767,I559903,I560019);
DFFARX1 I_32775 (I559937,I2859,I559790,I559782,);
not I_32776 (I560081,I28896);
nor I_32777 (I560098,I560081,I28902);
nor I_32778 (I560115,I560098,I559920);
DFFARX1 I_32779 (I560115,I2859,I559790,I559779,);
not I_32780 (I560146,I560098);
DFFARX1 I_32781 (I560146,I2859,I559790,I560172,);
not I_32782 (I560180,I560172);
nor I_32783 (I559776,I560180,I560098);
nor I_32784 (I560211,I560081,I28899);
and I_32785 (I560228,I560211,I28908);
or I_32786 (I560245,I560228,I28911);
DFFARX1 I_32787 (I560245,I2859,I559790,I560271,);
not I_32788 (I560279,I560271);
nand I_32789 (I560296,I560279,I560019);
not I_32790 (I559770,I560296);
nand I_32791 (I559764,I560296,I560036);
nand I_32792 (I559761,I560279,I559903);
not I_32793 (I560385,I2866);
DFFARX1 I_32794 (I515674,I2859,I560385,I560411,);
DFFARX1 I_32795 (I515677,I2859,I560385,I560428,);
not I_32796 (I560436,I560428);
nor I_32797 (I560353,I560411,I560436);
DFFARX1 I_32798 (I560436,I2859,I560385,I560368,);
nor I_32799 (I560481,I515677,I515692);
and I_32800 (I560498,I560481,I515686);
nor I_32801 (I560515,I560498,I515677);
not I_32802 (I560532,I515677);
and I_32803 (I560549,I560532,I515695);
nand I_32804 (I560566,I560549,I515683);
nor I_32805 (I560583,I560532,I560566);
DFFARX1 I_32806 (I560583,I2859,I560385,I560350,);
not I_32807 (I560614,I560566);
nand I_32808 (I560631,I560436,I560614);
nand I_32809 (I560362,I560498,I560614);
DFFARX1 I_32810 (I560532,I2859,I560385,I560377,);
not I_32811 (I560676,I515689);
nor I_32812 (I560693,I560676,I515695);
nor I_32813 (I560710,I560693,I560515);
DFFARX1 I_32814 (I560710,I2859,I560385,I560374,);
not I_32815 (I560741,I560693);
DFFARX1 I_32816 (I560741,I2859,I560385,I560767,);
not I_32817 (I560775,I560767);
nor I_32818 (I560371,I560775,I560693);
nor I_32819 (I560806,I560676,I515674);
and I_32820 (I560823,I560806,I515698);
or I_32821 (I560840,I560823,I515680);
DFFARX1 I_32822 (I560840,I2859,I560385,I560866,);
not I_32823 (I560874,I560866);
nand I_32824 (I560891,I560874,I560614);
not I_32825 (I560365,I560891);
nand I_32826 (I560359,I560891,I560631);
nand I_32827 (I560356,I560874,I560498);
not I_32828 (I560980,I2866);
DFFARX1 I_32829 (I231523,I2859,I560980,I561006,);
DFFARX1 I_32830 (I231517,I2859,I560980,I561023,);
not I_32831 (I561031,I561023);
nor I_32832 (I560948,I561006,I561031);
DFFARX1 I_32833 (I561031,I2859,I560980,I560963,);
nor I_32834 (I561076,I231514,I231505);
and I_32835 (I561093,I561076,I231502);
nor I_32836 (I561110,I561093,I231514);
not I_32837 (I561127,I231514);
and I_32838 (I561144,I561127,I231508);
nand I_32839 (I561161,I561144,I231520);
nor I_32840 (I561178,I561127,I561161);
DFFARX1 I_32841 (I561178,I2859,I560980,I560945,);
not I_32842 (I561209,I561161);
nand I_32843 (I561226,I561031,I561209);
nand I_32844 (I560957,I561093,I561209);
DFFARX1 I_32845 (I561127,I2859,I560980,I560972,);
not I_32846 (I561271,I231526);
nor I_32847 (I561288,I561271,I231508);
nor I_32848 (I561305,I561288,I561110);
DFFARX1 I_32849 (I561305,I2859,I560980,I560969,);
not I_32850 (I561336,I561288);
DFFARX1 I_32851 (I561336,I2859,I560980,I561362,);
not I_32852 (I561370,I561362);
nor I_32853 (I560966,I561370,I561288);
nor I_32854 (I561401,I561271,I231505);
and I_32855 (I561418,I561401,I231511);
or I_32856 (I561435,I561418,I231502);
DFFARX1 I_32857 (I561435,I2859,I560980,I561461,);
not I_32858 (I561469,I561461);
nand I_32859 (I561486,I561469,I561209);
not I_32860 (I560960,I561486);
nand I_32861 (I560954,I561486,I561226);
nand I_32862 (I560951,I561469,I561093);
not I_32863 (I561575,I2866);
DFFARX1 I_32864 (I507514,I2859,I561575,I561601,);
DFFARX1 I_32865 (I507517,I2859,I561575,I561618,);
not I_32866 (I561626,I561618);
nor I_32867 (I561543,I561601,I561626);
DFFARX1 I_32868 (I561626,I2859,I561575,I561558,);
nor I_32869 (I561671,I507517,I507532);
and I_32870 (I561688,I561671,I507526);
nor I_32871 (I561705,I561688,I507517);
not I_32872 (I561722,I507517);
and I_32873 (I561739,I561722,I507535);
nand I_32874 (I561756,I561739,I507523);
nor I_32875 (I561773,I561722,I561756);
DFFARX1 I_32876 (I561773,I2859,I561575,I561540,);
not I_32877 (I561804,I561756);
nand I_32878 (I561821,I561626,I561804);
nand I_32879 (I561552,I561688,I561804);
DFFARX1 I_32880 (I561722,I2859,I561575,I561567,);
not I_32881 (I561866,I507529);
nor I_32882 (I561883,I561866,I507535);
nor I_32883 (I561900,I561883,I561705);
DFFARX1 I_32884 (I561900,I2859,I561575,I561564,);
not I_32885 (I561931,I561883);
DFFARX1 I_32886 (I561931,I2859,I561575,I561957,);
not I_32887 (I561965,I561957);
nor I_32888 (I561561,I561965,I561883);
nor I_32889 (I561996,I561866,I507514);
and I_32890 (I562013,I561996,I507538);
or I_32891 (I562030,I562013,I507520);
DFFARX1 I_32892 (I562030,I2859,I561575,I562056,);
not I_32893 (I562064,I562056);
nand I_32894 (I562081,I562064,I561804);
not I_32895 (I561555,I562081);
nand I_32896 (I561549,I562081,I561821);
nand I_32897 (I561546,I562064,I561688);
not I_32898 (I562170,I2866);
DFFARX1 I_32899 (I1756,I2859,I562170,I562196,);
DFFARX1 I_32900 (I1500,I2859,I562170,I562213,);
not I_32901 (I562221,I562213);
nor I_32902 (I562138,I562196,I562221);
DFFARX1 I_32903 (I562221,I2859,I562170,I562153,);
nor I_32904 (I562266,I2604,I2428);
and I_32905 (I562283,I562266,I1596);
nor I_32906 (I562300,I562283,I2604);
not I_32907 (I562317,I2604);
and I_32908 (I562334,I562317,I1628);
nand I_32909 (I562351,I562334,I2332);
nor I_32910 (I562368,I562317,I562351);
DFFARX1 I_32911 (I562368,I2859,I562170,I562135,);
not I_32912 (I562399,I562351);
nand I_32913 (I562416,I562221,I562399);
nand I_32914 (I562147,I562283,I562399);
DFFARX1 I_32915 (I562317,I2859,I562170,I562162,);
not I_32916 (I562461,I2204);
nor I_32917 (I562478,I562461,I1628);
nor I_32918 (I562495,I562478,I562300);
DFFARX1 I_32919 (I562495,I2859,I562170,I562159,);
not I_32920 (I562526,I562478);
DFFARX1 I_32921 (I562526,I2859,I562170,I562552,);
not I_32922 (I562560,I562552);
nor I_32923 (I562156,I562560,I562478);
nor I_32924 (I562591,I562461,I2148);
and I_32925 (I562608,I562591,I2372);
or I_32926 (I562625,I562608,I1364);
DFFARX1 I_32927 (I562625,I2859,I562170,I562651,);
not I_32928 (I562659,I562651);
nand I_32929 (I562676,I562659,I562399);
not I_32930 (I562150,I562676);
nand I_32931 (I562144,I562676,I562416);
nand I_32932 (I562141,I562659,I562283);
not I_32933 (I562765,I2866);
DFFARX1 I_32934 (I144041,I2859,I562765,I562791,);
DFFARX1 I_32935 (I144035,I2859,I562765,I562808,);
not I_32936 (I562816,I562808);
nor I_32937 (I562733,I562791,I562816);
DFFARX1 I_32938 (I562816,I2859,I562765,I562748,);
nor I_32939 (I562861,I144023,I144044);
and I_32940 (I562878,I562861,I144038);
nor I_32941 (I562895,I562878,I144023);
not I_32942 (I562912,I144023);
and I_32943 (I562929,I562912,I144020);
nand I_32944 (I562946,I562929,I144032);
nor I_32945 (I562963,I562912,I562946);
DFFARX1 I_32946 (I562963,I2859,I562765,I562730,);
not I_32947 (I562994,I562946);
nand I_32948 (I563011,I562816,I562994);
nand I_32949 (I562742,I562878,I562994);
DFFARX1 I_32950 (I562912,I2859,I562765,I562757,);
not I_32951 (I563056,I144047);
nor I_32952 (I563073,I563056,I144020);
nor I_32953 (I563090,I563073,I562895);
DFFARX1 I_32954 (I563090,I2859,I562765,I562754,);
not I_32955 (I563121,I563073);
DFFARX1 I_32956 (I563121,I2859,I562765,I563147,);
not I_32957 (I563155,I563147);
nor I_32958 (I562751,I563155,I563073);
nor I_32959 (I563186,I563056,I144029);
and I_32960 (I563203,I563186,I144026);
or I_32961 (I563220,I563203,I144020);
DFFARX1 I_32962 (I563220,I2859,I562765,I563246,);
not I_32963 (I563254,I563246);
nand I_32964 (I563271,I563254,I562994);
not I_32965 (I562745,I563271);
nand I_32966 (I562739,I563271,I563011);
nand I_32967 (I562736,I563254,I562878);
not I_32968 (I563360,I2866);
DFFARX1 I_32969 (I186299,I2859,I563360,I563386,);
DFFARX1 I_32970 (I186305,I2859,I563360,I563403,);
not I_32971 (I563411,I563403);
nor I_32972 (I563328,I563386,I563411);
DFFARX1 I_32973 (I563411,I2859,I563360,I563343,);
nor I_32974 (I563456,I186314,I186299);
and I_32975 (I563473,I563456,I186326);
nor I_32976 (I563490,I563473,I186314);
not I_32977 (I563507,I186314);
and I_32978 (I563524,I563507,I186302);
nand I_32979 (I563541,I563524,I186323);
nor I_32980 (I563558,I563507,I563541);
DFFARX1 I_32981 (I563558,I2859,I563360,I563325,);
not I_32982 (I563589,I563541);
nand I_32983 (I563606,I563411,I563589);
nand I_32984 (I563337,I563473,I563589);
DFFARX1 I_32985 (I563507,I2859,I563360,I563352,);
not I_32986 (I563651,I186311);
nor I_32987 (I563668,I563651,I186302);
nor I_32988 (I563685,I563668,I563490);
DFFARX1 I_32989 (I563685,I2859,I563360,I563349,);
not I_32990 (I563716,I563668);
DFFARX1 I_32991 (I563716,I2859,I563360,I563742,);
not I_32992 (I563750,I563742);
nor I_32993 (I563346,I563750,I563668);
nor I_32994 (I563781,I563651,I186308);
and I_32995 (I563798,I563781,I186320);
or I_32996 (I563815,I563798,I186317);
DFFARX1 I_32997 (I563815,I2859,I563360,I563841,);
not I_32998 (I563849,I563841);
nand I_32999 (I563866,I563849,I563589);
not I_33000 (I563340,I563866);
nand I_33001 (I563334,I563866,I563606);
nand I_33002 (I563331,I563849,I563473);
not I_33003 (I563955,I2866);
DFFARX1 I_33004 (I298571,I2859,I563955,I563981,);
DFFARX1 I_33005 (I298553,I2859,I563955,I563998,);
not I_33006 (I564006,I563998);
nor I_33007 (I563923,I563981,I564006);
DFFARX1 I_33008 (I564006,I2859,I563955,I563938,);
nor I_33009 (I564051,I298559,I298562);
and I_33010 (I564068,I564051,I298550);
nor I_33011 (I564085,I564068,I298559);
not I_33012 (I564102,I298559);
and I_33013 (I564119,I564102,I298568);
nand I_33014 (I564136,I564119,I298556);
nor I_33015 (I564153,I564102,I564136);
DFFARX1 I_33016 (I564153,I2859,I563955,I563920,);
not I_33017 (I564184,I564136);
nand I_33018 (I564201,I564006,I564184);
nand I_33019 (I563932,I564068,I564184);
DFFARX1 I_33020 (I564102,I2859,I563955,I563947,);
not I_33021 (I564246,I298553);
nor I_33022 (I564263,I564246,I298568);
nor I_33023 (I564280,I564263,I564085);
DFFARX1 I_33024 (I564280,I2859,I563955,I563944,);
not I_33025 (I564311,I564263);
DFFARX1 I_33026 (I564311,I2859,I563955,I564337,);
not I_33027 (I564345,I564337);
nor I_33028 (I563941,I564345,I564263);
nor I_33029 (I564376,I564246,I298565);
and I_33030 (I564393,I564376,I298574);
or I_33031 (I564410,I564393,I298550);
DFFARX1 I_33032 (I564410,I2859,I563955,I564436,);
not I_33033 (I564444,I564436);
nand I_33034 (I564461,I564444,I564184);
not I_33035 (I563935,I564461);
nand I_33036 (I563929,I564461,I564201);
nand I_33037 (I563926,I564444,I564068);
not I_33038 (I564550,I2866);
DFFARX1 I_33039 (I533270,I2859,I564550,I564576,);
DFFARX1 I_33040 (I533261,I2859,I564550,I564593,);
not I_33041 (I564601,I564593);
nor I_33042 (I564518,I564576,I564601);
DFFARX1 I_33043 (I564601,I2859,I564550,I564533,);
nor I_33044 (I564646,I533252,I533267);
and I_33045 (I564663,I564646,I533255);
nor I_33046 (I564680,I564663,I533252);
not I_33047 (I564697,I533252);
and I_33048 (I564714,I564697,I533258);
nand I_33049 (I564731,I564714,I533276);
nor I_33050 (I564748,I564697,I564731);
DFFARX1 I_33051 (I564748,I2859,I564550,I564515,);
not I_33052 (I564779,I564731);
nand I_33053 (I564796,I564601,I564779);
nand I_33054 (I564527,I564663,I564779);
DFFARX1 I_33055 (I564697,I2859,I564550,I564542,);
not I_33056 (I564841,I533252);
nor I_33057 (I564858,I564841,I533258);
nor I_33058 (I564875,I564858,I564680);
DFFARX1 I_33059 (I564875,I2859,I564550,I564539,);
not I_33060 (I564906,I564858);
DFFARX1 I_33061 (I564906,I2859,I564550,I564932,);
not I_33062 (I564940,I564932);
nor I_33063 (I564536,I564940,I564858);
nor I_33064 (I564971,I564841,I533255);
and I_33065 (I564988,I564971,I533264);
or I_33066 (I565005,I564988,I533273);
DFFARX1 I_33067 (I565005,I2859,I564550,I565031,);
not I_33068 (I565039,I565031);
nand I_33069 (I565056,I565039,I564779);
not I_33070 (I564530,I565056);
nand I_33071 (I564524,I565056,I564796);
nand I_33072 (I564521,I565039,I564663);
not I_33073 (I565145,I2866);
DFFARX1 I_33074 (I364281,I2859,I565145,I565171,);
DFFARX1 I_33075 (I364278,I2859,I565145,I565188,);
not I_33076 (I565196,I565188);
nor I_33077 (I565113,I565171,I565196);
DFFARX1 I_33078 (I565196,I2859,I565145,I565128,);
nor I_33079 (I565241,I364293,I364275);
and I_33080 (I565258,I565241,I364272);
nor I_33081 (I565275,I565258,I364293);
not I_33082 (I565292,I364293);
and I_33083 (I565309,I565292,I364278);
nand I_33084 (I565326,I565309,I364290);
nor I_33085 (I565343,I565292,I565326);
DFFARX1 I_33086 (I565343,I2859,I565145,I565110,);
not I_33087 (I565374,I565326);
nand I_33088 (I565391,I565196,I565374);
nand I_33089 (I565122,I565258,I565374);
DFFARX1 I_33090 (I565292,I2859,I565145,I565137,);
not I_33091 (I565436,I364284);
nor I_33092 (I565453,I565436,I364278);
nor I_33093 (I565470,I565453,I565275);
DFFARX1 I_33094 (I565470,I2859,I565145,I565134,);
not I_33095 (I565501,I565453);
DFFARX1 I_33096 (I565501,I2859,I565145,I565527,);
not I_33097 (I565535,I565527);
nor I_33098 (I565131,I565535,I565453);
nor I_33099 (I565566,I565436,I364272);
and I_33100 (I565583,I565566,I364287);
or I_33101 (I565600,I565583,I364275);
DFFARX1 I_33102 (I565600,I2859,I565145,I565626,);
not I_33103 (I565634,I565626);
nand I_33104 (I565651,I565634,I565374);
not I_33105 (I565125,I565651);
nand I_33106 (I565119,I565651,I565391);
nand I_33107 (I565116,I565634,I565258);
not I_33108 (I565740,I2866);
DFFARX1 I_33109 (I197179,I2859,I565740,I565766,);
DFFARX1 I_33110 (I197185,I2859,I565740,I565783,);
not I_33111 (I565791,I565783);
nor I_33112 (I565708,I565766,I565791);
DFFARX1 I_33113 (I565791,I2859,I565740,I565723,);
nor I_33114 (I565836,I197194,I197179);
and I_33115 (I565853,I565836,I197206);
nor I_33116 (I565870,I565853,I197194);
not I_33117 (I565887,I197194);
and I_33118 (I565904,I565887,I197182);
nand I_33119 (I565921,I565904,I197203);
nor I_33120 (I565938,I565887,I565921);
DFFARX1 I_33121 (I565938,I2859,I565740,I565705,);
not I_33122 (I565969,I565921);
nand I_33123 (I565986,I565791,I565969);
nand I_33124 (I565717,I565853,I565969);
DFFARX1 I_33125 (I565887,I2859,I565740,I565732,);
not I_33126 (I566031,I197191);
nor I_33127 (I566048,I566031,I197182);
nor I_33128 (I566065,I566048,I565870);
DFFARX1 I_33129 (I566065,I2859,I565740,I565729,);
not I_33130 (I566096,I566048);
DFFARX1 I_33131 (I566096,I2859,I565740,I566122,);
not I_33132 (I566130,I566122);
nor I_33133 (I565726,I566130,I566048);
nor I_33134 (I566161,I566031,I197188);
and I_33135 (I566178,I566161,I197200);
or I_33136 (I566195,I566178,I197197);
DFFARX1 I_33137 (I566195,I2859,I565740,I566221,);
not I_33138 (I566229,I566221);
nand I_33139 (I566246,I566229,I565969);
not I_33140 (I565720,I566246);
nand I_33141 (I565714,I566246,I565986);
nand I_33142 (I565711,I566229,I565853);
not I_33143 (I566335,I2866);
DFFARX1 I_33144 (I154581,I2859,I566335,I566361,);
DFFARX1 I_33145 (I154575,I2859,I566335,I566378,);
not I_33146 (I566386,I566378);
nor I_33147 (I566303,I566361,I566386);
DFFARX1 I_33148 (I566386,I2859,I566335,I566318,);
nor I_33149 (I566431,I154563,I154584);
and I_33150 (I566448,I566431,I154578);
nor I_33151 (I566465,I566448,I154563);
not I_33152 (I566482,I154563);
and I_33153 (I566499,I566482,I154560);
nand I_33154 (I566516,I566499,I154572);
nor I_33155 (I566533,I566482,I566516);
DFFARX1 I_33156 (I566533,I2859,I566335,I566300,);
not I_33157 (I566564,I566516);
nand I_33158 (I566581,I566386,I566564);
nand I_33159 (I566312,I566448,I566564);
DFFARX1 I_33160 (I566482,I2859,I566335,I566327,);
not I_33161 (I566626,I154587);
nor I_33162 (I566643,I566626,I154560);
nor I_33163 (I566660,I566643,I566465);
DFFARX1 I_33164 (I566660,I2859,I566335,I566324,);
not I_33165 (I566691,I566643);
DFFARX1 I_33166 (I566691,I2859,I566335,I566717,);
not I_33167 (I566725,I566717);
nor I_33168 (I566321,I566725,I566643);
nor I_33169 (I566756,I566626,I154569);
and I_33170 (I566773,I566756,I154566);
or I_33171 (I566790,I566773,I154560);
DFFARX1 I_33172 (I566790,I2859,I566335,I566816,);
not I_33173 (I566824,I566816);
nand I_33174 (I566841,I566824,I566564);
not I_33175 (I566315,I566841);
nand I_33176 (I566309,I566841,I566581);
nand I_33177 (I566306,I566824,I566448);
not I_33178 (I566930,I2866);
DFFARX1 I_33179 (I73878,I2859,I566930,I566956,);
DFFARX1 I_33180 (I73881,I2859,I566930,I566973,);
not I_33181 (I566981,I566973);
nor I_33182 (I566898,I566956,I566981);
DFFARX1 I_33183 (I566981,I2859,I566930,I566913,);
nor I_33184 (I567026,I73887,I73881);
and I_33185 (I567043,I567026,I73884);
nor I_33186 (I567060,I567043,I73887);
not I_33187 (I567077,I73887);
and I_33188 (I567094,I567077,I73878);
nand I_33189 (I567111,I567094,I73896);
nor I_33190 (I567128,I567077,I567111);
DFFARX1 I_33191 (I567128,I2859,I566930,I566895,);
not I_33192 (I567159,I567111);
nand I_33193 (I567176,I566981,I567159);
nand I_33194 (I566907,I567043,I567159);
DFFARX1 I_33195 (I567077,I2859,I566930,I566922,);
not I_33196 (I567221,I73890);
nor I_33197 (I567238,I567221,I73878);
nor I_33198 (I567255,I567238,I567060);
DFFARX1 I_33199 (I567255,I2859,I566930,I566919,);
not I_33200 (I567286,I567238);
DFFARX1 I_33201 (I567286,I2859,I566930,I567312,);
not I_33202 (I567320,I567312);
nor I_33203 (I566916,I567320,I567238);
nor I_33204 (I567351,I567221,I73893);
and I_33205 (I567368,I567351,I73899);
or I_33206 (I567385,I567368,I73902);
DFFARX1 I_33207 (I567385,I2859,I566930,I567411,);
not I_33208 (I567419,I567411);
nand I_33209 (I567436,I567419,I567159);
not I_33210 (I566910,I567436);
nand I_33211 (I566904,I567436,I567176);
nand I_33212 (I566901,I567419,I567043);
not I_33213 (I567525,I2866);
DFFARX1 I_33214 (I343728,I2859,I567525,I567551,);
DFFARX1 I_33215 (I343725,I2859,I567525,I567568,);
not I_33216 (I567576,I567568);
nor I_33217 (I567493,I567551,I567576);
DFFARX1 I_33218 (I567576,I2859,I567525,I567508,);
nor I_33219 (I567621,I343740,I343722);
and I_33220 (I567638,I567621,I343719);
nor I_33221 (I567655,I567638,I343740);
not I_33222 (I567672,I343740);
and I_33223 (I567689,I567672,I343725);
nand I_33224 (I567706,I567689,I343737);
nor I_33225 (I567723,I567672,I567706);
DFFARX1 I_33226 (I567723,I2859,I567525,I567490,);
not I_33227 (I567754,I567706);
nand I_33228 (I567771,I567576,I567754);
nand I_33229 (I567502,I567638,I567754);
DFFARX1 I_33230 (I567672,I2859,I567525,I567517,);
not I_33231 (I567816,I343731);
nor I_33232 (I567833,I567816,I343725);
nor I_33233 (I567850,I567833,I567655);
DFFARX1 I_33234 (I567850,I2859,I567525,I567514,);
not I_33235 (I567881,I567833);
DFFARX1 I_33236 (I567881,I2859,I567525,I567907,);
not I_33237 (I567915,I567907);
nor I_33238 (I567511,I567915,I567833);
nor I_33239 (I567946,I567816,I343719);
and I_33240 (I567963,I567946,I343734);
or I_33241 (I567980,I567963,I343722);
DFFARX1 I_33242 (I567980,I2859,I567525,I568006,);
not I_33243 (I568014,I568006);
nand I_33244 (I568031,I568014,I567754);
not I_33245 (I567505,I568031);
nand I_33246 (I567499,I568031,I567771);
nand I_33247 (I567496,I568014,I567638);
not I_33248 (I568120,I2866);
DFFARX1 I_33249 (I280075,I2859,I568120,I568146,);
DFFARX1 I_33250 (I280057,I2859,I568120,I568163,);
not I_33251 (I568171,I568163);
nor I_33252 (I568088,I568146,I568171);
DFFARX1 I_33253 (I568171,I2859,I568120,I568103,);
nor I_33254 (I568216,I280063,I280066);
and I_33255 (I568233,I568216,I280054);
nor I_33256 (I568250,I568233,I280063);
not I_33257 (I568267,I280063);
and I_33258 (I568284,I568267,I280072);
nand I_33259 (I568301,I568284,I280060);
nor I_33260 (I568318,I568267,I568301);
DFFARX1 I_33261 (I568318,I2859,I568120,I568085,);
not I_33262 (I568349,I568301);
nand I_33263 (I568366,I568171,I568349);
nand I_33264 (I568097,I568233,I568349);
DFFARX1 I_33265 (I568267,I2859,I568120,I568112,);
not I_33266 (I568411,I280057);
nor I_33267 (I568428,I568411,I280072);
nor I_33268 (I568445,I568428,I568250);
DFFARX1 I_33269 (I568445,I2859,I568120,I568109,);
not I_33270 (I568476,I568428);
DFFARX1 I_33271 (I568476,I2859,I568120,I568502,);
not I_33272 (I568510,I568502);
nor I_33273 (I568106,I568510,I568428);
nor I_33274 (I568541,I568411,I280069);
and I_33275 (I568558,I568541,I280078);
or I_33276 (I568575,I568558,I280054);
DFFARX1 I_33277 (I568575,I2859,I568120,I568601,);
not I_33278 (I568609,I568601);
nand I_33279 (I568626,I568609,I568349);
not I_33280 (I568100,I568626);
nand I_33281 (I568094,I568626,I568366);
nand I_33282 (I568091,I568609,I568233);
not I_33283 (I568715,I2866);
DFFARX1 I_33284 (I145095,I2859,I568715,I568741,);
DFFARX1 I_33285 (I145089,I2859,I568715,I568758,);
not I_33286 (I568766,I568758);
nor I_33287 (I568683,I568741,I568766);
DFFARX1 I_33288 (I568766,I2859,I568715,I568698,);
nor I_33289 (I568811,I145077,I145098);
and I_33290 (I568828,I568811,I145092);
nor I_33291 (I568845,I568828,I145077);
not I_33292 (I568862,I145077);
and I_33293 (I568879,I568862,I145074);
nand I_33294 (I568896,I568879,I145086);
nor I_33295 (I568913,I568862,I568896);
DFFARX1 I_33296 (I568913,I2859,I568715,I568680,);
not I_33297 (I568944,I568896);
nand I_33298 (I568961,I568766,I568944);
nand I_33299 (I568692,I568828,I568944);
DFFARX1 I_33300 (I568862,I2859,I568715,I568707,);
not I_33301 (I569006,I145101);
nor I_33302 (I569023,I569006,I145074);
nor I_33303 (I569040,I569023,I568845);
DFFARX1 I_33304 (I569040,I2859,I568715,I568704,);
not I_33305 (I569071,I569023);
DFFARX1 I_33306 (I569071,I2859,I568715,I569097,);
not I_33307 (I569105,I569097);
nor I_33308 (I568701,I569105,I569023);
nor I_33309 (I569136,I569006,I145083);
and I_33310 (I569153,I569136,I145080);
or I_33311 (I569170,I569153,I145074);
DFFARX1 I_33312 (I569170,I2859,I568715,I569196,);
not I_33313 (I569204,I569196);
nand I_33314 (I569221,I569204,I568944);
not I_33315 (I568695,I569221);
nand I_33316 (I568689,I569221,I568961);
nand I_33317 (I568686,I569204,I568828);
not I_33318 (I569310,I2866);
DFFARX1 I_33319 (I116110,I2859,I569310,I569336,);
DFFARX1 I_33320 (I116104,I2859,I569310,I569353,);
not I_33321 (I569361,I569353);
nor I_33322 (I569278,I569336,I569361);
DFFARX1 I_33323 (I569361,I2859,I569310,I569293,);
nor I_33324 (I569406,I116092,I116113);
and I_33325 (I569423,I569406,I116107);
nor I_33326 (I569440,I569423,I116092);
not I_33327 (I569457,I116092);
and I_33328 (I569474,I569457,I116089);
nand I_33329 (I569491,I569474,I116101);
nor I_33330 (I569508,I569457,I569491);
DFFARX1 I_33331 (I569508,I2859,I569310,I569275,);
not I_33332 (I569539,I569491);
nand I_33333 (I569556,I569361,I569539);
nand I_33334 (I569287,I569423,I569539);
DFFARX1 I_33335 (I569457,I2859,I569310,I569302,);
not I_33336 (I569601,I116116);
nor I_33337 (I569618,I569601,I116089);
nor I_33338 (I569635,I569618,I569440);
DFFARX1 I_33339 (I569635,I2859,I569310,I569299,);
not I_33340 (I569666,I569618);
DFFARX1 I_33341 (I569666,I2859,I569310,I569692,);
not I_33342 (I569700,I569692);
nor I_33343 (I569296,I569700,I569618);
nor I_33344 (I569731,I569601,I116098);
and I_33345 (I569748,I569731,I116095);
or I_33346 (I569765,I569748,I116089);
DFFARX1 I_33347 (I569765,I2859,I569310,I569791,);
not I_33348 (I569799,I569791);
nand I_33349 (I569816,I569799,I569539);
not I_33350 (I569290,I569816);
nand I_33351 (I569284,I569816,I569556);
nand I_33352 (I569281,I569799,I569423);
not I_33353 (I569905,I2866);
DFFARX1 I_33354 (I268515,I2859,I569905,I569931,);
DFFARX1 I_33355 (I268497,I2859,I569905,I569948,);
not I_33356 (I569956,I569948);
nor I_33357 (I569873,I569931,I569956);
DFFARX1 I_33358 (I569956,I2859,I569905,I569888,);
nor I_33359 (I570001,I268503,I268506);
and I_33360 (I570018,I570001,I268494);
nor I_33361 (I570035,I570018,I268503);
not I_33362 (I570052,I268503);
and I_33363 (I570069,I570052,I268512);
nand I_33364 (I570086,I570069,I268500);
nor I_33365 (I570103,I570052,I570086);
DFFARX1 I_33366 (I570103,I2859,I569905,I569870,);
not I_33367 (I570134,I570086);
nand I_33368 (I570151,I569956,I570134);
nand I_33369 (I569882,I570018,I570134);
DFFARX1 I_33370 (I570052,I2859,I569905,I569897,);
not I_33371 (I570196,I268497);
nor I_33372 (I570213,I570196,I268512);
nor I_33373 (I570230,I570213,I570035);
DFFARX1 I_33374 (I570230,I2859,I569905,I569894,);
not I_33375 (I570261,I570213);
DFFARX1 I_33376 (I570261,I2859,I569905,I570287,);
not I_33377 (I570295,I570287);
nor I_33378 (I569891,I570295,I570213);
nor I_33379 (I570326,I570196,I268509);
and I_33380 (I570343,I570326,I268518);
or I_33381 (I570360,I570343,I268494);
DFFARX1 I_33382 (I570360,I2859,I569905,I570386,);
not I_33383 (I570394,I570386);
nand I_33384 (I570411,I570394,I570134);
not I_33385 (I569885,I570411);
nand I_33386 (I569879,I570411,I570151);
nand I_33387 (I569876,I570394,I570018);
endmodule


