module test_I15406(I12930,I1477,I1470,I12653,I15406);
input I12930,I1477,I1470,I12653;
output I15406;
wire I12619,I12670,I12602,I12584,I12783,I15047,I14982,I15389,I15064,I12596,I12587,I14965,I15372;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
not I_2(I12602,I12930);
and I_3(I12584,I12670,I12783);
DFFARX1 I_4(I1470,I12619,,,I12783,);
nor I_5(I15047,I14982,I12584);
not I_6(I14982,I12596);
not I_7(I15389,I15372);
nand I_8(I15064,I15047,I12587);
DFFARX1 I_9(I1470,I12619,,,I12596,);
nor I_10(I15406,I15064,I15389);
DFFARX1 I_11(I12670,I1470,I12619,,,I12587,);
not I_12(I14965,I1477);
DFFARX1 I_13(I12602,I1470,I14965,,,I15372,);
endmodule


