module test_I8896(I7122,I5085,I1477,I6975,I1470,I5642,I8896);
input I7122,I5085,I1477,I6975,I1470,I5642;
output I8896;
wire I7139,I6893,I5105,I7156,I6992,I6872,I5067,I6907,I7269,I5097,I7286;
or I_0(I7139,I7122,I5085);
nor I_1(I8896,I6893,I6872);
nand I_2(I6893,I7156,I7286);
not I_3(I5105,I1477);
DFFARX1 I_4(I7139,I1470,I6907,,,I7156,);
nand I_5(I6992,I6975,I5097);
DFFARX1 I_6(I7269,I1470,I6907,,,I6872,);
DFFARX1 I_7(I5642,I1470,I5105,,,I5067,);
not I_8(I6907,I1477);
DFFARX1 I_9(I5067,I1470,I6907,,,I7269,);
nand I_10(I5097,I5642);
nor I_11(I7286,I7269,I6992);
endmodule


