module test_I4068(I1447,I2929,I1477,I1263,I1470,I2861,I4068);
input I1447,I2929,I1477,I1263,I1470,I2861;
output I4068;
wire I2759,I2742,I3045,I3155,I2946,I3076,I2963,I3028,I2724;
not I_0(I2759,I1477);
or I_1(I2742,I3076,I2963);
and I_2(I3045,I2861,I3028);
or I_3(I3155,I3076,I3045);
or I_4(I2946,I2929,I1263);
DFFARX1 I_5(I1447,I1470,I2759,,,I3076,);
DFFARX1 I_6(I2946,I1470,I2759,,,I2963,);
nor I_7(I3028,I2963);
nor I_8(I4068,I2742,I2724);
DFFARX1 I_9(I3155,I1470,I2759,,,I2724,);
endmodule


