module test_I2072(I1518,I1215,I1423,I1207,I1295,I1470,I1455,I2072);
input I1518,I1215,I1423,I1207,I1295,I1470,I1455;
output I2072;
wire I2038,I2021,I1586,I1603,I1832,I1535,I2055;
not I_0(I2038,I2021);
and I_1(I2072,I1832,I2055);
DFFARX1 I_2(I1295,I1470,I1518,,,I2021,);
nor I_3(I1586,I1535,I1215);
nand I_4(I1603,I1586,I1423);
nand I_5(I1832,I1535,I1207);
not I_6(I1535,I1455);
nand I_7(I2055,I2038,I1603);
endmodule


