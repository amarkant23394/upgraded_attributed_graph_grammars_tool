module test_I6318(I3954,I1477,I1470,I3969,I6318);
input I3954,I1477,I1470,I3969;
output I6318;
wire I3963,I6346,I6329,I6380,I6363,I4181,I4034;
nor I_0(I3963,I4181,I4034);
nand I_1(I6346,I3969,I3954);
not I_2(I6329,I1477);
DFFARX1 I_3(I6363,I1470,I6329,,,I6380,);
and I_4(I6363,I6346,I3963);
not I_5(I6318,I6380);
DFFARX1 I_6(I1470,,,I4181,);
DFFARX1 I_7(I1470,,,I4034,);
endmodule


