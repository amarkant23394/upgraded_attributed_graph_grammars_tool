module test_I12687(I11167,I1477,I11057,I1470,I12687);
input I11167,I1477,I11057,I1470;
output I12687;
wire I12619,I12670,I10612,I10627,I10639,I12653,I12636;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
DFFARX1 I_2(I1470,,,I10612,);
not I_3(I12687,I12670);
nand I_4(I10627,I11167,I11057);
DFFARX1 I_5(I1470,,,I10639,);
and I_6(I12653,I12636,I10627);
nand I_7(I12636,I10612,I10639);
endmodule


