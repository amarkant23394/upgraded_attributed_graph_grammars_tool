module test_I16678(I14667,I1477,I13162,I14472,I1470,I16678);
input I14667,I1477,I13162,I14472,I1470;
output I16678;
wire I14338,I14856,I16339,I16644,I14605,I14356,I14537,I14808,I14370,I16356,I14347,I16240,I14353,I14777,I16661;
DFFARX1 I_0(I14605,I1470,I14370,,,I14338,);
nor I_1(I14856,I14808);
nor I_2(I16339,I14353,I14338);
DFFARX1 I_3(I14347,I1470,I16240,,,I16644,);
and I_4(I14605,I14537,I14472);
nand I_5(I14356,I14667,I14856);
DFFARX1 I_6(I1470,I14370,,,I14537,);
DFFARX1 I_7(I13162,I1470,I14370,,,I14808,);
not I_8(I14370,I1477);
DFFARX1 I_9(I14356,I1470,I16240,,,I16356,);
DFFARX1 I_10(I14777,I1470,I14370,,,I14347,);
not I_11(I16240,I1477);
not I_12(I14353,I14808);
or I_13(I14777,I14667);
nand I_14(I16661,I16644,I16356);
and I_15(I16678,I16339,I16661);
endmodule


