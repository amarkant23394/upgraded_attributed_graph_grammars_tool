module test_final(G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8,n_431_0_l_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_8,blif_clk_net_1_r_7,n8_7,G42_1_r_8,);
nor I_1(n_572_1_r_8,n39_8,n23_8);
and I_2(n_549_1_r_8,n38_8,n23_8);
nand I_3(n_569_1_r_8,n38_8,n24_8);
nor I_4(n_452_1_r_8,n25_8,n26_8);
nor I_5(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_6(N3_2_r_8,blif_clk_net_1_r_7,n8_7,G199_2_r_8,);
DFFARX1 I_7(N1_4_r_8,blif_clk_net_1_r_7,n8_7,G199_4_r_8,);
DFFARX1 I_8(G78_0_l_8,blif_clk_net_1_r_7,n8_7,G214_4_r_8,);
or I_9(n_431_0_l_8,IN_8_0_l_8,n29_8);
DFFARX1 I_10(n_431_0_l_8,blif_clk_net_1_r_7,n8_7,G78_0_l_8,);
not I_11(n19_8,G78_0_l_8);
DFFARX1 I_12(IN_2_5_l_8,blif_clk_net_1_r_7,n8_7,n39_8,);
not I_13(n22_8,n39_8);
DFFARX1 I_14(IN_1_5_l_8,blif_clk_net_1_r_7,n8_7,n38_8,);
nor I_15(n4_1_r_8,G78_0_l_8,n33_8);
nor I_16(N3_2_r_8,n22_8,n35_8);
nor I_17(N1_4_r_8,n27_8,n37_8);
nand I_18(n23_8,IN_7_0_l_8,n32_8);
not I_19(n24_8,n23_8);
nand I_20(n25_8,IN_11_0_l_8,n36_8);
nand I_21(n26_8,n27_8,n28_8);
nor I_22(n27_8,IN_5_0_l_8,n31_8);
not I_23(n28_8,G2_0_l_8);
and I_24(n29_8,IN_2_0_l_8,n30_8);
nor I_25(n30_8,IN_4_0_l_8,n31_8);
not I_26(n31_8,G1_0_l_8);
and I_27(n32_8,IN_5_0_l_8,n28_8);
nand I_28(n33_8,n28_8,n34_8);
not I_29(n34_8,n25_8);
nor I_30(n35_8,G2_0_l_8,n34_8);
not I_31(n36_8,IN_10_0_l_8);
nor I_32(n37_8,n19_8,n38_8);
DFFARX1 I_33(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_34(n_572_1_r_7,n30_7,n31_7);
nand I_35(n_573_1_r_7,n28_7,G42_1_r_8);
nor I_36(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_37(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_38(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_39(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_40(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_41(P6_5_r_7,P6_5_r_internal_7);
or I_42(n_431_0_l_7,n36_7,n_572_1_r_8);
not I_43(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_44(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_45(n27_7,n43_7);
DFFARX1 I_46(n_572_1_r_8,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_47(n_42_2_r_8,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_48(n4_1_r_7,n30_7,n38_7);
nor I_49(N1_4_r_7,n27_7,n40_7);
nand I_50(n26_7,n39_7,G214_4_r_8);
not I_51(n5_7,n_569_1_r_8);
DFFARX1 I_52(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_53(n28_7,n26_7,n29_7);
not I_54(n29_7,G199_2_r_8);
not I_55(n30_7,G42_1_r_8);
nand I_56(n31_7,n27_7,n29_7);
nor I_57(n32_7,ACVQN1_5_l_7,n34_7);
nor I_58(n33_7,n29_7,n_569_1_r_8);
not I_59(n34_7,G42_1_r_8);
nor I_60(n35_7,n43_7,n44_7);
and I_61(n36_7,n37_7,n_549_1_r_8);
nor I_62(n37_7,n30_7,n_452_1_r_8);
nand I_63(n38_7,n29_7,n_569_1_r_8);
nor I_64(n39_7,n_569_1_r_8,G199_4_r_8);
nor I_65(n40_7,n44_7,n41_7);
nor I_66(n41_7,n34_7,n42_7);
nand I_67(n42_7,n5_7,G199_2_r_8);
endmodule


