module test_I11378(I9320,I9179,I6887,I8896,I8981,I6884,I6992,I7057,I6878,I11378);
input I9320,I9179,I6887,I8896,I8981,I6884,I6992,I7057,I6878;
output I11378;
wire I8830,I8913,I8930,I9396,I6881,I8848,I9083,I9413,I8947,I9227,I8879,I11327;
nand I_0(I8830,I8913,I9227);
nand I_1(I8913,I8896,I6878);
nor I_2(I8930,I8879);
not I_3(I9396,I9320);
nand I_4(I6881,I6992,I7057);
nor I_5(I8848,I9083,I9413);
nand I_6(I9083,I8879,I6881);
and I_7(I9413,I8947,I9396);
nand I_8(I8947,I8930,I6884);
nor I_9(I11378,I11327,I8848);
nor I_10(I9227,I9179,I8981);
not I_11(I8879,I6887);
not I_12(I11327,I8830);
endmodule


