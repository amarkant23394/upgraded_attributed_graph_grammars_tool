module test_I15832(I12270,I1477,I1470,I11944,I15832);
input I12270,I1477,I1470,I11944;
output I15832;
wire I13908,I13743,I12239,I14162,I11938,I15628,I13749,I13891,I13775;
not I_0(I13908,I13891);
DFFARX1 I_1(I13891,I1470,I13775,,,I13743,);
DFFARX1 I_2(I1470,,,I12239,);
nand I_3(I15832,I15628,I13749);
DFFARX1 I_4(I11938,I1470,I13775,,,I14162,);
and I_5(I11938,I12270,I12239);
not I_6(I15628,I13743);
nand I_7(I13749,I14162,I13908);
DFFARX1 I_8(I11944,I1470,I13775,,,I13891,);
not I_9(I13775,I1477);
endmodule


