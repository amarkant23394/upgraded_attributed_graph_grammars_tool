module test_I8479(I1477,I5785,I8411,I6265,I1470,I8479);
input I1477,I5785,I8411,I6265,I1470;
output I8479;
wire I8428,I5802,I5833,I5728,I8216,I8298,I5719,I8315,I5751,I8445,I5734,I8462,I8233,I5740,I5722;
and I_0(I8428,I8411,I5734);
DFFARX1 I_1(I5785,I1470,I5751,,,I5802,);
DFFARX1 I_2(I5802,I1470,I5751,,,I5833,);
not I_3(I5728,I5833);
not I_4(I8216,I1477);
nor I_5(I8298,I8233,I5719);
DFFARX1 I_6(I6265,I1470,I5751,,,I5719,);
nand I_7(I8315,I8298,I5740);
not I_8(I5751,I1477);
or I_9(I8445,I8428,I5728);
DFFARX1 I_10(I1470,I5751,,,I5734,);
DFFARX1 I_11(I8445,I1470,I8216,,,I8462,);
nor I_12(I8479,I8462,I8315);
not I_13(I8233,I5722);
not I_14(I5740,I5802);
DFFARX1 I_15(I1470,I5751,,,I5722,);
endmodule


