module test_I12007(I10253,I7550,I1477,I1470,I10202,I10120,I12007);
input I10253,I7550,I1477,I1470,I10202,I10120;
output I12007;
wire I10349,I10270,I10029,I10219,I10154,I10020,I10137,I10052,I10287,I10332,I10459;
and I_0(I10349,I10332,I7550);
and I_1(I10270,I10120,I10253);
DFFARX1 I_2(I10459,I1470,I10052,,,I10029,);
DFFARX1 I_3(I10202,I1470,I10052,,,I10219,);
nand I_4(I10154,I10137,I10120);
nor I_5(I12007,I10020,I10029);
DFFARX1 I_6(I10287,I1470,I10052,,,I10020,);
DFFARX1 I_7(I1470,I10052,,,I10137,);
not I_8(I10052,I1477);
and I_9(I10287,I10219,I10154);
DFFARX1 I_10(I1470,I10052,,,I10332,);
or I_11(I10459,I10349,I10270);
endmodule


