module test_I4512(I1477,I1303,I1470,I4725,I4512);
input I1477,I1303,I1470,I4725;
output I4512;
wire I2540,I2143,I2181,I4544,I2170,I2557,I2232,I4674,I2155,I4742,I4807,I4824,I4790,I2633,I4773;
DFFARX1 I_0(I1470,I2181,,,I2540,);
DFFARX1 I_1(I2557,I1470,I2181,,,I2143,);
not I_2(I2181,I1477);
not I_3(I4544,I1477);
not I_4(I2170,I2232);
and I_5(I2557,I2540,I1303);
nand I_6(I4512,I4824,I4790);
DFFARX1 I_7(I1470,I2181,,,I2232,);
DFFARX1 I_8(I2155,I1470,I4544,,,I4674,);
DFFARX1 I_9(I2633,I1470,I2181,,,I2155,);
DFFARX1 I_10(I4725,I1470,I4544,,,I4742,);
DFFARX1 I_11(I2170,I1470,I4544,,,I4807,);
and I_12(I4824,I4807,I2143);
nor I_13(I4790,I4674,I4773);
DFFARX1 I_14(I1470,I2181,,,I2633,);
not I_15(I4773,I4742);
endmodule


