module test_I14227(I1477,I1470,I11990,I14227);
input I1477,I1470,I11990;
output I14227;
wire I12270,I12239,I14162,I11938,I10014,I12208,I13775,I11973;
nand I_0(I12270,I11990,I10014);
DFFARX1 I_1(I12208,I1470,I11973,,,I12239,);
DFFARX1 I_2(I11938,I1470,I13775,,,I14162,);
not I_3(I14227,I14162);
and I_4(I11938,I12270,I12239);
DFFARX1 I_5(I1470,,,I10014,);
DFFARX1 I_6(I1470,I11973,,,I12208,);
not I_7(I13775,I1477);
not I_8(I11973,I1477);
endmodule


