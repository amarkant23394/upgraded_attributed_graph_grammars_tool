module test_I3374(I1477,I1637,I1586,I1383,I1423,I1470,I3374);
input I1477,I1637,I1586,I1383,I1423,I1470;
output I3374;
wire I1486,I3470,I3747,I1897,I1483,I3388,I1492,I1767,I1518,I1668,I1504,I3620,I1880,I1603,I3877,I3453,I1501;
DFFARX1 I_0(I1470,I1518,,,I1486,);
not I_1(I3470,I3453);
DFFARX1 I_2(I1504,I1470,I3388,,,I3747,);
nor I_3(I1897,I1880,I1603);
DFFARX1 I_4(I1880,I1470,I1518,,,I1483,);
not I_5(I3388,I1477);
nand I_6(I1492,I1603,I1668);
DFFARX1 I_7(I1470,I1518,,,I1767,);
not I_8(I1518,I1477);
not I_9(I1668,I1637);
nand I_10(I1504,I1767,I1897);
nor I_11(I3620,I1492,I1483);
DFFARX1 I_12(I1383,I1470,I1518,,,I1880,);
nand I_13(I1603,I1586,I1423);
nor I_14(I3877,I3747,I3470);
nor I_15(I3453,I1486,I1501);
nand I_16(I3374,I3620,I3877);
not I_17(I1501,I1880);
endmodule


