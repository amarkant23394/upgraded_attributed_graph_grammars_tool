module test_I4536(I2173,I1477,I1470,I2678,I2311,I4536);
input I2173,I1477,I1470,I2678,I2311;
output I4536;
wire I2181,I4595,I4544,I4869,I2149,I4561,I2152,I2345,I4578,I2161,I2695;
not I_0(I2181,I1477);
nor I_1(I4536,I4869,I4595);
DFFARX1 I_2(I4578,I1470,I4544,,,I4595,);
not I_3(I4544,I1477);
DFFARX1 I_4(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_5(I2695,I1470,I2181,,,I2149,);
nand I_6(I4561,I2152,I2173);
DFFARX1 I_7(I1470,I2181,,,I2152,);
DFFARX1 I_8(I1470,I2181,,,I2345,);
and I_9(I4578,I4561,I2161);
nand I_10(I2161,I2345,I2311);
and I_11(I2695,I2345,I2678);
endmodule


