module test_I2039(I1322,I1294,I1492,I1301,I1639,I2039);
input I1322,I1294,I1492,I1301,I1639;
output I2039;
wire I1316,I1687,I2005,I1937,I2022,I1342,I1509,I1954,I1310,I1577;
nand I_0(I1316,I1509,I1687);
not I_1(I1687,I1639);
nor I_2(I2005,I1954,I1310);
not I_3(I1937,I1301);
nand I_4(I2022,I2005,I1316);
DFFARX1 I_5(I2022,I1294,I1937,,,I2039,);
not I_6(I1342,I1301);
DFFARX1 I_7(I1492,I1294,I1342,,,I1509,);
not I_8(I1954,I1322);
DFFARX1 I_9(I1577,I1294,I1342,,,I1310,);
and I_10(I1577,I1509);
endmodule


