module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_11,blif_reset_net_1_r_11,G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_11,blif_reset_net_1_r_11;
output G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,n_431_0_l_11,n9_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_11,n9_11,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_11,n9_11,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_11,n9_11,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_11,n9_11,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_11,n9_11,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_11,n9_11,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_11,n9_11,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_11,n9_11,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_11,n9_11,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_11,blif_clk_net_1_r_11,n9_11,G42_1_r_11,);
nor I_31(n_572_1_r_11,n29_11,n30_11);
nand I_32(n_573_1_r_11,n26_11,n28_11);
nor I_33(n_549_1_r_11,n27_11,n32_11);
nand I_34(n_569_1_r_11,n45_11,n28_11);
nor I_35(n_452_1_r_11,n43_11,n44_11);
nor I_36(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_37(N3_2_r_11,blif_clk_net_1_r_11,n9_11,G199_2_r_11,);
DFFARX1 I_38(n24_11,blif_clk_net_1_r_11,n9_11,ACVQN2_3_r_11,);
nor I_39(n_266_and_0_3_r_11,n20_11,n37_11);
or I_40(n_431_0_l_11,n33_11,G42_1_r_10);
not I_41(n9_11,blif_reset_net_1_r_11);
DFFARX1 I_42(n_431_0_l_11,blif_clk_net_1_r_11,n9_11,n43_11,);
not I_43(n26_11,n43_11);
DFFARX1 I_44(n_573_1_r_10,blif_clk_net_1_r_11,n9_11,n44_11,);
DFFARX1 I_45(n_572_1_r_10,blif_clk_net_1_r_11,n9_11,n45_11,);
not I_46(n27_11,n45_11);
nor I_47(n4_1_r_11,n44_11,n25_11);
nor I_48(N3_2_r_11,n45_11,n40_11);
nand I_49(n24_11,n39_11,n_572_1_r_10);
nand I_50(n25_11,n38_11,G42_1_r_10);
DFFARX1 I_51(n25_11,blif_clk_net_1_r_11,n9_11,n20_internal_11,);
not I_52(n20_11,n20_internal_11);
not I_53(n28_11,n25_11);
not I_54(n29_11,n_549_1_r_10);
nand I_55(n30_11,n26_11,n31_11);
not I_56(n31_11,ACVQN2_3_r_10);
and I_57(n32_11,n26_11,n44_11);
and I_58(n33_11,n34_11,n_266_and_0_3_r_10);
nor I_59(n34_11,n29_11,G199_2_r_10);
not I_60(n35_11,n_42_2_r_10);
nand I_61(n36_11,n31_11,n_549_1_r_10);
nor I_62(n37_11,n29_11,ACVQN2_3_r_10);
nor I_63(n38_11,n31_11,n_42_2_r_10);
nor I_64(n39_11,n_42_2_r_10,n_573_1_r_10);
nor I_65(n40_11,n41_11,n_42_2_r_10);
nor I_66(n41_11,n42_11,n_573_1_r_10);
not I_67(n42_11,n_572_1_r_10);
endmodule


