module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_7_r_4,n6_4,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_7_r_4,n6_4,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N1371_0_r_4,n25_4,N1372_1_r_16);
not I_41(N1508_0_r_4,n25_4);
nor I_42(N1507_6_r_4,n32_4,n33_4);
nor I_43(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_44(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_45(n_572_7_r_4,n_573_7_r_4);
nand I_46(n_573_7_r_4,n21_4,n22_4);
nor I_47(n_549_7_r_4,n24_4,N1372_1_r_16);
nand I_48(n_569_7_r_4,n22_4,n23_4);
nor I_49(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_50(N6147_9_r_4,n28_4);
nor I_51(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_52(I_BUFF_1_9_r_4,n21_4);
nor I_53(n4_7_r_4,N6147_9_r_4,N1372_1_r_16);
not I_54(n6_4,blif_reset_net_7_r_4);
nand I_55(n21_4,n39_4,n40_4);
or I_56(n22_4,n31_4,G42_7_r_16);
not I_57(n23_4,N1372_1_r_16);
nor I_58(n24_4,n25_4,n26_4);
nand I_59(n25_4,N1508_6_r_16,n_569_7_r_16);
nand I_60(n26_4,n21_4,n27_4);
nand I_61(n27_4,n36_4,n37_4);
nand I_62(n28_4,n38_4,n_573_7_r_16);
nand I_63(n29_4,N1508_0_r_4,n30_4);
nand I_64(n30_4,n34_4,n35_4);
nor I_65(n31_4,N1371_0_r_16,N6147_2_r_16);
not I_66(n32_4,n30_4);
nor I_67(n33_4,n21_4,n28_4);
nand I_68(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_69(n35_4,N1508_0_r_4,n27_4);
not I_70(n36_4,N1507_6_r_16);
nand I_71(n37_4,n_452_7_r_16,N1371_0_r_16);
or I_72(n38_4,N1371_0_r_16,N6147_2_r_16);
nor I_73(n39_4,N1508_1_r_16,N1508_0_r_16);
or I_74(n40_4,n41_4,N1372_1_r_16);
nor I_75(n41_4,N1508_0_r_16,n_572_7_r_16);
endmodule


