module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_5_r_11,n9_11,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
not I_34(N1372_1_r_11,n53_11);
nor I_35(N1508_1_r_11,n39_11,n53_11);
nor I_36(N6147_2_r_11,n48_11,n49_11);
nor I_37(N6147_3_r_11,n44_11,n45_11);
nand I_38(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_39(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_40(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_41(n_102_5_r_11,n39_11);
nand I_42(n_547_5_r_11,n36_11,n37_11);
nor I_43(N1507_6_r_11,n52_11,n57_11);
nor I_44(N1508_6_r_11,n46_11,n51_11);
nor I_45(N1372_10_r_11,n43_11,n47_11);
nor I_46(N1508_10_r_11,n55_11,n56_11);
nand I_47(n_431_5_r_11,n40_11,n41_11);
not I_48(n9_11,blif_reset_net_5_r_11);
nor I_49(n36_11,n38_11,n39_11);
not I_50(n37_11,n40_11);
nor I_51(n38_11,n60_11,G42_7_r_12);
nor I_52(n39_11,n54_11,n_572_7_r_12);
nand I_53(n40_11,G42_7_r_12,N1507_6_r_12);
nand I_54(n41_11,n_102_5_r_11,n42_11);
and I_55(n42_11,n58_11,N1507_6_r_12);
not I_56(n43_11,n44_11);
nor I_57(n44_11,n40_11,N1371_0_r_12);
nand I_58(n45_11,n46_11,n47_11);
not I_59(n46_11,n38_11);
nand I_60(n47_11,n59_11,n62_11);
and I_61(n48_11,n37_11,n47_11);
or I_62(n49_11,n44_11,n50_11);
nor I_63(n50_11,n60_11,n61_11);
or I_64(n51_11,n_102_5_r_11,n52_11);
nor I_65(n52_11,n42_11,n57_11);
nand I_66(n53_11,n37_11,n50_11);
or I_67(n54_11,N1371_0_r_12,N1508_0_r_12);
nor I_68(n55_11,n38_11,n42_11);
not I_69(n56_11,N1372_10_r_11);
and I_70(n57_11,n38_11,n50_11);
and I_71(n58_11,n59_11,N1508_0_r_12);
or I_72(n59_11,n63_11,N1508_6_r_12);
not I_73(n60_11,n_569_7_r_12);
nor I_74(n61_11,n_572_7_r_12,n_549_7_r_12);
nand I_75(n62_11,N1508_6_r_12,N6147_9_r_12);
and I_76(n63_11,N1508_6_r_12,N6147_9_r_12);
endmodule


