module test_I11768(I9320,I1477,I6881,I8947,I1470,I8879,I11768);
input I9320,I1477,I6881,I8947,I1470,I8879;
output I11768;
wire I8845,I8836,I9179,I8839,I11344,I9396,I9210,I8848,I9083,I9413,I11672,I11361,I11429,I9066,I11310,I11751;
or I_0(I8845,I9179,I9066);
nand I_1(I8836,I9320,I9210);
and I_2(I11768,I11429,I11751);
DFFARX1 I_3(I1470,,,I9179,);
DFFARX1 I_4(I1470,,,I8839,);
nor I_5(I11344,I8848,I8839);
not I_6(I9396,I9320);
nor I_7(I9210,I9179,I8947);
nor I_8(I8848,I9083,I9413);
nand I_9(I9083,I8879,I6881);
and I_10(I9413,I8947,I9396);
DFFARX1 I_11(I8836,I1470,I11310,,,I11672,);
nand I_12(I11361,I11344,I8845);
not I_13(I11429,I8848);
DFFARX1 I_14(I1470,,,I9066,);
not I_15(I11310,I1477);
nand I_16(I11751,I11672,I11361);
endmodule


