module test_I3447(I1911,I2022,I1294,I2344,I2702,I1301,I3447);
input I1911,I2022,I1294,I2344,I2702,I1301;
output I3447;
wire I2668,I2733,I1914,I2583,I3413,I2945,I2897,I2600,I2551,I2651,I2557,I1923,I3430,I2566;
nand I_0(I2668,I2651,I1914);
not I_1(I2733,I2702);
DFFARX1 I_2(I1294,,,I1914,);
not I_3(I2583,I1301);
not I_4(I3413,I2566);
DFFARX1 I_5(I1294,I2583,,,I2945,);
nand I_6(I2897,I2600,I1923);
not I_7(I2600,I1911);
and I_8(I3447,I3430,I2551);
DFFARX1 I_9(I2897,I1294,I2583,,,I2551,);
nor I_10(I2651,I2600);
nand I_11(I2557,I2668,I2733);
nand I_12(I1923,I2022,I2344);
nor I_13(I3430,I3413,I2557);
not I_14(I2566,I2945);
endmodule


