module test_I1359(I1263,I1359);
input I1263;
output I1359;
wire ;
not I_0(I1359,I1263);
endmodule


