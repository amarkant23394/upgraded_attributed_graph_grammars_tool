module test_I3951(I1477,I2980,I4164,I1470,I2844,I3951);
input I1477,I2980,I4164,I1470,I2844;
output I3951;
wire I2733,I3107,I3076,I2751,I3983,I3200,I4263,I3310,I4229,I2745,I3217,I4113,I4181,I4212,I4246;
nand I_0(I2733,I3217,I3107);
nor I_1(I3107,I3076,I2844);
DFFARX1 I_2(I1470,,,I3076,);
nor I_3(I2751,I3076,I3217);
not I_4(I3983,I1477);
DFFARX1 I_5(I1470,,,I3200,);
and I_6(I4263,I4246,I2733);
and I_7(I3310,I2844);
nor I_8(I4229,I4113,I4212);
nor I_9(I2745,I2980,I3310);
nand I_10(I3951,I4263,I4229);
not I_11(I3217,I3200);
DFFARX1 I_12(I2751,I1470,I3983,,,I4113,);
DFFARX1 I_13(I4164,I1470,I3983,,,I4181,);
not I_14(I4212,I4181);
DFFARX1 I_15(I2745,I1470,I3983,,,I4246,);
endmodule


