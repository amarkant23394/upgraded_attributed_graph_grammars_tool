module test_I11990(I10349,I10086,I1477,I1470,I8124,I11990);
input I10349,I10086,I1477,I1470,I8124;
output I11990;
wire I10032,I7570,I10414,I10397,I10137,I7553,I10052,I10103;
nand I_0(I10032,I10137,I10414);
not I_1(I7570,I1477);
nor I_2(I10414,I10103,I10397);
not I_3(I10397,I10349);
DFFARX1 I_4(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_5(I8124,I1470,I7570,,,I7553,);
not I_6(I11990,I10032);
not I_7(I10052,I1477);
DFFARX1 I_8(I10086,I1470,I10052,,,I10103,);
endmodule


