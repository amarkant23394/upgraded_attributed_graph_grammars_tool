module test_I14114(I12270,I1477,I10041,I1470,I14114);
input I12270,I1477,I10041,I1470;
output I14114;
wire I11935,I11956,I11950,I14004,I12349,I12208,I14049,I13987,I13775,I11973,I13970,I11962,I14066,I11941;
DFFARX1 I_0(I12208,I1470,I11973,,,I11935,);
not I_1(I11956,I12349);
DFFARX1 I_2(I1470,I11973,,,I11950,);
DFFARX1 I_3(I13987,I1470,I13775,,,I14004,);
nand I_4(I14114,I14066,I14004);
DFFARX1 I_5(I10041,I1470,I11973,,,I12349,);
DFFARX1 I_6(I1470,I11973,,,I12208,);
DFFARX1 I_7(I11962,I1470,I13775,,,I14049,);
and I_8(I13987,I13970,I11941);
not I_9(I13775,I1477);
not I_10(I11973,I1477);
nand I_11(I13970,I11935,I11950);
nor I_12(I11962,I12349,I12270);
and I_13(I14066,I14049,I11956);
DFFARX1 I_14(I12208,I1470,I11973,,,I11941,);
endmodule


