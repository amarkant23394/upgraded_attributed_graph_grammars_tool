module test_I1923(I1797,I1322,I1294,I1492,I1639,I1410,I1301,I1923);
input I1797,I1322,I1294,I1492,I1639,I1410,I1301;
output I1923;
wire I2005,I2313,I2022,I1316,I1971,I1334,I1310,I1577,I1319,I2344,I1331,I1954,I1687,I1937,I1342,I1988,I1509;
nor I_0(I2005,I1954,I1310);
DFFARX1 I_1(I1331,I1294,I1937,,,I2313,);
nand I_2(I2022,I2005,I1316);
nand I_3(I1316,I1509,I1687);
nor I_4(I1971,I1310,I1319);
DFFARX1 I_5(I1797,I1294,I1342,,,I1334,);
DFFARX1 I_6(I1577,I1294,I1342,,,I1310,);
and I_7(I1577,I1509);
DFFARX1 I_8(I1294,I1342,,,I1319,);
nor I_9(I2344,I2313,I1988);
nor I_10(I1331,I1639,I1410);
not I_11(I1954,I1322);
not I_12(I1687,I1639);
not I_13(I1937,I1301);
not I_14(I1342,I1301);
nand I_15(I1923,I2022,I2344);
nand I_16(I1988,I1971,I1334);
DFFARX1 I_17(I1492,I1294,I1342,,,I1509,);
endmodule


