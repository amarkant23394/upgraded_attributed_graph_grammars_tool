module test_I11938(I1477,I10414,I12174,I1470,I10202,I11938);
input I1477,I10414,I12174,I1470,I10202;
output I11938;
wire I12270,I10032,I10219,I12239,I10014,I12208,I10023,I11990,I10137,I11973,I10052,I12191;
nand I_0(I12270,I11990,I10014);
nand I_1(I10032,I10137,I10414);
DFFARX1 I_2(I10202,I1470,I10052,,,I10219,);
DFFARX1 I_3(I12208,I1470,I11973,,,I12239,);
DFFARX1 I_4(I10219,I1470,I10052,,,I10014,);
DFFARX1 I_5(I12191,I1470,I11973,,,I12208,);
and I_6(I11938,I12270,I12239);
DFFARX1 I_7(I10137,I1470,I10052,,,I10023,);
not I_8(I11990,I10032);
DFFARX1 I_9(I1470,I10052,,,I10137,);
not I_10(I11973,I1477);
not I_11(I10052,I1477);
or I_12(I12191,I12174,I10023);
endmodule


