module test_I2866(I2781,I1294,I2505,I2406,I1301,I2866);
input I2781,I1294,I2505,I2406,I1301;
output I2866;
wire I2815,I2798,I1917,I2583,I1899,I2832;
or I_0(I2815,I2798,I1917);
and I_1(I2798,I2781,I1899);
nand I_2(I1917,I2406,I2505);
DFFARX1 I_3(I2832,I1294,I2583,,,I2866,);
not I_4(I2583,I1301);
DFFARX1 I_5(I1294,,,I1899,);
DFFARX1 I_6(I2815,I1294,I2583,,,I2832,);
endmodule


