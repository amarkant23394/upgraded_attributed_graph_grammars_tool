module test_I4996(I1477,I2311,I1239,I1303,I4708,I1470,I2158,I4996);
input I1477,I2311,I1239,I1303,I4708,I1470,I2158;
output I4996;
wire I2167,I4979,I4629,I2328,I4544,I4869,I2149,I4962,I2633,I2540,I2458,I2173,I2181,I2509,I2557,I2232,I4742,I4725;
nand I_0(I2167,I2633,I2328);
nor I_1(I4979,I4742,I4962);
nor I_2(I4629,I2167,I2173);
nor I_3(I2328,I2232,I2311);
not I_4(I4544,I1477);
DFFARX1 I_5(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_6(I1470,I2181,,,I2149,);
not I_7(I4962,I4869);
DFFARX1 I_8(I1239,I1470,I2181,,,I2633,);
DFFARX1 I_9(I1470,I2181,,,I2540,);
DFFARX1 I_10(I1470,I2181,,,I2458,);
nand I_11(I2173,I2557,I2509);
not I_12(I2181,I1477);
nor I_13(I2509,I2458,I2232);
and I_14(I2557,I2540,I1303);
DFFARX1 I_15(I1470,I2181,,,I2232,);
DFFARX1 I_16(I4725,I1470,I4544,,,I4742,);
and I_17(I4725,I4708,I2158);
and I_18(I4996,I4629,I4979);
endmodule


