module test_I3702(I1637,I1477,I1603,I1470,I3702);
input I1637,I1477,I1603,I1470;
output I3702;
wire I3388,I1928,I1668,I3668,I2038,I1507,I2021,I1880,I1498,I3685;
not I_0(I3388,I1477);
DFFARX1 I_1(I3685,I1470,I3388,,,I3702,);
nor I_2(I1928,I1880,I1668);
not I_3(I1668,I1637);
DFFARX1 I_4(I1507,I1470,I3388,,,I3668,);
not I_5(I2038,I2021);
nor I_6(I1507,I1603,I1637);
DFFARX1 I_7(I1470,,,I2021,);
DFFARX1 I_8(I1470,,,I1880,);
nand I_9(I1498,I2038,I1928);
and I_10(I3685,I3668,I1498);
endmodule


