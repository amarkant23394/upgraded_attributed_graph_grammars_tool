module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_8_r_10,n11_10,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N1371_0_r_10,n37_10,n38_10);
nor I_37(N1508_0_r_10,n37_10,n58_10);
nand I_38(N6147_2_r_10,n39_10,n40_10);
not I_39(N6147_3_r_10,n39_10);
nor I_40(N1372_4_r_10,n46_10,n49_10);
nor I_41(N1508_4_r_10,n51_10,n52_10);
nor I_42(N1507_6_r_10,n49_10,n60_10);
nor I_43(N1508_6_r_10,n49_10,n50_10);
nor I_44(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_45(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_46(N6147_9_r_10,n36_10,n37_10);
nor I_47(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_48(I_BUFF_1_9_r_10,n48_10);
nor I_49(N3_8_r_10,n44_10,n47_10);
not I_50(n11_10,blif_reset_net_8_r_10);
not I_51(n35_10,n49_10);
nor I_52(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_53(n37_10,N1507_6_r_5);
not I_54(n38_10,n46_10);
nand I_55(n39_10,n43_10,n44_10);
nand I_56(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_57(n41_10,n42_10,N1507_6_r_5);
not I_58(n42_10,n44_10);
nor I_59(n43_10,n45_10,N1507_6_r_5);
nand I_60(n44_10,n54_10,N1508_0_r_5);
nor I_61(n45_10,n59_10,N1508_0_r_5);
nand I_62(n46_10,n61_10,N1371_0_r_5);
nor I_63(n47_10,n46_10,n48_10);
nand I_64(n48_10,n62_10,n63_10);
nand I_65(n49_10,n56_10,n_452_7_r_5);
not I_66(n50_10,n45_10);
nor I_67(n51_10,n42_10,n53_10);
not I_68(n52_10,N1372_4_r_10);
nor I_69(n53_10,n48_10,n50_10);
and I_70(n54_10,n55_10,N6147_2_r_5);
nand I_71(n55_10,n56_10,n57_10);
nand I_72(n56_10,N1508_1_r_5,N1371_0_r_5);
not I_73(n57_10,n_452_7_r_5);
nor I_74(n58_10,n35_10,n45_10);
nor I_75(n59_10,N1508_6_r_5,G42_7_r_5);
nor I_76(n60_10,n37_10,n46_10);
or I_77(n61_10,N1508_6_r_5,G42_7_r_5);
nor I_78(n62_10,N1372_1_r_5,N1508_1_r_5);
or I_79(n63_10,n64_10,n_572_7_r_5);
nor I_80(n64_10,n_573_7_r_5,n_569_7_r_5);
endmodule


