module test_I9474(I8527,I1477,I5737,I1470,I9474);
input I8527,I1477,I5737,I1470;
output I9474;
wire I8202,I8496,I9525,I9508,I9542,I8216,I8561,I5719,I8377,I8250,I9491,I8181,I8360,I8592,I8184,I8462,I9576,I8267,I8199;
nand I_0(I8202,I8267,I8496);
nor I_1(I8496,I8462,I8377);
or I_2(I9474,I9576,I9542);
and I_3(I9525,I9508,I8184);
nand I_4(I9508,I8199,I8202);
DFFARX1 I_5(I9525,I1470,I9491,,,I9542,);
not I_6(I8216,I1477);
and I_7(I8561,I8527);
DFFARX1 I_8(I1470,,,I5719,);
not I_9(I8377,I8360);
nor I_10(I8250,I5719);
not I_11(I9491,I1477);
and I_12(I8181,I8360,I8592);
not I_13(I8360,I5719);
DFFARX1 I_14(I8527,I1470,I8216,,,I8592,);
DFFARX1 I_15(I8561,I1470,I8216,,,I8184,);
DFFARX1 I_16(I1470,I8216,,,I8462,);
nor I_17(I9576,I8181,I8202);
nand I_18(I8267,I8250,I5737);
DFFARX1 I_19(I1470,I8216,,,I8199,);
endmodule


