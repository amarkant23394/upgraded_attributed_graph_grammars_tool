module test_I2557(I2440,I1911,I2234,I1294,I1301,I2557);
input I2440,I1911,I2234,I1294,I1301;
output I2557;
wire I2668,I2733,I2600,I1914,I2651,I1937,I2039,I1908,I2457,I2702;
nand I_0(I2668,I2651,I1914);
not I_1(I2733,I2702);
not I_2(I2600,I1911);
DFFARX1 I_3(I2457,I1294,I1937,,,I1914,);
nand I_4(I2557,I2668,I2733);
nor I_5(I2651,I2600,I1908);
not I_6(I1937,I1301);
DFFARX1 I_7(I1294,I1937,,,I2039,);
not I_8(I1908,I2039);
or I_9(I2457,I2234,I2440);
not I_10(I2702,I1908);
endmodule


