module test_final(G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_6,blif_reset_net_1_r_6,G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6);
input G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_6,blif_reset_net_1_r_6;
output G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6;
wire G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4,n_431_0_l_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,N3_2_l_6,n4_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6;
DFFARX1 I_0(n4_1_r_4,blif_clk_net_1_r_6,n4_6,G42_1_r_4,);
nor I_1(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_2(n_573_1_r_4,G2_0_l_4,n16_4);
nor I_3(n_549_1_r_4,n22_4,n23_4);
nand I_4(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_5(n19_4,blif_clk_net_1_r_6,n4_6,ACVQN2_3_r_4,);
nor I_6(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_7(n19_4,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_4,);
not I_8(P6_5_r_4,P6_5_r_internal_4);
or I_9(n_431_0_l_4,IN_8_0_l_4,n26_4);
DFFARX1 I_10(n_431_0_l_4,blif_clk_net_1_r_6,n4_6,G78_0_l_4,);
DFFARX1 I_11(IN_2_5_l_4,blif_clk_net_1_r_6,n4_6,ACVQN1_5_l_4,);
not I_12(n16_4,ACVQN1_5_l_4);
DFFARX1 I_13(IN_1_5_l_4,blif_clk_net_1_r_6,n4_6,n17_internal_4,);
not I_14(n17_4,n17_internal_4);
nor I_15(n4_1_r_4,n30_4,n31_4);
nand I_16(n19_4,G1_0_l_4,n33_4);
DFFARX1 I_17(G78_0_l_4,blif_clk_net_1_r_6,n4_6,n15_internal_4,);
not I_18(n15_4,n15_internal_4);
DFFARX1 I_19(ACVQN1_5_l_4,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_4,);
and I_20(n20_4,IN_11_0_l_4,n16_4);
nor I_21(n21_4,G2_0_l_4,IN_10_0_l_4);
nand I_22(n22_4,G78_0_l_4,n25_4);
nand I_23(n23_4,IN_11_0_l_4,n24_4);
not I_24(n24_4,G2_0_l_4);
not I_25(n25_4,IN_10_0_l_4);
and I_26(n26_4,IN_2_0_l_4,n27_4);
nor I_27(n27_4,IN_4_0_l_4,n28_4);
not I_28(n28_4,G1_0_l_4);
not I_29(n29_4,n30_4);
nand I_30(n30_4,IN_7_0_l_4,n32_4);
nand I_31(n31_4,IN_11_0_l_4,n25_4);
nor I_32(n32_4,G2_0_l_4,n33_4);
not I_33(n33_4,IN_5_0_l_4);
DFFARX1 I_34(n4_1_r_6,blif_clk_net_1_r_6,n4_6,G42_1_r_6,);
nor I_35(n_572_1_r_6,n27_6,n28_6);
nand I_36(n_573_1_r_6,n18_6,n19_6);
nor I_37(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_38(n_569_1_r_6,n19_6,n20_6);
nor I_39(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_40(N1_4_r_6,blif_clk_net_1_r_6,n4_6,G199_4_r_6,);
DFFARX1 I_41(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,G214_4_r_6,);
DFFARX1 I_42(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_6,);
not I_43(P6_5_r_6,P6_5_r_internal_6);
and I_44(N3_2_l_6,n23_6,n_572_1_r_4);
not I_45(n4_6,blif_reset_net_1_r_6);
DFFARX1 I_46(N3_2_l_6,blif_clk_net_1_r_6,n4_6,n27_6,);
not I_47(n17_6,n27_6);
DFFARX1 I_48(G42_1_r_4,blif_clk_net_1_r_6,n4_6,n28_6,);
DFFARX1 I_49(ACVQN1_5_r_4,blif_clk_net_1_r_6,n4_6,n26_6,);
and I_50(N1_4_l_6,n25_6,n_569_1_r_4);
DFFARX1 I_51(N1_4_l_6,blif_clk_net_1_r_6,n4_6,n29_6,);
not I_52(n18_6,n29_6);
DFFARX1 I_53(n_572_1_r_4,blif_clk_net_1_r_6,n4_6,G214_4_l_6,);
not I_54(n12_6,G214_4_l_6);
nor I_55(n4_1_r_6,n28_6,n22_6);
nor I_56(N1_4_r_6,n12_6,n24_6);
nor I_57(n_42_2_l_6,G42_1_r_4,P6_5_r_4);
DFFARX1 I_58(G214_4_l_6,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_6,);
nand I_59(n19_6,n26_6,ACVQN2_3_r_4);
not I_60(n20_6,n_42_2_l_6);
nor I_61(n21_6,n17_6,n28_6);
and I_62(n22_6,n26_6,ACVQN2_3_r_4);
nand I_63(n23_6,G42_1_r_4,n_573_1_r_4);
nor I_64(n24_6,n17_6,n18_6);
nand I_65(n25_6,n_549_1_r_4,n_266_and_0_3_r_4);
endmodule


