module test_I11150(I8360,I8267,I8496,I1477,I1470,I11150);
input I8360,I8267,I8496,I1477,I1470;
output I11150;
wire I10647,I9508,I9576,I9542,I8202,I8181,I9474,I8592,I8184,I9525,I9491;
not I_0(I10647,I1477);
nand I_1(I9508,I8202);
nor I_2(I9576,I8181,I8202);
DFFARX1 I_3(I9525,I1470,I9491,,,I9542,);
nand I_4(I8202,I8267,I8496);
and I_5(I8181,I8360,I8592);
or I_6(I9474,I9576,I9542);
DFFARX1 I_7(I1470,,,I8592,);
DFFARX1 I_8(I1470,,,I8184,);
DFFARX1 I_9(I9474,I1470,I10647,,,I11150,);
and I_10(I9525,I9508,I8184);
not I_11(I9491,I1477);
endmodule


