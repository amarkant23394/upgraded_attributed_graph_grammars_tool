module test_I6127(I1477,I2328,I2170,I2557,I2509,I1470,I6127);
input I1477,I2328,I2170,I2557,I2509,I1470;
output I6127;
wire I2167,I4629,I6110,I4544,I4824,I2633,I2143,I5751,I4533,I5013,I4807,I2173,I2181,I4996,I4509;
nand I_0(I2167,I2633,I2328);
nor I_1(I4629,I2167,I2173);
DFFARX1 I_2(I4509,I1470,I5751,,,I6110,);
not I_3(I4544,I1477);
and I_4(I4824,I4807,I2143);
DFFARX1 I_5(I1470,I2181,,,I2633,);
DFFARX1 I_6(I2557,I1470,I2181,,,I2143,);
not I_7(I5751,I1477);
or I_8(I4533,I4824,I4629);
or I_9(I5013,I4824,I4996);
DFFARX1 I_10(I2170,I1470,I4544,,,I4807,);
nand I_11(I2173,I2557,I2509);
not I_12(I2181,I1477);
and I_13(I6127,I6110,I4533);
and I_14(I4996,I4629);
DFFARX1 I_15(I5013,I1470,I4544,,,I4509,);
endmodule


