module test_I1911(I1444,I1328,I1294,I1301,I1911);
input I1444,I1328,I1294,I1301;
output I1911;
wire I1310,I1937,I1342,I2070,I1509,I2389,I2406,I1577,I2488;
nand I_0(I1911,I2070,I2488);
DFFARX1 I_1(I1577,I1294,I1342,,,I1310,);
not I_2(I1937,I1301);
not I_3(I1342,I1301);
not I_4(I2070,I1310);
DFFARX1 I_5(I1294,I1342,,,I1509,);
DFFARX1 I_6(I1328,I1294,I1937,,,I2389,);
not I_7(I2406,I2389);
and I_8(I1577,I1509,I1444);
not I_9(I2488,I2406);
endmodule


