module test_I11026(I1477,I9471,I9771,I8193,I9576,I1470,I11026);
input I1477,I9471,I9771,I8193,I9576,I1470;
output I11026;
wire I10647,I10664,I11009,I10715,I9638,I9816,I10732,I9491,I9477,I9468,I9833,I9465,I9621,I9864;
not I_0(I10647,I1477);
not I_1(I10664,I9471);
DFFARX1 I_2(I9468,I1470,I10647,,,I11009,);
nor I_3(I11026,I11009,I10732);
nor I_4(I10715,I10664,I9477);
nor I_5(I9638,I9621,I9576);
DFFARX1 I_6(I8193,I1470,I9491,,,I9816,);
nand I_7(I10732,I10715,I9465);
not I_8(I9491,I1477);
nor I_9(I9477,I9771,I9833);
DFFARX1 I_10(I9864,I1470,I9491,,,I9468,);
and I_11(I9833,I9816);
nand I_12(I9465,I9816,I9638);
DFFARX1 I_13(I1470,I9491,,,I9621,);
nor I_14(I9864,I9816,I9621);
endmodule


