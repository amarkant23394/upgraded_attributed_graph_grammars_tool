module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_12,blif_reset_net_1_r_12,G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_12,blif_reset_net_1_r_12;
output G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,n_431_0_l_12,n8_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_12,n8_12,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_12,n8_12,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_12,n8_12,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_12,n8_12,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_12,n8_12,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_12,n8_12,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_12,n8_12,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_12,n8_12,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_12,n8_12,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_12,blif_clk_net_1_r_12,n8_12,G42_1_r_12,);
nor I_31(n_572_1_r_12,n29_12,n30_12);
nand I_32(n_573_1_r_12,n26_12,n27_12);
nor I_33(n_549_1_r_12,n33_12,n34_12);
and I_34(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_35(N3_2_r_12,blif_clk_net_1_r_12,n8_12,G199_2_r_12,);
DFFARX1 I_36(n3_12,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_12,);
not I_37(P6_5_r_12,P6_5_r_internal_12);
or I_38(n_431_0_l_12,n36_12,G42_1_r_10);
not I_39(n8_12,blif_reset_net_1_r_12);
DFFARX1 I_40(n_431_0_l_12,blif_clk_net_1_r_12,n8_12,n41_12,);
DFFARX1 I_41(n_572_1_r_10,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_12,);
not I_42(n22_12,ACVQN1_5_l_12);
DFFARX1 I_43(ACVQN2_3_r_10,blif_clk_net_1_r_12,n8_12,n42_12,);
nor I_44(n4_1_r_12,n41_12,n31_12);
nor I_45(N3_2_r_12,n22_12,n40_12);
not I_46(n3_12,n39_12);
DFFARX1 I_47(ACVQN1_5_l_12,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_12,);
and I_48(n26_12,G42_1_r_10,n_572_1_r_10);
nor I_49(n27_12,n28_12,n29_12);
not I_50(n28_12,n_573_1_r_10);
nand I_51(n29_12,n31_12,n32_12);
nand I_52(n30_12,n42_12,n_573_1_r_10);
not I_53(n31_12,n_573_1_r_10);
not I_54(n32_12,G199_2_r_10);
nand I_55(n33_12,n31_12,n35_12);
nand I_56(n34_12,G42_1_r_10,n_572_1_r_10);
nand I_57(n35_12,n41_12,n42_12);
and I_58(n36_12,n37_12,n_266_and_0_3_r_10);
nor I_59(n37_12,n38_12,n_42_2_r_10);
not I_60(n38_12,n_549_1_r_10);
nor I_61(n39_12,n38_12,n_572_1_r_10);
nor I_62(n40_12,n39_12,n_573_1_r_10);
endmodule


