module test_I7122(I5659,I1477,I5122,I3380,I1470,I3453,I7122);
input I5659,I1477,I5122,I3380,I1470,I3453;
output I7122;
wire I5076,I5156,I5079,I5105,I7105,I5187,I3371,I3353,I5088,I5139,I3637,I7088,I5204;
DFFARX1 I_0(I5204,I1470,I5105,,,I5076,);
and I_1(I7122,I7105,I5076);
nand I_2(I5156,I5139,I3371);
DFFARX1 I_3(I5156,I1470,I5105,,,I5079,);
not I_4(I5105,I1477);
nor I_5(I7105,I7088,I5079);
nor I_6(I5187,I5122,I3380);
DFFARX1 I_7(I1470,,,I3371,);
and I_8(I3353,I3453,I3637);
DFFARX1 I_9(I5659,I1470,I5105,,,I5088,);
nor I_10(I5139,I3380);
DFFARX1 I_11(I1470,,,I3637,);
not I_12(I7088,I5088);
nand I_13(I5204,I5187,I3353);
endmodule


