module test_I17532(I13908,I13743,I14162,I13758,I16069,I17532);
input I13908,I13743,I14162,I13758,I16069;
output I17532;
wire I15597,I15696,I15832,I16145,I15628,I15679,I13749,I16162;
nor I_0(I15597,I15832,I16162);
nand I_1(I15696,I15679,I13758);
nand I_2(I15832,I15628,I13749);
not I_3(I17532,I15597);
not I_4(I16145,I16069);
not I_5(I15628,I13743);
nor I_6(I15679,I15628);
nand I_7(I13749,I14162,I13908);
and I_8(I16162,I15696,I16145);
endmodule


