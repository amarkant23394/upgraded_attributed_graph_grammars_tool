module test_I14777(I1477,I13296,I14404,I1470,I13508,I14777);
input I1477,I13296,I14404,I1470,I13508;
output I14777;
wire I14554,I14667,I14421,I13601,I13186,I14650,I13165,I14537,I14370,I13197,I13635,I13248,I13159,I13618,I14438,I13189,I14571,I14588;
not I_0(I14554,I14537);
and I_1(I14667,I14650,I13189);
DFFARX1 I_2(I14404,I1470,I14370,,,I14421,);
DFFARX1 I_3(I1470,I13197,,,I13601,);
nor I_4(I13186,I13601,I13508);
DFFARX1 I_5(I13165,I1470,I14370,,,I14650,);
DFFARX1 I_6(I13248,I1470,I13197,,,I13165,);
DFFARX1 I_7(I1470,I14370,,,I14537,);
not I_8(I14370,I1477);
not I_9(I13197,I1477);
and I_10(I13635,I13296,I13618);
DFFARX1 I_11(I1470,I13197,,,I13248,);
DFFARX1 I_12(I13508,I1470,I13197,,,I13159,);
nand I_13(I13618,I13601);
nor I_14(I14438,I13159,I13186);
DFFARX1 I_15(I13635,I1470,I13197,,,I13189,);
or I_16(I14777,I14667,I14588);
nor I_17(I14571,I14421,I14554);
and I_18(I14588,I14438,I14571);
endmodule


