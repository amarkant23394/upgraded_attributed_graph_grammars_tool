module test_I4034(I2878,I1447,I1477,I1470,I2980,I4034);
input I2878,I1447,I1477,I1470,I2980;
output I4034;
wire I2730,I2721,I2759,I4017,I3155,I4000,I3076,I2724,I3983;
not I_0(I2730,I3076);
nand I_1(I2721,I2980,I2878);
not I_2(I2759,I1477);
and I_3(I4017,I4000,I2730);
or I_4(I3155,I3076);
nand I_5(I4000,I2721,I2724);
DFFARX1 I_6(I1447,I1470,I2759,,,I3076,);
DFFARX1 I_7(I4017,I1470,I3983,,,I4034,);
DFFARX1 I_8(I3155,I1470,I2759,,,I2724,);
not I_9(I3983,I1477);
endmodule


