module test_final(G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_12,blif_reset_net_1_r_12,G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12);
input G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_12,blif_reset_net_1_r_12;
output G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12;
wire G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_569_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0,n4_1_l_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n_431_0_l_12,n8_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12;
DFFARX1 I_0(n4_1_r_0,blif_clk_net_1_r_12,n8_12,G42_1_r_0,);
nor I_1(n_572_1_r_0,IN_5_1_l_0,n23_0);
nand I_2(n_573_1_r_0,n21_0,n22_0);
nand I_3(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_4(n_569_1_r_0,n21_0,n26_0);
nor I_5(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_6(N3_2_r_0,blif_clk_net_1_r_12,n8_12,G199_2_r_0,);
DFFARX1 I_7(N1_4_r_0,blif_clk_net_1_r_12,n8_12,G199_4_r_0,);
DFFARX1 I_8(n2_0,blif_clk_net_1_r_12,n8_12,G214_4_r_0,);
nor I_9(n4_1_l_0,G18_1_l_0,IN_1_1_l_0);
DFFARX1 I_10(n4_1_l_0,blif_clk_net_1_r_12,n8_12,n37_0,);
DFFARX1 I_11(IN_1_3_l_0,blif_clk_net_1_r_12,n8_12,n38_0,);
not I_12(n20_0,n38_0);
DFFARX1 I_13(IN_2_3_l_0,blif_clk_net_1_r_12,n8_12,ACVQN1_3_l_0,);
nor I_14(n4_1_r_0,IN_10_1_l_0,n23_0);
nor I_15(N3_2_r_0,n31_0,n32_0);
nor I_16(N1_4_r_0,n29_0,n32_0);
not I_17(n2_0,n31_0);
nor I_18(n21_0,IN_9_1_l_0,n37_0);
not I_19(n22_0,IN_5_1_l_0);
nand I_20(n23_0,n20_0,n30_0);
nand I_21(n24_0,n38_0,n25_0);
nor I_22(n25_0,IN_9_1_l_0,IN_10_1_l_0);
not I_23(n26_0,IN_10_1_l_0);
not I_24(n27_0,n29_0);
nor I_25(n28_0,G15_1_l_0,IN_7_1_l_0);
nand I_26(n29_0,n26_0,n33_0);
not I_27(n30_0,IN_9_1_l_0);
nand I_28(n31_0,IN_4_3_l_0,ACVQN1_3_l_0);
and I_29(n32_0,n35_0,n36_0);
nand I_30(n33_0,IN_4_1_l_0,n34_0);
not I_31(n34_0,G15_1_l_0);
nor I_32(n35_0,G18_1_l_0,G15_1_l_0);
nor I_33(n36_0,IN_5_1_l_0,IN_7_1_l_0);
DFFARX1 I_34(n4_1_r_12,blif_clk_net_1_r_12,n8_12,G42_1_r_12,);
nor I_35(n_572_1_r_12,n29_12,n30_12);
nand I_36(n_573_1_r_12,n26_12,n27_12);
nor I_37(n_549_1_r_12,n33_12,n34_12);
and I_38(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_39(N3_2_r_12,blif_clk_net_1_r_12,n8_12,G199_2_r_12,);
DFFARX1 I_40(n3_12,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_12,);
not I_41(P6_5_r_12,P6_5_r_internal_12);
or I_42(n_431_0_l_12,n36_12,G199_4_r_0);
not I_43(n8_12,blif_reset_net_1_r_12);
DFFARX1 I_44(n_431_0_l_12,blif_clk_net_1_r_12,n8_12,n41_12,);
DFFARX1 I_45(n_573_1_r_0,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_12,);
not I_46(n22_12,ACVQN1_5_l_12);
DFFARX1 I_47(n_549_1_r_0,blif_clk_net_1_r_12,n8_12,n42_12,);
nor I_48(n4_1_r_12,n41_12,n31_12);
nor I_49(N3_2_r_12,n22_12,n40_12);
not I_50(n3_12,n39_12);
DFFARX1 I_51(ACVQN1_5_l_12,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_12,);
and I_52(n26_12,G42_1_r_0,G199_2_r_0);
nor I_53(n27_12,n28_12,n29_12);
not I_54(n28_12,G214_4_r_0);
nand I_55(n29_12,n31_12,n32_12);
nand I_56(n30_12,n42_12,G214_4_r_0);
not I_57(n31_12,n_572_1_r_0);
not I_58(n32_12,n_573_1_r_0);
nand I_59(n33_12,n31_12,n35_12);
nand I_60(n34_12,G42_1_r_0,G199_2_r_0);
nand I_61(n35_12,n41_12,n42_12);
and I_62(n36_12,n37_12,n_572_1_r_0);
nor I_63(n37_12,n38_12,G42_1_r_0);
not I_64(n38_12,n_42_2_r_0);
nor I_65(n39_12,n38_12,G199_2_r_0);
nor I_66(n40_12,n39_12,n_572_1_r_0);
endmodule


