module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_5_r_15,n9_15,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
and I_34(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_35(N1508_0_r_15,n55_15,N1371_0_r_12);
nor I_36(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_37(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_38(N1372_4_r_15,n39_15);
nor I_39(N1508_4_r_15,n39_15,n43_15);
nand I_40(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_41(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_42(n_576_5_r_15,n31_15,n32_15);
not I_43(n_102_5_r_15,n33_15);
nand I_44(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_45(N1507_6_r_15,n42_15,n46_15);
nand I_46(N1508_6_r_15,n39_15,n40_15);
nand I_47(n_431_5_r_15,n36_15,n37_15);
not I_48(n9_15,blif_reset_net_5_r_15);
nor I_49(n31_15,n33_15,n34_15);
nor I_50(n32_15,n44_15,N6147_9_r_12);
nor I_51(n33_15,n54_15,n55_15);
nand I_52(n34_15,n49_15,N1508_0_r_12);
nand I_53(n35_15,N1507_6_r_12,n_572_7_r_12);
not I_54(n36_15,n32_15);
nand I_55(n37_15,n34_15,n38_15);
not I_56(n38_15,n46_15);
nand I_57(n39_15,n38_15,n41_15);
nand I_58(n40_15,n41_15,n42_15);
and I_59(n41_15,n51_15,n_569_7_r_12);
and I_60(n42_15,n47_15,n_572_7_r_12);
and I_61(n43_15,n34_15,n36_15);
or I_62(n44_15,N1508_6_r_12,G42_7_r_12);
not I_63(n45_15,N1372_1_r_15);
nand I_64(n46_15,n53_15,n_572_7_r_12);
nor I_65(n47_15,n34_15,n48_15);
not I_66(n48_15,N1507_6_r_12);
and I_67(n49_15,n50_15,n_549_7_r_12);
nand I_68(n50_15,n51_15,n52_15);
nand I_69(n51_15,N1371_0_r_12,n_549_7_r_12);
not I_70(n52_15,n_569_7_r_12);
nor I_71(n53_15,n48_15,N1508_0_r_12);
nor I_72(n54_15,G42_7_r_12,n_572_7_r_12);
not I_73(n55_15,N1507_6_r_12);
endmodule


