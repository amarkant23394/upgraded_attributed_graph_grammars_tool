module test_I11296(I9320,I1477,I11508,I9083,I1470,I11327,I11296);
input I9320,I1477,I11508,I9083,I1470,I11327;
output I11296;
wire I8824,I8836,I9179,I11689,I11559,I11395,I11542,I9210,I8848,I11672,I11378,I9066,I11525,I8833,I11310,I8851;
nand I_0(I8824,I9083);
nand I_1(I11296,I11559,I11689);
nand I_2(I8836,I9320,I9210);
DFFARX1 I_3(I1470,,,I9179,);
nor I_4(I11689,I11672,I11395);
DFFARX1 I_5(I11542,I1470,I11310,,,I11559,);
nand I_6(I11395,I11378,I8851);
or I_7(I11542,I11525,I8833);
nor I_8(I9210,I9179);
nor I_9(I8848,I9083);
DFFARX1 I_10(I8836,I1470,I11310,,,I11672,);
nor I_11(I11378,I11327,I8848);
DFFARX1 I_12(I1470,,,I9066,);
and I_13(I11525,I11508,I8824);
not I_14(I8833,I9179);
not I_15(I11310,I1477);
or I_16(I8851,I9083,I9066);
endmodule


