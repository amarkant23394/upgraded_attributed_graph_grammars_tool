module test_I11576(I11508,I1477,I9083,I1470,I11327,I11576);
input I11508,I1477,I9083,I1470,I11327;
output I11576;
wire I11378,I8824,I11542,I11412,I8851,I9066,I11525,I8833,I11395,I9179,I8848,I11559,I11310;
nor I_0(I11576,I11559,I11412);
nor I_1(I11378,I11327,I8848);
nand I_2(I8824,I9083);
or I_3(I11542,I11525,I8833);
not I_4(I11412,I11395);
or I_5(I8851,I9083,I9066);
DFFARX1 I_6(I1470,,,I9066,);
and I_7(I11525,I11508,I8824);
not I_8(I8833,I9179);
nand I_9(I11395,I11378,I8851);
DFFARX1 I_10(I1470,,,I9179,);
nor I_11(I8848,I9083);
DFFARX1 I_12(I11542,I1470,I11310,,,I11559,);
not I_13(I11310,I1477);
endmodule


