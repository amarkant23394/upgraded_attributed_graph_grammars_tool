module test_I2268(I1444,I1322,I1294,I1797,I1301,I2268);
input I1444,I1322,I1294,I1797,I1301;
output I2268;
wire I1319,I1971,I2251,I1342,I2234,I2070,I1988,I1334,I1304,I1954,I1509,I1310,I1577;
and I_0(I2268,I2070,I2251);
DFFARX1 I_1(I1294,I1342,,,I1319,);
nor I_2(I1971,I1310,I1319);
nand I_3(I2251,I2234,I1988);
not I_4(I1342,I1301);
nand I_5(I2234,I1954,I1304);
not I_6(I2070,I1310);
nand I_7(I1988,I1971,I1334);
DFFARX1 I_8(I1797,I1294,I1342,,,I1334,);
DFFARX1 I_9(I1509,I1294,I1342,,,I1304,);
not I_10(I1954,I1322);
DFFARX1 I_11(I1294,I1342,,,I1509,);
DFFARX1 I_12(I1577,I1294,I1342,,,I1310,);
and I_13(I1577,I1509,I1444);
endmodule


