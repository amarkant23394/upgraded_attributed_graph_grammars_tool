module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_8_r_6,n9_6,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
nor I_44(N1371_0_r_6,n30_6,n33_6);
nor I_45(N1508_0_r_6,n33_6,n44_6);
not I_46(N1372_1_r_6,n41_6);
nor I_47(N1508_1_r_6,n40_6,n41_6);
nor I_48(N1507_6_r_6,n39_6,n45_6);
nor I_49(N1508_6_r_6,n37_6,n38_6);
nor I_50(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_51(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_52(N6147_9_r_6,n32_6,n33_6);
nor I_53(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_54(I_BUFF_1_9_r_6,n37_6);
not I_55(N1372_10_r_6,n43_6);
nor I_56(N1508_10_r_6,n42_6,n43_6);
nor I_57(N3_8_r_6,n36_6,N1507_6_r_10);
not I_58(n9_6,blif_reset_net_8_r_6);
nor I_59(n30_6,n53_6,N1508_0_r_10);
not I_60(n31_6,n36_6);
nor I_61(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_62(n33_6,N1507_6_r_10);
not I_63(n34_6,n35_6);
nand I_64(n35_6,n49_6,N1508_4_r_10);
nand I_65(n36_6,n51_6,N6147_9_r_10);
nand I_66(n37_6,n54_6,N6134_9_r_10);
or I_67(n38_6,n35_6,n39_6);
nor I_68(n39_6,n40_6,n45_6);
and I_69(n40_6,n46_6,n47_6);
nand I_70(n41_6,n30_6,n31_6);
nor I_71(n42_6,n34_6,n40_6);
nand I_72(n43_6,n30_6,N1507_6_r_10);
nor I_73(n44_6,n31_6,n40_6);
nor I_74(n45_6,n35_6,n36_6);
nor I_75(n46_6,N6147_3_r_10,N1508_4_r_10);
or I_76(n47_6,n48_6,G199_8_r_10);
nor I_77(n48_6,N1371_0_r_10,N1508_0_r_10);
and I_78(n49_6,n50_6,N6147_2_r_10);
nand I_79(n50_6,n51_6,n52_6);
nand I_80(n51_6,N6147_2_r_10,N1507_6_r_10);
not I_81(n52_6,N6147_9_r_10);
nor I_82(n53_6,N1508_6_r_10,n_42_8_r_10);
or I_83(n54_6,N1508_6_r_10,n_42_8_r_10);
endmodule


