module test_I5266(I3504,I1495,I3555,I3747,I5266);
input I3504,I1495,I3555,I3747;
output I5266;
wire I3846,I3521,I3380,I5249;
not I_0(I5266,I5249);
nor I_1(I3846,I3747,I3555);
nor I_2(I3521,I3504,I1495);
nand I_3(I3380,I3521,I3846);
not I_4(I5249,I3380);
endmodule


