module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14,I_BUFF_1_9_r_14,N3_8_l_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_14,n47_14,n30_14);
nor I_1(N1508_0_r_14,n30_14,n41_14);
nor I_2(N1507_6_r_14,n37_14,n44_14);
nor I_3(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_4(n4_7_r_14,blif_clk_net_7_r_1,n9_1,G42_7_r_14,);
nor I_5(n_572_7_r_14,n28_14,n29_14);
nand I_6(n_573_7_r_14,n26_14,n27_14);
nor I_7(n_549_7_r_14,n31_14,n32_14);
nand I_8(n_569_7_r_14,n26_14,n30_14);
nor I_9(n_452_7_r_14,n47_14,n28_14);
nor I_10(N6147_9_r_14,n36_14,n37_14);
nor I_11(N6134_9_r_14,n28_14,n36_14);
not I_12(I_BUFF_1_9_r_14,n26_14);
and I_13(N3_8_l_14,IN_6_8_l_14,n38_14);
DFFARX1 I_14(N3_8_l_14,blif_clk_net_7_r_1,n9_1,n47_14,);
nor I_15(n4_7_r_14,n47_14,n35_14);
nand I_16(n26_14,IN_1_10_l_14,IN_2_10_l_14);
not I_17(n27_14,n28_14);
nor I_18(n28_14,IN_2_0_l_14,n43_14);
not I_19(n29_14,n33_14);
not I_20(n30_14,n31_14);
nor I_21(n31_14,IN_1_3_l_14,n46_14);
and I_22(n32_14,n33_14,n34_14);
nand I_23(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_24(n34_14,n42_14,n43_14);
nor I_25(n35_14,IN_1_8_l_14,IN_3_8_l_14);
nor I_26(n36_14,n47_14,n34_14);
not I_27(n37_14,n35_14);
nand I_28(n38_14,IN_2_8_l_14,IN_3_8_l_14);
nand I_29(n39_14,n29_14,n40_14);
nand I_30(n40_14,n27_14,n37_14);
nor I_31(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_32(n42_14,IN_3_0_l_14,IN_4_0_l_14);
not I_33(n43_14,IN_1_0_l_14);
nor I_34(n44_14,n27_14,n33_14);
or I_35(n45_14,IN_3_10_l_14,IN_4_10_l_14);
or I_36(n46_14,IN_2_3_l_14,IN_3_3_l_14);
and I_37(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_38(N1508_0_r_1,n40_1,n44_1);
nor I_39(N1507_6_r_1,n43_1,n49_1);
nor I_40(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_41(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_42(n_572_7_r_1,n29_1,n30_1);
not I_43(n_573_7_r_1,n_452_7_r_1);
nor I_44(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_45(n_569_7_r_1,n30_1,n31_1);
nor I_46(n_452_7_r_1,n30_1,n32_1);
nor I_47(N6147_9_r_1,n35_1,n36_1);
nand I_48(N6134_9_r_1,n38_1,n39_1);
not I_49(I_BUFF_1_9_r_1,n40_1);
nor I_50(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_51(n9_1,blif_reset_net_7_r_1);
nor I_52(n29_1,n34_1,n_549_7_r_14);
nor I_53(n30_1,n33_1,n34_1);
nor I_54(n31_1,n54_1,N1508_6_r_14);
not I_55(n32_1,n48_1);
nor I_56(n33_1,N1508_0_r_14,n_572_7_r_14);
not I_57(n34_1,N1507_6_r_14);
nor I_58(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_59(n36_1,n29_1);
not I_60(n37_1,n41_1);
nand I_61(n38_1,I_BUFF_1_9_r_1,N1508_6_r_14);
nand I_62(n39_1,n37_1,n40_1);
nand I_63(n40_1,n_573_7_r_14,n_452_7_r_14);
nand I_64(n41_1,n52_1,N6147_9_r_14);
or I_65(n42_1,n36_1,n43_1);
nor I_66(n43_1,n32_1,n49_1);
nand I_67(n44_1,n45_1,n46_1);
nand I_68(n45_1,n47_1,n48_1);
not I_69(n46_1,N1508_6_r_14);
not I_70(n47_1,n31_1);
nand I_71(n48_1,n50_1,N6134_9_r_14);
nor I_72(n49_1,n41_1,n47_1);
and I_73(n50_1,n51_1,n_569_7_r_14);
nand I_74(n51_1,n52_1,n53_1);
nand I_75(n52_1,G42_7_r_14,N1507_6_r_14);
not I_76(n53_1,N6147_9_r_14);
or I_77(n54_1,N1371_0_r_14,N1508_0_r_14);
nor I_78(n55_1,n29_1,N1508_6_r_14);
endmodule


