module test_I10137(I8011,I1477,I1470,I10137);
input I8011,I1477,I1470;
output I10137;
wire I8107,I8090,I7570,I8028,I7553,I10052,I8124,I7977;
not I_0(I8107,I8090);
DFFARX1 I_1(I1470,I7570,,,I8090,);
not I_2(I7570,I1477);
and I_3(I8028,I7977,I8011);
DFFARX1 I_4(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_5(I8124,I1470,I7570,,,I7553,);
not I_6(I10052,I1477);
or I_7(I8124,I8107,I8028);
DFFARX1 I_8(I1470,I7570,,,I7977,);
endmodule


