module test_I13635(I1477,I11395,I11429,I1470,I11327,I13635);
input I1477,I11395,I11429,I1470,I11327;
output I13635;
wire I11302,I11278,I13601,I8827,I11847,I11624,I13313,I13197,I11299,I13296,I13618,I11672,I11293,I11310,I11864;
DFFARX1 I_0(I11864,I1470,I11310,,,I11302,);
DFFARX1 I_1(I11624,I1470,I11310,,,I11278,);
DFFARX1 I_2(I11299,I1470,I13197,,,I13601,);
DFFARX1 I_3(I1470,,,I8827,);
nand I_4(I11847,I11395);
nand I_5(I11624,I11327,I8827);
DFFARX1 I_6(I11293,I1470,I13197,,,I13313,);
not I_7(I13197,I1477);
nor I_8(I11299,I11395,I11429);
and I_9(I13635,I13296,I13618);
nor I_10(I13296,I11278,I11302);
nand I_11(I13618,I13601,I13313);
DFFARX1 I_12(I1470,I11310,,,I11672,);
not I_13(I11293,I11672);
not I_14(I11310,I1477);
and I_15(I11864,I11624,I11847);
endmodule


