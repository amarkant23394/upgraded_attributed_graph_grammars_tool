module test_I16818(I1477,I16818);
input I1477;
output I16818;
wire ;
not I_0(I16818,I1477);
endmodule


