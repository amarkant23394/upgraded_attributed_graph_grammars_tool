module test_I13165(I11720,I1477,I11830,I1470,I13165);
input I11720,I1477,I11830,I1470;
output I13165;
wire I13214,I13231,I11290,I13197,I11275,I11302,I13248;
nand I_0(I13214,I11275,I11302);
and I_1(I13231,I13214,I11290);
nand I_2(I11290,I11830,I11720);
not I_3(I13197,I1477);
DFFARX1 I_4(I1470,,,I11275,);
DFFARX1 I_5(I1470,,,I11302,);
DFFARX1 I_6(I13248,I1470,I13197,,,I13165,);
DFFARX1 I_7(I13231,I1470,I13197,,,I13248,);
endmodule


