module test_I14856(I13231,I1477,I1470,I13525,I14856);
input I13231,I1477,I1470,I13525;
output I14856;
wire I13361,I13313,I13601,I13162,I13183,I13197,I14404,I14387,I14421,I13186,I14808,I13171,I13248,I14370;
DFFARX1 I_0(I13313,I1470,I13197,,,I13361,);
DFFARX1 I_1(I1470,I13197,,,I13313,);
nor I_2(I14856,I14808,I14421);
DFFARX1 I_3(I1470,I13197,,,I13601,);
and I_4(I13162,I13248,I13361);
nand I_5(I13183,I13601,I13525);
not I_6(I13197,I1477);
and I_7(I14404,I14387,I13183);
nand I_8(I14387,I13171,I13186);
DFFARX1 I_9(I14404,I1470,I14370,,,I14421,);
nor I_10(I13186,I13601);
DFFARX1 I_11(I13162,I1470,I14370,,,I14808,);
nand I_12(I13171,I13248);
DFFARX1 I_13(I13231,I1470,I13197,,,I13248,);
not I_14(I14370,I1477);
endmodule


