module test_I17399(I1477,I15832,I17611,I16069,I17430,I1470,I17399);
input I1477,I15832,I17611,I16069,I17430,I1470;
output I17399;
wire I17413,I15585,I17792,I15582,I15600,I15815,I15959,I17498,I15928,I15597,I17628,I17775,I17662,I17645,I15573,I17481;
not I_0(I17413,I1477);
nand I_1(I15585,I16069,I15959);
nor I_2(I17792,I17775,I17498);
not I_3(I15582,I15928);
nand I_4(I17399,I17662,I17792);
or I_5(I15600,I15832,I15815);
DFFARX1 I_6(I1470,,,I15815,);
nor I_7(I15959,I15928);
nand I_8(I17498,I17481,I15600);
DFFARX1 I_9(I1470,,,I15928,);
nor I_10(I15597,I15832);
and I_11(I17628,I17611,I15573);
DFFARX1 I_12(I15585,I1470,I17413,,,I17775,);
DFFARX1 I_13(I17645,I1470,I17413,,,I17662,);
or I_14(I17645,I17628,I15582);
nand I_15(I15573,I15832);
nor I_16(I17481,I17430,I15597);
endmodule


