module Benchmark_testing100_removed(I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I163,I170,I735,I745,I755,I765,I775,I785,I795,I805,I815,I1437,I1447,I1457,I1467,I1477,I1487,I1497,I1507,I1517);
input I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I163,I170;
output I735,I745,I755,I765,I775,I785,I795,I805,I815,I1437,I1447,I1457,I1467,I1477,I1487,I1497,I1507,I1517;
wire I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I163,I170,I179,I206,I224,I233,I251,I269,I296,I314,I332,I350,I359,I377,I395,I422,I431,I449,I467,I485,I503,I530,I539,I566,I575,I593,I611,I629,I647,I674,I683,I701,I719,I827,I854,I863,I890,I908,I917,I935,I953,I971,I998,I1007,I1025,I1043,I1070,I1079,I1097,I1115,I1133,I1151,I1178,I1196,I1205,I1223,I1241,I1259,I1286,I1295,I1313,I1331,I1349,I1367,I1385,I1403,I1421;
not I_0 (I179,I170);
dffarx1 I_1 (I100,I163,I179,I206);
dffarx1 I_2 (I206,I163,I179,I224);
not I_3 (I233,I224);
nand I_4 (I251,I148,I124);
and I_5 (I269,I251,I92);
dffarx1 I_6 (I269,I163,I179,I296);
dffarx1 I_7 (I296,I163,I179,I314);
dffarx1 I_8 (I296,I163,I179,I332);
dffarx1 I_9 (I156,I163,I179,I350);
nand I_10 (I359,I350,I84);
not I_11 (I377,I359);
nor I_12 (I395,I206,I377);
dffarx1 I_13 (I132,I163,I179,I422);
not I_14 (I431,I422);
nor I_15 (I449,I431,I233);
nand I_16 (I467,I431,I359);
nand I_17 (I485,I116,I108);
and I_18 (I503,I485,I76);
dffarx1 I_19 (I503,I163,I179,I530);
nor I_20 (I539,I530,I206);
dffarx1 I_21 (I539,I163,I179,I566);
not I_22 (I575,I530);
nor I_23 (I593,I140,I108);
not I_24 (I611,I593);
nor I_25 (I629,I359,I611);
nor I_26 (I647,I575,I629);
dffarx1 I_27 (I647,I163,I179,I674);
nor I_28 (I683,I530,I611);
nor I_29 (I701,I377,I683);
nor I_30 (I719,I530,I593);
r I_31 (I735,I314);
r I_32 (I745,I332);
r I_33 (I755,I395);
r I_34 (I765,I449);
r I_35 (I775,I467);
r I_36 (I785,I566);
r I_37 (I795,I674);
r I_38 (I805,I701);
r I_39 (I815,I719);
not I_40 (I827,I170);
dffarx1 I_41 (I566,I163,I827,I854);
and I_42 (I863,I854,I719);
dffarx1 I_43 (I863,I163,I827,I890);
dffarx1 I_44 (I719,I163,I827,I908);
not I_45 (I917,I467);
not I_46 (I935,I674);
nand I_47 (I953,I935,I917);
nor I_48 (I971,I908,I953);
dffarx1 I_49 (I953,I163,I827,I998);
not I_50 (I1007,I998);
not I_51 (I1025,I332);
nand I_52 (I1043,I935,I1025);
dffarx1 I_53 (I1043,I163,I827,I1070);
not I_54 (I1079,I1070);
not I_55 (I1097,I449);
nand I_56 (I1115,I1097,I566);
and I_57 (I1133,I917,I1115);
nor I_58 (I1151,I1043,I1133);
dffarx1 I_59 (I1151,I163,I827,I1178);
dffarx1 I_60 (I1133,I163,I827,I1196);
nor I_61 (I1205,I449,I395);
nor I_62 (I1223,I1043,I1205);
or I_63 (I1241,I449,I395);
nor I_64 (I1259,I701,I314);
dffarx1 I_65 (I1259,I163,I827,I1286);
not I_66 (I1295,I1286);
nor I_67 (I1313,I1295,I1079);
nand I_68 (I1331,I1295,I908);
not I_69 (I1349,I701);
nand I_70 (I1367,I1349,I1025);
nand I_71 (I1385,I1295,I1367);
nand I_72 (I1403,I1385,I1331);
nand I_73 (I1421,I1367,I1241);
r I_74 (I1437,I1178);
r I_75 (I1447,I971);
r I_76 (I1457,I1421);
r I_77 (I1467,I1403);
r I_78 (I1477,I1223);
r I_79 (I1487,I890);
r I_80 (I1497,I1313);
r I_81 (I1507,I1196);
r I_82 (I1517,I1007);
endmodule


