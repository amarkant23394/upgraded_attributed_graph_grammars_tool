module test_final(IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5,N3_2_l_5,G199_2_l_5,ACVQN2_3_l_5,n13_5,ACVQN1_3_l_5,N1_4_l_5,n21_5,n15_5,n22_5,n4_1_r_5,n11_internal_5,n11_5,n_42_2_l_5,n1_5,P6_5_r_internal_5,n16_5,n17_5,n18_5,n19_5,n20_5,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n4_1_r_5,blif_clk_net_1_r_9,n5_9,G42_1_r_5,);
nor I_1(n_572_1_r_5,n21_5,n22_5);
nand I_2(n_573_1_r_5,n13_5,n16_5);
nor I_3(n_549_1_r_5,n21_5,n17_5);
nand I_4(n_569_1_r_5,n13_5,n15_5);
nor I_5(n_452_1_r_5,n22_5,n_42_2_l_5);
DFFARX1 I_6(G199_2_l_5,blif_clk_net_1_r_9,n5_9,ACVQN2_3_r_5,);
nor I_7(n_266_and_0_3_r_5,n11_5,n16_5);
DFFARX1 I_8(n_42_2_l_5,blif_clk_net_1_r_9,n5_9,ACVQN1_5_r_5,);
not I_9(P6_5_r_5,P6_5_r_internal_5);
and I_10(N3_2_l_5,IN_6_2_l_5,n19_5);
DFFARX1 I_11(N3_2_l_5,blif_clk_net_1_r_9,n5_9,G199_2_l_5,);
DFFARX1 I_12(IN_1_3_l_5,blif_clk_net_1_r_9,n5_9,ACVQN2_3_l_5,);
not I_13(n13_5,ACVQN2_3_l_5);
DFFARX1 I_14(IN_2_3_l_5,blif_clk_net_1_r_9,n5_9,ACVQN1_3_l_5,);
and I_15(N1_4_l_5,IN_6_4_l_5,n20_5);
DFFARX1 I_16(N1_4_l_5,blif_clk_net_1_r_9,n5_9,n21_5,);
not I_17(n15_5,n21_5);
DFFARX1 I_18(IN_3_4_l_5,blif_clk_net_1_r_9,n5_9,n22_5,);
nor I_19(n4_1_r_5,G199_2_l_5,n22_5);
DFFARX1 I_20(ACVQN2_3_l_5,blif_clk_net_1_r_9,n5_9,n11_internal_5,);
not I_21(n11_5,n11_internal_5);
nor I_22(n_42_2_l_5,IN_1_2_l_5,IN_3_2_l_5);
not I_23(n1_5,n18_5);
DFFARX1 I_24(n1_5,blif_clk_net_1_r_9,n5_9,P6_5_r_internal_5,);
not I_25(n16_5,n_42_2_l_5);
nor I_26(n17_5,n22_5,n18_5);
nand I_27(n18_5,IN_4_3_l_5,ACVQN1_3_l_5);
nand I_28(n19_5,IN_2_2_l_5,IN_3_2_l_5);
nand I_29(n20_5,IN_1_4_l_5,IN_2_4_l_5);
DFFARX1 I_30(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_31(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_32(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_33(n_549_1_r_9,n17_9,n18_9);
or I_34(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_35(n_452_1_r_9,n26_9,n25_9);
nor I_36(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_37(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_38(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_39(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_40(N3_2_l_9,n22_9,ACVQN2_3_r_5);
not I_41(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_42(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_43(n16_9,n27_9);
DFFARX1 I_44(n_549_1_r_5,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_45(n15_9,n26_9);
DFFARX1 I_46(G42_1_r_5,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_47(n29_9,n29_internal_9);
and I_48(N1_4_l_9,n24_9,G42_1_r_5);
DFFARX1 I_49(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_50(ACVQN1_5_r_5,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_51(n28_9,n28_internal_9);
nor I_52(n4_1_r_9,n27_9,n26_9);
nor I_53(N3_2_r_9,n15_9,n21_9);
nor I_54(N1_4_r_9,n16_9,n21_9);
nor I_55(n_42_2_l_9,n_452_1_r_5,n_266_and_0_3_r_5);
not I_56(n17_9,n_452_1_r_9);
nand I_57(n18_9,n27_9,n15_9);
nor I_58(n19_9,n29_9,n20_9);
not I_59(n20_9,n_573_1_r_5);
and I_60(n21_9,n23_9,n_573_1_r_5);
nand I_61(n22_9,n_569_1_r_5,n_266_and_0_3_r_5);
nor I_62(n23_9,n29_9,n28_9);
nand I_63(n24_9,n_572_1_r_5,P6_5_r_5);
endmodule


