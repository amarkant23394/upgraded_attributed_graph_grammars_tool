module test_final(IN_1_2_l_2,IN_2_2_l_2,G1_3_l_2,G2_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_5_3_l_2,IN_7_3_l_2,IN_8_3_l_2,IN_10_3_l_2,IN_11_3_l_2,blif_clk_net_3_r_0,blif_reset_net_3_r_0,n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0);
input IN_1_2_l_2,IN_2_2_l_2,G1_3_l_2,G2_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_5_3_l_2,IN_7_3_l_2,IN_8_3_l_2,IN_10_3_l_2,IN_11_3_l_2,blif_clk_net_3_r_0,blif_reset_net_3_r_0;
output n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0;
wire ACVQN2_0_r_2,n_266_and_0_0_r_2,G199_1_r_2,G214_1_r_2,n_429_or_0_3_r_2,G78_3_r_2,n_576_3_r_2,n_102_3_r_2,n_547_3_r_2,n_42_5_r_2,G199_5_r_2,ACVQN1_2_l_2,P6_2_l_2,P6_internal_2_l_2,n_429_or_0_3_l_2,n12_3_l_2,n_431_3_l_2,G78_3_l_2,n_576_3_l_2,n11_3_l_2,n_102_3_l_2,n_547_3_l_2,n13_3_l_2,n14_3_l_2,n15_3_l_2,n16_3_l_2,ACVQN1_0_r_2,N1_1_r_2,n3_1_r_2,n12_3_r_2,n_431_3_r_2,n11_3_r_2,n13_3_r_2,n14_3_r_2,n15_3_r_2,n16_3_r_2,N3_5_r_2,n3_5_r_2,n2_3_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0;
DFFARX1 I_0(P6_2_l_2,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_r_2,);
and I_1(n_266_and_0_0_r_2,n_102_3_l_2,ACVQN1_0_r_2);
DFFARX1 I_2(N1_1_r_2,blif_clk_net_3_r_0,n2_3_r_0,G199_1_r_2,);
DFFARX1 I_3(n_547_3_l_2,blif_clk_net_3_r_0,n2_3_r_0,G214_1_r_2,);
nand I_4(n_429_or_0_3_r_2,ACVQN1_2_l_2,n12_3_r_2);
DFFARX1 I_5(n_431_3_r_2,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_2,);
nand I_6(n_576_3_r_2,ACVQN1_2_l_2,n11_3_r_2);
not I_7(n_102_3_r_2,G78_3_l_2);
nand I_8(n_547_3_r_2,n_102_3_l_2,n13_3_r_2);
nor I_9(n_42_5_r_2,ACVQN1_2_l_2,P6_2_l_2);
DFFARX1 I_10(N3_5_r_2,blif_clk_net_3_r_0,n2_3_r_0,G199_5_r_2,);
DFFARX1 I_11(IN_2_2_l_2,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_2_l_2,);
not I_12(P6_2_l_2,P6_internal_2_l_2);
DFFARX1 I_13(IN_1_2_l_2,blif_clk_net_3_r_0,n2_3_r_0,P6_internal_2_l_2,);
nand I_14(n_429_or_0_3_l_2,G1_3_l_2,n12_3_l_2);
not I_15(n12_3_l_2,IN_5_3_l_2);
or I_16(n_431_3_l_2,IN_8_3_l_2,n14_3_l_2);
DFFARX1 I_17(n_431_3_l_2,blif_clk_net_3_r_0,n2_3_r_0,G78_3_l_2,);
nand I_18(n_576_3_l_2,IN_7_3_l_2,n11_3_l_2);
nor I_19(n11_3_l_2,G2_3_l_2,n12_3_l_2);
not I_20(n_102_3_l_2,G2_3_l_2);
nand I_21(n_547_3_l_2,IN_11_3_l_2,n13_3_l_2);
nor I_22(n13_3_l_2,G2_3_l_2,IN_10_3_l_2);
and I_23(n14_3_l_2,IN_2_3_l_2,n15_3_l_2);
nor I_24(n15_3_l_2,IN_4_3_l_2,n16_3_l_2);
not I_25(n16_3_l_2,G1_3_l_2);
DFFARX1 I_26(G78_3_l_2,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_r_2,);
and I_27(N1_1_r_2,G78_3_l_2,n3_1_r_2);
nand I_28(n3_1_r_2,n_576_3_l_2,n_547_3_l_2);
not I_29(n12_3_r_2,n_429_or_0_3_l_2);
or I_30(n_431_3_r_2,n_429_or_0_3_l_2,n14_3_r_2);
nor I_31(n11_3_r_2,G78_3_l_2,n12_3_r_2);
nor I_32(n13_3_r_2,G78_3_l_2,n_576_3_l_2);
and I_33(n14_3_r_2,n_576_3_l_2,n15_3_r_2);
nor I_34(n15_3_r_2,P6_2_l_2,n16_3_r_2);
not I_35(n16_3_r_2,ACVQN1_2_l_2);
and I_36(N3_5_r_2,n_102_3_l_2,n3_5_r_2);
nand I_37(n3_5_r_2,ACVQN1_2_l_2,n_429_or_0_3_l_2);
nand I_38(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_39(n_431_3_r_0,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_0,);
nand I_40(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_41(n_102_3_r_0,n_42_5_l_0);
nand I_42(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_43(n4_4_r_0,blif_clk_net_3_r_0,n2_3_r_0,G42_4_r_0,);
nor I_44(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_45(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_46(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_47(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_48(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
not I_49(n2_3_r_0,blif_reset_net_3_r_0);
DFFARX1 I_50(n_576_3_r_2,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_0,);
and I_51(n_266_and_0_0_l_0,ACVQN1_0_l_0,G199_5_r_2);
DFFARX1 I_52(n_547_3_r_2,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_0,);
and I_53(N1_1_l_0,n3_1_l_0,G78_3_r_2);
DFFARX1 I_54(N1_1_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_1_l_0,);
DFFARX1 I_55(n_102_3_r_2,blif_clk_net_3_r_0,n2_3_r_0,G214_1_l_0,);
nand I_56(n3_1_l_0,ACVQN2_0_r_2,n_429_or_0_3_r_2);
nor I_57(n_42_5_l_0,G199_1_r_2,n_42_5_r_2);
and I_58(N3_5_l_0,n3_5_l_0,n_266_and_0_0_r_2);
DFFARX1 I_59(N3_5_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_5_l_0,);
nand I_60(n3_5_l_0,G199_1_r_2,G214_1_r_2);
not I_61(n12_3_r_0,G199_1_l_0);
or I_62(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_63(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_64(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_65(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_66(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_67(n16_3_r_0,ACVQN2_0_l_0);
nor I_68(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_69(n_87_4_r_0,G199_5_l_0);
and I_70(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
endmodule


