module test_I1832(I1455,I1207,I1832);
input I1455,I1207;
output I1832;
wire I1535;
not I_0(I1535,I1455);
nand I_1(I1832,I1535,I1207);
endmodule


