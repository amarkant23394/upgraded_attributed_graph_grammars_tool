module test_I2739(I1415,I1431,I1477,I1470,I1407,I2739);
input I1415,I1431,I1477,I1470,I1407;
output I2739;
wire I3217,I2759,I3200,I2980,I2776;
not I_0(I3217,I3200);
not I_1(I2759,I1477);
DFFARX1 I_2(I1431,I1470,I2759,,,I3200,);
nor I_3(I2739,I3217,I2980);
nand I_4(I2980,I2776,I1415);
not I_5(I2776,I1407);
endmodule


