module test_final(G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11,n_431_0_l_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_11,blif_clk_net_1_r_7,n8_7,G42_1_r_11,);
nor I_1(n_572_1_r_11,n29_11,n30_11);
nand I_2(n_573_1_r_11,n26_11,n28_11);
nor I_3(n_549_1_r_11,n27_11,n32_11);
nand I_4(n_569_1_r_11,n45_11,n28_11);
nor I_5(n_452_1_r_11,n43_11,n44_11);
nor I_6(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_7(N3_2_r_11,blif_clk_net_1_r_7,n8_7,G199_2_r_11,);
DFFARX1 I_8(n24_11,blif_clk_net_1_r_7,n8_7,ACVQN2_3_r_11,);
nor I_9(n_266_and_0_3_r_11,n20_11,n37_11);
or I_10(n_431_0_l_11,IN_8_0_l_11,n33_11);
DFFARX1 I_11(n_431_0_l_11,blif_clk_net_1_r_7,n8_7,n43_11,);
not I_12(n26_11,n43_11);
DFFARX1 I_13(IN_2_5_l_11,blif_clk_net_1_r_7,n8_7,n44_11,);
DFFARX1 I_14(IN_1_5_l_11,blif_clk_net_1_r_7,n8_7,n45_11,);
not I_15(n27_11,n45_11);
nor I_16(n4_1_r_11,n44_11,n25_11);
nor I_17(N3_2_r_11,n45_11,n40_11);
nand I_18(n24_11,IN_11_0_l_11,n39_11);
nand I_19(n25_11,IN_7_0_l_11,n38_11);
DFFARX1 I_20(n25_11,blif_clk_net_1_r_7,n8_7,n20_internal_11,);
not I_21(n20_11,n20_internal_11);
not I_22(n28_11,n25_11);
not I_23(n29_11,G1_0_l_11);
nand I_24(n30_11,n26_11,n31_11);
not I_25(n31_11,IN_5_0_l_11);
and I_26(n32_11,n26_11,n44_11);
and I_27(n33_11,IN_2_0_l_11,n34_11);
nor I_28(n34_11,IN_4_0_l_11,n29_11);
not I_29(n35_11,G2_0_l_11);
nand I_30(n36_11,G1_0_l_11,n31_11);
nor I_31(n37_11,IN_5_0_l_11,n29_11);
nor I_32(n38_11,G2_0_l_11,n31_11);
nor I_33(n39_11,G2_0_l_11,IN_10_0_l_11);
nor I_34(n40_11,G2_0_l_11,n41_11);
nor I_35(n41_11,IN_10_0_l_11,n42_11);
not I_36(n42_11,IN_11_0_l_11);
DFFARX1 I_37(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_38(n_572_1_r_7,n30_7,n31_7);
nand I_39(n_573_1_r_7,n28_7,G42_1_r_11);
nor I_40(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_41(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_42(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_43(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_44(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_45(P6_5_r_7,P6_5_r_internal_7);
or I_46(n_431_0_l_7,n36_7,G42_1_r_11);
not I_47(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_48(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_49(n27_7,n43_7);
DFFARX1 I_50(n_452_1_r_11,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_51(n_572_1_r_11,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_52(n4_1_r_7,n30_7,n38_7);
nor I_53(N1_4_r_7,n27_7,n40_7);
nand I_54(n26_7,n39_7,G199_2_r_11);
not I_55(n5_7,n_549_1_r_11);
DFFARX1 I_56(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_57(n28_7,n26_7,n29_7);
not I_58(n29_7,n_569_1_r_11);
not I_59(n30_7,ACVQN2_3_r_11);
nand I_60(n31_7,n27_7,n29_7);
nor I_61(n32_7,ACVQN1_5_l_7,n34_7);
nor I_62(n33_7,n29_7,n_549_1_r_11);
not I_63(n34_7,G42_1_r_11);
nor I_64(n35_7,n43_7,n44_7);
and I_65(n36_7,n37_7,n_573_1_r_11);
nor I_66(n37_7,n30_7,n_266_and_0_3_r_11);
nand I_67(n38_7,n29_7,n_549_1_r_11);
nor I_68(n39_7,n_549_1_r_11,n_42_2_r_11);
nor I_69(n40_7,n44_7,n41_7);
nor I_70(n41_7,n34_7,n42_7);
nand I_71(n42_7,n5_7,n_569_1_r_11);
endmodule


