module test_I6869(I1477,I5091,I1470,I5249,I6869);
input I1477,I5091,I1470,I5249;
output I6869;
wire I7365,I6941,I5070,I7026,I5067,I6907,I7348,I7269,I5481,I6958;
and I_0(I7365,I7026,I7348);
nor I_1(I6941,I5070);
and I_2(I5070,I5249,I5481);
not I_3(I7026,I5070);
DFFARX1 I_4(I1470,,,I5067,);
not I_5(I6907,I1477);
nand I_6(I7348,I7269,I6958);
DFFARX1 I_7(I5067,I1470,I6907,,,I7269,);
DFFARX1 I_8(I7365,I1470,I6907,,,I6869,);
DFFARX1 I_9(I1470,,,I5481,);
nand I_10(I6958,I6941,I5091);
endmodule


