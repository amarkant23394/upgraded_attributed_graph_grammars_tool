module test_I1929(I1294,I1954,I1301,I1577,I1929);
input I1294,I1954,I1301,I1577;
output I1929;
wire I2268,I1971,I2251,I1937,I1342,I2234,I2070,I1988,I1304,I1334,I1310;
and I_0(I2268,I2070,I2251);
nor I_1(I1971,I1310);
nand I_2(I2251,I2234,I1988);
not I_3(I1937,I1301);
not I_4(I1342,I1301);
nand I_5(I2234,I1954,I1304);
not I_6(I2070,I1310);
nand I_7(I1988,I1971,I1334);
DFFARX1 I_8(I1294,I1342,,,I1304,);
DFFARX1 I_9(I2268,I1294,I1937,,,I1929,);
DFFARX1 I_10(I1294,I1342,,,I1334,);
DFFARX1 I_11(I1577,I1294,I1342,,,I1310,);
endmodule


