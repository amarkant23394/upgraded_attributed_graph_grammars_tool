module Benchmark_testing1000(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1470_clk,I1477_rst,I16208,I16211,I16205,I16214,I16220,I16223,I16202,I16232,I16229,I16217,I16226,I16801,I16804,I16786,I16807,I16798,I16789,I16780,I16810,I16795,I16792,I16783,I17402,I17387,I17384,I17381,I17399,I17396,I17375,I17378,I17405,I17390,I17393);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1470_clk,I1477_rst;
output I16208,I16211,I16205,I16214,I16220,I16223,I16202,I16232,I16229,I16217,I16226,I16801,I16804,I16786,I16807,I16798,I16789,I16780,I16810,I16795,I16792,I16783,I17402,I17387,I17384,I17381,I17399,I17396,I17375,I17378,I17405,I17390,I17393;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1470_clk,I1477_rst,I1518_rst,I1535,I1552,I1569,I1586,I1603,I1620,I1637,I1507,I1668,I1492,I1699,I1716,I1733,I1750,I1767,I1784,I1801,I1489,I1832,I1849,I1486,I1880,I1897,I1504,I1928,I1501,I1959,I1976,I1480,I1483,I2021,I2038,I2055,I2072,I1510,I2103,I1495,I1498,I2181_rst,I2198,I2215,I2232,I2170,I2263,I2158,I2294,I2311,I2328,I2345,I2362,I2161,I2393,I2146,I2424,I2441,I2458,I2475,I2492,I2509,I2152,I2540,I2557,I2574,I2164,I2173,I2143,I2633,I2167,I2155,I2678,I2695,I2149,I2759_rst,I2776,I2793,I2810,I2827,I2844,I2861,I2878,I2895,I2912,I2929,I2946,I2963,I2980,I2748,I3011,I3028,I3045,I2721,I3076,I2742,I3107,I3124,I2727,I3155,I2724,I2730,I3200,I3217,I3234,I2736,I2751,I2739,I3293,I3310,I2745,I2733,I3388_rst,I3405,I3422,I3362,I3453,I3470,I3487,I3504,I3521,I3538,I3555,I3572,I3589,I3356,I3620,I3637,I3353,I3668,I3685,I3702,I3365,I3350,I3747,I3764,I3781,I3798,I3815,I3371,I3846,I3380,I3877,I3374,I3377,I3368,I3359,I3983_rst,I4000,I4017,I4034,I4051,I4068,I3966,I3954,I4113,I4130,I4147,I4164,I4181,I3963,I4212,I4229,I4246,I4263,I3972,I3951,I4308,I4325,I3969,I4356,I3960,I3975,I4401,I4418,I4435,I4452,I3948,I3957,I3945,I4544_rst,I4561,I4578,I4595,I4612,I4629,I4527,I4515,I4674,I4691,I4708,I4725,I4742,I4524,I4773,I4790,I4807,I4824,I4533,I4512,I4869,I4886,I4530,I4917,I4521,I4536,I4962,I4979,I4996,I5013,I4509,I4518,I4506,I5105_rst,I5122,I5139,I5156,I5079,I5187,I5204,I5094,I5076,I5249,I5266,I5283,I5300,I5317,I5334,I5351,I5368,I5385,I5091,I5416,I5433,I5450,I5073,I5481,I5070,I5512,I5529,I5546,I5563,I5085,I5594,I5082,I5625,I5642,I5659,I5088,I5097,I5067,I5751_rst,I5768,I5785,I5802,I5740,I5833,I5728,I5864,I5881,I5898,I5915,I5932,I5731,I5963,I5716,I5994,I6011,I6028,I6045,I6062,I6079,I5722,I6110,I6127,I6144,I5734,I5743,I5713,I6203,I5737,I5725,I6248,I6265,I5719,I6329_rst,I6346,I6363,I6380,I6318,I6411,I6306,I6442,I6459,I6476,I6493,I6510,I6309,I6541,I6294,I6572,I6589,I6606,I6623,I6640,I6657,I6300,I6688,I6705,I6722,I6312,I6321,I6291,I6781,I6315,I6303,I6826,I6843,I6297,I6907_rst,I6924,I6941,I6958,I6975,I6992,I7009,I7026,I6896,I7057,I6881,I7088,I7105,I7122,I7139,I7156,I7173,I7190,I6878,I7221,I7238,I6875,I7269,I7286,I6893,I7317,I6890,I7348,I7365,I6869,I6872,I7410,I7427,I7444,I7461,I6899,I7492,I6884,I6887,I7570_rst,I7587,I7604,I7621,I7544,I7652,I7669,I7559,I7541,I7714,I7731,I7748,I7765,I7782,I7799,I7816,I7833,I7850,I7556,I7881,I7898,I7915,I7538,I7946,I7535,I7977,I7994,I8011,I8028,I7550,I8059,I7547,I8090,I8107,I8124,I7553,I7562,I7532,I8216_rst,I8233,I8250,I8267,I8190,I8298,I8315,I8205,I8187,I8360,I8377,I8394,I8411,I8428,I8445,I8462,I8479,I8496,I8202,I8527,I8544,I8561,I8184,I8592,I8181,I8623,I8640,I8657,I8674,I8196,I8705,I8193,I8736,I8753,I8770,I8199,I8208,I8178,I8862_rst,I8879,I8896,I8913,I8930,I8947,I8964,I8981,I8998,I9015,I9032,I9049,I9066,I9083,I8851,I9114,I9131,I9148,I8824,I9179,I8845,I9210,I9227,I8830,I9258,I8827,I8833,I9303,I9320,I9337,I8839,I8854,I8842,I9396,I9413,I8848,I8836,I9491_rst,I9508,I9525,I9542,I9559,I9576,I9474,I9462,I9621,I9638,I9655,I9672,I9689,I9471,I9720,I9737,I9754,I9771,I9480,I9459,I9816,I9833,I9477,I9864,I9468,I9483,I9909,I9926,I9943,I9960,I9456,I9465,I9453,I10052_rst,I10069,I10086,I10103,I10120,I10137,I10154,I10023,I10185,I10202,I10219,I10236,I10253,I10270,I10287,I10020,I10014,I10332,I10349,I10366,I10041,I10397,I10414,I10032,I10026,I10459,I10029,I10490,I10507,I10044,I10538,I10038,I10035,I10583,I10017,I10647,I10664,I10681,I10698,I10715,I10732,I10749,I10766,I10636,I10797,I10621,I10828,I10845,I10862,I10879,I10896,I10913,I10930,I10618,I10961,I10978,I10615,I11009,I11026,I10633,I11057,I10630,I11088,I11105,I10609,I10612,I11150,I11167,I11184,I11201,I10639,I11232,I10624,I10627,I11310_rst,I11327,I11344,I11361,I11378,I11395,I11412,I11429,I11299,I11460,I11284,I11491,I11508,I11525,I11542,I11559,I11576,I11593,I11281,I11624,I11641,I11278,I11672,I11689,I11296,I11720,I11293,I11751,I11768,I11272,I11275,I11813,I11830,I11847,I11864,I11302,I11895,I11287,I11290,I11973_rst,I11990,I12007,I12024,I12041,I12058,I12075,I11944,I12106,I12123,I12140,I12157,I12174,I12191,I12208,I11941,I12239,I11935,I12270,I12287,I12304,I11965,I11938,I12349,I11962,I12380,I11959,I11956,I12425,I12442,I12459,I12476,I12493,I11950,I12524,I12541,I11953,I11947,I12619_rst,I12636,I12653,I12670,I12687,I12587,I12718,I12735,I12752,I12590,I12783,I12584,I12814,I12831,I12848,I12865,I12882,I12593,I12913,I12930,I12947,I12964,I12599,I12602,I12581,I13023,I13040,I13057,I12611,I12608,I13102,I13119,I12596,I12605,I13197_rst,I13214,I13231,I13248,I13265,I13165,I13296,I13313,I13330,I13168,I13361,I13162,I13392,I13409,I13426,I13443,I13460,I13171,I13491,I13508,I13525,I13542,I13177,I13180,I13159,I13601,I13618,I13635,I13189,I13186,I13680,I13697,I13174,I13183,I13775_rst,I13792,I13809,I13826,I13843,I13860,I13758,I13891,I13908,I13925,I13761,I13743,I13970,I13987,I14004,I13764,I13755,I14049,I14066,I14083,I13746,I14114,I14131,I13737,I14162,I14179,I14196,I13767,I14227,I14244,I14261,I14278,I13752,I13749,I13740,I14370_rst,I14387,I14404,I14421,I14438,I14455,I14472,I14341,I14503,I14520,I14537,I14554,I14571,I14588,I14605,I14338,I14332,I14650,I14667,I14684,I14359,I14715,I14732,I14350,I14344,I14777,I14347,I14808,I14825,I14362,I14856,I14356,I14353,I14901,I14335,I14965_rst,I14982,I14999,I15016,I14939,I15047,I15064,I14954,I14936,I15109,I15126,I15143,I15160,I15177,I15194,I15211,I15228,I15245,I14951,I15276,I15293,I15310,I14933,I15341,I14930,I15372,I15389,I15406,I15423,I14945,I15454,I14942,I15485,I15502,I15519,I14948,I14957,I14927,I15611_rst,I15628,I15645,I15662,I15679,I15696,I15713,I15730,I15747,I15764,I15781,I15798,I15815,I15832,I15600,I15863,I15880,I15897,I15573,I15928,I15594,I15959,I15976,I15579,I16007,I15576,I15582,I16052,I16069,I16086,I15588,I15603,I15591,I16145,I16162,I15597,I15585,I16240_rst,I16257,I16274,I16291,I16308,I16339,I16356,I16373,I16404,I16435,I16452,I16469,I16486,I16503,I16534,I16551,I16568,I16585,I16644,I16661,I16678,I16723,I16740,I16818_rst,I16835,I16852,I16869,I16886,I16903,I16934,I16951,I16968,I17013,I17030,I17047,I17092,I17109,I17126,I17157,I17174,I17205,I17222,I17239,I17270,I17287,I17304,I17321,I17413_rst,I17430,I17447,I17464,I17481,I17498,I17515,I17532,I17563,I17594,I17611,I17628,I17645,I17662,I17679,I17696,I17727,I17744,I17775,I17792,I17823,I17854,I17871,I17916,I17933,I17950,I17967,I17998;
not I_0 (I1518_rst,I1477_rst);
not I_1 (I1535,I1455);
nor I_2 (I1552,I1215,I1399);
nand I_3 (I1569,I1552,I1463);
nor I_4 (I1586,I1535,I1215);
nand I_5 (I1603,I1586,I1423);
not I_6 (I1620,I1603);
not I_7 (I1637,I1215);
nor I_8 (I1507,I1603,I1637);
not I_9 (I1668,I1637);
nand I_10 (I1492,I1603,I1668);
not I_11 (I1699,I1207);
nor I_12 (I1716,I1699,I1367);
and I_13 (I1733,I1716,I1439);
or I_14 (I1750,I1733,I1279);
DFFARX1 I_15  ( .D(I1750), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I1767) );
nor I_16 (I1784,I1767,I1620);
DFFARX1 I_17  ( .D(I1767), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I1801) );
not I_18 (I1489,I1801);
nand I_19 (I1832,I1535,I1207);
and I_20 (I1849,I1832,I1784);
DFFARX1 I_21  ( .D(I1832), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I1486) );
DFFARX1 I_22  ( .D(I1383), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I1880) );
nor I_23 (I1897,I1880,I1603);
nand I_24 (I1504,I1767,I1897);
nor I_25 (I1928,I1880,I1668);
not I_26 (I1501,I1880);
nand I_27 (I1959,I1880,I1569);
and I_28 (I1976,I1637,I1959);
DFFARX1 I_29  ( .D(I1976), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I1480) );
DFFARX1 I_30  ( .D(I1880), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I1483) );
DFFARX1 I_31  ( .D(I1295), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I2021) );
not I_32 (I2038,I2021);
nand I_33 (I2055,I2038,I1603);
and I_34 (I2072,I1832,I2055);
DFFARX1 I_35  ( .D(I2072), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I1510) );
or I_36 (I2103,I2038,I1849);
DFFARX1 I_37  ( .D(I2103), .CLK(I1470_clk), .RSTB(I1518_rst), .Q(I1495) );
nand I_38 (I1498,I2038,I1928);
not I_39 (I2181_rst,I1477_rst);
nand I_40 (I2198,I1343,I1231);
and I_41 (I2215,I2198,I1271);
DFFARX1 I_42  ( .D(I2215), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2232) );
not I_43 (I2170,I2232);
DFFARX1 I_44  ( .D(I2232), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2263) );
not I_45 (I2158,I2263);
nor I_46 (I2294,I1287,I1231);
not I_47 (I2311,I2294);
nor I_48 (I2328,I2232,I2311);
DFFARX1 I_49  ( .D(I1375), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2345) );
not I_50 (I2362,I2345);
nand I_51 (I2161,I2345,I2311);
DFFARX1 I_52  ( .D(I2345), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2393) );
and I_53 (I2146,I2232,I2393);
nand I_54 (I2424,I1223,I1255);
and I_55 (I2441,I2424,I1327);
DFFARX1 I_56  ( .D(I2441), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2458) );
nor I_57 (I2475,I2458,I2362);
and I_58 (I2492,I2294,I2475);
nor I_59 (I2509,I2458,I2232);
DFFARX1 I_60  ( .D(I2458), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2152) );
DFFARX1 I_61  ( .D(I1247), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2540) );
and I_62 (I2557,I2540,I1303);
or I_63 (I2574,I2557,I2492);
DFFARX1 I_64  ( .D(I2574), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2164) );
nand I_65 (I2173,I2557,I2509);
DFFARX1 I_66  ( .D(I2557), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2143) );
DFFARX1 I_67  ( .D(I1239), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2633) );
nand I_68 (I2167,I2633,I2328);
DFFARX1 I_69  ( .D(I2633), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2155) );
nand I_70 (I2678,I2633,I2294);
and I_71 (I2695,I2345,I2678);
DFFARX1 I_72  ( .D(I2695), .CLK(I1470_clk), .RSTB(I2181_rst), .Q(I2149) );
not I_73 (I2759_rst,I1477_rst);
not I_74 (I2776,I1407);
nor I_75 (I2793,I1351,I1319);
nand I_76 (I2810,I2793,I1335);
nor I_77 (I2827,I2776,I1351);
nand I_78 (I2844,I2827,I1359);
not I_79 (I2861,I1351);
not I_80 (I2878,I2861);
not I_81 (I2895,I1415);
nor I_82 (I2912,I2895,I1311);
and I_83 (I2929,I2912,I1391);
or I_84 (I2946,I2929,I1263);
DFFARX1 I_85  ( .D(I2946), .CLK(I1470_clk), .RSTB(I2759_rst), .Q(I2963) );
nand I_86 (I2980,I2776,I1415);
or I_87 (I2748,I2980,I2963);
not I_88 (I3011,I2980);
nor I_89 (I3028,I2963,I3011);
and I_90 (I3045,I2861,I3028);
nand I_91 (I2721,I2980,I2878);
DFFARX1 I_92  ( .D(I1447), .CLK(I1470_clk), .RSTB(I2759_rst), .Q(I3076) );
or I_93 (I2742,I3076,I2963);
nor I_94 (I3107,I3076,I2844);
nor I_95 (I3124,I3076,I2878);
nand I_96 (I2727,I2810,I3124);
or I_97 (I3155,I3076,I3045);
DFFARX1 I_98  ( .D(I3155), .CLK(I1470_clk), .RSTB(I2759_rst), .Q(I2724) );
not I_99 (I2730,I3076);
DFFARX1 I_100  ( .D(I1431), .CLK(I1470_clk), .RSTB(I2759_rst), .Q(I3200) );
not I_101 (I3217,I3200);
nor I_102 (I3234,I3217,I2810);
DFFARX1 I_103  ( .D(I3234), .CLK(I1470_clk), .RSTB(I2759_rst), .Q(I2736) );
nor I_104 (I2751,I3076,I3217);
nor I_105 (I2739,I3217,I2980);
not I_106 (I3293,I3217);
and I_107 (I3310,I2844,I3293);
nor I_108 (I2745,I2980,I3310);
nand I_109 (I2733,I3217,I3107);
not I_110 (I3388_rst,I1477_rst);
or I_111 (I3405,I1480,I1495);
or I_112 (I3422,I1483,I1480);
DFFARX1 I_113  ( .D(I3422), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3362) );
nor I_114 (I3453,I1486,I1501);
not I_115 (I3470,I3453);
not I_116 (I3487,I1486);
and I_117 (I3504,I3487,I1489);
nor I_118 (I3521,I3504,I1495);
nor I_119 (I3538,I1492,I1510);
DFFARX1 I_120  ( .D(I3538), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3555) );
nand I_121 (I3572,I3555,I3405);
and I_122 (I3589,I3521,I3572);
DFFARX1 I_123  ( .D(I3589), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3356) );
nor I_124 (I3620,I1492,I1483);
DFFARX1 I_125  ( .D(I3620), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3637) );
and I_126 (I3353,I3453,I3637);
DFFARX1 I_127  ( .D(I1507), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3668) );
and I_128 (I3685,I3668,I1498);
DFFARX1 I_129  ( .D(I3685), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3702) );
not I_130 (I3365,I3702);
DFFARX1 I_131  ( .D(I3685), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3350) );
DFFARX1 I_132  ( .D(I1504), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3747) );
not I_133 (I3764,I3747);
nor I_134 (I3781,I3422,I3764);
and I_135 (I3798,I3685,I3781);
or I_136 (I3815,I3405,I3798);
DFFARX1 I_137  ( .D(I3815), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3371) );
nor I_138 (I3846,I3747,I3555);
nand I_139 (I3380,I3521,I3846);
nor I_140 (I3877,I3747,I3470);
nand I_141 (I3374,I3620,I3877);
not I_142 (I3377,I3747);
nand I_143 (I3368,I3747,I3470);
DFFARX1 I_144  ( .D(I3747), .CLK(I1470_clk), .RSTB(I3388_rst), .Q(I3359) );
not I_145 (I3983_rst,I1477_rst);
nand I_146 (I4000,I2721,I2724);
and I_147 (I4017,I4000,I2730);
DFFARX1 I_148  ( .D(I4017), .CLK(I1470_clk), .RSTB(I3983_rst), .Q(I4034) );
not I_149 (I4051,I4034);
nor I_150 (I4068,I2742,I2724);
or I_151 (I3966,I4068,I4034);
not I_152 (I3954,I4068);
DFFARX1 I_153  ( .D(I2751), .CLK(I1470_clk), .RSTB(I3983_rst), .Q(I4113) );
nor I_154 (I4130,I4113,I4068);
nand I_155 (I4147,I2739,I2736);
and I_156 (I4164,I4147,I2748);
DFFARX1 I_157  ( .D(I4164), .CLK(I1470_clk), .RSTB(I3983_rst), .Q(I4181) );
nor I_158 (I3963,I4181,I4034);
not I_159 (I4212,I4181);
nor I_160 (I4229,I4113,I4212);
DFFARX1 I_161  ( .D(I2745), .CLK(I1470_clk), .RSTB(I3983_rst), .Q(I4246) );
and I_162 (I4263,I4246,I2733);
or I_163 (I3972,I4263,I4068);
nand I_164 (I3951,I4263,I4229);
DFFARX1 I_165  ( .D(I2727), .CLK(I1470_clk), .RSTB(I3983_rst), .Q(I4308) );
and I_166 (I4325,I4308,I4051);
nor I_167 (I3969,I4263,I4325);
nor I_168 (I4356,I4308,I4113);
DFFARX1 I_169  ( .D(I4356), .CLK(I1470_clk), .RSTB(I3983_rst), .Q(I3960) );
nor I_170 (I3975,I4308,I4034);
not I_171 (I4401,I4308);
nor I_172 (I4418,I4181,I4401);
and I_173 (I4435,I4068,I4418);
or I_174 (I4452,I4263,I4435);
DFFARX1 I_175  ( .D(I4452), .CLK(I1470_clk), .RSTB(I3983_rst), .Q(I3948) );
nand I_176 (I3957,I4308,I4130);
nand I_177 (I3945,I4308,I4212);
not I_178 (I4544_rst,I1477_rst);
nand I_179 (I4561,I2152,I2173);
and I_180 (I4578,I4561,I2161);
DFFARX1 I_181  ( .D(I4578), .CLK(I1470_clk), .RSTB(I4544_rst), .Q(I4595) );
not I_182 (I4612,I4595);
nor I_183 (I4629,I2167,I2173);
or I_184 (I4527,I4629,I4595);
not I_185 (I4515,I4629);
DFFARX1 I_186  ( .D(I2155), .CLK(I1470_clk), .RSTB(I4544_rst), .Q(I4674) );
nor I_187 (I4691,I4674,I4629);
nand I_188 (I4708,I2146,I2164);
and I_189 (I4725,I4708,I2158);
DFFARX1 I_190  ( .D(I4725), .CLK(I1470_clk), .RSTB(I4544_rst), .Q(I4742) );
nor I_191 (I4524,I4742,I4595);
not I_192 (I4773,I4742);
nor I_193 (I4790,I4674,I4773);
DFFARX1 I_194  ( .D(I2170), .CLK(I1470_clk), .RSTB(I4544_rst), .Q(I4807) );
and I_195 (I4824,I4807,I2143);
or I_196 (I4533,I4824,I4629);
nand I_197 (I4512,I4824,I4790);
DFFARX1 I_198  ( .D(I2149), .CLK(I1470_clk), .RSTB(I4544_rst), .Q(I4869) );
and I_199 (I4886,I4869,I4612);
nor I_200 (I4530,I4824,I4886);
nor I_201 (I4917,I4869,I4674);
DFFARX1 I_202  ( .D(I4917), .CLK(I1470_clk), .RSTB(I4544_rst), .Q(I4521) );
nor I_203 (I4536,I4869,I4595);
not I_204 (I4962,I4869);
nor I_205 (I4979,I4742,I4962);
and I_206 (I4996,I4629,I4979);
or I_207 (I5013,I4824,I4996);
DFFARX1 I_208  ( .D(I5013), .CLK(I1470_clk), .RSTB(I4544_rst), .Q(I4509) );
nand I_209 (I4518,I4869,I4691);
nand I_210 (I4506,I4869,I4773);
not I_211 (I5105_rst,I1477_rst);
not I_212 (I5122,I3350);
nor I_213 (I5139,I3380,I3359);
nand I_214 (I5156,I5139,I3371);
DFFARX1 I_215  ( .D(I5156), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5079) );
nor I_216 (I5187,I5122,I3380);
nand I_217 (I5204,I5187,I3353);
not I_218 (I5094,I5204);
DFFARX1 I_219  ( .D(I5204), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5076) );
not I_220 (I5249,I3380);
not I_221 (I5266,I5249);
not I_222 (I5283,I3356);
nor I_223 (I5300,I5283,I3374);
and I_224 (I5317,I5300,I3365);
or I_225 (I5334,I5317,I3362);
DFFARX1 I_226  ( .D(I5334), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5351) );
nor I_227 (I5368,I5351,I5204);
nor I_228 (I5385,I5351,I5266);
nand I_229 (I5091,I5156,I5385);
nand I_230 (I5416,I5122,I3356);
nand I_231 (I5433,I5416,I5351);
and I_232 (I5450,I5416,I5433);
DFFARX1 I_233  ( .D(I5450), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5073) );
DFFARX1 I_234  ( .D(I5416), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5481) );
and I_235 (I5070,I5249,I5481);
DFFARX1 I_236  ( .D(I3368), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5512) );
not I_237 (I5529,I5512);
nor I_238 (I5546,I5204,I5529);
and I_239 (I5563,I5512,I5546);
nand I_240 (I5085,I5512,I5266);
DFFARX1 I_241  ( .D(I5512), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5594) );
not I_242 (I5082,I5594);
DFFARX1 I_243  ( .D(I3377), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5625) );
not I_244 (I5642,I5625);
or I_245 (I5659,I5642,I5563);
DFFARX1 I_246  ( .D(I5659), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5088) );
nand I_247 (I5097,I5642,I5368);
DFFARX1 I_248  ( .D(I5642), .CLK(I1470_clk), .RSTB(I5105_rst), .Q(I5067) );
not I_249 (I5751_rst,I1477_rst);
nand I_250 (I5768,I4530,I4515);
and I_251 (I5785,I5768,I4524);
DFFARX1 I_252  ( .D(I5785), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5802) );
not I_253 (I5740,I5802);
DFFARX1 I_254  ( .D(I5802), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5833) );
not I_255 (I5728,I5833);
nor I_256 (I5864,I4536,I4515);
not I_257 (I5881,I5864);
nor I_258 (I5898,I5802,I5881);
DFFARX1 I_259  ( .D(I4527), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5915) );
not I_260 (I5932,I5915);
nand I_261 (I5731,I5915,I5881);
DFFARX1 I_262  ( .D(I5915), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5963) );
and I_263 (I5716,I5802,I5963);
nand I_264 (I5994,I4512,I4506);
and I_265 (I6011,I5994,I4521);
DFFARX1 I_266  ( .D(I6011), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I6028) );
nor I_267 (I6045,I6028,I5932);
and I_268 (I6062,I5864,I6045);
nor I_269 (I6079,I6028,I5802);
DFFARX1 I_270  ( .D(I6028), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5722) );
DFFARX1 I_271  ( .D(I4509), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I6110) );
and I_272 (I6127,I6110,I4533);
or I_273 (I6144,I6127,I6062);
DFFARX1 I_274  ( .D(I6144), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5734) );
nand I_275 (I5743,I6127,I6079);
DFFARX1 I_276  ( .D(I6127), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5713) );
DFFARX1 I_277  ( .D(I4518), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I6203) );
nand I_278 (I5737,I6203,I5898);
DFFARX1 I_279  ( .D(I6203), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5725) );
nand I_280 (I6248,I6203,I5864);
and I_281 (I6265,I5915,I6248);
DFFARX1 I_282  ( .D(I6265), .CLK(I1470_clk), .RSTB(I5751_rst), .Q(I5719) );
not I_283 (I6329_rst,I1477_rst);
nand I_284 (I6346,I3969,I3954);
and I_285 (I6363,I6346,I3963);
DFFARX1 I_286  ( .D(I6363), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6380) );
not I_287 (I6318,I6380);
DFFARX1 I_288  ( .D(I6380), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6411) );
not I_289 (I6306,I6411);
nor I_290 (I6442,I3975,I3954);
not I_291 (I6459,I6442);
nor I_292 (I6476,I6380,I6459);
DFFARX1 I_293  ( .D(I3966), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6493) );
not I_294 (I6510,I6493);
nand I_295 (I6309,I6493,I6459);
DFFARX1 I_296  ( .D(I6493), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6541) );
and I_297 (I6294,I6380,I6541);
nand I_298 (I6572,I3951,I3945);
and I_299 (I6589,I6572,I3960);
DFFARX1 I_300  ( .D(I6589), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6606) );
nor I_301 (I6623,I6606,I6510);
and I_302 (I6640,I6442,I6623);
nor I_303 (I6657,I6606,I6380);
DFFARX1 I_304  ( .D(I6606), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6300) );
DFFARX1 I_305  ( .D(I3948), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6688) );
and I_306 (I6705,I6688,I3972);
or I_307 (I6722,I6705,I6640);
DFFARX1 I_308  ( .D(I6722), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6312) );
nand I_309 (I6321,I6705,I6657);
DFFARX1 I_310  ( .D(I6705), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6291) );
DFFARX1 I_311  ( .D(I3957), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6781) );
nand I_312 (I6315,I6781,I6476);
DFFARX1 I_313  ( .D(I6781), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6303) );
nand I_314 (I6826,I6781,I6442);
and I_315 (I6843,I6493,I6826);
DFFARX1 I_316  ( .D(I6843), .CLK(I1470_clk), .RSTB(I6329_rst), .Q(I6297) );
not I_317 (I6907_rst,I1477_rst);
not I_318 (I6924,I5073);
nor I_319 (I6941,I5070,I5094);
nand I_320 (I6958,I6941,I5091);
nor I_321 (I6975,I6924,I5070);
nand I_322 (I6992,I6975,I5097);
not I_323 (I7009,I6992);
not I_324 (I7026,I5070);
nor I_325 (I6896,I6992,I7026);
not I_326 (I7057,I7026);
nand I_327 (I6881,I6992,I7057);
not I_328 (I7088,I5088);
nor I_329 (I7105,I7088,I5079);
and I_330 (I7122,I7105,I5076);
or I_331 (I7139,I7122,I5085);
DFFARX1 I_332  ( .D(I7139), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I7156) );
nor I_333 (I7173,I7156,I7009);
DFFARX1 I_334  ( .D(I7156), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I7190) );
not I_335 (I6878,I7190);
nand I_336 (I7221,I6924,I5088);
and I_337 (I7238,I7221,I7173);
DFFARX1 I_338  ( .D(I7221), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I6875) );
DFFARX1 I_339  ( .D(I5067), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I7269) );
nor I_340 (I7286,I7269,I6992);
nand I_341 (I6893,I7156,I7286);
nor I_342 (I7317,I7269,I7057);
not I_343 (I6890,I7269);
nand I_344 (I7348,I7269,I6958);
and I_345 (I7365,I7026,I7348);
DFFARX1 I_346  ( .D(I7365), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I6869) );
DFFARX1 I_347  ( .D(I7269), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I6872) );
DFFARX1 I_348  ( .D(I5082), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I7410) );
not I_349 (I7427,I7410);
nand I_350 (I7444,I7427,I6992);
and I_351 (I7461,I7221,I7444);
DFFARX1 I_352  ( .D(I7461), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I6899) );
or I_353 (I7492,I7427,I7238);
DFFARX1 I_354  ( .D(I7492), .CLK(I1470_clk), .RSTB(I6907_rst), .Q(I6884) );
nand I_355 (I6887,I7427,I7317);
not I_356 (I7570_rst,I1477_rst);
not I_357 (I7587,I6300);
nor I_358 (I7604,I6297,I6294);
nand I_359 (I7621,I7604,I6315);
DFFARX1 I_360  ( .D(I7621), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I7544) );
nor I_361 (I7652,I7587,I6297);
nand I_362 (I7669,I7652,I6318);
not I_363 (I7559,I7669);
DFFARX1 I_364  ( .D(I7669), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I7541) );
not I_365 (I7714,I6297);
not I_366 (I7731,I7714);
not I_367 (I7748,I6291);
nor I_368 (I7765,I7748,I6303);
and I_369 (I7782,I7765,I6312);
or I_370 (I7799,I7782,I6306);
DFFARX1 I_371  ( .D(I7799), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I7816) );
nor I_372 (I7833,I7816,I7669);
nor I_373 (I7850,I7816,I7731);
nand I_374 (I7556,I7621,I7850);
nand I_375 (I7881,I7587,I6291);
nand I_376 (I7898,I7881,I7816);
and I_377 (I7915,I7881,I7898);
DFFARX1 I_378  ( .D(I7915), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I7538) );
DFFARX1 I_379  ( .D(I7881), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I7946) );
and I_380 (I7535,I7714,I7946);
DFFARX1 I_381  ( .D(I6321), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I7977) );
not I_382 (I7994,I7977);
nor I_383 (I8011,I7669,I7994);
and I_384 (I8028,I7977,I8011);
nand I_385 (I7550,I7977,I7731);
DFFARX1 I_386  ( .D(I7977), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I8059) );
not I_387 (I7547,I8059);
DFFARX1 I_388  ( .D(I6309), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I8090) );
not I_389 (I8107,I8090);
or I_390 (I8124,I8107,I8028);
DFFARX1 I_391  ( .D(I8124), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I7553) );
nand I_392 (I7562,I8107,I7833);
DFFARX1 I_393  ( .D(I8107), .CLK(I1470_clk), .RSTB(I7570_rst), .Q(I7532) );
not I_394 (I8216_rst,I1477_rst);
not I_395 (I8233,I5722);
nor I_396 (I8250,I5719,I5716);
nand I_397 (I8267,I8250,I5737);
DFFARX1 I_398  ( .D(I8267), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8190) );
nor I_399 (I8298,I8233,I5719);
nand I_400 (I8315,I8298,I5740);
not I_401 (I8205,I8315);
DFFARX1 I_402  ( .D(I8315), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8187) );
not I_403 (I8360,I5719);
not I_404 (I8377,I8360);
not I_405 (I8394,I5713);
nor I_406 (I8411,I8394,I5725);
and I_407 (I8428,I8411,I5734);
or I_408 (I8445,I8428,I5728);
DFFARX1 I_409  ( .D(I8445), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8462) );
nor I_410 (I8479,I8462,I8315);
nor I_411 (I8496,I8462,I8377);
nand I_412 (I8202,I8267,I8496);
nand I_413 (I8527,I8233,I5713);
nand I_414 (I8544,I8527,I8462);
and I_415 (I8561,I8527,I8544);
DFFARX1 I_416  ( .D(I8561), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8184) );
DFFARX1 I_417  ( .D(I8527), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8592) );
and I_418 (I8181,I8360,I8592);
DFFARX1 I_419  ( .D(I5743), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8623) );
not I_420 (I8640,I8623);
nor I_421 (I8657,I8315,I8640);
and I_422 (I8674,I8623,I8657);
nand I_423 (I8196,I8623,I8377);
DFFARX1 I_424  ( .D(I8623), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8705) );
not I_425 (I8193,I8705);
DFFARX1 I_426  ( .D(I5731), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8736) );
not I_427 (I8753,I8736);
or I_428 (I8770,I8753,I8674);
DFFARX1 I_429  ( .D(I8770), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8199) );
nand I_430 (I8208,I8753,I8479);
DFFARX1 I_431  ( .D(I8753), .CLK(I1470_clk), .RSTB(I8216_rst), .Q(I8178) );
not I_432 (I8862_rst,I1477_rst);
not I_433 (I8879,I6887);
nor I_434 (I8896,I6893,I6872);
nand I_435 (I8913,I8896,I6878);
nor I_436 (I8930,I8879,I6893);
nand I_437 (I8947,I8930,I6884);
not I_438 (I8964,I6893);
not I_439 (I8981,I8964);
not I_440 (I8998,I6881);
nor I_441 (I9015,I8998,I6899);
and I_442 (I9032,I9015,I6890);
or I_443 (I9049,I9032,I6869);
DFFARX1 I_444  ( .D(I9049), .CLK(I1470_clk), .RSTB(I8862_rst), .Q(I9066) );
nand I_445 (I9083,I8879,I6881);
or I_446 (I8851,I9083,I9066);
not I_447 (I9114,I9083);
nor I_448 (I9131,I9066,I9114);
and I_449 (I9148,I8964,I9131);
nand I_450 (I8824,I9083,I8981);
DFFARX1 I_451  ( .D(I6896), .CLK(I1470_clk), .RSTB(I8862_rst), .Q(I9179) );
or I_452 (I8845,I9179,I9066);
nor I_453 (I9210,I9179,I8947);
nor I_454 (I9227,I9179,I8981);
nand I_455 (I8830,I8913,I9227);
or I_456 (I9258,I9179,I9148);
DFFARX1 I_457  ( .D(I9258), .CLK(I1470_clk), .RSTB(I8862_rst), .Q(I8827) );
not I_458 (I8833,I9179);
DFFARX1 I_459  ( .D(I6875), .CLK(I1470_clk), .RSTB(I8862_rst), .Q(I9303) );
not I_460 (I9320,I9303);
nor I_461 (I9337,I9320,I8913);
DFFARX1 I_462  ( .D(I9337), .CLK(I1470_clk), .RSTB(I8862_rst), .Q(I8839) );
nor I_463 (I8854,I9179,I9320);
nor I_464 (I8842,I9320,I9083);
not I_465 (I9396,I9320);
and I_466 (I9413,I8947,I9396);
nor I_467 (I8848,I9083,I9413);
nand I_468 (I8836,I9320,I9210);
not I_469 (I9491_rst,I1477_rst);
nand I_470 (I9508,I8199,I8202);
and I_471 (I9525,I9508,I8184);
DFFARX1 I_472  ( .D(I9525), .CLK(I1470_clk), .RSTB(I9491_rst), .Q(I9542) );
not I_473 (I9559,I9542);
nor I_474 (I9576,I8181,I8202);
or I_475 (I9474,I9576,I9542);
not I_476 (I9462,I9576);
DFFARX1 I_477  ( .D(I8205), .CLK(I1470_clk), .RSTB(I9491_rst), .Q(I9621) );
nor I_478 (I9638,I9621,I9576);
nand I_479 (I9655,I8190,I8196);
and I_480 (I9672,I9655,I8208);
DFFARX1 I_481  ( .D(I9672), .CLK(I1470_clk), .RSTB(I9491_rst), .Q(I9689) );
nor I_482 (I9471,I9689,I9542);
not I_483 (I9720,I9689);
nor I_484 (I9737,I9621,I9720);
DFFARX1 I_485  ( .D(I8187), .CLK(I1470_clk), .RSTB(I9491_rst), .Q(I9754) );
and I_486 (I9771,I9754,I8178);
or I_487 (I9480,I9771,I9576);
nand I_488 (I9459,I9771,I9737);
DFFARX1 I_489  ( .D(I8193), .CLK(I1470_clk), .RSTB(I9491_rst), .Q(I9816) );
and I_490 (I9833,I9816,I9559);
nor I_491 (I9477,I9771,I9833);
nor I_492 (I9864,I9816,I9621);
DFFARX1 I_493  ( .D(I9864), .CLK(I1470_clk), .RSTB(I9491_rst), .Q(I9468) );
nor I_494 (I9483,I9816,I9542);
not I_495 (I9909,I9816);
nor I_496 (I9926,I9689,I9909);
and I_497 (I9943,I9576,I9926);
or I_498 (I9960,I9771,I9943);
DFFARX1 I_499  ( .D(I9960), .CLK(I1470_clk), .RSTB(I9491_rst), .Q(I9456) );
nand I_500 (I9465,I9816,I9638);
nand I_501 (I9453,I9816,I9720);
not I_502 (I10052_rst,I1477_rst);
nand I_503 (I10069,I7559,I7535);
and I_504 (I10086,I10069,I7544);
DFFARX1 I_505  ( .D(I10086), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10103) );
nor I_506 (I10120,I7538,I7535);
DFFARX1 I_507  ( .D(I7553), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10137) );
nand I_508 (I10154,I10137,I10120);
DFFARX1 I_509  ( .D(I10137), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10023) );
nand I_510 (I10185,I7547,I7562);
and I_511 (I10202,I10185,I7541);
DFFARX1 I_512  ( .D(I10202), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10219) );
not I_513 (I10236,I10219);
nor I_514 (I10253,I10103,I10236);
and I_515 (I10270,I10120,I10253);
and I_516 (I10287,I10219,I10154);
DFFARX1 I_517  ( .D(I10287), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10020) );
DFFARX1 I_518  ( .D(I10219), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10014) );
DFFARX1 I_519  ( .D(I7532), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10332) );
and I_520 (I10349,I10332,I7550);
nand I_521 (I10366,I10349,I10219);
nor I_522 (I10041,I10349,I10120);
not I_523 (I10397,I10349);
nor I_524 (I10414,I10103,I10397);
nand I_525 (I10032,I10137,I10414);
nand I_526 (I10026,I10219,I10397);
or I_527 (I10459,I10349,I10270);
DFFARX1 I_528  ( .D(I10459), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10029) );
DFFARX1 I_529  ( .D(I7556), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10490) );
and I_530 (I10507,I10490,I10366);
DFFARX1 I_531  ( .D(I10507), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10044) );
nor I_532 (I10538,I10490,I10103);
nand I_533 (I10038,I10349,I10538);
not I_534 (I10035,I10490);
DFFARX1 I_535  ( .D(I10490), .CLK(I1470_clk), .RSTB(I10052_rst), .Q(I10583) );
and I_536 (I10017,I10490,I10583);
not I_537 (I10647,I1477_rst);
not I_538 (I10664,I9471);
nor I_539 (I10681,I9477,I9480);
nand I_540 (I10698,I10681,I9456);
nor I_541 (I10715,I10664,I9477);
nand I_542 (I10732,I10715,I9465);
not I_543 (I10749,I10732);
not I_544 (I10766,I9477);
nor I_545 (I10636,I10732,I10766);
not I_546 (I10797,I10766);
nand I_547 (I10621,I10732,I10797);
not I_548 (I10828,I9459);
nor I_549 (I10845,I10828,I9483);
and I_550 (I10862,I10845,I9453);
or I_551 (I10879,I10862,I9462);
DFFARX1 I_552  ( .D(I10879), .CLK(I1470_clk), .RSTB(I10647), .Q(I10896) );
nor I_553 (I10913,I10896,I10749);
DFFARX1 I_554  ( .D(I10896), .CLK(I1470_clk), .RSTB(I10647), .Q(I10930) );
not I_555 (I10618,I10930);
nand I_556 (I10961,I10664,I9459);
and I_557 (I10978,I10961,I10913);
DFFARX1 I_558  ( .D(I10961), .CLK(I1470_clk), .RSTB(I10647), .Q(I10615) );
DFFARX1 I_559  ( .D(I9468), .CLK(I1470_clk), .RSTB(I10647), .Q(I11009) );
nor I_560 (I11026,I11009,I10732);
nand I_561 (I10633,I10896,I11026);
nor I_562 (I11057,I11009,I10797);
not I_563 (I10630,I11009);
nand I_564 (I11088,I11009,I10698);
and I_565 (I11105,I10766,I11088);
DFFARX1 I_566  ( .D(I11105), .CLK(I1470_clk), .RSTB(I10647), .Q(I10609) );
DFFARX1 I_567  ( .D(I11009), .CLK(I1470_clk), .RSTB(I10647), .Q(I10612) );
DFFARX1 I_568  ( .D(I9474), .CLK(I1470_clk), .RSTB(I10647), .Q(I11150) );
not I_569 (I11167,I11150);
nand I_570 (I11184,I11167,I10732);
and I_571 (I11201,I10961,I11184);
DFFARX1 I_572  ( .D(I11201), .CLK(I1470_clk), .RSTB(I10647), .Q(I10639) );
or I_573 (I11232,I11167,I10978);
DFFARX1 I_574  ( .D(I11232), .CLK(I1470_clk), .RSTB(I10647), .Q(I10624) );
nand I_575 (I10627,I11167,I11057);
not I_576 (I11310_rst,I1477_rst);
not I_577 (I11327,I8830);
nor I_578 (I11344,I8848,I8839);
nand I_579 (I11361,I11344,I8845);
nor I_580 (I11378,I11327,I8848);
nand I_581 (I11395,I11378,I8851);
not I_582 (I11412,I11395);
not I_583 (I11429,I8848);
nor I_584 (I11299,I11395,I11429);
not I_585 (I11460,I11429);
nand I_586 (I11284,I11395,I11460);
not I_587 (I11491,I8827);
nor I_588 (I11508,I11491,I8842);
and I_589 (I11525,I11508,I8824);
or I_590 (I11542,I11525,I8833);
DFFARX1 I_591  ( .D(I11542), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11559) );
nor I_592 (I11576,I11559,I11412);
DFFARX1 I_593  ( .D(I11559), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11593) );
not I_594 (I11281,I11593);
nand I_595 (I11624,I11327,I8827);
and I_596 (I11641,I11624,I11576);
DFFARX1 I_597  ( .D(I11624), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11278) );
DFFARX1 I_598  ( .D(I8836), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11672) );
nor I_599 (I11689,I11672,I11395);
nand I_600 (I11296,I11559,I11689);
nor I_601 (I11720,I11672,I11460);
not I_602 (I11293,I11672);
nand I_603 (I11751,I11672,I11361);
and I_604 (I11768,I11429,I11751);
DFFARX1 I_605  ( .D(I11768), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11272) );
DFFARX1 I_606  ( .D(I11672), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11275) );
DFFARX1 I_607  ( .D(I8854), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11813) );
not I_608 (I11830,I11813);
nand I_609 (I11847,I11830,I11395);
and I_610 (I11864,I11624,I11847);
DFFARX1 I_611  ( .D(I11864), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11302) );
or I_612 (I11895,I11830,I11641);
DFFARX1 I_613  ( .D(I11895), .CLK(I1470_clk), .RSTB(I11310_rst), .Q(I11287) );
nand I_614 (I11290,I11830,I11720);
not I_615 (I11973_rst,I1477_rst);
not I_616 (I11990,I10032);
nor I_617 (I12007,I10020,I10029);
nand I_618 (I12024,I12007,I10044);
nor I_619 (I12041,I11990,I10020);
nand I_620 (I12058,I12041,I10026);
DFFARX1 I_621  ( .D(I12058), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I12075) );
not I_622 (I11944,I12075);
not I_623 (I12106,I10020);
not I_624 (I12123,I12106);
not I_625 (I12140,I10014);
nor I_626 (I12157,I12140,I10035);
and I_627 (I12174,I12157,I10017);
or I_628 (I12191,I12174,I10023);
DFFARX1 I_629  ( .D(I12191), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I12208) );
DFFARX1 I_630  ( .D(I12208), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I11941) );
DFFARX1 I_631  ( .D(I12208), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I12239) );
DFFARX1 I_632  ( .D(I12208), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I11935) );
nand I_633 (I12270,I11990,I10014);
nand I_634 (I12287,I12270,I12024);
and I_635 (I12304,I12106,I12287);
DFFARX1 I_636  ( .D(I12304), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I11965) );
and I_637 (I11938,I12270,I12239);
DFFARX1 I_638  ( .D(I10041), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I12349) );
nor I_639 (I11962,I12349,I12270);
nor I_640 (I12380,I12349,I12024);
nand I_641 (I11959,I12058,I12380);
not I_642 (I11956,I12349);
DFFARX1 I_643  ( .D(I10038), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I12425) );
not I_644 (I12442,I12425);
nor I_645 (I12459,I12442,I12123);
and I_646 (I12476,I12349,I12459);
or I_647 (I12493,I12270,I12476);
DFFARX1 I_648  ( .D(I12493), .CLK(I1470_clk), .RSTB(I11973_rst), .Q(I11950) );
not I_649 (I12524,I12442);
nor I_650 (I12541,I12349,I12524);
nand I_651 (I11953,I12442,I12541);
nand I_652 (I11947,I12106,I12524);
not I_653 (I12619_rst,I1477_rst);
nand I_654 (I12636,I10612,I10639);
and I_655 (I12653,I12636,I10627);
DFFARX1 I_656  ( .D(I12653), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12670) );
not I_657 (I12687,I12670);
DFFARX1 I_658  ( .D(I12670), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12587) );
nor I_659 (I12718,I10615,I10639);
DFFARX1 I_660  ( .D(I10630), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12735) );
DFFARX1 I_661  ( .D(I12735), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12752) );
not I_662 (I12590,I12752);
DFFARX1 I_663  ( .D(I12735), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12783) );
and I_664 (I12584,I12670,I12783);
nand I_665 (I12814,I10624,I10621);
and I_666 (I12831,I12814,I10618);
DFFARX1 I_667  ( .D(I12831), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12848) );
nor I_668 (I12865,I12848,I12687);
not I_669 (I12882,I12848);
nand I_670 (I12593,I12670,I12882);
DFFARX1 I_671  ( .D(I10633), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12913) );
and I_672 (I12930,I12913,I10609);
nor I_673 (I12947,I12930,I12848);
nor I_674 (I12964,I12930,I12882);
nand I_675 (I12599,I12718,I12964);
not I_676 (I12602,I12930);
DFFARX1 I_677  ( .D(I12930), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12581) );
DFFARX1 I_678  ( .D(I10636), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I13023) );
nand I_679 (I13040,I13023,I12735);
and I_680 (I13057,I12718,I13040);
DFFARX1 I_681  ( .D(I13057), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12611) );
nor I_682 (I12608,I13023,I12930);
and I_683 (I13102,I13023,I12865);
or I_684 (I13119,I12718,I13102);
DFFARX1 I_685  ( .D(I13119), .CLK(I1470_clk), .RSTB(I12619_rst), .Q(I12596) );
nand I_686 (I12605,I13023,I12947);
not I_687 (I13197_rst,I1477_rst);
nand I_688 (I13214,I11275,I11302);
and I_689 (I13231,I13214,I11290);
DFFARX1 I_690  ( .D(I13231), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13248) );
not I_691 (I13265,I13248);
DFFARX1 I_692  ( .D(I13248), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13165) );
nor I_693 (I13296,I11278,I11302);
DFFARX1 I_694  ( .D(I11293), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13313) );
DFFARX1 I_695  ( .D(I13313), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13330) );
not I_696 (I13168,I13330);
DFFARX1 I_697  ( .D(I13313), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13361) );
and I_698 (I13162,I13248,I13361);
nand I_699 (I13392,I11287,I11284);
and I_700 (I13409,I13392,I11281);
DFFARX1 I_701  ( .D(I13409), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13426) );
nor I_702 (I13443,I13426,I13265);
not I_703 (I13460,I13426);
nand I_704 (I13171,I13248,I13460);
DFFARX1 I_705  ( .D(I11296), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13491) );
and I_706 (I13508,I13491,I11272);
nor I_707 (I13525,I13508,I13426);
nor I_708 (I13542,I13508,I13460);
nand I_709 (I13177,I13296,I13542);
not I_710 (I13180,I13508);
DFFARX1 I_711  ( .D(I13508), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13159) );
DFFARX1 I_712  ( .D(I11299), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13601) );
nand I_713 (I13618,I13601,I13313);
and I_714 (I13635,I13296,I13618);
DFFARX1 I_715  ( .D(I13635), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13189) );
nor I_716 (I13186,I13601,I13508);
and I_717 (I13680,I13601,I13443);
or I_718 (I13697,I13296,I13680);
DFFARX1 I_719  ( .D(I13697), .CLK(I1470_clk), .RSTB(I13197_rst), .Q(I13174) );
nand I_720 (I13183,I13601,I13525);
not I_721 (I13775_rst,I1477_rst);
nand I_722 (I13792,I11953,I11965);
and I_723 (I13809,I13792,I11947);
DFFARX1 I_724  ( .D(I13809), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I13826) );
nor I_725 (I13843,I11959,I11965);
nor I_726 (I13860,I13843,I13826);
not I_727 (I13758,I13843);
DFFARX1 I_728  ( .D(I11944), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I13891) );
not I_729 (I13908,I13891);
nor I_730 (I13925,I13843,I13908);
nand I_731 (I13761,I13891,I13860);
DFFARX1 I_732  ( .D(I13891), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I13743) );
nand I_733 (I13970,I11935,I11950);
and I_734 (I13987,I13970,I11941);
DFFARX1 I_735  ( .D(I13987), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I14004) );
nor I_736 (I13764,I14004,I13826);
nand I_737 (I13755,I14004,I13925);
DFFARX1 I_738  ( .D(I11962), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I14049) );
and I_739 (I14066,I14049,I11956);
DFFARX1 I_740  ( .D(I14066), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I14083) );
not I_741 (I13746,I14083);
nand I_742 (I14114,I14066,I14004);
and I_743 (I14131,I13826,I14114);
DFFARX1 I_744  ( .D(I14131), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I13737) );
DFFARX1 I_745  ( .D(I11938), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I14162) );
nand I_746 (I14179,I14162,I13826);
and I_747 (I14196,I14004,I14179);
DFFARX1 I_748  ( .D(I14196), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I13767) );
not I_749 (I14227,I14162);
nor I_750 (I14244,I13843,I14227);
and I_751 (I14261,I14162,I14244);
or I_752 (I14278,I14066,I14261);
DFFARX1 I_753  ( .D(I14278), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I13752) );
nand I_754 (I13749,I14162,I13908);
DFFARX1 I_755  ( .D(I14162), .CLK(I1470_clk), .RSTB(I13775_rst), .Q(I13740) );
not I_756 (I14370_rst,I1477_rst);
nand I_757 (I14387,I13171,I13186);
and I_758 (I14404,I14387,I13183);
DFFARX1 I_759  ( .D(I14404), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14421) );
nor I_760 (I14438,I13159,I13186);
DFFARX1 I_761  ( .D(I13177), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14455) );
nand I_762 (I14472,I14455,I14438);
DFFARX1 I_763  ( .D(I14455), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14341) );
nand I_764 (I14503,I13180,I13168);
and I_765 (I14520,I14503,I13174);
DFFARX1 I_766  ( .D(I14520), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14537) );
not I_767 (I14554,I14537);
nor I_768 (I14571,I14421,I14554);
and I_769 (I14588,I14438,I14571);
and I_770 (I14605,I14537,I14472);
DFFARX1 I_771  ( .D(I14605), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14338) );
DFFARX1 I_772  ( .D(I14537), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14332) );
DFFARX1 I_773  ( .D(I13165), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14650) );
and I_774 (I14667,I14650,I13189);
nand I_775 (I14684,I14667,I14537);
nor I_776 (I14359,I14667,I14438);
not I_777 (I14715,I14667);
nor I_778 (I14732,I14421,I14715);
nand I_779 (I14350,I14455,I14732);
nand I_780 (I14344,I14537,I14715);
or I_781 (I14777,I14667,I14588);
DFFARX1 I_782  ( .D(I14777), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14347) );
DFFARX1 I_783  ( .D(I13162), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14808) );
and I_784 (I14825,I14808,I14684);
DFFARX1 I_785  ( .D(I14825), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14362) );
nor I_786 (I14856,I14808,I14421);
nand I_787 (I14356,I14667,I14856);
not I_788 (I14353,I14808);
DFFARX1 I_789  ( .D(I14808), .CLK(I1470_clk), .RSTB(I14370_rst), .Q(I14901) );
and I_790 (I14335,I14808,I14901);
not I_791 (I14965_rst,I1477_rst);
not I_792 (I14982,I12596);
nor I_793 (I14999,I12584,I12590);
nand I_794 (I15016,I14999,I12581);
DFFARX1 I_795  ( .D(I15016), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I14939) );
nor I_796 (I15047,I14982,I12584);
nand I_797 (I15064,I15047,I12587);
not I_798 (I14954,I15064);
DFFARX1 I_799  ( .D(I15064), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I14936) );
not I_800 (I15109,I12584);
not I_801 (I15126,I15109);
not I_802 (I15143,I12599);
nor I_803 (I15160,I15143,I12611);
and I_804 (I15177,I15160,I12593);
or I_805 (I15194,I15177,I12608);
DFFARX1 I_806  ( .D(I15194), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I15211) );
nor I_807 (I15228,I15211,I15064);
nor I_808 (I15245,I15211,I15126);
nand I_809 (I14951,I15016,I15245);
nand I_810 (I15276,I14982,I12599);
nand I_811 (I15293,I15276,I15211);
and I_812 (I15310,I15276,I15293);
DFFARX1 I_813  ( .D(I15310), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I14933) );
DFFARX1 I_814  ( .D(I15276), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I15341) );
and I_815 (I14930,I15109,I15341);
DFFARX1 I_816  ( .D(I12602), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I15372) );
not I_817 (I15389,I15372);
nor I_818 (I15406,I15064,I15389);
and I_819 (I15423,I15372,I15406);
nand I_820 (I14945,I15372,I15126);
DFFARX1 I_821  ( .D(I15372), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I15454) );
not I_822 (I14942,I15454);
DFFARX1 I_823  ( .D(I12605), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I15485) );
not I_824 (I15502,I15485);
or I_825 (I15519,I15502,I15423);
DFFARX1 I_826  ( .D(I15519), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I14948) );
nand I_827 (I14957,I15502,I15228);
DFFARX1 I_828  ( .D(I15502), .CLK(I1470_clk), .RSTB(I14965_rst), .Q(I14927) );
not I_829 (I15611_rst,I1477_rst);
not I_830 (I15628,I13743);
nor I_831 (I15645,I13761,I13740);
nand I_832 (I15662,I15645,I13764);
nor I_833 (I15679,I15628,I13761);
nand I_834 (I15696,I15679,I13758);
not I_835 (I15713,I13761);
not I_836 (I15730,I15713);
not I_837 (I15747,I13749);
nor I_838 (I15764,I15747,I13737);
and I_839 (I15781,I15764,I13755);
or I_840 (I15798,I15781,I13767);
DFFARX1 I_841  ( .D(I15798), .CLK(I1470_clk), .RSTB(I15611_rst), .Q(I15815) );
nand I_842 (I15832,I15628,I13749);
or I_843 (I15600,I15832,I15815);
not I_844 (I15863,I15832);
nor I_845 (I15880,I15815,I15863);
and I_846 (I15897,I15713,I15880);
nand I_847 (I15573,I15832,I15730);
DFFARX1 I_848  ( .D(I13746), .CLK(I1470_clk), .RSTB(I15611_rst), .Q(I15928) );
or I_849 (I15594,I15928,I15815);
nor I_850 (I15959,I15928,I15696);
nor I_851 (I15976,I15928,I15730);
nand I_852 (I15579,I15662,I15976);
or I_853 (I16007,I15928,I15897);
DFFARX1 I_854  ( .D(I16007), .CLK(I1470_clk), .RSTB(I15611_rst), .Q(I15576) );
not I_855 (I15582,I15928);
DFFARX1 I_856  ( .D(I13752), .CLK(I1470_clk), .RSTB(I15611_rst), .Q(I16052) );
not I_857 (I16069,I16052);
nor I_858 (I16086,I16069,I15662);
DFFARX1 I_859  ( .D(I16086), .CLK(I1470_clk), .RSTB(I15611_rst), .Q(I15588) );
nor I_860 (I15603,I15928,I16069);
nor I_861 (I15591,I16069,I15832);
not I_862 (I16145,I16069);
and I_863 (I16162,I15696,I16145);
nor I_864 (I15597,I15832,I16162);
nand I_865 (I15585,I16069,I15959);
not I_866 (I16240_rst,I1477_rst);
nand I_867 (I16257,I14341,I14338);
and I_868 (I16274,I16257,I14332);
DFFARX1 I_869  ( .D(I16274), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16291) );
not I_870 (I16308,I16291);
DFFARX1 I_871  ( .D(I16291), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16208) );
nor I_872 (I16339,I14353,I14338);
DFFARX1 I_873  ( .D(I14356), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16356) );
DFFARX1 I_874  ( .D(I16356), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16373) );
not I_875 (I16211,I16373);
DFFARX1 I_876  ( .D(I16356), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16404) );
and I_877 (I16205,I16291,I16404);
nand I_878 (I16435,I14359,I14350);
and I_879 (I16452,I16435,I14362);
DFFARX1 I_880  ( .D(I16452), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16469) );
nor I_881 (I16486,I16469,I16308);
not I_882 (I16503,I16469);
nand I_883 (I16214,I16291,I16503);
DFFARX1 I_884  ( .D(I14335), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16534) );
and I_885 (I16551,I16534,I14344);
nor I_886 (I16568,I16551,I16469);
nor I_887 (I16585,I16551,I16503);
nand I_888 (I16220,I16339,I16585);
not I_889 (I16223,I16551);
DFFARX1 I_890  ( .D(I16551), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16202) );
DFFARX1 I_891  ( .D(I14347), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16644) );
nand I_892 (I16661,I16644,I16356);
and I_893 (I16678,I16339,I16661);
DFFARX1 I_894  ( .D(I16678), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16232) );
nor I_895 (I16229,I16644,I16551);
and I_896 (I16723,I16644,I16486);
or I_897 (I16740,I16339,I16723);
DFFARX1 I_898  ( .D(I16740), .CLK(I1470_clk), .RSTB(I16240_rst), .Q(I16217) );
nand I_899 (I16226,I16644,I16568);
not I_900 (I16818_rst,I1477_rst);
nand I_901 (I16835,I14936,I14948);
and I_902 (I16852,I16835,I14957);
DFFARX1 I_903  ( .D(I16852), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I16869) );
nor I_904 (I16886,I14951,I14948);
nor I_905 (I16903,I16886,I16869);
not I_906 (I16801,I16886);
DFFARX1 I_907  ( .D(I14945), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I16934) );
not I_908 (I16951,I16934);
nor I_909 (I16968,I16886,I16951);
nand I_910 (I16804,I16934,I16903);
DFFARX1 I_911  ( .D(I16934), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I16786) );
nand I_912 (I17013,I14942,I14939);
and I_913 (I17030,I17013,I14930);
DFFARX1 I_914  ( .D(I17030), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I17047) );
nor I_915 (I16807,I17047,I16869);
nand I_916 (I16798,I17047,I16968);
DFFARX1 I_917  ( .D(I14954), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I17092) );
and I_918 (I17109,I17092,I14933);
DFFARX1 I_919  ( .D(I17109), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I17126) );
not I_920 (I16789,I17126);
nand I_921 (I17157,I17109,I17047);
and I_922 (I17174,I16869,I17157);
DFFARX1 I_923  ( .D(I17174), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I16780) );
DFFARX1 I_924  ( .D(I14927), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I17205) );
nand I_925 (I17222,I17205,I16869);
and I_926 (I17239,I17047,I17222);
DFFARX1 I_927  ( .D(I17239), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I16810) );
not I_928 (I17270,I17205);
nor I_929 (I17287,I16886,I17270);
and I_930 (I17304,I17205,I17287);
or I_931 (I17321,I17109,I17304);
DFFARX1 I_932  ( .D(I17321), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I16795) );
nand I_933 (I16792,I17205,I16951);
DFFARX1 I_934  ( .D(I17205), .CLK(I1470_clk), .RSTB(I16818_rst), .Q(I16783) );
not I_935 (I17413_rst,I1477_rst);
not I_936 (I17430,I15579);
nor I_937 (I17447,I15597,I15588);
nand I_938 (I17464,I17447,I15594);
nor I_939 (I17481,I17430,I15597);
nand I_940 (I17498,I17481,I15600);
not I_941 (I17515,I17498);
not I_942 (I17532,I15597);
nor I_943 (I17402,I17498,I17532);
not I_944 (I17563,I17532);
nand I_945 (I17387,I17498,I17563);
not I_946 (I17594,I15576);
nor I_947 (I17611,I17594,I15591);
and I_948 (I17628,I17611,I15573);
or I_949 (I17645,I17628,I15582);
DFFARX1 I_950  ( .D(I17645), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17662) );
nor I_951 (I17679,I17662,I17515);
DFFARX1 I_952  ( .D(I17662), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17696) );
not I_953 (I17384,I17696);
nand I_954 (I17727,I17430,I15576);
and I_955 (I17744,I17727,I17679);
DFFARX1 I_956  ( .D(I17727), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17381) );
DFFARX1 I_957  ( .D(I15585), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17775) );
nor I_958 (I17792,I17775,I17498);
nand I_959 (I17399,I17662,I17792);
nor I_960 (I17823,I17775,I17563);
not I_961 (I17396,I17775);
nand I_962 (I17854,I17775,I17464);
and I_963 (I17871,I17532,I17854);
DFFARX1 I_964  ( .D(I17871), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17375) );
DFFARX1 I_965  ( .D(I17775), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17378) );
DFFARX1 I_966  ( .D(I15603), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17916) );
not I_967 (I17933,I17916);
nand I_968 (I17950,I17933,I17498);
and I_969 (I17967,I17727,I17950);
DFFARX1 I_970  ( .D(I17967), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17405) );
or I_971 (I17998,I17933,I17744);
DFFARX1 I_972  ( .D(I17998), .CLK(I1470_clk), .RSTB(I17413_rst), .Q(I17390) );
nand I_973 (I17393,I17933,I17823);
endmodule


