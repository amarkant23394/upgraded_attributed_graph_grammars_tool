module test_I11395(I9032,I1477,I6887,I8913,I9396,I6992,I7057,I8947,I1470,I9227,I11395);
input I9032,I1477,I6887,I8913,I9396,I6992,I7057,I8947,I1470,I9227;
output I11395;
wire I8830,I9049,I8862,I6881,I8848,I9083,I9413,I11378,I9066,I8879,I11327,I8851,I6869;
nand I_0(I8830,I8913,I9227);
nand I_1(I11395,I11378,I8851);
or I_2(I9049,I9032,I6869);
not I_3(I8862,I1477);
nand I_4(I6881,I6992,I7057);
nor I_5(I8848,I9083,I9413);
nand I_6(I9083,I8879,I6881);
and I_7(I9413,I8947,I9396);
nor I_8(I11378,I11327,I8848);
DFFARX1 I_9(I9049,I1470,I8862,,,I9066,);
not I_10(I8879,I6887);
not I_11(I11327,I8830);
or I_12(I8851,I9083,I9066);
DFFARX1 I_13(I1470,,,I6869,);
endmodule


