module test_I3368(I1750,I1477,I1603,I1470,I1832,I3368);
input I1750,I1477,I1603,I1470,I1832;
output I3368;
wire I1518,I3388,I1486,I1504,I3470,I1880,I1501,I3453,I3747,I1897,I1767;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
DFFARX1 I_2(I1832,I1470,I1518,,,I1486,);
nand I_3(I1504,I1767,I1897);
nand I_4(I3368,I3747,I3470);
not I_5(I3470,I3453);
DFFARX1 I_6(I1470,I1518,,,I1880,);
not I_7(I1501,I1880);
nor I_8(I3453,I1486,I1501);
DFFARX1 I_9(I1504,I1470,I3388,,,I3747,);
nor I_10(I1897,I1880,I1603);
DFFARX1 I_11(I1750,I1470,I1518,,,I1767,);
endmodule


