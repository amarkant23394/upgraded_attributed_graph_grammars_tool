module test_I1444(I1223,I1263,I1294,I1239,I1301,I1444);
input I1223,I1263,I1294,I1239,I1301;
output I1444;
wire I1410,I1342,I1427;
nand I_0(I1444,I1427,I1410);
nor I_1(I1410,I1223,I1239);
not I_2(I1342,I1301);
DFFARX1 I_3(I1263,I1294,I1342,,,I1427,);
endmodule


