module test_final(IN_1_0_l,IN_2_0_l,IN_3_0_l,IN_4_0_l,IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,blif_clk_net_5_r,blif_reset_net_5_r,N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N1372_4_r,N1508_4_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,N1507_6_r,N1508_6_r);
input IN_1_0_l,IN_2_0_l,IN_3_0_l,IN_4_0_l,IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,blif_clk_net_5_r,blif_reset_net_5_r;
output N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N1372_4_r,N1508_4_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,N1507_6_r,N1508_6_r;
wire N1371_0_l,N1508_0_l,n3_0_l,n4_0_l,N1372_1_l,N1508_1_l,n4_1_l,N6147_3_l,n3_3_l,N6138_3_l,N1507_6_l,N1508_6_l,n6_6_l,n7_6_l,n8_6_l,n9_6_l,n3_0_r,n4_0_r,n4_1_r,n6_4_r,n7_4_r,n8_4_r,n_431_5_r,n2_5_r,n11_5_r,n12_5_r,n13_5_r,n14_5_r,n15_5_r,n16_5_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r;
nor I_0(N1371_0_l,IN_2_0_l,n4_0_l);
nor I_1(N1508_0_l,n3_0_l,n4_0_l);
nor I_2(n3_0_l,IN_3_0_l,IN_4_0_l);
not I_3(n4_0_l,IN_1_0_l);
not I_4(N1372_1_l,n4_1_l);
nor I_5(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_6(n4_1_l,IN_1_1_l,IN_2_1_l);
nor I_7(N6147_3_l,IN_3_3_l,n3_3_l);
not I_8(n3_3_l,N6138_3_l);
nor I_9(N6138_3_l,IN_1_3_l,IN_2_3_l);
nor I_10(N1507_6_l,n8_6_l,n9_6_l);
and I_11(N1508_6_l,IN_2_6_l,n6_6_l);
nor I_12(n6_6_l,n7_6_l,n8_6_l);
not I_13(n7_6_l,IN_1_6_l);
nor I_14(n8_6_l,IN_5_6_l,n9_6_l);
and I_15(n9_6_l,IN_3_6_l,IN_4_6_l);
nor I_16(N1371_0_r,n4_0_r,N1508_0_l);
nor I_17(N1508_0_r,n3_0_r,n4_0_r);
nor I_18(n3_0_r,N1372_1_l,N1371_0_l);
not I_19(n4_0_r,N1371_0_l);
not I_20(N1372_1_r,n4_1_r);
nor I_21(N1508_1_r,n4_1_r,N1371_0_l);
nand I_22(n4_1_r,N1508_0_l,N1508_1_l);
not I_23(N1372_4_r,n7_4_r);
nor I_24(N1508_4_r,n6_4_r,n7_4_r);
nor I_25(n6_4_r,n8_4_r,N1508_6_l);
nand I_26(n7_4_r,N1508_1_l,N1507_6_l);
and I_27(n8_4_r,N6147_3_l,N1507_6_l);
nand I_28(n_429_or_0_5_r,n12_5_r,N1508_1_l);
DFFARX1 I_29(n_431_5_r,blif_clk_net_5_r,n2_5_r,G78_5_r,);
nand I_30(n_576_5_r,n11_5_r,N1508_6_l);
not I_31(n_102_5_r,N1508_0_l);
nand I_32(n_547_5_r,n13_5_r,N1371_0_l);
or I_33(n_431_5_r,n14_5_r,N6147_3_l);
not I_34(n2_5_r,blif_reset_net_5_r);
nor I_35(n11_5_r,n12_5_r,N1508_0_l);
not I_36(n12_5_r,N6147_3_l);
nor I_37(n13_5_r,N1508_0_l,N1372_1_l);
and I_38(n14_5_r,n15_5_r,N1372_1_l);
nor I_39(n15_5_r,n16_5_r,N1508_6_l);
not I_40(n16_5_r,N1508_1_l);
nor I_41(N1507_6_r,n8_6_r,n9_6_r);
and I_42(N1508_6_r,n6_6_r,N1507_6_l);
nor I_43(n6_6_r,n7_6_r,n8_6_r);
not I_44(n7_6_r,N1507_6_l);
nor I_45(n8_6_r,n9_6_r,N1508_1_l);
and I_46(n9_6_r,N1508_6_l,N1372_1_l);
endmodule


