module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_7,n8_7,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_7,n8_7,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_7,n8_7,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_7,n8_7,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_7,n8_7,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_32(n_572_1_r_7,n30_7,n31_7);
nand I_33(n_573_1_r_7,n28_7,P6_5_r_14);
nor I_34(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_35(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_36(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_37(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_38(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_39(P6_5_r_7,P6_5_r_internal_7);
or I_40(n_431_0_l_7,n36_7,n_572_1_r_14);
not I_41(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_42(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_43(n27_7,n43_7);
DFFARX1 I_44(G42_1_r_14,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_45(n_42_2_r_14,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_46(n4_1_r_7,n30_7,n38_7);
nor I_47(N1_4_r_7,n27_7,n40_7);
nand I_48(n26_7,n39_7,G199_2_r_14);
not I_49(n5_7,n_549_1_r_14);
DFFARX1 I_50(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_51(n28_7,n26_7,n29_7);
not I_52(n29_7,n_572_1_r_14);
not I_53(n30_7,G42_1_r_14);
nand I_54(n31_7,n27_7,n29_7);
nor I_55(n32_7,ACVQN1_5_l_7,n34_7);
nor I_56(n33_7,n29_7,n_549_1_r_14);
not I_57(n34_7,P6_5_r_14);
nor I_58(n35_7,n43_7,n44_7);
and I_59(n36_7,n37_7,n_573_1_r_14);
nor I_60(n37_7,n30_7,n_569_1_r_14);
nand I_61(n38_7,n29_7,n_549_1_r_14);
nor I_62(n39_7,n_549_1_r_14,ACVQN1_5_r_14);
nor I_63(n40_7,n44_7,n41_7);
nor I_64(n41_7,n34_7,n42_7);
nand I_65(n42_7,n5_7,n_572_1_r_14);
endmodule


