module test_I2727(I1351,I1319,I1447,I1477,I1470,I1335,I2727);
input I1351,I1319,I1447,I1477,I1470,I1335;
output I2727;
wire I2878,I2810,I2759,I3124,I3076,I2861,I2793;
not I_0(I2878,I2861);
nand I_1(I2810,I2793,I1335);
not I_2(I2759,I1477);
nor I_3(I3124,I3076,I2878);
nand I_4(I2727,I2810,I3124);
DFFARX1 I_5(I1447,I1470,I2759,,,I3076,);
not I_6(I2861,I1351);
nor I_7(I2793,I1351,I1319);
endmodule


