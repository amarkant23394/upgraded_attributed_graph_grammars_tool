module test_I10507(I1477,I10185,I6315,I7731,I7604,I1470,I10507);
input I1477,I10185,I6315,I7731,I7604,I1470;
output I10507;
wire I7816,I7850,I10202,I7621,I10219,I10490,I10052,I7977,I10366,I10349,I7541,I10332,I7556,I7550,I7532;
DFFARX1 I_0(I1470,,,I7816,);
nor I_1(I7850,I7816,I7731);
and I_2(I10507,I10490,I10366);
and I_3(I10202,I10185,I7541);
nand I_4(I7621,I7604,I6315);
DFFARX1 I_5(I10202,I1470,I10052,,,I10219,);
DFFARX1 I_6(I7556,I1470,I10052,,,I10490,);
not I_7(I10052,I1477);
DFFARX1 I_8(I1470,,,I7977,);
nand I_9(I10366,I10349,I10219);
and I_10(I10349,I10332,I7550);
DFFARX1 I_11(I1470,,,I7541,);
DFFARX1 I_12(I7532,I1470,I10052,,,I10332,);
nand I_13(I7556,I7621,I7850);
nand I_14(I7550,I7977,I7731);
DFFARX1 I_15(I1470,,,I7532,);
endmodule


