module test_I16274(I13177,I1477,I14503,I1470,I16274);
input I13177,I1477,I14503,I1470;
output I16274;
wire I14338,I16257,I14341,I14472,I14520,I14455,I13174,I14537,I14605,I14370,I14332;
DFFARX1 I_0(I14605,I1470,I14370,,,I14338,);
nand I_1(I16257,I14341,I14338);
DFFARX1 I_2(I14455,I1470,I14370,,,I14341,);
nand I_3(I14472,I14455);
and I_4(I14520,I14503,I13174);
DFFARX1 I_5(I13177,I1470,I14370,,,I14455,);
DFFARX1 I_6(I1470,,,I13174,);
and I_7(I16274,I16257,I14332);
DFFARX1 I_8(I14520,I1470,I14370,,,I14537,);
and I_9(I14605,I14537,I14472);
not I_10(I14370,I1477);
DFFARX1 I_11(I14537,I1470,I14370,,,I14332,);
endmodule


