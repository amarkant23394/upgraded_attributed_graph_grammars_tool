module test_final(G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,n_452_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15,n4_1_l_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n_452_1_r_15,blif_clk_net_1_r_4,n6_4,G42_1_r_15,);
and I_1(n_572_1_r_15,n17_15,n19_15);
nand I_2(n_573_1_r_15,n15_15,n18_15);
nor I_3(n_549_1_r_15,n21_15,n22_15);
nand I_4(n_569_1_r_15,n15_15,n20_15);
nor I_5(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_6(G42_1_l_15,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_15,);
nor I_7(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_8(N1_4_r_15,blif_clk_net_1_r_4,n6_4,G199_4_r_15,);
DFFARX1 I_9(n_573_1_l_15,blif_clk_net_1_r_4,n6_4,G214_4_r_15,);
nor I_10(n4_1_l_15,G18_1_l_15,IN_1_1_l_15);
DFFARX1 I_11(n4_1_l_15,blif_clk_net_1_r_4,n6_4,G42_1_l_15,);
not I_12(n15_15,G42_1_l_15);
DFFARX1 I_13(IN_1_3_l_15,blif_clk_net_1_r_4,n6_4,n17_internal_15,);
not I_14(n17_15,n17_internal_15);
DFFARX1 I_15(IN_2_3_l_15,blif_clk_net_1_r_4,n6_4,n30_15,);
nor I_16(n_572_1_l_15,G15_1_l_15,IN_7_1_l_15);
DFFARX1 I_17(n_572_1_l_15,blif_clk_net_1_r_4,n6_4,n14_internal_15,);
not I_18(n14_15,n14_internal_15);
nand I_19(N1_4_r_15,n25_15,n26_15);
or I_20(n_573_1_l_15,IN_5_1_l_15,IN_9_1_l_15);
nor I_21(n18_15,IN_9_1_l_15,IN_10_1_l_15);
nand I_22(n19_15,n27_15,n28_15);
nand I_23(n20_15,IN_4_3_l_15,n30_15);
not I_24(n21_15,n20_15);
and I_25(n22_15,n17_15,n_572_1_l_15);
nor I_26(n23_15,G18_1_l_15,IN_5_1_l_15);
or I_27(n24_15,IN_9_1_l_15,IN_10_1_l_15);
or I_28(n25_15,G18_1_l_15,n_573_1_l_15);
nand I_29(n26_15,n19_15,n23_15);
not I_30(n27_15,IN_10_1_l_15);
nand I_31(n28_15,IN_4_1_l_15,n29_15);
not I_32(n29_15,G15_1_l_15);
DFFARX1 I_33(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_34(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_35(n_573_1_r_4,n16_4,n_569_1_r_15);
nor I_36(n_549_1_r_4,n22_4,n23_4);
nand I_37(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_38(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_39(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_40(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_41(P6_5_r_4,P6_5_r_internal_4);
or I_42(n_431_0_l_4,n26_4,n_549_1_r_15);
not I_43(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_44(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_45(G199_4_r_15,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_46(n16_4,ACVQN1_5_l_4);
DFFARX1 I_47(G214_4_r_15,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_48(n17_4,n17_internal_4);
nor I_49(n4_1_r_4,n30_4,n31_4);
nand I_50(n19_4,n33_4,n_573_1_r_15);
DFFARX1 I_51(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_52(n15_4,n15_internal_4);
DFFARX1 I_53(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_54(n20_4,n16_4,n_572_1_r_15);
nor I_55(n21_4,G42_1_r_15,n_569_1_r_15);
nand I_56(n22_4,G78_0_l_4,n25_4);
nand I_57(n23_4,n24_4,n_572_1_r_15);
not I_58(n24_4,n_569_1_r_15);
not I_59(n25_4,G42_1_r_15);
and I_60(n26_4,n27_4,ACVQN2_3_r_15);
nor I_61(n27_4,n28_4,G42_1_r_15);
not I_62(n28_4,n_573_1_r_15);
not I_63(n29_4,n30_4);
nand I_64(n30_4,n32_4,n_572_1_r_15);
nand I_65(n31_4,n25_4,n_572_1_r_15);
nor I_66(n32_4,n33_4,n_569_1_r_15);
not I_67(n33_4,n_266_and_0_3_r_15);
endmodule


