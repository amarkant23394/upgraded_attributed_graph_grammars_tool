module test_final(IN_1_0_l_10,IN_2_0_l_10,IN_4_0_l_10,G18_4_l_10,G15_4_l_10,IN_1_4_l_10,IN_4_4_l_10,IN_5_4_l_10,IN_7_4_l_10,IN_9_4_l_10,IN_10_4_l_10,blif_reset_net_0_r_6,blif_clk_net_0_r_6,ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6);
input IN_1_0_l_10,IN_2_0_l_10,IN_4_0_l_10,G18_4_l_10,G15_4_l_10,IN_1_4_l_10,IN_4_4_l_10,IN_5_4_l_10,IN_7_4_l_10,IN_9_4_l_10,IN_10_4_l_10,blif_reset_net_0_r_6,blif_clk_net_0_r_6;
output ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6;
wire n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10,ACVQN2_0_l_10,n_266_and_0_0_l_10,ACVQN1_0_l_10,n4_4_l_10,G42_4_l_10,n_87_4_l_10,n_572_4_l_10,n_573_4_l_10,n_549_4_l_10,n7_4_l_10,n_569_4_l_10,n_452_4_l_10,n12_3_r_10,n_431_3_r_10,n11_3_r_10,n13_3_r_10,n14_3_r_10,n15_3_r_10,n16_3_r_10,n4_4_r_10,n_87_4_r_10,n7_4_r_10,n1_0_r_6,ACVQN1_2_l_6,P6_2_l_6,P6_internal_2_l_6,n_429_or_0_3_l_6,n12_3_l_6,n_431_3_l_6,G78_3_l_6,n_576_3_l_6,n11_3_l_6,n_102_3_l_6,n_547_3_l_6,n13_3_l_6,n14_3_l_6,n15_3_l_6,n16_3_l_6,ACVQN1_0_r_6,P6_internal_2_r_6,n12_3_r_6,n_431_3_r_6,n11_3_r_6,n13_3_r_6,n14_3_r_6,n15_3_r_6,n16_3_r_6,N3_5_r_6,n3_5_r_6;
nand I_0(n_429_or_0_3_r_10,n_266_and_0_0_l_10,n12_3_r_10);
DFFARX1 I_1(n_431_3_r_10,blif_clk_net_0_r_6,n1_0_r_6,G78_3_r_10,);
nand I_2(n_576_3_r_10,ACVQN2_0_l_10,n11_3_r_10);
not I_3(n_102_3_r_10,G42_4_l_10);
nand I_4(n_547_3_r_10,n_569_4_l_10,n13_3_r_10);
DFFARX1 I_5(n4_4_r_10,blif_clk_net_0_r_6,n1_0_r_6,G42_4_r_10,);
nor I_6(n_572_4_r_10,ACVQN2_0_l_10,n_573_4_l_10);
or I_7(n_573_4_r_10,n_569_4_l_10,n_452_4_l_10);
nor I_8(n_549_4_r_10,n_572_4_l_10,n7_4_r_10);
or I_9(n_569_4_r_10,n_572_4_l_10,n_569_4_l_10);
nor I_10(n_452_4_r_10,n_266_and_0_0_l_10,n_452_4_l_10);
DFFARX1 I_11(IN_1_0_l_10,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_l_10,);
and I_12(n_266_and_0_0_l_10,IN_4_0_l_10,ACVQN1_0_l_10);
DFFARX1 I_13(IN_2_0_l_10,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_l_10,);
nor I_14(n4_4_l_10,G18_4_l_10,IN_1_4_l_10);
DFFARX1 I_15(n4_4_l_10,blif_clk_net_0_r_6,n1_0_r_6,G42_4_l_10,);
not I_16(n_87_4_l_10,G15_4_l_10);
nor I_17(n_572_4_l_10,G15_4_l_10,IN_7_4_l_10);
or I_18(n_573_4_l_10,IN_5_4_l_10,IN_9_4_l_10);
nor I_19(n_549_4_l_10,IN_10_4_l_10,n7_4_l_10);
and I_20(n7_4_l_10,IN_4_4_l_10,n_87_4_l_10);
or I_21(n_569_4_l_10,IN_9_4_l_10,IN_10_4_l_10);
nor I_22(n_452_4_l_10,G18_4_l_10,IN_5_4_l_10);
not I_23(n12_3_r_10,n_549_4_l_10);
or I_24(n_431_3_r_10,n_572_4_l_10,n14_3_r_10);
nor I_25(n11_3_r_10,G42_4_l_10,n12_3_r_10);
nor I_26(n13_3_r_10,G42_4_l_10,n_549_4_l_10);
and I_27(n14_3_r_10,ACVQN2_0_l_10,n15_3_r_10);
nor I_28(n15_3_r_10,n_573_4_l_10,n16_3_r_10);
not I_29(n16_3_r_10,n_266_and_0_0_l_10);
nor I_30(n4_4_r_10,n_266_and_0_0_l_10,G42_4_l_10);
not I_31(n_87_4_r_10,ACVQN2_0_l_10);
and I_32(n7_4_r_10,n_452_4_l_10,n_87_4_r_10);
DFFARX1 I_33(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_r_6,);
and I_34(n_266_and_0_0_r_6,n_429_or_0_3_l_6,ACVQN1_0_r_6);
DFFARX1 I_35(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_r_6,);
not I_36(P6_2_r_6,P6_internal_2_r_6);
nand I_37(n_429_or_0_3_r_6,n_102_3_l_6,n12_3_r_6);
DFFARX1 I_38(n_431_3_r_6,blif_clk_net_0_r_6,n1_0_r_6,G78_3_r_6,);
nand I_39(n_576_3_r_6,P6_2_l_6,n11_3_r_6);
not I_40(n_102_3_r_6,ACVQN1_2_l_6);
nand I_41(n_547_3_r_6,n_576_3_l_6,n13_3_r_6);
nor I_42(n_42_5_r_6,ACVQN1_2_l_6,n_429_or_0_3_l_6);
DFFARX1 I_43(N3_5_r_6,blif_clk_net_0_r_6,n1_0_r_6,G199_5_r_6,);
not I_44(n1_0_r_6,blif_reset_net_0_r_6);
DFFARX1 I_45(n_576_3_r_10,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_l_6,);
not I_46(P6_2_l_6,P6_internal_2_l_6);
DFFARX1 I_47(n_547_3_r_10,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_l_6,);
nand I_48(n_429_or_0_3_l_6,n12_3_l_6,G42_4_r_10);
not I_49(n12_3_l_6,n_572_4_r_10);
or I_50(n_431_3_l_6,n14_3_l_6,n_429_or_0_3_r_10);
DFFARX1 I_51(n_431_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,G78_3_l_6,);
nand I_52(n_576_3_l_6,n11_3_l_6,n_452_4_r_10);
nor I_53(n11_3_l_6,n12_3_l_6,n_549_4_r_10);
not I_54(n_102_3_l_6,n_549_4_r_10);
nand I_55(n_547_3_l_6,n13_3_l_6,G78_3_r_10);
nor I_56(n13_3_l_6,n_102_3_r_10,n_549_4_r_10);
and I_57(n14_3_l_6,n15_3_l_6,n_569_4_r_10);
nor I_58(n15_3_l_6,n16_3_l_6,n_573_4_r_10);
not I_59(n16_3_l_6,G42_4_r_10);
DFFARX1 I_60(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_r_6,);
DFFARX1 I_61(n_576_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_r_6,);
not I_62(n12_3_r_6,P6_2_l_6);
or I_63(n_431_3_r_6,n_429_or_0_3_l_6,n14_3_r_6);
nor I_64(n11_3_r_6,ACVQN1_2_l_6,n12_3_r_6);
nor I_65(n13_3_r_6,ACVQN1_2_l_6,n_547_3_l_6);
and I_66(n14_3_r_6,ACVQN1_2_l_6,n15_3_r_6);
nor I_67(n15_3_r_6,P6_2_l_6,n16_3_r_6);
not I_68(n16_3_r_6,n_102_3_l_6);
and I_69(N3_5_r_6,n_102_3_l_6,n3_5_r_6);
nand I_70(n3_5_r_6,n_429_or_0_3_l_6,n_547_3_l_6);
endmodule


