module test_I3577(I3103,I1902,I1294,I2569,I1301,I3577);
input I3103,I1902,I1294,I2569,I1301;
output I3577;
wire I3263,I3560,I2563,I3379,I2548,I2583,I2560,I3280,I2993,I2566,I2945,I3543,I3297;
not I_0(I3263,I2569);
nand I_1(I3560,I3543,I3297);
nand I_2(I2563,I3103,I2993);
not I_3(I3379,I2548);
DFFARX1 I_4(I2945,I1294,I2583,,,I2548,);
not I_5(I2583,I1301);
DFFARX1 I_6(I1294,I2583,,,I2560,);
nor I_7(I3280,I2548,I2560);
and I_8(I3577,I3379,I3560);
nor I_9(I2993,I2945);
not I_10(I2566,I2945);
DFFARX1 I_11(I1902,I1294,I2583,,,I2945,);
nand I_12(I3543,I3263,I2566);
nand I_13(I3297,I3280,I2563);
endmodule


