module test_I8657(I6265,I1477,I6127,I5785,I1470,I8657);
input I6265,I1477,I6127,I5785,I1470;
output I8657;
wire I8233,I8640,I8216,I5751,I8623,I5743,I6079,I5802,I8298,I5719,I5740,I8315,I5722;
not I_0(I8233,I5722);
not I_1(I8640,I8623);
not I_2(I8216,I1477);
not I_3(I5751,I1477);
DFFARX1 I_4(I5743,I1470,I8216,,,I8623,);
nand I_5(I5743,I6127,I6079);
nor I_6(I8657,I8315,I8640);
nor I_7(I6079,I5802);
DFFARX1 I_8(I5785,I1470,I5751,,,I5802,);
nor I_9(I8298,I8233,I5719);
DFFARX1 I_10(I6265,I1470,I5751,,,I5719,);
not I_11(I5740,I5802);
nand I_12(I8315,I8298,I5740);
DFFARX1 I_13(I1470,I5751,,,I5722,);
endmodule


