module test_I2087(I1444,I1294,I1301,I2087);
input I1444,I1294,I1301;
output I2087;
wire I1342,I2070,I1509,I1310,I1577;
not I_0(I2087,I2070);
not I_1(I1342,I1301);
not I_2(I2070,I1310);
DFFARX1 I_3(I1294,I1342,,,I1509,);
DFFARX1 I_4(I1577,I1294,I1342,,,I1310,);
and I_5(I1577,I1509,I1444);
endmodule


