module test_I14370(I1477,I14370);
input I1477;
output I14370;
wire ;
not I_0(I14370,I1477);
endmodule


