module test_I3220(I2554,I1902,I1294,I1301,I3220);
input I2554,I1902,I1294,I1301;
output I3220;
wire I3379,I2548,I2583,I2945,I3246,I3797,I3715,I3698;
not I_0(I3379,I2548);
DFFARX1 I_1(I2945,I1294,I2583,,,I2548,);
not I_2(I2583,I1301);
DFFARX1 I_3(I1902,I1294,I2583,,,I2945,);
nand I_4(I3220,I3379,I3797);
not I_5(I3246,I1301);
not I_6(I3797,I3715);
not I_7(I3715,I3698);
DFFARX1 I_8(I2554,I1294,I3246,,,I3698,);
endmodule


