module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_7,n8_7,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_7,n8_7,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_7,n8_7,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_7,n8_7,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_7,n8_7,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_7,n8_7,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_33(n_572_1_r_7,n30_7,n31_7);
nand I_34(n_573_1_r_7,n28_7,ACVQN1_5_r_16);
nor I_35(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_36(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_37(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_38(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_39(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_40(P6_5_r_7,P6_5_r_internal_7);
or I_41(n_431_0_l_7,n36_7,n_572_1_r_16);
not I_42(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_43(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_44(n27_7,n43_7);
DFFARX1 I_45(n_452_1_r_16,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_46(G214_4_r_16,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_47(n4_1_r_7,n30_7,n38_7);
nor I_48(N1_4_r_7,n27_7,n40_7);
nand I_49(n26_7,n39_7,G42_1_r_16);
not I_50(n5_7,n_569_1_r_16);
DFFARX1 I_51(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_52(n28_7,n26_7,n29_7);
not I_53(n29_7,P6_5_r_16);
not I_54(n30_7,G42_1_r_16);
nand I_55(n31_7,n27_7,n29_7);
nor I_56(n32_7,ACVQN1_5_l_7,n34_7);
nor I_57(n33_7,n29_7,n_569_1_r_16);
not I_58(n34_7,ACVQN1_5_r_16);
nor I_59(n35_7,n43_7,n44_7);
and I_60(n36_7,n37_7,n_573_1_r_16);
nor I_61(n37_7,n30_7,n_549_1_r_16);
nand I_62(n38_7,n29_7,n_569_1_r_16);
nor I_63(n39_7,n_569_1_r_16,G199_4_r_16);
nor I_64(n40_7,n44_7,n41_7);
nor I_65(n41_7,n34_7,n42_7);
nand I_66(n42_7,n5_7,P6_5_r_16);
endmodule


