module test_final(IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_7_r,blif_reset_net_7_r,N1371_0_r,N1508_0_r,N1507_6_r,N1508_6_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r);
input IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_7_r,blif_reset_net_7_r;
output N1371_0_r,N1508_0_r,N1507_6_r,N1508_6_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r;
wire N6147_2_l,n5_2_l,n6_2_l,N6138_2_l,n7_2_l,N1507_6_l,N1508_6_l,n6_6_l,n7_6_l,n8_6_l,n9_6_l,N6150_9_l,N6147_9_l,N6134_9_l,n3_9_l,I_BUFF_1_9_l,n3_0_r,n4_0_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,n_87_7_r,n4_7_r,n2_7_r,n7_7_r,N6150_9_r,n3_9_r;
nor I_0(N6147_2_l,n5_2_l,n6_2_l);
nor I_1(n5_2_l,IN_5_2_l,n7_2_l);
not I_2(n6_2_l,N6138_2_l);
nor I_3(N6138_2_l,IN_1_2_l,IN_2_2_l);
nor I_4(n7_2_l,IN_3_2_l,IN_4_2_l);
nor I_5(N1507_6_l,n8_6_l,n9_6_l);
and I_6(N1508_6_l,IN_2_6_l,n6_6_l);
nor I_7(n6_6_l,n7_6_l,n8_6_l);
not I_8(n7_6_l,IN_1_6_l);
nor I_9(n8_6_l,IN_5_6_l,n9_6_l);
and I_10(n9_6_l,IN_3_6_l,IN_4_6_l);
not I_11(N6150_9_l,IN_2_9_l);
nor I_12(N6147_9_l,N6150_9_l,n3_9_l);
nor I_13(N6134_9_l,IN_5_9_l,n3_9_l);
nor I_14(n3_9_l,IN_3_9_l,IN_4_9_l);
buf I_15(I_BUFF_1_9_l,IN_1_9_l);
nor I_16(N1371_0_r,n4_0_r,N1507_6_l);
nor I_17(N1508_0_r,n3_0_r,n4_0_r);
nor I_18(n3_0_r,N6147_2_l,I_BUFF_1_9_l);
not I_19(n4_0_r,N6134_9_l);
nor I_20(N1507_6_r,n8_6_r,n9_6_r);
and I_21(N1508_6_r,n6_6_r,N1508_6_l);
nor I_22(n6_6_r,n7_6_r,n8_6_r);
not I_23(n7_6_r,N6134_9_l);
nor I_24(n8_6_r,n9_6_r,N1507_6_l);
and I_25(n9_6_r,N6147_2_l,N6147_9_l);
DFFARX1 I_26(n4_7_r,blif_clk_net_7_r,n2_7_r,G42_7_r,);
not I_27(n_87_7_r,N6147_9_l);
nor I_28(n_572_7_r,N1508_6_l,N6147_9_l);
or I_29(n_573_7_r,I_BUFF_1_9_l,N1507_6_l);
nor I_30(n_549_7_r,n7_7_r,N6147_2_l);
or I_31(n_569_7_r,N6147_2_l,N1507_6_l);
nor I_32(n_452_7_r,I_BUFF_1_9_l,N6147_9_l);
nor I_33(n4_7_r,N6147_9_l,N6147_2_l);
not I_34(n2_7_r,blif_reset_net_7_r);
and I_35(n7_7_r,n_87_7_r,N6134_9_l);
not I_36(N6150_9_r,N6134_9_l);
nor I_37(N6147_9_r,N6150_9_r,n3_9_r);
nor I_38(N6134_9_r,n3_9_r,I_BUFF_1_9_l);
nor I_39(n3_9_r,N1507_6_l,N1508_6_l);
buf I_40(I_BUFF_1_9_r,N6147_9_l);
endmodule


