module Benchmark_testing65000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2683,I2690,I6284,I6263,I6266,I6275,I6281,I6278,I6272,I6269,I8664,I8643,I8646,I8655,I8661,I8658,I8652,I8649,I11642,I11633,I11630,I11636,I11624,I11618,I11639,I11627,I11621,I147999,I147975,I147987,I147981,I147996,I147990,I147984,I147978,I147993,I229561,I229585,I229567,I229570,I229558,I229576,I229579,I229564,I229573,I229582,I424096,I424093,I424078,I424090,I424084,I424072,I424081,I424087,I424075,I468834,I468831,I468822,I468825,I468819,I468828,I468816,I468840,I468837,I476348,I476345,I476336,I476339,I476333,I476342,I476330,I476354,I476351,I508713,I508716,I508698,I508707,I508719,I508710,I508701,I508704,I508722,I541659,I541662,I541644,I541653,I541665,I541656,I541647,I541650,I541668,I550907,I550910,I550892,I550901,I550913,I550904,I550895,I550898,I550916,I552641,I552644,I552626,I552635,I552647,I552638,I552629,I552632,I552650,I910287,I910275,I910296,I910272,I910293,I910284,I910290,I910281,I910278,I1085222,I1085237,I1085219,I1085231,I1085246,I1085243,I1085240,I1085234,I1085228,I1085225,I1085817,I1085832,I1085814,I1085826,I1085841,I1085838,I1085835,I1085829,I1085823,I1085820);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2683,I2690;
output I6284,I6263,I6266,I6275,I6281,I6278,I6272,I6269,I8664,I8643,I8646,I8655,I8661,I8658,I8652,I8649,I11642,I11633,I11630,I11636,I11624,I11618,I11639,I11627,I11621,I147999,I147975,I147987,I147981,I147996,I147990,I147984,I147978,I147993,I229561,I229585,I229567,I229570,I229558,I229576,I229579,I229564,I229573,I229582,I424096,I424093,I424078,I424090,I424084,I424072,I424081,I424087,I424075,I468834,I468831,I468822,I468825,I468819,I468828,I468816,I468840,I468837,I476348,I476345,I476336,I476339,I476333,I476342,I476330,I476354,I476351,I508713,I508716,I508698,I508707,I508719,I508710,I508701,I508704,I508722,I541659,I541662,I541644,I541653,I541665,I541656,I541647,I541650,I541668,I550907,I550910,I550892,I550901,I550913,I550904,I550895,I550898,I550916,I552641,I552644,I552626,I552635,I552647,I552638,I552629,I552632,I552650,I910287,I910275,I910296,I910272,I910293,I910284,I910290,I910281,I910278,I1085222,I1085237,I1085219,I1085231,I1085246,I1085243,I1085240,I1085234,I1085228,I1085225,I1085817,I1085832,I1085814,I1085826,I1085841,I1085838,I1085835,I1085829,I1085823,I1085820;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2683,I2690,I2722,I630172,I2748,I2756,I630163,I2773,I2714,I630169,I2813,I2821,I2838,I2855,I630175,I2872,I2889,I2693,I2920,I2937,I2954,I630184,I630181,I2696,I2985,I3002,I3019,I630166,I3036,I3053,I3070,I2705,I3101,I3118,I3135,I2711,I3166,I2708,I3197,I630178,I3223,I3231,I3248,I2702,I2699,I3317,I600046,I3343,I3351,I600025,I3368,I3309,I600034,I3408,I3416,I3433,I600040,I3450,I600037,I3467,I3484,I3288,I3515,I3532,I3549,I600028,I600022,I3291,I3580,I3597,I600043,I3614,I3631,I3648,I3665,I3300,I3696,I600031,I3713,I3730,I3306,I3761,I3303,I3792,I3818,I3826,I3843,I3297,I3294,I3912,I1025430,I3938,I3946,I1025439,I3963,I3904,I1025445,I4003,I4011,I4028,I1025433,I4045,I1025442,I4062,I4079,I3883,I4110,I4127,I4144,I1025451,I1025448,I3886,I4175,I4192,I1025436,I4209,I1025454,I4226,I4243,I4260,I3895,I4291,I4308,I4325,I3901,I4356,I3898,I4387,I1025457,I4413,I4421,I4438,I3892,I3889,I4507,I482691,I4533,I4541,I482709,I4558,I4499,I482703,I4598,I4606,I4623,I482694,I4640,I4657,I4674,I4478,I4705,I4722,I4739,I482700,I482688,I4481,I4770,I4787,I482706,I4804,I482712,I4821,I4838,I4855,I4490,I4886,I4903,I4920,I4496,I4951,I4493,I4982,I482697,I5008,I5016,I5033,I4487,I4484,I5102,I527218,I5128,I5136,I527197,I5153,I5094,I527206,I5193,I5201,I5218,I527212,I5235,I527209,I5252,I5269,I5073,I5300,I5317,I5334,I527200,I527194,I5076,I5365,I5382,I527215,I5399,I5416,I5433,I5450,I5085,I5481,I527203,I5498,I5515,I5091,I5546,I5088,I5577,I5603,I5611,I5628,I5082,I5079,I5697,I388359,I5723,I5731,I388341,I5748,I5689,I388353,I5788,I5796,I5813,I388338,I5830,I388347,I5847,I5864,I5668,I5895,I5912,I5929,I388344,I388365,I5671,I5960,I5977,I388356,I5994,I388362,I6011,I6028,I6045,I5680,I6076,I6093,I6110,I5686,I6141,I5683,I6172,I388350,I6198,I6206,I6223,I5677,I5674,I6292,I74343,I6318,I6326,I74334,I6343,I74355,I6383,I6391,I6408,I74331,I6425,I6442,I6459,I6490,I6507,I6524,I74340,I6555,I6572,I74352,I6589,I74349,I6606,I6623,I6640,I6671,I74346,I6688,I6705,I6736,I6767,I74337,I6793,I6801,I6818,I6887,I287016,I6913,I6921,I287007,I6938,I6879,I287010,I6978,I6986,I7003,I287004,I7020,I287013,I7037,I7054,I6858,I7085,I7102,I7119,I287001,I287019,I6861,I7150,I7167,I7184,I287025,I7201,I7218,I7235,I6870,I7266,I287022,I7283,I7300,I6876,I7331,I6873,I7362,I287028,I7388,I7396,I7413,I6867,I6864,I7482,I364967,I7508,I7516,I364949,I7533,I7474,I364961,I7573,I7581,I7598,I364946,I7615,I364955,I7632,I7649,I7453,I7680,I7697,I7714,I364952,I364973,I7456,I7745,I7762,I364964,I7779,I364970,I7796,I7813,I7830,I7465,I7861,I7878,I7895,I7471,I7926,I7468,I7957,I364958,I7983,I7991,I8008,I7462,I7459,I8077,I1038229,I8103,I8111,I1038220,I8128,I8069,I1038223,I8168,I8176,I8193,I1038235,I8210,I1038226,I8227,I8244,I8048,I8275,I8292,I8309,I1038214,I8051,I8340,I8357,I1038238,I8374,I1038217,I8391,I8408,I8425,I8060,I8456,I1038232,I8473,I8490,I8066,I8521,I8063,I8552,I1038241,I8578,I8586,I8603,I8057,I8054,I8672,I858255,I8698,I8706,I8723,I858270,I8763,I8771,I8788,I858267,I8805,I858276,I8822,I8839,I8870,I8887,I8904,I858264,I858273,I8935,I8952,I858261,I8969,I858252,I8986,I9003,I9020,I9051,I858258,I9068,I9085,I9116,I9147,I9173,I9181,I9198,I9267,I444543,I9293,I9301,I444561,I9318,I9259,I444555,I9358,I9366,I9383,I444546,I9400,I9417,I9434,I9238,I9465,I9482,I9499,I444552,I444540,I9241,I9530,I9547,I444558,I9564,I444564,I9581,I9598,I9615,I9250,I9646,I9663,I9680,I9256,I9711,I9253,I9742,I444549,I9768,I9776,I9793,I9247,I9244,I9862,I699340,I9888,I9896,I699331,I9913,I9854,I699334,I9953,I9961,I9978,I699346,I9995,I699325,I10012,I10029,I9833,I10060,I10077,I10094,I699337,I699343,I9836,I10125,I10142,I699328,I10159,I699319,I10176,I10193,I10210,I9845,I10241,I10258,I10275,I9851,I10306,I9848,I10337,I699322,I10363,I10371,I10388,I9842,I9839,I10457,I912009,I10483,I10491,I10508,I10449,I912024,I10548,I10556,I10573,I912021,I10590,I912030,I10607,I10624,I10428,I10655,I10672,I10689,I912018,I912027,I10431,I10720,I10737,I912015,I10754,I912006,I10771,I10788,I10805,I10440,I10836,I912012,I10853,I10870,I10446,I10901,I10443,I10932,I10958,I10966,I10983,I10437,I10434,I11052,I851319,I11078,I11086,I11103,I11044,I851334,I11143,I11151,I11168,I851331,I11185,I851340,I11202,I11219,I11023,I11250,I11267,I11284,I851328,I851337,I11026,I11315,I11332,I851325,I11349,I851316,I11366,I11383,I11400,I11035,I11431,I851322,I11448,I11465,I11041,I11496,I11038,I11527,I11553,I11561,I11578,I11032,I11029,I11650,I93306,I11676,I11693,I11701,I11718,I93321,I11735,I93324,I11761,I93318,I11806,I11814,I93327,I11831,I93303,I11871,I11879,I11924,I93309,I11941,I93312,I11967,I11975,I12006,I12023,I93315,I12040,I12057,I12074,I12105,I12177,I1003617,I12203,I12220,I12228,I12245,I1003620,I1003614,I12262,I1003623,I12288,I12169,I12160,I1003611,I12333,I12341,I1003626,I12358,I12157,I1003602,I12398,I12406,I12163,I12151,I12451,I1003605,I12468,I12494,I12502,I12145,I12533,I12550,I1003608,I12567,I12584,I12601,I12166,I12632,I12154,I12148,I12704,I619632,I12730,I12747,I12755,I12772,I619623,I619644,I12789,I619626,I12815,I12696,I12687,I12860,I12868,I619641,I12885,I12684,I619635,I12925,I12933,I12690,I12678,I12978,I619629,I619638,I12995,I13021,I13029,I12672,I13060,I13077,I13094,I13111,I13128,I12693,I13159,I12681,I12675,I13231,I752315,I13257,I13274,I13282,I13299,I752291,I752318,I13316,I752303,I13342,I13223,I13214,I752309,I13387,I13395,I752294,I13412,I13211,I752312,I13452,I13460,I13217,I13205,I13505,I752297,I752300,I13522,I13548,I13556,I13199,I13587,I13604,I752306,I13621,I13638,I13655,I13220,I13686,I13208,I13202,I13758,I541072,I13784,I13801,I13809,I13826,I541087,I541090,I13843,I541069,I13869,I13750,I13741,I541075,I13914,I13922,I541081,I13939,I13738,I13979,I13987,I13744,I13732,I14032,I541084,I541066,I14049,I541078,I14075,I14083,I13726,I14114,I14131,I14148,I14165,I14182,I13747,I14213,I13735,I13729,I14285,I676021,I14311,I14328,I14336,I14353,I676012,I676033,I14370,I676015,I14396,I14277,I14268,I14441,I14449,I676030,I14466,I14265,I676024,I14506,I14514,I14271,I14259,I14559,I676018,I676027,I14576,I14602,I14610,I14253,I14641,I14658,I14675,I14692,I14709,I14274,I14740,I14262,I14256,I14812,I191416,I14838,I14855,I14863,I14880,I191434,I191419,I14897,I191422,I14923,I14804,I14795,I191410,I14968,I14976,I191413,I14993,I14792,I191425,I15033,I15041,I14798,I14786,I15086,I191431,I191428,I15103,I15129,I15137,I14780,I15168,I15185,I15202,I15219,I15236,I14801,I15267,I14789,I14783,I15339,I456115,I15365,I15382,I15390,I15407,I456100,I456118,I15424,I456112,I15450,I15331,I15322,I456109,I15495,I15503,I15520,I15319,I456103,I15560,I15568,I15325,I15313,I15613,I456124,I456106,I15630,I456121,I15656,I15664,I15307,I15695,I15712,I15729,I15746,I15763,I15328,I15794,I15316,I15310,I15866,I356786,I15892,I15909,I15917,I15934,I356789,I15951,I356810,I15977,I15858,I15849,I356798,I16022,I16030,I356801,I16047,I15846,I356807,I16087,I16095,I15852,I15840,I16140,I356804,I356792,I16157,I356795,I16183,I16191,I15834,I16222,I16239,I356813,I16256,I16273,I16290,I15855,I16321,I15843,I15837,I16393,I236963,I16419,I16436,I16444,I16461,I236960,I236954,I16478,I236948,I16504,I16385,I16376,I236936,I16549,I16557,I236945,I16574,I16373,I236942,I16614,I16622,I16379,I16367,I16667,I236939,I236957,I16684,I16710,I16718,I16361,I16749,I16766,I236951,I16783,I16800,I16817,I16382,I16848,I16370,I16364,I16920,I258043,I16946,I16963,I16971,I16988,I258040,I258034,I17005,I258028,I17031,I16912,I16903,I258016,I17076,I17084,I258025,I17101,I16900,I258022,I17141,I17149,I16906,I16894,I17194,I258019,I258037,I17211,I17237,I17245,I16888,I17276,I17293,I258031,I17310,I17327,I17344,I16909,I17375,I16897,I16891,I17447,I17473,I17490,I17498,I17515,I17532,I17558,I17439,I17430,I17603,I17611,I17628,I17427,I17668,I17676,I17433,I17421,I17721,I17738,I17764,I17772,I17415,I17803,I17820,I17837,I17854,I17871,I17436,I17902,I17424,I17418,I17974,I159286,I18000,I18017,I18025,I18042,I159304,I159289,I18059,I159292,I18085,I17966,I17957,I159280,I18130,I18138,I159283,I18155,I17954,I159295,I18195,I18203,I17960,I17948,I18248,I159301,I159298,I18265,I18291,I18299,I17942,I18330,I18347,I18364,I18381,I18398,I17963,I18429,I17951,I17945,I18501,I1045354,I18527,I18544,I18552,I18569,I1045357,I1045363,I18586,I1045372,I18612,I18493,I18484,I1045375,I18657,I18665,I1045366,I18682,I18481,I18722,I18730,I18487,I18475,I18775,I1045381,I1045360,I18792,I1045369,I18818,I18826,I18469,I18857,I18874,I1045378,I18891,I18908,I18925,I18490,I18956,I18478,I18472,I19028,I487327,I19054,I19071,I19079,I19096,I487312,I487330,I19113,I487324,I19139,I19020,I19011,I487321,I19184,I19192,I19209,I19008,I487315,I19249,I19257,I19014,I19002,I19302,I487336,I487318,I19319,I487333,I19345,I19353,I18996,I19384,I19401,I19418,I19435,I19452,I19017,I19483,I19005,I18999,I19555,I606386,I19581,I19598,I19606,I19623,I606401,I606404,I19640,I606383,I19666,I19547,I19538,I606389,I19711,I19719,I606395,I19736,I19535,I19776,I19784,I19541,I19529,I19829,I606398,I606380,I19846,I606392,I19872,I19880,I19523,I19911,I19928,I19945,I19962,I19979,I19544,I20010,I19532,I19526,I20082,I542228,I20108,I20125,I20133,I20150,I542243,I542246,I20167,I542225,I20193,I20074,I20065,I542231,I20238,I20246,I542237,I20263,I20062,I20303,I20311,I20068,I20056,I20356,I542240,I542222,I20373,I542234,I20399,I20407,I20050,I20438,I20455,I20472,I20489,I20506,I20071,I20537,I20059,I20053,I20609,I729705,I20635,I20652,I20660,I20677,I729681,I729708,I20694,I729693,I20720,I20601,I20592,I729699,I20765,I20773,I729684,I20790,I20589,I729702,I20830,I20838,I20595,I20583,I20883,I729687,I729690,I20900,I20926,I20934,I20577,I20965,I20982,I729696,I20999,I21016,I21033,I20598,I21064,I20586,I20580,I21136,I520842,I21162,I21179,I21187,I21204,I520857,I520860,I21221,I520839,I21247,I21128,I21119,I520845,I21292,I21300,I520851,I21317,I21116,I21357,I21365,I21122,I21110,I21410,I520854,I520836,I21427,I520848,I21453,I21461,I21104,I21492,I21509,I21526,I21543,I21560,I21125,I21591,I21113,I21107,I21663,I730997,I21689,I21706,I21714,I21731,I730973,I731000,I21748,I730985,I21774,I21655,I21646,I730991,I21819,I21827,I730976,I21844,I21643,I730994,I21884,I21892,I21649,I21637,I21937,I730979,I730982,I21954,I21980,I21988,I21631,I22019,I22036,I730988,I22053,I22070,I22087,I21652,I22118,I21640,I21634,I22190,I284920,I22216,I22233,I22241,I22258,I284917,I284911,I22275,I284905,I22301,I22182,I22173,I284893,I22346,I22354,I284902,I22371,I22170,I284899,I22411,I22419,I22176,I22164,I22464,I284896,I284914,I22481,I22507,I22515,I22158,I22546,I22563,I284908,I22580,I22597,I22614,I22179,I22645,I22167,I22161,I22717,I969534,I22743,I22760,I22768,I22785,I969552,I969546,I22802,I969555,I22828,I22709,I22700,I969540,I22873,I22881,I969549,I22898,I22697,I969537,I22938,I22946,I22703,I22691,I22991,I969558,I969543,I23008,I23034,I23042,I22685,I23073,I23090,I23107,I23124,I23141,I22706,I23172,I22694,I22688,I23244,I216937,I23270,I23287,I23295,I23312,I216934,I216928,I23329,I216922,I23355,I23236,I23227,I216910,I23400,I23408,I216919,I23425,I23224,I216916,I23465,I23473,I23230,I23218,I23518,I216913,I216931,I23535,I23561,I23569,I23212,I23600,I23617,I216925,I23634,I23651,I23668,I23233,I23699,I23221,I23215,I23771,I228531,I23797,I23814,I23822,I23839,I228528,I228522,I23856,I228516,I23882,I23763,I23754,I228504,I23927,I23935,I228513,I23952,I23751,I228510,I23992,I24000,I23757,I23745,I24045,I228507,I228525,I24062,I24088,I24096,I23739,I24127,I24144,I228519,I24161,I24178,I24195,I23760,I24226,I23748,I23742,I24298,I1020379,I24324,I24341,I24349,I24366,I1020382,I1020376,I24383,I1020385,I24409,I24290,I24281,I1020373,I24454,I24462,I1020388,I24479,I24278,I1020364,I24519,I24527,I24284,I24272,I24572,I1020367,I24589,I24615,I24623,I24266,I24654,I24671,I1020370,I24688,I24705,I24722,I24287,I24753,I24275,I24269,I24825,I744563,I24851,I24868,I24876,I24893,I744539,I744566,I24910,I744551,I24936,I24817,I24808,I744557,I24981,I24989,I744542,I25006,I24805,I744560,I25046,I25054,I24811,I24799,I25099,I744545,I744548,I25116,I25142,I25150,I24793,I25181,I25198,I744554,I25215,I25232,I25249,I24814,I25280,I24802,I24796,I25352,I79077,I25378,I25395,I25403,I25420,I79092,I25437,I79095,I25463,I25344,I25335,I79089,I25508,I25516,I79098,I25533,I25332,I79074,I25573,I25581,I25338,I25326,I25626,I79080,I25643,I79083,I25669,I25677,I25320,I25708,I25725,I79086,I25742,I25759,I25776,I25341,I25807,I25329,I25323,I25879,I808006,I25905,I25922,I25930,I25947,I808000,I808021,I25964,I25990,I25871,I25862,I808003,I26035,I26043,I808012,I26060,I25859,I26100,I26108,I25865,I25853,I26153,I808018,I26170,I808009,I26196,I26204,I25847,I26235,I26252,I808015,I26269,I26286,I26303,I25868,I26334,I25856,I25850,I26406,I471721,I26432,I26449,I26457,I26474,I471706,I471724,I26491,I471718,I26517,I26398,I26389,I471715,I26562,I26570,I26587,I26386,I471709,I26627,I26635,I26392,I26380,I26680,I471730,I471712,I26697,I471727,I26723,I26731,I26374,I26762,I26779,I26796,I26813,I26830,I26395,I26861,I26383,I26377,I26933,I114670,I26959,I26976,I26984,I27001,I114673,I114655,I27018,I114661,I27044,I26925,I26916,I114664,I27089,I27097,I27114,I26913,I114676,I27154,I27162,I26919,I26907,I27207,I114679,I114667,I27224,I114658,I27250,I27258,I26901,I27289,I27306,I114682,I27323,I27340,I27357,I26922,I27388,I26910,I26904,I27460,I69064,I27486,I27503,I27511,I27528,I69079,I27545,I69082,I27571,I27452,I27443,I69076,I27616,I27624,I69085,I27641,I27440,I69061,I27681,I27689,I27446,I27434,I27734,I69067,I27751,I69070,I27777,I27785,I27428,I27816,I27833,I69073,I27850,I27867,I27884,I27449,I27915,I27437,I27431,I27987,I500034,I28013,I28030,I28038,I28055,I500049,I500052,I28072,I500031,I28098,I27979,I27970,I500037,I28143,I28151,I500043,I28168,I27967,I28208,I28216,I27973,I27961,I28261,I500046,I500028,I28278,I500040,I28304,I28312,I27955,I28343,I28360,I28377,I28394,I28411,I27976,I28442,I27964,I27958,I28514,I598872,I28540,I28557,I28565,I28582,I598887,I598890,I28599,I598869,I28625,I28506,I28497,I598875,I28670,I28678,I598881,I28695,I28494,I28735,I28743,I28500,I28488,I28788,I598884,I598866,I28805,I598878,I28831,I28839,I28482,I28870,I28887,I28904,I28921,I28938,I28503,I28969,I28491,I28485,I29041,I1037024,I29067,I29084,I29092,I29109,I1037027,I1037033,I29126,I1037042,I29152,I29033,I29024,I1037045,I29197,I29205,I1037036,I29222,I29021,I29262,I29270,I29027,I29015,I29315,I1037051,I1037030,I29332,I1037039,I29358,I29366,I29009,I29397,I29414,I1037048,I29431,I29448,I29465,I29030,I29496,I29018,I29012,I29568,I1063799,I29594,I29611,I29619,I29636,I1063802,I1063808,I29653,I1063817,I29679,I29560,I29551,I1063820,I29724,I29732,I1063811,I29749,I29548,I29789,I29797,I29554,I29542,I29842,I1063826,I1063805,I29859,I1063814,I29885,I29893,I29536,I29924,I29941,I1063823,I29958,I29975,I29992,I29557,I30023,I29545,I29539,I30095,I335570,I30121,I30138,I30146,I30163,I335573,I30180,I335594,I30206,I30087,I30078,I335582,I30251,I30259,I335585,I30276,I30075,I335591,I30316,I30324,I30081,I30069,I30369,I335588,I335576,I30386,I335579,I30412,I30420,I30063,I30451,I30468,I335597,I30485,I30502,I30519,I30084,I30550,I30072,I30066,I30622,I115860,I30648,I30665,I30673,I30690,I115863,I115845,I30707,I115851,I30733,I30614,I30605,I115854,I30778,I30786,I30803,I30602,I115866,I30843,I30851,I30608,I30596,I30896,I115869,I115857,I30913,I115848,I30939,I30947,I30590,I30978,I30995,I115872,I31012,I31029,I31046,I30611,I31077,I30599,I30593,I31149,I960830,I31175,I31192,I31200,I31217,I960848,I960842,I31234,I960851,I31260,I31141,I31132,I960836,I31305,I31313,I960845,I31330,I31129,I960833,I31370,I31378,I31135,I31123,I31423,I960854,I960839,I31440,I31466,I31474,I31117,I31505,I31522,I31539,I31556,I31573,I31138,I31604,I31126,I31120,I31676,I537026,I31702,I31719,I31727,I31744,I537041,I537044,I31761,I537023,I31787,I31668,I31659,I537029,I31832,I31840,I537035,I31857,I31656,I31897,I31905,I31662,I31650,I31950,I537038,I537020,I31967,I537032,I31993,I32001,I31644,I32032,I32049,I32066,I32083,I32100,I31665,I32131,I31653,I31647,I32203,I990901,I32229,I32246,I32254,I32271,I990904,I990898,I32288,I990907,I32314,I32195,I32186,I990895,I32359,I32367,I990910,I32384,I32183,I990886,I32424,I32432,I32189,I32177,I32477,I990889,I32494,I32520,I32528,I32171,I32559,I32576,I990892,I32593,I32610,I32627,I32192,I32658,I32180,I32174,I32730,I489061,I32756,I32773,I32781,I32798,I489046,I489064,I32815,I489058,I32841,I32722,I32713,I489055,I32886,I32894,I32911,I32710,I489049,I32951,I32959,I32716,I32704,I33004,I489070,I489052,I33021,I489067,I33047,I33055,I32698,I33086,I33103,I33120,I33137,I33154,I32719,I33185,I32707,I32701,I33257,I307581,I33283,I33300,I33308,I33325,I307578,I307572,I33342,I307566,I33368,I33249,I33240,I307554,I33413,I33421,I307563,I33438,I33237,I307560,I33478,I33486,I33243,I33231,I33531,I307557,I307575,I33548,I33574,I33582,I33225,I33613,I33630,I307569,I33647,I33664,I33681,I33246,I33712,I33234,I33228,I33784,I561880,I33810,I33827,I33835,I33852,I561895,I561898,I33869,I561877,I33895,I33776,I33767,I561883,I33940,I33948,I561889,I33965,I33764,I34005,I34013,I33770,I33758,I34058,I561892,I561874,I34075,I561886,I34101,I34109,I33752,I34140,I34157,I34174,I34191,I34208,I33773,I34239,I33761,I33755,I34311,I951334,I34337,I34354,I34362,I34379,I951322,I951313,I34396,I951310,I34422,I34303,I34294,I951316,I34467,I34475,I951328,I34492,I34291,I951325,I34532,I34540,I34297,I34285,I34585,I951319,I34602,I951331,I34628,I34636,I34279,I34667,I34684,I34701,I34718,I34735,I34300,I34766,I34288,I34282,I34838,I649144,I34864,I34881,I34889,I34906,I649135,I649156,I34923,I649138,I34949,I34830,I34821,I34994,I35002,I649153,I35019,I34818,I649147,I35059,I35067,I34824,I34812,I35112,I649141,I649150,I35129,I35155,I35163,I34806,I35194,I35211,I35228,I35245,I35262,I34827,I35293,I34815,I34809,I35365,I521420,I35391,I35408,I35416,I35433,I521435,I521438,I35450,I521417,I35476,I35357,I35348,I521423,I35521,I35529,I521429,I35546,I35345,I35586,I35594,I35351,I35339,I35639,I521432,I521414,I35656,I521426,I35682,I35690,I35333,I35721,I35738,I35755,I35772,I35789,I35354,I35820,I35342,I35336,I35892,I342098,I35918,I35935,I35943,I35960,I342101,I35977,I342122,I36003,I35884,I35875,I342110,I36048,I36056,I342113,I36073,I35872,I342119,I36113,I36121,I35878,I35866,I36166,I342116,I342104,I36183,I342107,I36209,I36217,I35860,I36248,I36265,I342125,I36282,I36299,I36316,I35881,I36347,I35869,I35863,I36419,I293879,I36445,I36462,I36470,I36487,I293876,I293870,I36504,I293864,I36530,I36411,I36402,I293852,I36575,I36583,I293861,I36600,I36399,I293858,I36640,I36648,I36405,I36393,I36693,I293855,I293873,I36710,I36736,I36744,I36387,I36775,I36792,I293867,I36809,I36826,I36843,I36408,I36874,I36396,I36390,I36946,I914342,I36972,I36989,I36997,I37014,I914330,I914321,I37031,I914318,I37057,I36938,I36929,I914324,I37102,I37110,I914336,I37127,I36926,I914333,I37167,I37175,I36932,I36920,I37220,I914327,I37237,I914339,I37263,I37271,I36914,I37302,I37319,I37336,I37353,I37370,I36935,I37401,I36923,I36917,I37473,I935728,I37499,I37516,I37524,I37541,I935716,I935707,I37558,I935704,I37584,I37465,I37456,I935710,I37629,I37637,I935722,I37654,I37453,I935719,I37694,I37702,I37459,I37447,I37747,I935713,I37764,I935725,I37790,I37798,I37441,I37829,I37846,I37863,I37880,I37897,I37462,I37928,I37450,I37444,I38000,I117050,I38026,I38043,I38051,I38068,I117053,I117035,I38085,I117041,I38111,I37992,I37983,I117044,I38156,I38164,I38181,I37980,I117056,I38221,I38229,I37986,I37974,I38274,I117059,I117047,I38291,I117038,I38317,I38325,I37968,I38356,I38373,I117062,I38390,I38407,I38424,I37989,I38455,I37977,I37971,I38527,I729059,I38553,I38570,I38578,I38595,I729035,I729062,I38612,I729047,I38638,I38519,I38510,I729053,I38683,I38691,I729038,I38708,I38507,I729056,I38748,I38756,I38513,I38501,I38801,I729041,I729044,I38818,I38844,I38852,I38495,I38883,I38900,I729050,I38917,I38934,I38951,I38516,I38982,I38504,I38498,I39054,I251192,I39080,I39097,I39105,I39122,I251189,I251183,I39139,I251177,I39165,I39046,I39037,I251165,I39210,I39218,I251174,I39235,I39034,I251171,I39275,I39283,I39040,I39028,I39328,I251168,I251186,I39345,I39371,I39379,I39022,I39410,I39427,I251180,I39444,I39461,I39478,I39043,I39509,I39031,I39025,I39581,I595404,I39607,I39624,I39632,I39649,I595419,I595422,I39666,I595401,I39692,I39573,I39564,I595407,I39737,I39745,I595413,I39762,I39561,I39802,I39810,I39567,I39555,I39855,I595416,I595398,I39872,I595410,I39898,I39906,I39549,I39937,I39954,I39971,I39988,I40005,I39570,I40036,I39558,I39552,I40108,I925902,I40134,I40151,I40159,I40176,I925890,I925881,I40193,I925878,I40219,I40100,I40091,I925884,I40264,I40272,I925896,I40289,I40088,I925893,I40329,I40337,I40094,I40082,I40382,I925887,I40399,I925899,I40425,I40433,I40076,I40464,I40481,I40498,I40515,I40532,I40097,I40563,I40085,I40079,I40635,I736165,I40661,I40678,I40686,I40703,I736141,I736168,I40720,I736153,I40746,I40627,I40618,I736159,I40791,I40799,I736144,I40816,I40615,I736162,I40856,I40864,I40621,I40609,I40909,I736147,I736150,I40926,I40952,I40960,I40603,I40991,I41008,I736156,I41025,I41042,I41059,I40624,I41090,I40612,I40606,I41162,I690777,I41188,I41205,I41213,I41230,I690768,I690789,I41247,I690771,I41273,I41154,I41145,I41318,I41326,I690786,I41343,I41142,I690780,I41383,I41391,I41148,I41136,I41436,I690774,I690783,I41453,I41479,I41487,I41130,I41518,I41535,I41552,I41569,I41586,I41151,I41617,I41139,I41133,I41689,I695520,I41715,I41732,I41740,I41757,I695511,I695532,I41774,I695514,I41800,I41681,I41672,I41845,I41853,I695529,I41870,I41669,I695523,I41910,I41918,I41675,I41663,I41963,I695517,I695526,I41980,I42006,I42014,I41657,I42045,I42062,I42079,I42096,I42113,I41678,I42144,I41666,I41660,I42216,I399686,I42242,I42259,I42267,I42284,I399692,I399680,I42301,I399677,I42327,I42208,I42199,I399689,I42372,I42380,I399683,I42397,I42196,I399701,I42437,I42445,I42202,I42190,I42490,I399695,I399698,I42507,I42533,I42541,I42184,I42572,I42589,I42606,I42623,I42640,I42205,I42671,I42193,I42187,I42743,I871570,I42769,I42786,I42794,I42811,I871558,I871549,I42828,I871546,I42854,I42735,I42726,I871552,I42899,I42907,I871564,I42924,I42723,I871561,I42964,I42972,I42729,I42717,I43017,I871555,I43034,I871567,I43060,I43068,I42711,I43099,I43116,I43133,I43150,I43167,I42732,I43198,I42720,I42714,I43270,I895846,I43296,I43313,I43321,I43338,I895834,I895825,I43355,I895822,I43381,I43262,I43253,I895828,I43426,I43434,I895840,I43451,I43250,I895837,I43491,I43499,I43256,I43244,I43544,I895831,I43561,I895843,I43587,I43595,I43238,I43626,I43643,I43660,I43677,I43694,I43259,I43725,I43247,I43241,I43797,I814177,I43823,I43840,I43848,I43865,I814171,I814192,I43882,I43908,I43789,I43780,I814174,I43953,I43961,I814183,I43978,I43777,I44018,I44026,I43783,I43771,I44071,I814189,I44088,I814180,I44114,I44122,I43765,I44153,I44170,I814186,I44187,I44204,I44221,I43786,I44252,I43774,I43768,I44324,I397901,I44350,I44367,I44375,I44392,I397907,I397895,I44409,I397892,I44435,I44316,I44307,I397904,I44480,I44488,I397898,I44505,I44304,I397916,I44545,I44553,I44310,I44298,I44598,I397910,I397913,I44615,I44641,I44649,I44292,I44680,I44697,I44714,I44731,I44748,I44313,I44779,I44301,I44295,I44851,I62740,I44877,I44894,I44902,I44919,I62755,I44936,I62758,I44962,I44843,I44834,I62752,I45007,I45015,I62761,I45032,I44831,I62737,I45072,I45080,I44837,I44825,I45125,I62743,I45142,I62746,I45168,I45176,I44819,I45207,I45224,I62749,I45241,I45258,I45275,I44840,I45306,I44828,I44822,I45378,I583266,I45404,I45421,I45429,I45446,I583281,I583284,I45463,I583263,I45489,I45370,I45361,I583269,I45534,I45542,I583275,I45559,I45358,I45599,I45607,I45364,I45352,I45652,I583278,I583260,I45669,I583272,I45695,I45703,I45346,I45734,I45751,I45768,I45785,I45802,I45367,I45833,I45355,I45349,I45905,I738749,I45931,I45948,I45956,I45973,I738725,I738752,I45990,I738737,I46016,I45897,I45888,I738743,I46061,I46069,I738728,I46086,I45885,I738746,I46126,I46134,I45891,I45879,I46179,I738731,I738734,I46196,I46222,I46230,I45873,I46261,I46278,I738740,I46295,I46312,I46329,I45894,I46360,I45882,I45876,I46432,I176547,I46458,I46466,I46483,I176541,I176535,I46500,I176556,I46526,I176553,I46543,I46551,I176550,I46568,I46400,I46599,I46616,I46412,I46656,I46421,I46678,I176538,I46695,I176559,I46721,I46738,I46424,I46760,I46409,I46791,I176544,I46808,I46825,I46842,I46418,I46873,I46406,I46415,I46403,I46959,I46985,I46993,I47010,I47027,I47053,I47070,I47078,I47095,I46927,I47126,I47143,I46939,I47183,I46948,I47205,I47222,I47248,I47265,I46951,I47287,I46936,I47318,I47335,I47352,I47369,I46945,I47400,I46933,I46942,I46930,I47486,I689723,I47512,I47520,I47537,I689720,I689735,I47554,I689717,I47580,I689714,I47597,I47605,I47622,I47454,I47653,I47670,I47466,I47710,I47475,I47732,I689729,I47749,I689732,I47775,I47792,I47478,I47814,I47463,I47845,I689726,I47862,I47879,I47896,I47472,I47927,I47460,I47469,I47457,I48013,I960292,I48039,I48047,I48064,I960286,I960307,I48081,I960298,I48107,I960289,I48124,I48132,I960301,I48149,I47981,I48180,I48197,I47993,I48237,I48002,I48259,I960310,I960295,I48276,I48302,I48319,I48005,I48341,I47990,I48372,I960304,I48389,I48406,I48423,I47999,I48454,I47987,I47996,I47984,I48540,I594832,I48566,I48574,I48591,I594823,I594841,I48608,I594820,I48634,I48651,I48659,I594826,I48676,I48508,I48707,I48724,I48520,I48764,I48529,I48786,I594838,I594829,I48803,I594844,I48829,I48846,I48532,I48868,I48517,I48899,I594835,I48916,I48933,I48950,I48526,I48981,I48514,I48523,I48511,I49067,I114081,I49093,I49101,I49118,I114078,I114060,I49135,I114066,I49161,I114075,I49178,I49186,I114069,I49203,I49035,I49234,I49251,I49047,I114084,I49291,I49056,I49313,I114072,I114063,I49330,I49356,I49373,I49059,I49395,I49044,I49426,I114087,I49443,I49460,I49477,I49053,I49508,I49041,I49050,I49038,I49594,I421100,I49620,I49628,I49645,I421121,I421115,I49662,I421097,I49688,I49705,I49713,I421109,I49730,I49562,I49761,I49778,I49574,I421106,I49818,I49583,I49840,I421112,I421103,I49857,I49883,I49900,I49586,I49922,I49571,I49953,I421118,I49970,I49987,I50004,I49580,I50035,I49568,I49577,I49565,I50121,I634388,I50147,I50155,I50172,I634385,I634400,I50189,I634382,I50215,I634379,I50232,I50240,I50257,I50089,I50288,I50305,I50101,I50345,I50110,I50367,I634394,I50384,I634397,I50410,I50427,I50113,I50449,I50098,I50480,I634391,I50497,I50514,I50531,I50107,I50562,I50095,I50104,I50092,I50648,I680764,I50674,I50682,I50699,I680761,I680776,I50716,I680758,I50742,I680755,I50759,I50767,I50784,I50616,I50815,I50832,I50628,I50872,I50637,I50894,I680770,I50911,I680773,I50937,I50954,I50640,I50976,I50625,I51007,I680767,I51024,I51041,I51058,I50634,I51089,I50622,I50631,I50619,I51175,I225896,I51201,I51209,I51226,I225878,I225893,I51243,I225869,I51269,I225872,I51286,I51294,I225887,I51311,I51143,I51342,I51359,I51155,I225890,I51399,I51164,I51421,I225881,I51438,I225875,I51464,I51481,I51167,I51503,I51152,I51534,I225884,I51551,I51568,I51585,I51161,I51616,I51149,I51158,I51146,I51702,I330148,I51728,I51736,I51753,I330142,I330133,I51770,I330154,I51796,I330136,I51813,I51821,I330130,I51838,I51670,I51869,I51886,I51682,I51926,I51691,I51948,I330157,I330139,I51965,I330145,I51991,I52008,I51694,I52030,I51679,I52061,I330151,I52078,I52095,I52112,I51688,I52143,I51676,I51685,I51673,I52229,I52255,I52263,I52280,I52297,I52323,I52340,I52348,I52365,I52197,I52396,I52413,I52209,I52453,I52218,I52475,I52492,I52518,I52535,I52221,I52557,I52206,I52588,I52605,I52622,I52639,I52215,I52670,I52203,I52212,I52200,I52756,I300730,I52782,I52790,I52807,I300712,I300727,I52824,I300703,I52850,I300706,I52867,I52875,I300721,I52892,I52724,I52923,I52940,I52736,I300724,I52980,I52745,I53002,I300715,I53019,I300709,I53045,I53062,I52748,I53084,I52733,I53115,I300718,I53132,I53149,I53166,I52742,I53197,I52730,I52739,I52727,I53283,I544546,I53309,I53317,I53334,I544537,I544555,I53351,I544534,I53377,I53394,I53402,I544540,I53419,I53251,I53450,I53467,I53263,I53507,I53272,I53529,I544552,I544543,I53546,I544558,I53572,I53589,I53275,I53611,I53260,I53642,I544549,I53659,I53676,I53693,I53269,I53724,I53257,I53266,I53254,I53810,I464779,I53836,I53844,I53861,I464791,I464776,I53878,I464770,I53904,I464785,I53921,I53929,I464773,I53946,I53778,I53977,I53994,I53790,I464782,I54034,I53799,I54056,I464788,I464794,I54073,I54099,I54116,I53802,I54138,I53787,I54169,I54186,I54203,I54220,I53796,I54251,I53784,I53793,I53781,I54337,I268056,I54363,I54371,I54388,I268038,I268053,I54405,I268029,I54431,I268032,I54448,I54456,I268047,I54473,I54305,I54504,I54521,I54317,I268050,I54561,I54326,I54583,I268041,I54600,I268035,I54626,I54643,I54329,I54665,I54314,I54696,I268044,I54713,I54730,I54747,I54323,I54778,I54311,I54320,I54308,I54864,I526050,I54890,I54898,I54915,I526041,I526059,I54932,I526038,I54958,I54975,I54983,I526044,I55000,I54832,I55031,I55048,I54844,I55088,I54853,I55110,I526056,I526047,I55127,I526062,I55153,I55170,I54856,I55192,I54841,I55223,I526053,I55240,I55257,I55274,I54850,I55305,I54838,I54847,I54835,I55391,I1079876,I55417,I55425,I55442,I1079870,I1079891,I55459,I1079867,I55485,I1079888,I55502,I55510,I1079885,I55527,I55359,I55558,I55575,I55371,I1079873,I55615,I55380,I55637,I1079882,I1079879,I55654,I1079864,I55680,I55697,I55383,I55719,I55368,I55750,I55767,I55784,I55801,I55377,I55832,I55365,I55374,I55362,I55918,I774910,I55944,I55952,I55969,I774928,I774922,I55986,I774901,I56012,I774919,I56029,I56037,I774904,I56054,I55886,I56085,I56102,I55898,I774916,I56142,I55907,I56164,I774925,I774913,I56181,I774907,I56207,I56224,I55910,I56246,I55895,I56277,I56294,I56311,I56328,I55904,I56359,I55892,I55901,I55889,I56445,I855368,I56471,I56479,I56496,I855383,I855362,I56513,I855365,I56539,I855386,I56556,I56564,I56581,I56413,I56612,I56629,I56425,I56669,I56434,I56691,I855374,I855371,I56708,I855377,I56734,I56751,I56437,I56773,I56422,I56804,I855380,I56821,I56838,I56855,I56431,I56886,I56419,I56428,I56416,I56972,I486743,I56998,I57006,I57023,I486755,I486740,I57040,I486734,I57066,I486749,I57083,I57091,I486737,I57108,I56940,I57139,I57156,I56952,I486746,I57196,I56961,I57218,I486752,I486758,I57235,I57261,I57278,I56964,I57300,I56949,I57331,I57348,I57365,I57382,I56958,I57413,I56946,I56955,I56943,I57499,I524316,I57525,I57533,I57550,I524307,I524325,I57567,I524304,I57593,I57610,I57618,I524310,I57635,I57467,I57666,I57683,I57479,I57723,I57488,I57745,I524322,I524313,I57762,I524328,I57788,I57805,I57491,I57827,I57476,I57858,I524319,I57875,I57892,I57909,I57485,I57940,I57473,I57482,I57470,I58026,I518536,I58052,I58060,I58077,I518527,I518545,I58094,I518524,I58120,I58137,I58145,I518530,I58162,I57994,I58193,I58210,I58006,I58250,I58015,I58272,I518542,I518533,I58289,I518548,I58315,I58332,I58018,I58354,I58003,I58385,I518539,I58402,I58419,I58436,I58012,I58467,I58000,I58009,I57997,I58553,I240652,I58579,I58587,I58604,I240634,I240649,I58621,I240625,I58647,I240628,I58664,I58672,I240643,I58689,I58521,I58720,I58737,I58533,I240646,I58777,I58542,I58799,I240637,I58816,I240631,I58842,I58859,I58545,I58881,I58530,I58912,I240640,I58929,I58946,I58963,I58539,I58994,I58527,I58536,I58524,I59080,I59106,I59114,I59131,I59148,I59174,I59191,I59199,I59216,I59048,I59247,I59264,I59060,I59304,I59069,I59326,I59343,I59369,I59386,I59072,I59408,I59057,I59439,I59456,I59473,I59490,I59066,I59521,I59054,I59063,I59051,I59607,I602924,I59633,I59641,I59658,I602915,I602933,I59675,I602912,I59701,I59718,I59726,I602918,I59743,I59575,I59774,I59791,I59587,I59831,I59596,I59853,I602930,I602921,I59870,I602936,I59896,I59913,I59599,I59935,I59584,I59966,I602927,I59983,I60000,I60017,I59593,I60048,I59581,I59590,I59578,I60134,I368772,I60160,I60168,I60185,I368766,I368757,I60202,I368778,I60228,I368760,I60245,I60253,I368754,I60270,I60102,I60301,I60318,I60114,I60358,I60123,I60380,I368781,I368763,I60397,I368769,I60423,I60440,I60126,I60462,I60111,I60493,I368775,I60510,I60527,I60544,I60120,I60575,I60108,I60117,I60105,I60661,I829936,I60687,I60695,I60712,I829951,I829930,I60729,I829933,I60755,I829954,I60772,I60780,I60797,I60629,I60828,I60845,I60641,I60885,I60650,I60907,I829942,I829939,I60924,I829945,I60950,I60967,I60653,I60989,I60638,I61020,I829948,I61037,I61054,I61071,I60647,I61102,I60635,I60644,I60632,I61188,I355172,I61214,I61222,I61239,I355166,I355157,I61256,I355178,I61282,I355160,I61299,I61307,I355154,I61324,I61156,I61355,I61372,I61168,I61412,I61177,I61434,I355181,I355163,I61451,I355169,I61477,I61494,I61180,I61516,I61165,I61547,I355175,I61564,I61581,I61598,I61174,I61629,I61162,I61171,I61159,I61715,I61741,I61749,I61766,I61783,I61809,I61826,I61834,I61851,I61683,I61882,I61899,I61695,I61939,I61704,I61961,I61978,I62004,I62021,I61707,I62043,I61692,I62074,I62091,I62108,I62125,I61701,I62156,I61689,I61698,I61686,I62242,I847276,I62268,I62276,I62293,I847291,I847270,I62310,I847273,I62336,I847294,I62353,I62361,I62378,I62210,I62409,I62426,I62222,I62466,I62231,I62488,I847282,I847279,I62505,I847285,I62531,I62548,I62234,I62570,I62219,I62601,I847288,I62618,I62635,I62652,I62228,I62683,I62216,I62225,I62213,I62769,I844964,I62795,I62803,I62820,I844979,I844958,I62837,I844961,I62863,I844982,I62880,I62888,I62905,I62936,I62953,I62993,I63015,I844970,I844967,I63032,I844973,I63058,I63075,I63097,I63128,I844976,I63145,I63162,I63179,I63210,I63296,I63322,I63330,I63347,I63364,I63390,I63407,I63415,I63432,I63264,I63463,I63480,I63276,I63520,I63285,I63542,I63559,I63585,I63602,I63288,I63624,I63273,I63655,I63672,I63689,I63706,I63282,I63737,I63270,I63279,I63267,I63823,I465935,I63849,I63857,I63874,I465947,I465932,I63891,I465926,I63917,I465941,I63934,I63942,I465929,I63959,I63791,I63990,I64007,I63803,I465938,I64047,I63812,I64069,I465944,I465950,I64086,I64112,I64129,I63815,I64151,I63800,I64182,I64199,I64216,I64233,I63809,I64264,I63797,I63806,I63794,I64350,I244341,I64376,I64384,I64401,I244323,I244338,I64418,I244314,I64444,I244317,I64461,I64469,I244332,I64486,I64318,I64517,I64534,I64330,I244335,I64574,I64339,I64596,I244326,I64613,I244320,I64639,I64656,I64342,I64678,I64327,I64709,I244329,I64726,I64743,I64760,I64336,I64791,I64324,I64333,I64321,I64877,I605236,I64903,I64911,I64928,I605227,I605245,I64945,I605224,I64971,I64988,I64996,I605230,I65013,I64845,I65044,I65061,I64857,I65101,I64866,I65123,I605242,I605233,I65140,I605248,I65166,I65183,I64869,I65205,I64854,I65236,I605239,I65253,I65270,I65287,I64863,I65318,I64851,I64860,I64848,I65404,I438191,I65430,I65438,I65455,I438203,I438188,I65472,I438182,I65498,I438197,I65515,I65523,I438185,I65540,I65372,I65571,I65588,I65384,I438194,I65628,I65393,I65650,I438200,I438206,I65667,I65693,I65710,I65396,I65732,I65381,I65763,I65780,I65797,I65814,I65390,I65845,I65378,I65387,I65375,I65931,I394920,I65957,I65965,I65982,I394941,I394935,I65999,I394917,I66025,I66042,I66050,I394929,I66067,I65899,I66098,I66115,I65911,I394926,I66155,I65920,I66177,I394932,I394923,I66194,I66220,I66237,I65923,I66259,I65908,I66290,I394938,I66307,I66324,I66341,I65917,I66372,I65905,I65914,I65902,I66458,I586162,I66484,I66492,I66509,I586153,I586171,I66526,I586150,I66552,I66569,I66577,I586156,I66594,I66426,I66625,I66642,I66438,I66682,I66447,I66704,I586168,I586159,I66721,I586174,I66747,I66764,I66450,I66786,I66435,I66817,I586165,I66834,I66851,I66868,I66444,I66899,I66432,I66441,I66429,I66985,I1043581,I67011,I67019,I67036,I1043575,I1043596,I67053,I1043572,I67079,I1043593,I67096,I67104,I1043590,I67121,I66953,I67152,I67169,I66965,I1043578,I67209,I66974,I67231,I1043587,I1043584,I67248,I1043569,I67274,I67291,I66977,I67313,I66962,I67344,I67361,I67378,I67395,I66971,I67426,I66959,I66968,I66956,I67512,I406225,I67538,I67546,I67563,I406246,I406240,I67580,I406222,I67606,I67623,I67631,I406234,I67648,I67480,I67679,I67696,I67492,I406231,I67736,I67501,I67758,I406237,I406228,I67775,I67801,I67818,I67504,I67840,I67489,I67871,I406243,I67888,I67905,I67922,I67498,I67953,I67486,I67495,I67483,I68039,I919526,I68065,I68073,I68090,I919541,I919520,I68107,I919523,I68133,I919544,I68150,I68158,I68175,I68007,I68206,I68223,I68019,I68263,I68028,I68285,I919532,I919529,I68302,I919535,I68328,I68345,I68031,I68367,I68016,I68398,I919538,I68415,I68432,I68449,I68025,I68480,I68013,I68022,I68010,I68566,I958660,I68592,I68600,I68617,I958654,I958675,I68634,I958666,I68660,I958657,I68677,I68685,I958669,I68702,I68534,I68733,I68750,I68546,I68790,I68555,I68812,I958678,I958663,I68829,I68855,I68872,I68558,I68894,I68543,I68925,I958672,I68942,I68959,I68976,I68552,I69007,I68540,I68549,I68537,I69093,I797905,I69119,I69127,I69144,I797902,I797908,I69161,I69187,I69204,I69212,I69229,I69260,I69277,I797911,I69317,I69339,I797914,I797923,I69356,I797917,I69382,I69399,I69421,I69452,I797920,I69469,I69486,I69503,I69534,I69620,I1032871,I69646,I69654,I69671,I1032865,I1032886,I69688,I1032862,I69714,I1032883,I69731,I69739,I1032880,I69756,I69588,I69787,I69804,I69600,I1032868,I69844,I69609,I69866,I1032877,I1032874,I69883,I1032859,I69909,I69926,I69612,I69948,I69597,I69979,I69996,I70013,I70030,I69606,I70061,I69594,I69603,I69591,I70147,I1000155,I70173,I70181,I70198,I1000158,I1000152,I70215,I1000149,I70241,I1000134,I70258,I70266,I1000143,I70283,I70115,I70314,I70331,I70127,I70371,I70136,I70393,I1000137,I1000140,I70410,I1000146,I70436,I70453,I70139,I70475,I70124,I70506,I70523,I70540,I70557,I70133,I70588,I70121,I70130,I70118,I70674,I348644,I70700,I70708,I70725,I348638,I348629,I70742,I348650,I70768,I348632,I70785,I70793,I348626,I70810,I70642,I70841,I70858,I70654,I70898,I70663,I70920,I348653,I348635,I70937,I348641,I70963,I70980,I70666,I71002,I70651,I71033,I348647,I71050,I71067,I71084,I70660,I71115,I70648,I70657,I70645,I71201,I809125,I71227,I71235,I71252,I809122,I809128,I71269,I71295,I71312,I71320,I71337,I71169,I71368,I71385,I71181,I809131,I71425,I71190,I71447,I809134,I809143,I71464,I809137,I71490,I71507,I71193,I71529,I71178,I71560,I809140,I71577,I71594,I71611,I71187,I71642,I71175,I71184,I71172,I71728,I139062,I71754,I71762,I71779,I139056,I139050,I71796,I139071,I71822,I139068,I71839,I71847,I139065,I71864,I71696,I71895,I71912,I71708,I71952,I71717,I71974,I139053,I71991,I139074,I72017,I72034,I71720,I72056,I71705,I72087,I139059,I72104,I72121,I72138,I71714,I72169,I71702,I71711,I71699,I72255,I1001889,I72281,I72289,I72306,I1001892,I1001886,I72323,I1001883,I72349,I1001868,I72366,I72374,I1001877,I72391,I72223,I72422,I72439,I72235,I72479,I72244,I72501,I1001871,I1001874,I72518,I1001880,I72544,I72561,I72247,I72583,I72232,I72614,I72631,I72648,I72665,I72241,I72696,I72229,I72238,I72226,I72782,I283866,I72808,I72816,I72833,I283848,I283863,I72850,I283839,I72876,I283842,I72893,I72901,I283857,I72918,I72750,I72949,I72966,I72762,I283860,I73006,I72771,I73028,I283851,I73045,I283845,I73071,I73088,I72774,I73110,I72759,I73141,I283854,I73158,I73175,I73192,I72768,I73223,I72756,I72765,I72753,I73309,I703204,I73335,I73343,I73360,I703222,I703216,I73377,I703195,I73403,I703213,I73420,I73428,I703198,I73445,I73277,I73476,I73493,I73289,I703210,I73533,I73298,I73555,I703219,I703207,I73572,I703201,I73598,I73615,I73301,I73637,I73286,I73668,I73685,I73702,I73719,I73295,I73750,I73283,I73292,I73280,I73836,I1027674,I73862,I73870,I73887,I1027680,I1027698,I73904,I1027695,I73930,I1027692,I73947,I73955,I1027686,I73972,I73804,I74003,I74020,I73816,I74060,I73825,I74082,I1027689,I1027677,I74099,I1027701,I74125,I74142,I73828,I74164,I73813,I74195,I1027683,I74212,I74229,I74246,I73822,I74277,I73810,I73819,I73807,I74363,I865772,I74389,I74397,I74414,I865787,I865766,I74431,I865769,I74457,I865790,I74474,I74482,I74499,I74530,I74547,I74587,I74609,I865778,I865775,I74626,I865781,I74652,I74669,I74691,I74722,I865784,I74739,I74756,I74773,I74804,I74890,I402655,I74916,I74924,I74941,I402676,I402670,I74958,I402652,I74984,I75001,I75009,I402664,I75026,I74858,I75057,I75074,I74870,I402661,I75114,I74879,I75136,I402667,I402658,I75153,I75179,I75196,I74882,I75218,I74867,I75249,I402673,I75266,I75283,I75300,I74876,I75331,I74864,I74873,I74861,I75417,I758114,I75443,I75451,I75468,I758132,I758126,I75485,I758105,I75511,I758123,I75528,I75536,I758108,I75553,I75385,I75584,I75601,I75397,I758120,I75641,I75406,I75663,I758129,I758117,I75680,I758111,I75706,I75723,I75409,I75745,I75394,I75776,I75793,I75810,I75827,I75403,I75858,I75391,I75400,I75388,I75944,I75970,I75978,I75995,I76012,I76038,I76055,I76063,I76080,I75912,I76111,I76128,I75924,I76168,I75933,I76190,I76207,I76233,I76250,I75936,I76272,I75921,I76303,I76320,I76337,I76354,I75930,I76385,I75918,I75927,I75915,I76471,I806881,I76497,I76505,I76522,I806878,I806884,I76539,I76565,I76582,I76590,I76607,I76439,I76638,I76655,I76451,I806887,I76695,I76460,I76717,I806890,I806899,I76734,I806893,I76760,I76777,I76463,I76799,I76448,I76830,I806896,I76847,I76864,I76881,I76457,I76912,I76445,I76454,I76442,I76998,I379108,I77024,I77032,I77049,I379102,I379093,I77066,I379114,I77092,I379096,I77109,I77117,I379090,I77134,I76966,I77165,I77182,I76978,I77222,I76987,I77244,I379117,I379099,I77261,I379105,I77287,I77304,I76990,I77326,I76975,I77357,I379111,I77374,I77391,I77408,I76984,I77439,I76972,I76981,I76969,I77525,I600612,I77551,I77559,I77576,I600603,I600621,I77593,I600600,I77619,I77636,I77644,I600606,I77661,I77493,I77692,I77709,I77505,I77749,I77514,I77771,I600618,I600609,I77788,I600624,I77814,I77831,I77517,I77853,I77502,I77884,I600615,I77901,I77918,I77935,I77511,I77966,I77499,I77508,I77496,I78052,I657049,I78078,I78086,I78103,I657046,I657061,I78120,I657043,I78146,I657040,I78163,I78171,I78188,I78020,I78219,I78236,I78032,I78276,I78041,I78298,I657055,I78315,I657058,I78341,I78358,I78044,I78380,I78029,I78411,I657052,I78428,I78445,I78462,I78038,I78493,I78026,I78035,I78023,I78579,I502930,I78605,I78613,I78630,I502921,I502939,I78647,I502918,I78673,I78690,I78698,I502924,I78715,I78547,I78746,I78763,I78559,I78803,I78568,I78825,I502936,I502927,I78842,I502942,I78868,I78885,I78571,I78907,I78556,I78938,I502933,I78955,I78972,I78989,I78565,I79020,I78553,I78562,I78550,I79106,I563620,I79132,I79140,I79157,I563611,I563629,I79174,I563608,I79200,I79217,I79225,I563614,I79242,I79273,I79290,I79330,I79352,I563626,I563617,I79369,I563632,I79395,I79412,I79434,I79465,I563623,I79482,I79499,I79516,I79547,I79633,I262786,I79659,I79667,I79684,I262768,I262783,I79701,I262759,I79727,I262762,I79744,I79752,I262777,I79769,I79601,I79800,I79817,I79613,I262780,I79857,I79622,I79879,I262771,I79896,I262765,I79922,I79939,I79625,I79961,I79610,I79992,I262774,I80009,I80026,I80043,I79619,I80074,I79607,I79616,I79604,I80160,I321444,I80186,I80194,I80211,I321438,I321429,I80228,I321450,I80254,I321432,I80271,I80279,I321426,I80296,I80128,I80327,I80344,I80140,I80384,I80149,I80406,I321453,I321435,I80423,I321441,I80449,I80466,I80152,I80488,I80137,I80519,I321447,I80536,I80553,I80570,I80146,I80601,I80134,I80143,I80131,I80687,I144417,I80713,I80721,I80738,I144411,I144405,I80755,I144426,I80781,I144423,I80798,I80806,I144420,I80823,I80655,I80854,I80871,I80667,I80911,I80676,I80933,I144408,I80950,I144429,I80976,I80993,I80679,I81015,I80664,I81046,I144414,I81063,I81080,I81097,I80673,I81128,I80661,I80670,I80658,I81214,I400275,I81240,I81248,I81265,I400296,I400290,I81282,I400272,I81308,I81325,I81333,I400284,I81350,I81182,I81381,I81398,I81194,I400281,I81438,I81203,I81460,I400287,I400278,I81477,I81503,I81520,I81206,I81542,I81191,I81573,I400293,I81590,I81607,I81624,I81200,I81655,I81188,I81197,I81185,I81741,I745840,I81767,I81775,I81792,I745858,I745852,I81809,I745831,I81835,I745849,I81852,I81860,I745834,I81877,I81709,I81908,I81925,I81721,I745846,I81965,I81730,I81987,I745855,I745843,I82004,I745837,I82030,I82047,I81733,I82069,I81718,I82100,I82117,I82134,I82151,I81727,I82182,I81715,I81724,I81712,I82268,I237490,I82294,I82302,I82319,I237472,I237487,I82336,I237463,I82362,I237466,I82379,I82387,I237481,I82404,I82236,I82435,I82452,I82248,I237484,I82492,I82257,I82514,I237475,I82531,I237469,I82557,I82574,I82260,I82596,I82245,I82627,I237478,I82644,I82661,I82678,I82254,I82709,I82242,I82251,I82239,I82795,I903920,I82821,I82829,I82846,I903935,I903914,I82863,I903917,I82889,I903938,I82906,I82914,I82931,I82763,I82962,I82979,I82775,I83019,I82784,I83041,I903926,I903923,I83058,I903929,I83084,I83101,I82787,I83123,I82772,I83154,I903932,I83171,I83188,I83205,I82781,I83236,I82769,I82778,I82766,I83322,I500618,I83348,I83356,I83373,I500609,I500627,I83390,I500606,I83416,I83433,I83441,I500612,I83458,I83290,I83489,I83506,I83302,I83546,I83311,I83568,I500624,I500615,I83585,I500630,I83611,I83628,I83314,I83650,I83299,I83681,I500621,I83698,I83715,I83732,I83308,I83763,I83296,I83305,I83293,I83849,I822028,I83875,I83883,I83900,I822025,I822031,I83917,I83943,I83960,I83968,I83985,I83817,I84016,I84033,I83829,I822034,I84073,I83838,I84095,I822037,I822046,I84112,I822040,I84138,I84155,I83841,I84177,I83826,I84208,I822043,I84225,I84242,I84259,I83835,I84290,I83823,I83832,I83820,I84376,I172977,I84402,I84410,I84427,I172971,I172965,I84444,I172986,I84470,I172983,I84487,I84495,I172980,I84512,I84344,I84543,I84560,I84356,I84600,I84365,I84622,I172968,I84639,I172989,I84665,I84682,I84368,I84704,I84353,I84735,I172974,I84752,I84769,I84786,I84362,I84817,I84350,I84359,I84347,I84903,I1023747,I84929,I84937,I84954,I1023753,I1023771,I84971,I1023768,I84997,I1023765,I85014,I85022,I1023759,I85039,I84871,I85070,I85087,I84883,I85127,I84892,I85149,I1023762,I1023750,I85166,I1023774,I85192,I85209,I84895,I85231,I84880,I85262,I1023756,I85279,I85296,I85313,I84889,I85344,I84877,I84886,I84874,I85430,I797344,I85456,I85464,I85481,I797341,I797347,I85498,I85524,I85541,I85549,I85566,I85398,I85597,I85614,I85410,I797350,I85654,I85419,I85676,I797353,I797362,I85693,I797356,I85719,I85736,I85422,I85758,I85407,I85789,I797359,I85806,I85823,I85840,I85416,I85871,I85404,I85413,I85401,I85957,I617374,I85983,I85991,I86008,I617365,I617383,I86025,I617362,I86051,I86068,I86076,I617368,I86093,I85925,I86124,I86141,I85937,I86181,I85946,I86203,I617380,I617371,I86220,I617386,I86246,I86263,I85949,I86285,I85934,I86316,I617377,I86333,I86350,I86367,I85943,I86398,I85931,I85940,I85928,I86484,I966820,I86510,I86518,I86535,I966814,I966835,I86552,I966826,I86578,I966817,I86595,I86603,I966829,I86620,I86452,I86651,I86668,I86464,I86708,I86473,I86730,I966838,I966823,I86747,I86773,I86790,I86476,I86812,I86461,I86843,I966832,I86860,I86877,I86894,I86470,I86925,I86458,I86467,I86455,I87011,I243287,I87037,I87045,I87062,I243269,I243284,I87079,I243260,I87105,I243263,I87122,I87130,I243278,I87147,I86979,I87178,I87195,I86991,I243281,I87235,I87000,I87257,I243272,I87274,I243266,I87300,I87317,I87003,I87339,I86988,I87370,I243275,I87387,I87404,I87421,I86997,I87452,I86985,I86994,I86982,I87538,I367684,I87564,I87572,I87589,I367678,I367669,I87606,I367690,I87632,I367672,I87649,I87657,I367666,I87674,I87506,I87705,I87722,I87518,I87762,I87527,I87784,I367693,I367675,I87801,I367681,I87827,I87844,I87530,I87866,I87515,I87897,I367687,I87914,I87931,I87948,I87524,I87979,I87512,I87521,I87509,I88065,I608126,I88091,I88099,I88116,I608117,I608135,I88133,I608114,I88159,I88176,I88184,I608120,I88201,I88033,I88232,I88249,I88045,I88289,I88054,I88311,I608132,I608123,I88328,I608138,I88354,I88371,I88057,I88393,I88042,I88424,I608129,I88441,I88458,I88475,I88051,I88506,I88039,I88048,I88036,I88592,I860570,I88618,I88626,I88643,I860585,I860564,I88660,I860567,I88686,I860588,I88703,I88711,I88728,I88560,I88759,I88776,I88572,I88816,I88581,I88838,I860576,I860573,I88855,I860579,I88881,I88898,I88584,I88920,I88569,I88951,I860582,I88968,I88985,I89002,I88578,I89033,I88566,I88575,I88563,I89119,I658103,I89145,I89153,I89170,I658100,I658115,I89187,I658097,I89213,I658094,I89230,I89238,I89255,I89087,I89286,I89303,I89099,I89343,I89108,I89365,I658109,I89382,I658112,I89408,I89425,I89111,I89447,I89096,I89478,I658106,I89495,I89512,I89529,I89105,I89560,I89093,I89102,I89090,I89646,I809686,I89672,I89680,I89697,I809683,I809689,I89714,I89740,I89757,I89765,I89782,I89614,I89813,I89830,I89626,I809692,I89870,I89635,I89892,I809695,I809704,I89909,I809698,I89935,I89952,I89638,I89974,I89623,I90005,I809701,I90022,I90039,I90056,I89632,I90087,I89620,I89629,I89617,I90173,I167027,I90199,I90207,I90224,I167021,I167015,I90241,I167036,I90267,I167033,I90284,I90292,I167030,I90309,I90141,I90340,I90357,I90153,I90397,I90162,I90419,I167018,I90436,I167039,I90462,I90479,I90165,I90501,I90150,I90532,I167024,I90549,I90566,I90583,I90159,I90614,I90147,I90156,I90144,I90700,I325252,I90726,I90734,I90751,I325246,I325237,I90768,I325258,I90794,I325240,I90811,I90819,I325234,I90836,I90668,I90867,I90884,I90680,I90924,I90689,I90946,I325261,I325243,I90963,I325249,I90989,I91006,I90692,I91028,I90677,I91059,I325255,I91076,I91093,I91110,I90686,I91141,I90674,I90683,I90671,I91227,I258570,I91253,I91261,I91278,I258552,I258567,I91295,I258543,I91321,I258546,I91338,I91346,I258561,I91363,I91195,I91394,I91411,I91207,I258564,I91451,I91216,I91473,I258555,I91490,I258549,I91516,I91533,I91219,I91555,I91204,I91586,I258558,I91603,I91620,I91637,I91213,I91668,I91201,I91210,I91198,I91754,I725814,I91780,I91788,I91805,I725832,I725826,I91822,I725805,I91848,I725823,I91865,I91873,I725808,I91890,I91722,I91921,I91938,I91734,I725820,I91978,I91743,I92000,I725829,I725817,I92017,I725811,I92043,I92060,I91746,I92082,I91731,I92113,I92130,I92147,I92164,I91740,I92195,I91728,I91737,I91725,I92281,I149772,I92307,I92315,I92332,I149766,I149760,I92349,I149781,I92375,I149778,I92392,I92400,I149775,I92417,I92249,I92448,I92465,I92261,I92505,I92270,I92527,I149763,I92544,I149784,I92570,I92587,I92273,I92609,I92258,I92640,I149769,I92657,I92674,I92691,I92267,I92722,I92255,I92264,I92252,I92808,I1082256,I92834,I92842,I92859,I1082250,I1082271,I92876,I1082247,I92902,I1082268,I92919,I92927,I1082265,I92944,I92776,I92975,I92992,I92788,I1082253,I93032,I92797,I93054,I1082262,I1082259,I93071,I1082244,I93097,I93114,I92800,I93136,I92785,I93167,I93184,I93201,I93218,I92794,I93249,I92782,I92791,I92779,I93335,I621213,I93361,I93369,I93386,I621210,I621225,I93403,I621207,I93429,I621204,I93446,I93454,I93471,I93502,I93519,I93559,I93581,I621219,I93598,I621222,I93624,I93641,I93663,I93694,I621216,I93711,I93728,I93745,I93776,I93862,I1051911,I93888,I93896,I93913,I1051905,I1051926,I93930,I1051902,I93956,I1051923,I93973,I93981,I1051920,I93998,I93830,I94029,I94046,I93842,I1051908,I94086,I93851,I94108,I1051917,I1051914,I94125,I1051899,I94151,I94168,I93854,I94190,I93839,I94221,I94238,I94255,I94272,I93848,I94303,I93836,I93845,I93833,I94389,I219045,I94415,I94423,I94440,I219027,I219042,I94457,I219018,I94483,I219021,I94500,I94508,I219036,I94525,I94357,I94556,I94573,I94369,I219039,I94613,I94378,I94635,I219030,I94652,I219024,I94678,I94695,I94381,I94717,I94366,I94748,I219033,I94765,I94782,I94799,I94375,I94830,I94363,I94372,I94360,I94916,I215883,I94942,I94950,I94967,I215865,I215880,I94984,I215856,I95010,I215859,I95027,I95035,I215874,I95052,I94884,I95083,I95100,I94896,I215877,I95140,I94905,I95162,I215868,I95179,I215862,I95205,I95222,I94908,I95244,I94893,I95275,I215871,I95292,I95309,I95326,I94902,I95357,I94890,I94899,I94887,I95443,I407415,I95469,I95477,I95494,I407436,I407430,I95511,I407412,I95537,I95554,I95562,I407424,I95579,I95411,I95610,I95627,I95423,I407421,I95667,I95432,I95689,I407427,I407418,I95706,I95732,I95749,I95435,I95771,I95420,I95802,I407433,I95819,I95836,I95853,I95429,I95884,I95417,I95426,I95414,I95970,I938600,I95996,I96004,I96021,I938615,I938594,I96038,I938597,I96064,I938618,I96081,I96089,I96106,I95938,I96137,I96154,I95950,I96194,I95959,I96216,I938606,I938603,I96233,I938609,I96259,I96276,I95962,I96298,I95947,I96329,I938612,I96346,I96363,I96380,I95956,I96411,I95944,I95953,I95941,I96497,I193207,I96523,I96531,I96548,I193201,I193195,I96565,I193216,I96591,I193213,I96608,I96616,I193210,I96633,I96465,I96664,I96681,I96477,I96721,I96486,I96743,I193198,I96760,I193219,I96786,I96803,I96489,I96825,I96474,I96856,I193204,I96873,I96890,I96907,I96483,I96938,I96471,I96480,I96468,I97024,I983684,I97050,I97058,I97075,I983678,I983699,I97092,I983690,I97118,I983681,I97135,I97143,I983693,I97160,I96992,I97191,I97208,I97004,I97248,I97013,I97270,I983702,I983687,I97287,I97313,I97330,I97016,I97352,I97001,I97383,I983696,I97400,I97417,I97434,I97010,I97465,I96998,I97007,I96995,I97551,I515646,I97577,I97585,I97602,I515637,I515655,I97619,I515634,I97645,I97662,I97670,I515640,I97687,I97519,I97718,I97735,I97531,I97775,I97540,I97797,I515652,I515643,I97814,I515658,I97840,I97857,I97543,I97879,I97528,I97910,I515649,I97927,I97944,I97961,I97537,I97992,I97525,I97534,I97522,I98078,I863460,I98104,I98112,I98129,I863475,I863454,I98146,I863457,I98172,I863478,I98189,I98197,I98214,I98046,I98245,I98262,I98058,I98302,I98067,I98324,I863466,I863463,I98341,I863469,I98367,I98384,I98070,I98406,I98055,I98437,I863472,I98454,I98471,I98488,I98064,I98519,I98052,I98061,I98049,I98605,I421695,I98631,I98639,I98656,I421716,I421710,I98673,I421692,I98699,I98716,I98724,I421704,I98741,I98573,I98772,I98789,I98585,I421701,I98829,I98594,I98851,I421707,I421698,I98868,I98894,I98911,I98597,I98933,I98582,I98964,I421713,I98981,I98998,I99015,I98591,I99046,I98579,I98588,I98576,I99132,I549748,I99158,I99166,I99183,I549739,I549757,I99200,I549736,I99226,I99243,I99251,I549742,I99268,I99100,I99299,I99316,I99112,I99356,I99121,I99378,I549754,I549745,I99395,I549760,I99421,I99438,I99124,I99460,I99109,I99491,I549751,I99508,I99525,I99542,I99118,I99573,I99106,I99115,I99103,I99659,I99685,I99693,I99710,I99727,I99753,I99770,I99778,I99795,I99627,I99826,I99843,I99639,I99883,I99648,I99905,I99922,I99948,I99965,I99651,I99987,I99636,I100018,I100035,I100052,I100069,I99645,I100100,I99633,I99642,I99630,I100186,I599456,I100212,I100220,I100237,I599447,I599465,I100254,I599444,I100280,I100297,I100305,I599450,I100322,I100154,I100353,I100370,I100166,I100410,I100175,I100432,I599462,I599453,I100449,I599468,I100475,I100492,I100178,I100514,I100163,I100545,I599459,I100562,I100579,I100596,I100172,I100627,I100160,I100169,I100157,I100713,I1092371,I100739,I100747,I100764,I1092365,I1092386,I100781,I1092362,I100807,I1092383,I100824,I100832,I1092380,I100849,I100681,I100880,I100897,I100693,I1092368,I100937,I100702,I100959,I1092377,I1092374,I100976,I1092359,I101002,I101019,I100705,I101041,I100690,I101072,I101089,I101106,I101123,I100699,I101154,I100687,I100696,I100684,I101240,I903342,I101266,I101274,I101291,I903357,I903336,I101308,I903339,I101334,I903360,I101351,I101359,I101376,I101208,I101407,I101424,I101220,I101464,I101229,I101486,I903348,I903345,I101503,I903351,I101529,I101546,I101232,I101568,I101217,I101599,I903354,I101616,I101633,I101650,I101226,I101681,I101214,I101223,I101211,I101767,I1086421,I101793,I101801,I101818,I1086415,I1086436,I101835,I1086412,I101861,I1086433,I101878,I101886,I1086430,I101903,I101735,I101934,I101951,I101747,I1086418,I101991,I101756,I102013,I1086427,I1086424,I102030,I1086409,I102056,I102073,I101759,I102095,I101744,I102126,I102143,I102160,I102177,I101753,I102208,I101741,I101750,I101738,I102294,I1045961,I102320,I102328,I102345,I1045955,I1045976,I102362,I1045952,I102388,I1045973,I102405,I102413,I1045970,I102430,I102262,I102461,I102478,I102274,I1045958,I102518,I102283,I102540,I1045967,I1045964,I102557,I1045949,I102583,I102600,I102286,I102622,I102271,I102653,I102670,I102687,I102704,I102280,I102735,I102268,I102277,I102265,I102821,I467091,I102847,I102855,I102872,I467103,I467088,I102889,I467082,I102915,I467097,I102932,I102940,I467085,I102957,I102789,I102988,I103005,I102801,I467094,I103045,I102810,I103067,I467100,I467106,I103084,I103110,I103127,I102813,I103149,I102798,I103180,I103197,I103214,I103231,I102807,I103262,I102795,I102804,I102792,I103348,I178927,I103374,I103382,I103399,I178921,I178915,I103416,I178936,I103442,I178933,I103459,I103467,I178930,I103484,I103316,I103515,I103532,I103328,I103572,I103337,I103594,I178918,I103611,I178939,I103637,I103654,I103340,I103676,I103325,I103707,I178924,I103724,I103741,I103758,I103334,I103789,I103322,I103331,I103319,I103875,I696574,I103901,I103909,I103926,I696571,I696586,I103943,I696568,I103969,I696565,I103986,I103994,I104011,I103843,I104042,I104059,I103855,I104099,I103864,I104121,I696580,I104138,I696583,I104164,I104181,I103867,I104203,I103852,I104234,I696577,I104251,I104268,I104285,I103861,I104316,I103849,I103858,I103846,I104402,I104428,I104436,I104453,I104470,I104496,I104513,I104521,I104538,I104370,I104569,I104586,I104382,I104626,I104391,I104648,I104665,I104691,I104708,I104394,I104730,I104379,I104761,I104778,I104795,I104812,I104388,I104843,I104376,I104385,I104373,I104929,I1026552,I104955,I104963,I104980,I1026558,I1026576,I104997,I1026573,I105023,I1026570,I105040,I105048,I1026564,I105065,I104897,I105096,I105113,I104909,I105153,I104918,I105175,I1026567,I1026555,I105192,I1026579,I105218,I105235,I104921,I105257,I104906,I105288,I1026561,I105305,I105322,I105339,I104915,I105370,I104903,I104912,I104900,I105456,I785246,I105482,I105490,I105507,I785264,I785258,I105524,I785237,I105550,I785255,I105567,I105575,I785240,I105592,I105424,I105623,I105640,I105436,I785252,I105680,I105445,I105702,I785261,I785249,I105719,I785243,I105745,I105762,I105448,I105784,I105433,I105815,I105832,I105849,I105866,I105442,I105897,I105430,I105439,I105427,I105983,I285974,I106009,I106017,I106034,I285956,I285971,I106051,I285947,I106077,I285950,I106094,I106102,I285965,I106119,I105951,I106150,I106167,I105963,I285968,I106207,I105972,I106229,I285959,I106246,I285953,I106272,I106289,I105975,I106311,I105960,I106342,I285962,I106359,I106376,I106393,I105969,I106424,I105957,I105966,I105954,I106510,I149177,I106536,I106544,I106561,I149171,I149165,I106578,I149186,I106604,I149183,I106621,I106629,I149180,I106646,I106478,I106677,I106694,I106490,I106734,I106499,I106756,I149168,I106773,I149189,I106799,I106816,I106502,I106838,I106487,I106869,I149174,I106886,I106903,I106920,I106496,I106951,I106484,I106493,I106481,I107037,I902764,I107063,I107071,I107088,I902779,I902758,I107105,I902761,I107131,I902782,I107148,I107156,I107173,I107005,I107204,I107221,I107017,I107261,I107026,I107283,I902770,I902767,I107300,I902773,I107326,I107343,I107029,I107365,I107014,I107396,I902776,I107413,I107430,I107447,I107023,I107478,I107011,I107020,I107008,I107564,I408010,I107590,I107598,I107615,I408031,I408025,I107632,I408007,I107658,I107675,I107683,I408019,I107700,I107532,I107731,I107748,I107544,I408016,I107788,I107553,I107810,I408022,I408013,I107827,I107853,I107870,I107556,I107892,I107541,I107923,I408028,I107940,I107957,I107974,I107550,I108005,I107538,I107547,I107535,I108091,I584428,I108117,I108125,I108142,I584419,I584437,I108159,I584416,I108185,I108202,I108210,I584422,I108227,I108059,I108258,I108275,I108071,I108315,I108080,I108337,I584434,I584425,I108354,I584440,I108380,I108397,I108083,I108419,I108068,I108450,I584431,I108467,I108484,I108501,I108077,I108532,I108065,I108074,I108062,I108618,I820906,I108644,I108652,I108669,I820903,I820909,I108686,I108712,I108729,I108737,I108754,I108586,I108785,I108802,I108598,I820912,I108842,I108607,I108864,I820915,I820924,I108881,I820918,I108907,I108924,I108610,I108946,I108595,I108977,I820921,I108994,I109011,I109028,I108604,I109059,I108592,I108601,I108589,I109145,I515068,I109171,I109179,I109196,I515059,I515077,I109213,I515056,I109239,I109256,I109264,I515062,I109281,I109113,I109312,I109329,I109125,I109369,I109134,I109391,I515074,I515065,I109408,I515080,I109434,I109451,I109137,I109473,I109122,I109504,I515071,I109521,I109538,I109555,I109131,I109586,I109119,I109128,I109116,I109672,I411580,I109698,I109706,I109723,I411601,I411595,I109740,I411577,I109766,I109783,I109791,I411589,I109808,I109640,I109839,I109856,I109652,I411586,I109896,I109661,I109918,I411592,I411583,I109935,I109961,I109978,I109664,I110000,I109649,I110031,I411598,I110048,I110065,I110082,I109658,I110113,I109646,I109655,I109643,I110199,I613906,I110225,I110233,I110250,I613897,I613915,I110267,I613894,I110293,I110310,I110318,I613900,I110335,I110167,I110366,I110383,I110179,I110423,I110188,I110445,I613912,I613903,I110462,I613918,I110488,I110505,I110191,I110527,I110176,I110558,I613909,I110575,I110592,I110609,I110185,I110640,I110173,I110182,I110170,I110726,I897562,I110752,I110760,I110777,I897577,I897556,I110794,I897559,I110820,I897580,I110837,I110845,I110862,I110694,I110893,I110910,I110706,I110950,I110715,I110972,I897568,I897565,I110989,I897571,I111015,I111032,I110718,I111054,I110703,I111085,I897574,I111102,I111119,I111136,I110712,I111167,I110700,I110709,I110697,I111253,I931086,I111279,I111287,I111304,I931101,I931080,I111321,I931083,I111347,I931104,I111364,I111372,I111389,I111221,I111420,I111437,I111233,I111477,I111242,I111499,I931092,I931089,I111516,I931095,I111542,I111559,I111245,I111581,I111230,I111612,I931098,I111629,I111646,I111663,I111239,I111694,I111227,I111236,I111224,I111780,I263313,I111806,I111814,I111831,I263295,I263310,I111848,I263286,I111874,I263289,I111891,I111899,I263304,I111916,I111748,I111947,I111964,I111760,I263307,I112004,I111769,I112026,I263298,I112043,I263292,I112069,I112086,I111772,I112108,I111757,I112139,I263301,I112156,I112173,I112190,I111766,I112221,I111754,I111763,I111751,I112310,I286483,I112336,I112344,I286480,I112370,I112378,I286477,I112395,I286489,I112412,I112287,I112443,I286498,I112281,I112474,I286495,I112491,I112508,I286474,I112525,I112542,I112559,I112296,I112293,I112299,I112618,I112635,I112652,I286486,I286501,I112678,I112278,I112709,I112717,I286492,I112302,I112748,I112765,I112782,I112284,I112813,I112830,I112275,I112290,I112905,I434151,I112931,I112939,I434136,I112965,I112973,I434160,I112990,I434139,I113007,I112882,I113038,I434142,I112876,I113069,I434145,I113086,I113103,I434148,I434154,I113120,I113137,I113154,I112891,I112888,I112894,I113213,I113230,I113247,I434157,I113273,I112873,I113304,I113312,I112897,I113343,I113360,I113377,I112879,I113408,I113425,I112870,I112885,I113500,I945533,I113526,I113534,I945530,I113560,I113568,I945539,I113585,I113602,I113477,I113633,I945542,I113471,I113664,I945536,I113681,I113698,I945551,I113715,I113732,I113749,I113486,I113483,I113489,I113808,I113825,I113842,I945554,I945548,I113868,I113468,I113899,I113907,I945545,I113492,I113938,I113955,I113972,I113474,I114003,I114020,I113465,I113480,I114095,I491373,I114121,I114129,I491358,I114155,I114163,I491382,I114180,I491361,I114197,I114228,I491364,I114259,I491367,I114276,I114293,I491370,I491376,I114310,I114327,I114344,I114403,I114420,I114437,I491379,I114463,I114494,I114502,I114533,I114550,I114567,I114598,I114615,I114690,I875595,I114716,I114724,I875592,I114750,I114758,I875601,I114775,I114792,I114823,I875604,I114854,I875598,I114871,I114888,I875613,I114905,I114922,I114939,I114998,I115015,I115032,I875616,I875610,I115058,I115089,I115097,I875607,I115128,I115145,I115162,I115193,I115210,I115285,I259079,I115311,I115319,I259076,I115345,I115353,I259073,I115370,I259085,I115387,I115262,I115418,I259094,I115256,I115449,I259091,I115466,I115483,I259070,I115500,I115517,I115534,I115271,I115268,I115274,I115593,I115610,I115627,I259082,I259097,I115653,I115253,I115684,I115692,I259088,I115277,I115723,I115740,I115757,I115259,I115788,I115805,I115250,I115265,I115880,I678126,I115906,I115914,I115940,I115948,I678123,I115965,I678135,I115982,I116013,I678129,I116044,I678141,I116061,I116078,I678132,I678120,I116095,I116112,I116129,I116188,I116205,I116222,I116248,I116279,I116287,I678138,I116318,I116335,I116352,I116383,I116400,I116475,I973889,I116501,I116509,I973901,I116535,I116543,I973907,I116560,I973886,I116577,I116452,I116608,I973904,I116446,I116639,I116656,I116673,I973892,I116690,I116707,I116724,I116461,I116458,I116464,I116783,I116800,I116817,I973910,I973898,I116843,I116443,I116874,I116882,I973895,I116467,I116913,I116930,I116947,I116449,I116978,I116995,I116440,I116455,I117070,I298077,I117096,I117104,I298074,I117130,I117138,I298071,I117155,I298083,I117172,I117203,I298092,I117234,I298089,I117251,I117268,I298068,I117285,I117302,I117319,I117378,I117395,I117412,I298080,I298095,I117438,I117469,I117477,I298086,I117508,I117525,I117542,I117573,I117590,I117665,I976065,I117691,I117699,I976077,I117725,I117733,I976083,I117750,I976062,I117767,I117642,I117798,I976080,I117636,I117829,I117846,I117863,I976068,I117880,I117897,I117914,I117651,I117648,I117654,I117973,I117990,I118007,I976086,I976074,I118033,I117633,I118064,I118072,I976071,I117657,I118103,I118120,I118137,I117639,I118168,I118185,I117630,I117645,I118260,I662843,I118286,I118294,I118320,I118328,I662840,I118345,I662852,I118362,I118237,I118393,I662846,I118231,I118424,I662858,I118441,I118458,I662849,I662837,I118475,I118492,I118509,I118246,I118243,I118249,I118568,I118585,I118602,I118628,I118228,I118659,I118667,I662855,I118252,I118698,I118715,I118732,I118234,I118763,I118780,I118225,I118240,I118855,I212176,I118881,I118889,I212173,I118915,I118923,I212170,I118940,I212182,I118957,I118832,I118988,I212191,I118826,I119019,I212188,I119036,I119053,I212167,I119070,I119087,I119104,I118841,I118838,I118844,I119163,I119180,I119197,I212179,I212194,I119223,I118823,I119254,I119262,I212185,I118847,I119293,I119310,I119327,I118829,I119358,I119375,I118820,I118835,I119450,I360618,I119476,I119484,I360612,I119510,I119518,I360609,I119535,I360600,I119552,I119427,I119583,I360603,I119421,I119614,I360606,I119631,I119648,I360594,I360621,I119665,I119682,I119699,I119436,I119433,I119439,I119758,I119775,I119792,I360597,I119818,I119418,I119849,I119857,I360615,I119442,I119888,I119905,I119922,I119424,I119953,I119970,I119415,I119430,I120045,I701909,I120071,I120079,I701930,I120105,I120113,I701912,I120130,I701903,I120147,I120022,I120178,I701915,I120016,I120209,I701906,I120226,I120243,I701924,I701927,I120260,I120277,I120294,I120031,I120028,I120034,I120353,I120370,I120387,I701918,I701921,I120413,I120013,I120444,I120452,I120037,I120483,I120500,I120517,I120019,I120548,I120565,I120010,I120025,I120640,I767801,I120666,I120674,I767822,I120700,I120708,I767804,I120725,I767795,I120742,I120617,I120773,I767807,I120611,I120804,I767798,I120821,I120838,I767816,I767819,I120855,I120872,I120889,I120626,I120623,I120629,I120948,I120965,I120982,I767810,I767813,I121008,I120608,I121039,I121047,I120632,I121078,I121095,I121112,I120614,I121143,I121160,I120605,I120620,I121235,I888311,I121261,I121269,I888308,I121295,I121303,I888317,I121320,I121337,I121212,I121368,I888320,I121206,I121399,I888314,I121416,I121433,I888329,I121450,I121467,I121484,I121221,I121218,I121224,I121543,I121560,I121577,I888332,I888326,I121603,I121203,I121634,I121642,I888323,I121227,I121673,I121690,I121707,I121209,I121738,I121755,I121200,I121215,I121827,I760058,I121853,I121870,I121819,I121892,I760067,I121918,I121926,I121943,I760055,I121960,I760046,I121977,I121994,I760052,I122011,I760070,I122028,I760043,I122045,I121795,I122076,I122093,I122110,I122127,I121807,I121801,I122172,I760049,I121816,I121810,I122217,I122234,I760061,I122251,I122268,I760064,I122294,I122302,I121804,I121798,I122356,I122364,I121813,I122422,I276461,I122448,I122465,I122414,I122487,I276476,I122513,I122521,I122538,I276473,I122555,I122572,I122589,I276470,I122606,I276485,I122623,I276482,I122640,I122390,I122671,I122688,I122705,I122722,I122402,I122396,I122767,I276479,I122411,I122405,I122812,I122829,I276467,I122846,I276488,I122863,I276464,I122889,I122897,I122399,I122393,I122951,I122959,I122408,I123017,I952466,I123043,I123060,I123009,I123082,I123108,I123116,I123133,I952469,I123150,I952481,I123167,I123184,I952487,I123201,I952478,I123218,I952484,I123235,I122985,I123266,I123283,I123300,I123317,I122997,I122991,I123362,I952475,I123006,I123000,I123407,I123424,I952472,I123441,I952490,I123458,I123484,I123492,I122994,I122988,I123546,I123554,I123003,I123612,I123638,I123655,I123604,I123677,I123703,I123711,I123728,I123745,I123762,I123779,I123796,I123813,I123830,I123580,I123861,I123878,I123895,I123912,I123592,I123586,I123957,I123601,I123595,I124002,I124019,I124036,I124053,I124079,I124087,I123589,I123583,I124141,I124149,I123598,I124207,I490217,I124233,I124250,I124199,I124272,I490208,I124298,I124306,I124323,I490226,I124340,I490223,I124357,I124374,I490202,I124391,I490205,I124408,I490214,I124425,I124175,I124456,I124473,I124490,I124507,I124187,I124181,I124552,I490220,I124196,I124190,I124597,I124614,I124631,I490211,I124648,I124674,I124682,I124184,I124178,I124736,I124744,I124193,I124802,I922410,I124828,I124845,I124794,I124867,I124893,I124901,I124918,I922413,I124935,I922425,I124952,I124969,I922431,I124986,I922422,I125003,I922428,I125020,I124770,I125051,I125068,I125085,I125102,I124782,I124776,I125147,I922419,I124791,I124785,I125192,I125209,I922416,I125226,I922434,I125243,I125269,I125277,I124779,I124773,I125331,I125339,I124788,I125397,I535876,I125423,I125440,I125389,I125462,I535873,I125488,I125496,I125513,I535879,I125530,I535864,I125547,I125564,I535867,I125581,I535888,I125598,I535885,I125615,I125365,I125646,I125663,I125680,I125697,I125377,I125371,I125742,I125386,I125380,I125787,I125804,I535870,I125821,I535882,I125838,I125864,I125872,I125374,I125368,I125926,I125934,I125383,I125992,I629115,I126018,I126035,I125984,I126057,I629109,I126083,I126091,I126108,I629127,I126125,I126142,I126159,I126176,I629121,I126193,I629112,I126210,I125960,I126241,I126258,I126275,I126292,I125972,I125966,I126337,I629124,I125981,I125975,I126382,I126399,I629130,I126416,I126433,I629118,I126459,I126467,I125969,I125963,I126521,I126529,I125978,I126587,I509288,I126613,I126630,I126579,I126652,I509285,I126678,I126686,I126703,I509291,I126720,I509276,I126737,I126754,I509279,I126771,I509300,I126788,I509297,I126805,I126555,I126836,I126853,I126870,I126887,I126567,I126561,I126932,I126576,I126570,I126977,I126994,I509282,I127011,I509294,I127028,I127054,I127062,I126564,I126558,I127116,I127124,I126573,I127182,I234301,I127208,I127225,I127174,I127247,I234316,I127273,I127281,I127298,I234313,I127315,I127332,I127349,I234310,I127366,I234325,I127383,I234322,I127400,I127150,I127431,I127448,I127465,I127482,I127162,I127156,I127527,I234319,I127171,I127165,I127572,I127589,I234307,I127606,I234328,I127623,I234304,I127649,I127657,I127159,I127153,I127711,I127719,I127168,I127777,I127803,I127820,I127769,I127842,I127868,I127876,I127893,I127910,I127927,I127944,I127961,I127978,I127995,I127745,I128026,I128043,I128060,I128077,I127757,I127751,I128122,I127766,I127760,I128167,I128184,I128201,I128218,I128244,I128252,I127754,I127748,I128306,I128314,I127763,I128372,I601190,I128398,I128415,I128364,I128437,I601187,I128463,I128471,I128488,I601193,I128505,I601178,I128522,I128539,I601181,I128556,I601202,I128573,I601199,I128590,I128340,I128621,I128638,I128655,I128672,I128352,I128346,I128717,I128361,I128355,I128762,I128779,I601184,I128796,I601196,I128813,I128839,I128847,I128349,I128343,I128901,I128909,I128358,I128967,I1005339,I128993,I129010,I128959,I129032,I1005351,I129058,I129066,I129083,I1005345,I129100,I1005357,I129117,I129134,I1005342,I129151,I1005354,I129168,I1005336,I129185,I128935,I129216,I129233,I129250,I129267,I128947,I128941,I129312,I1005348,I128956,I128950,I129357,I129374,I129391,I129408,I1005360,I129434,I129442,I128944,I128938,I129496,I129504,I128953,I129562,I388906,I129588,I129605,I129554,I129627,I388894,I129653,I129661,I129678,I388903,I129695,I388900,I129712,I129729,I388891,I129746,I388897,I129763,I388882,I129780,I129530,I129811,I129828,I129845,I129862,I129542,I129536,I129907,I129551,I129545,I129952,I129969,I388888,I129986,I388885,I130003,I388909,I130029,I130037,I129539,I129533,I130091,I130099,I129548,I130157,I926456,I130183,I130200,I130149,I130222,I130248,I130256,I130273,I926459,I130290,I926471,I130307,I130324,I926477,I130341,I926468,I130358,I926474,I130375,I130125,I130406,I130423,I130440,I130457,I130137,I130131,I130502,I926465,I130146,I130140,I130547,I130564,I926462,I130581,I926480,I130598,I130624,I130632,I130134,I130128,I130686,I130694,I130143,I130752,I691828,I130778,I130795,I130744,I130817,I691822,I130843,I130851,I130868,I691840,I130885,I130902,I130919,I130936,I691834,I130953,I691825,I130970,I130720,I131001,I131018,I131035,I131052,I130732,I130726,I131097,I691837,I130741,I130735,I131142,I131159,I691843,I131176,I131193,I691831,I131219,I131227,I130729,I130723,I131281,I131289,I130738,I131347,I131373,I131390,I131339,I131412,I131438,I131446,I131463,I131480,I131497,I131514,I131531,I131548,I131565,I131315,I131596,I131613,I131630,I131647,I131327,I131321,I131692,I131336,I131330,I131737,I131754,I131771,I131788,I131814,I131822,I131324,I131318,I131876,I131884,I131333,I131942,I827638,I131968,I131985,I131934,I132007,I827647,I132033,I132041,I132058,I827641,I132075,I827635,I132092,I132109,I827650,I132126,I132143,I827644,I132160,I131910,I132191,I132208,I132225,I132242,I131922,I131916,I132287,I131931,I131925,I132332,I132349,I827656,I132366,I827653,I132383,I132409,I132417,I131919,I131913,I132471,I132479,I131928,I132537,I508132,I132563,I132580,I132529,I132602,I508129,I132628,I132636,I132653,I508135,I132670,I508120,I132687,I132704,I508123,I132721,I508144,I132738,I508141,I132755,I132505,I132786,I132803,I132820,I132837,I132517,I132511,I132882,I132526,I132520,I132927,I132944,I508126,I132961,I508138,I132978,I133004,I133012,I132514,I132508,I133066,I133074,I132523,I133132,I536454,I133158,I133175,I133124,I133197,I536451,I133223,I133231,I133248,I536457,I133265,I536442,I133282,I133299,I536445,I133316,I536466,I133333,I536463,I133350,I133100,I133381,I133398,I133415,I133432,I133112,I133106,I133477,I133121,I133115,I133522,I133539,I536448,I133556,I536460,I133573,I133599,I133607,I133109,I133103,I133661,I133669,I133118,I133727,I533564,I133753,I133770,I133719,I133792,I533561,I133818,I133826,I133843,I533567,I133860,I533552,I133877,I133894,I533555,I133911,I533576,I133928,I533573,I133945,I133695,I133976,I133993,I134010,I134027,I133707,I133701,I134072,I133716,I133710,I134117,I134134,I533558,I134151,I533570,I134168,I134194,I134202,I133704,I133698,I134256,I134264,I133713,I134322,I604658,I134348,I134365,I134314,I134387,I604655,I134413,I134421,I134438,I604661,I134455,I604646,I134472,I134489,I604649,I134506,I604670,I134523,I604667,I134540,I134290,I134571,I134588,I134605,I134622,I134302,I134296,I134667,I134311,I134305,I134712,I134729,I604652,I134746,I604664,I134763,I134789,I134797,I134299,I134293,I134851,I134859,I134308,I134917,I366602,I134943,I134960,I134909,I134982,I366590,I135008,I135016,I135033,I366599,I135050,I366596,I135067,I135084,I366587,I135101,I366593,I135118,I366578,I135135,I134885,I135166,I135183,I135200,I135217,I134897,I134891,I135262,I134906,I134900,I135307,I135324,I366584,I135341,I366581,I135358,I366605,I135384,I135392,I134894,I134888,I135446,I135454,I134903,I135512,I637020,I135538,I135555,I135504,I135577,I637014,I135603,I135611,I135628,I637032,I135645,I135662,I135679,I135696,I637026,I135713,I637017,I135730,I135480,I135761,I135778,I135795,I135812,I135492,I135486,I135857,I637029,I135501,I135495,I135902,I135919,I637035,I135936,I135953,I637023,I135979,I135987,I135489,I135483,I136041,I136049,I135498,I136107,I787836,I136133,I136150,I136099,I136172,I787845,I136198,I136206,I136223,I787833,I136240,I787824,I136257,I136274,I787830,I136291,I787848,I136308,I787821,I136325,I136075,I136356,I136373,I136390,I136407,I136087,I136081,I136452,I787827,I136096,I136090,I136497,I136514,I787839,I136531,I136548,I787842,I136574,I136582,I136084,I136078,I136636,I136644,I136093,I136702,I635439,I136728,I136745,I136694,I136767,I635433,I136793,I136801,I136818,I635451,I136835,I136852,I136869,I136886,I635445,I136903,I635436,I136920,I136670,I136951,I136968,I136985,I137002,I136682,I136676,I137047,I635448,I136691,I136685,I137092,I137109,I635454,I137126,I137143,I635442,I137169,I137177,I136679,I136673,I137231,I137239,I136688,I137297,I858830,I137323,I137340,I137289,I137362,I137388,I137396,I137413,I858833,I137430,I858845,I137447,I137464,I858851,I137481,I858842,I137498,I858848,I137515,I137265,I137546,I137563,I137580,I137597,I137277,I137271,I137642,I858839,I137286,I137280,I137687,I137704,I858836,I137721,I858854,I137738,I137764,I137772,I137274,I137268,I137826,I137834,I137283,I137892,I137918,I137935,I137884,I137957,I137983,I137991,I138008,I138025,I138042,I138059,I138076,I138093,I138110,I137860,I138141,I138158,I138175,I138192,I137872,I137866,I138237,I137881,I137875,I138282,I138299,I138316,I138333,I138359,I138367,I137869,I137863,I138421,I138429,I137878,I138487,I885996,I138513,I138530,I138479,I138552,I138578,I138586,I138603,I885999,I138620,I886011,I138637,I138654,I886017,I138671,I886008,I138688,I886014,I138705,I138455,I138736,I138753,I138770,I138787,I138467,I138461,I138832,I886005,I138476,I138470,I138877,I138894,I886002,I138911,I886020,I138928,I138954,I138962,I138464,I138458,I139016,I139024,I138473,I139082,I438775,I139108,I139125,I139147,I438766,I139173,I139181,I139198,I438784,I139215,I438781,I139232,I139249,I438760,I139266,I438763,I139283,I438772,I139300,I139331,I139348,I139365,I139382,I139427,I438778,I139472,I139489,I139506,I438769,I139523,I139549,I139557,I139611,I139619,I139677,I293325,I139703,I139720,I139669,I139742,I293340,I139768,I139776,I139793,I293337,I139810,I139827,I139844,I293334,I139861,I293349,I139878,I293346,I139895,I139645,I139926,I139943,I139960,I139977,I139657,I139651,I140022,I293343,I139666,I139660,I140067,I140084,I293331,I140101,I293352,I140118,I293328,I140144,I140152,I139654,I139648,I140206,I140214,I139663,I140272,I867500,I140298,I140315,I140264,I140337,I140363,I140371,I140388,I867503,I140405,I867515,I140422,I140439,I867521,I140456,I867512,I140473,I867518,I140490,I140240,I140521,I140538,I140555,I140572,I140252,I140246,I140617,I867509,I140261,I140255,I140662,I140679,I867506,I140696,I867524,I140713,I140739,I140747,I140249,I140243,I140801,I140809,I140258,I140867,I736802,I140893,I140910,I140859,I140932,I736811,I140958,I140966,I140983,I736799,I141000,I736790,I141017,I141034,I736796,I141051,I736814,I141068,I736787,I141085,I140835,I141116,I141133,I141150,I141167,I140847,I140841,I141212,I736793,I140856,I140850,I141257,I141274,I736805,I141291,I141308,I736808,I141334,I141342,I140844,I140838,I141396,I141404,I140853,I141462,I141488,I141505,I141454,I141527,I141553,I141561,I141578,I141595,I141612,I141629,I141646,I141663,I141680,I141430,I141711,I141728,I141745,I141762,I141442,I141436,I141807,I141451,I141445,I141852,I141869,I141886,I141903,I141929,I141937,I141439,I141433,I141991,I141999,I141448,I142057,I626480,I142083,I142100,I142049,I142122,I626474,I142148,I142156,I142173,I626492,I142190,I142207,I142224,I142241,I626486,I142258,I626477,I142275,I142025,I142306,I142323,I142340,I142357,I142037,I142031,I142402,I626489,I142046,I142040,I142447,I142464,I626495,I142481,I142498,I626483,I142524,I142532,I142034,I142028,I142586,I142594,I142043,I142652,I763934,I142678,I142695,I142644,I142717,I763943,I142743,I142751,I142768,I763931,I142785,I763922,I142802,I142819,I763928,I142836,I763946,I142853,I763919,I142870,I142620,I142901,I142918,I142935,I142952,I142632,I142626,I142997,I763925,I142641,I142635,I143042,I143059,I763937,I143076,I143093,I763940,I143119,I143127,I142629,I142623,I143181,I143189,I142638,I143247,I890042,I143273,I143290,I143239,I143312,I143338,I143346,I143363,I890045,I143380,I890057,I143397,I143414,I890063,I143431,I890054,I143448,I890060,I143465,I143215,I143496,I143513,I143530,I143547,I143227,I143221,I143592,I890051,I143236,I143230,I143637,I143654,I890048,I143671,I890066,I143688,I143714,I143722,I143224,I143218,I143776,I143784,I143233,I143842,I292798,I143868,I143885,I143834,I143907,I292813,I143933,I143941,I143958,I292810,I143975,I143992,I144009,I292807,I144026,I292822,I144043,I292819,I144060,I143810,I144091,I144108,I144125,I144142,I143822,I143816,I144187,I292816,I143831,I143825,I144232,I144249,I292804,I144266,I292825,I144283,I292801,I144309,I144317,I143819,I143813,I144371,I144379,I143828,I144437,I144463,I144480,I144502,I144528,I144536,I144553,I144570,I144587,I144604,I144621,I144638,I144655,I144686,I144703,I144720,I144737,I144782,I144827,I144844,I144861,I144878,I144904,I144912,I144966,I144974,I145032,I496572,I145058,I145075,I145024,I145097,I496569,I145123,I145131,I145148,I496575,I145165,I496560,I145182,I145199,I496563,I145216,I496584,I145233,I496581,I145250,I145000,I145281,I145298,I145315,I145332,I145012,I145006,I145377,I145021,I145015,I145422,I145439,I496566,I145456,I496578,I145473,I145499,I145507,I145009,I145003,I145561,I145569,I145018,I145627,I778792,I145653,I145670,I145619,I145692,I778801,I145718,I145726,I145743,I778789,I145760,I778780,I145777,I145794,I778786,I145811,I778804,I145828,I778777,I145845,I145595,I145876,I145893,I145910,I145927,I145607,I145601,I145972,I778783,I145616,I145610,I146017,I146034,I778795,I146051,I146068,I778798,I146094,I146102,I145604,I145598,I146156,I146164,I145613,I146222,I834554,I146248,I146265,I146214,I146287,I146313,I146321,I146338,I834557,I146355,I834569,I146372,I146389,I834575,I146406,I834566,I146423,I834572,I146440,I146190,I146471,I146488,I146505,I146522,I146202,I146196,I146567,I834563,I146211,I146205,I146612,I146629,I834560,I146646,I834578,I146663,I146689,I146697,I146199,I146193,I146751,I146759,I146208,I146817,I461317,I146843,I146860,I146809,I146882,I461308,I146908,I146916,I146933,I461326,I146950,I461323,I146967,I146984,I461302,I147001,I461305,I147018,I461314,I147035,I146785,I147066,I147083,I147100,I147117,I146797,I146791,I147162,I461320,I146806,I146800,I147207,I147224,I147241,I461311,I147258,I147284,I147292,I146794,I146788,I147346,I147354,I146803,I147412,I319818,I147438,I147455,I147404,I147477,I319806,I147503,I147511,I147528,I319815,I147545,I319812,I147562,I147579,I319803,I147596,I319809,I147613,I319794,I147630,I147380,I147661,I147678,I147695,I147712,I147392,I147386,I147757,I147401,I147395,I147802,I147819,I319800,I147836,I319797,I147853,I319821,I147879,I147887,I147389,I147383,I147941,I147949,I147398,I148007,I1042400,I148033,I148050,I148072,I1042391,I148098,I148106,I148123,I1042385,I148140,I1042379,I148157,I148174,I1042406,I148191,I148208,I1042403,I148225,I148256,I148273,I148290,I148307,I148352,I1042388,I148397,I148414,I1042394,I148431,I1042397,I148448,I1042382,I148474,I148482,I148536,I148544,I148602,I513334,I148628,I148645,I148594,I148667,I513331,I148693,I148701,I148718,I513337,I148735,I513322,I148752,I148769,I513325,I148786,I513346,I148803,I513343,I148820,I148570,I148851,I148868,I148885,I148902,I148582,I148576,I148947,I148591,I148585,I148992,I149009,I513328,I149026,I513340,I149043,I149069,I149077,I148579,I148573,I149131,I149139,I148588,I149197,I149223,I149240,I149262,I149288,I149296,I149313,I149330,I149347,I149364,I149381,I149398,I149415,I149446,I149463,I149480,I149497,I149542,I149587,I149604,I149621,I149638,I149664,I149672,I149726,I149734,I149792,I1094760,I149818,I149835,I149857,I1094751,I149883,I149891,I149908,I1094745,I149925,I1094739,I149942,I149959,I1094766,I149976,I149993,I1094763,I150010,I150041,I150058,I150075,I150092,I150137,I1094748,I150182,I150199,I1094754,I150216,I1094757,I150233,I1094742,I150259,I150267,I150321,I150329,I150387,I471143,I150413,I150430,I150379,I150452,I471134,I150478,I150486,I150503,I471152,I150520,I471149,I150537,I150554,I471128,I150571,I471131,I150588,I471140,I150605,I150355,I150636,I150653,I150670,I150687,I150367,I150361,I150732,I471146,I150376,I150370,I150777,I150794,I150811,I471137,I150828,I150854,I150862,I150364,I150358,I150916,I150924,I150373,I150982,I772332,I151008,I151025,I150974,I151047,I772341,I151073,I151081,I151098,I772329,I151115,I772320,I151132,I151149,I772326,I151166,I772344,I151183,I772317,I151200,I150950,I151231,I151248,I151265,I151282,I150962,I150956,I151327,I772323,I150971,I150965,I151372,I151389,I772335,I151406,I151423,I772338,I151449,I151457,I150959,I150953,I151511,I151519,I150968,I151577,I354634,I151603,I151620,I151569,I151642,I354622,I151668,I151676,I151693,I354631,I151710,I354628,I151727,I151744,I354619,I151761,I354625,I151778,I354610,I151795,I151545,I151826,I151843,I151860,I151877,I151557,I151551,I151922,I151566,I151560,I151967,I151984,I354616,I152001,I354613,I152018,I354637,I152044,I152052,I151554,I151548,I152106,I152114,I151563,I152172,I254854,I152198,I152215,I152164,I152237,I254869,I152263,I152271,I152288,I254866,I152305,I152322,I152339,I254863,I152356,I254878,I152373,I254875,I152390,I152140,I152421,I152438,I152455,I152472,I152152,I152146,I152517,I254872,I152161,I152155,I152562,I152579,I254860,I152596,I254881,I152613,I254857,I152639,I152647,I152149,I152143,I152701,I152709,I152158,I152767,I226396,I152793,I152810,I152759,I152832,I226411,I152858,I152866,I152883,I226408,I152900,I152917,I152934,I226405,I152951,I226420,I152968,I226417,I152985,I152735,I153016,I153033,I153050,I153067,I152747,I152741,I153112,I226414,I152756,I152750,I153157,I153174,I226402,I153191,I226423,I153208,I226399,I153234,I153242,I152744,I152738,I153296,I153304,I152753,I153362,I418134,I153388,I153405,I153354,I153427,I418128,I153453,I153461,I153478,I418143,I153495,I418140,I153512,I153529,I418131,I153546,I418122,I153563,I418125,I153580,I153330,I153611,I153628,I153645,I153662,I153342,I153336,I153707,I418146,I153351,I153345,I153752,I153769,I418137,I153786,I153803,I153829,I153837,I153339,I153333,I153891,I153899,I153348,I153957,I857674,I153983,I154000,I153949,I154022,I154048,I154056,I154073,I857677,I154090,I857689,I154107,I154124,I857695,I154141,I857686,I154158,I857692,I154175,I153925,I154206,I154223,I154240,I154257,I153937,I153931,I154302,I857683,I153946,I153940,I154347,I154364,I857680,I154381,I857698,I154398,I154424,I154432,I153934,I153928,I154486,I154494,I153943,I154552,I678653,I154578,I154595,I154544,I154617,I678647,I154643,I154651,I154668,I678665,I154685,I154702,I154719,I154736,I678659,I154753,I678650,I154770,I154520,I154801,I154818,I154835,I154852,I154532,I154526,I154897,I678662,I154541,I154535,I154942,I154959,I678668,I154976,I154993,I678656,I155019,I155027,I154529,I154523,I155081,I155089,I154538,I155147,I1006495,I155173,I155190,I155139,I155212,I1006507,I155238,I155246,I155263,I1006501,I155280,I1006513,I155297,I155314,I1006498,I155331,I1006510,I155348,I1006492,I155365,I155115,I155396,I155413,I155430,I155447,I155127,I155121,I155492,I1006504,I155136,I155130,I155537,I155554,I155571,I155588,I1006516,I155614,I155622,I155124,I155118,I155676,I155684,I155133,I155742,I1056085,I155768,I155785,I155734,I155807,I1056076,I155833,I155841,I155858,I1056070,I155875,I1056064,I155892,I155909,I1056091,I155926,I155943,I1056088,I155960,I155710,I155991,I156008,I156025,I156042,I155722,I155716,I156087,I1056073,I155731,I155725,I156132,I156149,I1056079,I156166,I1056082,I156183,I1056067,I156209,I156217,I155719,I155713,I156271,I156279,I155728,I156337,I320906,I156363,I156380,I156329,I156402,I320894,I156428,I156436,I156453,I320903,I156470,I320900,I156487,I156504,I320891,I156521,I320897,I156538,I320882,I156555,I156305,I156586,I156603,I156620,I156637,I156317,I156311,I156682,I156326,I156320,I156727,I156744,I320888,I156761,I320885,I156778,I320909,I156804,I156812,I156314,I156308,I156866,I156874,I156323,I156932,I967376,I156958,I156975,I156924,I156997,I967361,I157023,I157031,I157048,I967379,I157065,I157082,I157099,I967382,I157116,I967373,I157133,I967370,I157150,I156900,I157181,I157198,I157215,I157232,I156912,I156906,I157277,I967367,I156921,I156915,I157322,I157339,I967358,I157356,I967364,I157373,I157399,I157407,I156909,I156903,I157461,I157469,I156918,I157527,I412184,I157553,I157570,I157519,I157592,I412178,I157618,I157626,I157643,I412193,I157660,I412190,I157677,I157694,I412181,I157711,I412172,I157728,I412175,I157745,I157495,I157776,I157793,I157810,I157827,I157507,I157501,I157872,I412196,I157516,I157510,I157917,I157934,I412187,I157951,I157968,I157994,I158002,I157504,I157498,I158056,I158064,I157513,I158122,I708378,I158148,I158165,I158114,I158187,I708387,I158213,I158221,I158238,I708375,I158255,I708366,I158272,I158289,I708372,I158306,I708390,I158323,I708363,I158340,I158090,I158371,I158388,I158405,I158422,I158102,I158096,I158467,I708369,I158111,I158105,I158512,I158529,I708381,I158546,I158563,I708384,I158589,I158597,I158099,I158093,I158651,I158659,I158108,I158717,I375306,I158743,I158760,I158709,I158782,I375294,I158808,I158816,I158833,I375303,I158850,I375300,I158867,I158884,I375291,I158901,I375297,I158918,I375282,I158935,I158685,I158966,I158983,I159000,I159017,I158697,I158691,I159062,I158706,I158700,I159107,I159124,I375288,I159141,I375285,I159158,I375309,I159184,I159192,I158694,I158688,I159246,I159254,I158703,I159312,I994357,I159338,I159355,I159377,I994369,I159403,I159411,I159428,I994363,I159445,I994375,I159462,I159479,I994360,I159496,I994372,I159513,I994354,I159530,I159561,I159578,I159595,I159612,I159657,I994366,I159702,I159719,I159736,I159753,I994378,I159779,I159787,I159841,I159849,I159907,I1087620,I159933,I159950,I159899,I159972,I1087611,I159998,I160006,I160023,I1087605,I160040,I1087599,I160057,I160074,I1087626,I160091,I160108,I1087623,I160125,I159875,I160156,I160173,I160190,I160207,I159887,I159881,I160252,I1087608,I159896,I159890,I160297,I160314,I1087614,I160331,I1087617,I160348,I1087602,I160374,I160382,I159884,I159878,I160436,I160444,I159893,I160502,I160528,I160545,I160494,I160567,I160593,I160601,I160618,I160635,I160652,I160669,I160686,I160703,I160720,I160470,I160751,I160768,I160785,I160802,I160482,I160476,I160847,I160491,I160485,I160892,I160909,I160926,I160943,I160969,I160977,I160479,I160473,I161031,I161039,I160488,I161097,I465363,I161123,I161140,I161089,I161162,I465354,I161188,I161196,I161213,I465372,I161230,I465369,I161247,I161264,I465348,I161281,I465351,I161298,I465360,I161315,I161065,I161346,I161363,I161380,I161397,I161077,I161071,I161442,I465366,I161086,I161080,I161487,I161504,I161521,I465357,I161538,I161564,I161572,I161074,I161068,I161626,I161634,I161083,I161692,I698152,I161718,I161735,I161684,I161757,I698146,I161783,I161791,I161808,I698164,I161825,I161842,I161859,I161876,I698158,I161893,I698149,I161910,I161660,I161941,I161958,I161975,I161992,I161672,I161666,I162037,I698161,I161681,I161675,I162082,I162099,I698167,I162116,I162133,I698155,I162159,I162167,I161669,I161663,I162221,I162229,I161678,I162287,I931658,I162313,I162330,I162279,I162352,I162378,I162386,I162403,I931661,I162420,I931673,I162437,I162454,I931679,I162471,I931670,I162488,I931676,I162505,I162255,I162536,I162553,I162570,I162587,I162267,I162261,I162632,I931667,I162276,I162270,I162677,I162694,I931664,I162711,I931682,I162728,I162754,I162762,I162264,I162258,I162816,I162824,I162273,I162882,I925300,I162908,I162925,I162874,I162947,I162973,I162981,I162998,I925303,I163015,I925315,I163032,I163049,I925321,I163066,I925312,I163083,I925318,I163100,I162850,I163131,I163148,I163165,I163182,I162862,I162856,I163227,I925309,I162871,I162865,I163272,I163289,I925306,I163306,I925324,I163323,I163349,I163357,I162859,I162853,I163411,I163419,I162868,I163477,I294906,I163503,I163520,I163469,I163542,I294921,I163568,I163576,I163593,I294918,I163610,I163627,I163644,I294915,I163661,I294930,I163678,I294927,I163695,I163445,I163726,I163743,I163760,I163777,I163457,I163451,I163822,I294924,I163466,I163460,I163867,I163884,I294912,I163901,I294933,I163918,I294909,I163944,I163952,I163454,I163448,I164006,I164014,I163463,I164072,I975536,I164098,I164115,I164064,I164137,I975521,I164163,I164171,I164188,I975539,I164205,I164222,I164239,I975542,I164256,I975533,I164273,I975530,I164290,I164040,I164321,I164338,I164355,I164372,I164052,I164046,I164417,I975527,I164061,I164055,I164462,I164479,I975518,I164496,I975524,I164513,I164539,I164547,I164049,I164043,I164601,I164609,I164058,I164667,I526628,I164693,I164710,I164659,I164732,I526625,I164758,I164766,I164783,I526631,I164800,I526616,I164817,I164834,I526619,I164851,I526640,I164868,I526637,I164885,I164635,I164916,I164933,I164950,I164967,I164647,I164641,I165012,I164656,I164650,I165057,I165074,I526622,I165091,I526634,I165108,I165134,I165142,I164644,I164638,I165196,I165204,I164653,I165262,I165288,I165305,I165254,I165327,I165353,I165361,I165378,I165395,I165412,I165429,I165446,I165463,I165480,I165230,I165511,I165528,I165545,I165562,I165242,I165236,I165607,I165251,I165245,I165652,I165669,I165686,I165703,I165729,I165737,I165239,I165233,I165791,I165799,I165248,I165857,I881950,I165883,I165900,I165849,I165922,I165948,I165956,I165973,I881953,I165990,I881965,I166007,I166024,I881971,I166041,I881962,I166058,I881968,I166075,I165825,I166106,I166123,I166140,I166157,I165837,I165831,I166202,I881959,I165846,I165840,I166247,I166264,I881956,I166281,I881974,I166298,I166324,I166332,I165834,I165828,I166386,I166394,I165843,I166452,I280677,I166478,I166495,I166444,I166517,I280692,I166543,I166551,I166568,I280689,I166585,I166602,I166619,I280686,I166636,I280701,I166653,I280698,I166670,I166420,I166701,I166718,I166735,I166752,I166432,I166426,I166797,I280695,I166441,I166435,I166842,I166859,I280683,I166876,I280704,I166893,I280680,I166919,I166927,I166429,I166423,I166981,I166989,I166438,I167047,I611016,I167073,I167090,I167112,I611013,I167138,I167146,I167163,I611019,I167180,I611004,I167197,I167214,I611007,I167231,I611028,I167248,I611025,I167265,I167296,I167313,I167330,I167347,I167392,I167437,I167454,I611010,I167471,I611022,I167488,I167514,I167522,I167576,I167584,I167642,I269083,I167668,I167685,I167634,I167707,I269098,I167733,I167741,I167758,I269095,I167775,I167792,I167809,I269092,I167826,I269107,I167843,I269104,I167860,I167610,I167891,I167908,I167925,I167942,I167622,I167616,I167987,I269101,I167631,I167625,I168032,I168049,I269089,I168066,I269110,I168083,I269086,I168109,I168117,I167619,I167613,I168171,I168179,I167628,I168237,I957040,I168263,I168280,I168229,I168302,I957025,I168328,I168336,I168353,I957043,I168370,I168387,I168404,I957046,I168421,I957037,I168438,I957034,I168455,I168205,I168486,I168503,I168520,I168537,I168217,I168211,I168582,I957031,I168226,I168220,I168627,I168644,I957022,I168661,I957028,I168678,I168704,I168712,I168214,I168208,I168766,I168774,I168223,I168832,I347018,I168858,I168875,I168824,I168897,I347006,I168923,I168931,I168948,I347015,I168965,I347012,I168982,I168999,I347003,I169016,I347009,I169033,I346994,I169050,I168800,I169081,I169098,I169115,I169132,I168812,I168806,I169177,I168821,I168815,I169222,I169239,I347000,I169256,I346997,I169273,I347021,I169299,I169307,I168809,I168803,I169361,I169369,I168818,I169427,I632277,I169453,I169470,I169419,I169492,I632271,I169518,I169526,I169543,I632289,I169560,I169577,I169594,I169611,I632283,I169628,I632274,I169645,I169395,I169676,I169693,I169710,I169727,I169407,I169401,I169772,I632286,I169416,I169410,I169817,I169834,I632292,I169851,I169868,I632280,I169894,I169902,I169404,I169398,I169956,I169964,I169413,I170022,I615062,I170048,I170065,I170014,I170087,I615059,I170113,I170121,I170138,I615065,I170155,I615050,I170172,I170189,I615053,I170206,I615074,I170223,I615071,I170240,I169990,I170271,I170288,I170305,I170322,I170002,I169996,I170367,I170011,I170005,I170412,I170429,I615056,I170446,I615068,I170463,I170489,I170497,I169999,I169993,I170551,I170559,I170008,I170617,I170643,I170660,I170609,I170682,I170708,I170716,I170733,I170750,I170767,I170784,I170801,I170818,I170835,I170585,I170866,I170883,I170900,I170917,I170597,I170591,I170962,I170606,I170600,I171007,I171024,I171041,I171058,I171084,I171092,I170594,I170588,I171146,I171154,I170603,I171212,I171238,I171255,I171204,I171277,I171303,I171311,I171328,I171345,I171362,I171379,I171396,I171413,I171430,I171180,I171461,I171478,I171495,I171512,I171192,I171186,I171557,I171201,I171195,I171602,I171619,I171636,I171653,I171679,I171687,I171189,I171183,I171741,I171749,I171198,I171807,I485015,I171833,I171850,I171799,I171872,I485006,I171898,I171906,I171923,I485024,I171940,I485021,I171957,I171974,I485000,I171991,I485003,I172008,I485012,I172025,I171775,I172056,I172073,I172090,I172107,I171787,I171781,I172152,I485018,I171796,I171790,I172197,I172214,I172231,I485009,I172248,I172274,I172282,I171784,I171778,I172336,I172344,I171793,I172402,I652303,I172428,I172445,I172394,I172467,I652297,I172493,I172501,I172518,I652315,I172535,I172552,I172569,I172586,I652309,I172603,I652300,I172620,I172370,I172651,I172668,I172685,I172702,I172382,I172376,I172747,I652312,I172391,I172385,I172792,I172809,I652318,I172826,I172843,I652306,I172869,I172877,I172379,I172373,I172931,I172939,I172388,I172997,I173023,I173040,I173062,I173088,I173096,I173113,I173130,I173147,I173164,I173181,I173198,I173215,I173246,I173263,I173280,I173297,I173342,I173387,I173404,I173421,I173438,I173464,I173472,I173526,I173534,I173592,I173618,I173635,I173584,I173657,I173683,I173691,I173708,I173725,I173742,I173759,I173776,I173793,I173810,I173560,I173841,I173858,I173875,I173892,I173572,I173566,I173937,I173581,I173575,I173982,I173999,I174016,I174033,I174059,I174067,I173569,I173563,I174121,I174129,I173578,I174187,I802393,I174213,I174230,I174179,I174252,I802402,I174278,I174286,I174303,I802396,I174320,I802390,I174337,I174354,I802405,I174371,I174388,I802399,I174405,I174155,I174436,I174453,I174470,I174487,I174167,I174161,I174532,I174176,I174170,I174577,I174594,I802411,I174611,I802408,I174628,I174654,I174662,I174164,I174158,I174716,I174724,I174173,I174782,I663370,I174808,I174825,I174774,I174847,I663364,I174873,I174881,I174898,I663382,I174915,I174932,I174949,I174966,I663376,I174983,I663367,I175000,I174750,I175031,I175048,I175065,I175082,I174762,I174756,I175127,I663379,I174771,I174765,I175172,I175189,I663385,I175206,I175223,I663373,I175249,I175257,I174759,I174753,I175311,I175319,I174768,I175377,I175403,I175420,I175369,I175442,I175468,I175476,I175493,I175510,I175527,I175544,I175561,I175578,I175595,I175345,I175626,I175643,I175660,I175677,I175357,I175351,I175722,I175366,I175360,I175767,I175784,I175801,I175818,I175844,I175852,I175354,I175348,I175906,I175914,I175363,I175972,I859986,I175998,I176015,I175964,I176037,I176063,I176071,I176088,I859989,I176105,I860001,I176122,I176139,I860007,I176156,I859998,I176173,I860004,I176190,I175940,I176221,I176238,I176255,I176272,I175952,I175946,I176317,I859995,I175961,I175955,I176362,I176379,I859992,I176396,I860010,I176413,I176439,I176447,I175949,I175943,I176501,I176509,I175958,I176567,I909694,I176593,I176610,I176632,I176658,I176666,I176683,I909697,I176700,I909709,I176717,I176734,I909715,I176751,I909706,I176768,I909712,I176785,I176816,I176833,I176850,I176867,I176912,I909703,I176957,I176974,I909700,I176991,I909718,I177008,I177034,I177042,I177096,I177104,I177162,I751660,I177188,I177205,I177154,I177227,I751669,I177253,I177261,I177278,I751657,I177295,I751648,I177312,I177329,I751654,I177346,I751672,I177363,I751645,I177380,I177130,I177411,I177428,I177445,I177462,I177142,I177136,I177507,I751651,I177151,I177145,I177552,I177569,I751663,I177586,I177603,I751666,I177629,I177637,I177139,I177133,I177691,I177699,I177148,I177757,I628588,I177783,I177800,I177749,I177822,I628582,I177848,I177856,I177873,I628600,I177890,I177907,I177924,I177941,I628594,I177958,I628585,I177975,I177725,I178006,I178023,I178040,I178057,I177737,I177731,I178102,I628597,I177746,I177740,I178147,I178164,I628603,I178181,I178198,I628591,I178224,I178232,I177734,I177728,I178286,I178294,I177743,I178352,I732280,I178378,I178395,I178344,I178417,I732289,I178443,I178451,I178468,I732277,I178485,I732268,I178502,I178519,I732274,I178536,I732292,I178553,I732265,I178570,I178320,I178601,I178618,I178635,I178652,I178332,I178326,I178697,I732271,I178341,I178335,I178742,I178759,I732283,I178776,I178793,I732286,I178819,I178827,I178329,I178323,I178881,I178889,I178338,I178947,I531830,I178973,I178990,I179012,I531827,I179038,I179046,I179063,I531833,I179080,I531818,I179097,I179114,I531821,I179131,I531842,I179148,I531839,I179165,I179196,I179213,I179230,I179247,I179292,I179337,I179354,I531824,I179371,I531836,I179388,I179414,I179422,I179476,I179484,I179542,I938016,I179568,I179585,I179534,I179607,I179633,I179641,I179658,I938019,I179675,I938031,I179692,I179709,I938037,I179726,I938028,I179743,I938034,I179760,I179510,I179791,I179808,I179825,I179842,I179522,I179516,I179887,I938025,I179531,I179525,I179932,I179949,I938022,I179966,I938040,I179983,I180009,I180017,I179519,I179513,I180071,I180079,I179528,I180137,I650195,I180163,I180180,I180129,I180202,I650189,I180228,I180236,I180253,I650207,I180270,I180287,I180304,I180321,I650201,I180338,I650192,I180355,I180105,I180386,I180403,I180420,I180437,I180117,I180111,I180482,I650204,I180126,I180120,I180527,I180544,I650210,I180561,I180578,I650198,I180604,I180612,I180114,I180108,I180666,I180674,I180123,I180732,I313351,I180758,I180775,I180724,I180797,I313366,I180823,I180831,I180848,I313363,I180865,I180882,I180899,I313360,I180916,I313375,I180933,I313372,I180950,I180700,I180981,I180998,I181015,I181032,I180712,I180706,I181077,I313369,I180721,I180715,I181122,I181139,I313357,I181156,I313378,I181173,I313354,I181199,I181207,I180709,I180703,I181261,I181269,I180718,I181327,I901024,I181353,I181370,I181319,I181392,I181418,I181426,I181443,I901027,I181460,I901039,I181477,I181494,I901045,I181511,I901036,I181528,I901042,I181545,I181295,I181576,I181593,I181610,I181627,I181307,I181301,I181672,I901033,I181316,I181310,I181717,I181734,I901030,I181751,I901048,I181768,I181794,I181802,I181304,I181298,I181856,I181864,I181313,I181922,I785898,I181948,I181965,I181914,I181987,I785907,I182013,I182021,I182038,I785895,I182055,I785886,I182072,I182089,I785892,I182106,I785910,I182123,I785883,I182140,I181890,I182171,I182188,I182205,I182222,I181902,I181896,I182267,I785889,I181911,I181905,I182312,I182329,I785901,I182346,I182363,I785904,I182389,I182397,I181899,I181893,I182451,I182459,I181908,I182517,I430034,I182543,I182560,I182509,I182582,I430028,I182608,I182616,I182633,I430043,I182650,I430040,I182667,I182684,I430031,I182701,I430022,I182718,I430025,I182735,I182485,I182766,I182783,I182800,I182817,I182497,I182491,I182862,I430046,I182506,I182500,I182907,I182924,I430037,I182941,I182958,I182984,I182992,I182494,I182488,I183046,I183054,I182503,I183112,I183138,I183155,I183104,I183177,I183203,I183211,I183228,I183245,I183262,I183279,I183296,I183313,I183330,I183080,I183361,I183378,I183395,I183412,I183092,I183086,I183457,I183101,I183095,I183502,I183519,I183536,I183553,I183579,I183587,I183089,I183083,I183641,I183649,I183098,I183707,I898712,I183733,I183750,I183699,I183772,I183798,I183806,I183823,I898715,I183840,I898727,I183857,I183874,I898733,I183891,I898724,I183908,I898730,I183925,I183675,I183956,I183973,I183990,I184007,I183687,I183681,I184052,I898721,I183696,I183690,I184097,I184114,I898718,I184131,I898736,I184148,I184174,I184182,I183684,I183678,I184236,I184244,I183693,I184302,I944952,I184328,I184345,I184294,I184367,I184393,I184401,I184418,I944955,I184435,I944967,I184452,I184469,I944973,I184486,I944964,I184503,I944970,I184520,I184270,I184551,I184568,I184585,I184602,I184282,I184276,I184647,I944961,I184291,I184285,I184692,I184709,I944958,I184726,I944976,I184743,I184769,I184777,I184279,I184273,I184831,I184839,I184288,I184897,I548592,I184923,I184940,I184889,I184962,I548589,I184988,I184996,I185013,I548595,I185030,I548580,I185047,I185064,I548583,I185081,I548604,I185098,I548601,I185115,I184865,I185146,I185163,I185180,I185197,I184877,I184871,I185242,I184886,I184880,I185287,I185304,I548586,I185321,I548598,I185338,I185364,I185372,I184874,I184868,I185426,I185434,I184883,I185492,I586740,I185518,I185535,I185484,I185557,I586737,I185583,I185591,I185608,I586743,I185625,I586728,I185642,I185659,I586731,I185676,I586752,I185693,I586749,I185710,I185460,I185741,I185758,I185775,I185792,I185472,I185466,I185837,I185481,I185475,I185882,I185899,I586734,I185916,I586746,I185933,I185959,I185967,I185469,I185463,I186021,I186029,I185478,I186087,I462473,I186113,I186130,I186079,I186152,I462464,I186178,I186186,I186203,I462482,I186220,I462479,I186237,I186254,I462458,I186271,I462461,I186288,I462470,I186305,I186055,I186336,I186353,I186370,I186387,I186067,I186061,I186432,I462476,I186076,I186070,I186477,I186494,I186511,I462467,I186528,I186554,I186562,I186064,I186058,I186616,I186624,I186073,I186682,I1088810,I186708,I186725,I186674,I186747,I1088801,I186773,I186781,I186798,I1088795,I186815,I1088789,I186832,I186849,I1088816,I186866,I186883,I1088813,I186900,I186650,I186931,I186948,I186965,I186982,I186662,I186656,I187027,I1088798,I186671,I186665,I187072,I187089,I1088804,I187106,I1088807,I187123,I1088792,I187149,I187157,I186659,I186653,I187211,I187219,I186668,I187277,I964112,I187303,I187320,I187269,I187342,I964097,I187368,I187376,I187393,I964115,I187410,I187427,I187444,I964118,I187461,I964109,I187478,I964106,I187495,I187245,I187526,I187543,I187560,I187577,I187257,I187251,I187622,I964103,I187266,I187260,I187667,I187684,I964094,I187701,I964100,I187718,I187744,I187752,I187254,I187248,I187806,I187814,I187263,I187872,I737448,I187898,I187915,I187864,I187937,I737457,I187963,I187971,I187988,I737445,I188005,I737436,I188022,I188039,I737442,I188056,I737460,I188073,I737433,I188090,I187840,I188121,I188138,I188155,I188172,I187852,I187846,I188217,I737439,I187861,I187855,I188262,I188279,I737451,I188296,I188313,I737454,I188339,I188347,I187849,I187843,I188401,I188409,I187858,I188467,I771040,I188493,I188510,I188459,I188532,I771049,I188558,I188566,I188583,I771037,I188600,I771028,I188617,I188634,I771034,I188651,I771052,I188668,I771025,I188685,I188435,I188716,I188733,I188750,I188767,I188447,I188441,I188812,I771031,I188456,I188450,I188857,I188874,I771043,I188891,I188908,I771046,I188934,I188942,I188444,I188438,I188996,I189004,I188453,I189062,I529518,I189088,I189105,I189054,I189127,I529515,I189153,I189161,I189178,I529521,I189195,I529506,I189212,I189229,I529509,I189246,I529530,I189263,I529527,I189280,I189030,I189311,I189328,I189345,I189362,I189042,I189036,I189407,I189051,I189045,I189452,I189469,I529512,I189486,I529524,I189503,I189529,I189537,I189039,I189033,I189591,I189599,I189048,I189657,I354090,I189683,I189700,I189649,I189722,I354078,I189748,I189756,I189773,I354087,I189790,I354084,I189807,I189824,I354075,I189841,I354081,I189858,I354066,I189875,I189625,I189906,I189923,I189940,I189957,I189637,I189631,I190002,I189646,I189640,I190047,I190064,I354072,I190081,I354069,I190098,I354093,I190124,I190132,I189634,I189628,I190186,I190194,I189643,I190252,I435307,I190278,I190295,I190244,I190317,I435298,I190343,I190351,I190368,I435316,I190385,I435313,I190402,I190419,I435292,I190436,I435295,I190453,I435304,I190470,I190220,I190501,I190518,I190535,I190552,I190232,I190226,I190597,I435310,I190241,I190235,I190642,I190659,I190676,I435301,I190693,I190719,I190727,I190229,I190223,I190781,I190789,I190238,I190847,I877326,I190873,I190890,I190839,I190912,I190938,I190946,I190963,I877329,I190980,I877341,I190997,I191014,I877347,I191031,I877338,I191048,I877344,I191065,I190815,I191096,I191113,I191130,I191147,I190827,I190821,I191192,I877335,I190836,I190830,I191237,I191254,I877332,I191271,I877350,I191288,I191314,I191322,I190824,I190818,I191376,I191384,I190833,I191442,I289636,I191468,I191485,I191507,I289651,I191533,I191541,I191558,I289648,I191575,I191592,I191609,I289645,I191626,I289660,I191643,I289657,I191660,I191691,I191708,I191725,I191742,I191787,I289654,I191832,I191849,I289642,I191866,I289663,I191883,I289639,I191909,I191917,I191971,I191979,I192037,I791712,I192063,I192080,I192029,I192102,I791721,I192128,I192136,I192153,I791709,I192170,I791700,I192187,I192204,I791706,I192221,I791724,I192238,I791697,I192255,I192005,I192286,I192303,I192320,I192337,I192017,I192011,I192382,I791703,I192026,I192020,I192427,I192444,I791715,I192461,I192478,I791718,I192504,I192512,I192014,I192008,I192566,I192574,I192023,I192632,I1035855,I192658,I192675,I192624,I192697,I1035846,I192723,I192731,I192748,I1035840,I192765,I1035834,I192782,I192799,I1035861,I192816,I192833,I1035858,I192850,I192600,I192881,I192898,I192915,I192932,I192612,I192606,I192977,I1035843,I192621,I192615,I193022,I193039,I1035849,I193056,I1035852,I193073,I1035837,I193099,I193107,I192609,I192603,I193161,I193169,I192618,I193227,I214802,I193253,I193270,I193292,I214817,I193318,I193326,I193343,I214814,I193360,I193377,I193394,I214811,I193411,I214826,I193428,I214823,I193445,I193476,I193493,I193510,I193527,I193572,I214820,I193617,I193634,I214808,I193651,I214829,I193668,I214805,I193694,I193702,I193756,I193764,I193822,I1020969,I193848,I193865,I193814,I193887,I1020942,I193913,I193921,I193938,I1020966,I193955,I1020963,I193972,I193989,I194006,I1020960,I194023,I1020948,I194040,I193790,I194071,I194088,I194105,I194122,I193802,I193796,I194167,I1020954,I193811,I193805,I194212,I194229,I1020957,I194246,I1020945,I194263,I1020951,I194289,I194297,I193799,I193793,I194351,I194359,I193808,I194417,I738094,I194443,I194460,I194409,I194482,I738103,I194508,I194516,I194533,I738091,I194550,I738082,I194567,I194584,I738088,I194601,I738106,I194618,I738079,I194635,I194385,I194666,I194683,I194700,I194717,I194397,I194391,I194762,I738085,I194406,I194400,I194807,I194824,I738097,I194841,I194858,I738100,I194884,I194892,I194394,I194388,I194946,I194954,I194403,I195012,I994935,I195038,I195055,I195004,I195077,I994947,I195103,I195111,I195128,I994941,I195145,I994953,I195162,I195179,I994938,I195196,I994950,I195213,I994932,I195230,I194980,I195261,I195278,I195295,I195312,I194992,I194986,I195357,I994944,I195001,I194995,I195402,I195419,I195436,I195453,I994956,I195479,I195487,I194989,I194983,I195541,I195549,I194998,I195607,I365514,I195633,I195650,I195599,I195672,I365502,I195698,I195706,I195723,I365511,I195740,I365508,I195757,I195774,I365499,I195791,I365505,I195808,I365490,I195825,I195575,I195856,I195873,I195890,I195907,I195587,I195581,I195952,I195596,I195590,I195997,I196014,I365496,I196031,I365493,I196048,I365517,I196074,I196082,I195584,I195578,I196136,I196144,I195593,I196202,I196228,I196245,I196194,I196267,I196293,I196301,I196318,I196335,I196352,I196369,I196386,I196403,I196420,I196170,I196451,I196468,I196485,I196502,I196182,I196176,I196547,I196191,I196185,I196592,I196609,I196626,I196643,I196669,I196677,I196179,I196173,I196731,I196739,I196188,I196797,I670221,I196823,I196840,I196789,I196862,I670215,I196888,I196896,I196913,I670233,I196930,I196947,I196964,I196981,I670227,I196998,I670218,I197015,I196765,I197046,I197063,I197080,I197097,I196777,I196771,I197142,I670230,I196786,I196780,I197187,I197204,I670236,I197221,I197238,I670224,I197264,I197272,I196774,I196768,I197326,I197334,I196783,I197392,I514490,I197418,I197435,I197384,I197457,I514487,I197483,I197491,I197508,I514493,I197525,I514478,I197542,I197559,I514481,I197576,I514502,I197593,I514499,I197610,I197360,I197641,I197658,I197675,I197692,I197372,I197366,I197737,I197381,I197375,I197782,I197799,I514484,I197816,I514496,I197833,I197859,I197867,I197369,I197363,I197921,I197929,I197378,I197987,I264340,I198013,I198030,I197979,I198052,I264355,I198078,I198086,I198103,I264352,I198120,I198137,I198154,I264349,I198171,I264364,I198188,I264361,I198205,I197955,I198236,I198253,I198270,I198287,I197967,I197961,I198332,I264358,I197976,I197970,I198377,I198394,I264346,I198411,I264367,I198428,I264343,I198454,I198462,I197964,I197958,I198516,I198524,I197973,I198582,I1000715,I198608,I198625,I198574,I198647,I1000727,I198673,I198681,I198698,I1000721,I198715,I1000733,I198732,I198749,I1000718,I198766,I1000730,I198783,I1000712,I198800,I198550,I198831,I198848,I198865,I198882,I198562,I198556,I198927,I1000724,I198571,I198565,I198972,I198989,I199006,I199023,I1000736,I199049,I199057,I198559,I198553,I199111,I199119,I198568,I199177,I304919,I199203,I199220,I199169,I199242,I304934,I199268,I199276,I199293,I304931,I199310,I199327,I199344,I304928,I199361,I304943,I199378,I304940,I199395,I199145,I199426,I199443,I199460,I199477,I199157,I199151,I199522,I304937,I199166,I199160,I199567,I199584,I304925,I199601,I304946,I199618,I304922,I199644,I199652,I199154,I199148,I199706,I199714,I199163,I199772,I684450,I199798,I199815,I199764,I199837,I684444,I199863,I199871,I199888,I684462,I199905,I199922,I199939,I199956,I684456,I199973,I684447,I199990,I199740,I200021,I200038,I200055,I200072,I199752,I199746,I200117,I684459,I199761,I199755,I200162,I200179,I684465,I200196,I200213,I684453,I200239,I200247,I199749,I199743,I200301,I200309,I199758,I200367,I241679,I200393,I200410,I200359,I200432,I241694,I200458,I200466,I200483,I241691,I200500,I200517,I200534,I241688,I200551,I241703,I200568,I241700,I200585,I200335,I200616,I200633,I200650,I200667,I200347,I200341,I200712,I241697,I200356,I200350,I200757,I200774,I241685,I200791,I241706,I200808,I241682,I200834,I200842,I200344,I200338,I200896,I200904,I200353,I200962,I200988,I201005,I200954,I201027,I201053,I201061,I201078,I201095,I201112,I201129,I201146,I201163,I201180,I200930,I201211,I201228,I201245,I201262,I200942,I200936,I201307,I200951,I200945,I201352,I201369,I201386,I201403,I201429,I201437,I200939,I200933,I201491,I201499,I200948,I201557,I511022,I201583,I201600,I201549,I201622,I511019,I201648,I201656,I201673,I511025,I201690,I511010,I201707,I201724,I511013,I201741,I511034,I201758,I511031,I201775,I201525,I201806,I201823,I201840,I201857,I201537,I201531,I201902,I201546,I201540,I201947,I201964,I511016,I201981,I511028,I201998,I202024,I202032,I201534,I201528,I202086,I202094,I201543,I202152,I350282,I202178,I202195,I202144,I202217,I350270,I202243,I202251,I202268,I350279,I202285,I350276,I202302,I202319,I350267,I202336,I350273,I202353,I350258,I202370,I202120,I202401,I202418,I202435,I202452,I202132,I202126,I202497,I202141,I202135,I202542,I202559,I350264,I202576,I350261,I202593,I350285,I202619,I202627,I202129,I202123,I202681,I202689,I202138,I202747,I333418,I202773,I202790,I202739,I202812,I333406,I202838,I202846,I202863,I333415,I202880,I333412,I202897,I202914,I333403,I202931,I333409,I202948,I333394,I202965,I202715,I202996,I203013,I203030,I203047,I202727,I202721,I203092,I202736,I202730,I203137,I203154,I333400,I203171,I333397,I203188,I333421,I203214,I203222,I202724,I202718,I203276,I203284,I202733,I203342,I203368,I203385,I203334,I203407,I203433,I203441,I203458,I203475,I203492,I203509,I203526,I203543,I203560,I203310,I203591,I203608,I203625,I203642,I203322,I203316,I203687,I203331,I203325,I203732,I203749,I203766,I203783,I203809,I203817,I203319,I203313,I203871,I203879,I203328,I203937,I495419,I203963,I203980,I203929,I204002,I495410,I204028,I204036,I204053,I495428,I204070,I495425,I204087,I204104,I495404,I204121,I495407,I204138,I495416,I204155,I203905,I204186,I204203,I204220,I204237,I203917,I203911,I204282,I495422,I203926,I203920,I204327,I204344,I204361,I495413,I204378,I204404,I204412,I203914,I203908,I204466,I204474,I203923,I204532,I264867,I204558,I204575,I204524,I204597,I264882,I204623,I204631,I204648,I264879,I204665,I204682,I204699,I264876,I204716,I264891,I204733,I264888,I204750,I204500,I204781,I204798,I204815,I204832,I204512,I204506,I204877,I264885,I204521,I204515,I204922,I204939,I264873,I204956,I264894,I204973,I264870,I204999,I205007,I204509,I204503,I205061,I205069,I204518,I205127,I310716,I205153,I205170,I205119,I205192,I310731,I205218,I205226,I205243,I310728,I205260,I205277,I205294,I310725,I205311,I310740,I205328,I310737,I205345,I205095,I205376,I205393,I205410,I205427,I205107,I205101,I205472,I310734,I205116,I205110,I205517,I205534,I310722,I205551,I310743,I205568,I310719,I205594,I205602,I205104,I205098,I205656,I205664,I205113,I205722,I281204,I205748,I205765,I205714,I205787,I281219,I205813,I205821,I205838,I281216,I205855,I205872,I205889,I281213,I205906,I281228,I205923,I281225,I205940,I205690,I205971,I205988,I206005,I206022,I205702,I205696,I206067,I281222,I205711,I205705,I206112,I206129,I281210,I206146,I281231,I206163,I281207,I206189,I206197,I205699,I205693,I206251,I206259,I205708,I206317,I880216,I206343,I206360,I206309,I206382,I206408,I206416,I206433,I880219,I206450,I880231,I206467,I206484,I880237,I206501,I880228,I206518,I880234,I206535,I206285,I206566,I206583,I206600,I206617,I206297,I206291,I206662,I880225,I206306,I206300,I206707,I206724,I880222,I206741,I880240,I206758,I206784,I206792,I206294,I206288,I206846,I206854,I206303,I206912,I754890,I206938,I206955,I206904,I206977,I754899,I207003,I207011,I207028,I754887,I207045,I754878,I207062,I207079,I754884,I207096,I754902,I207113,I754875,I207130,I206880,I207161,I207178,I207195,I207212,I206892,I206886,I207257,I754881,I206901,I206895,I207302,I207319,I754893,I207336,I207353,I754896,I207379,I207387,I206889,I206883,I207441,I207449,I206898,I207507,I671275,I207533,I207550,I207499,I207572,I671269,I207598,I207606,I207623,I671287,I207640,I207657,I207674,I207691,I671281,I207708,I671272,I207725,I207475,I207756,I207773,I207790,I207807,I207487,I207481,I207852,I671284,I207496,I207490,I207897,I207914,I671290,I207931,I207948,I671278,I207974,I207982,I207484,I207478,I208036,I208044,I207493,I208102,I916630,I208128,I208145,I208094,I208167,I208193,I208201,I208218,I916633,I208235,I916645,I208252,I208269,I916651,I208286,I916642,I208303,I916648,I208320,I208070,I208351,I208368,I208385,I208402,I208082,I208076,I208447,I916639,I208091,I208085,I208492,I208509,I916636,I208526,I916654,I208543,I208569,I208577,I208079,I208073,I208631,I208639,I208088,I208697,I1012275,I208723,I208740,I208689,I208762,I1012287,I208788,I208796,I208813,I1012281,I208830,I1012293,I208847,I208864,I1012278,I208881,I1012290,I208898,I1012272,I208915,I208665,I208946,I208963,I208980,I208997,I208677,I208671,I209042,I1012284,I208686,I208680,I209087,I209104,I209121,I209138,I1012296,I209164,I209172,I208674,I208668,I209226,I209234,I208683,I209292,I474033,I209318,I209335,I209284,I209357,I474024,I209383,I209391,I209408,I474042,I209425,I474039,I209442,I209459,I474018,I209476,I474021,I209493,I474030,I209510,I209260,I209541,I209558,I209575,I209592,I209272,I209266,I209637,I474036,I209281,I209275,I209682,I209699,I209716,I474027,I209733,I209759,I209767,I209269,I209263,I209821,I209829,I209278,I209887,I847848,I209913,I209930,I209879,I209952,I209978,I209986,I210003,I847851,I210020,I847863,I210037,I210054,I847869,I210071,I847860,I210088,I847866,I210105,I209855,I210136,I210153,I210170,I210187,I209867,I209861,I210232,I847857,I209876,I209870,I210277,I210294,I847854,I210311,I847872,I210328,I210354,I210362,I209864,I209858,I210416,I210424,I209873,I210482,I380746,I210508,I210525,I210474,I210547,I380734,I210573,I210581,I210598,I380743,I210615,I380740,I210632,I210649,I380731,I210666,I380737,I210683,I380722,I210700,I210450,I210731,I210748,I210765,I210782,I210462,I210456,I210827,I210471,I210465,I210872,I210889,I380728,I210906,I380725,I210923,I380749,I210949,I210957,I210459,I210453,I211011,I211019,I210468,I211077,I651249,I211103,I211120,I211069,I211142,I651243,I211168,I211176,I211193,I651261,I211210,I211227,I211244,I211261,I651255,I211278,I651246,I211295,I211045,I211326,I211343,I211360,I211377,I211057,I211051,I211422,I651258,I211066,I211060,I211467,I211484,I651264,I211501,I211518,I651252,I211544,I211552,I211054,I211048,I211606,I211614,I211063,I211675,I506398,I211701,I211709,I506389,I506404,I211726,I506410,I211752,I211643,I211774,I506395,I211800,I211808,I211825,I211851,I211667,I211873,I211649,I506392,I211913,I211930,I211938,I211955,I211652,I211986,I506386,I506401,I212003,I212029,I212037,I211640,I211658,I212082,I506407,I212099,I211661,I211646,I211655,I211664,I212202,I666002,I212228,I212236,I666005,I665999,I212253,I666011,I212279,I212301,I666014,I212327,I212335,I212352,I212378,I212400,I666017,I212440,I212457,I212465,I212482,I212513,I666008,I212530,I212556,I212564,I212609,I666020,I212626,I212729,I315998,I212755,I212763,I316010,I315989,I212780,I316013,I212806,I212697,I212828,I316004,I212854,I212862,I315986,I212879,I212905,I212721,I212927,I212703,I316001,I212967,I212984,I212992,I213009,I212706,I213040,I315992,I213057,I315995,I213083,I213091,I212694,I212712,I213136,I316007,I213153,I212715,I212700,I212709,I212718,I213256,I982608,I213282,I213290,I982590,I982614,I213307,I982605,I213333,I213224,I213355,I982611,I213381,I213389,I982599,I213406,I213432,I213248,I213454,I213230,I213494,I213511,I213519,I213536,I213233,I213567,I982596,I982593,I213584,I982602,I213610,I213618,I213221,I213239,I213663,I213680,I213242,I213227,I213236,I213245,I213783,I213809,I213817,I213834,I213860,I213751,I213882,I213908,I213916,I213933,I213959,I213775,I213981,I213757,I214021,I214038,I214046,I214063,I213760,I214094,I214111,I214137,I214145,I213748,I213766,I214190,I214207,I213769,I213754,I213763,I213772,I214310,I214336,I214344,I214361,I214387,I214278,I214409,I214435,I214443,I214460,I214486,I214302,I214508,I214284,I214548,I214565,I214573,I214590,I214287,I214621,I214638,I214664,I214672,I214275,I214293,I214717,I214734,I214296,I214281,I214290,I214299,I214837,I597722,I214863,I214871,I597713,I597728,I214888,I597734,I214914,I214936,I597719,I214962,I214970,I214987,I215013,I215035,I597716,I215075,I215092,I215100,I215117,I215148,I597710,I597725,I215165,I215191,I215199,I215244,I597731,I215261,I215364,I326878,I215390,I215398,I326890,I326869,I215415,I326893,I215441,I215332,I215463,I326884,I215489,I215497,I326866,I215514,I215540,I215356,I215562,I215338,I326881,I215602,I215619,I215627,I215644,I215341,I215675,I326872,I215692,I326875,I215718,I215726,I215329,I215347,I215771,I326887,I215788,I215350,I215335,I215344,I215353,I215891,I215917,I215925,I215942,I215968,I215990,I216016,I216024,I216041,I216067,I216089,I216129,I216146,I216154,I216171,I216202,I216219,I216245,I216253,I216298,I216315,I216418,I962480,I216444,I216452,I962462,I962486,I216469,I962477,I216495,I216386,I216517,I962483,I216543,I216551,I962471,I216568,I216594,I216410,I216616,I216392,I216656,I216673,I216681,I216698,I216395,I216729,I962468,I962465,I216746,I962474,I216772,I216780,I216383,I216401,I216825,I216842,I216404,I216389,I216398,I216407,I216945,I499462,I216971,I216979,I499453,I499468,I216996,I499474,I217022,I217044,I499459,I217070,I217078,I217095,I217121,I217143,I499456,I217183,I217200,I217208,I217225,I217256,I499450,I499465,I217273,I217299,I217307,I217352,I499471,I217369,I217472,I396705,I217498,I217506,I396717,I217523,I396702,I217549,I217440,I217571,I396726,I217597,I217605,I396723,I217622,I217648,I217464,I217670,I217446,I396714,I217710,I217727,I217735,I217752,I217449,I217783,I396711,I217800,I396720,I217826,I217834,I217437,I217455,I217879,I396708,I217896,I217458,I217443,I217452,I217461,I217999,I1015755,I218025,I218033,I1015752,I1015743,I218050,I1015740,I218076,I217967,I218098,I1015749,I218124,I218132,I1015758,I218149,I218175,I217991,I218197,I217973,I1015761,I218237,I218254,I218262,I218279,I217976,I218310,I1015746,I218327,I1015764,I218353,I218361,I217964,I217982,I218406,I218423,I217985,I217970,I217979,I217988,I218526,I950154,I218552,I218560,I950169,I218577,I950172,I218603,I218494,I218625,I950178,I218651,I218659,I950160,I218676,I218702,I218518,I218724,I218500,I950157,I218764,I218781,I218789,I218806,I218503,I218837,I950163,I218854,I950175,I218880,I218888,I218491,I218509,I218933,I950166,I218950,I218512,I218497,I218506,I218515,I219053,I476923,I219079,I219087,I476908,I476911,I219104,I476926,I219130,I219152,I476920,I219178,I219186,I219203,I219229,I219251,I476917,I219291,I219308,I219316,I219333,I219364,I476932,I219381,I476929,I219407,I219415,I219460,I476914,I219477,I219580,I755524,I219606,I219614,I755521,I755539,I219631,I755530,I219657,I219548,I219679,I755545,I219705,I219713,I755527,I219730,I219756,I219572,I219778,I219554,I755533,I219818,I219835,I219843,I219860,I219557,I219891,I755548,I219908,I755536,I219934,I219942,I219545,I219563,I219987,I755542,I220004,I219566,I219551,I219560,I219569,I220107,I336670,I220133,I220141,I336682,I336661,I220158,I336685,I220184,I220075,I220206,I336676,I220232,I220240,I336658,I220257,I220283,I220099,I220305,I220081,I336673,I220345,I220362,I220370,I220387,I220084,I220418,I336664,I220435,I336667,I220461,I220469,I220072,I220090,I220514,I336679,I220531,I220093,I220078,I220087,I220096,I220634,I220660,I220668,I220685,I220711,I220602,I220733,I220759,I220767,I220784,I220810,I220626,I220832,I220608,I220872,I220889,I220897,I220914,I220611,I220945,I220962,I220988,I220996,I220599,I220617,I221041,I221058,I220620,I220605,I220614,I220623,I221161,I1062630,I221187,I221195,I1062609,I221212,I1062636,I221238,I221129,I221260,I1062624,I221286,I221294,I1062627,I221311,I221337,I221153,I221359,I221135,I1062618,I221399,I221416,I221424,I221441,I221138,I221472,I1062615,I1062612,I221489,I1062633,I221515,I221523,I221126,I221144,I221568,I1062621,I221585,I221147,I221132,I221141,I221150,I221688,I740666,I221714,I221722,I740663,I740681,I221739,I740672,I221765,I221656,I221787,I740687,I221813,I221821,I740669,I221838,I221864,I221680,I221886,I221662,I740675,I221926,I221943,I221951,I221968,I221665,I221999,I740690,I222016,I740678,I222042,I222050,I221653,I221671,I222095,I740684,I222112,I221674,I221659,I221668,I221677,I222215,I222241,I222249,I222266,I222292,I222183,I222314,I222340,I222348,I222365,I222391,I222207,I222413,I222189,I222453,I222470,I222478,I222495,I222192,I222526,I222543,I222569,I222577,I222180,I222198,I222622,I222639,I222201,I222186,I222195,I222204,I222742,I222768,I222776,I222793,I222819,I222710,I222841,I222867,I222875,I222892,I222918,I222734,I222940,I222716,I222980,I222997,I223005,I223022,I222719,I223053,I223070,I223096,I223104,I222707,I222725,I223149,I223166,I222728,I222713,I222722,I222731,I223269,I578648,I223295,I223303,I578639,I578654,I223320,I578660,I223346,I223237,I223368,I578645,I223394,I223402,I223419,I223445,I223261,I223467,I223243,I578642,I223507,I223524,I223532,I223549,I223246,I223580,I578636,I578651,I223597,I223623,I223631,I223234,I223252,I223676,I578657,I223693,I223255,I223240,I223249,I223258,I223796,I391070,I223822,I223830,I391082,I391061,I223847,I391085,I223873,I223764,I223895,I391076,I223921,I223929,I391058,I223946,I223972,I223788,I223994,I223770,I391073,I224034,I224051,I224059,I224076,I223773,I224107,I391064,I224124,I391067,I224150,I224158,I223761,I223779,I224203,I391079,I224220,I223782,I223767,I223776,I223785,I224323,I224349,I224357,I224374,I224400,I224291,I224422,I224448,I224456,I224473,I224499,I224315,I224521,I224297,I224561,I224578,I224586,I224603,I224300,I224634,I224651,I224677,I224685,I224288,I224306,I224730,I224747,I224309,I224294,I224303,I224312,I224850,I592520,I224876,I224884,I592511,I592526,I224901,I592532,I224927,I224818,I224949,I592517,I224975,I224983,I225000,I225026,I224842,I225048,I224824,I592514,I225088,I225105,I225113,I225130,I224827,I225161,I592508,I592523,I225178,I225204,I225212,I224815,I224833,I225257,I592529,I225274,I224836,I224821,I224830,I224839,I225377,I1002461,I225403,I225411,I1002458,I1002449,I225428,I1002446,I225454,I225345,I225476,I1002455,I225502,I225510,I1002464,I225527,I225553,I225369,I225575,I225351,I1002467,I225615,I225632,I225640,I225657,I225354,I225688,I1002452,I225705,I1002470,I225731,I225739,I225342,I225360,I225784,I225801,I225363,I225348,I225357,I225366,I225904,I819223,I225930,I225938,I819220,I225955,I819232,I225981,I226003,I226029,I226037,I819238,I226054,I226080,I226102,I819226,I226142,I226159,I226167,I226184,I226215,I819235,I819241,I226232,I226258,I226266,I226311,I819229,I226328,I226431,I226457,I226465,I226482,I226508,I226530,I226556,I226564,I226581,I226607,I226629,I226669,I226686,I226694,I226711,I226742,I226759,I226785,I226793,I226838,I226855,I226958,I226984,I226992,I227009,I227035,I226926,I227057,I227083,I227091,I227108,I227134,I226950,I227156,I226932,I227196,I227213,I227221,I227238,I226935,I227269,I227286,I227312,I227320,I226923,I226941,I227365,I227382,I226944,I226929,I226938,I226947,I227485,I545124,I227511,I227519,I545115,I545130,I227536,I545136,I227562,I227453,I227584,I545121,I227610,I227618,I227635,I227661,I227477,I227683,I227459,I545118,I227723,I227740,I227748,I227765,I227462,I227796,I545112,I545127,I227813,I227839,I227847,I227450,I227468,I227892,I545133,I227909,I227471,I227456,I227465,I227474,I228012,I900446,I228038,I228046,I900461,I228063,I900464,I228089,I227980,I228111,I900470,I228137,I228145,I900452,I228162,I228188,I228004,I228210,I227986,I900449,I228250,I228267,I228275,I228292,I227989,I228323,I900455,I228340,I900467,I228366,I228374,I227977,I227995,I228419,I900458,I228436,I227998,I227983,I227992,I228001,I228539,I228565,I228573,I228590,I228616,I228638,I228664,I228672,I228689,I228715,I228737,I228777,I228794,I228802,I228819,I228850,I228867,I228893,I228901,I228946,I228963,I229066,I418720,I229092,I229100,I418732,I229117,I418717,I229143,I229034,I229165,I418741,I229191,I229199,I418738,I229216,I229242,I229058,I229264,I229040,I418729,I229304,I229321,I229329,I229346,I229043,I229377,I418726,I229394,I418735,I229420,I229428,I229031,I229049,I229473,I418723,I229490,I229052,I229037,I229046,I229055,I229593,I806320,I229619,I229627,I806317,I229644,I806329,I229670,I229692,I229718,I229726,I806335,I229743,I229769,I229791,I806323,I229831,I229848,I229856,I229873,I229904,I806332,I806338,I229921,I229947,I229955,I230000,I806326,I230017,I230120,I498884,I230146,I230154,I498875,I498890,I230171,I498896,I230197,I230088,I230219,I498881,I230245,I230253,I230270,I230296,I230112,I230318,I230094,I498878,I230358,I230375,I230383,I230400,I230097,I230431,I498872,I498887,I230448,I230474,I230482,I230085,I230103,I230527,I498893,I230544,I230106,I230091,I230100,I230109,I230647,I878482,I230673,I230681,I878497,I230698,I878500,I230724,I230615,I230746,I878506,I230772,I230780,I878488,I230797,I230823,I230639,I230845,I230621,I878485,I230885,I230902,I230910,I230927,I230624,I230958,I878491,I230975,I878503,I231001,I231009,I230612,I230630,I231054,I878494,I231071,I230633,I230618,I230627,I230636,I231174,I231200,I231208,I231225,I231251,I231142,I231273,I231299,I231307,I231324,I231350,I231166,I231372,I231148,I231412,I231429,I231437,I231454,I231151,I231485,I231502,I231528,I231536,I231139,I231157,I231581,I231598,I231160,I231145,I231154,I231163,I231701,I845536,I231727,I231735,I845551,I231752,I845554,I231778,I231669,I231800,I845560,I231826,I231834,I845542,I231851,I231877,I231693,I231899,I231675,I845539,I231939,I231956,I231964,I231981,I231678,I232012,I845545,I232029,I845557,I232055,I232063,I231666,I231684,I232108,I845548,I232125,I231687,I231672,I231681,I231690,I232228,I645449,I232254,I232262,I645452,I645446,I232279,I645458,I232305,I232196,I232327,I645461,I232353,I232361,I232378,I232404,I232220,I232426,I232202,I645464,I232466,I232483,I232491,I232508,I232205,I232539,I645455,I232556,I232582,I232590,I232193,I232211,I232635,I645467,I232652,I232214,I232199,I232208,I232217,I232755,I723870,I232781,I232789,I723867,I723885,I232806,I723876,I232832,I232723,I232854,I723891,I232880,I232888,I723873,I232905,I232931,I232747,I232953,I232729,I723879,I232993,I233010,I233018,I233035,I232732,I233066,I723894,I233083,I723882,I233109,I233117,I232720,I232738,I233162,I723888,I233179,I232741,I232726,I232735,I232744,I233282,I997837,I233308,I233316,I997834,I997825,I233333,I997822,I233359,I233250,I233381,I997831,I233407,I233415,I997840,I233432,I233458,I233274,I233480,I233256,I997843,I233520,I233537,I233545,I233562,I233259,I233593,I997828,I233610,I997846,I233636,I233644,I233247,I233265,I233689,I233706,I233268,I233253,I233262,I233271,I233809,I667056,I233835,I233843,I667059,I667053,I233860,I667065,I233886,I233777,I233908,I667068,I233934,I233942,I233959,I233985,I233801,I234007,I233783,I667071,I234047,I234064,I234072,I234089,I233786,I234120,I667062,I234137,I234163,I234171,I233774,I233792,I234216,I667074,I234233,I233795,I233780,I233789,I233798,I234336,I1044185,I234362,I234370,I1044164,I234387,I1044191,I234413,I234435,I1044179,I234461,I234469,I1044182,I234486,I234512,I234534,I1044173,I234574,I234591,I234599,I234616,I234647,I1044170,I1044167,I234664,I1044188,I234690,I234698,I234743,I1044176,I234760,I234863,I479813,I234889,I234897,I479798,I479801,I234914,I479816,I234940,I234831,I234962,I479810,I234988,I234996,I235013,I235039,I234855,I235061,I234837,I479807,I235101,I235118,I235126,I235143,I234840,I235174,I479822,I235191,I479819,I235217,I235225,I234828,I234846,I235270,I479804,I235287,I234849,I234834,I234843,I234852,I235390,I1078695,I235416,I235424,I1078674,I235441,I1078701,I235467,I235358,I235489,I1078689,I235515,I235523,I1078692,I235540,I235566,I235382,I235588,I235364,I1078683,I235628,I235645,I235653,I235670,I235367,I235701,I1078680,I1078677,I235718,I1078698,I235744,I235752,I235355,I235373,I235797,I1078686,I235814,I235376,I235361,I235370,I235379,I235917,I235943,I235951,I235968,I235994,I235885,I236016,I236042,I236050,I236067,I236093,I235909,I236115,I235891,I236155,I236172,I236180,I236197,I235894,I236228,I236245,I236271,I236279,I235882,I235900,I236324,I236341,I235903,I235888,I235897,I235906,I236444,I660732,I236470,I236478,I660735,I660729,I236495,I660741,I236521,I236412,I236543,I660744,I236569,I236577,I236594,I236620,I236436,I236642,I236418,I660747,I236682,I236699,I236707,I236724,I236421,I236755,I660738,I236772,I236798,I236806,I236409,I236427,I236851,I660750,I236868,I236430,I236415,I236424,I236433,I236971,I369854,I236997,I237005,I369866,I369845,I237022,I369869,I237048,I237070,I369860,I237096,I237104,I369842,I237121,I237147,I237169,I369857,I237209,I237226,I237234,I237251,I237282,I369848,I237299,I369851,I237325,I237333,I237378,I369863,I237395,I237498,I389982,I237524,I237532,I389994,I389973,I237549,I389997,I237575,I237597,I389988,I237623,I237631,I389970,I237648,I237674,I237696,I389985,I237736,I237753,I237761,I237778,I237809,I389976,I237826,I389979,I237852,I237860,I237905,I389991,I237922,I238025,I238051,I238059,I238076,I238102,I237993,I238124,I238150,I238158,I238175,I238201,I238017,I238223,I237999,I238263,I238280,I238288,I238305,I238002,I238336,I238353,I238379,I238387,I237990,I238008,I238432,I238449,I238011,I237996,I238005,I238014,I238552,I238578,I238586,I238603,I238629,I238520,I238651,I238677,I238685,I238702,I238728,I238544,I238750,I238526,I238790,I238807,I238815,I238832,I238529,I238863,I238880,I238906,I238914,I238517,I238535,I238959,I238976,I238538,I238523,I238532,I238541,I239079,I805198,I239105,I239113,I805195,I239130,I805207,I239156,I239047,I239178,I239204,I239212,I805213,I239229,I239255,I239071,I239277,I239053,I805201,I239317,I239334,I239342,I239359,I239056,I239390,I805210,I805216,I239407,I239433,I239441,I239044,I239062,I239486,I805204,I239503,I239065,I239050,I239059,I239068,I239606,I589630,I239632,I239640,I589621,I589636,I239657,I589642,I239683,I239574,I239705,I589627,I239731,I239739,I239756,I239782,I239598,I239804,I239580,I589624,I239844,I239861,I239869,I239886,I239583,I239917,I589618,I589633,I239934,I239960,I239968,I239571,I239589,I240013,I589639,I240030,I239592,I239577,I239586,I239595,I240133,I240159,I240167,I240184,I240210,I240101,I240232,I240258,I240266,I240283,I240309,I240125,I240331,I240107,I240371,I240388,I240396,I240413,I240110,I240444,I240461,I240487,I240495,I240098,I240116,I240540,I240557,I240119,I240104,I240113,I240122,I240660,I494841,I240686,I240694,I494826,I494829,I240711,I494844,I240737,I240759,I494838,I240785,I240793,I240810,I240836,I240858,I494835,I240898,I240915,I240923,I240940,I240971,I494850,I240988,I494847,I241014,I241022,I241067,I494832,I241084,I241187,I640706,I241213,I241221,I640709,I640703,I241238,I640715,I241264,I241155,I241286,I640718,I241312,I241320,I241337,I241363,I241179,I241385,I241161,I640721,I241425,I241442,I241450,I241467,I241164,I241498,I640712,I241515,I241541,I241549,I241152,I241170,I241594,I640724,I241611,I241173,I241158,I241167,I241176,I241714,I325790,I241740,I241748,I325802,I325781,I241765,I325805,I241791,I241813,I325796,I241839,I241847,I325778,I241864,I241890,I241912,I325793,I241952,I241969,I241977,I241994,I242025,I325784,I242042,I325787,I242068,I242076,I242121,I325799,I242138,I242241,I391614,I242267,I242275,I391626,I391605,I242292,I391629,I242318,I242209,I242340,I391620,I242366,I242374,I391602,I242391,I242417,I242233,I242439,I242215,I391617,I242479,I242496,I242504,I242521,I242218,I242552,I391608,I242569,I391611,I242595,I242603,I242206,I242224,I242648,I391623,I242665,I242227,I242212,I242221,I242230,I242768,I696041,I242794,I242802,I696044,I696038,I242819,I696050,I242845,I242736,I242867,I696053,I242893,I242901,I242918,I242944,I242760,I242966,I242742,I696056,I243006,I243023,I243031,I243048,I242745,I243079,I696047,I243096,I243122,I243130,I242733,I242751,I243175,I696059,I243192,I242754,I242739,I242748,I242757,I243295,I243321,I243329,I243346,I243372,I243394,I243420,I243428,I243445,I243471,I243493,I243533,I243550,I243558,I243575,I243606,I243623,I243649,I243657,I243702,I243719,I243822,I537610,I243848,I243856,I537601,I537616,I243873,I537622,I243899,I243790,I243921,I537607,I243947,I243955,I243972,I243998,I243814,I244020,I243796,I537604,I244060,I244077,I244085,I244102,I243799,I244133,I537598,I537613,I244150,I244176,I244184,I243787,I243805,I244229,I537619,I244246,I243808,I243793,I243802,I243811,I244349,I244375,I244383,I244400,I244426,I244448,I244474,I244482,I244499,I244525,I244547,I244587,I244604,I244612,I244629,I244660,I244677,I244703,I244711,I244756,I244773,I244876,I564198,I244902,I244910,I564189,I564204,I244927,I564210,I244953,I244844,I244975,I564195,I245001,I245009,I245026,I245052,I244868,I245074,I244850,I564192,I245114,I245131,I245139,I245156,I244853,I245187,I564186,I564201,I245204,I245230,I245238,I244841,I244859,I245283,I564207,I245300,I244862,I244847,I244856,I244865,I245403,I245429,I245437,I245454,I245480,I245371,I245502,I245528,I245536,I245553,I245579,I245395,I245601,I245377,I245641,I245658,I245666,I245683,I245380,I245714,I245731,I245757,I245765,I245368,I245386,I245810,I245827,I245389,I245374,I245383,I245392,I245930,I245956,I245964,I245981,I246007,I245898,I246029,I246055,I246063,I246080,I246106,I245922,I246128,I245904,I246168,I246185,I246193,I246210,I245907,I246241,I246258,I246284,I246292,I245895,I245913,I246337,I246354,I245916,I245901,I245910,I245919,I246457,I951888,I246483,I246491,I951903,I246508,I951906,I246534,I246425,I246556,I951912,I246582,I246590,I951894,I246607,I246633,I246449,I246655,I246431,I951891,I246695,I246712,I246720,I246737,I246434,I246768,I951897,I246785,I951909,I246811,I246819,I246422,I246440,I246864,I951900,I246881,I246443,I246428,I246437,I246446,I246984,I1101305,I247010,I247018,I1101284,I247035,I1101311,I247061,I246952,I247083,I1101299,I247109,I247117,I1101302,I247134,I247160,I246976,I247182,I246958,I1101293,I247222,I247239,I247247,I247264,I246961,I247295,I1101290,I1101287,I247312,I1101308,I247338,I247346,I246949,I246967,I247391,I1101296,I247408,I246970,I246955,I246964,I246973,I247511,I419315,I247537,I247545,I419327,I247562,I419312,I247588,I247479,I247610,I419336,I247636,I247644,I419333,I247661,I247687,I247503,I247709,I247485,I419324,I247749,I247766,I247774,I247791,I247488,I247822,I419321,I247839,I419330,I247865,I247873,I247476,I247494,I247918,I419318,I247935,I247497,I247482,I247491,I247500,I248038,I876748,I248064,I248072,I876763,I248089,I876766,I248115,I248006,I248137,I876772,I248163,I248171,I876754,I248188,I248214,I248030,I248236,I248012,I876751,I248276,I248293,I248301,I248318,I248015,I248349,I876757,I248366,I876769,I248392,I248400,I248003,I248021,I248445,I876760,I248462,I248024,I248009,I248018,I248027,I248565,I949576,I248591,I248599,I949591,I248616,I949594,I248642,I248533,I248664,I949600,I248690,I248698,I949582,I248715,I248741,I248557,I248763,I248539,I949579,I248803,I248820,I248828,I248845,I248542,I248876,I949585,I248893,I949597,I248919,I248927,I248530,I248548,I248972,I949588,I248989,I248551,I248536,I248545,I248554,I249092,I605814,I249118,I249126,I605805,I605820,I249143,I605826,I249169,I249060,I249191,I605811,I249217,I249225,I249242,I249268,I249084,I249290,I249066,I605808,I249330,I249347,I249355,I249372,I249069,I249403,I605802,I605817,I249420,I249446,I249454,I249057,I249075,I249499,I605823,I249516,I249078,I249063,I249072,I249081,I249619,I722578,I249645,I249653,I722575,I722593,I249670,I722584,I249696,I249587,I249718,I722599,I249744,I249752,I722581,I249769,I249795,I249611,I249817,I249593,I722587,I249857,I249874,I249882,I249899,I249596,I249930,I722602,I249947,I722590,I249973,I249981,I249584,I249602,I250026,I722596,I250043,I249605,I249590,I249599,I249608,I250146,I924722,I250172,I250180,I924737,I250197,I924740,I250223,I250114,I250245,I924746,I250271,I250279,I924728,I250296,I250322,I250138,I250344,I250120,I924725,I250384,I250401,I250409,I250426,I250123,I250457,I924731,I250474,I924743,I250500,I250508,I250111,I250129,I250553,I924734,I250570,I250132,I250117,I250126,I250135,I250673,I792346,I250699,I250707,I792343,I792361,I250724,I792352,I250750,I250641,I250772,I792367,I250798,I250806,I792349,I250823,I250849,I250665,I250871,I250647,I792355,I250911,I250928,I250936,I250953,I250650,I250984,I792370,I251001,I792358,I251027,I251035,I250638,I250656,I251080,I792364,I251097,I250659,I250644,I250653,I250662,I251200,I610438,I251226,I251234,I610429,I610444,I251251,I610450,I251277,I251299,I610435,I251325,I251333,I251350,I251376,I251398,I610432,I251438,I251455,I251463,I251480,I251511,I610426,I610441,I251528,I251554,I251562,I251607,I610447,I251624,I251727,I251753,I251761,I251778,I251804,I251695,I251826,I251852,I251860,I251877,I251903,I251719,I251925,I251701,I251965,I251982,I251990,I252007,I251704,I252038,I252055,I252081,I252089,I251692,I251710,I252134,I252151,I251713,I251698,I251707,I251716,I252254,I568244,I252280,I252288,I568235,I568250,I252305,I568256,I252331,I252222,I252353,I568241,I252379,I252387,I252404,I252430,I252246,I252452,I252228,I568238,I252492,I252509,I252517,I252534,I252231,I252565,I568232,I568247,I252582,I252608,I252616,I252219,I252237,I252661,I568253,I252678,I252240,I252225,I252234,I252243,I252781,I487905,I252807,I252815,I487890,I487893,I252832,I487908,I252858,I252749,I252880,I487902,I252906,I252914,I252931,I252957,I252773,I252979,I252755,I487899,I253019,I253036,I253044,I253061,I252758,I253092,I487914,I253109,I487911,I253135,I253143,I252746,I252764,I253188,I487896,I253205,I252767,I252752,I252761,I252770,I253308,I507554,I253334,I253342,I507545,I507560,I253359,I507566,I253385,I253276,I253407,I507551,I253433,I253441,I253458,I253484,I253300,I253506,I253282,I507548,I253546,I253563,I253571,I253588,I253285,I253619,I507542,I507557,I253636,I253662,I253670,I253273,I253291,I253715,I507563,I253732,I253294,I253279,I253288,I253297,I253835,I721286,I253861,I253869,I721283,I721301,I253886,I721292,I253912,I253803,I253934,I721307,I253960,I253968,I721289,I253985,I254011,I253827,I254033,I253809,I721295,I254073,I254090,I254098,I254115,I253812,I254146,I721310,I254163,I721298,I254189,I254197,I253800,I253818,I254242,I721304,I254259,I253821,I253806,I253815,I253824,I254362,I658624,I254388,I254396,I658627,I658621,I254413,I658633,I254439,I254330,I254461,I658636,I254487,I254495,I254512,I254538,I254354,I254560,I254336,I658639,I254600,I254617,I254625,I254642,I254339,I254673,I658630,I254690,I254716,I254724,I254327,I254345,I254769,I658642,I254786,I254348,I254333,I254342,I254351,I254889,I531252,I254915,I254923,I531243,I531258,I254940,I531264,I254966,I254988,I531249,I255014,I255022,I255039,I255065,I255087,I531246,I255127,I255144,I255152,I255169,I255200,I531240,I531255,I255217,I255243,I255251,I255296,I531261,I255313,I255416,I971728,I255442,I255450,I971710,I971734,I255467,I971725,I255493,I255384,I255515,I971731,I255541,I255549,I971719,I255566,I255592,I255408,I255614,I255390,I255654,I255671,I255679,I255696,I255393,I255727,I971716,I971713,I255744,I971722,I255770,I255778,I255381,I255399,I255823,I255840,I255402,I255387,I255396,I255405,I255943,I641760,I255969,I255977,I641763,I641757,I255994,I641769,I256020,I255911,I256042,I641772,I256068,I256076,I256093,I256119,I255935,I256141,I255917,I641775,I256181,I256198,I256206,I256223,I255920,I256254,I641766,I256271,I256297,I256305,I255908,I255926,I256350,I641778,I256367,I255929,I255914,I255923,I255932,I256470,I579226,I256496,I256504,I579217,I579232,I256521,I579238,I256547,I256438,I256569,I579223,I256595,I256603,I256620,I256646,I256462,I256668,I256444,I579220,I256708,I256725,I256733,I256750,I256447,I256781,I579214,I579229,I256798,I256824,I256832,I256435,I256453,I256877,I579235,I256894,I256456,I256441,I256450,I256459,I256997,I257023,I257031,I257048,I257074,I256965,I257096,I257122,I257130,I257147,I257173,I256989,I257195,I256971,I257235,I257252,I257260,I257277,I256974,I257308,I257325,I257351,I257359,I256962,I256980,I257404,I257421,I256983,I256968,I256977,I256986,I257524,I882528,I257550,I257558,I882543,I257575,I882546,I257601,I257492,I257623,I882552,I257649,I257657,I882534,I257674,I257700,I257516,I257722,I257498,I882531,I257762,I257779,I257787,I257804,I257501,I257835,I882537,I257852,I882549,I257878,I257886,I257489,I257507,I257931,I882540,I257948,I257510,I257495,I257504,I257513,I258051,I571712,I258077,I258085,I571703,I571718,I258102,I571724,I258128,I258150,I571709,I258176,I258184,I258201,I258227,I258249,I571706,I258289,I258306,I258314,I258331,I258362,I571700,I571715,I258379,I258405,I258413,I258458,I571721,I258475,I258578,I603502,I258604,I258612,I603493,I603508,I258629,I603514,I258655,I258677,I603499,I258703,I258711,I258728,I258754,I258776,I603496,I258816,I258833,I258841,I258858,I258889,I603490,I603505,I258906,I258932,I258940,I258985,I603511,I259002,I259105,I818662,I259131,I259139,I818659,I259156,I818671,I259182,I259204,I259230,I259238,I818677,I259255,I259281,I259303,I818665,I259343,I259360,I259368,I259385,I259416,I818674,I818680,I259433,I259459,I259467,I259512,I818668,I259529,I259632,I392158,I259658,I259666,I392170,I392149,I259683,I392173,I259709,I259600,I259731,I392164,I259757,I259765,I392146,I259782,I259808,I259624,I259830,I259606,I392161,I259870,I259887,I259895,I259912,I259609,I259943,I392152,I259960,I392155,I259986,I259994,I259597,I259615,I260039,I392167,I260056,I259618,I259603,I259612,I259621,I260159,I1057275,I260185,I260193,I1057254,I260210,I1057281,I260236,I260127,I260258,I1057269,I260284,I260292,I1057272,I260309,I260335,I260151,I260357,I260133,I1057263,I260397,I260414,I260422,I260439,I260136,I260470,I1057260,I1057257,I260487,I1057278,I260513,I260521,I260124,I260142,I260566,I1057266,I260583,I260145,I260130,I260139,I260148,I260686,I802954,I260712,I260720,I802951,I260737,I802963,I260763,I260654,I260785,I260811,I260819,I802969,I260836,I260862,I260678,I260884,I260660,I802957,I260924,I260941,I260949,I260966,I260663,I260997,I802966,I802972,I261014,I261040,I261048,I260651,I260669,I261093,I802960,I261110,I260672,I260657,I260666,I260675,I261213,I261239,I261247,I261264,I261290,I261181,I261312,I261338,I261346,I261363,I261389,I261205,I261411,I261187,I261451,I261468,I261476,I261493,I261190,I261524,I261541,I261567,I261575,I261178,I261196,I261620,I261637,I261199,I261184,I261193,I261202,I261740,I458427,I261766,I261774,I458412,I458415,I261791,I458430,I261817,I261708,I261839,I458424,I261865,I261873,I261890,I261916,I261732,I261938,I261714,I458421,I261978,I261995,I262003,I262020,I261717,I262051,I458436,I262068,I458433,I262094,I262102,I261705,I261723,I262147,I458418,I262164,I261726,I261711,I261720,I261729,I262267,I387262,I262293,I262301,I387274,I387253,I262318,I387277,I262344,I262235,I262366,I387268,I262392,I262400,I387250,I262417,I262443,I262259,I262465,I262241,I387265,I262505,I262522,I262530,I262547,I262244,I262578,I387256,I262595,I387259,I262621,I262629,I262232,I262250,I262674,I387271,I262691,I262253,I262238,I262247,I262256,I262794,I262820,I262828,I262845,I262871,I262893,I262919,I262927,I262944,I262970,I262992,I263032,I263049,I263057,I263074,I263105,I263122,I263148,I263156,I263201,I263218,I263321,I734206,I263347,I263355,I734203,I734221,I263372,I734212,I263398,I263420,I734227,I263446,I263454,I734209,I263471,I263497,I263519,I734215,I263559,I263576,I263584,I263601,I263632,I734230,I263649,I734218,I263675,I263683,I263728,I734224,I263745,I263848,I741312,I263874,I263882,I741309,I741327,I263899,I741318,I263925,I263816,I263947,I741333,I263973,I263981,I741315,I263998,I264024,I263840,I264046,I263822,I741321,I264086,I264103,I264111,I264128,I263825,I264159,I741336,I264176,I741324,I264202,I264210,I263813,I263831,I264255,I741330,I264272,I263834,I263819,I263828,I263837,I264375,I501196,I264401,I264409,I501187,I501202,I264426,I501208,I264452,I264474,I501193,I264500,I264508,I264525,I264551,I264573,I501190,I264613,I264630,I264638,I264655,I264686,I501184,I501199,I264703,I264729,I264737,I264782,I501205,I264799,I264902,I264928,I264936,I264953,I264979,I265001,I265027,I265035,I265052,I265078,I265100,I265140,I265157,I265165,I265182,I265213,I265230,I265256,I265264,I265309,I265326,I265429,I265455,I265463,I265480,I265506,I265397,I265528,I265554,I265562,I265579,I265605,I265421,I265627,I265403,I265667,I265684,I265692,I265709,I265406,I265740,I265757,I265783,I265791,I265394,I265412,I265836,I265853,I265415,I265400,I265409,I265418,I265956,I807442,I265982,I265990,I807439,I266007,I807451,I266033,I265924,I266055,I266081,I266089,I807457,I266106,I266132,I265948,I266154,I265930,I807445,I266194,I266211,I266219,I266236,I265933,I266267,I807454,I807460,I266284,I266310,I266318,I265921,I265939,I266363,I807448,I266380,I265942,I265927,I265936,I265945,I266483,I778134,I266509,I266517,I778131,I778149,I266534,I778140,I266560,I266451,I266582,I778155,I266608,I266616,I778137,I266633,I266659,I266475,I266681,I266457,I778143,I266721,I266738,I266746,I266763,I266460,I266794,I778158,I266811,I778146,I266837,I266845,I266448,I266466,I266890,I778152,I266907,I266469,I266454,I266463,I266472,I267010,I567666,I267036,I267044,I567657,I567672,I267061,I567678,I267087,I266978,I267109,I567663,I267135,I267143,I267160,I267186,I267002,I267208,I266984,I567660,I267248,I267265,I267273,I267290,I266987,I267321,I567654,I567669,I267338,I267364,I267372,I266975,I266993,I267417,I567675,I267434,I266996,I266981,I266990,I266999,I267537,I791054,I267563,I267571,I791051,I791069,I267588,I791060,I267614,I267505,I267636,I791075,I267662,I267670,I791057,I267687,I267713,I267529,I267735,I267511,I791063,I267775,I267792,I267800,I267817,I267514,I267848,I791078,I267865,I791066,I267891,I267899,I267502,I267520,I267944,I791072,I267961,I267523,I267508,I267517,I267526,I268064,I1084645,I268090,I268098,I1084624,I268115,I1084651,I268141,I268163,I1084639,I268189,I268197,I1084642,I268214,I268240,I268262,I1084633,I268302,I268319,I268327,I268344,I268375,I1084630,I1084627,I268392,I1084648,I268418,I268426,I268471,I1084636,I268488,I268591,I1037640,I268617,I268625,I1037619,I268642,I1037646,I268668,I268559,I268690,I1037634,I268716,I268724,I1037637,I268741,I268767,I268583,I268789,I268565,I1037628,I268829,I268846,I268854,I268871,I268568,I268902,I1037625,I1037622,I268919,I1037643,I268945,I268953,I268556,I268574,I268998,I1037631,I269015,I268577,I268562,I268571,I268580,I269118,I972272,I269144,I269152,I972254,I972278,I269169,I972269,I269195,I269217,I972275,I269243,I269251,I972263,I269268,I269294,I269316,I269356,I269373,I269381,I269398,I269429,I972260,I972257,I269446,I972266,I269472,I269480,I269525,I269542,I269645,I634909,I269671,I269679,I634912,I634906,I269696,I634918,I269722,I269613,I269744,I634921,I269770,I269778,I269795,I269821,I269637,I269843,I269619,I634924,I269883,I269900,I269908,I269925,I269622,I269956,I634915,I269973,I269999,I270007,I269610,I269628,I270052,I634927,I270069,I269631,I269616,I269625,I269634,I270172,I339390,I270198,I270206,I339402,I339381,I270223,I339405,I270249,I270140,I270271,I339396,I270297,I270305,I339378,I270322,I270348,I270164,I270370,I270146,I339393,I270410,I270427,I270435,I270452,I270149,I270483,I339384,I270500,I339387,I270526,I270534,I270137,I270155,I270579,I339399,I270596,I270158,I270143,I270152,I270161,I270699,I479235,I270725,I270733,I479220,I479223,I270750,I479238,I270776,I270667,I270798,I479232,I270824,I270832,I270849,I270875,I270691,I270897,I270673,I479229,I270937,I270954,I270962,I270979,I270676,I271010,I479244,I271027,I479241,I271053,I271061,I270664,I270682,I271106,I479226,I271123,I270685,I270670,I270679,I270688,I271226,I440509,I271252,I271260,I440494,I440497,I271277,I440512,I271303,I271194,I271325,I440506,I271351,I271359,I271376,I271402,I271218,I271424,I271200,I440503,I271464,I271481,I271489,I271506,I271203,I271537,I440518,I271554,I440515,I271580,I271588,I271191,I271209,I271633,I440500,I271650,I271212,I271197,I271206,I271215,I271753,I690244,I271779,I271787,I690247,I690241,I271804,I690253,I271830,I271721,I271852,I690256,I271878,I271886,I271903,I271929,I271745,I271951,I271727,I690259,I271991,I272008,I272016,I272033,I271730,I272064,I690250,I272081,I272107,I272115,I271718,I271736,I272160,I690262,I272177,I271739,I271724,I271733,I271742,I272280,I272306,I272314,I272331,I272357,I272248,I272379,I272405,I272413,I272430,I272456,I272272,I272478,I272254,I272518,I272535,I272543,I272560,I272257,I272591,I272608,I272634,I272642,I272245,I272263,I272687,I272704,I272266,I272251,I272260,I272269,I272807,I741958,I272833,I272841,I741955,I741973,I272858,I741964,I272884,I272775,I272906,I741979,I272932,I272940,I741961,I272957,I272983,I272799,I273005,I272781,I741967,I273045,I273062,I273070,I273087,I272784,I273118,I741982,I273135,I741970,I273161,I273169,I272772,I272790,I273214,I741976,I273231,I272793,I272778,I272787,I272796,I273334,I370942,I273360,I273368,I370954,I370933,I273385,I370957,I273411,I273302,I273433,I370948,I273459,I273467,I370930,I273484,I273510,I273326,I273532,I273308,I370945,I273572,I273589,I273597,I273614,I273311,I273645,I370936,I273662,I370939,I273688,I273696,I273299,I273317,I273741,I370951,I273758,I273320,I273305,I273314,I273323,I273861,I983152,I273887,I273895,I983134,I983158,I273912,I983149,I273938,I273829,I273960,I983155,I273986,I273994,I983143,I274011,I274037,I273853,I274059,I273835,I274099,I274116,I274124,I274141,I273838,I274172,I983140,I983137,I274189,I983146,I274215,I274223,I273826,I273844,I274268,I274285,I273847,I273832,I273841,I273850,I274388,I743896,I274414,I274422,I743893,I743911,I274439,I743902,I274465,I274356,I274487,I743917,I274513,I274521,I743899,I274538,I274564,I274380,I274586,I274362,I743905,I274626,I274643,I274651,I274668,I274365,I274699,I743920,I274716,I743908,I274742,I274750,I274353,I274371,I274795,I743914,I274812,I274374,I274359,I274368,I274377,I274915,I874436,I274941,I274949,I874451,I274966,I874454,I274992,I274883,I275014,I874460,I275040,I275048,I874442,I275065,I275091,I274907,I275113,I274889,I874439,I275153,I275170,I275178,I275195,I274892,I275226,I874445,I275243,I874457,I275269,I275277,I274880,I274898,I275322,I874448,I275339,I274901,I274886,I274895,I274904,I275442,I543390,I275468,I275476,I543381,I543396,I275493,I543402,I275519,I275410,I275541,I543387,I275567,I275575,I275592,I275618,I275434,I275640,I275416,I543384,I275680,I275697,I275705,I275722,I275419,I275753,I543378,I543393,I275770,I275796,I275804,I275407,I275425,I275849,I543399,I275866,I275428,I275413,I275422,I275431,I275969,I622788,I275995,I276003,I622791,I622785,I276020,I622797,I276046,I275937,I276068,I622800,I276094,I276102,I276119,I276145,I275961,I276167,I275943,I622803,I276207,I276224,I276232,I276249,I275946,I276280,I622794,I276297,I276323,I276331,I275934,I275952,I276376,I622806,I276393,I275955,I275940,I275949,I275958,I276496,I877904,I276522,I276530,I877919,I276547,I877922,I276573,I276595,I877928,I276621,I276629,I877910,I276646,I276672,I276694,I877907,I276734,I276751,I276759,I276776,I276807,I877913,I276824,I877925,I276850,I276858,I276903,I877916,I276920,I277023,I403845,I277049,I277057,I403857,I277074,I403842,I277100,I276991,I277122,I403866,I277148,I277156,I403863,I277173,I277199,I277015,I277221,I276997,I403854,I277261,I277278,I277286,I277303,I277000,I277334,I403851,I277351,I403860,I277377,I277385,I276988,I277006,I277430,I403848,I277447,I277009,I276994,I277003,I277012,I277550,I680231,I277576,I277584,I680234,I680228,I277601,I680240,I277627,I277518,I277649,I680243,I277675,I277683,I277700,I277726,I277542,I277748,I277524,I680246,I277788,I277805,I277813,I277830,I277527,I277861,I680237,I277878,I277904,I277912,I277515,I277533,I277957,I680249,I277974,I277536,I277521,I277530,I277539,I278077,I352990,I278103,I278111,I353002,I352981,I278128,I353005,I278154,I278045,I278176,I352996,I278202,I278210,I352978,I278227,I278253,I278069,I278275,I278051,I352993,I278315,I278332,I278340,I278357,I278054,I278388,I352984,I278405,I352987,I278431,I278439,I278042,I278060,I278484,I352999,I278501,I278063,I278048,I278057,I278066,I278604,I958128,I278630,I278638,I958110,I958134,I278655,I958125,I278681,I278572,I278703,I958131,I278729,I278737,I958119,I278754,I278780,I278596,I278802,I278578,I278842,I278859,I278867,I278884,I278581,I278915,I958116,I958113,I278932,I958122,I278958,I278966,I278569,I278587,I279011,I279028,I278590,I278575,I278584,I278593,I279131,I279157,I279165,I279182,I279208,I279099,I279230,I279256,I279264,I279281,I279307,I279123,I279329,I279105,I279369,I279386,I279394,I279411,I279108,I279442,I279459,I279485,I279493,I279096,I279114,I279538,I279555,I279117,I279102,I279111,I279120,I279658,I279684,I279692,I279709,I279735,I279626,I279757,I279783,I279791,I279808,I279834,I279650,I279856,I279632,I279896,I279913,I279921,I279938,I279635,I279969,I279986,I280012,I280020,I279623,I279641,I280065,I280082,I279644,I279629,I279638,I279647,I280185,I280211,I280219,I280236,I280262,I280153,I280284,I280310,I280318,I280335,I280361,I280177,I280383,I280159,I280423,I280440,I280448,I280465,I280162,I280496,I280513,I280539,I280547,I280150,I280168,I280592,I280609,I280171,I280156,I280165,I280174,I280712,I668637,I280738,I280746,I668640,I668634,I280763,I668646,I280789,I280811,I668649,I280837,I280845,I280862,I280888,I280910,I668652,I280950,I280967,I280975,I280992,I281023,I668643,I281040,I281066,I281074,I281119,I668655,I281136,I281239,I823150,I281265,I281273,I823147,I281290,I823159,I281316,I281338,I281364,I281372,I823165,I281389,I281415,I281437,I823153,I281477,I281494,I281502,I281519,I281550,I823162,I823168,I281567,I281593,I281601,I281646,I823156,I281663,I281766,I961936,I281792,I281800,I961918,I961942,I281817,I961933,I281843,I281734,I281865,I961939,I281891,I281899,I961927,I281916,I281942,I281758,I281964,I281740,I282004,I282021,I282029,I282046,I281743,I282077,I961924,I961921,I282094,I961930,I282120,I282128,I281731,I281749,I282173,I282190,I281752,I281737,I281746,I281755,I282293,I282319,I282327,I282344,I282370,I282261,I282392,I282418,I282426,I282443,I282469,I282285,I282491,I282267,I282531,I282548,I282556,I282573,I282270,I282604,I282621,I282647,I282655,I282258,I282276,I282700,I282717,I282279,I282264,I282273,I282282,I282820,I753586,I282846,I282854,I753583,I753601,I282871,I753592,I282897,I282788,I282919,I753607,I282945,I282953,I753589,I282970,I282996,I282812,I283018,I282794,I753595,I283058,I283075,I283083,I283100,I282797,I283131,I753610,I283148,I753598,I283174,I283182,I282785,I282803,I283227,I753604,I283244,I282806,I282791,I282800,I282809,I283347,I824272,I283373,I283381,I824269,I283398,I824281,I283424,I283315,I283446,I283472,I283480,I824287,I283497,I283523,I283339,I283545,I283321,I824275,I283585,I283602,I283610,I283627,I283324,I283658,I824284,I824290,I283675,I283701,I283709,I283312,I283330,I283754,I824278,I283771,I283333,I283318,I283327,I283336,I283874,I1013443,I283900,I283908,I1013440,I1013431,I283925,I1013428,I283951,I283973,I1013437,I283999,I284007,I1013446,I284024,I284050,I284072,I1013449,I284112,I284129,I284137,I284154,I284185,I1013434,I284202,I1013452,I284228,I284236,I284281,I284298,I284401,I575180,I284427,I284435,I575171,I575186,I284452,I575192,I284478,I284369,I284500,I575177,I284526,I284534,I284551,I284577,I284393,I284599,I284375,I575174,I284639,I284656,I284664,I284681,I284378,I284712,I575168,I575183,I284729,I284755,I284763,I284366,I284384,I284808,I575189,I284825,I284387,I284372,I284381,I284390,I284928,I284954,I284962,I284979,I285005,I285027,I285053,I285061,I285078,I285104,I285126,I285166,I285183,I285191,I285208,I285239,I285256,I285282,I285290,I285335,I285352,I285455,I831086,I285481,I285489,I831101,I285506,I831104,I285532,I285423,I285554,I831110,I285580,I285588,I831092,I285605,I285631,I285447,I285653,I285429,I831089,I285693,I285710,I285718,I285735,I285432,I285766,I831095,I285783,I831107,I285809,I285817,I285420,I285438,I285862,I831098,I285879,I285441,I285426,I285435,I285444,I285982,I286008,I286016,I286033,I286059,I286081,I286107,I286115,I286132,I286158,I286180,I286220,I286237,I286245,I286262,I286293,I286310,I286336,I286344,I286389,I286406,I286509,I713534,I286535,I286543,I713531,I713549,I286560,I713540,I286586,I286608,I713555,I286634,I286642,I713537,I286659,I286685,I286707,I713543,I286747,I286764,I286772,I286789,I286820,I713558,I286837,I713546,I286863,I286871,I286916,I713552,I286933,I287036,I679177,I287062,I287070,I679180,I679174,I287087,I679186,I287113,I287135,I679189,I287161,I287169,I287186,I287212,I287234,I679192,I287274,I287291,I287299,I287316,I287347,I679183,I287364,I287390,I287398,I287443,I679195,I287460,I287563,I287589,I287597,I287614,I287640,I287531,I287662,I287688,I287696,I287713,I287739,I287555,I287761,I287537,I287801,I287818,I287826,I287843,I287540,I287874,I287891,I287917,I287925,I287528,I287546,I287970,I287987,I287549,I287534,I287543,I287552,I288090,I861720,I288116,I288124,I861735,I288141,I861738,I288167,I288058,I288189,I861744,I288215,I288223,I861726,I288240,I288266,I288082,I288288,I288064,I861723,I288328,I288345,I288353,I288370,I288067,I288401,I861729,I288418,I861741,I288444,I288452,I288055,I288073,I288497,I861732,I288514,I288076,I288061,I288070,I288079,I288617,I899868,I288643,I288651,I899883,I288668,I899886,I288694,I288585,I288716,I899892,I288742,I288750,I899874,I288767,I288793,I288609,I288815,I288591,I899871,I288855,I288872,I288880,I288897,I288594,I288928,I899877,I288945,I899889,I288971,I288979,I288582,I288600,I289024,I899880,I289041,I288603,I288588,I288597,I288606,I289144,I851894,I289170,I289178,I851909,I289195,I851912,I289221,I289112,I289243,I851918,I289269,I289277,I851900,I289294,I289320,I289136,I289342,I289118,I851897,I289382,I289399,I289407,I289424,I289121,I289455,I851903,I289472,I851915,I289498,I289506,I289109,I289127,I289551,I851906,I289568,I289130,I289115,I289124,I289133,I289671,I955356,I289697,I289705,I955371,I289722,I955374,I289748,I289770,I955380,I289796,I289804,I955362,I289821,I289847,I289869,I955359,I289909,I289926,I289934,I289951,I289982,I955365,I289999,I955377,I290025,I290033,I290078,I955368,I290095,I290198,I456693,I290224,I290232,I456678,I456681,I290249,I456696,I290275,I290166,I290297,I456690,I290323,I290331,I290348,I290374,I290190,I290396,I290172,I456687,I290436,I290453,I290461,I290478,I290175,I290509,I456702,I290526,I456699,I290552,I290560,I290163,I290181,I290605,I456684,I290622,I290184,I290169,I290178,I290187,I290725,I290751,I290759,I290776,I290802,I290693,I290824,I290850,I290858,I290875,I290901,I290717,I290923,I290699,I290963,I290980,I290988,I291005,I290702,I291036,I291053,I291079,I291087,I290690,I290708,I291132,I291149,I290711,I290696,I290705,I290714,I291252,I291278,I291286,I291303,I291329,I291220,I291351,I291377,I291385,I291402,I291428,I291244,I291450,I291226,I291490,I291507,I291515,I291532,I291229,I291563,I291580,I291606,I291614,I291217,I291235,I291659,I291676,I291238,I291223,I291232,I291241,I291779,I914896,I291805,I291813,I914911,I291830,I914914,I291856,I291747,I291878,I914920,I291904,I291912,I914902,I291929,I291955,I291771,I291977,I291753,I914899,I292017,I292034,I292042,I292059,I291756,I292090,I914905,I292107,I914917,I292133,I292141,I291744,I291762,I292186,I914908,I292203,I291765,I291750,I291759,I291768,I292306,I410985,I292332,I292340,I410997,I292357,I410982,I292383,I292274,I292405,I411006,I292431,I292439,I411003,I292456,I292482,I292298,I292504,I292280,I410994,I292544,I292561,I292569,I292586,I292283,I292617,I410991,I292634,I411000,I292660,I292668,I292271,I292289,I292713,I410988,I292730,I292292,I292277,I292286,I292295,I292833,I292859,I292867,I292884,I292910,I292932,I292958,I292966,I292983,I293009,I293031,I293071,I293088,I293096,I293113,I293144,I293161,I293187,I293195,I293240,I293257,I293360,I986416,I293386,I293394,I986398,I986422,I293411,I986413,I293437,I293459,I986419,I293485,I293493,I986407,I293510,I293536,I293558,I293598,I293615,I293623,I293640,I293671,I986404,I986401,I293688,I986410,I293714,I293722,I293767,I293784,I293887,I701260,I293913,I293921,I701257,I701275,I293938,I701266,I293964,I293986,I701281,I294012,I294020,I701263,I294037,I294063,I294085,I701269,I294125,I294142,I294150,I294167,I294198,I701284,I294215,I701272,I294241,I294249,I294294,I701278,I294311,I294414,I872124,I294440,I294448,I872139,I294465,I872142,I294491,I294382,I294513,I872148,I294539,I294547,I872130,I294564,I294590,I294406,I294612,I294388,I872127,I294652,I294669,I294677,I294694,I294391,I294725,I872133,I294742,I872145,I294768,I294776,I294379,I294397,I294821,I872136,I294838,I294400,I294385,I294394,I294403,I294941,I554950,I294967,I294975,I554941,I554956,I294992,I554962,I295018,I295040,I554947,I295066,I295074,I295091,I295117,I295139,I554944,I295179,I295196,I295204,I295221,I295252,I554938,I554953,I295269,I295295,I295303,I295348,I554959,I295365,I295468,I594254,I295494,I295502,I594245,I594260,I295519,I594266,I295545,I295436,I295567,I594251,I295593,I295601,I295618,I295644,I295460,I295666,I295442,I594248,I295706,I295723,I295731,I295748,I295445,I295779,I594242,I594257,I295796,I295822,I295830,I295433,I295451,I295875,I594263,I295892,I295454,I295439,I295448,I295457,I295995,I752940,I296021,I296029,I752937,I752955,I296046,I752946,I296072,I295963,I296094,I752961,I296120,I296128,I752943,I296145,I296171,I295987,I296193,I295969,I752949,I296233,I296250,I296258,I296275,I295972,I296306,I752964,I296323,I752952,I296349,I296357,I295960,I295978,I296402,I752958,I296419,I295981,I295966,I295975,I295984,I296522,I408605,I296548,I296556,I408617,I296573,I408602,I296599,I296490,I296621,I408626,I296647,I296655,I408623,I296672,I296698,I296514,I296720,I296496,I408614,I296760,I296777,I296785,I296802,I296499,I296833,I408611,I296850,I408620,I296876,I296884,I296487,I296505,I296929,I408608,I296946,I296508,I296493,I296502,I296511,I297049,I905648,I297075,I297083,I905663,I297100,I905666,I297126,I297017,I297148,I905672,I297174,I297182,I905654,I297199,I297225,I297041,I297247,I297023,I905651,I297287,I297304,I297312,I297329,I297026,I297360,I905657,I297377,I905669,I297403,I297411,I297014,I297032,I297456,I905660,I297473,I297035,I297020,I297029,I297038,I297576,I711596,I297602,I297610,I711593,I711611,I297627,I711602,I297653,I297544,I297675,I711617,I297701,I297709,I711599,I297726,I297752,I297568,I297774,I297550,I711605,I297814,I297831,I297839,I297856,I297553,I297887,I711620,I297904,I711608,I297930,I297938,I297541,I297559,I297983,I711614,I298000,I297562,I297547,I297556,I297565,I298103,I991479,I298129,I298137,I991476,I991467,I298154,I991464,I298180,I298202,I991473,I298228,I298236,I991482,I298253,I298279,I298301,I991485,I298341,I298358,I298366,I298383,I298414,I991470,I298431,I991488,I298457,I298465,I298510,I298527,I298630,I840334,I298656,I298664,I840349,I298681,I840352,I298707,I298598,I298729,I840358,I298755,I298763,I840340,I298780,I298806,I298622,I298828,I298604,I840337,I298868,I298885,I298893,I298910,I298607,I298941,I840343,I298958,I840355,I298984,I298992,I298595,I298613,I299037,I840346,I299054,I298616,I298601,I298610,I298619,I299157,I299183,I299191,I299208,I299234,I299125,I299256,I299282,I299290,I299307,I299333,I299149,I299355,I299131,I299395,I299412,I299420,I299437,I299134,I299468,I299485,I299511,I299519,I299122,I299140,I299564,I299581,I299143,I299128,I299137,I299146,I299684,I959760,I299710,I299718,I959742,I959766,I299735,I959757,I299761,I299652,I299783,I959763,I299809,I299817,I959751,I299834,I299860,I299676,I299882,I299658,I299922,I299939,I299947,I299964,I299661,I299995,I959748,I959745,I300012,I959754,I300038,I300046,I299649,I299667,I300091,I300108,I299670,I299655,I299664,I299673,I300211,I300237,I300245,I300262,I300288,I300179,I300310,I300336,I300344,I300361,I300387,I300203,I300409,I300185,I300449,I300466,I300474,I300491,I300188,I300522,I300539,I300565,I300573,I300176,I300194,I300618,I300635,I300197,I300182,I300191,I300200,I300738,I300764,I300772,I300789,I300815,I300837,I300863,I300871,I300888,I300914,I300936,I300976,I300993,I301001,I301018,I301049,I301066,I301092,I301100,I301145,I301162,I301265,I693933,I301291,I301299,I693936,I693930,I301316,I693942,I301342,I301233,I301364,I693945,I301390,I301398,I301415,I301441,I301257,I301463,I301239,I693948,I301503,I301520,I301528,I301545,I301242,I301576,I693939,I301593,I301619,I301627,I301230,I301248,I301672,I693951,I301689,I301251,I301236,I301245,I301254,I301792,I1095950,I301818,I301826,I1095929,I301843,I1095956,I301869,I301760,I301891,I1095944,I301917,I301925,I1095947,I301942,I301968,I301784,I301990,I301766,I1095938,I302030,I302047,I302055,I302072,I301769,I302103,I1095935,I1095932,I302120,I1095953,I302146,I302154,I301757,I301775,I302199,I1095941,I302216,I301778,I301763,I301772,I301781,I302319,I811930,I302345,I302353,I811927,I302370,I811939,I302396,I302287,I302418,I302444,I302452,I811945,I302469,I302495,I302311,I302517,I302293,I811933,I302557,I302574,I302582,I302599,I302296,I302630,I811942,I811948,I302647,I302673,I302681,I302284,I302302,I302726,I811936,I302743,I302305,I302290,I302299,I302308,I302846,I448023,I302872,I302880,I448008,I448011,I302897,I448026,I302923,I302814,I302945,I448020,I302971,I302979,I302996,I303022,I302838,I303044,I302820,I448017,I303084,I303101,I303109,I303126,I302823,I303157,I448032,I303174,I448029,I303200,I303208,I302811,I302829,I303253,I448014,I303270,I302832,I302817,I302826,I302835,I303373,I492529,I303399,I303407,I492514,I492517,I303424,I492532,I303450,I303341,I303472,I492526,I303498,I303506,I303523,I303549,I303365,I303571,I303347,I492523,I303611,I303628,I303636,I303653,I303350,I303684,I492538,I303701,I492535,I303727,I303735,I303338,I303356,I303780,I492520,I303797,I303359,I303344,I303353,I303362,I303900,I825394,I303926,I303934,I825391,I303951,I825403,I303977,I303868,I303999,I304025,I304033,I825409,I304050,I304076,I303892,I304098,I303874,I825397,I304138,I304155,I304163,I304180,I303877,I304211,I825406,I825412,I304228,I304254,I304262,I303865,I303883,I304307,I825400,I304324,I303886,I303871,I303880,I303889,I304427,I813613,I304453,I304461,I813610,I304478,I813622,I304504,I304395,I304526,I304552,I304560,I813628,I304577,I304603,I304419,I304625,I304401,I813616,I304665,I304682,I304690,I304707,I304404,I304738,I813625,I813631,I304755,I304781,I304789,I304392,I304410,I304834,I813619,I304851,I304413,I304398,I304407,I304416,I304954,I1030500,I304980,I304988,I1030479,I305005,I1030506,I305031,I305053,I1030494,I305079,I305087,I1030497,I305104,I305130,I305152,I1030488,I305192,I305209,I305217,I305234,I305265,I1030485,I1030482,I305282,I1030503,I305308,I305316,I305361,I1030491,I305378,I305481,I305507,I305515,I305532,I305558,I305449,I305580,I305606,I305614,I305631,I305657,I305473,I305679,I305455,I305719,I305736,I305744,I305761,I305458,I305792,I305809,I305835,I305843,I305446,I305464,I305888,I305905,I305467,I305452,I305461,I305470,I306008,I650719,I306034,I306042,I650722,I650716,I306059,I650728,I306085,I305976,I306107,I650731,I306133,I306141,I306158,I306184,I306000,I306206,I305982,I650734,I306246,I306263,I306271,I306288,I305985,I306319,I650725,I306336,I306362,I306370,I305973,I305991,I306415,I650737,I306432,I305994,I305979,I305988,I305997,I306535,I1029918,I306561,I306569,I1029945,I1029921,I306586,I1029930,I306612,I306503,I306634,I306660,I306668,I1029942,I306685,I306711,I306527,I306733,I306509,I1029924,I306773,I306790,I306798,I306815,I306512,I306846,I1029939,I1029927,I306863,I1029933,I306889,I306897,I306500,I306518,I306942,I1029936,I306959,I306521,I306506,I306515,I306524,I307062,I661786,I307088,I307096,I661789,I661783,I307113,I661795,I307139,I307030,I307161,I661798,I307187,I307195,I307212,I307238,I307054,I307260,I307036,I661801,I307300,I307317,I307325,I307342,I307039,I307373,I661792,I307390,I307416,I307424,I307027,I307045,I307469,I661804,I307486,I307048,I307033,I307042,I307051,I307589,I307615,I307623,I307640,I307666,I307688,I307714,I307722,I307739,I307765,I307787,I307827,I307844,I307852,I307869,I307900,I307917,I307943,I307951,I307996,I308013,I308116,I723224,I308142,I308150,I723221,I723239,I308167,I723230,I308193,I308084,I308215,I723245,I308241,I308249,I723227,I308266,I308292,I308108,I308314,I308090,I723233,I308354,I308371,I308379,I308396,I308093,I308427,I723248,I308444,I723236,I308470,I308478,I308081,I308099,I308523,I723242,I308540,I308102,I308087,I308096,I308105,I308643,I329054,I308669,I308677,I329066,I329045,I308694,I329069,I308720,I308611,I308742,I329060,I308768,I308776,I329042,I308793,I308819,I308635,I308841,I308617,I329057,I308881,I308898,I308906,I308923,I308620,I308954,I329048,I308971,I329051,I308997,I309005,I308608,I308626,I309050,I329063,I309067,I308629,I308614,I308623,I308632,I309170,I309196,I309204,I309221,I309247,I309138,I309269,I309295,I309303,I309320,I309346,I309162,I309368,I309144,I309408,I309425,I309433,I309450,I309147,I309481,I309498,I309524,I309532,I309135,I309153,I309577,I309594,I309156,I309141,I309150,I309159,I309697,I309723,I309731,I309748,I309774,I309665,I309796,I309822,I309830,I309847,I309873,I309689,I309895,I309671,I309935,I309952,I309960,I309977,I309674,I310008,I310025,I310051,I310059,I309662,I309680,I310104,I310121,I309683,I309668,I309677,I309686,I310224,I489639,I310250,I310258,I489624,I489627,I310275,I489642,I310301,I310192,I310323,I489636,I310349,I310357,I310374,I310400,I310216,I310422,I310198,I489633,I310462,I310479,I310487,I310504,I310201,I310535,I489648,I310552,I489645,I310578,I310586,I310189,I310207,I310631,I489630,I310648,I310210,I310195,I310204,I310213,I310751,I965744,I310777,I310785,I965726,I965750,I310802,I965741,I310828,I310850,I965747,I310876,I310884,I965735,I310901,I310927,I310949,I310989,I311006,I311014,I311031,I311062,I965732,I965729,I311079,I965738,I311105,I311113,I311158,I311175,I311278,I988589,I311304,I311312,I988586,I988577,I311329,I988574,I311355,I311246,I311377,I988583,I311403,I311411,I988592,I311428,I311454,I311270,I311476,I311252,I988595,I311516,I311533,I311541,I311558,I311255,I311589,I988580,I311606,I988598,I311632,I311640,I311243,I311261,I311685,I311702,I311264,I311249,I311258,I311267,I311805,I637544,I311831,I311839,I637547,I637541,I311856,I637553,I311882,I311773,I311904,I637556,I311930,I311938,I311955,I311981,I311797,I312003,I311779,I637559,I312043,I312060,I312068,I312085,I311782,I312116,I637550,I312133,I312159,I312167,I311770,I311788,I312212,I637562,I312229,I311791,I311776,I311785,I311794,I312332,I1096545,I312358,I312366,I1096524,I312383,I1096551,I312409,I312300,I312431,I1096539,I312457,I312465,I1096542,I312482,I312508,I312324,I312530,I312306,I1096533,I312570,I312587,I312595,I312612,I312309,I312643,I1096530,I1096527,I312660,I1096548,I312686,I312694,I312297,I312315,I312739,I1096536,I312756,I312318,I312303,I312312,I312321,I312859,I446867,I312885,I312893,I446852,I446855,I312910,I446870,I312936,I312827,I312958,I446864,I312984,I312992,I313009,I313035,I312851,I313057,I312833,I446861,I313097,I313114,I313122,I313139,I312836,I313170,I446876,I313187,I446873,I313213,I313221,I312824,I312842,I313266,I446858,I313283,I312845,I312830,I312839,I312848,I313386,I313412,I313420,I313437,I313463,I313485,I313511,I313519,I313536,I313562,I313584,I313624,I313641,I313649,I313666,I313697,I313714,I313740,I313748,I313793,I313810,I313913,I1066795,I313939,I313947,I1066774,I313964,I1066801,I313990,I313881,I314012,I1066789,I314038,I314046,I1066792,I314063,I314089,I313905,I314111,I313887,I1066783,I314151,I314168,I314176,I314193,I313890,I314224,I1066780,I1066777,I314241,I1066798,I314267,I314275,I313878,I313896,I314320,I1066786,I314337,I313899,I313884,I313893,I313902,I314440,I473455,I314466,I314474,I473440,I473443,I314491,I473458,I314517,I314408,I314539,I473452,I314565,I314573,I314590,I314616,I314432,I314638,I314414,I473449,I314678,I314695,I314703,I314720,I314417,I314751,I473464,I314768,I473461,I314794,I314802,I314405,I314423,I314847,I473446,I314864,I314426,I314411,I314420,I314429,I314967,I314993,I315001,I315018,I315044,I314935,I315066,I315092,I315100,I315117,I315143,I314959,I315165,I314941,I315205,I315222,I315230,I315247,I314944,I315278,I315295,I315321,I315329,I314932,I314950,I315374,I315391,I314953,I314938,I314947,I314956,I315494,I315520,I315528,I315545,I315571,I315462,I315593,I315619,I315627,I315644,I315670,I315486,I315692,I315468,I315732,I315749,I315757,I315774,I315471,I315805,I315822,I315848,I315856,I315459,I315477,I315901,I315918,I315480,I315465,I315474,I315483,I316021,I395515,I316047,I316064,I316086,I316103,I395518,I395536,I316120,I395524,I316146,I316154,I316180,I316188,I395533,I316205,I395527,I316245,I316253,I316298,I395530,I395512,I316315,I395521,I316341,I316363,I316380,I316397,I316428,I316445,I316476,I316565,I673916,I316591,I316608,I316557,I316630,I316647,I673910,I673907,I316664,I673922,I316690,I316698,I316724,I316732,I673904,I316749,I316536,I316789,I316797,I316530,I316545,I316842,I673919,I673913,I316859,I316885,I316533,I316907,I316924,I316941,I316548,I316972,I316989,I673925,I316539,I317020,I316542,I316554,I316551,I317109,I432983,I317135,I317152,I317101,I317174,I317191,I432980,I433001,I317208,I433004,I317234,I317242,I432989,I317268,I317276,I432992,I317293,I317080,I432995,I317333,I317341,I317074,I317089,I317386,I432986,I317403,I432998,I317429,I317077,I317451,I317468,I317485,I317092,I317516,I317533,I317083,I317564,I317086,I317098,I317095,I317653,I981505,I317679,I317696,I317645,I317718,I317735,I981517,I981520,I317752,I981523,I317778,I317786,I981508,I317812,I317820,I981514,I317837,I317624,I981502,I317877,I317885,I317618,I317633,I317930,I981526,I317947,I981511,I317973,I317621,I317995,I318012,I318029,I317636,I318060,I318077,I317627,I318108,I317630,I317642,I317639,I318197,I998418,I318223,I318240,I318189,I318262,I318279,I998415,I998412,I318296,I998400,I318322,I318330,I998424,I318356,I318364,I998409,I318381,I318168,I998403,I318421,I318429,I318162,I318177,I318474,I998406,I318491,I998421,I318517,I318165,I318539,I318556,I318573,I318180,I318604,I318621,I318171,I318652,I318174,I318186,I318183,I318741,I318767,I318784,I318733,I318806,I318823,I318840,I318866,I318874,I318900,I318908,I318925,I318712,I318965,I318973,I318706,I318721,I319018,I319035,I319061,I318709,I319083,I319100,I319117,I318724,I319148,I319165,I318715,I319196,I318718,I318730,I318727,I319285,I709661,I319311,I319328,I319277,I319350,I319367,I709676,I709664,I319384,I709655,I319410,I319418,I709667,I319444,I319452,I709658,I319469,I319256,I709673,I319509,I319517,I319250,I319265,I319562,I709682,I709670,I319579,I709679,I319605,I319253,I319627,I319644,I319661,I319268,I319692,I319709,I319259,I319740,I319262,I319274,I319271,I319829,I394325,I319855,I319872,I319894,I319911,I394328,I394346,I319928,I394334,I319954,I319962,I319988,I319996,I394343,I320013,I394337,I320053,I320061,I320106,I394340,I394322,I320123,I394331,I320149,I320171,I320188,I320205,I320236,I320253,I320284,I320373,I320399,I320416,I320365,I320438,I320455,I320472,I320498,I320506,I320532,I320540,I320557,I320344,I320597,I320605,I320338,I320353,I320650,I320667,I320693,I320341,I320715,I320732,I320749,I320356,I320780,I320797,I320347,I320828,I320350,I320362,I320359,I320917,I724519,I320943,I320960,I320982,I320999,I724534,I724522,I321016,I724513,I321042,I321050,I724525,I321076,I321084,I724516,I321101,I724531,I321141,I321149,I321194,I724540,I724528,I321211,I724537,I321237,I321259,I321276,I321293,I321324,I321341,I321372,I321461,I843227,I321487,I321504,I321526,I321543,I843239,I321560,I843230,I321586,I321594,I843248,I321620,I321628,I843224,I321645,I843242,I321685,I321693,I321738,I843236,I843233,I321755,I843245,I321781,I321803,I321820,I321837,I321868,I321885,I321916,I322005,I322031,I322048,I321997,I322070,I322087,I322104,I322130,I322138,I322164,I322172,I322189,I321976,I322229,I322237,I321970,I321985,I322282,I322299,I322325,I321973,I322347,I322364,I322381,I321988,I322412,I322429,I321979,I322460,I321982,I321994,I321991,I322549,I892935,I322575,I322592,I322541,I322614,I322631,I892947,I322648,I892938,I322674,I322682,I892956,I322708,I322716,I892932,I322733,I322520,I892950,I322773,I322781,I322514,I322529,I322826,I892944,I892941,I322843,I892953,I322869,I322517,I322891,I322908,I322925,I322532,I322956,I322973,I322523,I323004,I322526,I322538,I322535,I323093,I714829,I323119,I323136,I323085,I323158,I323175,I714844,I714832,I323192,I714823,I323218,I323226,I714835,I323252,I323260,I714826,I323277,I323064,I714841,I323317,I323325,I323058,I323073,I323370,I714850,I714838,I323387,I714847,I323413,I323061,I323435,I323452,I323469,I323076,I323500,I323517,I323067,I323548,I323070,I323082,I323079,I323637,I964641,I323663,I323680,I323629,I323702,I323719,I964653,I964656,I323736,I964659,I323762,I323770,I964644,I323796,I323804,I964650,I323821,I323608,I964638,I323861,I323869,I323602,I323617,I323914,I964662,I323931,I964647,I323957,I323605,I323979,I323996,I324013,I323620,I324044,I324061,I323611,I324092,I323614,I323626,I323623,I324181,I1003042,I324207,I324224,I324173,I324246,I324263,I1003039,I1003036,I324280,I1003024,I324306,I324314,I1003048,I324340,I324348,I1003033,I324365,I324152,I1003027,I324405,I324413,I324146,I324161,I324458,I1003030,I324475,I1003045,I324501,I324149,I324523,I324540,I324557,I324164,I324588,I324605,I324155,I324636,I324158,I324170,I324167,I324725,I324751,I324768,I324717,I324790,I324807,I324824,I324850,I324858,I324884,I324892,I324909,I324696,I324949,I324957,I324690,I324705,I325002,I325019,I325045,I324693,I325067,I325084,I325101,I324708,I325132,I325149,I324699,I325180,I324702,I324714,I324711,I325269,I739377,I325295,I325312,I325334,I325351,I739392,I739380,I325368,I739371,I325394,I325402,I739383,I325428,I325436,I739374,I325453,I739389,I325493,I325501,I325546,I739398,I739386,I325563,I739395,I325589,I325611,I325628,I325645,I325676,I325693,I325724,I325813,I718705,I325839,I325856,I325878,I325895,I718720,I718708,I325912,I718699,I325938,I325946,I718711,I325972,I325980,I718702,I325997,I718717,I326037,I326045,I326090,I718726,I718714,I326107,I718723,I326133,I326155,I326172,I326189,I326220,I326237,I326268,I326357,I1057876,I326383,I326400,I326349,I326422,I326439,I1057852,I1057873,I326456,I1057870,I326482,I326490,I1057849,I326516,I326524,I1057861,I326541,I326328,I1057864,I326581,I326589,I326322,I326337,I326634,I1057867,I1057855,I326651,I1057858,I326677,I326325,I326699,I326716,I326733,I326340,I326764,I326781,I326331,I326812,I326334,I326346,I326343,I326901,I772969,I326927,I326944,I326966,I326983,I772984,I772972,I327000,I772963,I327026,I327034,I772975,I327060,I327068,I772966,I327085,I772981,I327125,I327133,I327178,I772990,I772978,I327195,I772987,I327221,I327243,I327260,I327277,I327308,I327325,I327356,I327445,I435873,I327471,I327488,I327437,I327510,I327527,I435870,I435891,I327544,I435894,I327570,I327578,I435879,I327604,I327612,I435882,I327629,I327416,I435885,I327669,I327677,I327410,I327425,I327722,I435876,I327739,I435888,I327765,I327413,I327787,I327804,I327821,I327428,I327852,I327869,I327419,I327900,I327422,I327434,I327431,I327989,I1033481,I328015,I328032,I327981,I328054,I328071,I1033457,I1033478,I328088,I1033475,I328114,I328122,I1033454,I328148,I328156,I1033466,I328173,I327960,I1033469,I328213,I328221,I327954,I327969,I328266,I1033472,I1033460,I328283,I1033463,I328309,I327957,I328331,I328348,I328365,I327972,I328396,I328413,I327963,I328444,I327966,I327978,I327975,I328533,I328559,I328576,I328525,I328598,I328615,I328632,I328658,I328666,I328692,I328700,I328717,I328504,I328757,I328765,I328498,I328513,I328810,I328827,I328853,I328501,I328875,I328892,I328909,I328516,I328940,I328957,I328507,I328988,I328510,I328522,I328519,I329077,I1098931,I329103,I329120,I329142,I329159,I1098907,I1098928,I329176,I1098925,I329202,I329210,I1098904,I329236,I329244,I1098916,I329261,I1098919,I329301,I329309,I329354,I1098922,I1098910,I329371,I1098913,I329397,I329419,I329436,I329453,I329484,I329501,I329532,I329621,I669700,I329647,I329664,I329613,I329686,I329703,I669694,I669691,I329720,I669706,I329746,I329754,I329780,I329788,I669688,I329805,I329592,I329845,I329853,I329586,I329601,I329898,I669703,I669697,I329915,I329941,I329589,I329963,I329980,I329997,I329604,I330028,I330045,I669709,I329595,I330076,I329598,I329610,I329607,I330165,I876173,I330191,I330208,I330230,I330247,I876185,I330264,I876176,I330290,I330298,I876194,I330324,I330332,I876170,I330349,I876188,I330389,I330397,I330442,I876182,I876179,I330459,I876191,I330485,I330507,I330524,I330541,I330572,I330589,I330620,I330709,I330735,I330752,I330701,I330774,I330791,I330808,I330834,I330842,I330868,I330876,I330893,I330680,I330933,I330941,I330674,I330689,I330986,I331003,I331029,I330677,I331051,I331068,I331085,I330692,I331116,I331133,I330683,I331164,I330686,I330698,I330695,I331253,I825952,I331279,I331296,I331245,I331318,I331335,I825970,I331352,I825964,I331378,I331386,I825958,I331412,I331420,I825967,I331437,I331224,I825955,I331477,I331485,I331218,I331233,I331530,I825973,I331547,I331573,I331221,I331595,I331612,I331629,I331236,I331660,I331677,I825961,I331227,I331708,I331230,I331242,I331239,I331797,I331823,I331840,I331789,I331862,I331879,I331896,I331922,I331930,I331956,I331964,I331981,I331768,I332021,I332029,I331762,I331777,I332074,I332091,I332117,I331765,I332139,I332156,I332173,I331780,I332204,I332221,I331771,I332252,I331774,I331786,I331783,I332341,I332367,I332384,I332333,I332406,I332423,I332440,I332466,I332474,I332500,I332508,I332525,I332312,I332565,I332573,I332306,I332321,I332618,I332635,I332661,I332309,I332683,I332700,I332717,I332324,I332748,I332765,I332315,I332796,I332318,I332330,I332327,I332885,I332911,I332928,I332877,I332950,I332967,I332984,I333010,I333018,I333044,I333052,I333069,I332856,I333109,I333117,I332850,I332865,I333162,I333179,I333205,I332853,I333227,I333244,I333261,I332868,I333292,I333309,I332859,I333340,I332862,I332874,I332871,I333429,I727103,I333455,I333472,I333494,I333511,I727118,I727106,I333528,I727097,I333554,I333562,I727109,I333588,I333596,I727100,I333613,I727115,I333653,I333661,I333706,I727124,I727112,I333723,I727121,I333749,I333771,I333788,I333805,I333836,I333853,I333884,I333973,I894091,I333999,I334016,I333965,I334038,I334055,I894103,I334072,I894094,I334098,I334106,I894112,I334132,I334140,I894088,I334157,I333944,I894106,I334197,I334205,I333938,I333953,I334250,I894100,I894097,I334267,I894109,I334293,I333941,I334315,I334332,I334349,I333956,I334380,I334397,I333947,I334428,I333950,I333962,I333959,I334517,I1097146,I334543,I334560,I334509,I334582,I334599,I1097122,I1097143,I334616,I1097140,I334642,I334650,I1097119,I334676,I334684,I1097131,I334701,I334488,I1097134,I334741,I334749,I334482,I334497,I334794,I1097137,I1097125,I334811,I1097128,I334837,I334485,I334859,I334876,I334893,I334500,I334924,I334941,I334491,I334972,I334494,I334506,I334503,I335061,I335087,I335104,I335053,I335126,I335143,I335160,I335186,I335194,I335220,I335228,I335245,I335032,I335285,I335293,I335026,I335041,I335338,I335355,I335381,I335029,I335403,I335420,I335437,I335044,I335468,I335485,I335035,I335516,I335038,I335050,I335047,I335605,I579795,I335631,I335648,I335670,I335687,I579816,I579807,I335704,I335730,I335738,I579801,I335764,I335772,I579798,I335789,I579792,I335829,I335837,I335882,I579804,I335899,I579813,I335925,I335947,I335964,I335981,I336012,I336029,I579810,I336060,I336149,I336175,I336192,I336141,I336214,I336231,I336248,I336274,I336282,I336308,I336316,I336333,I336120,I336373,I336381,I336114,I336129,I336426,I336443,I336469,I336117,I336491,I336508,I336525,I336132,I336556,I336573,I336123,I336604,I336126,I336138,I336135,I336693,I1032291,I336719,I336736,I336758,I336775,I1032267,I1032288,I336792,I1032285,I336818,I336826,I1032264,I336852,I336860,I1032276,I336877,I1032279,I336917,I336925,I336970,I1032282,I1032270,I336987,I1032273,I337013,I337035,I337052,I337069,I337100,I337117,I337148,I337237,I1060851,I337263,I337280,I337229,I337302,I337319,I1060827,I1060848,I337336,I1060845,I337362,I337370,I1060824,I337396,I337404,I1060836,I337421,I337208,I1060839,I337461,I337469,I337202,I337217,I337514,I1060842,I1060830,I337531,I1060833,I337557,I337205,I337579,I337596,I337613,I337220,I337644,I337661,I337211,I337692,I337214,I337226,I337223,I337781,I583841,I337807,I337824,I337773,I337846,I337863,I583862,I583853,I337880,I337906,I337914,I583847,I337940,I337948,I583844,I337965,I337752,I583838,I338005,I338013,I337746,I337761,I338058,I583850,I338075,I583859,I338101,I337749,I338123,I338140,I338157,I337764,I338188,I338205,I583856,I337755,I338236,I337758,I337770,I337767,I338325,I1054306,I338351,I338368,I338317,I338390,I338407,I1054282,I1054303,I338424,I1054300,I338450,I338458,I1054279,I338484,I338492,I1054291,I338509,I338296,I1054294,I338549,I338557,I338290,I338305,I338602,I1054297,I1054285,I338619,I1054288,I338645,I338293,I338667,I338684,I338701,I338308,I338732,I338749,I338299,I338780,I338302,I338314,I338311,I338869,I338895,I338912,I338861,I338934,I338951,I338968,I338994,I339002,I339028,I339036,I339053,I338840,I339093,I339101,I338834,I338849,I339146,I339163,I339189,I338837,I339211,I339228,I339245,I338852,I339276,I339293,I338843,I339324,I338846,I338858,I338855,I339413,I1009400,I339439,I339456,I339478,I339495,I1009397,I1009394,I339512,I1009382,I339538,I339546,I1009406,I339572,I339580,I1009391,I339597,I1009385,I339637,I339645,I339690,I1009388,I339707,I1009403,I339733,I339755,I339772,I339789,I339820,I339837,I339868,I339957,I1081676,I339983,I340000,I339949,I340022,I340039,I1081652,I1081673,I340056,I1081670,I340082,I340090,I1081649,I340116,I340124,I1081661,I340141,I339928,I1081664,I340181,I340189,I339922,I339937,I340234,I1081667,I1081655,I340251,I1081658,I340277,I339925,I340299,I340316,I340333,I339940,I340364,I340381,I339931,I340412,I339934,I339946,I339943,I340501,I340527,I340544,I340493,I340566,I340583,I340600,I340626,I340634,I340660,I340668,I340685,I340472,I340725,I340733,I340466,I340481,I340778,I340795,I340821,I340469,I340843,I340860,I340877,I340484,I340908,I340925,I340475,I340956,I340478,I340490,I340487,I341045,I669173,I341071,I341088,I341037,I341110,I341127,I669167,I669164,I341144,I669179,I341170,I341178,I341204,I341212,I669161,I341229,I341016,I341269,I341277,I341010,I341025,I341322,I669176,I669170,I341339,I341365,I341013,I341387,I341404,I341421,I341028,I341452,I341469,I669182,I341019,I341500,I341022,I341034,I341031,I341589,I341615,I341632,I341581,I341654,I341671,I341688,I341714,I341722,I341748,I341756,I341773,I341560,I341813,I341821,I341554,I341569,I341866,I341883,I341909,I341557,I341931,I341948,I341965,I341572,I341996,I342013,I341563,I342044,I341566,I341578,I341575,I342133,I342159,I342176,I342198,I342215,I342232,I342258,I342266,I342292,I342300,I342317,I342357,I342365,I342410,I342427,I342453,I342475,I342492,I342509,I342540,I342557,I342588,I342677,I459571,I342703,I342720,I342669,I342742,I342759,I459568,I459589,I342776,I459592,I342802,I342810,I459577,I342836,I342844,I459580,I342861,I342648,I459583,I342901,I342909,I342642,I342657,I342954,I459574,I342971,I459586,I342997,I342645,I343019,I343036,I343053,I342660,I343084,I343101,I342651,I343132,I342654,I342666,I342663,I343221,I343247,I343264,I343213,I343286,I343303,I343320,I343346,I343354,I343380,I343388,I343405,I343192,I343445,I343453,I343186,I343201,I343498,I343515,I343541,I343189,I343563,I343580,I343597,I343204,I343628,I343645,I343195,I343676,I343198,I343210,I343207,I343765,I584997,I343791,I343808,I343757,I343830,I343847,I585018,I585009,I343864,I343890,I343898,I585003,I343924,I343932,I585000,I343949,I343736,I584994,I343989,I343997,I343730,I343745,I344042,I585006,I344059,I585015,I344085,I343733,I344107,I344124,I344141,I343748,I344172,I344189,I585012,I343739,I344220,I343742,I343754,I343751,I344309,I906229,I344335,I344352,I344301,I344374,I344391,I906241,I344408,I906232,I344434,I344442,I906250,I344468,I344476,I906226,I344493,I344280,I906244,I344533,I344541,I344274,I344289,I344586,I906238,I906235,I344603,I906247,I344629,I344277,I344651,I344668,I344685,I344292,I344716,I344733,I344283,I344764,I344286,I344298,I344295,I344853,I344879,I344896,I344845,I344918,I344935,I344952,I344978,I344986,I345012,I345020,I345037,I344824,I345077,I345085,I344818,I344833,I345130,I345147,I345173,I344821,I345195,I345212,I345229,I344836,I345260,I345277,I344827,I345308,I344830,I344842,I344839,I345397,I345423,I345440,I345389,I345462,I345479,I345496,I345522,I345530,I345556,I345564,I345581,I345368,I345621,I345629,I345362,I345377,I345674,I345691,I345717,I345365,I345739,I345756,I345773,I345380,I345804,I345821,I345371,I345852,I345374,I345386,I345383,I345941,I942643,I345967,I345984,I345933,I346006,I346023,I942655,I346040,I942646,I346066,I346074,I942664,I346100,I346108,I942640,I346125,I345912,I942658,I346165,I346173,I345906,I345921,I346218,I942652,I942649,I346235,I942661,I346261,I345909,I346283,I346300,I346317,I345924,I346348,I346365,I345915,I346396,I345918,I345930,I345927,I346485,I346511,I346528,I346477,I346550,I346567,I346584,I346610,I346618,I346644,I346652,I346669,I346456,I346709,I346717,I346450,I346465,I346762,I346779,I346805,I346453,I346827,I346844,I346861,I346468,I346892,I346909,I346459,I346940,I346462,I346474,I346471,I347029,I557831,I347055,I347072,I347094,I347111,I557852,I557843,I347128,I347154,I347162,I557837,I347188,I347196,I557834,I347213,I557828,I347253,I347261,I347306,I557840,I347323,I557849,I347349,I347371,I347388,I347405,I347436,I347453,I557846,I347484,I347573,I538757,I347599,I347616,I347565,I347638,I347655,I538778,I538769,I347672,I347698,I347706,I538763,I347732,I347740,I538760,I347757,I347544,I538754,I347797,I347805,I347538,I347553,I347850,I538766,I347867,I538775,I347893,I347541,I347915,I347932,I347949,I347556,I347980,I347997,I538772,I347547,I348028,I347550,I347562,I347559,I348117,I766509,I348143,I348160,I348109,I348182,I348199,I766524,I766512,I348216,I766503,I348242,I348250,I766515,I348276,I348284,I766506,I348301,I348088,I766521,I348341,I348349,I348082,I348097,I348394,I766530,I766518,I348411,I766527,I348437,I348085,I348459,I348476,I348493,I348100,I348524,I348541,I348091,I348572,I348094,I348106,I348103,I348661,I655998,I348687,I348704,I348726,I348743,I655992,I655989,I348760,I656004,I348786,I348794,I348820,I348828,I655986,I348845,I348885,I348893,I348938,I656001,I655995,I348955,I348981,I349003,I349020,I349037,I349068,I349085,I656007,I349116,I349205,I349231,I349248,I349197,I349270,I349287,I349304,I349330,I349338,I349364,I349372,I349389,I349176,I349429,I349437,I349170,I349185,I349482,I349499,I349525,I349173,I349547,I349564,I349581,I349188,I349612,I349629,I349179,I349660,I349182,I349194,I349191,I349749,I779429,I349775,I349792,I349741,I349814,I349831,I779444,I779432,I349848,I779423,I349874,I349882,I779435,I349908,I349916,I779426,I349933,I349720,I779441,I349973,I349981,I349714,I349729,I350026,I779450,I779438,I350043,I779447,I350069,I349717,I350091,I350108,I350125,I349732,I350156,I350173,I349723,I350204,I349726,I349738,I349735,I350293,I350319,I350336,I350358,I350375,I350392,I350418,I350426,I350452,I350460,I350477,I350517,I350525,I350570,I350587,I350613,I350635,I350652,I350669,I350700,I350717,I350748,I350837,I350863,I350880,I350829,I350902,I350919,I350936,I350962,I350970,I350996,I351004,I351021,I350808,I351061,I351069,I350802,I350817,I351114,I351131,I351157,I350805,I351179,I351196,I351213,I350820,I351244,I351261,I350811,I351292,I350814,I350826,I350823,I351381,I351407,I351424,I351373,I351446,I351463,I351480,I351506,I351514,I351540,I351548,I351565,I351352,I351605,I351613,I351346,I351361,I351658,I351675,I351701,I351349,I351723,I351740,I351757,I351364,I351788,I351805,I351355,I351836,I351358,I351370,I351367,I351925,I836291,I351951,I351968,I351917,I351990,I352007,I836303,I352024,I836294,I352050,I352058,I836312,I352084,I352092,I836288,I352109,I351896,I836306,I352149,I352157,I351890,I351905,I352202,I836300,I836297,I352219,I836309,I352245,I351893,I352267,I352284,I352301,I351908,I352332,I352349,I351899,I352380,I351902,I351914,I351911,I352469,I625432,I352495,I352512,I352461,I352534,I352551,I625426,I625423,I352568,I625438,I352594,I352602,I352628,I352636,I625420,I352653,I352440,I352693,I352701,I352434,I352449,I352746,I625435,I625429,I352763,I352789,I352437,I352811,I352828,I352845,I352452,I352876,I352893,I625441,I352443,I352924,I352446,I352458,I352455,I353013,I353039,I353056,I353078,I353095,I353112,I353138,I353146,I353172,I353180,I353197,I353237,I353245,I353290,I353307,I353333,I353355,I353372,I353389,I353420,I353437,I353468,I353557,I632810,I353583,I353600,I353549,I353622,I353639,I632804,I632801,I353656,I632816,I353682,I353690,I353716,I353724,I632798,I353741,I353528,I353781,I353789,I353522,I353537,I353834,I632813,I632807,I353851,I353877,I353525,I353899,I353916,I353933,I353540,I353964,I353981,I632819,I353531,I354012,I353534,I353546,I353543,I354101,I710953,I354127,I354144,I354166,I354183,I710968,I710956,I354200,I710947,I354226,I354234,I710959,I354260,I354268,I710950,I354285,I710965,I354325,I354333,I354378,I710974,I710962,I354395,I710971,I354421,I354443,I354460,I354477,I354508,I354525,I354556,I354645,I354671,I354688,I354710,I354727,I354744,I354770,I354778,I354804,I354812,I354829,I354869,I354877,I354922,I354939,I354965,I354987,I355004,I355021,I355052,I355069,I355100,I355189,I907963,I355215,I355232,I355254,I355271,I907975,I355288,I907966,I355314,I355322,I907984,I355348,I355356,I907960,I355373,I907978,I355413,I355421,I355466,I907972,I907969,I355483,I907981,I355509,I355531,I355548,I355565,I355596,I355613,I355644,I355733,I710307,I355759,I355776,I355725,I355798,I355815,I710322,I710310,I355832,I710301,I355858,I355866,I710313,I355892,I355900,I710304,I355917,I355704,I710319,I355957,I355965,I355698,I355713,I356010,I710328,I710316,I356027,I710325,I356053,I355701,I356075,I356092,I356109,I355716,I356140,I356157,I355707,I356188,I355710,I355722,I355719,I356277,I356303,I356320,I356269,I356342,I356359,I356376,I356402,I356410,I356436,I356444,I356461,I356248,I356501,I356509,I356242,I356257,I356554,I356571,I356597,I356245,I356619,I356636,I356653,I356260,I356684,I356701,I356251,I356732,I356254,I356266,I356263,I356821,I1093576,I356847,I356864,I356886,I356903,I1093552,I1093573,I356920,I1093570,I356946,I356954,I1093549,I356980,I356988,I1093561,I357005,I1093564,I357045,I357053,I357098,I1093567,I1093555,I357115,I1093558,I357141,I357163,I357180,I357197,I357228,I357245,I357276,I357365,I838603,I357391,I357408,I357357,I357430,I357447,I838615,I357464,I838606,I357490,I357498,I838624,I357524,I357532,I838600,I357549,I357336,I838618,I357589,I357597,I357330,I357345,I357642,I838612,I838609,I357659,I838621,I357685,I357333,I357707,I357724,I357741,I357348,I357772,I357789,I357339,I357820,I357342,I357354,I357351,I357909,I357935,I357952,I357901,I357974,I357991,I358008,I358034,I358042,I358068,I358076,I358093,I357880,I358133,I358141,I357874,I357889,I358186,I358203,I358229,I357877,I358251,I358268,I358285,I357892,I358316,I358333,I357883,I358364,I357886,I357898,I357895,I358453,I358479,I358496,I358445,I358518,I358535,I358552,I358578,I358586,I358612,I358620,I358637,I358424,I358677,I358685,I358418,I358433,I358730,I358747,I358773,I358421,I358795,I358812,I358829,I358436,I358860,I358877,I358427,I358908,I358430,I358442,I358439,I358997,I754235,I359023,I359040,I358989,I359062,I359079,I754250,I754238,I359096,I754229,I359122,I359130,I754241,I359156,I359164,I754232,I359181,I358968,I754247,I359221,I359229,I358962,I358977,I359274,I754256,I754244,I359291,I754253,I359317,I358965,I359339,I359356,I359373,I358980,I359404,I359421,I358971,I359452,I358974,I358986,I358983,I359541,I359567,I359584,I359533,I359606,I359623,I359640,I359666,I359674,I359700,I359708,I359725,I359512,I359765,I359773,I359506,I359521,I359818,I359835,I359861,I359509,I359883,I359900,I359917,I359524,I359948,I359965,I359515,I359996,I359518,I359530,I359527,I360085,I971169,I360111,I360128,I360077,I360150,I360167,I971181,I971184,I360184,I971187,I360210,I360218,I971172,I360244,I360252,I971178,I360269,I360056,I971166,I360309,I360317,I360050,I360065,I360362,I971190,I360379,I971175,I360405,I360053,I360427,I360444,I360461,I360068,I360492,I360509,I360059,I360540,I360062,I360074,I360071,I360629,I360655,I360672,I360694,I360711,I360728,I360754,I360762,I360788,I360796,I360813,I360853,I360861,I360906,I360923,I360949,I360971,I360988,I361005,I361036,I361053,I361084,I361173,I936285,I361199,I361216,I361165,I361238,I361255,I936297,I361272,I936288,I361298,I361306,I936306,I361332,I361340,I936282,I361357,I361144,I936300,I361397,I361405,I361138,I361153,I361450,I936294,I936291,I361467,I936303,I361493,I361141,I361515,I361532,I361549,I361156,I361580,I361597,I361147,I361628,I361150,I361162,I361159,I361717,I484425,I361743,I361760,I361709,I361782,I361799,I484422,I484443,I361816,I484446,I361842,I361850,I484431,I361876,I361884,I484434,I361901,I361688,I484437,I361941,I361949,I361682,I361697,I361994,I484428,I362011,I484440,I362037,I361685,I362059,I362076,I362093,I361700,I362124,I362141,I361691,I362172,I361694,I361706,I361703,I362261,I838025,I362287,I362304,I362253,I362326,I362343,I838037,I362360,I838028,I362386,I362394,I838046,I362420,I362428,I838022,I362445,I362232,I838040,I362485,I362493,I362226,I362241,I362538,I838034,I838031,I362555,I838043,I362581,I362229,I362603,I362620,I362637,I362244,I362668,I362685,I362235,I362716,I362238,I362250,I362247,I362805,I672335,I362831,I362848,I362797,I362870,I362887,I672329,I672326,I362904,I672341,I362930,I362938,I362964,I362972,I672323,I362989,I362776,I363029,I363037,I362770,I362785,I363082,I672338,I672332,I363099,I363125,I362773,I363147,I363164,I363181,I362788,I363212,I363229,I672344,I362779,I363260,I362782,I362794,I362791,I363349,I642296,I363375,I363392,I363341,I363414,I363431,I642290,I642287,I363448,I642302,I363474,I363482,I363508,I363516,I642284,I363533,I363320,I363573,I363581,I363314,I363329,I363626,I642299,I642293,I363643,I363669,I363317,I363691,I363708,I363725,I363332,I363756,I363773,I642305,I363323,I363804,I363326,I363338,I363335,I363893,I820342,I363919,I363936,I363885,I363958,I363975,I820360,I363992,I820354,I364018,I364026,I820348,I364052,I364060,I820357,I364077,I363864,I820345,I364117,I364125,I363858,I363873,I364170,I820363,I364187,I364213,I363861,I364235,I364252,I364269,I363876,I364300,I364317,I820351,I363867,I364348,I363870,I363882,I363879,I364437,I719997,I364463,I364480,I364429,I364502,I364519,I720012,I720000,I364536,I719991,I364562,I364570,I720003,I364596,I364604,I719994,I364621,I364408,I720009,I364661,I364669,I364402,I364417,I364714,I720018,I720006,I364731,I720015,I364757,I364405,I364779,I364796,I364813,I364420,I364844,I364861,I364411,I364892,I364414,I364426,I364423,I364981,I760695,I365007,I365024,I365046,I365063,I760710,I760698,I365080,I760689,I365106,I365114,I760701,I365140,I365148,I760692,I365165,I760707,I365205,I365213,I365258,I760716,I760704,I365275,I760713,I365301,I365323,I365340,I365357,I365388,I365405,I365436,I365525,I607539,I365551,I365568,I365590,I365607,I607560,I607551,I365624,I365650,I365658,I607545,I365684,I365692,I607542,I365709,I607536,I365749,I365757,I365802,I607548,I365819,I607557,I365845,I365867,I365884,I365901,I365932,I365949,I607554,I365980,I366069,I577483,I366095,I366112,I366061,I366134,I366151,I577504,I577495,I366168,I366194,I366202,I577489,I366228,I366236,I577486,I366253,I366040,I577480,I366293,I366301,I366034,I366049,I366346,I577492,I366363,I577501,I366389,I366037,I366411,I366428,I366445,I366052,I366476,I366493,I577498,I366043,I366524,I366046,I366058,I366055,I366613,I841493,I366639,I366656,I366678,I366695,I841505,I366712,I841496,I366738,I366746,I841514,I366772,I366780,I841490,I366797,I841508,I366837,I366845,I366890,I841502,I841499,I366907,I841511,I366933,I366955,I366972,I366989,I367020,I367037,I367068,I367157,I367183,I367200,I367149,I367222,I367239,I367256,I367282,I367290,I367316,I367324,I367341,I367128,I367381,I367389,I367122,I367137,I367434,I367451,I367477,I367125,I367499,I367516,I367533,I367140,I367564,I367581,I367131,I367612,I367134,I367146,I367143,I367701,I749713,I367727,I367744,I367766,I367783,I749728,I749716,I367800,I749707,I367826,I367834,I749719,I367860,I367868,I749710,I367885,I749725,I367925,I367933,I367978,I749734,I749722,I367995,I749731,I368021,I368043,I368060,I368077,I368108,I368125,I368156,I368245,I368271,I368288,I368237,I368310,I368327,I368344,I368370,I368378,I368404,I368412,I368429,I368216,I368469,I368477,I368210,I368225,I368522,I368539,I368565,I368213,I368587,I368604,I368621,I368228,I368652,I368669,I368219,I368700,I368222,I368234,I368231,I368789,I368815,I368832,I368854,I368871,I368888,I368914,I368922,I368948,I368956,I368973,I369013,I369021,I369066,I369083,I369109,I369131,I369148,I369165,I369196,I369213,I369244,I369333,I984769,I369359,I369376,I369325,I369398,I369415,I984781,I984784,I369432,I984787,I369458,I369466,I984772,I369492,I369500,I984778,I369517,I369304,I984766,I369557,I369565,I369298,I369313,I369610,I984790,I369627,I984775,I369653,I369301,I369675,I369692,I369709,I369316,I369740,I369757,I369307,I369788,I369310,I369322,I369319,I369877,I620689,I369903,I369920,I369942,I369959,I620683,I620680,I369976,I620695,I370002,I370010,I370036,I370044,I620677,I370061,I370101,I370109,I370154,I620692,I620686,I370171,I370197,I370219,I370236,I370253,I370284,I370301,I620698,I370332,I370421,I557253,I370447,I370464,I370413,I370486,I370503,I557274,I557265,I370520,I370546,I370554,I557259,I370580,I370588,I557256,I370605,I370392,I557250,I370645,I370653,I370386,I370401,I370698,I557262,I370715,I557271,I370741,I370389,I370763,I370780,I370797,I370404,I370828,I370845,I557268,I370395,I370876,I370398,I370410,I370407,I370965,I504077,I370991,I371008,I371030,I371047,I504098,I504089,I371064,I371090,I371098,I504083,I371124,I371132,I504080,I371149,I504074,I371189,I371197,I371242,I504086,I371259,I504095,I371285,I371307,I371324,I371341,I371372,I371389,I504092,I371420,I371509,I371535,I371552,I371501,I371574,I371591,I371608,I371634,I371642,I371668,I371676,I371693,I371480,I371733,I371741,I371474,I371489,I371786,I371803,I371829,I371477,I371851,I371868,I371885,I371492,I371916,I371933,I371483,I371964,I371486,I371498,I371495,I372053,I1014024,I372079,I372096,I372045,I372118,I372135,I1014021,I1014018,I372152,I1014006,I372178,I372186,I1014030,I372212,I372220,I1014015,I372237,I372024,I1014009,I372277,I372285,I372018,I372033,I372330,I1014012,I372347,I1014027,I372373,I372021,I372395,I372412,I372429,I372036,I372460,I372477,I372027,I372508,I372030,I372042,I372039,I372597,I1048356,I372623,I372640,I372589,I372662,I372679,I1048332,I1048353,I372696,I1048350,I372722,I372730,I1048329,I372756,I372764,I1048341,I372781,I372568,I1048344,I372821,I372829,I372562,I372577,I372874,I1048347,I1048335,I372891,I1048338,I372917,I372565,I372939,I372956,I372973,I372580,I373004,I373021,I372571,I373052,I372574,I372586,I372583,I373141,I1040026,I373167,I373184,I373133,I373206,I373223,I1040002,I1040023,I373240,I1040020,I373266,I373274,I1039999,I373300,I373308,I1040011,I373325,I373112,I1040014,I373365,I373373,I373106,I373121,I373418,I1040017,I1040005,I373435,I1040008,I373461,I373109,I373483,I373500,I373517,I373124,I373548,I373565,I373115,I373596,I373118,I373130,I373127,I373685,I687618,I373711,I373728,I373677,I373750,I373767,I687612,I687609,I373784,I687624,I373810,I373818,I373844,I373852,I687606,I373869,I373656,I373909,I373917,I373650,I373665,I373962,I687621,I687615,I373979,I374005,I373653,I374027,I374044,I374061,I373668,I374092,I374109,I687627,I373659,I374140,I373662,I373674,I373671,I374229,I896403,I374255,I374272,I374221,I374294,I374311,I896415,I374328,I896406,I374354,I374362,I896424,I374388,I374396,I896400,I374413,I374200,I896418,I374453,I374461,I374194,I374209,I374506,I896412,I896409,I374523,I896421,I374549,I374197,I374571,I374588,I374605,I374212,I374636,I374653,I374203,I374684,I374206,I374218,I374215,I374773,I615631,I374799,I374816,I374765,I374838,I374855,I615652,I615643,I374872,I374898,I374906,I615637,I374932,I374940,I615634,I374957,I374744,I615628,I374997,I375005,I374738,I374753,I375050,I615640,I375067,I615649,I375093,I374741,I375115,I375132,I375149,I374756,I375180,I375197,I615646,I374747,I375228,I374750,I374762,I374759,I375317,I375343,I375360,I375382,I375399,I375416,I375442,I375450,I375476,I375484,I375501,I375541,I375549,I375594,I375611,I375637,I375659,I375676,I375693,I375724,I375741,I375772,I375861,I941487,I375887,I375904,I375853,I375926,I375943,I941499,I375960,I941490,I375986,I375994,I941508,I376020,I376028,I941484,I376045,I375832,I941502,I376085,I376093,I375826,I375841,I376138,I941496,I941493,I376155,I941505,I376181,I375829,I376203,I376220,I376237,I375844,I376268,I376285,I375835,I376316,I375838,I375850,I375847,I376405,I636499,I376431,I376448,I376397,I376470,I376487,I636493,I636490,I376504,I636505,I376530,I376538,I376564,I376572,I636487,I376589,I376376,I376629,I376637,I376370,I376385,I376682,I636502,I636496,I376699,I376725,I376373,I376747,I376764,I376781,I376388,I376812,I376829,I636508,I376379,I376860,I376382,I376394,I376391,I376949,I376975,I376992,I376941,I377014,I377031,I377048,I377074,I377082,I377108,I377116,I377133,I376920,I377173,I377181,I376914,I376929,I377226,I377243,I377269,I376917,I377291,I377308,I377325,I376932,I377356,I377373,I376923,I377404,I376926,I376938,I376935,I377493,I718059,I377519,I377536,I377485,I377558,I377575,I718074,I718062,I377592,I718053,I377618,I377626,I718065,I377652,I377660,I718056,I377677,I377464,I718071,I377717,I377725,I377458,I377473,I377770,I718080,I718068,I377787,I718077,I377813,I377461,I377835,I377852,I377869,I377476,I377900,I377917,I377467,I377948,I377470,I377482,I377479,I378037,I1015180,I378063,I378080,I378029,I378102,I378119,I1015177,I1015174,I378136,I1015162,I378162,I378170,I1015186,I378196,I378204,I1015171,I378221,I378008,I1015165,I378261,I378269,I378002,I378017,I378314,I1015168,I378331,I1015183,I378357,I378005,I378379,I378396,I378413,I378020,I378444,I378461,I378011,I378492,I378014,I378026,I378023,I378581,I832823,I378607,I378624,I378573,I378646,I378663,I832835,I378680,I832826,I378706,I378714,I832844,I378740,I378748,I832820,I378765,I378552,I832838,I378805,I378813,I378546,I378561,I378858,I832832,I832829,I378875,I832841,I378901,I378549,I378923,I378940,I378957,I378564,I378988,I379005,I378555,I379036,I378558,I378570,I378567,I379125,I974977,I379151,I379168,I379190,I379207,I974989,I974992,I379224,I974995,I379250,I379258,I974980,I379284,I379292,I974986,I379309,I974974,I379349,I379357,I379402,I974998,I379419,I974983,I379445,I379467,I379484,I379501,I379532,I379549,I379580,I379669,I379695,I379712,I379661,I379734,I379751,I379768,I379794,I379802,I379828,I379836,I379853,I379640,I379893,I379901,I379634,I379649,I379946,I379963,I379989,I379637,I380011,I380028,I380045,I379652,I380076,I380093,I379643,I380124,I379646,I379658,I379655,I380213,I1014602,I380239,I380256,I380205,I380278,I380295,I1014599,I1014596,I380312,I1014584,I380338,I380346,I1014608,I380372,I380380,I1014593,I380397,I380184,I1014587,I380437,I380445,I380178,I380193,I380490,I1014590,I380507,I1014605,I380533,I380181,I380555,I380572,I380589,I380196,I380620,I380637,I380187,I380668,I380190,I380202,I380199,I380757,I380783,I380800,I380822,I380839,I380856,I380882,I380890,I380916,I380924,I380941,I380981,I380989,I381034,I381051,I381077,I381099,I381116,I381133,I381164,I381181,I381212,I381301,I475755,I381327,I381344,I381293,I381366,I381383,I475752,I475773,I381400,I475776,I381426,I381434,I475761,I381460,I381468,I475764,I381485,I381272,I475767,I381525,I381533,I381266,I381281,I381578,I475758,I381595,I475770,I381621,I381269,I381643,I381660,I381677,I381284,I381708,I381725,I381275,I381756,I381278,I381290,I381287,I381845,I381871,I381888,I381837,I381910,I381927,I381944,I381970,I381978,I382004,I382012,I382029,I381816,I382069,I382077,I381810,I381825,I382122,I382139,I382165,I381813,I382187,I382204,I382221,I381828,I382252,I382269,I381819,I382300,I381822,I381834,I381831,I382389,I382415,I382432,I382381,I382454,I382471,I382488,I382514,I382522,I382548,I382556,I382573,I382360,I382613,I382621,I382354,I382369,I382666,I382683,I382709,I382357,I382731,I382748,I382765,I382372,I382796,I382813,I382363,I382844,I382366,I382378,I382375,I382933,I382959,I382976,I382925,I382998,I383015,I383032,I383058,I383066,I383092,I383100,I383117,I382904,I383157,I383165,I382898,I382913,I383210,I383227,I383253,I382901,I383275,I383292,I383309,I382916,I383340,I383357,I382907,I383388,I382910,I382922,I382919,I383477,I480957,I383503,I383520,I383469,I383542,I383559,I480954,I480975,I383576,I480978,I383602,I383610,I480963,I383636,I383644,I480966,I383661,I383448,I480969,I383701,I383709,I383442,I383457,I383754,I480960,I383771,I480972,I383797,I383445,I383819,I383836,I383853,I383460,I383884,I383901,I383451,I383932,I383454,I383466,I383463,I384021,I384047,I384064,I384013,I384086,I384103,I384120,I384146,I384154,I384180,I384188,I384205,I383992,I384245,I384253,I383986,I384001,I384298,I384315,I384341,I383989,I384363,I384380,I384397,I384004,I384428,I384445,I383995,I384476,I383998,I384010,I384007,I384565,I384591,I384608,I384557,I384630,I384647,I384664,I384690,I384698,I384724,I384732,I384749,I384536,I384789,I384797,I384530,I384545,I384842,I384859,I384885,I384533,I384907,I384924,I384941,I384548,I384972,I384989,I384539,I385020,I384542,I384554,I384551,I385109,I638607,I385135,I385152,I385101,I385174,I385191,I638601,I638598,I385208,I638613,I385234,I385242,I385268,I385276,I638595,I385293,I385080,I385333,I385341,I385074,I385089,I385386,I638610,I638604,I385403,I385429,I385077,I385451,I385468,I385485,I385092,I385516,I385533,I638616,I385083,I385564,I385086,I385098,I385095,I385653,I676551,I385679,I385696,I385645,I385718,I385735,I676545,I676542,I385752,I676557,I385778,I385786,I385812,I385820,I676539,I385837,I385624,I385877,I385885,I385618,I385633,I385930,I676554,I676548,I385947,I385973,I385621,I385995,I386012,I386029,I385636,I386060,I386077,I676560,I385627,I386108,I385630,I385642,I385639,I386197,I657579,I386223,I386240,I386189,I386262,I386279,I657573,I657570,I386296,I657585,I386322,I386330,I386356,I386364,I657567,I386381,I386168,I386421,I386429,I386162,I386177,I386474,I657582,I657576,I386491,I386517,I386165,I386539,I386556,I386573,I386180,I386604,I386621,I657588,I386171,I386652,I386174,I386186,I386183,I386741,I558987,I386767,I386784,I386733,I386806,I386823,I559008,I558999,I386840,I386866,I386874,I558993,I386900,I386908,I558990,I386925,I386712,I558984,I386965,I386973,I386706,I386721,I387018,I558996,I387035,I559005,I387061,I386709,I387083,I387100,I387117,I386724,I387148,I387165,I559002,I386715,I387196,I386718,I386730,I386727,I387285,I387311,I387328,I387350,I387367,I387384,I387410,I387418,I387444,I387452,I387469,I387509,I387517,I387562,I387579,I387605,I387627,I387644,I387661,I387692,I387709,I387740,I387829,I387855,I387872,I387821,I387894,I387911,I387928,I387954,I387962,I387988,I387996,I388013,I387800,I388053,I388061,I387794,I387809,I388106,I388123,I388149,I387797,I388171,I388188,I388205,I387812,I388236,I388253,I387803,I388284,I387806,I387818,I387815,I388373,I837447,I388399,I388416,I388438,I388455,I837459,I388472,I837450,I388498,I388506,I837468,I388532,I388540,I837444,I388557,I837462,I388597,I388605,I388650,I837456,I837453,I388667,I837465,I388693,I388715,I388732,I388749,I388780,I388797,I388828,I388917,I870393,I388943,I388960,I388982,I388999,I870405,I389016,I870396,I389042,I389050,I870414,I389076,I389084,I870390,I389101,I870408,I389141,I389149,I389194,I870402,I870399,I389211,I870411,I389237,I389259,I389276,I389293,I389324,I389341,I389372,I389461,I389487,I389504,I389453,I389526,I389543,I389560,I389586,I389594,I389620,I389628,I389645,I389432,I389685,I389693,I389426,I389441,I389738,I389755,I389781,I389429,I389803,I389820,I389837,I389444,I389868,I389885,I389435,I389916,I389438,I389450,I389447,I390005,I692888,I390031,I390048,I390070,I390087,I692882,I692879,I390104,I692894,I390130,I390138,I390164,I390172,I692876,I390189,I390229,I390237,I390282,I692891,I692885,I390299,I390325,I390347,I390364,I390381,I390412,I390429,I692897,I390460,I390549,I789765,I390575,I390592,I390541,I390614,I390631,I789780,I789768,I390648,I789759,I390674,I390682,I789771,I390708,I390716,I789762,I390733,I390520,I789777,I390773,I390781,I390514,I390529,I390826,I789786,I789774,I390843,I789783,I390869,I390517,I390891,I390908,I390925,I390532,I390956,I390973,I390523,I391004,I390526,I390538,I390535,I391093,I747775,I391119,I391136,I391158,I391175,I747790,I747778,I391192,I747769,I391218,I391226,I747781,I391252,I391260,I747772,I391277,I747787,I391317,I391325,I391370,I747796,I747784,I391387,I747793,I391413,I391435,I391452,I391469,I391500,I391517,I391548,I391637,I560721,I391663,I391680,I391702,I391719,I560742,I560733,I391736,I391762,I391770,I560727,I391796,I391804,I560724,I391821,I560718,I391861,I391869,I391914,I560730,I391931,I560739,I391957,I391979,I391996,I392013,I392044,I392061,I560736,I392092,I392181,I425265,I392207,I392224,I392246,I392263,I425268,I425286,I392280,I425274,I392306,I392314,I392340,I392348,I425283,I392365,I425277,I392405,I392413,I392458,I425280,I425262,I392475,I425271,I392501,I392523,I392540,I392557,I392588,I392605,I392636,I392725,I987489,I392751,I392768,I392717,I392790,I392807,I987501,I987504,I392824,I987507,I392850,I392858,I987492,I392884,I392892,I987498,I392909,I392696,I987486,I392949,I392957,I392690,I392705,I393002,I987510,I393019,I987495,I393045,I392693,I393067,I393084,I393101,I392708,I393132,I393149,I392699,I393180,I392702,I392714,I392711,I393269,I393295,I393312,I393261,I393334,I393351,I393368,I393394,I393402,I393428,I393436,I393453,I393240,I393493,I393501,I393234,I393249,I393546,I393563,I393589,I393237,I393611,I393628,I393645,I393252,I393676,I393693,I393243,I393724,I393246,I393258,I393255,I393813,I643877,I393839,I393856,I393805,I393878,I393895,I643871,I643868,I393912,I643883,I393938,I393946,I393972,I393980,I643865,I393997,I393784,I394037,I394045,I393778,I393793,I394090,I643880,I643874,I394107,I394133,I393781,I394155,I394172,I394189,I393796,I394220,I394237,I643886,I393787,I394268,I393790,I393802,I393799,I394354,I394380,I394397,I394428,I394436,I394453,I394470,I394487,I394504,I394521,I394538,I394569,I394586,I394603,I394648,I394665,I394696,I394713,I394744,I394761,I394778,I394804,I394812,I394843,I394860,I394891,I394949,I394975,I394992,I395023,I395031,I395048,I395065,I395082,I395099,I395116,I395133,I395164,I395181,I395198,I395243,I395260,I395291,I395308,I395339,I395356,I395373,I395399,I395407,I395438,I395455,I395486,I395544,I395570,I395587,I395618,I395626,I395643,I395660,I395677,I395694,I395711,I395728,I395759,I395776,I395793,I395838,I395855,I395886,I395903,I395934,I395951,I395968,I395994,I396002,I396033,I396050,I396081,I396139,I573443,I396165,I396182,I396131,I573437,I396213,I396221,I573434,I396238,I396255,I573446,I396272,I573449,I396289,I396306,I396323,I396128,I396354,I573458,I396371,I573452,I396388,I396113,I396125,I396433,I396450,I396119,I396481,I573440,I396498,I396107,I396529,I573455,I396546,I396563,I396589,I396597,I396116,I396628,I396645,I396122,I396676,I396110,I396734,I692358,I396760,I396777,I692355,I396808,I396816,I396833,I396850,I692352,I396867,I692367,I396884,I396901,I396918,I396949,I692361,I396966,I692349,I396983,I397028,I397045,I397076,I692370,I397093,I397124,I397141,I692364,I397158,I397184,I397192,I397223,I397240,I397271,I397329,I397355,I397372,I397321,I397403,I397411,I397428,I397445,I397462,I397479,I397496,I397513,I397318,I397544,I397561,I397578,I397303,I397315,I397623,I397640,I397309,I397671,I397688,I397297,I397719,I397736,I397753,I397779,I397787,I397306,I397818,I397835,I397312,I397866,I397300,I397924,I908556,I397950,I397967,I908538,I397998,I398006,I908544,I398023,I398040,I908559,I398057,I908550,I398074,I398091,I398108,I398139,I908562,I398156,I908541,I398173,I398218,I398235,I398266,I908547,I398283,I398314,I908553,I398331,I398348,I398374,I398382,I398413,I398430,I398461,I398519,I928208,I398545,I398562,I398511,I928190,I398593,I398601,I928196,I398618,I398635,I928211,I398652,I928202,I398669,I398686,I398703,I398508,I398734,I928214,I398751,I928193,I398768,I398493,I398505,I398813,I398830,I398499,I398861,I928199,I398878,I398487,I398909,I928205,I398926,I398943,I398969,I398977,I398496,I399008,I399025,I398502,I399056,I398490,I399114,I954218,I399140,I399157,I399106,I954200,I399188,I399196,I954206,I399213,I399230,I954221,I399247,I954212,I399264,I399281,I399298,I399103,I399329,I954224,I399346,I954203,I399363,I399088,I399100,I399408,I399425,I399094,I399456,I954209,I399473,I399082,I399504,I954215,I399521,I399538,I399564,I399572,I399091,I399603,I399620,I399097,I399651,I399085,I399709,I399735,I399752,I399783,I399791,I399808,I399825,I399842,I399859,I399876,I399893,I399924,I399941,I399958,I400003,I400020,I400051,I400068,I400099,I400116,I400133,I400159,I400167,I400198,I400215,I400246,I400304,I400330,I400347,I400378,I400386,I400403,I400420,I400437,I400454,I400471,I400488,I400519,I400536,I400553,I400598,I400615,I400646,I400663,I400694,I400711,I400728,I400754,I400762,I400793,I400810,I400841,I400899,I560149,I400925,I400942,I400891,I560143,I400973,I400981,I560140,I400998,I401015,I560152,I401032,I560155,I401049,I401066,I401083,I400888,I401114,I560164,I401131,I560158,I401148,I400873,I400885,I401193,I401210,I400879,I401241,I560146,I401258,I400867,I401289,I560161,I401306,I401323,I401349,I401357,I400876,I401388,I401405,I400882,I401436,I400870,I401494,I401520,I401537,I401486,I401568,I401576,I401593,I401610,I401627,I401644,I401661,I401678,I401483,I401709,I401726,I401743,I401468,I401480,I401788,I401805,I401474,I401836,I401853,I401462,I401884,I401901,I401918,I401944,I401952,I401471,I401983,I402000,I401477,I402031,I401465,I402089,I889482,I402115,I402132,I402081,I889464,I402163,I402171,I889470,I402188,I402205,I889485,I402222,I889476,I402239,I402256,I402273,I402078,I402304,I889488,I402321,I889467,I402338,I402063,I402075,I402383,I402400,I402069,I402431,I889473,I402448,I402057,I402479,I889479,I402496,I402513,I402539,I402547,I402066,I402578,I402595,I402072,I402626,I402060,I402684,I402710,I402727,I402758,I402766,I402783,I402800,I402817,I402834,I402851,I402868,I402899,I402916,I402933,I402978,I402995,I403026,I403043,I403074,I403091,I403108,I403134,I403142,I403173,I403190,I403221,I403279,I933988,I403305,I403322,I403271,I933970,I403353,I403361,I933976,I403378,I403395,I933991,I403412,I933982,I403429,I403446,I403463,I403268,I403494,I933994,I403511,I933973,I403528,I403253,I403265,I403573,I403590,I403259,I403621,I933979,I403638,I403247,I403669,I933985,I403686,I403703,I403729,I403737,I403256,I403768,I403785,I403262,I403816,I403250,I403874,I775562,I403900,I403917,I775550,I403948,I403956,I775547,I403973,I403990,I775559,I404007,I775556,I404024,I404041,I404058,I404089,I775565,I404106,I775568,I404123,I404168,I404185,I404216,I775571,I404233,I404264,I775574,I404281,I775553,I404298,I404324,I404332,I404363,I404380,I404411,I404469,I1081054,I404495,I404512,I404461,I1081060,I404543,I404551,I1081075,I404568,I404585,I1081066,I404602,I1081063,I404619,I404636,I404653,I404458,I404684,I404701,I1081078,I404718,I404443,I404455,I404763,I404780,I404449,I404811,I1081072,I404828,I404437,I404859,I1081057,I404876,I1081069,I404893,I1081081,I404919,I404927,I404446,I404958,I404975,I404452,I405006,I404440,I405064,I1065584,I405090,I405107,I405056,I1065590,I405138,I405146,I1065605,I405163,I405180,I1065596,I405197,I1065593,I405214,I405231,I405248,I405053,I405279,I405296,I1065608,I405313,I405038,I405050,I405358,I405375,I405044,I405406,I1065602,I405423,I405032,I405454,I1065587,I405471,I1065599,I405488,I1065611,I405514,I405522,I405041,I405553,I405570,I405047,I405601,I405035,I405659,I582113,I405685,I405702,I405651,I582107,I405733,I405741,I582104,I405758,I405775,I582116,I405792,I582119,I405809,I405826,I405843,I405648,I405874,I582128,I405891,I582122,I405908,I405633,I405645,I405953,I405970,I405639,I406001,I582110,I406018,I405627,I406049,I582125,I406066,I406083,I406109,I406117,I405636,I406148,I406165,I405642,I406196,I405630,I406254,I565929,I406280,I406297,I565923,I406328,I406336,I565920,I406353,I406370,I565932,I406387,I565935,I406404,I406421,I406438,I406469,I565944,I406486,I565938,I406503,I406548,I406565,I406596,I565926,I406613,I406644,I565941,I406661,I406678,I406704,I406712,I406743,I406760,I406791,I406849,I406875,I406892,I406841,I406923,I406931,I406948,I406965,I406982,I406999,I407016,I407033,I406838,I407064,I407081,I407098,I406823,I406835,I407143,I407160,I406829,I407191,I407208,I406817,I407239,I407256,I407273,I407299,I407307,I406826,I407338,I407355,I406832,I407386,I406820,I407444,I407470,I407487,I407518,I407526,I407543,I407560,I407577,I407594,I407611,I407628,I407659,I407676,I407693,I407738,I407755,I407786,I407803,I407834,I407851,I407868,I407894,I407902,I407933,I407950,I407981,I408039,I556103,I408065,I408082,I556097,I408113,I408121,I556094,I408138,I408155,I556106,I408172,I556109,I408189,I408206,I408223,I408254,I556118,I408271,I556112,I408288,I408333,I408350,I408381,I556100,I408398,I408429,I556115,I408446,I408463,I408489,I408497,I408528,I408545,I408576,I408634,I784606,I408660,I408677,I784594,I408708,I408716,I784591,I408733,I408750,I784603,I408767,I784600,I408784,I408801,I408818,I408849,I784609,I408866,I784612,I408883,I408928,I408945,I408976,I784615,I408993,I409024,I784618,I409041,I784597,I409058,I409084,I409092,I409123,I409140,I409171,I409229,I460727,I409255,I409272,I409221,I460739,I409303,I409311,I460724,I409328,I409345,I460742,I409362,I460733,I409379,I409396,I409413,I409218,I409444,I460745,I409461,I460748,I409478,I409203,I409215,I409523,I409540,I409209,I409571,I409588,I409197,I409619,I460736,I409636,I460730,I409653,I409679,I409687,I409206,I409718,I409735,I409212,I409766,I409200,I409824,I675494,I409850,I409867,I409816,I675491,I409898,I409906,I409923,I409940,I675488,I409957,I675503,I409974,I409991,I410008,I409813,I410039,I675497,I410056,I675485,I410073,I409798,I409810,I410118,I410135,I409804,I410166,I675506,I410183,I409792,I410214,I410231,I675500,I410248,I410274,I410282,I409801,I410313,I410330,I409807,I410361,I409795,I410419,I410445,I410462,I410411,I410493,I410501,I410518,I410535,I410552,I410569,I410586,I410603,I410408,I410634,I410651,I410668,I410393,I410405,I410713,I410730,I410399,I410761,I410778,I410387,I410809,I410826,I410843,I410869,I410877,I410396,I410908,I410925,I410402,I410956,I410390,I411014,I463039,I411040,I411057,I463051,I411088,I411096,I463036,I411113,I411130,I463054,I411147,I463045,I411164,I411181,I411198,I411229,I463057,I411246,I463060,I411263,I411308,I411325,I411356,I411373,I411404,I463048,I411421,I463042,I411438,I411464,I411472,I411503,I411520,I411551,I411609,I910868,I411635,I411652,I910850,I411683,I411691,I910856,I411708,I411725,I910871,I411742,I910862,I411759,I411776,I411793,I411824,I910874,I411841,I910853,I411858,I411903,I411920,I411951,I910859,I411968,I411999,I910865,I412016,I412033,I412059,I412067,I412098,I412115,I412146,I412204,I412230,I412247,I412278,I412286,I412303,I412320,I412337,I412354,I412371,I412388,I412419,I412436,I412453,I412498,I412515,I412546,I412563,I412594,I412611,I412628,I412654,I412662,I412693,I412710,I412741,I412799,I412825,I412842,I412791,I412873,I412881,I412898,I412915,I412932,I412949,I412966,I412983,I412788,I413014,I413031,I413048,I412773,I412785,I413093,I413110,I412779,I413141,I413158,I412767,I413189,I413206,I413223,I413249,I413257,I412776,I413288,I413305,I412782,I413336,I412770,I413394,I827074,I413420,I413437,I413386,I827077,I413468,I413476,I827080,I413493,I413510,I827092,I413527,I827083,I413544,I413561,I413578,I413383,I413609,I827089,I413626,I413643,I413368,I413380,I413688,I413705,I413374,I413736,I413753,I413362,I413784,I827086,I413801,I413818,I827095,I413844,I413852,I413371,I413883,I413900,I413377,I413931,I413365,I413989,I816976,I414015,I414032,I413981,I816979,I414063,I414071,I816982,I414088,I414105,I816994,I414122,I816985,I414139,I414156,I414173,I413978,I414204,I816991,I414221,I414238,I413963,I413975,I414283,I414300,I413969,I414331,I414348,I413957,I414379,I816988,I414396,I414413,I816997,I414439,I414447,I413966,I414478,I414495,I413972,I414526,I413960,I414584,I932254,I414610,I414627,I414576,I932236,I414658,I414666,I932242,I414683,I414700,I932257,I414717,I932248,I414734,I414751,I414768,I414573,I414799,I932260,I414816,I932239,I414833,I414558,I414570,I414878,I414895,I414564,I414926,I932245,I414943,I414552,I414974,I932251,I414991,I415008,I415034,I415042,I414561,I415073,I415090,I414567,I415121,I414555,I415179,I659684,I415205,I415222,I415171,I659681,I415253,I415261,I415278,I415295,I659678,I415312,I659693,I415329,I415346,I415363,I415168,I415394,I659687,I415411,I659675,I415428,I415153,I415165,I415473,I415490,I415159,I415521,I659696,I415538,I415147,I415569,I415586,I659690,I415603,I415629,I415637,I415156,I415668,I415685,I415162,I415716,I415150,I415774,I415800,I415817,I415766,I415848,I415856,I415873,I415890,I415907,I415924,I415941,I415958,I415763,I415989,I416006,I416023,I415748,I415760,I416068,I416085,I415754,I416116,I416133,I415742,I416164,I416181,I416198,I416224,I416232,I415751,I416263,I416280,I415757,I416311,I415745,I416369,I556681,I416395,I416412,I416361,I556675,I416443,I416451,I556672,I416468,I416485,I556684,I416502,I556687,I416519,I416536,I416553,I416358,I416584,I556696,I416601,I556690,I416618,I416343,I416355,I416663,I416680,I416349,I416711,I556678,I416728,I416337,I416759,I556693,I416776,I416793,I416819,I416827,I416346,I416858,I416875,I416352,I416906,I416340,I416964,I416990,I417007,I416956,I417038,I417046,I417063,I417080,I417097,I417114,I417131,I417148,I416953,I417179,I417196,I417213,I416938,I416950,I417258,I417275,I416944,I417306,I417323,I416932,I417354,I417371,I417388,I417414,I417422,I416941,I417453,I417470,I416947,I417501,I416935,I417559,I828792,I417585,I417602,I417551,I828774,I417633,I417641,I828780,I417658,I417675,I828795,I417692,I828786,I417709,I417726,I417743,I417548,I417774,I828798,I417791,I828777,I417808,I417533,I417545,I417853,I417870,I417539,I417901,I828783,I417918,I417527,I417949,I828789,I417966,I417983,I418009,I418017,I417536,I418048,I418065,I417542,I418096,I417530,I418154,I418180,I418197,I418228,I418236,I418253,I418270,I418287,I418304,I418321,I418338,I418369,I418386,I418403,I418448,I418465,I418496,I418513,I418544,I418561,I418578,I418604,I418612,I418643,I418660,I418691,I418749,I748430,I418775,I418792,I748418,I418823,I418831,I748415,I418848,I418865,I748427,I418882,I748424,I418899,I418916,I418933,I418964,I748433,I418981,I748436,I418998,I419043,I419060,I419091,I748439,I419108,I419139,I748442,I419156,I748421,I419173,I419199,I419207,I419238,I419255,I419286,I419344,I939190,I419370,I419387,I939172,I419418,I419426,I939178,I419443,I419460,I939193,I419477,I939184,I419494,I419511,I419528,I419559,I939196,I419576,I939175,I419593,I419638,I419655,I419686,I939181,I419703,I419734,I939187,I419751,I419768,I419794,I419802,I419833,I419850,I419881,I419939,I866940,I419965,I419982,I419931,I866922,I420013,I420021,I866928,I420038,I420055,I866943,I420072,I866934,I420089,I420106,I420123,I419928,I420154,I866946,I420171,I866925,I420188,I419913,I419925,I420233,I420250,I419919,I420281,I866931,I420298,I419907,I420329,I866937,I420346,I420363,I420389,I420397,I419916,I420428,I420445,I419922,I420476,I419910,I420534,I420560,I420577,I420526,I420608,I420616,I420633,I420650,I420667,I420684,I420701,I420718,I420523,I420749,I420766,I420783,I420508,I420520,I420828,I420845,I420514,I420876,I420893,I420502,I420924,I420941,I420958,I420984,I420992,I420511,I421023,I421040,I420517,I421071,I420505,I421129,I1019795,I421155,I421172,I1019801,I421203,I421211,I1019789,I421228,I421245,I1019792,I421262,I1019798,I421279,I421296,I421313,I421344,I421361,I1019807,I421378,I421423,I421440,I421471,I1019786,I421488,I421519,I1019810,I421536,I421553,I1019804,I421579,I421587,I421618,I421635,I421666,I421724,I996097,I421750,I421767,I996103,I421798,I421806,I996091,I421823,I421840,I996094,I421857,I996100,I421874,I421891,I421908,I421939,I421956,I996109,I421973,I422018,I422035,I422066,I996088,I422083,I422114,I996112,I422131,I422148,I996106,I422174,I422182,I422213,I422230,I422261,I422319,I442231,I422345,I422362,I422311,I442243,I422393,I422401,I442228,I422418,I422435,I442246,I422452,I442237,I422469,I422486,I422503,I422308,I422534,I442249,I422551,I442252,I422568,I422293,I422305,I422613,I422630,I422299,I422661,I422678,I422287,I422709,I442240,I422726,I442234,I422743,I422769,I422777,I422296,I422808,I422825,I422302,I422856,I422290,I422914,I422940,I422957,I422906,I422988,I422996,I423013,I423030,I423047,I423064,I423081,I423098,I422903,I423129,I423146,I423163,I422888,I422900,I423208,I423225,I422894,I423256,I423273,I422882,I423304,I423321,I423338,I423364,I423372,I422891,I423403,I423420,I422897,I423451,I422885,I423509,I423535,I423552,I423501,I423583,I423591,I423608,I423625,I423642,I423659,I423676,I423693,I423498,I423724,I423741,I423758,I423483,I423495,I423803,I423820,I423489,I423851,I423868,I423477,I423899,I423916,I423933,I423959,I423967,I423486,I423998,I424015,I423492,I424046,I423480,I424104,I534139,I424130,I424147,I534133,I424178,I424186,I534130,I424203,I424220,I534142,I424237,I534145,I424254,I424271,I424288,I424319,I534154,I424336,I534148,I424353,I424398,I424415,I424446,I534136,I424463,I424494,I534151,I424511,I424528,I424554,I424562,I424593,I424610,I424641,I424699,I424725,I424742,I424691,I424773,I424781,I424798,I424815,I424832,I424849,I424866,I424883,I424688,I424914,I424931,I424948,I424673,I424685,I424993,I425010,I424679,I425041,I425058,I424667,I425089,I425106,I425123,I425149,I425157,I424676,I425188,I425205,I424682,I425236,I424670,I425294,I425320,I425337,I425368,I425376,I425393,I425410,I425427,I425444,I425461,I425478,I425509,I425526,I425543,I425588,I425605,I425636,I425653,I425684,I425701,I425718,I425744,I425752,I425783,I425800,I425831,I425889,I762642,I425915,I425932,I425881,I762630,I425963,I425971,I762627,I425988,I426005,I762639,I426022,I762636,I426039,I426056,I426073,I425878,I426104,I762645,I426121,I762648,I426138,I425863,I425875,I426183,I426200,I425869,I426231,I762651,I426248,I425857,I426279,I762654,I426296,I762633,I426313,I426339,I426347,I425866,I426378,I426395,I425872,I426426,I425860,I426484,I426510,I426527,I426476,I426558,I426566,I426583,I426600,I426617,I426634,I426651,I426668,I426473,I426699,I426716,I426733,I426458,I426470,I426778,I426795,I426464,I426826,I426843,I426452,I426874,I426891,I426908,I426934,I426942,I426461,I426973,I426990,I426467,I427021,I426455,I427079,I707732,I427105,I427122,I427071,I707720,I427153,I427161,I707717,I427178,I427195,I707729,I427212,I707726,I427229,I427246,I427263,I427068,I427294,I707735,I427311,I707738,I427328,I427053,I427065,I427373,I427390,I427059,I427421,I707741,I427438,I427047,I427469,I707744,I427486,I707723,I427503,I427529,I427537,I427056,I427568,I427585,I427062,I427616,I427050,I427674,I427700,I427717,I427666,I427748,I427756,I427773,I427790,I427807,I427824,I427841,I427858,I427663,I427889,I427906,I427923,I427648,I427660,I427968,I427985,I427654,I428016,I428033,I427642,I428064,I428081,I428098,I428124,I428132,I427651,I428163,I428180,I427657,I428211,I427645,I428269,I667589,I428295,I428312,I428261,I667586,I428343,I428351,I428368,I428385,I667583,I428402,I667598,I428419,I428436,I428453,I428258,I428484,I667592,I428501,I667580,I428518,I428243,I428255,I428563,I428580,I428249,I428611,I667601,I428628,I428237,I428659,I428676,I667595,I428693,I428719,I428727,I428246,I428758,I428775,I428252,I428806,I428240,I428864,I528937,I428890,I428907,I428856,I528931,I428938,I428946,I528928,I428963,I428980,I528940,I428997,I528943,I429014,I429031,I429048,I428853,I429079,I528952,I429096,I528946,I429113,I428838,I428850,I429158,I429175,I428844,I429206,I528934,I429223,I428832,I429254,I528949,I429271,I429288,I429314,I429322,I428841,I429353,I429370,I428847,I429401,I428835,I429459,I687088,I429485,I429502,I429451,I687085,I429533,I429541,I429558,I429575,I687082,I429592,I687097,I429609,I429626,I429643,I429448,I429674,I687091,I429691,I687079,I429708,I429433,I429445,I429753,I429770,I429439,I429801,I687100,I429818,I429427,I429849,I429866,I687094,I429883,I429909,I429917,I429436,I429948,I429965,I429442,I429996,I429430,I430054,I430080,I430097,I430128,I430136,I430153,I430170,I430187,I430204,I430221,I430238,I430269,I430286,I430303,I430348,I430365,I430396,I430413,I430444,I430461,I430478,I430504,I430512,I430543,I430560,I430591,I430649,I887170,I430675,I430692,I430641,I887152,I430723,I430731,I887158,I430748,I430765,I887173,I430782,I887164,I430799,I430816,I430833,I430638,I430864,I887176,I430881,I887155,I430898,I430623,I430635,I430943,I430960,I430629,I430991,I887161,I431008,I430617,I431039,I887167,I431056,I431073,I431099,I431107,I430626,I431138,I431155,I430632,I431186,I430620,I431244,I431270,I431287,I431236,I431318,I431326,I431343,I431360,I431377,I431394,I431411,I431428,I431233,I431459,I431476,I431493,I431218,I431230,I431538,I431555,I431224,I431586,I431603,I431212,I431634,I431651,I431668,I431694,I431702,I431221,I431733,I431750,I431227,I431781,I431215,I431839,I431865,I431882,I431831,I431913,I431921,I431938,I431955,I431972,I431989,I432006,I432023,I431828,I432054,I432071,I432088,I431813,I431825,I432133,I432150,I431819,I432181,I432198,I431807,I432229,I432246,I432263,I432289,I432297,I431816,I432328,I432345,I431822,I432376,I431810,I432434,I968464,I432460,I432468,I968458,I432494,I432502,I968467,I432519,I968446,I432536,I432553,I968455,I432570,I432420,I432601,I432618,I432635,I968470,I432652,I968449,I432417,I432408,I432697,I432411,I432405,I432742,I968452,I432759,I432776,I432414,I432807,I968461,I432824,I432841,I432867,I432875,I432402,I432426,I432920,I432937,I432954,I432423,I433012,I433038,I433046,I433072,I433080,I433097,I433114,I433131,I433148,I433179,I433196,I433213,I433230,I433275,I433320,I433337,I433354,I433385,I433402,I433419,I433445,I433453,I433498,I433515,I433532,I433590,I817558,I433616,I433624,I817549,I433650,I433658,I817543,I433675,I817555,I433692,I433709,I817546,I433726,I433576,I433757,I433774,I433791,I817552,I433808,I817537,I433573,I433564,I433853,I433567,I433561,I433898,I433915,I433932,I433570,I433963,I817540,I433980,I433997,I434023,I434031,I433558,I433582,I434076,I434093,I434110,I433579,I434168,I664951,I434194,I434202,I434228,I434236,I664948,I434253,I664963,I434270,I434287,I664957,I434304,I434335,I434352,I434369,I664954,I434386,I664945,I434431,I434476,I664966,I434493,I434510,I434541,I434558,I434575,I664960,I434601,I434609,I434654,I434671,I434688,I434746,I434772,I434780,I434806,I434814,I434831,I434848,I434865,I434882,I434732,I434913,I434930,I434947,I434964,I434729,I434720,I435009,I434723,I434717,I435054,I435071,I435088,I434726,I435119,I435136,I435153,I435179,I435187,I434714,I434738,I435232,I435249,I435266,I434735,I435324,I435350,I435358,I435384,I435392,I435409,I435426,I435443,I435460,I435491,I435508,I435525,I435542,I435587,I435632,I435649,I435666,I435697,I435714,I435731,I435757,I435765,I435810,I435827,I435844,I435902,I435928,I435936,I435962,I435970,I435987,I436004,I436021,I436038,I436069,I436086,I436103,I436120,I436165,I436210,I436227,I436244,I436275,I436292,I436309,I436335,I436343,I436388,I436405,I436422,I436480,I436506,I436514,I436540,I436548,I436565,I436582,I436599,I436616,I436466,I436647,I436664,I436681,I436698,I436463,I436454,I436743,I436457,I436451,I436788,I436805,I436822,I436460,I436853,I436870,I436887,I436913,I436921,I436448,I436472,I436966,I436983,I437000,I436469,I437058,I1027113,I437084,I437092,I1027131,I437118,I437126,I1027128,I437143,I1027119,I437160,I437177,I1027116,I437194,I437044,I437225,I437242,I437259,I1027122,I437276,I1027137,I437041,I437032,I437321,I437035,I437029,I437366,I437383,I437400,I437038,I437431,I1027134,I437448,I1027125,I437465,I1027140,I437491,I437499,I437026,I437050,I437544,I437561,I437578,I437047,I437636,I587306,I437662,I437670,I587318,I437696,I437704,I587309,I437721,I587312,I437738,I437755,I587315,I437772,I437622,I437803,I437820,I437837,I437854,I587321,I437619,I437610,I437899,I437613,I437607,I437944,I587327,I437961,I437978,I437616,I438009,I438026,I587324,I438043,I587330,I438069,I438077,I437604,I437628,I438122,I438139,I438156,I437625,I438214,I923566,I438240,I438248,I923572,I438274,I438282,I438299,I923569,I438316,I438333,I923587,I438350,I438381,I438398,I438415,I923590,I438432,I438477,I438522,I923575,I438539,I438556,I438587,I923581,I438604,I923578,I438621,I923584,I438647,I438655,I438700,I438717,I438734,I438792,I846114,I438818,I438826,I846120,I438852,I438860,I438877,I846117,I438894,I438911,I846135,I438928,I438959,I438976,I438993,I846138,I439010,I439055,I439100,I846123,I439117,I439134,I439165,I846129,I439182,I846126,I439199,I846132,I439225,I439233,I439278,I439295,I439312,I439370,I980432,I439396,I439404,I980426,I439430,I439438,I980435,I439455,I980414,I439472,I439489,I980423,I439506,I439356,I439537,I439554,I439571,I980438,I439588,I980417,I439353,I439344,I439633,I439347,I439341,I439678,I980420,I439695,I439712,I439350,I439743,I980429,I439760,I439777,I439803,I439811,I439338,I439362,I439856,I439873,I439890,I439359,I439948,I948420,I439974,I439982,I948426,I440008,I440016,I440033,I948423,I440050,I440067,I948441,I440084,I439934,I440115,I440132,I440149,I948444,I440166,I439931,I439922,I440211,I439925,I439919,I440256,I948429,I440273,I440290,I439928,I440321,I948435,I440338,I948432,I440355,I948438,I440381,I440389,I439916,I439940,I440434,I440451,I440468,I439937,I440526,I1021503,I440552,I440560,I1021521,I440586,I440594,I1021518,I440611,I1021509,I440628,I440645,I1021506,I440662,I440693,I440710,I440727,I1021512,I440744,I1021527,I440789,I440834,I440851,I440868,I440899,I1021524,I440916,I1021515,I440933,I1021530,I440959,I440967,I441012,I441029,I441046,I441104,I441130,I441138,I441164,I441172,I441189,I441206,I441223,I441240,I441090,I441271,I441288,I441305,I441322,I441087,I441078,I441367,I441081,I441075,I441412,I441429,I441446,I441084,I441477,I441494,I441511,I441537,I441545,I441072,I441096,I441590,I441607,I441624,I441093,I441682,I523148,I441708,I441716,I523160,I441742,I441750,I523151,I441767,I523154,I441784,I441801,I523157,I441818,I441668,I441849,I441866,I441883,I441900,I523163,I441665,I441656,I441945,I441659,I441653,I441990,I523169,I442007,I442024,I441662,I442055,I442072,I523166,I442089,I523172,I442115,I442123,I441650,I441674,I442168,I442185,I442202,I441671,I442260,I442286,I442294,I442320,I442328,I442345,I442362,I442379,I442396,I442427,I442444,I442461,I442478,I442523,I442568,I442585,I442602,I442633,I442650,I442667,I442693,I442701,I442746,I442763,I442780,I442838,I953044,I442864,I442872,I953050,I442898,I442906,I442923,I953047,I442940,I442957,I953065,I442974,I442824,I443005,I443022,I443039,I953068,I443056,I442821,I442812,I443101,I442815,I442809,I443146,I953053,I443163,I443180,I442818,I443211,I953059,I443228,I953056,I443245,I953062,I443271,I443279,I442806,I442830,I443324,I443341,I443358,I442827,I443416,I913740,I443442,I443450,I913746,I443476,I443484,I443501,I913743,I443518,I443535,I913761,I443552,I443402,I443583,I443600,I443617,I913764,I443634,I443399,I443390,I443679,I443393,I443387,I443724,I913749,I443741,I443758,I443396,I443789,I913755,I443806,I913752,I443823,I913758,I443849,I443857,I443384,I443408,I443902,I443919,I443936,I443405,I443994,I854206,I444020,I444028,I854212,I444054,I444062,I444079,I854209,I444096,I444113,I854227,I444130,I443980,I444161,I444178,I444195,I854230,I444212,I443977,I443968,I444257,I443971,I443965,I444302,I854215,I444319,I444336,I443974,I444367,I854221,I444384,I854218,I444401,I854224,I444427,I444435,I443962,I443986,I444480,I444497,I444514,I443983,I444572,I979344,I444598,I444606,I979338,I444632,I444640,I979347,I444657,I979326,I444674,I444691,I979335,I444708,I444739,I444756,I444773,I979350,I444790,I979329,I444835,I444880,I979332,I444897,I444914,I444945,I979341,I444962,I444979,I445005,I445013,I445058,I445075,I445092,I445150,I1034644,I445176,I445184,I445210,I445218,I1034668,I445235,I1034650,I445252,I445269,I1034665,I445286,I445136,I445317,I445334,I445351,I1034647,I445368,I1034656,I445133,I445124,I445413,I445127,I445121,I445458,I1034653,I445475,I445492,I445130,I445523,I1034662,I445540,I1034671,I445557,I1034659,I445583,I445591,I445118,I445142,I445636,I445653,I445670,I445139,I445728,I861142,I445754,I445762,I861148,I445788,I445796,I445813,I861145,I445830,I445847,I861163,I445864,I445714,I445895,I445912,I445929,I861166,I445946,I445711,I445702,I445991,I445705,I445699,I446036,I861151,I446053,I446070,I445708,I446101,I861157,I446118,I861154,I446135,I861160,I446161,I446169,I445696,I445720,I446214,I446231,I446248,I445717,I446306,I699971,I446332,I446340,I699968,I446366,I446374,I699965,I446391,I699992,I446408,I446425,I699980,I446442,I446292,I446473,I446490,I446507,I699986,I446524,I699977,I446289,I446280,I446569,I446283,I446277,I446614,I699974,I446631,I446648,I446286,I446679,I699989,I446696,I699983,I446713,I446739,I446747,I446274,I446298,I446792,I446809,I446826,I446295,I446884,I857096,I446910,I446918,I857102,I446944,I446952,I446969,I857099,I446986,I447003,I857117,I447020,I447051,I447068,I447085,I857120,I447102,I447147,I447192,I857105,I447209,I447226,I447257,I857111,I447274,I857108,I447291,I857114,I447317,I447325,I447370,I447387,I447404,I447462,I818119,I447488,I447496,I818110,I447522,I447530,I818104,I447547,I818116,I447564,I447581,I818107,I447598,I447448,I447629,I447646,I447663,I818113,I447680,I818098,I447445,I447436,I447725,I447439,I447433,I447770,I447787,I447804,I447442,I447835,I818101,I447852,I447869,I447895,I447903,I447430,I447454,I447948,I447965,I447982,I447451,I448040,I448066,I448074,I448100,I448108,I448125,I448142,I448159,I448176,I448207,I448224,I448241,I448258,I448303,I448348,I448365,I448382,I448413,I448430,I448447,I448473,I448481,I448526,I448543,I448560,I448618,I448644,I448652,I448678,I448686,I448703,I448720,I448737,I448754,I448604,I448785,I448802,I448819,I448836,I448601,I448592,I448881,I448595,I448589,I448926,I448943,I448960,I448598,I448991,I449008,I449025,I449051,I449059,I448586,I448610,I449104,I449121,I449138,I448607,I449196,I574012,I449222,I449230,I574024,I449256,I449264,I574015,I449281,I574018,I449298,I449315,I574021,I449332,I449182,I449363,I449380,I449397,I449414,I574027,I449179,I449170,I449459,I449173,I449167,I449504,I574033,I449521,I449538,I449176,I449569,I449586,I574030,I449603,I574036,I449629,I449637,I449164,I449188,I449682,I449699,I449716,I449185,I449774,I449800,I449808,I449834,I449842,I449859,I449876,I449893,I449910,I449760,I449941,I449958,I449975,I449992,I449757,I449748,I450037,I449751,I449745,I450082,I450099,I450116,I449754,I450147,I450164,I450181,I450207,I450215,I449742,I449766,I450260,I450277,I450294,I449763,I450352,I1036429,I450378,I450386,I450412,I450420,I1036453,I450437,I1036435,I450454,I450471,I1036450,I450488,I450338,I450519,I450536,I450553,I1036432,I450570,I1036441,I450335,I450326,I450615,I450329,I450323,I450660,I1036438,I450677,I450694,I450332,I450725,I1036447,I450742,I1036456,I450759,I1036444,I450785,I450793,I450320,I450344,I450838,I450855,I450872,I450341,I450930,I511588,I450956,I450964,I511600,I450990,I450998,I511591,I451015,I511594,I451032,I451049,I511597,I451066,I450916,I451097,I451114,I451131,I451148,I511603,I450913,I450904,I451193,I450907,I450901,I451238,I511609,I451255,I451272,I450910,I451303,I451320,I511606,I451337,I511612,I451363,I451371,I450898,I450922,I451416,I451433,I451450,I450919,I451508,I659154,I451534,I451542,I451568,I451576,I659151,I451593,I659166,I451610,I451627,I659160,I451644,I451494,I451675,I451692,I451709,I659157,I451726,I659148,I451491,I451482,I451771,I451485,I451479,I451816,I659169,I451833,I451850,I451488,I451881,I451898,I451915,I659163,I451941,I451949,I451476,I451500,I451994,I452011,I452028,I451497,I452086,I707077,I452112,I452120,I707074,I452146,I452154,I707071,I452171,I707098,I452188,I452205,I707086,I452222,I452072,I452253,I452270,I452287,I707092,I452304,I707083,I452069,I452060,I452349,I452063,I452057,I452394,I707080,I452411,I452428,I452066,I452459,I707095,I452476,I707089,I452493,I452519,I452527,I452054,I452078,I452572,I452589,I452606,I452075,I452664,I635966,I452690,I452698,I452724,I452732,I635963,I452749,I635978,I452766,I452783,I635972,I452800,I452650,I452831,I452848,I452865,I635969,I452882,I635960,I452647,I452638,I452927,I452641,I452635,I452972,I635981,I452989,I453006,I452644,I453037,I453054,I453071,I635975,I453097,I453105,I452632,I452656,I453150,I453167,I453184,I452653,I453242,I978800,I453268,I453276,I978794,I453302,I453310,I978803,I453327,I978782,I453344,I453361,I978791,I453378,I453228,I453409,I453426,I453443,I978806,I453460,I978785,I453225,I453216,I453505,I453219,I453213,I453550,I978788,I453567,I453584,I453222,I453615,I978797,I453632,I453649,I453675,I453683,I453210,I453234,I453728,I453745,I453762,I453231,I453820,I453846,I453854,I453880,I453888,I453905,I453922,I453939,I453956,I453806,I453987,I454004,I454021,I454038,I453803,I453794,I454083,I453797,I453791,I454128,I454145,I454162,I453800,I454193,I454210,I454227,I454253,I454261,I453788,I453812,I454306,I454323,I454340,I453809,I454398,I963568,I454424,I454432,I963562,I454458,I454466,I963571,I454483,I963550,I454500,I454517,I963559,I454534,I454384,I454565,I454582,I454599,I963574,I454616,I963553,I454381,I454372,I454661,I454375,I454369,I454706,I963556,I454723,I454740,I454378,I454771,I963565,I454788,I454805,I454831,I454839,I454366,I454390,I454884,I454901,I454918,I454387,I454976,I735501,I455002,I455010,I735498,I455036,I455044,I735495,I455061,I735522,I455078,I455095,I735510,I455112,I454962,I455143,I455160,I455177,I735516,I455194,I735507,I454959,I454950,I455239,I454953,I454947,I455284,I735504,I455301,I455318,I454956,I455349,I735519,I455366,I735513,I455383,I455409,I455417,I454944,I454968,I455462,I455479,I455496,I454965,I455554,I524882,I455580,I455588,I524894,I455614,I455622,I524885,I455639,I524888,I455656,I455673,I524891,I455690,I455540,I455721,I455738,I455755,I455772,I524897,I455537,I455528,I455817,I455531,I455525,I455862,I524903,I455879,I455896,I455534,I455927,I455944,I524900,I455961,I524906,I455987,I455995,I455522,I455546,I456040,I456057,I456074,I455543,I456132,I1052494,I456158,I456166,I456192,I456200,I1052518,I456217,I1052500,I456234,I456251,I1052515,I456268,I456299,I456316,I456333,I1052497,I456350,I1052506,I456395,I456440,I1052503,I456457,I456474,I456505,I1052512,I456522,I1052521,I456539,I1052509,I456565,I456573,I456618,I456635,I456652,I456710,I456736,I456744,I456770,I456778,I456795,I456812,I456829,I456846,I456877,I456894,I456911,I456928,I456973,I457018,I457035,I457052,I457083,I457100,I457117,I457143,I457151,I457196,I457213,I457230,I457288,I895244,I457314,I457322,I895250,I457348,I457356,I457373,I895247,I457390,I457407,I895265,I457424,I457274,I457455,I457472,I457489,I895268,I457506,I457271,I457262,I457551,I457265,I457259,I457596,I895253,I457613,I457630,I457268,I457661,I895259,I457678,I895256,I457695,I895262,I457721,I457729,I457256,I457280,I457774,I457791,I457808,I457277,I457866,I457892,I457900,I457926,I457934,I457951,I457968,I457985,I458002,I457852,I458033,I458050,I458067,I458084,I457849,I457840,I458129,I457843,I457837,I458174,I458191,I458208,I457846,I458239,I458256,I458273,I458299,I458307,I457834,I457858,I458352,I458369,I458386,I457855,I458444,I873280,I458470,I458478,I873286,I458504,I458512,I458529,I873283,I458546,I458563,I873301,I458580,I458611,I458628,I458645,I873304,I458662,I458707,I458752,I873289,I458769,I458786,I458817,I873295,I458834,I873292,I458851,I873298,I458877,I458885,I458930,I458947,I458964,I459022,I1010550,I459048,I459056,I1010562,I459082,I459090,I1010553,I459107,I1010541,I459124,I459141,I1010538,I459158,I459008,I459189,I459206,I459223,I1010544,I459240,I459005,I458996,I459285,I458999,I458993,I459330,I1010559,I459347,I459364,I459002,I459395,I1010547,I459412,I459429,I1010556,I459455,I459463,I458990,I459014,I459508,I459525,I459542,I459011,I459600,I459626,I459634,I459660,I459668,I459685,I459702,I459719,I459736,I459767,I459784,I459801,I459818,I459863,I459908,I459925,I459942,I459973,I459990,I460007,I460033,I460041,I460086,I460103,I460120,I460178,I460204,I460212,I460238,I460246,I460263,I460280,I460297,I460314,I460164,I460345,I460362,I460379,I460396,I460161,I460152,I460441,I460155,I460149,I460486,I460503,I460520,I460158,I460551,I460568,I460585,I460611,I460619,I460146,I460170,I460664,I460681,I460698,I460167,I460756,I884262,I460782,I460790,I884268,I460816,I460824,I460841,I884265,I460858,I460875,I884283,I460892,I460923,I460940,I460957,I884286,I460974,I461019,I461064,I884271,I461081,I461098,I461129,I884277,I461146,I884274,I461163,I884280,I461189,I461197,I461242,I461259,I461276,I461334,I712245,I461360,I461368,I712242,I461394,I461402,I712239,I461419,I712266,I461436,I461453,I712254,I461470,I461501,I461518,I461535,I712260,I461552,I712251,I461597,I461642,I712248,I461659,I461676,I461707,I712263,I461724,I712257,I461741,I461767,I461775,I461820,I461837,I461854,I461912,I461938,I461946,I461972,I461980,I461997,I462014,I462031,I462048,I461898,I462079,I462096,I462113,I462130,I461895,I461886,I462175,I461889,I461883,I462220,I462237,I462254,I461892,I462285,I462302,I462319,I462345,I462353,I461880,I461904,I462398,I462415,I462432,I461901,I462490,I1056659,I462516,I462524,I462550,I462558,I1056683,I462575,I1056665,I462592,I462609,I1056680,I462626,I462657,I462674,I462691,I1056662,I462708,I1056671,I462753,I462798,I1056668,I462815,I462832,I462863,I1056677,I462880,I1056686,I462897,I1056674,I462923,I462931,I462976,I462993,I463010,I463068,I463094,I463102,I463128,I463136,I463153,I463170,I463187,I463204,I463235,I463252,I463269,I463286,I463331,I463376,I463393,I463410,I463441,I463458,I463475,I463501,I463509,I463554,I463571,I463588,I463646,I1047139,I463672,I463680,I463706,I463714,I1047163,I463731,I1047145,I463748,I463765,I1047160,I463782,I463632,I463813,I463830,I463847,I1047142,I463864,I1047151,I463629,I463620,I463909,I463623,I463617,I463954,I1047148,I463971,I463988,I463626,I464019,I1047157,I464036,I1047166,I464053,I1047154,I464079,I464087,I463614,I463638,I464132,I464149,I464166,I463635,I464224,I554360,I464250,I464258,I554372,I464284,I464292,I554363,I464309,I554366,I464326,I464343,I554369,I464360,I464210,I464391,I464408,I464425,I464442,I554375,I464207,I464198,I464487,I464201,I464195,I464532,I554381,I464549,I464566,I464204,I464597,I464614,I554378,I464631,I554384,I464657,I464665,I464192,I464216,I464710,I464727,I464744,I464213,I464802,I464828,I464836,I464862,I464870,I464887,I464904,I464921,I464938,I464969,I464986,I465003,I465020,I465065,I465110,I465127,I465144,I465175,I465192,I465209,I465235,I465243,I465288,I465305,I465322,I465380,I1041784,I465406,I465414,I465440,I465448,I1041808,I465465,I1041790,I465482,I465499,I1041805,I465516,I465547,I465564,I465581,I1041787,I465598,I1041796,I465643,I465688,I1041793,I465705,I465722,I465753,I1041802,I465770,I1041811,I465787,I1041799,I465813,I465821,I465866,I465883,I465900,I465958,I590196,I465984,I465992,I590208,I466018,I466026,I590199,I466043,I590202,I466060,I466077,I590205,I466094,I466125,I466142,I466159,I466176,I590211,I466221,I466266,I590217,I466283,I466300,I466331,I466348,I590214,I466365,I590220,I466391,I466399,I466444,I466461,I466478,I466536,I539332,I466562,I466570,I539344,I466596,I466604,I539335,I466621,I539338,I466638,I466655,I539341,I466672,I466522,I466703,I466720,I466737,I466754,I539347,I466519,I466510,I466799,I466513,I466507,I466844,I539353,I466861,I466878,I466516,I466909,I466926,I539350,I466943,I539356,I466969,I466977,I466504,I466528,I467022,I467039,I467056,I466525,I467114,I467140,I467148,I467174,I467182,I467199,I467216,I467233,I467250,I467281,I467298,I467315,I467332,I467377,I467422,I467439,I467456,I467487,I467504,I467521,I467547,I467555,I467600,I467617,I467634,I467692,I467718,I467726,I467752,I467760,I467777,I467794,I467811,I467828,I467678,I467859,I467876,I467893,I467910,I467675,I467666,I467955,I467669,I467663,I468000,I468017,I468034,I467672,I468065,I468082,I468099,I468125,I468133,I467660,I467684,I468178,I468195,I468212,I467681,I468270,I468296,I468304,I468330,I468338,I468355,I468372,I468389,I468406,I468256,I468437,I468454,I468471,I468488,I468253,I468244,I468533,I468247,I468241,I468578,I468595,I468612,I468250,I468643,I468660,I468677,I468703,I468711,I468238,I468262,I468756,I468773,I468790,I468259,I468848,I880794,I468874,I468882,I880800,I468908,I468916,I468933,I880797,I468950,I468967,I880815,I468984,I469015,I469032,I469049,I880818,I469066,I469111,I469156,I880803,I469173,I469190,I469221,I880809,I469238,I880806,I469255,I880812,I469281,I469289,I469334,I469351,I469368,I469426,I469452,I469460,I469486,I469494,I469511,I469528,I469545,I469562,I469412,I469593,I469610,I469627,I469644,I469409,I469400,I469689,I469403,I469397,I469734,I469751,I469768,I469406,I469799,I469816,I469833,I469859,I469867,I469394,I469418,I469912,I469929,I469946,I469415,I470004,I470030,I470038,I470064,I470072,I470089,I470106,I470123,I470140,I469990,I470171,I470188,I470205,I470222,I469987,I469978,I470267,I469981,I469975,I470312,I470329,I470346,I469984,I470377,I470394,I470411,I470437,I470445,I469972,I469996,I470490,I470507,I470524,I469993,I470582,I470608,I470616,I470642,I470650,I470667,I470684,I470701,I470718,I470568,I470749,I470766,I470783,I470800,I470565,I470556,I470845,I470559,I470553,I470890,I470907,I470924,I470562,I470955,I470972,I470989,I471015,I471023,I470550,I470574,I471068,I471085,I471102,I470571,I471160,I471186,I471194,I471220,I471228,I471245,I471262,I471279,I471296,I471327,I471344,I471361,I471378,I471423,I471468,I471485,I471502,I471533,I471550,I471567,I471593,I471601,I471646,I471663,I471680,I471738,I471764,I471772,I471798,I471806,I471823,I471840,I471857,I471874,I471905,I471922,I471939,I471956,I472001,I472046,I472063,I472080,I472111,I472128,I472145,I472171,I472179,I472224,I472241,I472258,I472316,I946686,I472342,I472350,I946692,I472376,I472384,I472401,I946689,I472418,I472435,I946707,I472452,I472302,I472483,I472500,I472517,I946710,I472534,I472299,I472290,I472579,I472293,I472287,I472624,I946695,I472641,I472658,I472296,I472689,I946701,I472706,I946698,I472723,I946704,I472749,I472757,I472284,I472308,I472802,I472819,I472836,I472305,I472894,I472920,I472928,I472954,I472962,I472979,I472996,I473013,I473030,I472880,I473061,I473078,I473095,I473112,I472877,I472868,I473157,I472871,I472865,I473202,I473219,I473236,I472874,I473267,I473284,I473301,I473327,I473335,I472862,I472886,I473380,I473397,I473414,I472883,I473472,I974448,I473498,I473506,I974442,I473532,I473540,I974451,I473557,I974430,I473574,I473591,I974439,I473608,I473639,I473656,I473673,I974454,I473690,I974433,I473735,I473780,I974436,I473797,I473814,I473845,I974445,I473862,I473879,I473905,I473913,I473958,I473975,I473992,I474050,I732917,I474076,I474084,I732914,I474110,I474118,I732911,I474135,I732938,I474152,I474169,I732926,I474186,I474217,I474234,I474251,I732932,I474268,I732923,I474313,I474358,I732920,I474375,I474392,I474423,I732935,I474440,I732929,I474457,I474483,I474491,I474536,I474553,I474570,I474628,I474654,I474662,I474688,I474696,I474713,I474730,I474747,I474764,I474614,I474795,I474812,I474829,I474846,I474611,I474602,I474891,I474605,I474599,I474936,I474953,I474970,I474608,I475001,I475018,I475035,I475061,I475069,I474596,I474620,I475114,I475131,I475148,I474617,I475206,I475232,I475240,I475266,I475274,I475291,I475308,I475325,I475342,I475192,I475373,I475390,I475407,I475424,I475189,I475180,I475469,I475183,I475177,I475514,I475531,I475548,I475186,I475579,I475596,I475613,I475639,I475647,I475174,I475198,I475692,I475709,I475726,I475195,I475784,I475810,I475818,I475844,I475852,I475869,I475886,I475903,I475920,I475951,I475968,I475985,I476002,I476047,I476092,I476109,I476126,I476157,I476174,I476191,I476217,I476225,I476270,I476287,I476304,I476362,I1023186,I476388,I476396,I1023204,I476422,I476430,I1023201,I476447,I1023192,I476464,I476481,I1023189,I476498,I476529,I476546,I476563,I1023195,I476580,I1023210,I476625,I476670,I476687,I476704,I476735,I1023207,I476752,I1023198,I476769,I1023213,I476795,I476803,I476848,I476865,I476882,I476940,I476966,I476974,I477000,I477008,I477025,I477042,I477059,I477076,I477107,I477124,I477141,I477158,I477203,I477248,I477265,I477282,I477313,I477330,I477347,I477373,I477381,I477426,I477443,I477460,I477518,I714183,I477544,I477552,I714180,I477578,I477586,I714177,I477603,I714204,I477620,I477637,I714192,I477654,I477504,I477685,I477702,I477719,I714198,I477736,I714189,I477501,I477492,I477781,I477495,I477489,I477826,I714186,I477843,I477860,I477498,I477891,I714201,I477908,I714195,I477925,I477951,I477959,I477486,I477510,I478004,I478021,I478038,I477507,I478096,I478122,I478130,I478156,I478164,I478181,I478198,I478215,I478232,I478082,I478263,I478280,I478297,I478314,I478079,I478070,I478359,I478073,I478067,I478404,I478421,I478438,I478076,I478469,I478486,I478503,I478529,I478537,I478064,I478088,I478582,I478599,I478616,I478085,I478674,I602334,I478700,I478708,I602346,I478734,I478742,I602337,I478759,I602340,I478776,I478793,I602343,I478810,I478660,I478841,I478858,I478875,I478892,I602349,I478657,I478648,I478937,I478651,I478645,I478982,I602355,I478999,I479016,I478654,I479047,I479064,I602352,I479081,I602358,I479107,I479115,I478642,I478666,I479160,I479177,I479194,I478663,I479252,I705139,I479278,I479286,I705136,I479312,I479320,I705133,I479337,I705160,I479354,I479371,I705148,I479388,I479419,I479436,I479453,I705154,I479470,I705145,I479515,I479560,I705142,I479577,I479594,I479625,I705157,I479642,I705151,I479659,I479685,I479693,I479738,I479755,I479772,I479830,I479856,I479864,I479890,I479898,I479915,I479932,I479949,I479966,I479997,I480014,I480031,I480048,I480093,I480138,I480155,I480172,I480203,I480220,I480237,I480263,I480271,I480316,I480333,I480350,I480408,I1022625,I480434,I480442,I1022643,I480468,I480476,I1022640,I480493,I1022631,I480510,I480527,I1022628,I480544,I480394,I480575,I480592,I480609,I1022634,I480626,I1022649,I480391,I480382,I480671,I480385,I480379,I480716,I480733,I480750,I480388,I480781,I1022646,I480798,I1022637,I480815,I1022652,I480841,I480849,I480376,I480400,I480894,I480911,I480928,I480397,I480986,I481012,I481020,I481046,I481054,I481071,I481088,I481105,I481122,I481153,I481170,I481187,I481204,I481249,I481294,I481311,I481328,I481359,I481376,I481393,I481419,I481427,I481472,I481489,I481506,I481564,I1073319,I481590,I481598,I481624,I481632,I1073343,I481649,I1073325,I481666,I481683,I1073340,I481700,I481550,I481731,I481748,I481765,I1073322,I481782,I1073331,I481547,I481538,I481827,I481541,I481535,I481872,I1073328,I481889,I481906,I481544,I481937,I1073337,I481954,I1073346,I481971,I1073334,I481997,I482005,I481532,I481556,I482050,I482067,I482084,I481553,I482142,I482168,I482176,I482202,I482210,I482227,I482244,I482261,I482278,I482128,I482309,I482326,I482343,I482360,I482125,I482116,I482405,I482119,I482113,I482450,I482467,I482484,I482122,I482515,I482532,I482549,I482575,I482583,I482110,I482134,I482628,I482645,I482662,I482131,I482720,I482746,I482754,I482780,I482788,I482805,I482822,I482839,I482856,I482887,I482904,I482921,I482938,I482983,I483028,I483045,I483062,I483093,I483110,I483127,I483153,I483161,I483206,I483223,I483240,I483298,I516790,I483324,I483332,I516802,I483358,I483366,I516793,I483383,I516796,I483400,I483417,I516799,I483434,I483284,I483465,I483482,I483499,I483516,I516805,I483281,I483272,I483561,I483275,I483269,I483606,I516811,I483623,I483640,I483278,I483671,I483688,I516808,I483705,I516814,I483731,I483739,I483266,I483290,I483784,I483801,I483818,I483287,I483876,I633331,I483902,I483910,I483936,I483944,I633328,I483961,I633343,I483978,I483995,I633337,I484012,I483862,I484043,I484060,I484077,I633334,I484094,I633325,I483859,I483850,I484139,I483853,I483847,I484184,I633346,I484201,I484218,I483856,I484249,I484266,I484283,I633340,I484309,I484317,I483844,I483868,I484362,I484379,I484396,I483865,I484454,I484480,I484488,I484514,I484522,I484539,I484556,I484573,I484590,I484621,I484638,I484655,I484672,I484717,I484762,I484779,I484796,I484827,I484844,I484861,I484887,I484895,I484940,I484957,I484974,I485032,I989164,I485058,I485066,I989176,I485092,I485100,I989167,I485117,I989155,I485134,I485151,I989152,I485168,I485199,I485216,I485233,I989158,I485250,I485295,I485340,I989173,I485357,I485374,I485405,I989161,I485422,I485439,I989170,I485465,I485473,I485518,I485535,I485552,I485610,I485636,I485644,I485670,I485678,I485695,I485712,I485729,I485746,I485596,I485777,I485794,I485811,I485828,I485593,I485584,I485873,I485587,I485581,I485918,I485935,I485952,I485590,I485983,I486000,I486017,I486043,I486051,I485578,I485602,I486096,I486113,I486130,I485599,I486188,I486214,I486222,I486248,I486256,I486273,I486290,I486307,I486324,I486174,I486355,I486372,I486389,I486406,I486171,I486162,I486451,I486165,I486159,I486496,I486513,I486530,I486168,I486561,I486578,I486595,I486621,I486629,I486156,I486180,I486674,I486691,I486708,I486177,I486766,I486792,I486800,I486826,I486834,I486851,I486868,I486885,I486902,I486933,I486950,I486967,I486984,I487029,I487074,I487091,I487108,I487139,I487156,I487173,I487199,I487207,I487252,I487269,I487286,I487344,I677072,I487370,I487378,I487404,I487412,I677069,I487429,I677084,I487446,I487463,I677078,I487480,I487511,I487528,I487545,I677075,I487562,I677066,I487607,I487652,I677087,I487669,I487686,I487717,I487734,I487751,I677081,I487777,I487785,I487830,I487847,I487864,I487922,I487948,I487956,I487982,I487990,I488007,I488024,I488041,I488058,I488089,I488106,I488123,I488140,I488185,I488230,I488247,I488264,I488295,I488312,I488329,I488355,I488363,I488408,I488425,I488442,I488500,I488526,I488534,I488560,I488568,I488585,I488602,I488619,I488636,I488486,I488667,I488684,I488701,I488718,I488483,I488474,I488763,I488477,I488471,I488808,I488825,I488842,I488480,I488873,I488890,I488907,I488933,I488941,I488468,I488492,I488986,I489003,I489020,I488489,I489078,I489104,I489112,I489138,I489146,I489163,I489180,I489197,I489214,I489245,I489262,I489279,I489296,I489341,I489386,I489403,I489420,I489451,I489468,I489485,I489511,I489519,I489564,I489581,I489598,I489656,I1083434,I489682,I489690,I489716,I489724,I1083458,I489741,I1083440,I489758,I489775,I1083455,I489792,I489823,I489840,I489857,I1083437,I489874,I1083446,I489919,I489964,I1083443,I489981,I489998,I490029,I1083452,I490046,I1083461,I490063,I1083449,I490089,I490097,I490142,I490159,I490176,I490234,I490260,I490268,I490294,I490302,I490319,I490336,I490353,I490370,I490401,I490418,I490435,I490452,I490497,I490542,I490559,I490576,I490607,I490624,I490641,I490667,I490675,I490720,I490737,I490754,I490812,I1007082,I490838,I490846,I1007094,I490872,I490880,I1007085,I490897,I1007073,I490914,I490931,I1007070,I490948,I490798,I490979,I490996,I491013,I1007076,I491030,I490795,I490786,I491075,I490789,I490783,I491120,I1007091,I491137,I491154,I490792,I491185,I1007079,I491202,I491219,I1007088,I491245,I491253,I490780,I490804,I491298,I491315,I491332,I490801,I491390,I548002,I491416,I491424,I548014,I491450,I491458,I548005,I491475,I548008,I491492,I491509,I548011,I491526,I491557,I491574,I491591,I491608,I548017,I491653,I491698,I548023,I491715,I491732,I491763,I491780,I548020,I491797,I548026,I491823,I491831,I491876,I491893,I491910,I491968,I491994,I492002,I492028,I492036,I492053,I492070,I492087,I492104,I491954,I492135,I492152,I492169,I492186,I491951,I491942,I492231,I491945,I491939,I492276,I492293,I492310,I491948,I492341,I492358,I492375,I492401,I492409,I491936,I491960,I492454,I492471,I492488,I491957,I492546,I613316,I492572,I492580,I613328,I492606,I492614,I613319,I492631,I613322,I492648,I492665,I613325,I492682,I492713,I492730,I492747,I492764,I613331,I492809,I492854,I613337,I492871,I492888,I492919,I492936,I613334,I492953,I613340,I492979,I492987,I493032,I493049,I493066,I493124,I493150,I493158,I493184,I493192,I493209,I493226,I493243,I493260,I493110,I493291,I493308,I493325,I493342,I493107,I493098,I493387,I493101,I493095,I493432,I493449,I493466,I493104,I493497,I493514,I493531,I493557,I493565,I493092,I493116,I493610,I493627,I493644,I493113,I493702,I587884,I493728,I493736,I587896,I493762,I493770,I587887,I493787,I587890,I493804,I493821,I587893,I493838,I493688,I493869,I493886,I493903,I493920,I587899,I493685,I493676,I493965,I493679,I493673,I494010,I587905,I494027,I494044,I493682,I494075,I494092,I587902,I494109,I587908,I494135,I494143,I493670,I493694,I494188,I494205,I494222,I493691,I494280,I869234,I494306,I494314,I869240,I494340,I494348,I494365,I869237,I494382,I494399,I869255,I494416,I494266,I494447,I494464,I494481,I869258,I494498,I494263,I494254,I494543,I494257,I494251,I494588,I869243,I494605,I494622,I494260,I494653,I869249,I494670,I869246,I494687,I869252,I494713,I494721,I494248,I494272,I494766,I494783,I494800,I494269,I494858,I799045,I494884,I494892,I799036,I494918,I494926,I799030,I494943,I799042,I494960,I494977,I799033,I494994,I495025,I495042,I495059,I799039,I495076,I799024,I495121,I495166,I495183,I495200,I495231,I799027,I495248,I495265,I495291,I495299,I495344,I495361,I495378,I495436,I495462,I495470,I495496,I495504,I495521,I495538,I495555,I495572,I495603,I495620,I495637,I495654,I495699,I495744,I495761,I495778,I495809,I495826,I495843,I495869,I495877,I495922,I495939,I495956,I496014,I496040,I496048,I496074,I496082,I496099,I496116,I496133,I496150,I496000,I496181,I496198,I496215,I496232,I495997,I495988,I496277,I495991,I495985,I496322,I496339,I496356,I495994,I496387,I496404,I496421,I496447,I496455,I495982,I496006,I496500,I496517,I496534,I496003,I496592,I892372,I496618,I496626,I496643,I892354,I892366,I496660,I892369,I496686,I496694,I892363,I892360,I496720,I496728,I496745,I496762,I496779,I892378,I496819,I496827,I496844,I496861,I496878,I496909,I892357,I496926,I496952,I496960,I496991,I497022,I497039,I497070,I892375,I497170,I497196,I497204,I497221,I497238,I497264,I497272,I497298,I497306,I497323,I497340,I497357,I497153,I497397,I497405,I497422,I497439,I497456,I497156,I497487,I497504,I497530,I497538,I497138,I497569,I497147,I497600,I497617,I497159,I497648,I497150,I497141,I497144,I497162,I497748,I497774,I497782,I497799,I497816,I497842,I497850,I497876,I497884,I497901,I497918,I497935,I497731,I497975,I497983,I498000,I498017,I498034,I497734,I498065,I498082,I498108,I498116,I497716,I498147,I497725,I498178,I498195,I497737,I498226,I497728,I497719,I497722,I497740,I498326,I1089411,I498352,I498360,I498377,I1089396,I1089384,I498394,I1089399,I498420,I498428,I1089402,I498454,I498462,I498479,I498496,I498513,I498309,I1089390,I498553,I498561,I498578,I498595,I498612,I498312,I498643,I1089387,I1089393,I498660,I1089408,I498686,I498694,I498294,I498725,I498303,I498756,I498773,I498315,I498804,I1089405,I498306,I498297,I498300,I498318,I498904,I891794,I498930,I498938,I498955,I891776,I891788,I498972,I891791,I498998,I499006,I891785,I891782,I499032,I499040,I499057,I499074,I499091,I891800,I499131,I499139,I499156,I499173,I499190,I499221,I891779,I499238,I499264,I499272,I499303,I499334,I499351,I499382,I891797,I499482,I499508,I499516,I499533,I499550,I499576,I499584,I499610,I499618,I499635,I499652,I499669,I499709,I499717,I499734,I499751,I499768,I499799,I499816,I499842,I499850,I499881,I499912,I499929,I499960,I500060,I869830,I500086,I500094,I500111,I869812,I869824,I500128,I869827,I500154,I500162,I869821,I869818,I500188,I500196,I500213,I500230,I500247,I869836,I500287,I500295,I500312,I500329,I500346,I500377,I869815,I500394,I500420,I500428,I500459,I500490,I500507,I500538,I869833,I500638,I500664,I500672,I500689,I500706,I500732,I500740,I500766,I500774,I500791,I500808,I500825,I500865,I500873,I500890,I500907,I500924,I500955,I500972,I500998,I501006,I501037,I501068,I501085,I501116,I501216,I501242,I501250,I501267,I501284,I501310,I501318,I501344,I501352,I501369,I501386,I501403,I501443,I501451,I501468,I501485,I501502,I501533,I501550,I501576,I501584,I501615,I501646,I501663,I501694,I501794,I501820,I501828,I501845,I501862,I501888,I501896,I501922,I501930,I501947,I501964,I501981,I501777,I502021,I502029,I502046,I502063,I502080,I501780,I502111,I502128,I502154,I502162,I501762,I502193,I501771,I502224,I502241,I501783,I502272,I501774,I501765,I501768,I501786,I502372,I828214,I502398,I502406,I502423,I828196,I828208,I502440,I828211,I502466,I502474,I828205,I828202,I502500,I502508,I502525,I502542,I502559,I502355,I828220,I502599,I502607,I502624,I502641,I502658,I502358,I502689,I828199,I502706,I502732,I502740,I502340,I502771,I502349,I502802,I502819,I502361,I502850,I828217,I502352,I502343,I502346,I502364,I502950,I1076916,I502976,I502984,I503001,I1076901,I1076889,I503018,I1076904,I503044,I503052,I1076907,I503078,I503086,I503103,I503120,I503137,I1076895,I503177,I503185,I503202,I503219,I503236,I503267,I1076892,I1076898,I503284,I1076913,I503310,I503318,I503349,I503380,I503397,I503428,I1076910,I503528,I503554,I503562,I503579,I503596,I503622,I503630,I503656,I503664,I503681,I503698,I503715,I503511,I503755,I503763,I503780,I503797,I503814,I503514,I503845,I503862,I503888,I503896,I503496,I503927,I503505,I503958,I503975,I503517,I504006,I503508,I503499,I503502,I503520,I504106,I504132,I504140,I504157,I504174,I504200,I504208,I504234,I504242,I504259,I504276,I504293,I504333,I504341,I504358,I504375,I504392,I504423,I504440,I504466,I504474,I504505,I504536,I504553,I504584,I504684,I504710,I504718,I504735,I504752,I504778,I504786,I504812,I504820,I504837,I504854,I504871,I504667,I504911,I504919,I504936,I504953,I504970,I504670,I505001,I505018,I505044,I505052,I504652,I505083,I504661,I505114,I505131,I504673,I505162,I504664,I504655,I504658,I504676,I505262,I505288,I505296,I505313,I505330,I505356,I505364,I505390,I505398,I505415,I505432,I505449,I505245,I505489,I505497,I505514,I505531,I505548,I505248,I505579,I505596,I505622,I505630,I505230,I505661,I505239,I505692,I505709,I505251,I505740,I505242,I505233,I505236,I505254,I505840,I505866,I505874,I505891,I505908,I505934,I505942,I505968,I505976,I505993,I506010,I506027,I505823,I506067,I506075,I506092,I506109,I506126,I505826,I506157,I506174,I506200,I506208,I505808,I506239,I505817,I506270,I506287,I505829,I506318,I505820,I505811,I505814,I505832,I506418,I506444,I506452,I506469,I506486,I506512,I506520,I506546,I506554,I506571,I506588,I506605,I506645,I506653,I506670,I506687,I506704,I506735,I506752,I506778,I506786,I506817,I506848,I506865,I506896,I506996,I801835,I507022,I507030,I507047,I801832,I801850,I507064,I801847,I507090,I507098,I801829,I507124,I507132,I507149,I507166,I507183,I506979,I801841,I507223,I507231,I507248,I507265,I507282,I506982,I507313,I801844,I507330,I507356,I507364,I506964,I507395,I506973,I507426,I507443,I506985,I507474,I801838,I506976,I506967,I506970,I506988,I507574,I833994,I507600,I507608,I507625,I833976,I833988,I507642,I833991,I507668,I507676,I833985,I833982,I507702,I507710,I507727,I507744,I507761,I834000,I507801,I507809,I507826,I507843,I507860,I507891,I833979,I507908,I507934,I507942,I507973,I508004,I508021,I508052,I833997,I508152,I508178,I508186,I508203,I508220,I508246,I508254,I508280,I508288,I508305,I508322,I508339,I508379,I508387,I508404,I508421,I508438,I508469,I508486,I508512,I508520,I508551,I508582,I508599,I508630,I508730,I508756,I508764,I508781,I508798,I508824,I508832,I508858,I508866,I508883,I508900,I508917,I508957,I508965,I508982,I508999,I509016,I509047,I509064,I509090,I509098,I509129,I509160,I509177,I509208,I509308,I509334,I509342,I509359,I509376,I509402,I509410,I509436,I509444,I509461,I509478,I509495,I509535,I509543,I509560,I509577,I509594,I509625,I509642,I509668,I509676,I509707,I509738,I509755,I509786,I509886,I918960,I509912,I509920,I509937,I918942,I918954,I509954,I918957,I509980,I509988,I918951,I918948,I510014,I510022,I510039,I510056,I510073,I509869,I918966,I510113,I510121,I510138,I510155,I510172,I509872,I510203,I918945,I510220,I510246,I510254,I509854,I510285,I509863,I510316,I510333,I509875,I510364,I918963,I509866,I509857,I509860,I509878,I510464,I956478,I510490,I510498,I510515,I956481,I956490,I510532,I956493,I510558,I510566,I956502,I956484,I510592,I510600,I510617,I510634,I510651,I510447,I510691,I510699,I510716,I510733,I510750,I510450,I510781,I956499,I510798,I956496,I510824,I510832,I510432,I510863,I510441,I510894,I510911,I510453,I510942,I956487,I510444,I510435,I510438,I510456,I511042,I511068,I511076,I511093,I511110,I511136,I511144,I511170,I511178,I511195,I511212,I511229,I511269,I511277,I511294,I511311,I511328,I511359,I511376,I511402,I511410,I511441,I511472,I511489,I511520,I511620,I511646,I511654,I511671,I511688,I511714,I511722,I511748,I511756,I511773,I511790,I511807,I511847,I511855,I511872,I511889,I511906,I511937,I511954,I511980,I511988,I512019,I512050,I512067,I512098,I512198,I512224,I512232,I512249,I512266,I512292,I512300,I512326,I512334,I512351,I512368,I512385,I512181,I512425,I512433,I512450,I512467,I512484,I512184,I512515,I512532,I512558,I512566,I512166,I512597,I512175,I512628,I512645,I512187,I512676,I512178,I512169,I512172,I512190,I512776,I512802,I512810,I512827,I512844,I512870,I512878,I512904,I512912,I512929,I512946,I512963,I512759,I513003,I513011,I513028,I513045,I513062,I512762,I513093,I513110,I513136,I513144,I512744,I513175,I512753,I513206,I513223,I512765,I513254,I512756,I512747,I512750,I512768,I513354,I513380,I513388,I513405,I513422,I513448,I513456,I513482,I513490,I513507,I513524,I513541,I513581,I513589,I513606,I513623,I513640,I513671,I513688,I513714,I513722,I513753,I513784,I513801,I513832,I513932,I513958,I513966,I513983,I514000,I514026,I514034,I514060,I514068,I514085,I514102,I514119,I513915,I514159,I514167,I514184,I514201,I514218,I513918,I514249,I514266,I514292,I514300,I513900,I514331,I513909,I514362,I514379,I513921,I514410,I513912,I513903,I513906,I513924,I514510,I514536,I514544,I514561,I514578,I514604,I514612,I514638,I514646,I514663,I514680,I514697,I514737,I514745,I514762,I514779,I514796,I514827,I514844,I514870,I514878,I514909,I514940,I514957,I514988,I515088,I830526,I515114,I515122,I515139,I830508,I830520,I515156,I830523,I515182,I515190,I830517,I830514,I515216,I515224,I515241,I515258,I515275,I830532,I515315,I515323,I515340,I515357,I515374,I515405,I830511,I515422,I515448,I515456,I515487,I515518,I515535,I515566,I830529,I515666,I1094171,I515692,I515700,I515717,I1094156,I1094144,I515734,I1094159,I515760,I515768,I1094162,I515794,I515802,I515819,I515836,I515853,I1094150,I515893,I515901,I515918,I515935,I515952,I515983,I1094147,I1094153,I516000,I1094168,I516026,I516034,I516065,I516096,I516113,I516144,I1094165,I516244,I516270,I516278,I516295,I516312,I516338,I516346,I516372,I516380,I516397,I516414,I516431,I516227,I516471,I516479,I516496,I516513,I516530,I516230,I516561,I516578,I516604,I516612,I516212,I516643,I516221,I516674,I516691,I516233,I516722,I516224,I516215,I516218,I516236,I516822,I643353,I516848,I516856,I516873,I643341,I643359,I516890,I643356,I516916,I516924,I643347,I643344,I516950,I516958,I516975,I516992,I517009,I643338,I517049,I517057,I517074,I517091,I517108,I517139,I517156,I517182,I517190,I517221,I517252,I517269,I517300,I643350,I517400,I757483,I517426,I517434,I517451,I757459,I757474,I517468,I757486,I517494,I517502,I757471,I757462,I517528,I517536,I517553,I517570,I517587,I517383,I517627,I517635,I517652,I517669,I517686,I517386,I517717,I757477,I757468,I517734,I757480,I517760,I517768,I517368,I517799,I517377,I517830,I517847,I517389,I517878,I757465,I517380,I517371,I517374,I517392,I517978,I930520,I518004,I518012,I518029,I930502,I930514,I518046,I930517,I518072,I518080,I930511,I930508,I518106,I518114,I518131,I518148,I518165,I517961,I930526,I518205,I518213,I518230,I518247,I518264,I517964,I518295,I930505,I518312,I518338,I518346,I517946,I518377,I517955,I518408,I518425,I517967,I518456,I930523,I517958,I517949,I517952,I517970,I518556,I518582,I518590,I518607,I518624,I518650,I518658,I518684,I518692,I518709,I518726,I518743,I518783,I518791,I518808,I518825,I518842,I518873,I518890,I518916,I518924,I518955,I518986,I519003,I519034,I519134,I519160,I519168,I519185,I519202,I519228,I519236,I519262,I519270,I519287,I519304,I519321,I519117,I519361,I519369,I519386,I519403,I519420,I519120,I519451,I519468,I519494,I519502,I519102,I519533,I519111,I519564,I519581,I519123,I519612,I519114,I519105,I519108,I519126,I519712,I758775,I519738,I519746,I519763,I758751,I758766,I519780,I758778,I519806,I519814,I758763,I758754,I519840,I519848,I519865,I519882,I519899,I519695,I519939,I519947,I519964,I519981,I519998,I519698,I520029,I758769,I758760,I520046,I758772,I520072,I520080,I519680,I520111,I519689,I520142,I520159,I519701,I520190,I758757,I519692,I519683,I519686,I519704,I520290,I520316,I520324,I520341,I520358,I520384,I520392,I520418,I520426,I520443,I520460,I520477,I520273,I520517,I520525,I520542,I520559,I520576,I520276,I520607,I520624,I520650,I520658,I520258,I520689,I520267,I520720,I520737,I520279,I520768,I520270,I520261,I520264,I520282,I520868,I520894,I520902,I520919,I520936,I520962,I520970,I520996,I521004,I521021,I521038,I521055,I521095,I521103,I521120,I521137,I521154,I521185,I521202,I521228,I521236,I521267,I521298,I521315,I521346,I521446,I842086,I521472,I521480,I521497,I842068,I842080,I521514,I842083,I521540,I521548,I842077,I842074,I521574,I521582,I521599,I521616,I521633,I842092,I521673,I521681,I521698,I521715,I521732,I521763,I842071,I521780,I521806,I521814,I521845,I521876,I521893,I521924,I842089,I522024,I932832,I522050,I522058,I522075,I932814,I932826,I522092,I932829,I522118,I522126,I932823,I932820,I522152,I522160,I522177,I522194,I522211,I522007,I932838,I522251,I522259,I522276,I522293,I522310,I522010,I522341,I932817,I522358,I522384,I522392,I521992,I522423,I522001,I522454,I522471,I522013,I522502,I932835,I522004,I521995,I521998,I522016,I522602,I522628,I522636,I522653,I522670,I522696,I522704,I522730,I522738,I522755,I522772,I522789,I522585,I522829,I522837,I522854,I522871,I522888,I522588,I522919,I522936,I522962,I522970,I522570,I523001,I522579,I523032,I523049,I522591,I523080,I522582,I522573,I522576,I522594,I523180,I523206,I523214,I523231,I523248,I523274,I523282,I523308,I523316,I523333,I523350,I523367,I523407,I523415,I523432,I523449,I523466,I523497,I523514,I523540,I523548,I523579,I523610,I523627,I523658,I523758,I653893,I523784,I523792,I523809,I653881,I653899,I523826,I653896,I523852,I523860,I653887,I653884,I523886,I523894,I523911,I523928,I523945,I523741,I653878,I523985,I523993,I524010,I524027,I524044,I523744,I524075,I524092,I524118,I524126,I523726,I524157,I523735,I524188,I524205,I523747,I524236,I653890,I523738,I523729,I523732,I523750,I524336,I909134,I524362,I524370,I524387,I909116,I909128,I524404,I909131,I524430,I524438,I909125,I909122,I524464,I524472,I524489,I524506,I524523,I909140,I524563,I524571,I524588,I524605,I524622,I524653,I909119,I524670,I524696,I524704,I524735,I524766,I524783,I524814,I909137,I524914,I992620,I524940,I524948,I524965,I992644,I992626,I524982,I992632,I525008,I525016,I992638,I992623,I525042,I525050,I525067,I525084,I525101,I992635,I525141,I525149,I525166,I525183,I525200,I525231,I992641,I992629,I525248,I525274,I525282,I525313,I525344,I525361,I525392,I525492,I525518,I525526,I525543,I525560,I525586,I525594,I525620,I525628,I525645,I525662,I525679,I525475,I525719,I525727,I525744,I525761,I525778,I525478,I525809,I525826,I525852,I525860,I525460,I525891,I525469,I525922,I525939,I525481,I525970,I525472,I525463,I525466,I525484,I526070,I526096,I526104,I526121,I526138,I526164,I526172,I526198,I526206,I526223,I526240,I526257,I526297,I526305,I526322,I526339,I526356,I526387,I526404,I526430,I526438,I526469,I526500,I526517,I526548,I526648,I526674,I526682,I526699,I526716,I526742,I526750,I526776,I526784,I526801,I526818,I526835,I526875,I526883,I526900,I526917,I526934,I526965,I526982,I527008,I527016,I527047,I527078,I527095,I527126,I527226,I527252,I527260,I527277,I527294,I527320,I527328,I527354,I527362,I527379,I527396,I527413,I527453,I527461,I527478,I527495,I527512,I527543,I527560,I527586,I527594,I527625,I527656,I527673,I527704,I527804,I698697,I527830,I527838,I527855,I698673,I698688,I527872,I698700,I527898,I527906,I698685,I698676,I527932,I527940,I527957,I527974,I527991,I527787,I528031,I528039,I528056,I528073,I528090,I527790,I528121,I698691,I698682,I528138,I698694,I528164,I528172,I527772,I528203,I527781,I528234,I528251,I527793,I528282,I698679,I527784,I527775,I527778,I527796,I528382,I929942,I528408,I528416,I528433,I929924,I929936,I528450,I929939,I528476,I528484,I929933,I929930,I528510,I528518,I528535,I528552,I528569,I528365,I929948,I528609,I528617,I528634,I528651,I528668,I528368,I528699,I929927,I528716,I528742,I528750,I528350,I528781,I528359,I528812,I528829,I528371,I528860,I929945,I528362,I528353,I528356,I528374,I528960,I749085,I528986,I528994,I529011,I749061,I749076,I529028,I749088,I529054,I529062,I749073,I749064,I529088,I529096,I529113,I529130,I529147,I529187,I529195,I529212,I529229,I529246,I529277,I749079,I749070,I529294,I749082,I529320,I529328,I529359,I529390,I529407,I529438,I749067,I529538,I529564,I529572,I529589,I529606,I529632,I529640,I529666,I529674,I529691,I529708,I529725,I529765,I529773,I529790,I529807,I529824,I529855,I529872,I529898,I529906,I529937,I529968,I529985,I530016,I530116,I920116,I530142,I530150,I530167,I920098,I920110,I530184,I920113,I530210,I530218,I920107,I920104,I530244,I530252,I530269,I530286,I530303,I530099,I920122,I530343,I530351,I530368,I530385,I530402,I530102,I530433,I920101,I530450,I530476,I530484,I530084,I530515,I530093,I530546,I530563,I530105,I530594,I920119,I530096,I530087,I530090,I530108,I530694,I530720,I530728,I530745,I530762,I530788,I530796,I530822,I530830,I530847,I530864,I530881,I530677,I530921,I530929,I530946,I530963,I530980,I530680,I531011,I531028,I531054,I531062,I530662,I531093,I530671,I531124,I531141,I530683,I531172,I530674,I530665,I530668,I530686,I531272,I531298,I531306,I531323,I531340,I531366,I531374,I531400,I531408,I531425,I531442,I531459,I531499,I531507,I531524,I531541,I531558,I531589,I531606,I531632,I531640,I531671,I531702,I531719,I531750,I531850,I780739,I531876,I531884,I531901,I780715,I780730,I531918,I780742,I531944,I531952,I780727,I780718,I531978,I531986,I532003,I532020,I532037,I532077,I532085,I532102,I532119,I532136,I532167,I780733,I780724,I532184,I780736,I532210,I532218,I532249,I532280,I532297,I532328,I780721,I532428,I780093,I532454,I532462,I532479,I780069,I780084,I532496,I780096,I532522,I532530,I780081,I780072,I532556,I532564,I532581,I532598,I532615,I532411,I532655,I532663,I532680,I532697,I532714,I532414,I532745,I780087,I780078,I532762,I780090,I532788,I532796,I532396,I532827,I532405,I532858,I532875,I532417,I532906,I780075,I532408,I532399,I532402,I532420,I533006,I836884,I533032,I533040,I533057,I836866,I836878,I533074,I836881,I533100,I533108,I836875,I836872,I533134,I533142,I533159,I533176,I533193,I532989,I836890,I533233,I533241,I533258,I533275,I533292,I532992,I533323,I836869,I533340,I533366,I533374,I532974,I533405,I532983,I533436,I533453,I532995,I533484,I836887,I532986,I532977,I532980,I532998,I533584,I875032,I533610,I533618,I533635,I875014,I875026,I533652,I875029,I533678,I533686,I875023,I875020,I533712,I533720,I533737,I533754,I533771,I875038,I533811,I533819,I533836,I533853,I533870,I533901,I875017,I533918,I533944,I533952,I533983,I534014,I534031,I534062,I875035,I534162,I534188,I534196,I534213,I534230,I534256,I534264,I534290,I534298,I534315,I534332,I534349,I534389,I534397,I534414,I534431,I534448,I534479,I534496,I534522,I534530,I534561,I534592,I534609,I534640,I534740,I686567,I534766,I534774,I534791,I686555,I686573,I534808,I686570,I534834,I534842,I686561,I686558,I534868,I534876,I534893,I534910,I534927,I534723,I686552,I534967,I534975,I534992,I535009,I535026,I534726,I535057,I535074,I535100,I535108,I534708,I535139,I534717,I535170,I535187,I534729,I535218,I686564,I534720,I534711,I534714,I534732,I535318,I535344,I535352,I535369,I535386,I535412,I535420,I535446,I535454,I535471,I535488,I535505,I535301,I535545,I535553,I535570,I535587,I535604,I535304,I535635,I535652,I535678,I535686,I535286,I535717,I535295,I535748,I535765,I535307,I535796,I535298,I535289,I535292,I535310,I535896,I961374,I535922,I535930,I535947,I961377,I961386,I535964,I961389,I535990,I535998,I961398,I961380,I536024,I536032,I536049,I536066,I536083,I536123,I536131,I536148,I536165,I536182,I536213,I961395,I536230,I961392,I536256,I536264,I536295,I536326,I536343,I536374,I961383,I536474,I536500,I536508,I536525,I536542,I536568,I536576,I536602,I536610,I536627,I536644,I536661,I536701,I536709,I536726,I536743,I536760,I536791,I536808,I536834,I536842,I536873,I536904,I536921,I536952,I537052,I1035266,I537078,I537086,I537103,I1035251,I1035239,I537120,I1035254,I537146,I537154,I1035257,I537180,I537188,I537205,I537222,I537239,I1035245,I537279,I537287,I537304,I537321,I537338,I537369,I1035242,I1035248,I537386,I1035263,I537412,I537420,I537451,I537482,I537499,I537530,I1035260,I537630,I537656,I537664,I537681,I537698,I537724,I537732,I537758,I537766,I537783,I537800,I537817,I537857,I537865,I537882,I537899,I537916,I537947,I537964,I537990,I537998,I538029,I538060,I538077,I538108,I538208,I538234,I538242,I538259,I538276,I538302,I538310,I538336,I538344,I538361,I538378,I538395,I538191,I538435,I538443,I538460,I538477,I538494,I538194,I538525,I538542,I538568,I538576,I538176,I538607,I538185,I538638,I538655,I538197,I538686,I538188,I538179,I538182,I538200,I538786,I538812,I538820,I538837,I538854,I538880,I538888,I538914,I538922,I538939,I538956,I538973,I539013,I539021,I539038,I539055,I539072,I539103,I539120,I539146,I539154,I539185,I539216,I539233,I539264,I539364,I539390,I539398,I539415,I539432,I539458,I539466,I539492,I539500,I539517,I539534,I539551,I539591,I539599,I539616,I539633,I539650,I539681,I539698,I539724,I539732,I539763,I539794,I539811,I539842,I539942,I539968,I539976,I539993,I540010,I540036,I540044,I540070,I540078,I540095,I540112,I540129,I539925,I540169,I540177,I540194,I540211,I540228,I539928,I540259,I540276,I540302,I540310,I539910,I540341,I539919,I540372,I540389,I539931,I540420,I539922,I539913,I539916,I539934,I540520,I668122,I540546,I540554,I540571,I668110,I668128,I540588,I668125,I540614,I540622,I668116,I668113,I540648,I540656,I540673,I540690,I540707,I540503,I668107,I540747,I540755,I540772,I540789,I540806,I540506,I540837,I540854,I540880,I540888,I540488,I540919,I540497,I540950,I540967,I540509,I540998,I668119,I540500,I540491,I540494,I540512,I541098,I541124,I541132,I541149,I541166,I541192,I541200,I541226,I541234,I541251,I541268,I541285,I541325,I541333,I541350,I541367,I541384,I541415,I541432,I541458,I541466,I541497,I541528,I541545,I541576,I541676,I672865,I541702,I541710,I541727,I672853,I672871,I541744,I672868,I541770,I541778,I672859,I672856,I541804,I541812,I541829,I541846,I541863,I672850,I541903,I541911,I541928,I541945,I541962,I541993,I542010,I542036,I542044,I542075,I542106,I542123,I542154,I672862,I542254,I542280,I542288,I542305,I542322,I542348,I542356,I542382,I542390,I542407,I542424,I542441,I542481,I542489,I542506,I542523,I542540,I542571,I542588,I542614,I542622,I542653,I542684,I542701,I542732,I542832,I1039431,I542858,I542866,I542883,I1039416,I1039404,I542900,I1039419,I542926,I542934,I1039422,I542960,I542968,I542985,I543002,I543019,I542815,I1039410,I543059,I543067,I543084,I543101,I543118,I542818,I543149,I1039407,I1039413,I543166,I1039428,I543192,I543200,I542800,I543231,I542809,I543262,I543279,I542821,I543310,I1039425,I542812,I542803,I542806,I542824,I543410,I543436,I543444,I543461,I543478,I543504,I543512,I543538,I543546,I543563,I543580,I543597,I543637,I543645,I543662,I543679,I543696,I543727,I543744,I543770,I543778,I543809,I543840,I543857,I543888,I543988,I633867,I544014,I544022,I544039,I633855,I633873,I544056,I633870,I544082,I544090,I633861,I633858,I544116,I544124,I544141,I544158,I544175,I543971,I633852,I544215,I544223,I544240,I544257,I544274,I543974,I544305,I544322,I544348,I544356,I543956,I544387,I543965,I544418,I544435,I543977,I544466,I633864,I543968,I543959,I543962,I543980,I544566,I1011116,I544592,I544600,I544617,I1011140,I1011122,I544634,I1011128,I544660,I544668,I1011134,I1011119,I544694,I544702,I544719,I544736,I544753,I1011131,I544793,I544801,I544818,I544835,I544852,I544883,I1011137,I1011125,I544900,I544926,I544934,I544965,I544996,I545013,I545044,I545144,I1084056,I545170,I545178,I545195,I1084041,I1084029,I545212,I1084044,I545238,I545246,I1084047,I545272,I545280,I545297,I545314,I545331,I1084035,I545371,I545379,I545396,I545413,I545430,I545461,I1084032,I1084038,I545478,I1084053,I545504,I545512,I545543,I545574,I545591,I545622,I1084050,I545722,I545748,I545756,I545773,I545790,I545816,I545824,I545850,I545858,I545875,I545892,I545909,I545705,I545949,I545957,I545974,I545991,I546008,I545708,I546039,I546056,I546082,I546090,I545690,I546121,I545699,I546152,I546169,I545711,I546200,I545702,I545693,I545696,I545714,I546300,I546326,I546334,I546351,I546368,I546394,I546402,I546428,I546436,I546453,I546470,I546487,I546283,I546527,I546535,I546552,I546569,I546586,I546286,I546617,I546634,I546660,I546668,I546268,I546699,I546277,I546730,I546747,I546289,I546778,I546280,I546271,I546274,I546292,I546878,I546904,I546912,I546929,I546946,I546972,I546980,I547006,I547014,I547031,I547048,I547065,I546861,I547105,I547113,I547130,I547147,I547164,I546864,I547195,I547212,I547238,I547246,I546846,I547277,I546855,I547308,I547325,I546867,I547356,I546858,I546849,I546852,I546870,I547456,I547482,I547490,I547507,I547524,I547550,I547558,I547584,I547592,I547609,I547626,I547643,I547439,I547683,I547691,I547708,I547725,I547742,I547442,I547773,I547790,I547816,I547824,I547424,I547855,I547433,I547886,I547903,I547445,I547934,I547436,I547427,I547430,I547448,I548034,I548060,I548068,I548085,I548102,I548128,I548136,I548162,I548170,I548187,I548204,I548221,I548261,I548269,I548286,I548303,I548320,I548351,I548368,I548394,I548402,I548433,I548464,I548481,I548512,I548612,I548638,I548646,I548663,I548680,I548706,I548714,I548740,I548748,I548765,I548782,I548799,I548839,I548847,I548864,I548881,I548898,I548929,I548946,I548972,I548980,I549011,I549042,I549059,I549090,I549190,I549216,I549224,I549241,I549258,I549284,I549292,I549318,I549326,I549343,I549360,I549377,I549173,I549417,I549425,I549442,I549459,I549476,I549176,I549507,I549524,I549550,I549558,I549158,I549589,I549167,I549620,I549637,I549179,I549668,I549170,I549161,I549164,I549182,I549768,I924162,I549794,I549802,I549819,I924144,I924156,I549836,I924159,I549862,I549870,I924153,I924150,I549896,I549904,I549921,I549938,I549955,I924168,I549995,I550003,I550020,I550037,I550054,I550085,I924147,I550102,I550128,I550136,I550167,I550198,I550215,I550246,I924165,I550346,I550372,I550380,I550397,I550414,I550440,I550448,I550474,I550482,I550499,I550516,I550533,I550329,I550573,I550581,I550598,I550615,I550632,I550332,I550663,I550680,I550706,I550714,I550314,I550745,I550323,I550776,I550793,I550335,I550824,I550326,I550317,I550320,I550338,I550924,I904510,I550950,I550958,I550975,I904492,I904504,I550992,I904507,I551018,I551026,I904501,I904498,I551052,I551060,I551077,I551094,I551111,I904516,I551151,I551159,I551176,I551193,I551210,I551241,I904495,I551258,I551284,I551292,I551323,I551354,I551371,I551402,I904513,I551502,I551528,I551536,I551553,I551570,I551596,I551604,I551630,I551638,I551655,I551672,I551689,I551485,I551729,I551737,I551754,I551771,I551788,I551488,I551819,I551836,I551862,I551870,I551470,I551901,I551479,I551932,I551949,I551491,I551980,I551482,I551473,I551476,I551494,I552080,I552106,I552114,I552131,I552148,I552174,I552182,I552208,I552216,I552233,I552250,I552267,I552063,I552307,I552315,I552332,I552349,I552366,I552066,I552397,I552414,I552440,I552448,I552048,I552479,I552057,I552510,I552527,I552069,I552558,I552060,I552051,I552054,I552072,I552658,I552684,I552692,I552709,I552726,I552752,I552760,I552786,I552794,I552811,I552828,I552845,I552885,I552893,I552910,I552927,I552944,I552975,I552992,I553018,I553026,I553057,I553088,I553105,I553136,I553236,I553262,I553270,I553287,I553304,I553330,I553338,I553364,I553372,I553389,I553406,I553423,I553219,I553463,I553471,I553488,I553505,I553522,I553222,I553553,I553570,I553596,I553604,I553204,I553635,I553213,I553666,I553683,I553225,I553714,I553216,I553207,I553210,I553228,I553814,I859426,I553840,I553848,I553865,I859408,I859420,I553882,I859423,I553908,I553916,I859417,I859414,I553942,I553950,I553967,I553984,I554001,I553797,I859432,I554041,I554049,I554066,I554083,I554100,I553800,I554131,I859411,I554148,I554174,I554182,I553782,I554213,I553791,I554244,I554261,I553803,I554292,I859429,I553794,I553785,I553788,I553806,I554392,I984222,I554418,I554426,I554443,I984225,I984234,I554460,I984237,I554486,I554494,I984246,I984228,I554520,I554528,I554545,I554562,I554579,I554619,I554627,I554644,I554661,I554678,I554709,I984243,I554726,I984240,I554752,I554760,I554791,I554822,I554839,I554870,I984231,I554970,I913180,I554996,I555004,I555021,I913162,I913174,I555038,I913177,I555064,I555072,I913171,I913168,I555098,I555106,I555123,I555140,I555157,I913186,I555197,I555205,I555222,I555239,I555256,I555287,I913165,I555304,I555330,I555338,I555369,I555400,I555417,I555448,I913183,I555548,I555574,I555582,I555599,I555616,I555642,I555650,I555676,I555684,I555701,I555718,I555735,I555531,I555775,I555783,I555800,I555817,I555834,I555534,I555865,I555882,I555908,I555916,I555516,I555947,I555525,I555978,I555995,I555537,I556026,I555528,I555519,I555522,I555540,I556126,I652839,I556152,I556160,I556177,I652827,I652845,I556194,I652842,I556220,I556228,I652833,I652830,I556254,I556262,I556279,I556296,I556313,I652824,I556353,I556361,I556378,I556395,I556412,I556443,I556460,I556486,I556494,I556525,I556556,I556573,I556604,I652836,I556704,I556730,I556738,I556755,I556772,I556798,I556806,I556832,I556840,I556857,I556874,I556891,I556931,I556939,I556956,I556973,I556990,I557021,I557038,I557064,I557072,I557103,I557134,I557151,I557182,I557282,I557308,I557316,I557333,I557350,I557376,I557384,I557410,I557418,I557435,I557452,I557469,I557509,I557517,I557534,I557551,I557568,I557599,I557616,I557642,I557650,I557681,I557712,I557729,I557760,I557860,I972798,I557886,I557894,I557911,I972801,I972810,I557928,I972813,I557954,I557962,I972822,I972804,I557988,I557996,I558013,I558030,I558047,I558087,I558095,I558112,I558129,I558146,I558177,I972819,I558194,I972816,I558220,I558228,I558259,I558290,I558307,I558338,I972807,I558438,I558464,I558472,I558489,I558506,I558532,I558540,I558566,I558574,I558591,I558608,I558625,I558421,I558665,I558673,I558690,I558707,I558724,I558424,I558755,I558772,I558798,I558806,I558406,I558837,I558415,I558868,I558885,I558427,I558916,I558418,I558409,I558412,I558430,I559016,I773633,I559042,I559050,I559067,I773609,I773624,I559084,I773636,I559110,I559118,I773621,I773612,I559144,I559152,I559169,I559186,I559203,I559243,I559251,I559268,I559285,I559302,I559333,I773627,I773618,I559350,I773630,I559376,I559384,I559415,I559446,I559463,I559494,I773615,I559594,I559620,I559628,I559645,I559662,I559688,I559696,I559722,I559730,I559747,I559764,I559781,I559577,I559821,I559829,I559846,I559863,I559880,I559580,I559911,I559928,I559954,I559962,I559562,I559993,I559571,I560024,I560041,I559583,I560072,I559574,I559565,I559568,I559586,I560172,I560198,I560206,I560223,I560240,I560266,I560274,I560300,I560308,I560325,I560342,I560359,I560399,I560407,I560424,I560441,I560458,I560489,I560506,I560532,I560540,I560571,I560602,I560619,I560650,I560750,I688675,I560776,I560784,I560801,I688663,I688681,I560818,I688678,I560844,I560852,I688669,I688666,I560878,I560886,I560903,I560920,I560937,I688660,I560977,I560985,I561002,I561019,I561036,I561067,I561084,I561110,I561118,I561149,I561180,I561197,I561228,I688672,I561328,I561354,I561362,I561379,I561396,I561422,I561430,I561456,I561464,I561481,I561498,I561515,I561311,I561555,I561563,I561580,I561597,I561614,I561314,I561645,I561662,I561688,I561696,I561296,I561727,I561305,I561758,I561775,I561317,I561806,I561308,I561299,I561302,I561320,I561906,I561932,I561940,I561957,I561974,I562000,I562008,I562034,I562042,I562059,I562076,I562093,I562133,I562141,I562158,I562175,I562192,I562223,I562240,I562266,I562274,I562305,I562336,I562353,I562384,I562484,I562510,I562518,I562535,I562552,I562578,I562586,I562612,I562620,I562637,I562654,I562671,I562467,I562711,I562719,I562736,I562753,I562770,I562470,I562801,I562818,I562844,I562852,I562452,I562883,I562461,I562914,I562931,I562473,I562962,I562464,I562455,I562458,I562476,I563062,I896996,I563088,I563096,I563113,I896978,I896990,I563130,I896993,I563156,I563164,I896987,I896984,I563190,I563198,I563215,I563232,I563249,I563045,I897002,I563289,I563297,I563314,I563331,I563348,I563048,I563379,I896981,I563396,I563422,I563430,I563030,I563461,I563039,I563492,I563509,I563051,I563540,I896999,I563042,I563033,I563036,I563054,I563640,I1017474,I563666,I563674,I563691,I1017498,I1017480,I563708,I1017486,I563734,I563742,I1017492,I1017477,I563768,I563776,I563793,I563810,I563827,I1017489,I563867,I563875,I563892,I563909,I563926,I563957,I1017495,I1017483,I563974,I564000,I564008,I564039,I564070,I564087,I564118,I564218,I819787,I564244,I564252,I564269,I819784,I819802,I564286,I819799,I564312,I564320,I819781,I564346,I564354,I564371,I564388,I564405,I819793,I564445,I564453,I564470,I564487,I564504,I564535,I819796,I564552,I564578,I564586,I564617,I564648,I564665,I564696,I819790,I564796,I564822,I564830,I564847,I564864,I564890,I564898,I564924,I564932,I564949,I564966,I564983,I564779,I565023,I565031,I565048,I565065,I565082,I564782,I565113,I565130,I565156,I565164,I564764,I565195,I564773,I565226,I565243,I564785,I565274,I564776,I564767,I564770,I564788,I565374,I565400,I565408,I565425,I565442,I565468,I565476,I565502,I565510,I565527,I565544,I565561,I565357,I565601,I565609,I565626,I565643,I565660,I565360,I565691,I565708,I565734,I565742,I565342,I565773,I565351,I565804,I565821,I565363,I565852,I565354,I565345,I565348,I565366,I565952,I666541,I565978,I565986,I566003,I666529,I666547,I566020,I666544,I566046,I566054,I666535,I666532,I566080,I566088,I566105,I566122,I566139,I666526,I566179,I566187,I566204,I566221,I566238,I566269,I566286,I566312,I566320,I566351,I566382,I566399,I566430,I666538,I566530,I566556,I566564,I566581,I566598,I566624,I566632,I566658,I566666,I566683,I566700,I566717,I566513,I566757,I566765,I566782,I566799,I566816,I566516,I566847,I566864,I566890,I566898,I566498,I566929,I566507,I566960,I566977,I566519,I567008,I566510,I566501,I566504,I566522,I567108,I567134,I567142,I567159,I567176,I567202,I567210,I567236,I567244,I567261,I567278,I567295,I567091,I567335,I567343,I567360,I567377,I567394,I567094,I567425,I567442,I567468,I567476,I567076,I567507,I567085,I567538,I567555,I567097,I567586,I567088,I567079,I567082,I567100,I567686,I989730,I567712,I567720,I567737,I989754,I989736,I567754,I989742,I567780,I567788,I989748,I989733,I567814,I567822,I567839,I567856,I567873,I989745,I567913,I567921,I567938,I567955,I567972,I568003,I989751,I989739,I568020,I568046,I568054,I568085,I568116,I568133,I568164,I568264,I716139,I568290,I568298,I568315,I716115,I716130,I568332,I716142,I568358,I568366,I716127,I716118,I568392,I568400,I568417,I568434,I568451,I568491,I568499,I568516,I568533,I568550,I568581,I716133,I716124,I568598,I716136,I568624,I568632,I568663,I568694,I568711,I568742,I716121,I568842,I568868,I568876,I568893,I568910,I568936,I568944,I568970,I568978,I568995,I569012,I569029,I568825,I569069,I569077,I569094,I569111,I569128,I568828,I569159,I569176,I569202,I569210,I568810,I569241,I568819,I569272,I569289,I568831,I569320,I568822,I568813,I568816,I568834,I569420,I569446,I569454,I569471,I569488,I569514,I569522,I569548,I569556,I569573,I569590,I569607,I569403,I569647,I569655,I569672,I569689,I569706,I569406,I569737,I569754,I569780,I569788,I569388,I569819,I569397,I569850,I569867,I569409,I569898,I569400,I569391,I569394,I569412,I569998,I570024,I570032,I570049,I570066,I570092,I570100,I570126,I570134,I570151,I570168,I570185,I569981,I570225,I570233,I570250,I570267,I570284,I569984,I570315,I570332,I570358,I570366,I569966,I570397,I569975,I570428,I570445,I569987,I570476,I569978,I569969,I569972,I569990,I570576,I570602,I570610,I570627,I570644,I570670,I570678,I570704,I570712,I570729,I570746,I570763,I570559,I570803,I570811,I570828,I570845,I570862,I570562,I570893,I570910,I570936,I570944,I570544,I570975,I570553,I571006,I571023,I570565,I571054,I570556,I570547,I570550,I570568,I571154,I630705,I571180,I571188,I571205,I630693,I630711,I571222,I630708,I571248,I571256,I630699,I630696,I571282,I571290,I571307,I571324,I571341,I571137,I630690,I571381,I571389,I571406,I571423,I571440,I571140,I571471,I571488,I571514,I571522,I571122,I571553,I571131,I571584,I571601,I571143,I571632,I630702,I571134,I571125,I571128,I571146,I571732,I1038836,I571758,I571766,I571783,I1038821,I1038809,I571800,I1038824,I571826,I571834,I1038827,I571860,I571868,I571885,I571902,I571919,I1038815,I571959,I571967,I571984,I572001,I572018,I572049,I1038812,I1038818,I572066,I1038833,I572092,I572100,I572131,I572162,I572179,I572210,I1038830,I572310,I881390,I572336,I572344,I572361,I881372,I881384,I572378,I881387,I572404,I572412,I881381,I881378,I572438,I572446,I572463,I572480,I572497,I572293,I881396,I572537,I572545,I572562,I572579,I572596,I572296,I572627,I881375,I572644,I572670,I572678,I572278,I572709,I572287,I572740,I572757,I572299,I572788,I881393,I572290,I572281,I572284,I572302,I572888,I572914,I572922,I572939,I572956,I572982,I572990,I573016,I573024,I573041,I573058,I573075,I572871,I573115,I573123,I573140,I573157,I573174,I572874,I573205,I573222,I573248,I573256,I572856,I573287,I572865,I573318,I573335,I572877,I573366,I572868,I572859,I572862,I572880,I573466,I573492,I573500,I573517,I573534,I573560,I573568,I573594,I573602,I573619,I573636,I573653,I573693,I573701,I573718,I573735,I573752,I573783,I573800,I573826,I573834,I573865,I573896,I573913,I573944,I574044,I686040,I574070,I574078,I574095,I686028,I686046,I574112,I686043,I574138,I574146,I686034,I686031,I574172,I574180,I574197,I574214,I574231,I686025,I574271,I574279,I574296,I574313,I574330,I574361,I574378,I574404,I574412,I574443,I574474,I574491,I574522,I686037,I574622,I716785,I574648,I574656,I574673,I716761,I716776,I574690,I716788,I574716,I574724,I716773,I716764,I574750,I574758,I574775,I574792,I574809,I574605,I574849,I574857,I574874,I574891,I574908,I574608,I574939,I716779,I716770,I574956,I716782,I574982,I574990,I574590,I575021,I574599,I575052,I575069,I574611,I575100,I716767,I574602,I574593,I574596,I574614,I575200,I575226,I575234,I575251,I575268,I575294,I575302,I575328,I575336,I575353,I575370,I575387,I575427,I575435,I575452,I575469,I575486,I575517,I575534,I575560,I575568,I575599,I575630,I575647,I575678,I575778,I883124,I575804,I575812,I575829,I883106,I883118,I575846,I883121,I575872,I575880,I883115,I883112,I575906,I575914,I575931,I575948,I575965,I575761,I883130,I576005,I576013,I576030,I576047,I576064,I575764,I576095,I883109,I576112,I576138,I576146,I575746,I576177,I575755,I576208,I576225,I575767,I576256,I883127,I575758,I575749,I575752,I575770,I576356,I1012850,I576382,I576390,I576407,I1012874,I1012856,I576424,I1012862,I576450,I576458,I1012868,I1012853,I576484,I576492,I576509,I576526,I576543,I576339,I1012865,I576583,I576591,I576608,I576625,I576642,I576342,I576673,I1012871,I1012859,I576690,I576716,I576724,I576324,I576755,I576333,I576786,I576803,I576345,I576834,I576336,I576327,I576330,I576348,I576934,I1072156,I576960,I576968,I576985,I1072141,I1072129,I577002,I1072144,I577028,I577036,I1072147,I577062,I577070,I577087,I577104,I577121,I576917,I1072135,I577161,I577169,I577186,I577203,I577220,I576920,I577251,I1072132,I1072138,I577268,I1072153,I577294,I577302,I576902,I577333,I576911,I577364,I577381,I576923,I577412,I1072150,I576914,I576905,I576908,I576926,I577512,I577538,I577546,I577563,I577580,I577606,I577614,I577640,I577648,I577665,I577682,I577699,I577739,I577747,I577764,I577781,I577798,I577829,I577846,I577872,I577880,I577911,I577942,I577959,I577990,I578090,I578116,I578124,I578141,I578158,I578184,I578192,I578218,I578226,I578243,I578260,I578277,I578073,I578317,I578325,I578342,I578359,I578376,I578076,I578407,I578424,I578450,I578458,I578058,I578489,I578067,I578520,I578537,I578079,I578568,I578070,I578061,I578064,I578082,I578668,I578694,I578702,I578719,I578736,I578762,I578770,I578796,I578804,I578821,I578838,I578855,I578895,I578903,I578920,I578937,I578954,I578985,I579002,I579028,I579036,I579067,I579098,I579115,I579146,I579246,I957566,I579272,I579280,I579297,I957569,I957578,I579314,I957581,I579340,I579348,I957590,I957572,I579374,I579382,I579399,I579416,I579433,I579473,I579481,I579498,I579515,I579532,I579563,I957587,I579580,I957584,I579606,I579614,I579645,I579676,I579693,I579724,I957575,I579824,I934566,I579850,I579858,I579875,I934548,I934560,I579892,I934563,I579918,I579926,I934557,I934554,I579952,I579960,I579977,I579994,I580011,I934572,I580051,I580059,I580076,I580093,I580110,I580141,I934551,I580158,I580184,I580192,I580223,I580254,I580271,I580302,I934569,I580402,I580428,I580436,I580453,I580470,I580496,I580504,I580530,I580538,I580555,I580572,I580589,I580385,I580629,I580637,I580654,I580671,I580688,I580388,I580719,I580736,I580762,I580770,I580370,I580801,I580379,I580832,I580849,I580391,I580880,I580382,I580373,I580376,I580394,I580980,I629651,I581006,I581014,I581031,I629639,I629657,I581048,I629654,I581074,I581082,I629645,I629642,I581108,I581116,I581133,I581150,I581167,I580963,I629636,I581207,I581215,I581232,I581249,I581266,I580966,I581297,I581314,I581340,I581348,I580948,I581379,I580957,I581410,I581427,I580969,I581458,I629648,I580960,I580951,I580954,I580972,I581558,I581584,I581592,I581609,I581626,I581652,I581660,I581686,I581694,I581711,I581728,I581745,I581541,I581785,I581793,I581810,I581827,I581844,I581544,I581875,I581892,I581918,I581926,I581526,I581957,I581535,I581988,I582005,I581547,I582036,I581538,I581529,I581532,I581550,I582136,I582162,I582170,I582187,I582204,I582230,I582238,I582264,I582272,I582289,I582306,I582323,I582363,I582371,I582388,I582405,I582422,I582453,I582470,I582496,I582504,I582535,I582566,I582583,I582614,I582714,I582740,I582748,I582765,I582782,I582808,I582816,I582842,I582850,I582867,I582884,I582901,I582697,I582941,I582949,I582966,I582983,I583000,I582700,I583031,I583048,I583074,I583082,I582682,I583113,I582691,I583144,I583161,I582703,I583192,I582694,I582685,I582688,I582706,I583292,I583318,I583326,I583343,I583360,I583386,I583394,I583420,I583428,I583445,I583462,I583479,I583519,I583527,I583544,I583561,I583578,I583609,I583626,I583652,I583660,I583691,I583722,I583739,I583770,I583870,I583896,I583904,I583921,I583938,I583964,I583972,I583998,I584006,I584023,I584040,I584057,I584097,I584105,I584122,I584139,I584156,I584187,I584204,I584230,I584238,I584269,I584300,I584317,I584348,I584448,I627543,I584474,I584482,I584499,I627531,I627549,I584516,I627546,I584542,I584550,I627537,I627534,I584576,I584584,I584601,I584618,I584635,I627528,I584675,I584683,I584700,I584717,I584734,I584765,I584782,I584808,I584816,I584847,I584878,I584895,I584926,I627540,I585026,I585052,I585060,I585077,I585094,I585120,I585128,I585154,I585162,I585179,I585196,I585213,I585253,I585261,I585278,I585295,I585312,I585343,I585360,I585386,I585394,I585425,I585456,I585473,I585504,I585604,I585630,I585638,I585655,I585672,I585698,I585706,I585732,I585740,I585757,I585774,I585791,I585587,I585831,I585839,I585856,I585873,I585890,I585590,I585921,I585938,I585964,I585972,I585572,I586003,I585581,I586034,I586051,I585593,I586082,I585584,I585575,I585578,I585596,I586182,I623854,I586208,I586216,I586233,I623842,I623860,I586250,I623857,I586276,I586284,I623848,I623845,I586310,I586318,I586335,I586352,I586369,I623839,I586409,I586417,I586434,I586451,I586468,I586499,I586516,I586542,I586550,I586581,I586612,I586629,I586660,I623851,I586760,I759421,I586786,I586794,I586811,I759397,I759412,I586828,I759424,I586854,I586862,I759409,I759400,I586888,I586896,I586913,I586930,I586947,I586987,I586995,I587012,I587029,I587046,I587077,I759415,I759406,I587094,I759418,I587120,I587128,I587159,I587190,I587207,I587238,I759403,I587338,I587364,I587372,I587389,I587406,I587432,I587440,I587466,I587474,I587491,I587508,I587525,I587565,I587573,I587590,I587607,I587624,I587655,I587672,I587698,I587706,I587737,I587768,I587785,I587816,I587916,I587942,I587950,I587967,I587984,I588010,I588018,I588044,I588052,I588069,I588086,I588103,I588143,I588151,I588168,I588185,I588202,I588233,I588250,I588276,I588284,I588315,I588346,I588363,I588394,I588494,I588520,I588528,I588545,I588562,I588588,I588596,I588622,I588630,I588647,I588664,I588681,I588477,I588721,I588729,I588746,I588763,I588780,I588480,I588811,I588828,I588854,I588862,I588462,I588893,I588471,I588924,I588941,I588483,I588972,I588474,I588465,I588468,I588486,I589072,I883702,I589098,I589106,I589123,I883684,I883696,I589140,I883699,I589166,I589174,I883693,I883690,I589200,I589208,I589225,I589242,I589259,I589055,I883708,I589299,I589307,I589324,I589341,I589358,I589058,I589389,I883687,I589406,I589432,I589440,I589040,I589471,I589049,I589502,I589519,I589061,I589550,I883705,I589052,I589043,I589046,I589064,I589650,I746501,I589676,I589684,I589701,I746477,I746492,I589718,I746504,I589744,I589752,I746489,I746480,I589778,I589786,I589803,I589820,I589837,I589877,I589885,I589902,I589919,I589936,I589967,I746495,I746486,I589984,I746498,I590010,I590018,I590049,I590080,I590097,I590128,I746483,I590228,I590254,I590262,I590279,I590296,I590322,I590330,I590356,I590364,I590381,I590398,I590415,I590455,I590463,I590480,I590497,I590514,I590545,I590562,I590588,I590596,I590627,I590658,I590675,I590706,I590806,I849022,I590832,I590840,I590857,I849004,I849016,I590874,I849019,I590900,I590908,I849013,I849010,I590934,I590942,I590959,I590976,I590993,I590789,I849028,I591033,I591041,I591058,I591075,I591092,I590792,I591123,I849007,I591140,I591166,I591174,I590774,I591205,I590783,I591236,I591253,I590795,I591284,I849025,I590786,I590777,I590780,I590798,I591384,I993198,I591410,I591418,I591435,I993222,I993204,I591452,I993210,I591478,I591486,I993216,I993201,I591512,I591520,I591537,I591554,I591571,I591367,I993213,I591611,I591619,I591636,I591653,I591670,I591370,I591701,I993219,I993207,I591718,I591744,I591752,I591352,I591783,I591361,I591814,I591831,I591373,I591862,I591364,I591355,I591358,I591376,I591962,I879078,I591988,I591996,I592013,I879060,I879072,I592030,I879075,I592056,I592064,I879069,I879066,I592090,I592098,I592115,I592132,I592149,I591945,I879084,I592189,I592197,I592214,I592231,I592248,I591948,I592279,I879063,I592296,I592322,I592330,I591930,I592361,I591939,I592392,I592409,I591951,I592440,I879081,I591942,I591933,I591936,I591954,I592540,I592566,I592574,I592591,I592608,I592634,I592642,I592668,I592676,I592693,I592710,I592727,I592767,I592775,I592792,I592809,I592826,I592857,I592874,I592900,I592908,I592939,I592970,I592987,I593018,I593118,I593144,I593152,I593169,I593186,I593212,I593220,I593246,I593254,I593271,I593288,I593305,I593101,I593345,I593353,I593370,I593387,I593404,I593104,I593435,I593452,I593478,I593486,I593086,I593517,I593095,I593548,I593565,I593107,I593596,I593098,I593089,I593092,I593110,I593696,I990308,I593722,I593730,I593747,I990332,I990314,I593764,I990320,I593790,I593798,I990326,I990311,I593824,I593832,I593849,I593866,I593883,I593679,I990323,I593923,I593931,I593948,I593965,I593982,I593682,I594013,I990329,I990317,I594030,I594056,I594064,I593664,I594095,I593673,I594126,I594143,I593685,I594174,I593676,I593667,I593670,I593688,I594274,I594300,I594308,I594325,I594342,I594368,I594376,I594402,I594410,I594427,I594444,I594461,I594501,I594509,I594526,I594543,I594560,I594591,I594608,I594634,I594642,I594673,I594704,I594721,I594752,I594852,I594878,I594886,I594903,I594920,I594946,I594954,I594980,I594988,I595005,I595022,I595039,I595079,I595087,I595104,I595121,I595138,I595169,I595186,I595212,I595220,I595251,I595282,I595299,I595330,I595430,I595456,I595464,I595481,I595498,I595524,I595532,I595558,I595566,I595583,I595600,I595617,I595657,I595665,I595682,I595699,I595716,I595747,I595764,I595790,I595798,I595829,I595860,I595877,I595908,I596008,I648623,I596034,I596042,I596059,I648611,I648629,I596076,I648626,I596102,I596110,I648617,I648614,I596136,I596144,I596161,I596178,I596195,I595991,I648608,I596235,I596243,I596260,I596277,I596294,I595994,I596325,I596342,I596368,I596376,I595976,I596407,I595985,I596438,I596455,I595997,I596486,I648620,I595988,I595979,I595982,I596000,I596586,I596612,I596620,I596637,I596654,I596680,I596688,I596714,I596722,I596739,I596756,I596773,I596569,I596813,I596821,I596838,I596855,I596872,I596572,I596903,I596920,I596946,I596954,I596554,I596985,I596563,I597016,I597033,I596575,I597064,I596566,I596557,I596560,I596578,I597164,I683932,I597190,I597198,I597215,I683920,I683938,I597232,I683935,I597258,I597266,I683926,I683923,I597292,I597300,I597317,I597334,I597351,I597147,I683917,I597391,I597399,I597416,I597433,I597450,I597150,I597481,I597498,I597524,I597532,I597132,I597563,I597141,I597594,I597611,I597153,I597642,I683929,I597144,I597135,I597138,I597156,I597742,I835728,I597768,I597776,I597793,I835710,I835722,I597810,I835725,I597836,I597844,I835719,I835716,I597870,I597878,I597895,I597912,I597929,I835734,I597969,I597977,I597994,I598011,I598028,I598059,I835713,I598076,I598102,I598110,I598141,I598172,I598189,I598220,I835731,I598320,I598346,I598354,I598371,I598388,I598414,I598422,I598448,I598456,I598473,I598490,I598507,I598303,I598547,I598555,I598572,I598589,I598606,I598306,I598637,I598654,I598680,I598688,I598288,I598719,I598297,I598750,I598767,I598309,I598798,I598300,I598291,I598294,I598312,I598898,I598924,I598932,I598949,I598966,I598992,I599000,I599026,I599034,I599051,I599068,I599085,I599125,I599133,I599150,I599167,I599184,I599215,I599232,I599258,I599266,I599297,I599328,I599345,I599376,I599476,I599502,I599510,I599527,I599544,I599570,I599578,I599604,I599612,I599629,I599646,I599663,I599703,I599711,I599728,I599745,I599762,I599793,I599810,I599836,I599844,I599875,I599906,I599923,I599954,I600054,I600080,I600088,I600105,I600122,I600148,I600156,I600182,I600190,I600207,I600224,I600241,I600281,I600289,I600306,I600323,I600340,I600371,I600388,I600414,I600422,I600453,I600484,I600501,I600532,I600632,I731643,I600658,I600666,I600683,I731619,I731634,I600700,I731646,I600726,I600734,I731631,I731622,I600760,I600768,I600785,I600802,I600819,I600859,I600867,I600884,I600901,I600918,I600949,I731637,I731628,I600966,I731640,I600992,I601000,I601031,I601062,I601079,I601110,I731625,I601210,I601236,I601244,I601261,I601278,I601304,I601312,I601338,I601346,I601363,I601380,I601397,I601437,I601445,I601462,I601479,I601496,I601527,I601544,I601570,I601578,I601609,I601640,I601657,I601688,I601788,I601814,I601822,I601839,I601856,I601882,I601890,I601916,I601924,I601941,I601958,I601975,I601771,I602015,I602023,I602040,I602057,I602074,I601774,I602105,I602122,I602148,I602156,I601756,I602187,I601765,I602218,I602235,I601777,I602266,I601768,I601759,I601762,I601780,I602366,I602392,I602400,I602417,I602434,I602460,I602468,I602494,I602502,I602519,I602536,I602553,I602593,I602601,I602618,I602635,I602652,I602683,I602700,I602726,I602734,I602765,I602796,I602813,I602844,I602944,I783323,I602970,I602978,I602995,I783299,I783314,I603012,I783326,I603038,I603046,I783311,I783302,I603072,I603080,I603097,I603114,I603131,I603171,I603179,I603196,I603213,I603230,I603261,I783317,I783308,I603278,I783320,I603304,I603312,I603343,I603374,I603391,I603422,I783305,I603522,I603548,I603556,I603573,I603590,I603616,I603624,I603650,I603658,I603675,I603692,I603709,I603749,I603757,I603774,I603791,I603808,I603839,I603856,I603882,I603890,I603921,I603952,I603969,I604000,I604100,I747147,I604126,I604134,I604151,I747123,I747138,I604168,I747150,I604194,I604202,I747135,I747126,I604228,I604236,I604253,I604270,I604287,I604083,I604327,I604335,I604352,I604369,I604386,I604086,I604417,I747141,I747132,I604434,I747144,I604460,I604468,I604068,I604499,I604077,I604530,I604547,I604089,I604578,I747129,I604080,I604071,I604074,I604092,I604678,I604704,I604712,I604729,I604746,I604772,I604780,I604806,I604814,I604831,I604848,I604865,I604905,I604913,I604930,I604947,I604964,I604995,I605012,I605038,I605046,I605077,I605108,I605125,I605156,I605256,I694472,I605282,I605290,I605307,I694460,I694478,I605324,I694475,I605350,I605358,I694466,I694463,I605384,I605392,I605409,I605426,I605443,I694457,I605483,I605491,I605508,I605525,I605542,I605573,I605590,I605616,I605624,I605655,I605686,I605703,I605734,I694469,I605834,I605860,I605868,I605885,I605902,I605928,I605936,I605962,I605970,I605987,I606004,I606021,I606061,I606069,I606086,I606103,I606120,I606151,I606168,I606194,I606202,I606233,I606264,I606281,I606312,I606412,I606438,I606446,I606463,I606480,I606506,I606514,I606540,I606548,I606565,I606582,I606599,I606639,I606647,I606664,I606681,I606698,I606729,I606746,I606772,I606780,I606811,I606842,I606859,I606890,I606990,I813055,I607016,I607024,I607041,I813052,I813070,I607058,I813067,I607084,I607092,I813049,I607118,I607126,I607143,I607160,I607177,I606973,I813061,I607217,I607225,I607242,I607259,I607276,I606976,I607307,I813064,I607324,I607350,I607358,I606958,I607389,I606967,I607420,I607437,I606979,I607468,I813058,I606970,I606961,I606964,I606982,I607568,I607594,I607602,I607619,I607636,I607662,I607670,I607696,I607704,I607721,I607738,I607755,I607795,I607803,I607820,I607837,I607854,I607885,I607902,I607928,I607936,I607967,I607998,I608015,I608046,I608146,I712909,I608172,I608180,I608197,I712885,I712900,I608214,I712912,I608240,I608248,I712897,I712888,I608274,I608282,I608299,I608316,I608333,I608373,I608381,I608398,I608415,I608432,I608463,I712903,I712894,I608480,I712906,I608506,I608514,I608545,I608576,I608593,I608624,I712891,I608724,I608750,I608758,I608775,I608792,I608818,I608826,I608852,I608860,I608877,I608894,I608911,I608707,I608951,I608959,I608976,I608993,I609010,I608710,I609041,I609058,I609084,I609092,I608692,I609123,I608701,I609154,I609171,I608713,I609202,I608704,I608695,I608698,I608716,I609302,I1059066,I609328,I609336,I609353,I1059051,I1059039,I609370,I1059054,I609396,I609404,I1059057,I609430,I609438,I609455,I609472,I609489,I609285,I1059045,I609529,I609537,I609554,I609571,I609588,I609288,I609619,I1059042,I1059048,I609636,I1059063,I609662,I609670,I609270,I609701,I609279,I609732,I609749,I609291,I609780,I1059060,I609282,I609273,I609276,I609294,I609880,I1082866,I609906,I609914,I609931,I1082851,I1082839,I609948,I1082854,I609974,I609982,I1082857,I610008,I610016,I610033,I610050,I610067,I609863,I1082845,I610107,I610115,I610132,I610149,I610166,I609866,I610197,I1082842,I1082848,I610214,I1082863,I610240,I610248,I609848,I610279,I609857,I610310,I610327,I609869,I610358,I1082860,I609860,I609851,I609854,I609872,I610458,I725183,I610484,I610492,I610509,I725159,I725174,I610526,I725186,I610552,I610560,I725171,I725162,I610586,I610594,I610611,I610628,I610645,I610685,I610693,I610710,I610727,I610744,I610775,I725177,I725168,I610792,I725180,I610818,I610826,I610857,I610888,I610905,I610936,I725165,I611036,I611062,I611070,I611087,I611104,I611130,I611138,I611164,I611172,I611189,I611206,I611223,I611263,I611271,I611288,I611305,I611322,I611353,I611370,I611396,I611404,I611435,I611466,I611483,I611514,I611614,I855958,I611640,I611648,I611665,I855940,I855952,I611682,I855955,I611708,I611716,I855949,I855946,I611742,I611750,I611767,I611784,I611801,I611597,I855964,I611841,I611849,I611866,I611883,I611900,I611600,I611931,I855943,I611948,I611974,I611982,I611582,I612013,I611591,I612044,I612061,I611603,I612092,I855961,I611594,I611585,I611588,I611606,I612192,I612218,I612226,I612243,I612260,I612286,I612294,I612320,I612328,I612345,I612362,I612379,I612175,I612419,I612427,I612444,I612461,I612478,I612178,I612509,I612526,I612552,I612560,I612160,I612591,I612169,I612622,I612639,I612181,I612670,I612172,I612163,I612166,I612184,I612770,I612796,I612804,I612821,I612838,I612864,I612872,I612898,I612906,I612923,I612940,I612957,I612753,I612997,I613005,I613022,I613039,I613056,I612756,I613087,I613104,I613130,I613138,I612738,I613169,I612747,I613200,I613217,I612759,I613248,I612750,I612741,I612744,I612762,I613348,I691310,I613374,I613382,I613399,I691298,I691316,I613416,I691313,I613442,I613450,I691304,I691301,I613476,I613484,I613501,I613518,I613535,I691295,I613575,I613583,I613600,I613617,I613634,I613665,I613682,I613708,I613716,I613747,I613778,I613795,I613826,I691307,I613926,I854802,I613952,I613960,I613977,I854784,I854796,I613994,I854799,I614020,I614028,I854793,I854790,I614054,I614062,I614079,I614096,I614113,I854808,I614153,I614161,I614178,I614195,I614212,I614243,I854787,I614260,I614286,I614294,I614325,I614356,I614373,I614404,I854805,I614504,I1076321,I614530,I614538,I614555,I1076306,I1076294,I614572,I1076309,I614598,I614606,I1076312,I614632,I614640,I614657,I614674,I614691,I614487,I1076300,I614731,I614739,I614756,I614773,I614790,I614490,I614821,I1076297,I1076303,I614838,I1076318,I614864,I614872,I614472,I614903,I614481,I614934,I614951,I614493,I614982,I1076315,I614484,I614475,I614478,I614496,I615082,I615108,I615116,I615133,I615150,I615176,I615184,I615210,I615218,I615235,I615252,I615269,I615309,I615317,I615334,I615351,I615368,I615399,I615416,I615442,I615450,I615481,I615512,I615529,I615560,I615660,I615686,I615694,I615711,I615728,I615754,I615762,I615788,I615796,I615813,I615830,I615847,I615887,I615895,I615912,I615929,I615946,I615977,I615994,I616020,I616028,I616059,I616090,I616107,I616138,I616238,I1098336,I616264,I616272,I616289,I1098321,I1098309,I616306,I1098324,I616332,I616340,I1098327,I616366,I616374,I616391,I616408,I616425,I616221,I1098315,I616465,I616473,I616490,I616507,I616524,I616224,I616555,I1098312,I1098318,I616572,I1098333,I616598,I616606,I616206,I616637,I616215,I616668,I616685,I616227,I616716,I1098330,I616218,I616209,I616212,I616230,I616816,I616842,I616850,I616867,I616884,I616910,I616918,I616944,I616952,I616969,I616986,I617003,I616799,I617043,I617051,I617068,I617085,I617102,I616802,I617133,I617150,I617176,I617184,I616784,I617215,I616793,I617246,I617263,I616805,I617294,I616796,I616787,I616790,I616808,I617394,I832260,I617420,I617428,I617445,I832242,I832254,I617462,I832257,I617488,I617496,I832251,I832248,I617522,I617530,I617547,I617564,I617581,I832266,I617621,I617629,I617646,I617663,I617680,I617711,I832245,I617728,I617754,I617762,I617793,I617824,I617841,I617872,I832263,I617972,I617998,I618006,I618023,I618040,I618066,I618074,I618100,I618108,I618125,I618142,I618159,I617955,I618199,I618207,I618224,I618241,I618258,I617958,I618289,I618306,I618332,I618340,I617940,I618371,I617949,I618402,I618419,I617961,I618450,I617952,I617943,I617946,I617964,I618550,I985310,I618576,I618584,I618601,I985313,I985322,I618618,I985325,I618644,I618652,I985334,I985316,I618678,I618686,I618703,I618720,I618737,I618533,I618777,I618785,I618802,I618819,I618836,I618536,I618867,I985331,I618884,I985328,I618910,I618918,I618518,I618949,I618527,I618980,I618997,I618539,I619028,I985319,I618530,I618521,I618524,I618542,I619125,I1075714,I619151,I619159,I619176,I1075711,I1075720,I619193,I1075699,I619219,I619114,I1075702,I619250,I619258,I1075717,I619275,I619301,I619309,I619117,I1075723,I619349,I619108,I619099,I619385,I1075705,I1075726,I619402,I1075708,I619428,I619436,I619453,I619102,I619484,I619501,I619518,I619111,I619549,I619096,I619580,I619597,I619105,I619652,I619678,I619686,I619703,I619720,I619746,I619777,I619785,I619802,I619828,I619836,I619876,I619912,I619929,I619955,I619963,I619980,I620011,I620028,I620045,I620076,I620107,I620124,I620179,I1090589,I620205,I620213,I620230,I1090586,I1090595,I620247,I1090574,I620273,I620168,I1090577,I620304,I620312,I1090592,I620329,I620355,I620363,I620171,I1090598,I620403,I620162,I620153,I620439,I1090580,I1090601,I620456,I1090583,I620482,I620490,I620507,I620156,I620538,I620555,I620572,I620165,I620603,I620150,I620634,I620651,I620159,I620706,I1053699,I620732,I620740,I620757,I1053696,I1053705,I620774,I1053684,I620800,I1053687,I620831,I620839,I1053702,I620856,I620882,I620890,I1053708,I620930,I620966,I1053690,I1053711,I620983,I1053693,I621009,I621017,I621034,I621065,I621082,I621099,I621130,I621161,I621178,I621233,I621259,I621267,I621284,I621301,I621327,I621358,I621366,I621383,I621409,I621417,I621457,I621493,I621510,I621536,I621544,I621561,I621592,I621609,I621626,I621657,I621688,I621705,I621760,I917226,I621786,I621794,I621811,I917208,I621828,I917214,I621854,I621749,I917211,I621885,I621893,I917220,I621910,I621936,I621944,I621752,I917232,I621984,I621743,I621734,I622020,I917223,I917217,I622037,I622063,I622071,I622088,I621737,I622119,I917229,I622136,I622153,I621746,I622184,I621731,I622215,I622232,I621740,I622287,I912602,I622313,I622321,I622338,I912584,I622355,I912590,I622381,I622276,I912587,I622412,I622420,I912596,I622437,I622463,I622471,I622279,I912608,I622511,I622270,I622261,I622547,I912599,I912593,I622564,I622590,I622598,I622615,I622264,I622646,I912605,I622663,I622680,I622273,I622711,I622258,I622742,I622759,I622267,I622814,I982058,I622840,I622848,I622865,I982064,I982046,I622882,I982055,I622908,I982061,I622939,I622947,I982049,I622964,I622990,I622998,I982067,I623038,I623074,I982052,I623091,I982070,I623117,I623125,I623142,I623173,I623190,I623207,I623238,I623269,I623286,I623341,I623367,I623375,I623392,I623409,I623435,I623330,I623466,I623474,I623491,I623517,I623525,I623333,I623565,I623324,I623315,I623601,I623618,I623644,I623652,I623669,I623318,I623700,I623717,I623734,I623327,I623765,I623312,I623796,I623813,I623321,I623868,I623894,I623902,I623919,I623936,I623962,I623993,I624001,I624018,I624044,I624052,I624092,I624128,I624145,I624171,I624179,I624196,I624227,I624244,I624261,I624292,I624323,I624340,I624395,I624421,I624429,I624446,I624463,I624489,I624384,I624520,I624528,I624545,I624571,I624579,I624387,I624619,I624378,I624369,I624655,I624672,I624698,I624706,I624723,I624372,I624754,I624771,I624788,I624381,I624819,I624366,I624850,I624867,I624375,I624922,I624948,I624956,I624973,I624990,I625016,I624911,I625047,I625055,I625072,I625098,I625106,I624914,I625146,I624905,I624896,I625182,I625199,I625225,I625233,I625250,I624899,I625281,I625298,I625315,I624908,I625346,I624893,I625377,I625394,I624902,I625449,I625475,I625483,I625500,I625517,I625543,I625574,I625582,I625599,I625625,I625633,I625673,I625709,I625726,I625752,I625760,I625777,I625808,I625825,I625842,I625873,I625904,I625921,I625976,I626002,I626010,I626027,I626044,I626070,I625965,I626101,I626109,I626126,I626152,I626160,I625968,I626200,I625959,I625950,I626236,I626253,I626279,I626287,I626304,I625953,I626335,I626352,I626369,I625962,I626400,I625947,I626431,I626448,I625956,I626503,I626529,I626537,I626554,I626571,I626597,I626628,I626636,I626653,I626679,I626687,I626727,I626763,I626780,I626806,I626814,I626831,I626862,I626879,I626896,I626927,I626958,I626975,I627030,I1099514,I627056,I627064,I627081,I1099511,I1099520,I627098,I1099499,I627124,I627019,I1099502,I627155,I627163,I1099517,I627180,I627206,I627214,I627022,I1099523,I627254,I627013,I627004,I627290,I1099505,I1099526,I627307,I1099508,I627333,I627341,I627358,I627007,I627389,I627406,I627423,I627016,I627454,I627001,I627485,I627502,I627010,I627557,I953640,I627583,I627591,I627608,I953622,I627625,I953628,I627651,I953625,I627682,I627690,I953634,I627707,I627733,I627741,I953646,I627781,I627817,I953637,I953631,I627834,I627860,I627868,I627885,I627916,I953643,I627933,I627950,I627981,I628012,I628029,I628084,I628110,I628118,I628135,I628152,I628178,I628073,I628209,I628217,I628234,I628260,I628268,I628076,I628308,I628067,I628058,I628344,I628361,I628387,I628395,I628412,I628061,I628443,I628460,I628477,I628070,I628508,I628055,I628539,I628556,I628064,I628611,I628637,I628645,I628662,I628679,I628705,I628736,I628744,I628761,I628787,I628795,I628835,I628871,I628888,I628914,I628922,I628939,I628970,I628987,I629004,I629035,I629066,I629083,I629138,I629164,I629172,I629189,I629206,I629232,I629263,I629271,I629288,I629314,I629322,I629362,I629398,I629415,I629441,I629449,I629466,I629497,I629514,I629531,I629562,I629593,I629610,I629665,I629691,I629699,I629716,I629733,I629759,I629790,I629798,I629815,I629841,I629849,I629889,I629925,I629942,I629968,I629976,I629993,I630024,I630041,I630058,I630089,I630120,I630137,I630192,I978250,I630218,I630226,I630243,I978256,I978238,I630260,I978247,I630286,I978253,I630317,I630325,I978241,I630342,I630368,I630376,I978259,I630416,I630452,I978244,I630469,I978262,I630495,I630503,I630520,I630551,I630568,I630585,I630616,I630647,I630664,I630719,I1068574,I630745,I630753,I630770,I1068571,I1068580,I630787,I1068559,I630813,I1068562,I630844,I630852,I1068577,I630869,I630895,I630903,I1068583,I630943,I630979,I1068565,I1068586,I630996,I1068568,I631022,I631030,I631047,I631078,I631095,I631112,I631143,I631174,I631191,I631246,I631272,I631280,I631297,I631314,I631340,I631235,I631371,I631379,I631396,I631422,I631430,I631238,I631470,I631229,I631220,I631506,I631523,I631549,I631557,I631574,I631223,I631605,I631622,I631639,I631232,I631670,I631217,I631701,I631718,I631226,I631773,I631799,I631807,I631824,I631841,I631867,I631762,I631898,I631906,I631923,I631949,I631957,I631765,I631997,I631756,I631747,I632033,I632050,I632076,I632084,I632101,I631750,I632132,I632149,I632166,I631759,I632197,I631744,I632228,I632245,I631753,I632300,I632326,I632334,I632351,I632368,I632394,I632425,I632433,I632450,I632476,I632484,I632524,I632560,I632577,I632603,I632611,I632628,I632659,I632676,I632693,I632724,I632755,I632772,I632827,I632853,I632861,I632878,I632895,I632921,I632952,I632960,I632977,I633003,I633011,I633051,I633087,I633104,I633130,I633138,I633155,I633186,I633203,I633220,I633251,I633282,I633299,I633354,I1042989,I633380,I633388,I633405,I1042986,I1042995,I633422,I1042974,I633448,I1042977,I633479,I633487,I1042992,I633504,I633530,I633538,I1042998,I633578,I633614,I1042980,I1043001,I633631,I1042983,I633657,I633665,I633682,I633713,I633730,I633747,I633778,I633809,I633826,I633881,I823717,I633907,I633915,I633932,I823726,I823714,I633949,I823711,I633975,I634006,I634014,I823708,I634031,I634057,I634065,I634105,I634141,I823729,I823720,I634158,I823723,I634184,I634192,I634209,I634240,I634257,I634274,I634305,I634336,I634353,I634408,I634434,I634442,I634459,I634476,I634502,I634533,I634541,I634558,I634584,I634592,I634632,I634668,I634685,I634711,I634719,I634736,I634767,I634784,I634801,I634832,I634863,I634880,I634935,I822595,I634961,I634969,I634986,I822604,I822592,I635003,I822589,I635029,I635060,I635068,I822586,I635085,I635111,I635119,I635159,I635195,I822607,I822598,I635212,I822601,I635238,I635246,I635263,I635294,I635311,I635328,I635359,I635390,I635407,I635462,I635488,I635496,I635513,I635530,I635556,I635587,I635595,I635612,I635638,I635646,I635686,I635722,I635739,I635765,I635773,I635790,I635821,I635838,I635855,I635886,I635917,I635934,I635989,I636015,I636023,I636040,I636057,I636083,I636114,I636122,I636139,I636165,I636173,I636213,I636249,I636266,I636292,I636300,I636317,I636348,I636365,I636382,I636413,I636444,I636461,I636516,I636542,I636550,I636567,I636584,I636610,I636641,I636649,I636666,I636692,I636700,I636740,I636776,I636793,I636819,I636827,I636844,I636875,I636892,I636909,I636940,I636971,I636988,I637043,I637069,I637077,I637094,I637111,I637137,I637168,I637176,I637193,I637219,I637227,I637267,I637303,I637320,I637346,I637354,I637371,I637402,I637419,I637436,I637467,I637498,I637515,I637570,I637596,I637604,I637621,I637638,I637664,I637695,I637703,I637720,I637746,I637754,I637794,I637830,I637847,I637873,I637881,I637898,I637929,I637946,I637963,I637994,I638025,I638042,I638097,I943236,I638123,I638131,I638148,I943218,I638165,I943224,I638191,I638086,I943221,I638222,I638230,I943230,I638247,I638273,I638281,I638089,I943242,I638321,I638080,I638071,I638357,I943233,I943227,I638374,I638400,I638408,I638425,I638074,I638456,I943239,I638473,I638490,I638083,I638521,I638068,I638552,I638569,I638077,I638624,I733560,I638650,I638658,I638675,I733575,I733557,I638692,I638718,I733566,I638749,I638757,I733584,I638774,I638800,I638808,I733581,I638848,I638884,I733578,I733569,I638901,I733563,I638927,I638935,I638952,I638983,I733572,I639000,I639017,I639048,I639079,I639096,I639151,I986954,I639177,I639185,I639202,I986960,I986942,I639219,I986951,I639245,I639140,I986957,I639276,I639284,I986945,I639301,I639327,I639335,I639143,I986963,I639375,I639134,I639125,I639411,I986948,I639428,I986966,I639454,I639462,I639479,I639128,I639510,I639527,I639544,I639137,I639575,I639122,I639606,I639623,I639131,I639678,I769090,I639704,I639712,I639729,I769105,I769087,I639746,I639772,I639667,I769096,I639803,I639811,I769114,I639828,I639854,I639862,I639670,I769111,I639902,I639661,I639652,I639938,I769108,I769099,I639955,I769093,I639981,I639989,I640006,I639655,I640037,I769102,I640054,I640071,I639664,I640102,I639649,I640133,I640150,I639658,I640205,I640231,I640239,I640256,I640273,I640299,I640194,I640330,I640338,I640355,I640381,I640389,I640197,I640429,I640188,I640179,I640465,I640482,I640508,I640516,I640533,I640182,I640564,I640581,I640598,I640191,I640629,I640176,I640660,I640677,I640185,I640732,I640758,I640766,I640783,I640800,I640826,I640857,I640865,I640882,I640908,I640916,I640956,I640992,I641009,I641035,I641043,I641060,I641091,I641108,I641125,I641156,I641187,I641204,I641259,I641285,I641293,I641310,I641327,I641353,I641248,I641384,I641392,I641409,I641435,I641443,I641251,I641483,I641242,I641233,I641519,I641536,I641562,I641570,I641587,I641236,I641618,I641635,I641652,I641245,I641683,I641230,I641714,I641731,I641239,I641786,I641812,I641820,I641837,I641854,I641880,I641911,I641919,I641936,I641962,I641970,I642010,I642046,I642063,I642089,I642097,I642114,I642145,I642162,I642179,I642210,I642241,I642258,I642313,I946126,I642339,I642347,I642364,I946108,I642381,I946114,I642407,I946111,I642438,I642446,I946120,I642463,I642489,I642497,I946132,I642537,I642573,I946123,I946117,I642590,I642616,I642624,I642641,I642672,I946129,I642689,I642706,I642737,I642768,I642785,I642840,I810253,I642866,I642874,I642891,I810262,I810250,I642908,I810247,I642934,I642829,I642965,I642973,I810244,I642990,I643016,I643024,I642832,I643064,I642823,I642814,I643100,I810265,I810256,I643117,I810259,I643143,I643151,I643168,I642817,I643199,I643216,I643233,I642826,I643264,I642811,I643295,I643312,I642820,I643367,I643393,I643401,I643418,I643435,I643461,I643492,I643500,I643517,I643543,I643551,I643591,I643627,I643644,I643670,I643678,I643695,I643726,I643743,I643760,I643791,I643822,I643839,I643894,I643920,I643928,I643945,I643962,I643988,I644019,I644027,I644044,I644070,I644078,I644118,I644154,I644171,I644197,I644205,I644222,I644253,I644270,I644287,I644318,I644349,I644366,I644421,I644447,I644455,I644472,I644489,I644515,I644410,I644546,I644554,I644571,I644597,I644605,I644413,I644645,I644404,I644395,I644681,I644698,I644724,I644732,I644749,I644398,I644780,I644797,I644814,I644407,I644845,I644392,I644876,I644893,I644401,I644948,I783948,I644974,I644982,I644999,I783963,I783945,I645016,I645042,I644937,I783954,I645073,I645081,I783972,I645098,I645124,I645132,I644940,I783969,I645172,I644931,I644922,I645208,I783966,I783957,I645225,I783951,I645251,I645259,I645276,I644925,I645307,I783960,I645324,I645341,I644934,I645372,I644919,I645403,I645420,I644928,I645475,I1079284,I645501,I645509,I645526,I1079281,I1079290,I645543,I1079269,I645569,I1079272,I645600,I645608,I1079287,I645625,I645651,I645659,I1079293,I645699,I645735,I1079275,I1079296,I645752,I1079278,I645778,I645786,I645803,I645834,I645851,I645868,I645899,I645930,I645947,I646002,I646028,I646036,I646053,I646070,I646096,I645991,I646127,I646135,I646152,I646178,I646186,I645994,I646226,I645985,I645976,I646262,I646279,I646305,I646313,I646330,I645979,I646361,I646378,I646395,I645988,I646426,I645973,I646457,I646474,I645982,I646529,I646555,I646563,I646580,I646597,I646623,I646518,I646654,I646662,I646679,I646705,I646713,I646521,I646753,I646512,I646503,I646789,I646806,I646832,I646840,I646857,I646506,I646888,I646905,I646922,I646515,I646953,I646500,I646984,I647001,I646509,I647056,I647082,I647090,I647107,I647124,I647150,I647045,I647181,I647189,I647206,I647232,I647240,I647048,I647280,I647039,I647030,I647316,I647333,I647359,I647367,I647384,I647033,I647415,I647432,I647449,I647042,I647480,I647027,I647511,I647528,I647036,I647583,I647609,I647617,I647634,I647651,I647677,I647572,I647708,I647716,I647733,I647759,I647767,I647575,I647807,I647566,I647557,I647843,I647860,I647886,I647894,I647911,I647560,I647942,I647959,I647976,I647569,I648007,I647554,I648038,I648055,I647563,I648110,I648136,I648144,I648161,I648178,I648204,I648099,I648235,I648243,I648260,I648286,I648294,I648102,I648334,I648093,I648084,I648370,I648387,I648413,I648421,I648438,I648087,I648469,I648486,I648503,I648096,I648534,I648081,I648565,I648582,I648090,I648637,I1028241,I648663,I648671,I648688,I1028235,I1028253,I648705,I1028238,I648731,I1028259,I648762,I648770,I1028244,I648787,I648813,I648821,I1028256,I648861,I648897,I1028247,I1028262,I648914,I1028250,I648940,I648948,I648965,I648996,I649013,I649030,I649061,I649092,I649109,I649164,I649190,I649198,I649215,I649232,I649258,I649289,I649297,I649314,I649340,I649348,I649388,I649424,I649441,I649467,I649475,I649492,I649523,I649540,I649557,I649588,I649619,I649636,I649691,I954796,I649717,I649725,I649742,I954778,I649759,I954784,I649785,I649680,I954781,I649816,I649824,I954790,I649841,I649867,I649875,I649683,I954802,I649915,I649674,I649665,I649951,I954793,I954787,I649968,I649994,I650002,I650019,I649668,I650050,I954799,I650067,I650084,I649677,I650115,I649662,I650146,I650163,I649671,I650218,I917804,I650244,I650252,I650269,I917786,I650286,I917792,I650312,I917789,I650343,I650351,I917798,I650368,I650394,I650402,I917810,I650442,I650478,I917801,I917795,I650495,I650521,I650529,I650546,I650577,I917807,I650594,I650611,I650642,I650673,I650690,I650745,I852490,I650771,I650779,I650796,I852472,I650813,I852478,I650839,I852475,I650870,I650878,I852484,I650895,I650921,I650929,I852496,I650969,I651005,I852487,I852481,I651022,I651048,I651056,I651073,I651104,I852493,I651121,I651138,I651169,I651200,I651217,I651272,I651298,I651306,I651323,I651340,I651366,I651397,I651405,I651422,I651448,I651456,I651496,I651532,I651549,I651575,I651583,I651600,I651631,I651648,I651665,I651696,I651727,I651744,I651799,I816424,I651825,I651833,I651850,I816433,I816421,I651867,I816418,I651893,I651788,I651924,I651932,I816415,I651949,I651975,I651983,I651791,I652023,I651782,I651773,I652059,I816436,I816427,I652076,I816430,I652102,I652110,I652127,I651776,I652158,I652175,I652192,I651785,I652223,I651770,I652254,I652271,I651779,I652326,I652352,I652360,I652377,I652394,I652420,I652451,I652459,I652476,I652502,I652510,I652550,I652586,I652603,I652629,I652637,I652654,I652685,I652702,I652719,I652750,I652781,I652798,I652853,I1050129,I652879,I652887,I652904,I1050126,I1050135,I652921,I1050114,I652947,I1050117,I652978,I652986,I1050132,I653003,I653029,I653037,I1050138,I653077,I653113,I1050120,I1050141,I653130,I1050123,I653156,I653164,I653181,I653212,I653229,I653246,I653277,I653308,I653325,I653380,I653406,I653414,I653431,I653448,I653474,I653369,I653505,I653513,I653530,I653556,I653564,I653372,I653604,I653363,I653354,I653640,I653657,I653683,I653691,I653708,I653357,I653739,I653756,I653773,I653366,I653804,I653351,I653835,I653852,I653360,I653907,I653933,I653941,I653958,I653975,I654001,I654032,I654040,I654057,I654083,I654091,I654131,I654167,I654184,I654210,I654218,I654235,I654266,I654283,I654300,I654331,I654362,I654379,I654434,I654460,I654468,I654485,I654502,I654528,I654423,I654559,I654567,I654584,I654610,I654618,I654426,I654658,I654417,I654408,I654694,I654711,I654737,I654745,I654762,I654411,I654793,I654810,I654827,I654420,I654858,I654405,I654889,I654906,I654414,I654961,I654987,I654995,I655012,I655029,I655055,I654950,I655086,I655094,I655111,I655137,I655145,I654953,I655185,I654944,I654935,I655221,I655238,I655264,I655272,I655289,I654938,I655320,I655337,I655354,I654947,I655385,I654932,I655416,I655433,I654941,I655488,I1011712,I655514,I655522,I655539,I1011694,I1011697,I655556,I1011709,I655582,I655477,I1011718,I655613,I655621,I1011703,I655638,I655664,I655672,I655480,I1011715,I655712,I655471,I655462,I655748,I1011706,I1011700,I655765,I655791,I655799,I655816,I655465,I655847,I655864,I655881,I655474,I655912,I655459,I655943,I655960,I655468,I656015,I656041,I656049,I656066,I656083,I656109,I656140,I656148,I656165,I656191,I656199,I656239,I656275,I656292,I656318,I656326,I656343,I656374,I656391,I656408,I656439,I656470,I656487,I656542,I840930,I656568,I656576,I656593,I840912,I656610,I840918,I656636,I656531,I840915,I656667,I656675,I840924,I656692,I656718,I656726,I656534,I840936,I656766,I656525,I656516,I656802,I840927,I840921,I656819,I656845,I656853,I656870,I656519,I656901,I840933,I656918,I656935,I656528,I656966,I656513,I656997,I657014,I656522,I657069,I657095,I657103,I657120,I657137,I657163,I657194,I657202,I657219,I657245,I657253,I657293,I657329,I657346,I657372,I657380,I657397,I657428,I657445,I657462,I657493,I657524,I657541,I657596,I657622,I657630,I657647,I657664,I657690,I657721,I657729,I657746,I657772,I657780,I657820,I657856,I657873,I657899,I657907,I657924,I657955,I657972,I657989,I658020,I658051,I658068,I658123,I658149,I658157,I658174,I658191,I658217,I658248,I658256,I658273,I658299,I658307,I658347,I658383,I658400,I658426,I658434,I658451,I658482,I658499,I658516,I658547,I658578,I658595,I658650,I658676,I658684,I658701,I658718,I658744,I658775,I658783,I658800,I658826,I658834,I658874,I658910,I658927,I658953,I658961,I658978,I659009,I659026,I659043,I659074,I659105,I659122,I659177,I1051319,I659203,I659211,I659228,I1051316,I1051325,I659245,I1051304,I659271,I1051307,I659302,I659310,I1051322,I659327,I659353,I659361,I1051328,I659401,I659437,I1051310,I1051331,I659454,I1051313,I659480,I659488,I659505,I659536,I659553,I659570,I659601,I659632,I659649,I659704,I659730,I659738,I659755,I659772,I659798,I659829,I659837,I659854,I659880,I659888,I659928,I659964,I659981,I660007,I660015,I660032,I660063,I660080,I660097,I660128,I660159,I660176,I660231,I906822,I660257,I660265,I660282,I906804,I660299,I906810,I660325,I660220,I906807,I660356,I660364,I906816,I660381,I660407,I660415,I660223,I906828,I660455,I660214,I660205,I660491,I906819,I906813,I660508,I660534,I660542,I660559,I660208,I660590,I906825,I660607,I660624,I660217,I660655,I660202,I660686,I660703,I660211,I660758,I844398,I660784,I660792,I660809,I844380,I660826,I844386,I660852,I844383,I660883,I660891,I844392,I660908,I660934,I660942,I844404,I660982,I661018,I844395,I844389,I661035,I661061,I661069,I661086,I661117,I844401,I661134,I661151,I661182,I661213,I661230,I661285,I661311,I661319,I661336,I661353,I661379,I661274,I661410,I661418,I661435,I661461,I661469,I661277,I661509,I661268,I661259,I661545,I661562,I661588,I661596,I661613,I661262,I661644,I661661,I661678,I661271,I661709,I661256,I661740,I661757,I661265,I661812,I848444,I661838,I661846,I661863,I848426,I661880,I848432,I661906,I848429,I661937,I661945,I848438,I661962,I661988,I661996,I848450,I662036,I662072,I848441,I848435,I662089,I662115,I662123,I662140,I662171,I848447,I662188,I662205,I662236,I662267,I662284,I662339,I726454,I662365,I662373,I662390,I726469,I726451,I662407,I662433,I662328,I726460,I662464,I662472,I726478,I662489,I662515,I662523,I662331,I726475,I662563,I662322,I662313,I662599,I726472,I726463,I662616,I726457,I662642,I662650,I662667,I662316,I662698,I726466,I662715,I662732,I662325,I662763,I662310,I662794,I662811,I662319,I662866,I662892,I662900,I662917,I662934,I662960,I662991,I662999,I663016,I663042,I663050,I663090,I663126,I663143,I663169,I663177,I663194,I663225,I663242,I663259,I663290,I663321,I663338,I663393,I663419,I663427,I663444,I663461,I663487,I663518,I663526,I663543,I663569,I663577,I663617,I663653,I663670,I663696,I663704,I663721,I663752,I663769,I663786,I663817,I663848,I663865,I663920,I856536,I663946,I663954,I663971,I856518,I663988,I856524,I664014,I663909,I856521,I664045,I664053,I856530,I664070,I664096,I664104,I663912,I856542,I664144,I663903,I663894,I664180,I856533,I856527,I664197,I664223,I664231,I664248,I663897,I664279,I856539,I664296,I664313,I663906,I664344,I663891,I664375,I664392,I663900,I664447,I702552,I664473,I664481,I664498,I702567,I702549,I664515,I664541,I664436,I702558,I664572,I664580,I702576,I664597,I664623,I664631,I664439,I702573,I664671,I664430,I664421,I664707,I702570,I702561,I664724,I702555,I664750,I664758,I664775,I664424,I664806,I702564,I664823,I664840,I664433,I664871,I664418,I664902,I664919,I664427,I664974,I665000,I665008,I665025,I665042,I665068,I665099,I665107,I665124,I665150,I665158,I665198,I665234,I665251,I665277,I665285,I665302,I665333,I665350,I665367,I665398,I665429,I665446,I665501,I750356,I665527,I665535,I665552,I750371,I750353,I665569,I665595,I665490,I750362,I665626,I665634,I750380,I665651,I665677,I665685,I665493,I750377,I665725,I665484,I665475,I665761,I750374,I750365,I665778,I750359,I665804,I665812,I665829,I665478,I665860,I750368,I665877,I665894,I665487,I665925,I665472,I665956,I665973,I665481,I666028,I811375,I666054,I666062,I666079,I811384,I811372,I666096,I811369,I666122,I666153,I666161,I811366,I666178,I666204,I666212,I666252,I666288,I811387,I811378,I666305,I811381,I666331,I666339,I666356,I666387,I666404,I666421,I666452,I666483,I666500,I666555,I666581,I666589,I666606,I666623,I666649,I666680,I666688,I666705,I666731,I666739,I666779,I666815,I666832,I666858,I666866,I666883,I666914,I666931,I666948,I666979,I667010,I667027,I667082,I667108,I667116,I667133,I667150,I667176,I667207,I667215,I667232,I667258,I667266,I667306,I667342,I667359,I667385,I667393,I667410,I667441,I667458,I667475,I667506,I667537,I667554,I667609,I1055484,I667635,I667643,I667660,I1055481,I1055490,I667677,I1055469,I667703,I1055472,I667734,I667742,I1055487,I667759,I667785,I667793,I1055493,I667833,I667869,I1055475,I1055496,I667886,I1055478,I667912,I667920,I667937,I667968,I667985,I668002,I668033,I668064,I668081,I668136,I1074524,I668162,I668170,I668187,I1074521,I1074530,I668204,I1074509,I668230,I1074512,I668261,I668269,I1074527,I668286,I668312,I668320,I1074533,I668360,I668396,I1074515,I1074536,I668413,I1074518,I668439,I668447,I668464,I668495,I668512,I668529,I668560,I668591,I668608,I668663,I668689,I668697,I668714,I668731,I668757,I668788,I668796,I668813,I668839,I668847,I668887,I668923,I668940,I668966,I668974,I668991,I669022,I669039,I669056,I669087,I669118,I669135,I669190,I669216,I669224,I669241,I669258,I669284,I669315,I669323,I669340,I669366,I669374,I669414,I669450,I669467,I669493,I669501,I669518,I669549,I669566,I669583,I669614,I669645,I669662,I669717,I1073929,I669743,I669751,I669768,I1073926,I1073935,I669785,I1073914,I669811,I1073917,I669842,I669850,I1073932,I669867,I669893,I669901,I1073938,I669941,I669977,I1073920,I1073941,I669994,I1073923,I670020,I670028,I670045,I670076,I670093,I670110,I670141,I670172,I670189,I670244,I796228,I670270,I670278,I670295,I796237,I796225,I670312,I796222,I670338,I670369,I670377,I796219,I670394,I670420,I670428,I670468,I670504,I796240,I796231,I670521,I796234,I670547,I670555,I670572,I670603,I670620,I670637,I670668,I670699,I670716,I670771,I849600,I670797,I670805,I670822,I849582,I670839,I849588,I670865,I670760,I849585,I670896,I670904,I849594,I670921,I670947,I670955,I670763,I849606,I670995,I670754,I670745,I671031,I849597,I849591,I671048,I671074,I671082,I671099,I670748,I671130,I849603,I671147,I671164,I670757,I671195,I670742,I671226,I671243,I670751,I671298,I671324,I671332,I671349,I671366,I671392,I671423,I671431,I671448,I671474,I671482,I671522,I671558,I671575,I671601,I671609,I671626,I671657,I671674,I671691,I671722,I671753,I671770,I671825,I864050,I671851,I671859,I671876,I864032,I671893,I864038,I671919,I671814,I864035,I671950,I671958,I864044,I671975,I672001,I672009,I671817,I864056,I672049,I671808,I671799,I672085,I864047,I864041,I672102,I672128,I672136,I672153,I671802,I672184,I864053,I672201,I672218,I671811,I672249,I671796,I672280,I672297,I671805,I672352,I862316,I672378,I672386,I672403,I862298,I672420,I862304,I672446,I862301,I672477,I672485,I862310,I672502,I672528,I672536,I862322,I672576,I672612,I862313,I862307,I672629,I672655,I672663,I672680,I672711,I862319,I672728,I672745,I672776,I672807,I672824,I672879,I829370,I672905,I672913,I672930,I829352,I672947,I829358,I672973,I829355,I673004,I673012,I829364,I673029,I673055,I673063,I829376,I673103,I673139,I829367,I829361,I673156,I673182,I673190,I673207,I673238,I829373,I673255,I673272,I673303,I673334,I673351,I673406,I1097729,I673432,I673440,I673457,I1097726,I1097735,I673474,I1097714,I673500,I673395,I1097717,I673531,I673539,I1097732,I673556,I673582,I673590,I673398,I1097738,I673630,I673389,I673380,I673666,I1097720,I1097741,I673683,I1097723,I673709,I673717,I673734,I673383,I673765,I673782,I673799,I673392,I673830,I673377,I673861,I673878,I673386,I673933,I715472,I673959,I673967,I673984,I715487,I715469,I674001,I674027,I715478,I674058,I674066,I715496,I674083,I674109,I674117,I715493,I674157,I674193,I715490,I715481,I674210,I715475,I674236,I674244,I674261,I674292,I715484,I674309,I674326,I674357,I674388,I674405,I674460,I868096,I674486,I674494,I674511,I868078,I674528,I868084,I674554,I674449,I868081,I674585,I674593,I868090,I674610,I674636,I674644,I674452,I868102,I674684,I674443,I674434,I674720,I868093,I868087,I674737,I674763,I674771,I674788,I674437,I674819,I868099,I674836,I674853,I674446,I674884,I674431,I674915,I674932,I674440,I674987,I675013,I675021,I675038,I675055,I675081,I674976,I675112,I675120,I675137,I675163,I675171,I674979,I675211,I674970,I674961,I675247,I675264,I675290,I675298,I675315,I674964,I675346,I675363,I675380,I674973,I675411,I674958,I675442,I675459,I674967,I675514,I888904,I675540,I675548,I675565,I888886,I675582,I888892,I675608,I888889,I675639,I675647,I888898,I675664,I675690,I675698,I888910,I675738,I675774,I888901,I888895,I675791,I675817,I675825,I675842,I675873,I888907,I675890,I675907,I675938,I675969,I675986,I676041,I898152,I676067,I676075,I676092,I898134,I676109,I898140,I676135,I898137,I676166,I676174,I898146,I676191,I676217,I676225,I898158,I676265,I676301,I898149,I898143,I676318,I676344,I676352,I676369,I676400,I898155,I676417,I676434,I676465,I676496,I676513,I676568,I676594,I676602,I676619,I676636,I676662,I676693,I676701,I676718,I676744,I676752,I676792,I676828,I676845,I676871,I676879,I676896,I676927,I676944,I676961,I676992,I677023,I677040,I677095,I677121,I677129,I677146,I677163,I677189,I677220,I677228,I677245,I677271,I677279,I677319,I677355,I677372,I677398,I677406,I677423,I677454,I677471,I677488,I677519,I677550,I677567,I677622,I677648,I677656,I677673,I677690,I677716,I677611,I677747,I677755,I677772,I677798,I677806,I677614,I677846,I677605,I677596,I677882,I677899,I677925,I677933,I677950,I677599,I677981,I677998,I678015,I677608,I678046,I677593,I678077,I678094,I677602,I678149,I1041204,I678175,I678183,I678200,I1041201,I1041210,I678217,I1041189,I678243,I1041192,I678274,I678282,I1041207,I678299,I678325,I678333,I1041213,I678373,I678409,I1041195,I1041216,I678426,I1041198,I678452,I678460,I678477,I678508,I678525,I678542,I678573,I678604,I678621,I678676,I678702,I678710,I678727,I678744,I678770,I678801,I678809,I678826,I678852,I678860,I678900,I678936,I678953,I678979,I678987,I679004,I679035,I679052,I679069,I679100,I679131,I679148,I679203,I776842,I679229,I679237,I679254,I776857,I776839,I679271,I679297,I776848,I679328,I679336,I776866,I679353,I679379,I679387,I776863,I679427,I679463,I776860,I776851,I679480,I776845,I679506,I679514,I679531,I679562,I776854,I679579,I679596,I679627,I679658,I679675,I679730,I679756,I679764,I679781,I679798,I679824,I679719,I679855,I679863,I679880,I679906,I679914,I679722,I679954,I679713,I679704,I679990,I680007,I680033,I680041,I680058,I679707,I680089,I680106,I680123,I679716,I680154,I679701,I680185,I680202,I679710,I680257,I850756,I680283,I680291,I680308,I850738,I680325,I850744,I680351,I850741,I680382,I680390,I850750,I680407,I680433,I680441,I850762,I680481,I680517,I850753,I850747,I680534,I680560,I680568,I680585,I680616,I850759,I680633,I680650,I680681,I680712,I680729,I680784,I1080474,I680810,I680818,I680835,I1080471,I1080480,I680852,I1080459,I680878,I1080462,I680909,I680917,I1080477,I680934,I680960,I680968,I1080483,I681008,I681044,I1080465,I1080486,I681061,I1080468,I681087,I681095,I681112,I681143,I681160,I681177,I681208,I681239,I681256,I681311,I681337,I681345,I681362,I681379,I681405,I681300,I681436,I681444,I681461,I681487,I681495,I681303,I681535,I681294,I681285,I681571,I681588,I681614,I681622,I681639,I681288,I681670,I681687,I681704,I681297,I681735,I681282,I681766,I681783,I681291,I681838,I792992,I681864,I681872,I681889,I793007,I792989,I681906,I681932,I681827,I792998,I681963,I681971,I793016,I681988,I682014,I682022,I681830,I793013,I682062,I681821,I681812,I682098,I793010,I793001,I682115,I792995,I682141,I682149,I682166,I681815,I682197,I793004,I682214,I682231,I681824,I682262,I681809,I682293,I682310,I681818,I682365,I1029363,I682391,I682399,I682416,I1029357,I1029375,I682433,I1029360,I682459,I682354,I1029381,I682490,I682498,I1029366,I682515,I682541,I682549,I682357,I1029378,I682589,I682348,I682339,I682625,I1029369,I1029384,I682642,I1029372,I682668,I682676,I682693,I682342,I682724,I682741,I682758,I682351,I682789,I682336,I682820,I682837,I682345,I682892,I682918,I682926,I682943,I682960,I682986,I682881,I683017,I683025,I683042,I683068,I683076,I682884,I683116,I682875,I682866,I683152,I683169,I683195,I683203,I683220,I682869,I683251,I683268,I683285,I682878,I683316,I682863,I683347,I683364,I682872,I683419,I937456,I683445,I683453,I683470,I937438,I683487,I937444,I683513,I683408,I937441,I683544,I683552,I937450,I683569,I683595,I683603,I683411,I937462,I683643,I683402,I683393,I683679,I937453,I937447,I683696,I683722,I683730,I683747,I683396,I683778,I937459,I683795,I683812,I683405,I683843,I683390,I683874,I683891,I683399,I683946,I683972,I683980,I683997,I684014,I684040,I684071,I684079,I684096,I684122,I684130,I684170,I684206,I684223,I684249,I684257,I684274,I684305,I684322,I684339,I684370,I684401,I684418,I684473,I684499,I684507,I684524,I684541,I684567,I684598,I684606,I684623,I684649,I684657,I684697,I684733,I684750,I684776,I684784,I684801,I684832,I684849,I684866,I684897,I684928,I684945,I685000,I970090,I685026,I685034,I685051,I970096,I970078,I685068,I970087,I685094,I684989,I970093,I685125,I685133,I970081,I685150,I685176,I685184,I684992,I970099,I685224,I684983,I684974,I685260,I970084,I685277,I970102,I685303,I685311,I685328,I684977,I685359,I685376,I685393,I684986,I685424,I684971,I685455,I685472,I684980,I685527,I1004776,I685553,I685561,I685578,I1004758,I1004761,I685595,I1004773,I685621,I685516,I1004782,I685652,I685660,I1004767,I685677,I685703,I685711,I685519,I1004779,I685751,I685510,I685501,I685787,I1004770,I1004764,I685804,I685830,I685838,I685855,I685504,I685886,I685903,I685920,I685513,I685951,I685498,I685982,I685999,I685507,I686054,I686080,I686088,I686105,I686122,I686148,I686179,I686187,I686204,I686230,I686238,I686278,I686314,I686331,I686357,I686365,I686382,I686413,I686430,I686447,I686478,I686509,I686526,I686581,I686607,I686615,I686632,I686649,I686675,I686706,I686714,I686731,I686757,I686765,I686805,I686841,I686858,I686884,I686892,I686909,I686940,I686957,I686974,I687005,I687036,I687053,I687108,I687134,I687142,I687159,I687176,I687202,I687233,I687241,I687258,I687284,I687292,I687332,I687368,I687385,I687411,I687419,I687436,I687467,I687484,I687501,I687532,I687563,I687580,I687635,I687661,I687669,I687686,I687703,I687729,I687760,I687768,I687785,I687811,I687819,I687859,I687895,I687912,I687938,I687946,I687963,I687994,I688011,I688028,I688059,I688090,I688107,I688162,I688188,I688196,I688213,I688230,I688256,I688151,I688287,I688295,I688312,I688338,I688346,I688154,I688386,I688145,I688136,I688422,I688439,I688465,I688473,I688490,I688139,I688521,I688538,I688555,I688148,I688586,I688133,I688617,I688634,I688142,I688689,I782010,I688715,I688723,I688740,I782025,I782007,I688757,I688783,I782016,I688814,I688822,I782034,I688839,I688865,I688873,I782031,I688913,I688949,I782028,I782019,I688966,I782013,I688992,I689000,I689017,I689048,I782022,I689065,I689082,I689113,I689144,I689161,I689216,I689242,I689250,I689267,I689284,I689310,I689205,I689341,I689349,I689366,I689392,I689400,I689208,I689440,I689199,I689190,I689476,I689493,I689519,I689527,I689544,I689193,I689575,I689592,I689609,I689202,I689640,I689187,I689671,I689688,I689196,I689743,I689769,I689777,I689794,I689811,I689837,I689868,I689876,I689893,I689919,I689927,I689967,I690003,I690020,I690046,I690054,I690071,I690102,I690119,I690136,I690167,I690198,I690215,I690270,I690296,I690304,I690321,I690338,I690364,I690395,I690403,I690420,I690446,I690454,I690494,I690530,I690547,I690573,I690581,I690598,I690629,I690646,I690663,I690694,I690725,I690742,I690797,I1100109,I690823,I690831,I690848,I1100106,I1100115,I690865,I1100094,I690891,I1100097,I690922,I690930,I1100112,I690947,I690973,I690981,I1100118,I691021,I691057,I1100100,I1100121,I691074,I1100103,I691100,I691108,I691125,I691156,I691173,I691190,I691221,I691252,I691269,I691324,I691350,I691358,I691375,I691392,I691418,I691449,I691457,I691474,I691500,I691508,I691548,I691584,I691601,I691627,I691635,I691652,I691683,I691700,I691717,I691748,I691779,I691796,I691851,I691877,I691885,I691902,I691919,I691945,I691976,I691984,I692001,I692027,I692035,I692075,I692111,I692128,I692154,I692162,I692179,I692210,I692227,I692244,I692275,I692306,I692323,I692378,I692404,I692412,I692429,I692446,I692472,I692503,I692511,I692528,I692554,I692562,I692602,I692638,I692655,I692681,I692689,I692706,I692737,I692754,I692771,I692802,I692833,I692850,I692905,I1088209,I692931,I692939,I692956,I1088206,I1088215,I692973,I1088194,I692999,I1088197,I693030,I693038,I1088212,I693055,I693081,I693089,I1088218,I693129,I693165,I1088200,I1088221,I693182,I1088203,I693208,I693216,I693233,I693264,I693281,I693298,I693329,I693360,I693377,I693432,I717410,I693458,I693466,I693483,I717425,I717407,I693500,I693526,I693421,I717416,I693557,I693565,I717434,I693582,I693608,I693616,I693424,I717431,I693656,I693415,I693406,I693692,I717428,I717419,I693709,I717413,I693735,I693743,I693760,I693409,I693791,I717422,I693808,I693825,I693418,I693856,I693403,I693887,I693904,I693412,I693959,I879656,I693985,I693993,I694010,I879638,I694027,I879644,I694053,I879641,I694084,I694092,I879650,I694109,I694135,I694143,I879662,I694183,I694219,I879653,I879647,I694236,I694262,I694270,I694287,I694318,I879659,I694335,I694352,I694383,I694414,I694431,I694486,I694512,I694520,I694537,I694554,I694580,I694611,I694619,I694636,I694662,I694670,I694710,I694746,I694763,I694789,I694797,I694814,I694845,I694862,I694879,I694910,I694941,I694958,I695013,I850178,I695039,I695047,I695064,I850160,I695081,I850166,I695107,I695002,I850163,I695138,I695146,I850172,I695163,I695189,I695197,I695005,I850184,I695237,I694996,I694987,I695273,I850175,I850169,I695290,I695316,I695324,I695341,I694990,I695372,I850181,I695389,I695406,I694999,I695437,I694984,I695468,I695485,I694993,I695540,I695566,I695574,I695591,I695608,I695634,I695665,I695673,I695690,I695716,I695724,I695764,I695800,I695817,I695843,I695851,I695868,I695899,I695916,I695933,I695964,I695995,I696012,I696067,I835150,I696093,I696101,I696118,I835132,I696135,I835138,I696161,I835135,I696192,I696200,I835144,I696217,I696243,I696251,I835156,I696291,I696327,I835147,I835141,I696344,I696370,I696378,I696395,I696426,I835153,I696443,I696460,I696491,I696522,I696539,I696594,I696620,I696628,I696645,I696662,I696688,I696719,I696727,I696744,I696770,I696778,I696818,I696854,I696871,I696897,I696905,I696922,I696953,I696970,I696987,I697018,I697049,I697066,I697121,I789116,I697147,I697155,I697172,I789131,I789113,I697189,I697215,I697110,I789122,I697246,I697254,I789140,I697271,I697297,I697305,I697113,I789137,I697345,I697104,I697095,I697381,I789134,I789125,I697398,I789119,I697424,I697432,I697449,I697098,I697480,I789128,I697497,I697514,I697107,I697545,I697092,I697576,I697593,I697101,I697648,I697674,I697682,I697699,I697716,I697742,I697637,I697773,I697781,I697798,I697824,I697832,I697640,I697872,I697631,I697622,I697908,I697925,I697951,I697959,I697976,I697625,I698007,I698024,I698041,I697634,I698072,I697619,I698103,I698120,I697628,I698175,I764568,I698201,I698209,I698226,I764583,I764565,I698243,I698269,I764574,I698300,I698308,I764592,I698325,I698351,I698359,I764589,I698399,I698435,I764586,I764577,I698452,I764571,I698478,I698486,I698503,I698534,I764580,I698551,I698568,I698599,I698630,I698647,I698708,I698734,I698751,I698759,I698776,I698793,I698810,I698827,I698844,I698875,I698892,I698923,I698940,I698957,I698988,I699028,I699036,I699053,I699070,I699087,I699118,I699135,I699152,I699178,I699200,I699217,I699248,I699293,I699354,I699380,I699397,I699405,I699422,I699439,I699456,I699473,I699490,I699521,I699538,I699569,I699586,I699603,I699634,I699674,I699682,I699699,I699716,I699733,I699764,I699781,I699798,I699824,I699846,I699863,I699894,I699939,I700000,I700026,I700043,I700051,I700068,I700085,I700102,I700119,I700136,I700167,I700184,I700215,I700232,I700249,I700280,I700320,I700328,I700345,I700362,I700379,I700410,I700427,I700444,I700470,I700492,I700509,I700540,I700585,I700646,I700672,I700689,I700697,I700714,I700731,I700748,I700765,I700782,I700632,I700813,I700830,I700635,I700861,I700878,I700895,I700611,I700926,I700623,I700966,I700974,I700991,I701008,I701025,I700638,I701056,I701073,I701090,I701116,I700626,I701138,I701155,I700620,I701186,I700614,I700617,I701231,I700629,I701292,I701318,I701335,I701343,I701360,I701377,I701394,I701411,I701428,I701459,I701476,I701507,I701524,I701541,I701572,I701612,I701620,I701637,I701654,I701671,I701702,I701719,I701736,I701762,I701784,I701801,I701832,I701877,I701938,I939768,I701964,I939750,I701981,I701989,I702006,I939759,I702023,I939771,I702040,I939753,I702057,I939762,I702074,I702105,I702122,I702153,I702170,I939774,I702187,I702218,I702258,I702266,I702283,I702300,I702317,I702348,I939756,I702365,I939765,I702382,I702408,I702430,I702447,I702478,I702523,I702584,I702610,I702627,I702635,I702652,I702669,I702686,I702703,I702720,I702751,I702768,I702799,I702816,I702833,I702864,I702904,I702912,I702929,I702946,I702963,I702994,I703011,I703028,I703054,I703076,I703093,I703124,I703169,I703230,I703256,I703273,I703281,I703298,I703315,I703332,I703349,I703366,I703397,I703414,I703445,I703462,I703479,I703510,I703550,I703558,I703575,I703592,I703609,I703640,I703657,I703674,I703700,I703722,I703739,I703770,I703815,I703876,I866362,I703902,I866344,I703919,I703927,I703944,I866353,I703961,I866365,I703978,I866347,I703995,I866356,I704012,I703862,I704043,I704060,I703865,I704091,I704108,I866368,I704125,I703841,I704156,I703853,I704196,I704204,I704221,I704238,I704255,I703868,I704286,I866350,I704303,I866359,I704320,I704346,I703856,I704368,I704385,I703850,I704416,I703844,I703847,I704461,I703859,I704522,I704548,I704565,I704573,I704590,I704607,I704624,I704641,I704658,I704508,I704689,I704706,I704511,I704737,I704754,I704771,I704487,I704802,I704499,I704842,I704850,I704867,I704884,I704901,I704514,I704932,I704949,I704966,I704992,I704502,I705014,I705031,I704496,I705062,I704490,I704493,I705107,I704505,I705168,I705194,I705211,I705219,I705236,I705253,I705270,I705287,I705304,I705335,I705352,I705383,I705400,I705417,I705448,I705488,I705496,I705513,I705530,I705547,I705578,I705595,I705612,I705638,I705660,I705677,I705708,I705753,I705814,I705840,I705857,I705865,I705882,I705899,I705916,I705933,I705950,I705800,I705981,I705998,I705803,I706029,I706046,I706063,I705779,I706094,I705791,I706134,I706142,I706159,I706176,I706193,I705806,I706224,I706241,I706258,I706284,I705794,I706306,I706323,I705788,I706354,I705782,I705785,I706399,I705797,I706460,I706486,I706503,I706511,I706528,I706545,I706562,I706579,I706596,I706446,I706627,I706644,I706449,I706675,I706692,I706709,I706425,I706740,I706437,I706780,I706788,I706805,I706822,I706839,I706452,I706870,I706887,I706904,I706930,I706440,I706952,I706969,I706434,I707000,I706428,I706431,I707045,I706443,I707106,I707132,I707149,I707157,I707174,I707191,I707208,I707225,I707242,I707273,I707290,I707321,I707338,I707355,I707386,I707426,I707434,I707451,I707468,I707485,I707516,I707533,I707550,I707576,I707598,I707615,I707646,I707691,I707752,I707778,I707795,I707803,I707820,I707837,I707854,I707871,I707888,I707919,I707936,I707967,I707984,I708001,I708032,I708072,I708080,I708097,I708114,I708131,I708162,I708179,I708196,I708222,I708244,I708261,I708292,I708337,I708398,I708424,I708441,I708449,I708466,I708483,I708500,I708517,I708534,I708565,I708582,I708613,I708630,I708647,I708678,I708718,I708726,I708743,I708760,I708777,I708808,I708825,I708842,I708868,I708890,I708907,I708938,I708983,I709044,I709070,I709087,I709095,I709112,I709129,I709146,I709163,I709180,I709030,I709211,I709228,I709033,I709259,I709276,I709293,I709009,I709324,I709021,I709364,I709372,I709389,I709406,I709423,I709036,I709454,I709471,I709488,I709514,I709024,I709536,I709553,I709018,I709584,I709012,I709015,I709629,I709027,I709690,I709716,I709733,I709741,I709758,I709775,I709792,I709809,I709826,I709857,I709874,I709905,I709922,I709939,I709970,I710010,I710018,I710035,I710052,I710069,I710100,I710117,I710134,I710160,I710182,I710199,I710230,I710275,I710336,I710362,I710379,I710387,I710404,I710421,I710438,I710455,I710472,I710503,I710520,I710551,I710568,I710585,I710616,I710656,I710664,I710681,I710698,I710715,I710746,I710763,I710780,I710806,I710828,I710845,I710876,I710921,I710982,I711008,I711025,I711033,I711050,I711067,I711084,I711101,I711118,I711149,I711166,I711197,I711214,I711231,I711262,I711302,I711310,I711327,I711344,I711361,I711392,I711409,I711426,I711452,I711474,I711491,I711522,I711567,I711628,I711654,I711671,I711679,I711696,I711713,I711730,I711747,I711764,I711795,I711812,I711843,I711860,I711877,I711908,I711948,I711956,I711973,I711990,I712007,I712038,I712055,I712072,I712098,I712120,I712137,I712168,I712213,I712274,I1077484,I712300,I1077508,I712317,I712325,I712342,I1077490,I712359,I1077499,I712376,I712393,I1077505,I712410,I712441,I712458,I712489,I712506,I1077502,I712523,I712554,I712594,I712602,I712619,I712636,I1077496,I712653,I712684,I1077487,I712701,I1077511,I712718,I1077493,I712744,I712766,I712783,I712814,I712859,I712920,I1070344,I712946,I1070368,I712963,I712971,I712988,I1070350,I713005,I1070359,I713022,I713039,I1070365,I713056,I713087,I713104,I713135,I713152,I1070362,I713169,I713200,I713240,I713248,I713265,I713282,I1070356,I713299,I713330,I1070347,I713347,I1070371,I713364,I1070353,I713390,I713412,I713429,I713460,I713505,I713566,I988048,I713592,I988054,I713609,I713617,I713634,I988051,I713651,I988030,I713668,I988033,I713685,I988039,I713702,I713733,I713750,I713781,I713798,I713815,I713846,I713886,I713894,I713911,I713928,I988042,I713945,I713976,I713993,I988036,I714010,I988045,I714036,I714058,I714075,I714106,I714151,I714212,I714238,I714255,I714263,I714280,I714297,I714314,I714331,I714348,I714379,I714396,I714427,I714444,I714461,I714492,I714532,I714540,I714557,I714574,I714591,I714622,I714639,I714656,I714682,I714704,I714721,I714752,I714797,I714858,I714884,I714901,I714909,I714926,I714943,I714960,I714977,I714994,I715025,I715042,I715073,I715090,I715107,I715138,I715178,I715186,I715203,I715220,I715237,I715268,I715285,I715302,I715328,I715350,I715367,I715398,I715443,I715504,I715530,I715547,I715555,I715572,I715589,I715606,I715623,I715640,I715671,I715688,I715719,I715736,I715753,I715784,I715824,I715832,I715849,I715866,I715883,I715914,I715931,I715948,I715974,I715996,I716013,I716044,I716089,I716150,I716176,I716193,I716201,I716218,I716235,I716252,I716269,I716286,I716317,I716334,I716365,I716382,I716399,I716430,I716470,I716478,I716495,I716512,I716529,I716560,I716577,I716594,I716620,I716642,I716659,I716690,I716735,I716796,I716822,I716839,I716847,I716864,I716881,I716898,I716915,I716932,I716963,I716980,I717011,I717028,I717045,I717076,I717116,I717124,I717141,I717158,I717175,I717206,I717223,I717240,I717266,I717288,I717305,I717336,I717381,I717442,I1067964,I717468,I1067988,I717485,I717493,I717510,I1067970,I717527,I1067979,I717544,I717561,I1067985,I717578,I717609,I717626,I717657,I717674,I1067982,I717691,I717722,I717762,I717770,I717787,I717804,I1067976,I717821,I717852,I1067967,I717869,I1067991,I717886,I1067973,I717912,I717934,I717951,I717982,I718027,I718088,I718114,I718131,I718139,I718156,I718173,I718190,I718207,I718224,I718255,I718272,I718303,I718320,I718337,I718368,I718408,I718416,I718433,I718450,I718467,I718498,I718515,I718532,I718558,I718580,I718597,I718628,I718673,I718734,I718760,I718777,I718785,I718802,I718819,I718836,I718853,I718870,I718901,I718918,I718949,I718966,I718983,I719014,I719054,I719062,I719079,I719096,I719113,I719144,I719161,I719178,I719204,I719226,I719243,I719274,I719319,I719380,I719406,I719423,I719431,I719448,I719465,I719482,I719499,I719516,I719366,I719547,I719564,I719369,I719595,I719612,I719629,I719345,I719660,I719357,I719700,I719708,I719725,I719742,I719759,I719372,I719790,I719807,I719824,I719850,I719360,I719872,I719889,I719354,I719920,I719348,I719351,I719965,I719363,I720026,I720052,I720069,I720077,I720094,I720111,I720128,I720145,I720162,I720193,I720210,I720241,I720258,I720275,I720306,I720346,I720354,I720371,I720388,I720405,I720436,I720453,I720470,I720496,I720518,I720535,I720566,I720611,I720672,I720698,I720715,I720723,I720740,I720757,I720774,I720791,I720808,I720658,I720839,I720856,I720661,I720887,I720904,I720921,I720637,I720952,I720649,I720992,I721000,I721017,I721034,I721051,I720664,I721082,I721099,I721116,I721142,I720652,I721164,I721181,I720646,I721212,I720640,I720643,I721257,I720655,I721318,I721344,I721361,I721369,I721386,I721403,I721420,I721437,I721454,I721485,I721502,I721533,I721550,I721567,I721598,I721638,I721646,I721663,I721680,I721697,I721728,I721745,I721762,I721788,I721810,I721827,I721858,I721903,I721964,I1063204,I721990,I1063228,I722007,I722015,I722032,I1063210,I722049,I1063219,I722066,I722083,I1063225,I722100,I721950,I722131,I722148,I721953,I722179,I722196,I1063222,I722213,I721929,I722244,I721941,I722284,I722292,I722309,I722326,I1063216,I722343,I721956,I722374,I1063207,I722391,I1063231,I722408,I1063213,I722434,I721944,I722456,I722473,I721938,I722504,I721932,I721935,I722549,I721947,I722610,I722636,I722653,I722661,I722678,I722695,I722712,I722729,I722746,I722777,I722794,I722825,I722842,I722859,I722890,I722930,I722938,I722955,I722972,I722989,I723020,I723037,I723054,I723080,I723102,I723119,I723150,I723195,I723256,I723282,I723299,I723307,I723324,I723341,I723358,I723375,I723392,I723423,I723440,I723471,I723488,I723505,I723536,I723576,I723584,I723601,I723618,I723635,I723666,I723683,I723700,I723726,I723748,I723765,I723796,I723841,I723902,I1095334,I723928,I1095358,I723945,I723953,I723970,I1095340,I723987,I1095349,I724004,I724021,I1095355,I724038,I724069,I724086,I724117,I724134,I1095352,I724151,I724182,I724222,I724230,I724247,I724264,I1095346,I724281,I724312,I1095337,I724329,I1095361,I724346,I1095343,I724372,I724394,I724411,I724442,I724487,I724548,I724574,I724591,I724599,I724616,I724633,I724650,I724667,I724684,I724715,I724732,I724763,I724780,I724797,I724828,I724868,I724876,I724893,I724910,I724927,I724958,I724975,I724992,I725018,I725040,I725057,I725088,I725133,I725194,I864628,I725220,I864610,I725237,I725245,I725262,I864619,I725279,I864631,I725296,I864613,I725313,I864622,I725330,I725361,I725378,I725409,I725426,I864634,I725443,I725474,I725514,I725522,I725539,I725556,I725573,I725604,I864616,I725621,I864625,I725638,I725664,I725686,I725703,I725734,I725779,I725840,I992051,I725866,I992045,I725883,I725891,I725908,I992054,I725925,I992066,I725942,I992048,I725959,I725976,I726007,I726024,I726055,I726072,I992042,I726089,I726120,I726160,I726168,I726185,I726202,I992063,I726219,I726250,I992057,I726267,I726284,I992060,I726310,I726332,I726349,I726380,I726425,I726486,I726512,I726529,I726537,I726554,I726571,I726588,I726605,I726622,I726653,I726670,I726701,I726718,I726735,I726766,I726806,I726814,I726831,I726848,I726865,I726896,I726913,I726930,I726956,I726978,I726995,I727026,I727071,I727132,I727158,I727175,I727183,I727200,I727217,I727234,I727251,I727268,I727299,I727316,I727347,I727364,I727381,I727412,I727452,I727460,I727477,I727494,I727511,I727542,I727559,I727576,I727602,I727624,I727641,I727672,I727717,I727778,I727804,I727821,I727829,I727846,I727863,I727880,I727897,I727914,I727764,I727945,I727962,I727767,I727993,I728010,I728027,I727743,I728058,I727755,I728098,I728106,I728123,I728140,I728157,I727770,I728188,I728205,I728222,I728248,I727758,I728270,I728287,I727752,I728318,I727746,I727749,I728363,I727761,I728424,I728450,I728467,I728475,I728492,I728509,I728526,I728543,I728560,I728410,I728591,I728608,I728413,I728639,I728656,I728673,I728389,I728704,I728401,I728744,I728752,I728769,I728786,I728803,I728416,I728834,I728851,I728868,I728894,I728404,I728916,I728933,I728398,I728964,I728392,I728395,I729009,I728407,I729070,I729096,I729113,I729121,I729138,I729155,I729172,I729189,I729206,I729237,I729254,I729285,I729302,I729319,I729350,I729390,I729398,I729415,I729432,I729449,I729480,I729497,I729514,I729540,I729562,I729579,I729610,I729655,I729716,I729742,I729759,I729767,I729784,I729801,I729818,I729835,I729852,I729883,I729900,I729931,I729948,I729965,I729996,I730036,I730044,I730061,I730078,I730095,I730126,I730143,I730160,I730186,I730208,I730225,I730256,I730301,I730362,I730388,I730405,I730413,I730430,I730447,I730464,I730481,I730498,I730348,I730529,I730546,I730351,I730577,I730594,I730611,I730327,I730642,I730339,I730682,I730690,I730707,I730724,I730741,I730354,I730772,I730789,I730806,I730832,I730342,I730854,I730871,I730336,I730902,I730330,I730333,I730947,I730345,I731008,I731034,I731051,I731059,I731076,I731093,I731110,I731127,I731144,I731175,I731192,I731223,I731240,I731257,I731288,I731328,I731336,I731353,I731370,I731387,I731418,I731435,I731452,I731478,I731500,I731517,I731548,I731593,I731654,I843820,I731680,I843802,I731697,I731705,I731722,I843811,I731739,I843823,I731756,I843805,I731773,I843814,I731790,I731821,I731838,I731869,I731886,I843826,I731903,I731934,I731974,I731982,I731999,I732016,I732033,I732064,I843808,I732081,I843817,I732098,I732124,I732146,I732163,I732194,I732239,I732300,I732326,I732343,I732351,I732368,I732385,I732402,I732419,I732436,I732467,I732484,I732515,I732532,I732549,I732580,I732620,I732628,I732645,I732662,I732679,I732710,I732727,I732744,I732770,I732792,I732809,I732840,I732885,I732946,I732972,I732989,I732997,I733014,I733031,I733048,I733065,I733082,I733113,I733130,I733161,I733178,I733195,I733226,I733266,I733274,I733291,I733308,I733325,I733356,I733373,I733390,I733416,I733438,I733455,I733486,I733531,I733592,I973360,I733618,I973366,I733635,I733643,I733660,I973363,I733677,I973342,I733694,I973345,I733711,I973351,I733728,I733759,I733776,I733807,I733824,I733841,I733872,I733912,I733920,I733937,I733954,I973354,I733971,I734002,I734019,I973348,I734036,I973357,I734062,I734084,I734101,I734132,I734177,I734238,I734264,I734281,I734289,I734306,I734323,I734340,I734357,I734374,I734405,I734422,I734453,I734470,I734487,I734518,I734558,I734566,I734583,I734600,I734617,I734648,I734665,I734682,I734708,I734730,I734747,I734778,I734823,I734884,I734910,I734927,I734935,I734952,I734969,I734986,I735003,I735020,I734870,I735051,I735068,I734873,I735099,I735116,I735133,I734849,I735164,I734861,I735204,I735212,I735229,I735246,I735263,I734876,I735294,I735311,I735328,I735354,I734864,I735376,I735393,I734858,I735424,I734852,I734855,I735469,I734867,I735530,I735556,I735573,I735581,I735598,I735615,I735632,I735649,I735666,I735697,I735714,I735745,I735762,I735779,I735810,I735850,I735858,I735875,I735892,I735909,I735940,I735957,I735974,I736000,I736022,I736039,I736070,I736115,I736176,I1054874,I736202,I1054898,I736219,I736227,I736244,I1054880,I736261,I1054889,I736278,I736295,I1054895,I736312,I736343,I736360,I736391,I736408,I1054892,I736425,I736456,I736496,I736504,I736521,I736538,I1054886,I736555,I736586,I1054877,I736603,I1054901,I736620,I1054883,I736646,I736668,I736685,I736716,I736761,I736822,I736848,I736865,I736873,I736890,I736907,I736924,I736941,I736958,I736989,I737006,I737037,I737054,I737071,I737102,I737142,I737150,I737167,I737184,I737201,I737232,I737249,I737266,I737292,I737314,I737331,I737362,I737407,I737468,I737494,I737511,I737519,I737536,I737553,I737570,I737587,I737604,I737635,I737652,I737683,I737700,I737717,I737748,I737788,I737796,I737813,I737830,I737847,I737878,I737895,I737912,I737938,I737960,I737977,I738008,I738053,I738114,I803512,I738140,I803515,I738157,I738165,I738182,I738199,I803524,I738216,I803533,I738233,I803521,I738250,I738281,I738298,I738329,I738346,I803527,I738363,I738394,I738434,I738442,I738459,I738476,I803518,I738493,I738524,I803530,I738541,I738558,I738584,I738606,I738623,I738654,I738699,I738760,I738786,I738803,I738811,I738828,I738845,I738862,I738879,I738896,I738927,I738944,I738975,I738992,I739009,I739040,I739080,I739088,I739105,I739122,I739139,I739170,I739187,I739204,I739230,I739252,I739269,I739300,I739345,I739406,I739432,I739449,I739457,I739474,I739491,I739508,I739525,I739542,I739573,I739590,I739621,I739638,I739655,I739686,I739726,I739734,I739751,I739768,I739785,I739816,I739833,I739850,I739876,I739898,I739915,I739946,I739991,I740052,I740078,I740095,I740103,I740120,I740137,I740154,I740171,I740188,I740038,I740219,I740236,I740041,I740267,I740284,I740301,I740017,I740332,I740029,I740372,I740380,I740397,I740414,I740431,I740044,I740462,I740479,I740496,I740522,I740032,I740544,I740561,I740026,I740592,I740020,I740023,I740637,I740035,I740698,I740724,I740741,I740749,I740766,I740783,I740800,I740817,I740834,I740865,I740882,I740913,I740930,I740947,I740978,I741018,I741026,I741043,I741060,I741077,I741108,I741125,I741142,I741168,I741190,I741207,I741238,I741283,I741344,I741370,I741387,I741395,I741412,I741429,I741446,I741463,I741480,I741511,I741528,I741559,I741576,I741593,I741624,I741664,I741672,I741689,I741706,I741723,I741754,I741771,I741788,I741814,I741836,I741853,I741884,I741929,I741990,I742016,I742033,I742041,I742058,I742075,I742092,I742109,I742126,I742157,I742174,I742205,I742222,I742239,I742270,I742310,I742318,I742335,I742352,I742369,I742400,I742417,I742434,I742460,I742482,I742499,I742530,I742575,I742636,I742662,I742679,I742687,I742704,I742721,I742738,I742755,I742772,I742622,I742803,I742820,I742625,I742851,I742868,I742885,I742601,I742916,I742613,I742956,I742964,I742981,I742998,I743015,I742628,I743046,I743063,I743080,I743106,I742616,I743128,I743145,I742610,I743176,I742604,I742607,I743221,I742619,I743282,I743308,I743325,I743333,I743350,I743367,I743384,I743401,I743418,I743268,I743449,I743466,I743271,I743497,I743514,I743531,I743247,I743562,I743259,I743602,I743610,I743627,I743644,I743661,I743274,I743692,I743709,I743726,I743752,I743262,I743774,I743791,I743256,I743822,I743250,I743253,I743867,I743265,I743928,I743954,I743971,I743979,I743996,I744013,I744030,I744047,I744064,I744095,I744112,I744143,I744160,I744177,I744208,I744248,I744256,I744273,I744290,I744307,I744338,I744355,I744372,I744398,I744420,I744437,I744468,I744513,I744574,I1061419,I744600,I1061443,I744617,I744625,I744642,I1061425,I744659,I1061434,I744676,I744693,I1061440,I744710,I744741,I744758,I744789,I744806,I1061437,I744823,I744854,I744894,I744902,I744919,I744936,I1061431,I744953,I744984,I1061422,I745001,I1061446,I745018,I1061428,I745044,I745066,I745083,I745114,I745159,I745220,I745246,I745263,I745271,I745288,I745305,I745322,I745339,I745356,I745206,I745387,I745404,I745209,I745435,I745452,I745469,I745185,I745500,I745197,I745540,I745548,I745565,I745582,I745599,I745212,I745630,I745647,I745664,I745690,I745200,I745712,I745729,I745194,I745760,I745188,I745191,I745805,I745203,I745866,I884858,I745892,I884840,I745909,I745917,I745934,I884849,I745951,I884861,I745968,I884843,I745985,I884852,I746002,I746033,I746050,I746081,I746098,I884864,I746115,I746146,I746186,I746194,I746211,I746228,I746245,I746276,I884846,I746293,I884855,I746310,I746336,I746358,I746375,I746406,I746451,I746512,I746538,I746555,I746563,I746580,I746597,I746614,I746631,I746648,I746679,I746696,I746727,I746744,I746761,I746792,I746832,I746840,I746857,I746874,I746891,I746922,I746939,I746956,I746982,I747004,I747021,I747052,I747097,I747158,I747184,I747201,I747209,I747226,I747243,I747260,I747277,I747294,I747325,I747342,I747373,I747390,I747407,I747438,I747478,I747486,I747503,I747520,I747537,I747568,I747585,I747602,I747628,I747650,I747667,I747698,I747743,I747804,I747830,I747847,I747855,I747872,I747889,I747906,I747923,I747940,I747971,I747988,I748019,I748036,I748053,I748084,I748124,I748132,I748149,I748166,I748183,I748214,I748231,I748248,I748274,I748296,I748313,I748344,I748389,I748450,I748476,I748493,I748501,I748518,I748535,I748552,I748569,I748586,I748617,I748634,I748665,I748682,I748699,I748730,I748770,I748778,I748795,I748812,I748829,I748860,I748877,I748894,I748920,I748942,I748959,I748990,I749035,I749096,I749122,I749139,I749147,I749164,I749181,I749198,I749215,I749232,I749263,I749280,I749311,I749328,I749345,I749376,I749416,I749424,I749441,I749458,I749475,I749506,I749523,I749540,I749566,I749588,I749605,I749636,I749681,I749742,I749768,I749785,I749793,I749810,I749827,I749844,I749861,I749878,I749909,I749926,I749957,I749974,I749991,I750022,I750062,I750070,I750087,I750104,I750121,I750152,I750169,I750186,I750212,I750234,I750251,I750282,I750327,I750388,I750414,I750431,I750439,I750456,I750473,I750490,I750507,I750524,I750555,I750572,I750603,I750620,I750637,I750668,I750708,I750716,I750733,I750750,I750767,I750798,I750815,I750832,I750858,I750880,I750897,I750928,I750973,I751034,I751060,I751077,I751085,I751102,I751119,I751136,I751153,I751170,I751020,I751201,I751218,I751023,I751249,I751266,I751283,I750999,I751314,I751011,I751354,I751362,I751379,I751396,I751413,I751026,I751444,I751461,I751478,I751504,I751014,I751526,I751543,I751008,I751574,I751002,I751005,I751619,I751017,I751680,I933410,I751706,I933392,I751723,I751731,I751748,I933401,I751765,I933413,I751782,I933395,I751799,I933404,I751816,I751847,I751864,I751895,I751912,I933416,I751929,I751960,I752000,I752008,I752025,I752042,I752059,I752090,I933398,I752107,I933407,I752124,I752150,I752172,I752189,I752220,I752265,I752326,I752352,I752369,I752377,I752394,I752411,I752428,I752445,I752462,I752493,I752510,I752541,I752558,I752575,I752606,I752646,I752654,I752671,I752688,I752705,I752736,I752753,I752770,I752796,I752818,I752835,I752866,I752911,I752972,I752998,I753015,I753023,I753040,I753057,I753074,I753091,I753108,I753139,I753156,I753187,I753204,I753221,I753252,I753292,I753300,I753317,I753334,I753351,I753382,I753399,I753416,I753442,I753464,I753481,I753512,I753557,I753618,I753644,I753661,I753669,I753686,I753703,I753720,I753737,I753754,I753785,I753802,I753833,I753850,I753867,I753898,I753938,I753946,I753963,I753980,I753997,I754028,I754045,I754062,I754088,I754110,I754127,I754158,I754203,I754264,I754290,I754307,I754315,I754332,I754349,I754366,I754383,I754400,I754431,I754448,I754479,I754496,I754513,I754544,I754584,I754592,I754609,I754626,I754643,I754674,I754691,I754708,I754734,I754756,I754773,I754804,I754849,I754910,I754936,I754953,I754961,I754978,I754995,I755012,I755029,I755046,I755077,I755094,I755125,I755142,I755159,I755190,I755230,I755238,I755255,I755272,I755289,I755320,I755337,I755354,I755380,I755402,I755419,I755450,I755495,I755556,I755582,I755599,I755607,I755624,I755641,I755658,I755675,I755692,I755723,I755740,I755771,I755788,I755805,I755836,I755876,I755884,I755901,I755918,I755935,I755966,I755983,I756000,I756026,I756048,I756065,I756096,I756141,I756202,I842664,I756228,I842646,I756245,I756253,I756270,I842655,I756287,I842667,I756304,I842649,I756321,I842658,I756338,I756188,I756369,I756386,I756191,I756417,I756434,I842670,I756451,I756167,I756482,I756179,I756522,I756530,I756547,I756564,I756581,I756194,I756612,I842652,I756629,I842661,I756646,I756672,I756182,I756694,I756711,I756176,I756742,I756170,I756173,I756787,I756185,I756848,I756874,I756891,I756899,I756916,I756933,I756950,I756967,I756984,I756834,I757015,I757032,I756837,I757063,I757080,I757097,I756813,I757128,I756825,I757168,I757176,I757193,I757210,I757227,I756840,I757258,I757275,I757292,I757318,I756828,I757340,I757357,I756822,I757388,I756816,I756819,I757433,I756831,I757494,I757520,I757537,I757545,I757562,I757579,I757596,I757613,I757630,I757661,I757678,I757709,I757726,I757743,I757774,I757814,I757822,I757839,I757856,I757873,I757904,I757921,I757938,I757964,I757986,I758003,I758034,I758079,I758140,I758166,I758183,I758191,I758208,I758225,I758242,I758259,I758276,I758307,I758324,I758355,I758372,I758389,I758420,I758460,I758468,I758485,I758502,I758519,I758550,I758567,I758584,I758610,I758632,I758649,I758680,I758725,I758786,I758812,I758829,I758837,I758854,I758871,I758888,I758905,I758922,I758953,I758970,I759001,I759018,I759035,I759066,I759106,I759114,I759131,I759148,I759165,I759196,I759213,I759230,I759256,I759278,I759295,I759326,I759371,I759432,I1031669,I759458,I1031693,I759475,I759483,I759500,I1031675,I759517,I1031684,I759534,I759551,I1031690,I759568,I759599,I759616,I759647,I759664,I1031687,I759681,I759712,I759752,I759760,I759777,I759794,I1031681,I759811,I759842,I1031672,I759859,I1031696,I759876,I1031678,I759902,I759924,I759941,I759972,I760017,I760078,I853646,I760104,I853628,I760121,I760129,I760146,I853637,I760163,I853649,I760180,I853631,I760197,I853640,I760214,I760245,I760262,I760293,I760310,I853652,I760327,I760358,I760398,I760406,I760423,I760440,I760457,I760488,I853634,I760505,I853643,I760522,I760548,I760570,I760587,I760618,I760663,I760724,I872720,I760750,I872702,I760767,I760775,I760792,I872711,I760809,I872723,I760826,I872705,I760843,I872714,I760860,I760891,I760908,I760939,I760956,I872726,I760973,I761004,I761044,I761052,I761069,I761086,I761103,I761134,I872708,I761151,I872717,I761168,I761194,I761216,I761233,I761264,I761309,I761370,I808561,I761396,I808564,I761413,I761421,I761438,I761455,I808573,I761472,I808582,I761489,I808570,I761506,I761356,I761537,I761554,I761359,I761585,I761602,I808576,I761619,I761335,I761650,I761347,I761690,I761698,I761715,I761732,I808567,I761749,I761362,I761780,I808579,I761797,I761814,I761840,I761350,I761862,I761879,I761344,I761910,I761338,I761341,I761955,I761353,I762016,I762042,I762059,I762067,I762084,I762101,I762118,I762135,I762152,I762002,I762183,I762200,I762005,I762231,I762248,I762265,I761981,I762296,I761993,I762336,I762344,I762361,I762378,I762395,I762008,I762426,I762443,I762460,I762486,I761996,I762508,I762525,I761990,I762556,I761984,I761987,I762601,I761999,I762662,I1031074,I762688,I1031098,I762705,I762713,I762730,I1031080,I762747,I1031089,I762764,I762781,I1031095,I762798,I762829,I762846,I762877,I762894,I1031092,I762911,I762942,I762982,I762990,I763007,I763024,I1031086,I763041,I763072,I1031077,I763089,I1031101,I763106,I1031083,I763132,I763154,I763171,I763202,I763247,I763308,I763334,I763351,I763359,I763376,I763393,I763410,I763427,I763444,I763294,I763475,I763492,I763297,I763523,I763540,I763557,I763273,I763588,I763285,I763628,I763636,I763653,I763670,I763687,I763300,I763718,I763735,I763752,I763778,I763288,I763800,I763817,I763282,I763848,I763276,I763279,I763893,I763291,I763954,I763980,I763997,I764005,I764022,I764039,I764056,I764073,I764090,I764121,I764138,I764169,I764186,I764203,I764234,I764274,I764282,I764299,I764316,I764333,I764364,I764381,I764398,I764424,I764446,I764463,I764494,I764539,I764600,I764626,I764643,I764651,I764668,I764685,I764702,I764719,I764736,I764767,I764784,I764815,I764832,I764849,I764880,I764920,I764928,I764945,I764962,I764979,I765010,I765027,I765044,I765070,I765092,I765109,I765140,I765185,I765246,I765272,I765289,I765297,I765314,I765331,I765348,I765365,I765382,I765232,I765413,I765430,I765235,I765461,I765478,I765495,I765211,I765526,I765223,I765566,I765574,I765591,I765608,I765625,I765238,I765656,I765673,I765690,I765716,I765226,I765738,I765755,I765220,I765786,I765214,I765217,I765831,I765229,I765892,I765918,I765935,I765943,I765960,I765977,I765994,I766011,I766028,I765878,I766059,I766076,I765881,I766107,I766124,I766141,I765857,I766172,I765869,I766212,I766220,I766237,I766254,I766271,I765884,I766302,I766319,I766336,I766362,I765872,I766384,I766401,I765866,I766432,I765860,I765863,I766477,I765875,I766538,I893528,I766564,I893510,I766581,I766589,I766606,I893519,I766623,I893531,I766640,I893513,I766657,I893522,I766674,I766705,I766722,I766753,I766770,I893534,I766787,I766818,I766858,I766866,I766883,I766900,I766917,I766948,I893516,I766965,I893525,I766982,I767008,I767030,I767047,I767078,I767123,I767184,I1071534,I767210,I1071558,I767227,I767235,I767252,I1071540,I767269,I1071549,I767286,I767303,I1071555,I767320,I767170,I767351,I767368,I767173,I767399,I767416,I1071552,I767433,I767149,I767464,I767161,I767504,I767512,I767529,I767546,I1071546,I767563,I767176,I767594,I1071537,I767611,I1071561,I767628,I1071543,I767654,I767164,I767676,I767693,I767158,I767724,I767152,I767155,I767769,I767167,I767830,I810805,I767856,I810808,I767873,I767881,I767898,I767915,I810817,I767932,I810826,I767949,I810814,I767966,I767997,I768014,I768045,I768062,I810820,I768079,I768110,I768150,I768158,I768175,I768192,I810811,I768209,I768240,I810823,I768257,I768274,I768300,I768322,I768339,I768370,I768415,I768476,I768502,I768519,I768527,I768544,I768561,I768578,I768595,I768612,I768462,I768643,I768660,I768465,I768691,I768708,I768725,I768441,I768756,I768453,I768796,I768804,I768821,I768838,I768855,I768468,I768886,I768903,I768920,I768946,I768456,I768968,I768985,I768450,I769016,I768444,I768447,I769061,I768459,I769122,I769148,I769165,I769173,I769190,I769207,I769224,I769241,I769258,I769289,I769306,I769337,I769354,I769371,I769402,I769442,I769450,I769467,I769484,I769501,I769532,I769549,I769566,I769592,I769614,I769631,I769662,I769707,I769768,I769794,I769811,I769819,I769836,I769853,I769870,I769887,I769904,I769754,I769935,I769952,I769757,I769983,I770000,I770017,I769733,I770048,I769745,I770088,I770096,I770113,I770130,I770147,I769760,I770178,I770195,I770212,I770238,I769748,I770260,I770277,I769742,I770308,I769736,I769739,I770353,I769751,I770414,I1072724,I770440,I1072748,I770457,I770465,I770482,I1072730,I770499,I1072739,I770516,I770533,I1072745,I770550,I770400,I770581,I770598,I770403,I770629,I770646,I1072742,I770663,I770379,I770694,I770391,I770734,I770742,I770759,I770776,I1072736,I770793,I770406,I770824,I1072727,I770841,I1072751,I770858,I1072733,I770884,I770394,I770906,I770923,I770388,I770954,I770382,I770385,I770999,I770397,I771060,I1019217,I771086,I1019211,I771103,I771111,I771128,I1019220,I771145,I1019232,I771162,I1019214,I771179,I771196,I771227,I771244,I771275,I771292,I1019208,I771309,I771340,I771380,I771388,I771405,I771422,I1019229,I771439,I771470,I1019223,I771487,I771504,I1019226,I771530,I771552,I771569,I771600,I771645,I771706,I771732,I771749,I771757,I771774,I771791,I771808,I771825,I771842,I771692,I771873,I771890,I771695,I771921,I771938,I771955,I771671,I771986,I771683,I772026,I772034,I772051,I772068,I772085,I771698,I772116,I772133,I772150,I772176,I771686,I772198,I772215,I771680,I772246,I771674,I771677,I772291,I771689,I772352,I772378,I772395,I772403,I772420,I772437,I772454,I772471,I772488,I772519,I772536,I772567,I772584,I772601,I772632,I772672,I772680,I772697,I772714,I772731,I772762,I772779,I772796,I772822,I772844,I772861,I772892,I772937,I772998,I1034049,I773024,I1034073,I773041,I773049,I773066,I1034055,I773083,I1034064,I773100,I773117,I1034070,I773134,I773165,I773182,I773213,I773230,I1034067,I773247,I773278,I773318,I773326,I773343,I773360,I1034061,I773377,I773408,I1034052,I773425,I1034076,I773442,I1034058,I773468,I773490,I773507,I773538,I773583,I773644,I773670,I773687,I773695,I773712,I773729,I773746,I773763,I773780,I773811,I773828,I773859,I773876,I773893,I773924,I773964,I773972,I773989,I774006,I774023,I774054,I774071,I774088,I774114,I774136,I774153,I774184,I774229,I774290,I774316,I774333,I774341,I774358,I774375,I774392,I774409,I774426,I774276,I774457,I774474,I774279,I774505,I774522,I774539,I774255,I774570,I774267,I774610,I774618,I774635,I774652,I774669,I774282,I774700,I774717,I774734,I774760,I774270,I774782,I774799,I774264,I774830,I774258,I774261,I774875,I774273,I774936,I1022079,I774962,I1022076,I774979,I774987,I775004,I1022073,I775021,I1022064,I775038,I1022085,I775055,I775072,I775103,I775120,I775151,I775168,I1022088,I775185,I775216,I775256,I775264,I775281,I775298,I1022067,I775315,I775346,I1022070,I775363,I1022091,I775380,I1022082,I775406,I775428,I775445,I775476,I775521,I775582,I929364,I775608,I929346,I775625,I775633,I775650,I929355,I775667,I929367,I775684,I929349,I775701,I929358,I775718,I775749,I775766,I775797,I775814,I929370,I775831,I775862,I775902,I775910,I775927,I775944,I775961,I775992,I929352,I776009,I929361,I776026,I776052,I776074,I776091,I776122,I776167,I776228,I776254,I776271,I776279,I776296,I776313,I776330,I776347,I776364,I776214,I776395,I776412,I776217,I776443,I776460,I776477,I776193,I776508,I776205,I776548,I776556,I776573,I776590,I776607,I776220,I776638,I776655,I776672,I776698,I776208,I776720,I776737,I776202,I776768,I776196,I776199,I776813,I776211,I776874,I776900,I776917,I776925,I776942,I776959,I776976,I776993,I777010,I777041,I777058,I777089,I777106,I777123,I777154,I777194,I777202,I777219,I777236,I777253,I777284,I777301,I777318,I777344,I777366,I777383,I777414,I777459,I777520,I777546,I777563,I777571,I777588,I777605,I777622,I777639,I777656,I777506,I777687,I777704,I777509,I777735,I777752,I777769,I777485,I777800,I777497,I777840,I777848,I777865,I777882,I777899,I777512,I777930,I777947,I777964,I777990,I777500,I778012,I778029,I777494,I778060,I777488,I777491,I778105,I777503,I778166,I1066179,I778192,I1066203,I778209,I778217,I778234,I1066185,I778251,I1066194,I778268,I778285,I1066200,I778302,I778333,I778350,I778381,I778398,I1066197,I778415,I778446,I778486,I778494,I778511,I778528,I1066191,I778545,I778576,I1066182,I778593,I1066206,I778610,I1066188,I778636,I778658,I778675,I778706,I778751,I778812,I947860,I778838,I947842,I778855,I778863,I778880,I947851,I778897,I947863,I778914,I947845,I778931,I947854,I778948,I778979,I778996,I779027,I779044,I947866,I779061,I779092,I779132,I779140,I779157,I779174,I779191,I779222,I947848,I779239,I947857,I779256,I779282,I779304,I779321,I779352,I779397,I779458,I886592,I779484,I886574,I779501,I779509,I779526,I886583,I779543,I886595,I779560,I886577,I779577,I886586,I779594,I779625,I779642,I779673,I779690,I886598,I779707,I779738,I779778,I779786,I779803,I779820,I779837,I779868,I886580,I779885,I886589,I779902,I779928,I779950,I779967,I779998,I780043,I780104,I780130,I780147,I780155,I780172,I780189,I780206,I780223,I780240,I780271,I780288,I780319,I780336,I780353,I780384,I780424,I780432,I780449,I780466,I780483,I780514,I780531,I780548,I780574,I780596,I780613,I780644,I780689,I780750,I891216,I780776,I891198,I780793,I780801,I780818,I891207,I780835,I891219,I780852,I891201,I780869,I891210,I780886,I780917,I780934,I780965,I780982,I891222,I780999,I781030,I781070,I781078,I781095,I781112,I781129,I781160,I891204,I781177,I891213,I781194,I781220,I781242,I781259,I781290,I781335,I781396,I781422,I781439,I781447,I781464,I781481,I781498,I781515,I781532,I781382,I781563,I781580,I781385,I781611,I781628,I781645,I781361,I781676,I781373,I781716,I781724,I781741,I781758,I781775,I781388,I781806,I781823,I781840,I781866,I781376,I781888,I781905,I781370,I781936,I781364,I781367,I781981,I781379,I782042,I853068,I782068,I853050,I782085,I782093,I782110,I853059,I782127,I853071,I782144,I853053,I782161,I853062,I782178,I782209,I782226,I782257,I782274,I853074,I782291,I782322,I782362,I782370,I782387,I782404,I782421,I782452,I853056,I782469,I853065,I782486,I782512,I782534,I782551,I782582,I782627,I782688,I873876,I782714,I873858,I782731,I782739,I782756,I873867,I782773,I873879,I782790,I873861,I782807,I873870,I782824,I782674,I782855,I782872,I782677,I782903,I782920,I873882,I782937,I782653,I782968,I782665,I783008,I783016,I783033,I783050,I783067,I782680,I783098,I873864,I783115,I873873,I783132,I783158,I782668,I783180,I783197,I782662,I783228,I782656,I782659,I783273,I782671,I783334,I783360,I783377,I783385,I783402,I783419,I783436,I783453,I783470,I783501,I783518,I783549,I783566,I783583,I783614,I783654,I783662,I783679,I783696,I783713,I783744,I783761,I783778,I783804,I783826,I783843,I783874,I783919,I783980,I784006,I784023,I784031,I784048,I784065,I784082,I784099,I784116,I784147,I784164,I784195,I784212,I784229,I784260,I784300,I784308,I784325,I784342,I784359,I784390,I784407,I784424,I784450,I784472,I784489,I784520,I784565,I784626,I940346,I784652,I940328,I784669,I784677,I784694,I940337,I784711,I940349,I784728,I940331,I784745,I940340,I784762,I784793,I784810,I784841,I784858,I940352,I784875,I784906,I784946,I784954,I784971,I784988,I785005,I785036,I940334,I785053,I940343,I785070,I785096,I785118,I785135,I785166,I785211,I785272,I785298,I785315,I785323,I785340,I785357,I785374,I785391,I785408,I785439,I785456,I785487,I785504,I785521,I785552,I785592,I785600,I785617,I785634,I785651,I785682,I785699,I785716,I785742,I785764,I785781,I785812,I785857,I785918,I785944,I785961,I785969,I785986,I786003,I786020,I786037,I786054,I786085,I786102,I786133,I786150,I786167,I786198,I786238,I786246,I786263,I786280,I786297,I786328,I786345,I786362,I786388,I786410,I786427,I786458,I786503,I786564,I786590,I786607,I786615,I786632,I786649,I786666,I786683,I786700,I786550,I786731,I786748,I786553,I786779,I786796,I786813,I786529,I786844,I786541,I786884,I786892,I786909,I786926,I786943,I786556,I786974,I786991,I787008,I787034,I786544,I787056,I787073,I786538,I787104,I786532,I786535,I787149,I786547,I787210,I787236,I787253,I787261,I787278,I787295,I787312,I787329,I787346,I787196,I787377,I787394,I787199,I787425,I787442,I787459,I787175,I787490,I787187,I787530,I787538,I787555,I787572,I787589,I787202,I787620,I787637,I787654,I787680,I787190,I787702,I787719,I787184,I787750,I787178,I787181,I787795,I787193,I787856,I787882,I787899,I787907,I787924,I787941,I787958,I787975,I787992,I788023,I788040,I788071,I788088,I788105,I788136,I788176,I788184,I788201,I788218,I788235,I788266,I788283,I788300,I788326,I788348,I788365,I788396,I788441,I788502,I927052,I788528,I927034,I788545,I788553,I788570,I927043,I788587,I927055,I788604,I927037,I788621,I927046,I788638,I788488,I788669,I788686,I788491,I788717,I788734,I927058,I788751,I788467,I788782,I788479,I788822,I788830,I788847,I788864,I788881,I788494,I788912,I927040,I788929,I927049,I788946,I788972,I788482,I788994,I789011,I788476,I789042,I788470,I788473,I789087,I788485,I789148,I1018061,I789174,I1018055,I789191,I789199,I789216,I1018064,I789233,I1018076,I789250,I1018058,I789267,I789284,I789315,I789332,I789363,I789380,I1018052,I789397,I789428,I789468,I789476,I789493,I789510,I1018073,I789527,I789558,I1018067,I789575,I789592,I1018070,I789618,I789640,I789657,I789688,I789733,I789794,I789820,I789837,I789845,I789862,I789879,I789896,I789913,I789930,I789961,I789978,I790009,I790026,I790043,I790074,I790114,I790122,I790139,I790156,I790173,I790204,I790221,I790238,I790264,I790286,I790303,I790334,I790379,I790440,I790466,I790483,I790491,I790508,I790525,I790542,I790559,I790576,I790426,I790607,I790624,I790429,I790655,I790672,I790689,I790405,I790720,I790417,I790760,I790768,I790785,I790802,I790819,I790432,I790850,I790867,I790884,I790910,I790420,I790932,I790949,I790414,I790980,I790408,I790411,I791025,I790423,I791086,I791112,I791129,I791137,I791154,I791171,I791188,I791205,I791222,I791253,I791270,I791301,I791318,I791335,I791366,I791406,I791414,I791431,I791448,I791465,I791496,I791513,I791530,I791556,I791578,I791595,I791626,I791671,I791732,I915492,I791758,I915474,I791775,I791783,I791800,I915483,I791817,I915495,I791834,I915477,I791851,I915486,I791868,I791899,I791916,I791947,I791964,I915498,I791981,I792012,I792052,I792060,I792077,I792094,I792111,I792142,I915480,I792159,I915489,I792176,I792202,I792224,I792241,I792272,I792317,I792378,I792404,I792421,I792429,I792446,I792463,I792480,I792497,I792514,I792545,I792562,I792593,I792610,I792627,I792658,I792698,I792706,I792723,I792740,I792757,I792788,I792805,I792822,I792848,I792870,I792887,I792918,I792963,I793024,I793050,I793067,I793075,I793092,I793109,I793126,I793143,I793160,I793191,I793208,I793239,I793256,I793273,I793304,I793344,I793352,I793369,I793386,I793403,I793434,I793451,I793468,I793494,I793516,I793533,I793564,I793609,I793670,I793696,I793713,I793721,I793738,I793755,I793772,I793789,I793806,I793656,I793837,I793854,I793659,I793885,I793902,I793919,I793635,I793950,I793647,I793990,I793998,I794015,I794032,I794049,I793662,I794080,I794097,I794114,I794140,I793650,I794162,I794179,I793644,I794210,I793638,I793641,I794255,I793653,I794316,I794342,I794359,I794367,I794384,I794401,I794418,I794435,I794452,I794302,I794483,I794500,I794305,I794531,I794548,I794565,I794281,I794596,I794293,I794636,I794644,I794661,I794678,I794695,I794308,I794726,I794743,I794760,I794786,I794296,I794808,I794825,I794290,I794856,I794284,I794287,I794901,I794299,I794962,I794988,I795005,I795013,I795030,I795047,I795064,I795081,I795098,I794948,I795129,I795146,I794951,I795177,I795194,I795211,I794927,I795242,I794939,I795282,I795290,I795307,I795324,I795341,I794954,I795372,I795389,I795406,I795432,I794942,I795454,I795471,I794936,I795502,I794930,I794933,I795547,I794945,I795608,I1091764,I795634,I1091788,I795651,I795659,I795676,I1091770,I795693,I1091779,I795710,I795727,I1091785,I795744,I795594,I795775,I795792,I795597,I795823,I795840,I1091782,I795857,I795573,I795888,I795585,I795928,I795936,I795953,I795970,I1091776,I795987,I795600,I796018,I1091767,I796035,I1091791,I796052,I1091773,I796078,I795588,I796100,I796117,I795582,I796148,I795576,I795579,I796193,I795591,I796248,I796274,I796291,I796313,I796339,I796347,I796364,I796381,I796398,I796415,I796432,I796449,I796480,I796511,I796528,I796545,I796562,I796593,I796638,I796655,I796672,I796698,I796706,I796737,I796754,I796809,I1008807,I796835,I796852,I796801,I796874,I1008804,I796900,I796908,I1008810,I796925,I796942,I1008819,I796959,I1008813,I796976,I796993,I1008825,I797010,I796783,I797041,I796786,I797072,I1008822,I797089,I797106,I797123,I796795,I797154,I796798,I796792,I797199,I1008816,I797216,I1008828,I797233,I797259,I797267,I796780,I797298,I797315,I796789,I797370,I839193,I797396,I797413,I797435,I839184,I797461,I797469,I839181,I797486,I797503,I839190,I797520,I839199,I797537,I797554,I839178,I797571,I797602,I797633,I839187,I797650,I797667,I797684,I797715,I797760,I839202,I797777,I797794,I839196,I797820,I797828,I797859,I797876,I797931,I797957,I797974,I797996,I798022,I798030,I798047,I798064,I798081,I798098,I798115,I798132,I798163,I798194,I798211,I798228,I798245,I798276,I798321,I798338,I798355,I798381,I798389,I798420,I798437,I798492,I798518,I798535,I798484,I798557,I798583,I798591,I798608,I798625,I798642,I798659,I798676,I798693,I798466,I798724,I798469,I798755,I798772,I798789,I798806,I798478,I798837,I798481,I798475,I798882,I798899,I798916,I798942,I798950,I798463,I798981,I798998,I798472,I799053,I799079,I799096,I799118,I799144,I799152,I799169,I799186,I799203,I799220,I799237,I799254,I799285,I799316,I799333,I799350,I799367,I799398,I799443,I799460,I799477,I799503,I799511,I799542,I799559,I799614,I979876,I799640,I799657,I799606,I799679,I979882,I799705,I799713,I979891,I799730,I799747,I979870,I799764,I979873,I799781,I799798,I979885,I799815,I799588,I799846,I799591,I799877,I979879,I799894,I799911,I799928,I799600,I799959,I799603,I799597,I800004,I979894,I800021,I800038,I979888,I800064,I800072,I799585,I800103,I800120,I799594,I800175,I800201,I800218,I800167,I800240,I800266,I800274,I800291,I800308,I800325,I800342,I800359,I800376,I800149,I800407,I800152,I800438,I800455,I800472,I800489,I800161,I800520,I800164,I800158,I800565,I800582,I800599,I800625,I800633,I800146,I800664,I800681,I800155,I800736,I800762,I800779,I800728,I800801,I800827,I800835,I800852,I800869,I800886,I800903,I800920,I800937,I800710,I800968,I800713,I800999,I801016,I801033,I801050,I800722,I801081,I800725,I800719,I801126,I801143,I801160,I801186,I801194,I800707,I801225,I801242,I800716,I801297,I1028817,I801323,I801340,I801289,I801362,I1028802,I801388,I801396,I1028811,I801413,I801430,I1028805,I801447,I1028823,I1028820,I801464,I801481,I1028796,I801498,I801271,I801529,I801274,I801560,I1028799,I801577,I801594,I801611,I801283,I801642,I801286,I801280,I801687,I801704,I1028814,I801721,I1028808,I801747,I801755,I801268,I801786,I801803,I801277,I801858,I801884,I801901,I801923,I801949,I801957,I801974,I801991,I802008,I802025,I802042,I802059,I802090,I802121,I802138,I802155,I802172,I802203,I802248,I802265,I802282,I802308,I802316,I802347,I802364,I802419,I802445,I802462,I802484,I802510,I802518,I802535,I802552,I802569,I802586,I802603,I802620,I802651,I802682,I802699,I802716,I802733,I802764,I802809,I802826,I802843,I802869,I802877,I802908,I802925,I802980,I803006,I803023,I803045,I803071,I803079,I803096,I803113,I803130,I803147,I803164,I803181,I803212,I803243,I803260,I803277,I803294,I803325,I803370,I803387,I803404,I803430,I803438,I803469,I803486,I803541,I1058459,I803567,I803584,I803606,I1058453,I803632,I803640,I1058444,I803657,I803674,I1058471,I803691,I1058456,I1058465,I803708,I803725,I1058450,I803742,I803773,I803804,I1058468,I803821,I803838,I803855,I803886,I803931,I1058462,I803948,I803965,I1058447,I803991,I803999,I804030,I804047,I804102,I996669,I804128,I804145,I804094,I804167,I996666,I804193,I804201,I996672,I804218,I804235,I996681,I804252,I996675,I804269,I804286,I996687,I804303,I804076,I804334,I804079,I804365,I996684,I804382,I804399,I804416,I804088,I804447,I804091,I804085,I804492,I996678,I804509,I996690,I804526,I804552,I804560,I804073,I804591,I804608,I804082,I804663,I804689,I804706,I804655,I804728,I804754,I804762,I804779,I804796,I804813,I804830,I804847,I804864,I804637,I804895,I804640,I804926,I804943,I804960,I804977,I804649,I805008,I804652,I804646,I805053,I805070,I805087,I805113,I805121,I804634,I805152,I805169,I804643,I805224,I805250,I805267,I805289,I805315,I805323,I805340,I805357,I805374,I805391,I805408,I805425,I805456,I805487,I805504,I805521,I805538,I805569,I805614,I805631,I805648,I805674,I805682,I805713,I805730,I805785,I805811,I805828,I805777,I805850,I805876,I805884,I805901,I805918,I805935,I805952,I805969,I805986,I805759,I806017,I805762,I806048,I806065,I806082,I806099,I805771,I806130,I805774,I805768,I806175,I806192,I806209,I806235,I806243,I805756,I806274,I806291,I805765,I806346,I806372,I806389,I806411,I806437,I806445,I806462,I806479,I806496,I806513,I806530,I806547,I806578,I806609,I806626,I806643,I806660,I806691,I806736,I806753,I806770,I806796,I806804,I806835,I806852,I806907,I806933,I806950,I806972,I806998,I807006,I807023,I807040,I807057,I807074,I807091,I807108,I807139,I807170,I807187,I807204,I807221,I807252,I807297,I807314,I807331,I807357,I807365,I807396,I807413,I807468,I918379,I807494,I807511,I807533,I918370,I807559,I807567,I918367,I807584,I807601,I918376,I807618,I918385,I807635,I807652,I918364,I807669,I807700,I807731,I918373,I807748,I807765,I807782,I807813,I807858,I918388,I807875,I807892,I918382,I807918,I807926,I807957,I807974,I808029,I808055,I808072,I808094,I808120,I808128,I808145,I808162,I808179,I808196,I808213,I808230,I808261,I808292,I808309,I808326,I808343,I808374,I808419,I808436,I808453,I808479,I808487,I808518,I808535,I808590,I1075119,I808616,I808633,I808655,I1075113,I808681,I808689,I1075104,I808706,I808723,I1075131,I808740,I1075116,I1075125,I808757,I808774,I1075110,I808791,I808822,I808853,I1075128,I808870,I808887,I808904,I808935,I808980,I1075122,I808997,I809014,I1075107,I809040,I809048,I809079,I809096,I809151,I921847,I809177,I809194,I809216,I921838,I809242,I809250,I921835,I809267,I809284,I921844,I809301,I921853,I809318,I809335,I921832,I809352,I809383,I809414,I921841,I809431,I809448,I809465,I809496,I809541,I921856,I809558,I809575,I921850,I809601,I809609,I809640,I809657,I809712,I809738,I809755,I809777,I809803,I809811,I809828,I809845,I809862,I809879,I809896,I809913,I809944,I809975,I809992,I810009,I810026,I810057,I810102,I810119,I810136,I810162,I810170,I810201,I810218,I810273,I810299,I810316,I810338,I810364,I810372,I810389,I810406,I810423,I810440,I810457,I810474,I810505,I810536,I810553,I810570,I810587,I810618,I810663,I810680,I810697,I810723,I810731,I810762,I810779,I810834,I810860,I810877,I810899,I810925,I810933,I810950,I810967,I810984,I811001,I811018,I811035,I811066,I811097,I811114,I811131,I811148,I811179,I811224,I811241,I811258,I811284,I811292,I811323,I811340,I811395,I811421,I811438,I811460,I811486,I811494,I811511,I811528,I811545,I811562,I811579,I811596,I811627,I811658,I811675,I811692,I811709,I811740,I811785,I811802,I811819,I811845,I811853,I811884,I811901,I811956,I811982,I811999,I812021,I812047,I812055,I812072,I812089,I812106,I812123,I812140,I812157,I812188,I812219,I812236,I812253,I812270,I812301,I812346,I812363,I812380,I812406,I812414,I812445,I812462,I812517,I963012,I812543,I812560,I812509,I812582,I963018,I812608,I812616,I963027,I812633,I812650,I963006,I812667,I963009,I812684,I812701,I963021,I812718,I812491,I812749,I812494,I812780,I963015,I812797,I812814,I812831,I812503,I812862,I812506,I812500,I812907,I963030,I812924,I812941,I963024,I812967,I812975,I812488,I813006,I813023,I812497,I813078,I813104,I813121,I813143,I813169,I813177,I813194,I813211,I813228,I813245,I813262,I813279,I813310,I813341,I813358,I813375,I813392,I813423,I813468,I813485,I813502,I813528,I813536,I813567,I813584,I813639,I1065004,I813665,I813682,I813704,I1064998,I813730,I813738,I1064989,I813755,I813772,I1065016,I813789,I1065001,I1065010,I813806,I813823,I1064995,I813840,I813871,I813902,I1065013,I813919,I813936,I813953,I813984,I814029,I1065007,I814046,I814063,I1064992,I814089,I814097,I814128,I814145,I814200,I814226,I814243,I814265,I814291,I814299,I814316,I814333,I814350,I814367,I814384,I814401,I814432,I814463,I814480,I814497,I814514,I814545,I814590,I814607,I814624,I814650,I814658,I814689,I814706,I814761,I814787,I814804,I814753,I814826,I814852,I814860,I814877,I814894,I814911,I814928,I814945,I814962,I814735,I814993,I814738,I815024,I815041,I815058,I815075,I814747,I815106,I814750,I814744,I815151,I815168,I815185,I815211,I815219,I814732,I815250,I815267,I814741,I815322,I815348,I815365,I815314,I815387,I815413,I815421,I815438,I815455,I815472,I815489,I815506,I815523,I815296,I815554,I815299,I815585,I815602,I815619,I815636,I815308,I815667,I815311,I815305,I815712,I815729,I815746,I815772,I815780,I815293,I815811,I815828,I815302,I815883,I1046559,I815909,I815926,I815875,I815948,I1046553,I815974,I815982,I1046544,I815999,I816016,I1046571,I816033,I1046556,I1046565,I816050,I816067,I1046550,I816084,I815857,I816115,I815860,I816146,I1046568,I816163,I816180,I816197,I815869,I816228,I815872,I815866,I816273,I1046562,I816290,I816307,I1046547,I816333,I816341,I815854,I816372,I816389,I815863,I816444,I816470,I816487,I816509,I816535,I816543,I816560,I816577,I816594,I816611,I816628,I816645,I816676,I816707,I816724,I816741,I816758,I816789,I816834,I816851,I816868,I816894,I816902,I816933,I816950,I817005,I817031,I817048,I817070,I817096,I817104,I817121,I817138,I817155,I817172,I817189,I817206,I817237,I817268,I817285,I817302,I817319,I817350,I817395,I817412,I817429,I817455,I817463,I817494,I817511,I817566,I817592,I817609,I817631,I817657,I817665,I817682,I817699,I817716,I817733,I817750,I817767,I817798,I817829,I817846,I817863,I817880,I817911,I817956,I817973,I817990,I818016,I818024,I818055,I818072,I818127,I901617,I818153,I818170,I818192,I901608,I818218,I818226,I901605,I818243,I818260,I901614,I818277,I901623,I818294,I818311,I901602,I818328,I818359,I818390,I901611,I818407,I818424,I818441,I818472,I818517,I901626,I818534,I818551,I901620,I818577,I818585,I818616,I818633,I818688,I818714,I818731,I818753,I818779,I818787,I818804,I818821,I818838,I818855,I818872,I818889,I818920,I818951,I818968,I818985,I819002,I819033,I819078,I819095,I819112,I819138,I819146,I819177,I819194,I819249,I831679,I819275,I819292,I819314,I831670,I819340,I819348,I831667,I819365,I819382,I831676,I819399,I831685,I819416,I819433,I831664,I819450,I819481,I819512,I831673,I819529,I819546,I819563,I819594,I819639,I831688,I819656,I819673,I831682,I819699,I819707,I819738,I819755,I819810,I819836,I819853,I819875,I819901,I819909,I819926,I819943,I819960,I819977,I819994,I820011,I820042,I820073,I820090,I820107,I820124,I820155,I820200,I820217,I820234,I820260,I820268,I820299,I820316,I820371,I820397,I820414,I820436,I820462,I820470,I820487,I820504,I820521,I820538,I820555,I820572,I820603,I820634,I820651,I820668,I820685,I820716,I820761,I820778,I820795,I820821,I820829,I820860,I820877,I820932,I820958,I820975,I820997,I821023,I821031,I821048,I821065,I821082,I821099,I821116,I821133,I821164,I821195,I821212,I821229,I821246,I821277,I821322,I821339,I821356,I821382,I821390,I821421,I821438,I821493,I943811,I821519,I821536,I821485,I821558,I943802,I821584,I821592,I943799,I821609,I821626,I943808,I821643,I943817,I821660,I821677,I943796,I821694,I821467,I821725,I821470,I821756,I943805,I821773,I821790,I821807,I821479,I821838,I821482,I821476,I821883,I943820,I821900,I821917,I943814,I821943,I821951,I821464,I821982,I821999,I821473,I822054,I822080,I822097,I822119,I822145,I822153,I822170,I822187,I822204,I822221,I822238,I822255,I822286,I822317,I822334,I822351,I822368,I822399,I822444,I822461,I822478,I822504,I822512,I822543,I822560,I822615,I822641,I822658,I822680,I822706,I822714,I822731,I822748,I822765,I822782,I822799,I822816,I822847,I822878,I822895,I822912,I822929,I822960,I823005,I823022,I823039,I823065,I823073,I823104,I823121,I823176,I823202,I823219,I823241,I823267,I823275,I823292,I823309,I823326,I823343,I823360,I823377,I823408,I823439,I823456,I823473,I823490,I823521,I823566,I823583,I823600,I823626,I823634,I823665,I823682,I823737,I823763,I823780,I823802,I823828,I823836,I823853,I823870,I823887,I823904,I823921,I823938,I823969,I824000,I824017,I824034,I824051,I824082,I824127,I824144,I824161,I824187,I824195,I824226,I824243,I824298,I824324,I824341,I824363,I824389,I824397,I824414,I824431,I824448,I824465,I824482,I824499,I824530,I824561,I824578,I824595,I824612,I824643,I824688,I824705,I824722,I824748,I824756,I824787,I824804,I824859,I824885,I824902,I824851,I824924,I824950,I824958,I824975,I824992,I825009,I825026,I825043,I825060,I824833,I825091,I824836,I825122,I825139,I825156,I825173,I824845,I825204,I824848,I824842,I825249,I825266,I825283,I825309,I825317,I824830,I825348,I825365,I824839,I825420,I1070954,I825446,I825463,I825485,I1070948,I825511,I825519,I1070939,I825536,I825553,I1070966,I825570,I1070951,I1070960,I825587,I825604,I1070945,I825621,I825652,I825683,I1070963,I825700,I825717,I825734,I825765,I825810,I1070957,I825827,I825844,I1070942,I825870,I825878,I825909,I825926,I825981,I1024890,I826007,I826024,I826046,I1024875,I826072,I826080,I1024884,I826097,I826114,I1024878,I826131,I1024896,I1024893,I826148,I826165,I1024869,I826182,I826213,I826244,I1024872,I826261,I826278,I826295,I826326,I826371,I826388,I1024887,I826405,I1024881,I826431,I826439,I826470,I826487,I826542,I1005917,I826568,I826585,I826534,I826607,I1005914,I826633,I826641,I1005920,I826658,I826675,I1005929,I826692,I1005923,I826709,I826726,I1005935,I826743,I826516,I826774,I826519,I826805,I1005932,I826822,I826839,I826856,I826528,I826887,I826531,I826525,I826932,I1005926,I826949,I1005938,I826966,I826992,I827000,I826513,I827031,I827048,I826522,I827103,I827129,I827146,I827168,I827194,I827202,I827219,I827236,I827253,I827270,I827287,I827304,I827335,I827366,I827383,I827400,I827417,I827448,I827493,I827510,I827527,I827553,I827561,I827592,I827609,I827664,I833413,I827690,I827707,I827729,I833404,I827755,I827763,I833401,I827780,I827797,I833410,I827814,I833419,I827831,I827848,I833398,I827865,I827896,I827927,I833407,I827944,I827961,I827978,I828009,I828054,I833422,I828071,I828088,I833416,I828114,I828122,I828153,I828170,I828228,I828254,I828262,I828302,I828310,I828327,I828344,I828384,I828406,I828423,I828449,I828457,I828474,I828491,I828508,I828525,I828570,I828601,I828618,I828644,I828652,I828683,I828700,I828717,I828734,I828806,I828832,I828840,I828880,I828888,I828905,I828922,I828962,I828984,I829001,I829027,I829035,I829052,I829069,I829086,I829103,I829148,I829179,I829196,I829222,I829230,I829261,I829278,I829295,I829312,I829384,I829410,I829418,I829458,I829466,I829483,I829500,I829540,I829562,I829579,I829605,I829613,I829630,I829647,I829664,I829681,I829726,I829757,I829774,I829800,I829808,I829839,I829856,I829873,I829890,I829962,I829988,I829996,I830036,I830044,I830061,I830078,I830118,I830140,I830157,I830183,I830191,I830208,I830225,I830242,I830259,I830304,I830335,I830352,I830378,I830386,I830417,I830434,I830451,I830468,I830540,I965203,I830566,I830574,I965197,I965182,I830614,I830622,I965188,I830639,I965200,I830656,I830696,I830718,I830735,I830761,I830769,I830786,I965206,I830803,I965194,I830820,I830837,I830882,I965185,I830913,I830930,I965191,I830956,I830964,I830995,I831012,I831029,I831046,I831118,I831144,I831152,I831192,I831200,I831217,I831234,I831274,I831296,I831313,I831339,I831347,I831364,I831381,I831398,I831415,I831460,I831491,I831508,I831534,I831542,I831573,I831590,I831607,I831624,I831696,I831722,I831730,I831770,I831778,I831795,I831812,I831852,I831874,I831891,I831917,I831925,I831942,I831959,I831976,I831993,I832038,I832069,I832086,I832112,I832120,I832151,I832168,I832185,I832202,I832274,I832300,I832308,I832348,I832356,I832373,I832390,I832430,I832452,I832469,I832495,I832503,I832520,I832537,I832554,I832571,I832616,I832647,I832664,I832690,I832698,I832729,I832746,I832763,I832780,I832852,I832878,I832886,I832926,I832934,I832951,I832968,I833008,I833030,I833047,I833073,I833081,I833098,I833115,I833132,I833149,I833194,I833225,I833242,I833268,I833276,I833307,I833324,I833341,I833358,I833430,I833456,I833464,I833504,I833512,I833529,I833546,I833586,I833608,I833625,I833651,I833659,I833676,I833693,I833710,I833727,I833772,I833803,I833820,I833846,I833854,I833885,I833902,I833919,I833936,I834008,I834034,I834042,I834082,I834090,I834107,I834124,I834164,I834186,I834203,I834229,I834237,I834254,I834271,I834288,I834305,I834350,I834381,I834398,I834424,I834432,I834463,I834480,I834497,I834514,I834586,I834612,I834620,I834660,I834668,I834685,I834702,I834742,I834764,I834781,I834807,I834815,I834832,I834849,I834866,I834883,I834928,I834959,I834976,I835002,I835010,I835041,I835058,I835075,I835092,I835164,I835190,I835198,I835238,I835246,I835263,I835280,I835320,I835342,I835359,I835385,I835393,I835410,I835427,I835444,I835461,I835506,I835537,I835554,I835580,I835588,I835619,I835636,I835653,I835670,I835742,I985875,I835768,I835776,I985869,I985854,I835816,I835824,I985860,I835841,I985872,I835858,I835898,I835920,I835937,I835963,I835971,I835988,I985878,I836005,I985866,I836022,I836039,I836084,I985857,I836115,I836132,I985863,I836158,I836166,I836197,I836214,I836231,I836248,I836320,I836346,I836354,I836394,I836402,I836419,I836436,I836476,I836498,I836515,I836541,I836549,I836566,I836583,I836600,I836617,I836662,I836693,I836710,I836736,I836744,I836775,I836792,I836809,I836826,I836898,I836924,I836932,I836972,I836980,I836997,I837014,I837054,I837076,I837093,I837119,I837127,I837144,I837161,I837178,I837195,I837240,I837271,I837288,I837314,I837322,I837353,I837370,I837387,I837404,I837476,I837502,I837510,I837550,I837558,I837575,I837592,I837632,I837654,I837671,I837697,I837705,I837722,I837739,I837756,I837773,I837818,I837849,I837866,I837892,I837900,I837931,I837948,I837965,I837982,I838054,I838080,I838088,I838128,I838136,I838153,I838170,I838210,I838232,I838249,I838275,I838283,I838300,I838317,I838334,I838351,I838396,I838427,I838444,I838470,I838478,I838509,I838526,I838543,I838560,I838632,I838658,I838666,I838706,I838714,I838731,I838748,I838788,I838810,I838827,I838853,I838861,I838878,I838895,I838912,I838929,I838974,I839005,I839022,I839048,I839056,I839087,I839104,I839121,I839138,I839210,I839236,I839244,I839284,I839292,I839309,I839326,I839366,I839388,I839405,I839431,I839439,I839456,I839473,I839490,I839507,I839552,I839583,I839600,I839626,I839634,I839665,I839682,I839699,I839716,I839788,I839814,I839822,I839771,I839862,I839870,I839887,I839904,I839759,I839944,I839780,I839966,I839983,I840009,I840017,I840034,I840051,I840068,I840085,I839756,I839777,I840130,I839768,I840161,I840178,I840204,I840212,I839774,I840243,I840260,I840277,I840294,I839765,I839762,I840366,I840392,I840400,I840440,I840448,I840465,I840482,I840522,I840544,I840561,I840587,I840595,I840612,I840629,I840646,I840663,I840708,I840739,I840756,I840782,I840790,I840821,I840838,I840855,I840872,I840944,I840970,I840978,I841018,I841026,I841043,I841060,I841100,I841122,I841139,I841165,I841173,I841190,I841207,I841224,I841241,I841286,I841317,I841334,I841360,I841368,I841399,I841416,I841433,I841450,I841522,I841548,I841556,I841596,I841604,I841621,I841638,I841678,I841700,I841717,I841743,I841751,I841768,I841785,I841802,I841819,I841864,I841895,I841912,I841938,I841946,I841977,I841994,I842011,I842028,I842100,I842126,I842134,I842174,I842182,I842199,I842216,I842256,I842278,I842295,I842321,I842329,I842346,I842363,I842380,I842397,I842442,I842473,I842490,I842516,I842524,I842555,I842572,I842589,I842606,I842678,I842704,I842712,I842752,I842760,I842777,I842794,I842834,I842856,I842873,I842899,I842907,I842924,I842941,I842958,I842975,I843020,I843051,I843068,I843094,I843102,I843133,I843150,I843167,I843184,I843256,I843282,I843290,I843330,I843338,I843355,I843372,I843412,I843434,I843451,I843477,I843485,I843502,I843519,I843536,I843553,I843598,I843629,I843646,I843672,I843680,I843711,I843728,I843745,I843762,I843834,I843860,I843868,I843908,I843916,I843933,I843950,I843990,I844012,I844029,I844055,I844063,I844080,I844097,I844114,I844131,I844176,I844207,I844224,I844250,I844258,I844289,I844306,I844323,I844340,I844412,I844438,I844446,I844486,I844494,I844511,I844528,I844568,I844590,I844607,I844633,I844641,I844658,I844675,I844692,I844709,I844754,I844785,I844802,I844828,I844836,I844867,I844884,I844901,I844918,I844990,I845016,I845024,I845064,I845072,I845089,I845106,I845146,I845168,I845185,I845211,I845219,I845236,I845253,I845270,I845287,I845332,I845363,I845380,I845406,I845414,I845445,I845462,I845479,I845496,I845568,I845594,I845602,I845642,I845650,I845667,I845684,I845724,I845746,I845763,I845789,I845797,I845814,I845831,I845848,I845865,I845910,I845941,I845958,I845984,I845992,I846023,I846040,I846057,I846074,I846146,I846172,I846180,I846220,I846228,I846245,I846262,I846302,I846324,I846341,I846367,I846375,I846392,I846409,I846426,I846443,I846488,I846519,I846536,I846562,I846570,I846601,I846618,I846635,I846652,I846724,I846750,I846758,I846707,I846798,I846806,I846823,I846840,I846695,I846880,I846716,I846902,I846919,I846945,I846953,I846970,I846987,I847004,I847021,I846692,I846713,I847066,I846704,I847097,I847114,I847140,I847148,I846710,I847179,I847196,I847213,I847230,I846701,I846698,I847302,I847328,I847336,I847376,I847384,I847401,I847418,I847458,I847480,I847497,I847523,I847531,I847548,I847565,I847582,I847599,I847644,I847675,I847692,I847718,I847726,I847757,I847774,I847791,I847808,I847880,I847906,I847914,I847954,I847962,I847979,I847996,I848036,I848058,I848075,I848101,I848109,I848126,I848143,I848160,I848177,I848222,I848253,I848270,I848296,I848304,I848335,I848352,I848369,I848386,I848458,I1062041,I848484,I848492,I1062023,I1062014,I848532,I848540,I1062029,I848557,I1062017,I848574,I848614,I848636,I1062026,I848653,I848679,I848687,I848704,I1062035,I848721,I848738,I848755,I848800,I1062038,I848831,I848848,I1062032,I1062020,I848874,I848882,I848913,I848930,I848947,I848964,I849036,I970643,I849062,I849070,I970637,I970622,I849110,I849118,I970628,I849135,I970640,I849152,I849192,I849214,I849231,I849257,I849265,I849282,I970646,I849299,I970634,I849316,I849333,I849378,I970625,I849409,I849426,I970631,I849452,I849460,I849491,I849508,I849525,I849542,I849614,I976627,I849640,I849648,I976621,I976606,I849688,I849696,I976612,I849713,I976624,I849730,I849770,I849792,I849809,I849835,I849843,I849860,I976630,I849877,I976618,I849894,I849911,I849956,I976609,I849987,I850004,I976615,I850030,I850038,I850069,I850086,I850103,I850120,I850192,I850218,I850226,I850266,I850274,I850291,I850308,I850348,I850370,I850387,I850413,I850421,I850438,I850455,I850472,I850489,I850534,I850565,I850582,I850608,I850616,I850647,I850664,I850681,I850698,I850770,I850796,I850804,I850844,I850852,I850869,I850886,I850926,I850948,I850965,I850991,I850999,I851016,I851033,I851050,I851067,I851112,I851143,I851160,I851186,I851194,I851225,I851242,I851259,I851276,I851348,I851374,I851382,I851422,I851430,I851447,I851464,I851504,I851526,I851543,I851569,I851577,I851594,I851611,I851628,I851645,I851690,I851721,I851738,I851764,I851772,I851803,I851820,I851837,I851854,I851926,I851952,I851960,I852000,I852008,I852025,I852042,I852082,I852104,I852121,I852147,I852155,I852172,I852189,I852206,I852223,I852268,I852299,I852316,I852342,I852350,I852381,I852398,I852415,I852432,I852504,I852530,I852538,I852578,I852586,I852603,I852620,I852660,I852682,I852699,I852725,I852733,I852750,I852767,I852784,I852801,I852846,I852877,I852894,I852920,I852928,I852959,I852976,I852993,I853010,I853082,I853108,I853116,I853156,I853164,I853181,I853198,I853238,I853260,I853277,I853303,I853311,I853328,I853345,I853362,I853379,I853424,I853455,I853472,I853498,I853506,I853537,I853554,I853571,I853588,I853660,I853686,I853694,I853734,I853742,I853759,I853776,I853816,I853838,I853855,I853881,I853889,I853906,I853923,I853940,I853957,I854002,I854033,I854050,I854076,I854084,I854115,I854132,I854149,I854166,I854238,I854264,I854272,I854312,I854320,I854337,I854354,I854394,I854416,I854433,I854459,I854467,I854484,I854501,I854518,I854535,I854580,I854611,I854628,I854654,I854662,I854693,I854710,I854727,I854744,I854816,I854842,I854850,I854890,I854898,I854915,I854932,I854972,I854994,I855011,I855037,I855045,I855062,I855079,I855096,I855113,I855158,I855189,I855206,I855232,I855240,I855271,I855288,I855305,I855322,I855394,I855420,I855428,I855468,I855476,I855493,I855510,I855550,I855572,I855589,I855615,I855623,I855640,I855657,I855674,I855691,I855736,I855767,I855784,I855810,I855818,I855849,I855866,I855883,I855900,I855972,I855998,I856006,I856046,I856054,I856071,I856088,I856128,I856150,I856167,I856193,I856201,I856218,I856235,I856252,I856269,I856314,I856345,I856362,I856388,I856396,I856427,I856444,I856461,I856478,I856550,I856576,I856584,I856624,I856632,I856649,I856666,I856706,I856728,I856745,I856771,I856779,I856796,I856813,I856830,I856847,I856892,I856923,I856940,I856966,I856974,I857005,I857022,I857039,I857056,I857128,I857154,I857162,I857202,I857210,I857227,I857244,I857284,I857306,I857323,I857349,I857357,I857374,I857391,I857408,I857425,I857470,I857501,I857518,I857544,I857552,I857583,I857600,I857617,I857634,I857706,I857732,I857740,I857780,I857788,I857805,I857822,I857862,I857884,I857901,I857927,I857935,I857952,I857969,I857986,I858003,I858048,I858079,I858096,I858122,I858130,I858161,I858178,I858195,I858212,I858284,I858310,I858318,I858358,I858366,I858383,I858400,I858440,I858462,I858479,I858505,I858513,I858530,I858547,I858564,I858581,I858626,I858657,I858674,I858700,I858708,I858739,I858756,I858773,I858790,I858862,I858888,I858896,I858936,I858944,I858961,I858978,I859018,I859040,I859057,I859083,I859091,I859108,I859125,I859142,I859159,I859204,I859235,I859252,I859278,I859286,I859317,I859334,I859351,I859368,I859440,I859466,I859474,I859514,I859522,I859539,I859556,I859596,I859618,I859635,I859661,I859669,I859686,I859703,I859720,I859737,I859782,I859813,I859830,I859856,I859864,I859895,I859912,I859929,I859946,I860018,I860044,I860052,I860092,I860100,I860117,I860134,I860174,I860196,I860213,I860239,I860247,I860264,I860281,I860298,I860315,I860360,I860391,I860408,I860434,I860442,I860473,I860490,I860507,I860524,I860596,I860622,I860630,I860670,I860678,I860695,I860712,I860752,I860774,I860791,I860817,I860825,I860842,I860859,I860876,I860893,I860938,I860969,I860986,I861012,I861020,I861051,I861068,I861085,I861102,I861174,I861200,I861208,I861248,I861256,I861273,I861290,I861330,I861352,I861369,I861395,I861403,I861420,I861437,I861454,I861471,I861516,I861547,I861564,I861590,I861598,I861629,I861646,I861663,I861680,I861752,I861778,I861786,I861826,I861834,I861851,I861868,I861908,I861930,I861947,I861973,I861981,I861998,I862015,I862032,I862049,I862094,I862125,I862142,I862168,I862176,I862207,I862224,I862241,I862258,I862330,I862356,I862364,I862404,I862412,I862429,I862446,I862486,I862508,I862525,I862551,I862559,I862576,I862593,I862610,I862627,I862672,I862703,I862720,I862746,I862754,I862785,I862802,I862819,I862836,I862908,I862934,I862942,I862891,I862982,I862990,I863007,I863024,I862879,I863064,I862900,I863086,I863103,I863129,I863137,I863154,I863171,I863188,I863205,I862876,I862897,I863250,I862888,I863281,I863298,I863324,I863332,I862894,I863363,I863380,I863397,I863414,I862885,I862882,I863486,I863512,I863520,I863560,I863568,I863585,I863602,I863642,I863664,I863681,I863707,I863715,I863732,I863749,I863766,I863783,I863828,I863859,I863876,I863902,I863910,I863941,I863958,I863975,I863992,I864064,I864090,I864098,I864138,I864146,I864163,I864180,I864220,I864242,I864259,I864285,I864293,I864310,I864327,I864344,I864361,I864406,I864437,I864454,I864480,I864488,I864519,I864536,I864553,I864570,I864642,I864668,I864676,I864716,I864724,I864741,I864758,I864798,I864820,I864837,I864863,I864871,I864888,I864905,I864922,I864939,I864984,I865015,I865032,I865058,I865066,I865097,I865114,I865131,I865148,I865220,I865246,I865254,I865203,I865294,I865302,I865319,I865336,I865191,I865376,I865212,I865398,I865415,I865441,I865449,I865466,I865483,I865500,I865517,I865188,I865209,I865562,I865200,I865593,I865610,I865636,I865644,I865206,I865675,I865692,I865709,I865726,I865197,I865194,I865798,I865824,I865832,I865872,I865880,I865897,I865914,I865954,I865976,I865993,I866019,I866027,I866044,I866061,I866078,I866095,I866140,I866171,I866188,I866214,I866222,I866253,I866270,I866287,I866304,I866376,I866402,I866410,I866450,I866458,I866475,I866492,I866532,I866554,I866571,I866597,I866605,I866622,I866639,I866656,I866673,I866718,I866749,I866766,I866792,I866800,I866831,I866848,I866865,I866882,I866954,I866980,I866988,I867028,I867036,I867053,I867070,I867110,I867132,I867149,I867175,I867183,I867200,I867217,I867234,I867251,I867296,I867327,I867344,I867370,I867378,I867409,I867426,I867443,I867460,I867532,I1067396,I867558,I867566,I1067378,I1067369,I867606,I867614,I1067384,I867631,I1067372,I867648,I867688,I867710,I1067381,I867727,I867753,I867761,I867778,I1067390,I867795,I867812,I867829,I867874,I1067393,I867905,I867922,I1067387,I1067375,I867948,I867956,I867987,I868004,I868021,I868038,I868110,I868136,I868144,I868184,I868192,I868209,I868226,I868266,I868288,I868305,I868331,I868339,I868356,I868373,I868390,I868407,I868452,I868483,I868500,I868526,I868534,I868565,I868582,I868599,I868616,I868688,I868714,I868722,I868671,I868762,I868770,I868787,I868804,I868659,I868844,I868680,I868866,I868883,I868909,I868917,I868934,I868951,I868968,I868985,I868656,I868677,I869030,I868668,I869061,I869078,I869104,I869112,I868674,I869143,I869160,I869177,I869194,I868665,I868662,I869266,I869292,I869300,I869340,I869348,I869365,I869382,I869422,I869444,I869461,I869487,I869495,I869512,I869529,I869546,I869563,I869608,I869639,I869656,I869682,I869690,I869721,I869738,I869755,I869772,I869844,I869870,I869878,I869918,I869926,I869943,I869960,I870000,I870022,I870039,I870065,I870073,I870090,I870107,I870124,I870141,I870186,I870217,I870234,I870260,I870268,I870299,I870316,I870333,I870350,I870422,I870448,I870456,I870496,I870504,I870521,I870538,I870578,I870600,I870617,I870643,I870651,I870668,I870685,I870702,I870719,I870764,I870795,I870812,I870838,I870846,I870877,I870894,I870911,I870928,I871000,I871026,I871034,I870983,I871074,I871082,I871099,I871116,I870971,I871156,I870992,I871178,I871195,I871221,I871229,I871246,I871263,I871280,I871297,I870968,I870989,I871342,I870980,I871373,I871390,I871416,I871424,I870986,I871455,I871472,I871489,I871506,I870977,I870974,I871578,I871604,I871612,I871652,I871660,I871677,I871694,I871734,I871756,I871773,I871799,I871807,I871824,I871841,I871858,I871875,I871920,I871951,I871968,I871994,I872002,I872033,I872050,I872067,I872084,I872156,I872182,I872190,I872230,I872238,I872255,I872272,I872312,I872334,I872351,I872377,I872385,I872402,I872419,I872436,I872453,I872498,I872529,I872546,I872572,I872580,I872611,I872628,I872645,I872662,I872734,I872760,I872768,I872808,I872816,I872833,I872850,I872890,I872912,I872929,I872955,I872963,I872980,I872997,I873014,I873031,I873076,I873107,I873124,I873150,I873158,I873189,I873206,I873223,I873240,I873312,I873338,I873346,I873386,I873394,I873411,I873428,I873468,I873490,I873507,I873533,I873541,I873558,I873575,I873592,I873609,I873654,I873685,I873702,I873728,I873736,I873767,I873784,I873801,I873818,I873890,I873916,I873924,I873964,I873972,I873989,I874006,I874046,I874068,I874085,I874111,I874119,I874136,I874153,I874170,I874187,I874232,I874263,I874280,I874306,I874314,I874345,I874362,I874379,I874396,I874468,I874494,I874502,I874542,I874550,I874567,I874584,I874624,I874646,I874663,I874689,I874697,I874714,I874731,I874748,I874765,I874810,I874841,I874858,I874884,I874892,I874923,I874940,I874957,I874974,I875046,I999580,I875072,I875080,I999562,I999571,I875120,I875128,I999556,I875145,I999568,I875162,I875202,I875224,I999559,I875241,I875267,I875275,I875292,I875309,I875326,I875343,I875388,I999577,I875419,I875436,I999565,I999574,I875462,I875470,I875501,I875518,I875535,I875552,I875624,I875650,I875658,I875698,I875706,I875723,I875740,I875780,I875802,I875819,I875845,I875853,I875870,I875887,I875904,I875921,I875966,I875997,I876014,I876040,I876048,I876079,I876096,I876113,I876130,I876202,I876228,I876236,I876276,I876284,I876301,I876318,I876358,I876380,I876397,I876423,I876431,I876448,I876465,I876482,I876499,I876544,I876575,I876592,I876618,I876626,I876657,I876674,I876691,I876708,I876780,I876806,I876814,I876854,I876862,I876879,I876896,I876936,I876958,I876975,I877001,I877009,I877026,I877043,I877060,I877077,I877122,I877153,I877170,I877196,I877204,I877235,I877252,I877269,I877286,I877358,I877384,I877392,I877432,I877440,I877457,I877474,I877514,I877536,I877553,I877579,I877587,I877604,I877621,I877638,I877655,I877700,I877731,I877748,I877774,I877782,I877813,I877830,I877847,I877864,I877936,I1016342,I877962,I877970,I1016324,I1016333,I878010,I878018,I1016318,I878035,I1016330,I878052,I878092,I878114,I1016321,I878131,I878157,I878165,I878182,I878199,I878216,I878233,I878278,I1016339,I878309,I878326,I1016327,I1016336,I878352,I878360,I878391,I878408,I878425,I878442,I878514,I878540,I878548,I878588,I878596,I878613,I878630,I878670,I878692,I878709,I878735,I878743,I878760,I878777,I878794,I878811,I878856,I878887,I878904,I878930,I878938,I878969,I878986,I879003,I879020,I879092,I879118,I879126,I879166,I879174,I879191,I879208,I879248,I879270,I879287,I879313,I879321,I879338,I879355,I879372,I879389,I879434,I879465,I879482,I879508,I879516,I879547,I879564,I879581,I879598,I879670,I879696,I879704,I879744,I879752,I879769,I879786,I879826,I879848,I879865,I879891,I879899,I879916,I879933,I879950,I879967,I880012,I880043,I880060,I880086,I880094,I880125,I880142,I880159,I880176,I880248,I880274,I880282,I880322,I880330,I880347,I880364,I880404,I880426,I880443,I880469,I880477,I880494,I880511,I880528,I880545,I880590,I880621,I880638,I880664,I880672,I880703,I880720,I880737,I880754,I880826,I880852,I880860,I880900,I880908,I880925,I880942,I880982,I881004,I881021,I881047,I881055,I881072,I881089,I881106,I881123,I881168,I881199,I881216,I881242,I881250,I881281,I881298,I881315,I881332,I881404,I881430,I881438,I881478,I881486,I881503,I881520,I881560,I881582,I881599,I881625,I881633,I881650,I881667,I881684,I881701,I881746,I881777,I881794,I881820,I881828,I881859,I881876,I881893,I881910,I881982,I882008,I882016,I882056,I882064,I882081,I882098,I882138,I882160,I882177,I882203,I882211,I882228,I882245,I882262,I882279,I882324,I882355,I882372,I882398,I882406,I882437,I882454,I882471,I882488,I882560,I882586,I882594,I882634,I882642,I882659,I882676,I882716,I882738,I882755,I882781,I882789,I882806,I882823,I882840,I882857,I882902,I882933,I882950,I882976,I882984,I883015,I883032,I883049,I883066,I883138,I883164,I883172,I883212,I883220,I883237,I883254,I883294,I883316,I883333,I883359,I883367,I883384,I883401,I883418,I883435,I883480,I883511,I883528,I883554,I883562,I883593,I883610,I883627,I883644,I883716,I883742,I883750,I883790,I883798,I883815,I883832,I883872,I883894,I883911,I883937,I883945,I883962,I883979,I883996,I884013,I884058,I884089,I884106,I884132,I884140,I884171,I884188,I884205,I884222,I884294,I884320,I884328,I884368,I884376,I884393,I884410,I884450,I884472,I884489,I884515,I884523,I884540,I884557,I884574,I884591,I884636,I884667,I884684,I884710,I884718,I884749,I884766,I884783,I884800,I884872,I884898,I884906,I884946,I884954,I884971,I884988,I885028,I885050,I885067,I885093,I885101,I885118,I885135,I885152,I885169,I885214,I885245,I885262,I885288,I885296,I885327,I885344,I885361,I885378,I885450,I885476,I885484,I885433,I885524,I885532,I885549,I885566,I885421,I885606,I885442,I885628,I885645,I885671,I885679,I885696,I885713,I885730,I885747,I885418,I885439,I885792,I885430,I885823,I885840,I885866,I885874,I885436,I885905,I885922,I885939,I885956,I885427,I885424,I886028,I886054,I886062,I886102,I886110,I886127,I886144,I886184,I886206,I886223,I886249,I886257,I886274,I886291,I886308,I886325,I886370,I886401,I886418,I886444,I886452,I886483,I886500,I886517,I886534,I886606,I886632,I886640,I886680,I886688,I886705,I886722,I886762,I886784,I886801,I886827,I886835,I886852,I886869,I886886,I886903,I886948,I886979,I886996,I887022,I887030,I887061,I887078,I887095,I887112,I887184,I887210,I887218,I887258,I887266,I887283,I887300,I887340,I887362,I887379,I887405,I887413,I887430,I887447,I887464,I887481,I887526,I887557,I887574,I887600,I887608,I887639,I887656,I887673,I887690,I887762,I887788,I887796,I887745,I887836,I887844,I887861,I887878,I887733,I887918,I887754,I887940,I887957,I887983,I887991,I888008,I888025,I888042,I888059,I887730,I887751,I888104,I887742,I888135,I888152,I888178,I888186,I887748,I888217,I888234,I888251,I888268,I887739,I887736,I888340,I888366,I888374,I888414,I888422,I888439,I888456,I888496,I888518,I888535,I888561,I888569,I888586,I888603,I888620,I888637,I888682,I888713,I888730,I888756,I888764,I888795,I888812,I888829,I888846,I888918,I1078106,I888944,I888952,I1078088,I1078079,I888992,I889000,I1078094,I889017,I1078082,I889034,I889074,I889096,I1078091,I889113,I889139,I889147,I889164,I1078100,I889181,I889198,I889215,I889260,I1078103,I889291,I889308,I1078097,I1078085,I889334,I889342,I889373,I889390,I889407,I889424,I889496,I889522,I889530,I889570,I889578,I889595,I889612,I889652,I889674,I889691,I889717,I889725,I889742,I889759,I889776,I889793,I889838,I889869,I889886,I889912,I889920,I889951,I889968,I889985,I890002,I890074,I890100,I890108,I890148,I890156,I890173,I890190,I890230,I890252,I890269,I890295,I890303,I890320,I890337,I890354,I890371,I890416,I890447,I890464,I890490,I890498,I890529,I890546,I890563,I890580,I890652,I1025991,I890678,I890686,I1026018,I890635,I1026000,I890726,I890734,I1026009,I890751,I1026012,I890768,I890623,I890808,I890644,I890830,I1026006,I890847,I890873,I890881,I890898,I1025994,I890915,I1025997,I890932,I890949,I890620,I890641,I890994,I1026015,I890632,I891025,I891042,I1026003,I891068,I891076,I890638,I891107,I891124,I891141,I891158,I890629,I890626,I891230,I891256,I891264,I891304,I891312,I891329,I891346,I891386,I891408,I891425,I891451,I891459,I891476,I891493,I891510,I891527,I891572,I891603,I891620,I891646,I891654,I891685,I891702,I891719,I891736,I891808,I891834,I891842,I891882,I891890,I891907,I891924,I891964,I891986,I892003,I892029,I892037,I892054,I892071,I892088,I892105,I892150,I892181,I892198,I892224,I892232,I892263,I892280,I892297,I892314,I892386,I1087031,I892412,I892420,I1087013,I1087004,I892460,I892468,I1087019,I892485,I1087007,I892502,I892542,I892564,I1087016,I892581,I892607,I892615,I892632,I1087025,I892649,I892666,I892683,I892728,I1087028,I892759,I892776,I1087022,I1087010,I892802,I892810,I892841,I892858,I892875,I892892,I892964,I892990,I892998,I893038,I893046,I893063,I893080,I893120,I893142,I893159,I893185,I893193,I893210,I893227,I893244,I893261,I893306,I893337,I893354,I893380,I893388,I893419,I893436,I893453,I893470,I893542,I893568,I893576,I893616,I893624,I893641,I893658,I893698,I893720,I893737,I893763,I893771,I893788,I893805,I893822,I893839,I893884,I893915,I893932,I893958,I893966,I893997,I894014,I894031,I894048,I894120,I894146,I894154,I894194,I894202,I894219,I894236,I894276,I894298,I894315,I894341,I894349,I894366,I894383,I894400,I894417,I894462,I894493,I894510,I894536,I894544,I894575,I894592,I894609,I894626,I894698,I894724,I894732,I894681,I894772,I894780,I894797,I894814,I894669,I894854,I894690,I894876,I894893,I894919,I894927,I894944,I894961,I894978,I894995,I894666,I894687,I895040,I894678,I895071,I895088,I895114,I895122,I894684,I895153,I895170,I895187,I895204,I894675,I894672,I895276,I895302,I895310,I895350,I895358,I895375,I895392,I895432,I895454,I895471,I895497,I895505,I895522,I895539,I895556,I895573,I895618,I895649,I895666,I895692,I895700,I895731,I895748,I895765,I895782,I895854,I895880,I895888,I895928,I895936,I895953,I895970,I896010,I896032,I896049,I896075,I896083,I896100,I896117,I896134,I896151,I896196,I896227,I896244,I896270,I896278,I896309,I896326,I896343,I896360,I896432,I1040621,I896458,I896466,I1040603,I1040594,I896506,I896514,I1040609,I896531,I1040597,I896548,I896588,I896610,I1040606,I896627,I896653,I896661,I896678,I1040615,I896695,I896712,I896729,I896774,I1040618,I896805,I896822,I1040612,I1040600,I896848,I896856,I896887,I896904,I896921,I896938,I897010,I1091196,I897036,I897044,I1091178,I1091169,I897084,I897092,I1091184,I897109,I1091172,I897126,I897166,I897188,I1091181,I897205,I897231,I897239,I897256,I1091190,I897273,I897290,I897307,I897352,I1091193,I897383,I897400,I1091187,I1091175,I897426,I897434,I897465,I897482,I897499,I897516,I897588,I897614,I897622,I897662,I897670,I897687,I897704,I897744,I897766,I897783,I897809,I897817,I897834,I897851,I897868,I897885,I897930,I897961,I897978,I898004,I898012,I898043,I898060,I898077,I898094,I898166,I959219,I898192,I898200,I959213,I959198,I898240,I898248,I959204,I898265,I959216,I898282,I898322,I898344,I898361,I898387,I898395,I898412,I959222,I898429,I959210,I898446,I898463,I898508,I959201,I898539,I898556,I959207,I898582,I898590,I898621,I898638,I898655,I898672,I898744,I898770,I898778,I898818,I898826,I898843,I898860,I898900,I898922,I898939,I898965,I898973,I898990,I899007,I899024,I899041,I899086,I899117,I899134,I899160,I899168,I899199,I899216,I899233,I899250,I899322,I899348,I899356,I899305,I899396,I899404,I899421,I899438,I899293,I899478,I899314,I899500,I899517,I899543,I899551,I899568,I899585,I899602,I899619,I899290,I899311,I899664,I899302,I899695,I899712,I899738,I899746,I899308,I899777,I899794,I899811,I899828,I899299,I899296,I899900,I899926,I899934,I899974,I899982,I899999,I900016,I900056,I900078,I900095,I900121,I900129,I900146,I900163,I900180,I900197,I900242,I900273,I900290,I900316,I900324,I900355,I900372,I900389,I900406,I900478,I900504,I900512,I900552,I900560,I900577,I900594,I900634,I900656,I900673,I900699,I900707,I900724,I900741,I900758,I900775,I900820,I900851,I900868,I900894,I900902,I900933,I900950,I900967,I900984,I901056,I901082,I901090,I901130,I901138,I901155,I901172,I901212,I901234,I901251,I901277,I901285,I901302,I901319,I901336,I901353,I901398,I901429,I901446,I901472,I901480,I901511,I901528,I901545,I901562,I901634,I901660,I901668,I901708,I901716,I901733,I901750,I901790,I901812,I901829,I901855,I901863,I901880,I901897,I901914,I901931,I901976,I902007,I902024,I902050,I902058,I902089,I902106,I902123,I902140,I902212,I902238,I902246,I902195,I902286,I902294,I902311,I902328,I902183,I902368,I902204,I902390,I902407,I902433,I902441,I902458,I902475,I902492,I902509,I902180,I902201,I902554,I902192,I902585,I902602,I902628,I902636,I902198,I902667,I902684,I902701,I902718,I902189,I902186,I902790,I902816,I902824,I902864,I902872,I902889,I902906,I902946,I902968,I902985,I903011,I903019,I903036,I903053,I903070,I903087,I903132,I903163,I903180,I903206,I903214,I903245,I903262,I903279,I903296,I903368,I903394,I903402,I903442,I903450,I903467,I903484,I903524,I903546,I903563,I903589,I903597,I903614,I903631,I903648,I903665,I903710,I903741,I903758,I903784,I903792,I903823,I903840,I903857,I903874,I903946,I967923,I903972,I903980,I967917,I967902,I904020,I904028,I967908,I904045,I967920,I904062,I904102,I904124,I904141,I904167,I904175,I904192,I967926,I904209,I967914,I904226,I904243,I904288,I967905,I904319,I904336,I967911,I904362,I904370,I904401,I904418,I904435,I904452,I904524,I904550,I904558,I904598,I904606,I904623,I904640,I904680,I904702,I904719,I904745,I904753,I904770,I904787,I904804,I904821,I904866,I904897,I904914,I904940,I904948,I904979,I904996,I905013,I905030,I905102,I905128,I905136,I905085,I905176,I905184,I905201,I905218,I905073,I905258,I905094,I905280,I905297,I905323,I905331,I905348,I905365,I905382,I905399,I905070,I905091,I905444,I905082,I905475,I905492,I905518,I905526,I905088,I905557,I905574,I905591,I905608,I905079,I905076,I905680,I905706,I905714,I905754,I905762,I905779,I905796,I905836,I905858,I905875,I905901,I905909,I905926,I905943,I905960,I905977,I906022,I906053,I906070,I906096,I906104,I906135,I906152,I906169,I906186,I906258,I906284,I906292,I906332,I906340,I906357,I906374,I906414,I906436,I906453,I906479,I906487,I906504,I906521,I906538,I906555,I906600,I906631,I906648,I906674,I906682,I906713,I906730,I906747,I906764,I906836,I906862,I906870,I906910,I906918,I906935,I906952,I906992,I907014,I907031,I907057,I907065,I907082,I907099,I907116,I907133,I907178,I907209,I907226,I907252,I907260,I907291,I907308,I907325,I907342,I907414,I907440,I907448,I907397,I907488,I907496,I907513,I907530,I907385,I907570,I907406,I907592,I907609,I907635,I907643,I907660,I907677,I907694,I907711,I907382,I907403,I907756,I907394,I907787,I907804,I907830,I907838,I907400,I907869,I907886,I907903,I907920,I907391,I907388,I907992,I908018,I908026,I908066,I908074,I908091,I908108,I908148,I908170,I908187,I908213,I908221,I908238,I908255,I908272,I908289,I908334,I908365,I908382,I908408,I908416,I908447,I908464,I908481,I908498,I908570,I908596,I908604,I908644,I908652,I908669,I908686,I908726,I908748,I908765,I908791,I908799,I908816,I908833,I908850,I908867,I908912,I908943,I908960,I908986,I908994,I909025,I909042,I909059,I909076,I909148,I909174,I909182,I909222,I909230,I909247,I909264,I909304,I909326,I909343,I909369,I909377,I909394,I909411,I909428,I909445,I909490,I909521,I909538,I909564,I909572,I909603,I909620,I909637,I909654,I909726,I909752,I909760,I909800,I909808,I909825,I909842,I909882,I909904,I909921,I909947,I909955,I909972,I909989,I910006,I910023,I910068,I910099,I910116,I910142,I910150,I910181,I910198,I910215,I910232,I910304,I969011,I910330,I910338,I969005,I968990,I910378,I910386,I968996,I910403,I969008,I910420,I910460,I910482,I910499,I910525,I910533,I910550,I969014,I910567,I969002,I910584,I910601,I910646,I968993,I910677,I910694,I968999,I910720,I910728,I910759,I910776,I910793,I910810,I910882,I910908,I910916,I910956,I910964,I910981,I910998,I911038,I911060,I911077,I911103,I911111,I911128,I911145,I911162,I911179,I911224,I911255,I911272,I911298,I911306,I911337,I911354,I911371,I911388,I911460,I911486,I911494,I911443,I911534,I911542,I911559,I911576,I911431,I911616,I911452,I911638,I911655,I911681,I911689,I911706,I911723,I911740,I911757,I911428,I911449,I911802,I911440,I911833,I911850,I911876,I911884,I911446,I911915,I911932,I911949,I911966,I911437,I911434,I912038,I912064,I912072,I912112,I912120,I912137,I912154,I912194,I912216,I912233,I912259,I912267,I912284,I912301,I912318,I912335,I912380,I912411,I912428,I912454,I912462,I912493,I912510,I912527,I912544,I912616,I912642,I912650,I912690,I912698,I912715,I912732,I912772,I912794,I912811,I912837,I912845,I912862,I912879,I912896,I912913,I912958,I912989,I913006,I913032,I913040,I913071,I913088,I913105,I913122,I913194,I993800,I913220,I913228,I993782,I993791,I913268,I913276,I993776,I913293,I993788,I913310,I913350,I913372,I993779,I913389,I913415,I913423,I913440,I913457,I913474,I913491,I913536,I993797,I913567,I913584,I993785,I993794,I913610,I913618,I913649,I913666,I913683,I913700,I913772,I913798,I913806,I913846,I913854,I913871,I913888,I913928,I913950,I913967,I913993,I914001,I914018,I914035,I914052,I914069,I914114,I914145,I914162,I914188,I914196,I914227,I914244,I914261,I914278,I914350,I914376,I914384,I914424,I914432,I914449,I914466,I914506,I914528,I914545,I914571,I914579,I914596,I914613,I914630,I914647,I914692,I914723,I914740,I914766,I914774,I914805,I914822,I914839,I914856,I914928,I914954,I914962,I915002,I915010,I915027,I915044,I915084,I915106,I915123,I915149,I915157,I915174,I915191,I915208,I915225,I915270,I915301,I915318,I915344,I915352,I915383,I915400,I915417,I915434,I915506,I915532,I915540,I915580,I915588,I915605,I915622,I915662,I915684,I915701,I915727,I915735,I915752,I915769,I915786,I915803,I915848,I915879,I915896,I915922,I915930,I915961,I915978,I915995,I916012,I916084,I916110,I916118,I916067,I916158,I916166,I916183,I916200,I916055,I916240,I916076,I916262,I916279,I916305,I916313,I916330,I916347,I916364,I916381,I916052,I916073,I916426,I916064,I916457,I916474,I916500,I916508,I916070,I916539,I916556,I916573,I916590,I916061,I916058,I916662,I916688,I916696,I916736,I916744,I916761,I916778,I916818,I916840,I916857,I916883,I916891,I916908,I916925,I916942,I916959,I917004,I917035,I917052,I917078,I917086,I917117,I917134,I917151,I917168,I917240,I917266,I917274,I917314,I917322,I917339,I917356,I917396,I917418,I917435,I917461,I917469,I917486,I917503,I917520,I917537,I917582,I917613,I917630,I917656,I917664,I917695,I917712,I917729,I917746,I917818,I977171,I917844,I917852,I977165,I977150,I917892,I917900,I977156,I917917,I977168,I917934,I917974,I917996,I918013,I918039,I918047,I918064,I977174,I918081,I977162,I918098,I918115,I918160,I977153,I918191,I918208,I977159,I918234,I918242,I918273,I918290,I918307,I918324,I918396,I918422,I918430,I918470,I918478,I918495,I918512,I918552,I918574,I918591,I918617,I918625,I918642,I918659,I918676,I918693,I918738,I918769,I918786,I918812,I918820,I918851,I918868,I918885,I918902,I918974,I919000,I919008,I919048,I919056,I919073,I919090,I919130,I919152,I919169,I919195,I919203,I919220,I919237,I919254,I919271,I919316,I919347,I919364,I919390,I919398,I919429,I919446,I919463,I919480,I919552,I919578,I919586,I919626,I919634,I919651,I919668,I919708,I919730,I919747,I919773,I919781,I919798,I919815,I919832,I919849,I919894,I919925,I919942,I919968,I919976,I920007,I920024,I920041,I920058,I920130,I1009984,I920156,I920164,I1009966,I1009975,I920204,I920212,I1009960,I920229,I1009972,I920246,I920286,I920308,I1009963,I920325,I920351,I920359,I920376,I920393,I920410,I920427,I920472,I1009981,I920503,I920520,I1009969,I1009978,I920546,I920554,I920585,I920602,I920619,I920636,I920708,I920734,I920742,I920691,I920782,I920790,I920807,I920824,I920679,I920864,I920700,I920886,I920903,I920929,I920937,I920954,I920971,I920988,I921005,I920676,I920697,I921050,I920688,I921081,I921098,I921124,I921132,I920694,I921163,I921180,I921197,I921214,I920685,I920682,I921286,I921312,I921320,I921269,I921360,I921368,I921385,I921402,I921257,I921442,I921278,I921464,I921481,I921507,I921515,I921532,I921549,I921566,I921583,I921254,I921275,I921628,I921266,I921659,I921676,I921702,I921710,I921272,I921741,I921758,I921775,I921792,I921263,I921260,I921864,I921890,I921898,I921938,I921946,I921963,I921980,I922020,I922042,I922059,I922085,I922093,I922110,I922127,I922144,I922161,I922206,I922237,I922254,I922280,I922288,I922319,I922336,I922353,I922370,I922442,I922468,I922476,I922516,I922524,I922541,I922558,I922598,I922620,I922637,I922663,I922671,I922688,I922705,I922722,I922739,I922784,I922815,I922832,I922858,I922866,I922897,I922914,I922931,I922948,I923020,I923046,I923054,I923003,I923094,I923102,I923119,I923136,I922991,I923176,I923012,I923198,I923215,I923241,I923249,I923266,I923283,I923300,I923317,I922988,I923009,I923362,I923000,I923393,I923410,I923436,I923444,I923006,I923475,I923492,I923509,I923526,I922997,I922994,I923598,I1100716,I923624,I923632,I1100698,I1100689,I923672,I923680,I1100704,I923697,I1100692,I923714,I923754,I923776,I1100701,I923793,I923819,I923827,I923844,I1100710,I923861,I923878,I923895,I923940,I1100713,I923971,I923988,I1100707,I1100695,I924014,I924022,I924053,I924070,I924087,I924104,I924176,I924202,I924210,I924250,I924258,I924275,I924292,I924332,I924354,I924371,I924397,I924405,I924422,I924439,I924456,I924473,I924518,I924549,I924566,I924592,I924600,I924631,I924648,I924665,I924682,I924754,I1008250,I924780,I924788,I1008232,I1008241,I924828,I924836,I1008226,I924853,I1008238,I924870,I924910,I924932,I1008229,I924949,I924975,I924983,I925000,I925017,I925034,I925051,I925096,I1008247,I925127,I925144,I1008235,I1008244,I925170,I925178,I925209,I925226,I925243,I925260,I925332,I925358,I925366,I925406,I925414,I925431,I925448,I925488,I925510,I925527,I925553,I925561,I925578,I925595,I925612,I925629,I925674,I925705,I925722,I925748,I925756,I925787,I925804,I925821,I925838,I925910,I925936,I925944,I925984,I925992,I926009,I926026,I926066,I926088,I926105,I926131,I926139,I926156,I926173,I926190,I926207,I926252,I926283,I926300,I926326,I926334,I926365,I926382,I926399,I926416,I926488,I926514,I926522,I926562,I926570,I926587,I926604,I926644,I926666,I926683,I926709,I926717,I926734,I926751,I926768,I926785,I926830,I926861,I926878,I926904,I926912,I926943,I926960,I926977,I926994,I927066,I927092,I927100,I927140,I927148,I927165,I927182,I927222,I927244,I927261,I927287,I927295,I927312,I927329,I927346,I927363,I927408,I927439,I927456,I927482,I927490,I927521,I927538,I927555,I927572,I927644,I927670,I927678,I927627,I927718,I927726,I927743,I927760,I927615,I927800,I927636,I927822,I927839,I927865,I927873,I927890,I927907,I927924,I927941,I927612,I927633,I927986,I927624,I928017,I928034,I928060,I928068,I927630,I928099,I928116,I928133,I928150,I927621,I927618,I928222,I928248,I928256,I928296,I928304,I928321,I928338,I928378,I928400,I928417,I928443,I928451,I928468,I928485,I928502,I928519,I928564,I928595,I928612,I928638,I928646,I928677,I928694,I928711,I928728,I928800,I928826,I928834,I928783,I928874,I928882,I928899,I928916,I928771,I928956,I928792,I928978,I928995,I929021,I929029,I929046,I929063,I929080,I929097,I928768,I928789,I929142,I928780,I929173,I929190,I929216,I929224,I928786,I929255,I929272,I929289,I929306,I928777,I928774,I929378,I929404,I929412,I929452,I929460,I929477,I929494,I929534,I929556,I929573,I929599,I929607,I929624,I929641,I929658,I929675,I929720,I929751,I929768,I929794,I929802,I929833,I929850,I929867,I929884,I929956,I929982,I929990,I930030,I930038,I930055,I930072,I930112,I930134,I930151,I930177,I930185,I930202,I930219,I930236,I930253,I930298,I930329,I930346,I930372,I930380,I930411,I930428,I930445,I930462,I930534,I930560,I930568,I930608,I930616,I930633,I930650,I930690,I930712,I930729,I930755,I930763,I930780,I930797,I930814,I930831,I930876,I930907,I930924,I930950,I930958,I930989,I931006,I931023,I931040,I931112,I1007672,I931138,I931146,I1007654,I1007663,I931186,I931194,I1007648,I931211,I1007660,I931228,I931268,I931290,I1007651,I931307,I931333,I931341,I931358,I931375,I931392,I931409,I931454,I1007669,I931485,I931502,I1007657,I1007666,I931528,I931536,I931567,I931584,I931601,I931618,I931690,I931716,I931724,I931764,I931772,I931789,I931806,I931846,I931868,I931885,I931911,I931919,I931936,I931953,I931970,I931987,I932032,I932063,I932080,I932106,I932114,I932145,I932162,I932179,I932196,I932268,I932294,I932302,I932342,I932350,I932367,I932384,I932424,I932446,I932463,I932489,I932497,I932514,I932531,I932548,I932565,I932610,I932641,I932658,I932684,I932692,I932723,I932740,I932757,I932774,I932846,I932872,I932880,I932920,I932928,I932945,I932962,I933002,I933024,I933041,I933067,I933075,I933092,I933109,I933126,I933143,I933188,I933219,I933236,I933262,I933270,I933301,I933318,I933335,I933352,I933424,I933450,I933458,I933498,I933506,I933523,I933540,I933580,I933602,I933619,I933645,I933653,I933670,I933687,I933704,I933721,I933766,I933797,I933814,I933840,I933848,I933879,I933896,I933913,I933930,I934002,I934028,I934036,I934076,I934084,I934101,I934118,I934158,I934180,I934197,I934223,I934231,I934248,I934265,I934282,I934299,I934344,I934375,I934392,I934418,I934426,I934457,I934474,I934491,I934508,I934580,I1044786,I934606,I934614,I1044768,I1044759,I934654,I934662,I1044774,I934679,I1044762,I934696,I934736,I934758,I1044771,I934775,I934801,I934809,I934826,I1044780,I934843,I934860,I934877,I934922,I1044783,I934953,I934970,I1044777,I1044765,I934996,I935004,I935035,I935052,I935069,I935086,I935158,I977715,I935184,I935192,I977709,I935141,I977694,I935232,I935240,I977700,I935257,I977712,I935274,I935129,I935314,I935150,I935336,I935353,I935379,I935387,I935404,I977718,I935421,I977706,I935438,I935455,I935126,I935147,I935500,I977697,I935138,I935531,I935548,I977703,I935574,I935582,I935144,I935613,I935630,I935647,I935664,I935135,I935132,I935736,I955955,I935762,I935770,I955949,I955934,I935810,I935818,I955940,I935835,I955952,I935852,I935892,I935914,I935931,I935957,I935965,I935982,I955958,I935999,I955946,I936016,I936033,I936078,I955937,I936109,I936126,I955943,I936152,I936160,I936191,I936208,I936225,I936242,I936314,I936340,I936348,I936388,I936396,I936413,I936430,I936470,I936492,I936509,I936535,I936543,I936560,I936577,I936594,I936611,I936656,I936687,I936704,I936730,I936738,I936769,I936786,I936803,I936820,I936892,I936918,I936926,I936875,I936966,I936974,I936991,I937008,I936863,I937048,I936884,I937070,I937087,I937113,I937121,I937138,I937155,I937172,I937189,I936860,I936881,I937234,I936872,I937265,I937282,I937308,I937316,I936878,I937347,I937364,I937381,I937398,I936869,I936866,I937470,I937496,I937504,I937544,I937552,I937569,I937586,I937626,I937648,I937665,I937691,I937699,I937716,I937733,I937750,I937767,I937812,I937843,I937860,I937886,I937894,I937925,I937942,I937959,I937976,I938048,I995534,I938074,I938082,I995516,I995525,I938122,I938130,I995510,I938147,I995522,I938164,I938204,I938226,I995513,I938243,I938269,I938277,I938294,I938311,I938328,I938345,I938390,I995531,I938421,I938438,I995519,I995528,I938464,I938472,I938503,I938520,I938537,I938554,I938626,I938652,I938660,I938700,I938708,I938725,I938742,I938782,I938804,I938821,I938847,I938855,I938872,I938889,I938906,I938923,I938968,I938999,I939016,I939042,I939050,I939081,I939098,I939115,I939132,I939204,I939230,I939238,I939278,I939286,I939303,I939320,I939360,I939382,I939399,I939425,I939433,I939450,I939467,I939484,I939501,I939546,I939577,I939594,I939620,I939628,I939659,I939676,I939693,I939710,I939782,I939808,I939816,I939856,I939864,I939881,I939898,I939938,I939960,I939977,I940003,I940011,I940028,I940045,I940062,I940079,I940124,I940155,I940172,I940198,I940206,I940237,I940254,I940271,I940288,I940360,I940386,I940394,I940434,I940442,I940459,I940476,I940516,I940538,I940555,I940581,I940589,I940606,I940623,I940640,I940657,I940702,I940733,I940750,I940776,I940784,I940815,I940832,I940849,I940866,I940938,I940964,I940972,I940921,I941012,I941020,I941037,I941054,I940909,I941094,I940930,I941116,I941133,I941159,I941167,I941184,I941201,I941218,I941235,I940906,I940927,I941280,I940918,I941311,I941328,I941354,I941362,I940924,I941393,I941410,I941427,I941444,I940915,I940912,I941516,I941542,I941550,I941590,I941598,I941615,I941632,I941672,I941694,I941711,I941737,I941745,I941762,I941779,I941796,I941813,I941858,I941889,I941906,I941932,I941940,I941971,I941988,I942005,I942022,I942094,I1060256,I942120,I942128,I1060238,I942077,I1060229,I942168,I942176,I1060244,I942193,I1060232,I942210,I942065,I942250,I942086,I942272,I1060241,I942289,I942315,I942323,I942340,I1060250,I942357,I942374,I942391,I942062,I942083,I942436,I1060253,I942074,I942467,I942484,I1060247,I1060235,I942510,I942518,I942080,I942549,I942566,I942583,I942600,I942071,I942068,I942672,I942698,I942706,I942746,I942754,I942771,I942788,I942828,I942850,I942867,I942893,I942901,I942918,I942935,I942952,I942969,I943014,I943045,I943062,I943088,I943096,I943127,I943144,I943161,I943178,I943250,I1069181,I943276,I943284,I1069163,I1069154,I943324,I943332,I1069169,I943349,I1069157,I943366,I943406,I943428,I1069166,I943445,I943471,I943479,I943496,I1069175,I943513,I943530,I943547,I943592,I1069178,I943623,I943640,I1069172,I1069160,I943666,I943674,I943705,I943722,I943739,I943756,I943828,I943854,I943862,I943902,I943910,I943927,I943944,I943984,I944006,I944023,I944049,I944057,I944074,I944091,I944108,I944125,I944170,I944201,I944218,I944244,I944252,I944283,I944300,I944317,I944334,I944406,I944432,I944440,I944389,I944480,I944488,I944505,I944522,I944377,I944562,I944398,I944584,I944601,I944627,I944635,I944652,I944669,I944686,I944703,I944374,I944395,I944748,I944386,I944779,I944796,I944822,I944830,I944392,I944861,I944878,I944895,I944912,I944383,I944380,I944984,I945010,I945018,I945058,I945066,I945083,I945100,I945140,I945162,I945179,I945205,I945213,I945230,I945247,I945264,I945281,I945326,I945357,I945374,I945400,I945408,I945439,I945456,I945473,I945490,I945562,I945588,I945596,I945636,I945644,I945661,I945678,I945718,I945740,I945757,I945783,I945791,I945808,I945825,I945842,I945859,I945904,I945935,I945952,I945978,I945986,I946017,I946034,I946051,I946068,I946140,I946166,I946174,I946214,I946222,I946239,I946256,I946296,I946318,I946335,I946361,I946369,I946386,I946403,I946420,I946437,I946482,I946513,I946530,I946556,I946564,I946595,I946612,I946629,I946646,I946718,I946744,I946752,I946792,I946800,I946817,I946834,I946874,I946896,I946913,I946939,I946947,I946964,I946981,I946998,I947015,I947060,I947091,I947108,I947134,I947142,I947173,I947190,I947207,I947224,I947296,I947322,I947330,I947279,I947370,I947378,I947395,I947412,I947267,I947452,I947288,I947474,I947491,I947517,I947525,I947542,I947559,I947576,I947593,I947264,I947285,I947638,I947276,I947669,I947686,I947712,I947720,I947282,I947751,I947768,I947785,I947802,I947273,I947270,I947874,I947900,I947908,I947948,I947956,I947973,I947990,I948030,I948052,I948069,I948095,I948103,I948120,I948137,I948154,I948171,I948216,I948247,I948264,I948290,I948298,I948329,I948346,I948363,I948380,I948452,I948478,I948486,I948526,I948534,I948551,I948568,I948608,I948630,I948647,I948673,I948681,I948698,I948715,I948732,I948749,I948794,I948825,I948842,I948868,I948876,I948907,I948924,I948941,I948958,I949030,I949056,I949064,I949013,I949104,I949112,I949129,I949146,I949001,I949186,I949022,I949208,I949225,I949251,I949259,I949276,I949293,I949310,I949327,I948998,I949019,I949372,I949010,I949403,I949420,I949446,I949454,I949016,I949485,I949502,I949519,I949536,I949007,I949004,I949608,I949634,I949642,I949682,I949690,I949707,I949724,I949764,I949786,I949803,I949829,I949837,I949854,I949871,I949888,I949905,I949950,I949981,I949998,I950024,I950032,I950063,I950080,I950097,I950114,I950186,I950212,I950220,I950260,I950268,I950285,I950302,I950342,I950364,I950381,I950407,I950415,I950432,I950449,I950466,I950483,I950528,I950559,I950576,I950602,I950610,I950641,I950658,I950675,I950692,I950764,I950790,I950798,I950747,I950838,I950846,I950863,I950880,I950735,I950920,I950756,I950942,I950959,I950985,I950993,I951010,I951027,I951044,I951061,I950732,I950753,I951106,I950744,I951137,I951154,I951180,I951188,I950750,I951219,I951236,I951253,I951270,I950741,I950738,I951342,I951368,I951376,I951416,I951424,I951441,I951458,I951498,I951520,I951537,I951563,I951571,I951588,I951605,I951622,I951639,I951684,I951715,I951732,I951758,I951766,I951797,I951814,I951831,I951848,I951920,I951946,I951954,I951994,I952002,I952019,I952036,I952076,I952098,I952115,I952141,I952149,I952166,I952183,I952200,I952217,I952262,I952293,I952310,I952336,I952344,I952375,I952392,I952409,I952426,I952498,I952524,I952532,I952572,I952580,I952597,I952614,I952654,I952676,I952693,I952719,I952727,I952744,I952761,I952778,I952795,I952840,I952871,I952888,I952914,I952922,I952953,I952970,I952987,I953004,I953076,I953102,I953110,I953150,I953158,I953175,I953192,I953232,I953254,I953271,I953297,I953305,I953322,I953339,I953356,I953373,I953418,I953449,I953466,I953492,I953500,I953531,I953548,I953565,I953582,I953654,I953680,I953688,I953728,I953736,I953753,I953770,I953810,I953832,I953849,I953875,I953883,I953900,I953917,I953934,I953951,I953996,I954027,I954044,I954070,I954078,I954109,I954126,I954143,I954160,I954232,I954258,I954266,I954306,I954314,I954331,I954348,I954388,I954410,I954427,I954453,I954461,I954478,I954495,I954512,I954529,I954574,I954605,I954622,I954648,I954656,I954687,I954704,I954721,I954738,I954810,I954836,I954844,I954884,I954892,I954909,I954926,I954966,I954988,I955005,I955031,I955039,I955056,I955073,I955090,I955107,I955152,I955183,I955200,I955226,I955234,I955265,I955282,I955299,I955316,I955388,I955414,I955422,I955462,I955470,I955487,I955504,I955544,I955566,I955583,I955609,I955617,I955634,I955651,I955668,I955685,I955730,I955761,I955778,I955804,I955812,I955843,I955860,I955877,I955894,I955966,I955992,I956000,I956026,I956043,I956065,I956082,I956099,I956116,I956133,I956164,I956181,I956198,I956215,I956260,I956277,I956294,I956353,I956379,I956387,I956404,I956421,I956452,I956510,I956536,I956544,I956570,I956587,I956609,I956626,I956643,I956660,I956677,I956708,I956725,I956742,I956759,I956804,I956821,I956838,I956897,I956923,I956931,I956948,I956965,I956996,I957054,I1092981,I957080,I957088,I1092966,I1092960,I957114,I957131,I957153,I1092954,I957170,I1092975,I957187,I1092963,I957204,I957221,I957252,I1092972,I957269,I1092978,I957286,I1092969,I957303,I957348,I1092957,I957365,I957382,I957441,I957467,I957475,I957492,I957509,I957540,I957598,I1024335,I957624,I957632,I1024320,I1024332,I957658,I957675,I957697,I1024326,I957714,I1024317,I957731,I1024311,I957748,I957765,I957796,I1024323,I957813,I1024308,I957830,I1024329,I957847,I957892,I1024314,I957909,I957926,I957985,I958011,I958019,I958036,I958053,I958084,I958142,I958168,I958176,I958202,I958219,I958241,I958258,I958275,I958292,I958309,I958340,I958357,I958374,I958391,I958436,I958453,I958470,I958529,I958555,I958563,I958580,I958597,I958628,I958686,I958712,I958720,I958746,I958763,I958785,I958802,I958819,I958836,I958853,I958884,I958901,I958918,I958935,I958980,I958997,I959014,I959073,I959099,I959107,I959124,I959141,I959172,I959230,I959256,I959264,I959290,I959307,I959329,I959346,I959363,I959380,I959397,I959428,I959445,I959462,I959479,I959524,I959541,I959558,I959617,I959643,I959651,I959668,I959685,I959716,I959774,I959800,I959808,I959834,I959851,I959873,I959890,I959907,I959924,I959941,I959972,I959989,I960006,I960023,I960068,I960085,I960102,I960161,I960187,I960195,I960212,I960229,I960260,I960318,I960344,I960352,I960378,I960395,I960417,I960434,I960451,I960468,I960485,I960516,I960533,I960550,I960567,I960612,I960629,I960646,I960705,I960731,I960739,I960756,I960773,I960804,I960862,I1059661,I960888,I960896,I1059646,I1059640,I960922,I960939,I960961,I1059634,I960978,I1059655,I960995,I1059643,I961012,I961029,I961060,I1059652,I961077,I1059658,I961094,I1059649,I961111,I961156,I1059637,I961173,I961190,I961249,I961275,I961283,I961300,I961317,I961348,I961406,I961432,I961440,I961466,I961483,I961505,I961522,I961539,I961556,I961573,I961604,I961621,I961638,I961655,I961700,I961717,I961734,I961793,I961819,I961827,I961844,I961861,I961892,I961950,I961976,I961984,I962010,I962027,I962049,I962066,I962083,I962100,I962117,I962148,I962165,I962182,I962199,I962244,I962261,I962278,I962337,I962363,I962371,I962388,I962405,I962436,I962494,I962520,I962528,I962554,I962571,I962593,I962610,I962627,I962644,I962661,I962692,I962709,I962726,I962743,I962788,I962805,I962822,I962881,I962907,I962915,I962932,I962949,I962980,I963038,I1053116,I963064,I963072,I1053101,I1053095,I963098,I963115,I963137,I1053089,I963154,I1053110,I963171,I1053098,I963188,I963205,I963236,I1053107,I963253,I1053113,I963270,I1053104,I963287,I963332,I1053092,I963349,I963366,I963425,I963451,I963459,I963476,I963493,I963524,I963582,I963608,I963616,I963642,I963659,I963681,I963698,I963715,I963732,I963749,I963780,I963797,I963814,I963831,I963876,I963893,I963910,I963969,I963995,I964003,I964020,I964037,I964068,I964126,I964152,I964160,I964186,I964203,I964225,I964242,I964259,I964276,I964293,I964324,I964341,I964358,I964375,I964420,I964437,I964454,I964513,I964539,I964547,I964564,I964581,I964612,I964670,I964696,I964704,I964730,I964747,I964769,I964786,I964803,I964820,I964837,I964868,I964885,I964902,I964919,I964964,I964981,I964998,I965057,I965083,I965091,I965108,I965125,I965156,I965214,I965240,I965248,I965274,I965291,I965313,I965330,I965347,I965364,I965381,I965412,I965429,I965446,I965463,I965508,I965525,I965542,I965601,I965627,I965635,I965652,I965669,I965700,I965758,I965784,I965792,I965818,I965835,I965857,I965874,I965891,I965908,I965925,I965956,I965973,I965990,I966007,I966052,I966069,I966086,I966145,I966171,I966179,I966196,I966213,I966244,I966302,I966328,I966336,I966362,I966379,I966294,I966401,I966418,I966435,I966452,I966469,I966273,I966500,I966517,I966534,I966551,I966276,I966291,I966596,I966613,I966630,I966288,I966285,I966282,I966689,I966715,I966723,I966740,I966757,I966270,I966788,I966279,I966846,I966872,I966880,I966906,I966923,I966945,I966962,I966979,I966996,I967013,I967044,I967061,I967078,I967095,I967140,I967157,I967174,I967233,I967259,I967267,I967284,I967301,I967332,I967390,I967416,I967424,I967450,I967467,I967489,I967506,I967523,I967540,I967557,I967588,I967605,I967622,I967639,I967684,I967701,I967718,I967777,I967803,I967811,I967828,I967845,I967876,I967934,I967960,I967968,I967994,I968011,I968033,I968050,I968067,I968084,I968101,I968132,I968149,I968166,I968183,I968228,I968245,I968262,I968321,I968347,I968355,I968372,I968389,I968420,I968478,I968504,I968512,I968538,I968555,I968577,I968594,I968611,I968628,I968645,I968676,I968693,I968710,I968727,I968772,I968789,I968806,I968865,I968891,I968899,I968916,I968933,I968964,I969022,I969048,I969056,I969082,I969099,I969121,I969138,I969155,I969172,I969189,I969220,I969237,I969254,I969271,I969316,I969333,I969350,I969409,I969435,I969443,I969460,I969477,I969508,I969566,I969592,I969600,I969626,I969643,I969665,I969682,I969699,I969716,I969733,I969764,I969781,I969798,I969815,I969860,I969877,I969894,I969953,I969979,I969987,I970004,I970021,I970052,I970110,I970136,I970144,I970170,I970187,I970209,I970226,I970243,I970260,I970277,I970308,I970325,I970342,I970359,I970404,I970421,I970438,I970497,I970523,I970531,I970548,I970565,I970596,I970654,I970680,I970688,I970714,I970731,I970753,I970770,I970787,I970804,I970821,I970852,I970869,I970886,I970903,I970948,I970965,I970982,I971041,I971067,I971075,I971092,I971109,I971140,I971198,I971224,I971232,I971258,I971275,I971297,I971314,I971331,I971348,I971365,I971396,I971413,I971430,I971447,I971492,I971509,I971526,I971585,I971611,I971619,I971636,I971653,I971684,I971742,I971768,I971776,I971802,I971819,I971841,I971858,I971875,I971892,I971909,I971940,I971957,I971974,I971991,I972036,I972053,I972070,I972129,I972155,I972163,I972180,I972197,I972228,I972286,I972312,I972320,I972346,I972363,I972385,I972402,I972419,I972436,I972453,I972484,I972501,I972518,I972535,I972580,I972597,I972614,I972673,I972699,I972707,I972724,I972741,I972772,I972830,I972856,I972864,I972890,I972907,I972929,I972946,I972963,I972980,I972997,I973028,I973045,I973062,I973079,I973124,I973141,I973158,I973217,I973243,I973251,I973268,I973285,I973316,I973374,I973400,I973408,I973434,I973451,I973473,I973490,I973507,I973524,I973541,I973572,I973589,I973606,I973623,I973668,I973685,I973702,I973761,I973787,I973795,I973812,I973829,I973860,I973918,I973944,I973952,I973978,I973995,I974017,I974034,I974051,I974068,I974085,I974116,I974133,I974150,I974167,I974212,I974229,I974246,I974305,I974331,I974339,I974356,I974373,I974404,I974462,I974488,I974496,I974522,I974539,I974561,I974578,I974595,I974612,I974629,I974660,I974677,I974694,I974711,I974756,I974773,I974790,I974849,I974875,I974883,I974900,I974917,I974948,I975006,I975032,I975040,I975066,I975083,I975105,I975122,I975139,I975156,I975173,I975204,I975221,I975238,I975255,I975300,I975317,I975334,I975393,I975419,I975427,I975444,I975461,I975492,I975550,I975576,I975584,I975610,I975627,I975649,I975666,I975683,I975700,I975717,I975748,I975765,I975782,I975799,I975844,I975861,I975878,I975937,I975963,I975971,I975988,I976005,I976036,I976094,I976120,I976128,I976154,I976171,I976193,I976210,I976227,I976244,I976261,I976292,I976309,I976326,I976343,I976388,I976405,I976422,I976481,I976507,I976515,I976532,I976549,I976580,I976638,I976664,I976672,I976698,I976715,I976737,I976754,I976771,I976788,I976805,I976836,I976853,I976870,I976887,I976932,I976949,I976966,I977025,I977051,I977059,I977076,I977093,I977124,I977182,I977208,I977216,I977242,I977259,I977281,I977298,I977315,I977332,I977349,I977380,I977397,I977414,I977431,I977476,I977493,I977510,I977569,I977595,I977603,I977620,I977637,I977668,I977726,I1064421,I977752,I977760,I1064406,I1064400,I977786,I977803,I977825,I1064394,I977842,I1064415,I977859,I1064403,I977876,I977893,I977924,I1064412,I977941,I1064418,I977958,I1064409,I977975,I978020,I1064397,I978037,I978054,I978113,I978139,I978147,I978164,I978181,I978212,I978270,I978296,I978304,I978330,I978347,I978369,I978386,I978403,I978420,I978437,I978468,I978485,I978502,I978519,I978564,I978581,I978598,I978657,I978683,I978691,I978708,I978725,I978756,I978814,I978840,I978848,I978874,I978891,I978913,I978930,I978947,I978964,I978981,I979012,I979029,I979046,I979063,I979108,I979125,I979142,I979201,I979227,I979235,I979252,I979269,I979300,I979358,I979384,I979392,I979418,I979435,I979457,I979474,I979491,I979508,I979525,I979556,I979573,I979590,I979607,I979652,I979669,I979686,I979745,I979771,I979779,I979796,I979813,I979844,I979902,I979928,I979936,I979962,I979979,I980001,I980018,I980035,I980052,I980069,I980100,I980117,I980134,I980151,I980196,I980213,I980230,I980289,I980315,I980323,I980340,I980357,I980388,I980446,I980472,I980480,I980506,I980523,I980545,I980562,I980579,I980596,I980613,I980644,I980661,I980678,I980695,I980740,I980757,I980774,I980833,I980859,I980867,I980884,I980901,I980932,I980990,I981016,I981024,I981050,I981067,I980982,I981089,I981106,I981123,I981140,I981157,I980961,I981188,I981205,I981222,I981239,I980964,I980979,I981284,I981301,I981318,I980976,I980973,I980970,I981377,I981403,I981411,I981428,I981445,I980958,I981476,I980967,I981534,I981560,I981568,I981594,I981611,I981633,I981650,I981667,I981684,I981701,I981732,I981749,I981766,I981783,I981828,I981845,I981862,I981921,I981947,I981955,I981972,I981989,I982020,I982078,I1050736,I982104,I982112,I1050721,I1050715,I982138,I982155,I982177,I1050709,I982194,I1050730,I982211,I1050718,I982228,I982245,I982276,I1050727,I982293,I1050733,I982310,I1050724,I982327,I982372,I1050712,I982389,I982406,I982465,I982491,I982499,I982516,I982533,I982564,I982622,I982648,I982656,I982682,I982699,I982721,I982738,I982755,I982772,I982789,I982820,I982837,I982854,I982871,I982916,I982933,I982950,I983009,I983035,I983043,I983060,I983077,I983108,I983166,I983192,I983200,I983226,I983243,I983265,I983282,I983299,I983316,I983333,I983364,I983381,I983398,I983415,I983460,I983477,I983494,I983553,I983579,I983587,I983604,I983621,I983652,I983710,I983736,I983744,I983770,I983787,I983809,I983826,I983843,I983860,I983877,I983908,I983925,I983942,I983959,I984004,I984021,I984038,I984097,I984123,I984131,I984148,I984165,I984196,I984254,I984280,I984288,I984314,I984331,I984353,I984370,I984387,I984404,I984421,I984452,I984469,I984486,I984503,I984548,I984565,I984582,I984641,I984667,I984675,I984692,I984709,I984740,I984798,I984824,I984832,I984858,I984875,I984897,I984914,I984931,I984948,I984965,I984996,I985013,I985030,I985047,I985092,I985109,I985126,I985185,I985211,I985219,I985236,I985253,I985284,I985342,I1049546,I985368,I985376,I1049531,I1049525,I985402,I985419,I985441,I1049519,I985458,I1049540,I985475,I1049528,I985492,I985509,I985540,I1049537,I985557,I1049543,I985574,I1049534,I985591,I985636,I1049522,I985653,I985670,I985729,I985755,I985763,I985780,I985797,I985828,I985886,I985912,I985920,I985946,I985963,I985985,I986002,I986019,I986036,I986053,I986084,I986101,I986118,I986135,I986180,I986197,I986214,I986273,I986299,I986307,I986324,I986341,I986372,I986430,I986456,I986464,I986490,I986507,I986529,I986546,I986563,I986580,I986597,I986628,I986645,I986662,I986679,I986724,I986741,I986758,I986817,I986843,I986851,I986868,I986885,I986916,I986974,I987000,I987008,I987034,I987051,I987073,I987090,I987107,I987124,I987141,I987172,I987189,I987206,I987223,I987268,I987285,I987302,I987361,I987387,I987395,I987412,I987429,I987460,I987518,I987544,I987552,I987578,I987595,I987617,I987634,I987651,I987668,I987685,I987716,I987733,I987750,I987767,I987812,I987829,I987846,I987905,I987931,I987939,I987956,I987973,I988004,I988062,I988088,I988096,I988122,I988139,I988161,I988178,I988195,I988212,I988229,I988260,I988277,I988294,I988311,I988356,I988373,I988390,I988449,I988475,I988483,I988500,I988517,I988548,I988606,I1048948,I988632,I988640,I1048939,I988657,I1048924,I988683,I988691,I988708,I1048927,I988725,I1048936,I988742,I988759,I1048933,I988790,I1048945,I988807,I988824,I988855,I1048930,I988872,I988912,I988920,I988951,I1048951,I988968,I988985,I989002,I989033,I989064,I1048942,I989090,I989112,I989184,I989210,I989218,I989235,I989261,I989269,I989286,I989303,I989320,I989337,I989368,I989385,I989402,I989433,I989450,I989490,I989498,I989529,I989546,I989563,I989580,I989611,I989642,I989668,I989690,I989762,I989788,I989796,I989813,I989839,I989847,I989864,I989881,I989898,I989915,I989946,I989963,I989980,I990011,I990028,I990068,I990076,I990107,I990124,I990141,I990158,I990189,I990220,I990246,I990268,I990340,I990366,I990374,I990391,I990417,I990425,I990442,I990459,I990476,I990493,I990524,I990541,I990558,I990589,I990606,I990646,I990654,I990685,I990702,I990719,I990736,I990767,I990798,I990824,I990846,I990918,I990944,I990952,I990969,I990995,I991003,I991020,I991037,I991054,I991071,I991102,I991119,I991136,I991167,I991184,I991224,I991232,I991263,I991280,I991297,I991314,I991345,I991376,I991402,I991424,I991496,I991522,I991530,I991547,I991573,I991581,I991598,I991615,I991632,I991649,I991680,I991697,I991714,I991745,I991762,I991802,I991810,I991841,I991858,I991875,I991892,I991923,I991954,I991980,I992002,I992074,I992100,I992108,I992125,I992151,I992159,I992176,I992193,I992210,I992227,I992258,I992275,I992292,I992323,I992340,I992380,I992388,I992419,I992436,I992453,I992470,I992501,I992532,I992558,I992580,I992652,I992678,I992686,I992703,I992729,I992737,I992754,I992771,I992788,I992805,I992836,I992853,I992870,I992901,I992918,I992958,I992966,I992997,I993014,I993031,I993048,I993079,I993110,I993136,I993158,I993230,I993256,I993264,I993281,I993307,I993315,I993332,I993349,I993366,I993383,I993414,I993431,I993448,I993479,I993496,I993536,I993544,I993575,I993592,I993609,I993626,I993657,I993688,I993714,I993736,I993808,I993834,I993842,I993859,I993885,I993893,I993910,I993927,I993944,I993961,I993992,I994009,I994026,I994057,I994074,I994114,I994122,I994153,I994170,I994187,I994204,I994235,I994266,I994292,I994314,I994386,I1069773,I994412,I994420,I1069764,I994437,I1069749,I994463,I994471,I994488,I1069752,I994505,I1069761,I994522,I994539,I1069758,I994570,I1069770,I994587,I994604,I994635,I1069755,I994652,I994692,I994700,I994731,I1069776,I994748,I994765,I994782,I994813,I994844,I1069767,I994870,I994892,I994964,I994990,I994998,I995015,I995041,I995049,I995066,I995083,I995100,I995117,I995148,I995165,I995182,I995213,I995230,I995270,I995278,I995309,I995326,I995343,I995360,I995391,I995422,I995448,I995470,I995542,I995568,I995576,I995593,I995619,I995627,I995644,I995661,I995678,I995695,I995726,I995743,I995760,I995791,I995808,I995848,I995856,I995887,I995904,I995921,I995938,I995969,I996000,I996026,I996048,I996120,I996146,I996154,I996171,I996197,I996205,I996222,I996239,I996256,I996273,I996304,I996321,I996338,I996369,I996386,I996426,I996434,I996465,I996482,I996499,I996516,I996547,I996578,I996604,I996626,I996698,I996724,I996732,I996749,I996775,I996783,I996800,I996817,I996834,I996851,I996882,I996899,I996916,I996947,I996964,I997004,I997012,I997043,I997060,I997077,I997094,I997125,I997156,I997182,I997204,I997276,I997302,I997310,I997327,I997353,I997361,I997378,I997395,I997412,I997429,I997268,I997460,I997477,I997494,I997247,I997525,I997542,I997253,I997582,I997590,I997262,I997621,I997638,I997655,I997672,I997265,I997703,I997244,I997734,I997760,I997259,I997782,I997256,I997250,I997854,I997880,I997888,I997905,I997931,I997939,I997956,I997973,I997990,I998007,I998038,I998055,I998072,I998103,I998120,I998160,I998168,I998199,I998216,I998233,I998250,I998281,I998312,I998338,I998360,I998432,I998458,I998466,I998483,I998509,I998517,I998534,I998551,I998568,I998585,I998616,I998633,I998650,I998681,I998698,I998738,I998746,I998777,I998794,I998811,I998828,I998859,I998890,I998916,I998938,I999010,I999036,I999044,I999061,I999087,I999095,I999112,I999129,I999146,I999163,I999002,I999194,I999211,I999228,I998981,I999259,I999276,I998987,I999316,I999324,I998996,I999355,I999372,I999389,I999406,I998999,I999437,I998978,I999468,I999494,I998993,I999516,I998990,I998984,I999588,I999614,I999622,I999639,I999665,I999673,I999690,I999707,I999724,I999741,I999772,I999789,I999806,I999837,I999854,I999894,I999902,I999933,I999950,I999967,I999984,I1000015,I1000046,I1000072,I1000094,I1000166,I1000192,I1000200,I1000217,I1000243,I1000251,I1000268,I1000285,I1000302,I1000319,I1000350,I1000367,I1000384,I1000415,I1000432,I1000472,I1000480,I1000511,I1000528,I1000545,I1000562,I1000593,I1000624,I1000650,I1000672,I1000744,I1000770,I1000778,I1000795,I1000821,I1000829,I1000846,I1000863,I1000880,I1000897,I1000928,I1000945,I1000962,I1000993,I1001010,I1001050,I1001058,I1001089,I1001106,I1001123,I1001140,I1001171,I1001202,I1001228,I1001250,I1001322,I1001348,I1001356,I1001373,I1001399,I1001407,I1001424,I1001441,I1001458,I1001475,I1001314,I1001506,I1001523,I1001540,I1001293,I1001571,I1001588,I1001299,I1001628,I1001636,I1001308,I1001667,I1001684,I1001701,I1001718,I1001311,I1001749,I1001290,I1001780,I1001806,I1001305,I1001828,I1001302,I1001296,I1001900,I1001926,I1001934,I1001951,I1001977,I1001985,I1002002,I1002019,I1002036,I1002053,I1002084,I1002101,I1002118,I1002149,I1002166,I1002206,I1002214,I1002245,I1002262,I1002279,I1002296,I1002327,I1002358,I1002384,I1002406,I1002478,I1002504,I1002512,I1002529,I1002555,I1002563,I1002580,I1002597,I1002614,I1002631,I1002662,I1002679,I1002696,I1002727,I1002744,I1002784,I1002792,I1002823,I1002840,I1002857,I1002874,I1002905,I1002936,I1002962,I1002984,I1003056,I1003082,I1003090,I1003107,I1003133,I1003141,I1003158,I1003175,I1003192,I1003209,I1003240,I1003257,I1003274,I1003305,I1003322,I1003362,I1003370,I1003401,I1003418,I1003435,I1003452,I1003483,I1003514,I1003540,I1003562,I1003634,I1003660,I1003668,I1003685,I1003711,I1003719,I1003736,I1003753,I1003770,I1003787,I1003818,I1003835,I1003852,I1003883,I1003900,I1003940,I1003948,I1003979,I1003996,I1004013,I1004030,I1004061,I1004092,I1004118,I1004140,I1004212,I1004238,I1004246,I1004263,I1004289,I1004297,I1004314,I1004331,I1004348,I1004365,I1004204,I1004396,I1004413,I1004430,I1004183,I1004461,I1004478,I1004189,I1004518,I1004526,I1004198,I1004557,I1004574,I1004591,I1004608,I1004201,I1004639,I1004180,I1004670,I1004696,I1004195,I1004718,I1004192,I1004186,I1004790,I1004816,I1004824,I1004841,I1004867,I1004875,I1004892,I1004909,I1004926,I1004943,I1004974,I1004991,I1005008,I1005039,I1005056,I1005096,I1005104,I1005135,I1005152,I1005169,I1005186,I1005217,I1005248,I1005274,I1005296,I1005368,I1005394,I1005402,I1005419,I1005445,I1005453,I1005470,I1005487,I1005504,I1005521,I1005552,I1005569,I1005586,I1005617,I1005634,I1005674,I1005682,I1005713,I1005730,I1005747,I1005764,I1005795,I1005826,I1005852,I1005874,I1005946,I1005972,I1005980,I1005997,I1006023,I1006031,I1006048,I1006065,I1006082,I1006099,I1006130,I1006147,I1006164,I1006195,I1006212,I1006252,I1006260,I1006291,I1006308,I1006325,I1006342,I1006373,I1006404,I1006430,I1006452,I1006524,I1006550,I1006558,I1006575,I1006601,I1006609,I1006626,I1006643,I1006660,I1006677,I1006708,I1006725,I1006742,I1006773,I1006790,I1006830,I1006838,I1006869,I1006886,I1006903,I1006920,I1006951,I1006982,I1007008,I1007030,I1007102,I1007128,I1007136,I1007153,I1007179,I1007187,I1007204,I1007221,I1007238,I1007255,I1007286,I1007303,I1007320,I1007351,I1007368,I1007408,I1007416,I1007447,I1007464,I1007481,I1007498,I1007529,I1007560,I1007586,I1007608,I1007680,I1007706,I1007714,I1007731,I1007757,I1007765,I1007782,I1007799,I1007816,I1007833,I1007864,I1007881,I1007898,I1007929,I1007946,I1007986,I1007994,I1008025,I1008042,I1008059,I1008076,I1008107,I1008138,I1008164,I1008186,I1008258,I1008284,I1008292,I1008309,I1008335,I1008343,I1008360,I1008377,I1008394,I1008411,I1008442,I1008459,I1008476,I1008507,I1008524,I1008564,I1008572,I1008603,I1008620,I1008637,I1008654,I1008685,I1008716,I1008742,I1008764,I1008836,I1008862,I1008870,I1008887,I1008913,I1008921,I1008938,I1008955,I1008972,I1008989,I1009020,I1009037,I1009054,I1009085,I1009102,I1009142,I1009150,I1009181,I1009198,I1009215,I1009232,I1009263,I1009294,I1009320,I1009342,I1009414,I1009440,I1009448,I1009465,I1009491,I1009499,I1009516,I1009533,I1009550,I1009567,I1009598,I1009615,I1009632,I1009663,I1009680,I1009720,I1009728,I1009759,I1009776,I1009793,I1009810,I1009841,I1009872,I1009898,I1009920,I1009992,I1010018,I1010026,I1010043,I1010069,I1010077,I1010094,I1010111,I1010128,I1010145,I1010176,I1010193,I1010210,I1010241,I1010258,I1010298,I1010306,I1010337,I1010354,I1010371,I1010388,I1010419,I1010450,I1010476,I1010498,I1010570,I1010596,I1010604,I1010621,I1010647,I1010655,I1010672,I1010689,I1010706,I1010723,I1010754,I1010771,I1010788,I1010819,I1010836,I1010876,I1010884,I1010915,I1010932,I1010949,I1010966,I1010997,I1011028,I1011054,I1011076,I1011148,I1047758,I1011174,I1011182,I1047749,I1011199,I1047734,I1011225,I1011233,I1011250,I1047737,I1011267,I1047746,I1011284,I1011301,I1047743,I1011332,I1047755,I1011349,I1011366,I1011397,I1047740,I1011414,I1011454,I1011462,I1011493,I1047761,I1011510,I1011527,I1011544,I1011575,I1011606,I1047752,I1011632,I1011654,I1011726,I1011752,I1011760,I1011777,I1011803,I1011811,I1011828,I1011845,I1011862,I1011879,I1011910,I1011927,I1011944,I1011975,I1011992,I1012032,I1012040,I1012071,I1012088,I1012105,I1012122,I1012153,I1012184,I1012210,I1012232,I1012304,I1012330,I1012338,I1012355,I1012381,I1012389,I1012406,I1012423,I1012440,I1012457,I1012488,I1012505,I1012522,I1012553,I1012570,I1012610,I1012618,I1012649,I1012666,I1012683,I1012700,I1012731,I1012762,I1012788,I1012810,I1012882,I1012908,I1012916,I1012933,I1012959,I1012967,I1012984,I1013001,I1013018,I1013035,I1013066,I1013083,I1013100,I1013131,I1013148,I1013188,I1013196,I1013227,I1013244,I1013261,I1013278,I1013309,I1013340,I1013366,I1013388,I1013460,I1013486,I1013494,I1013511,I1013537,I1013545,I1013562,I1013579,I1013596,I1013613,I1013644,I1013661,I1013678,I1013709,I1013726,I1013766,I1013774,I1013805,I1013822,I1013839,I1013856,I1013887,I1013918,I1013944,I1013966,I1014038,I1014064,I1014072,I1014089,I1014115,I1014123,I1014140,I1014157,I1014174,I1014191,I1014222,I1014239,I1014256,I1014287,I1014304,I1014344,I1014352,I1014383,I1014400,I1014417,I1014434,I1014465,I1014496,I1014522,I1014544,I1014616,I1014642,I1014650,I1014667,I1014693,I1014701,I1014718,I1014735,I1014752,I1014769,I1014800,I1014817,I1014834,I1014865,I1014882,I1014922,I1014930,I1014961,I1014978,I1014995,I1015012,I1015043,I1015074,I1015100,I1015122,I1015194,I1015220,I1015228,I1015245,I1015271,I1015279,I1015296,I1015313,I1015330,I1015347,I1015378,I1015395,I1015412,I1015443,I1015460,I1015500,I1015508,I1015539,I1015556,I1015573,I1015590,I1015621,I1015652,I1015678,I1015700,I1015772,I1015798,I1015806,I1015823,I1015849,I1015857,I1015874,I1015891,I1015908,I1015925,I1015956,I1015973,I1015990,I1016021,I1016038,I1016078,I1016086,I1016117,I1016134,I1016151,I1016168,I1016199,I1016230,I1016256,I1016278,I1016350,I1016376,I1016384,I1016401,I1016427,I1016435,I1016452,I1016469,I1016486,I1016503,I1016534,I1016551,I1016568,I1016599,I1016616,I1016656,I1016664,I1016695,I1016712,I1016729,I1016746,I1016777,I1016808,I1016834,I1016856,I1016928,I1016954,I1016962,I1016979,I1017005,I1017013,I1017030,I1017047,I1017064,I1017081,I1016920,I1017112,I1017129,I1017146,I1016899,I1017177,I1017194,I1016905,I1017234,I1017242,I1016914,I1017273,I1017290,I1017307,I1017324,I1016917,I1017355,I1016896,I1017386,I1017412,I1016911,I1017434,I1016908,I1016902,I1017506,I1017532,I1017540,I1017557,I1017583,I1017591,I1017608,I1017625,I1017642,I1017659,I1017690,I1017707,I1017724,I1017755,I1017772,I1017812,I1017820,I1017851,I1017868,I1017885,I1017902,I1017933,I1017964,I1017990,I1018012,I1018084,I1018110,I1018118,I1018135,I1018161,I1018169,I1018186,I1018203,I1018220,I1018237,I1018268,I1018285,I1018302,I1018333,I1018350,I1018390,I1018398,I1018429,I1018446,I1018463,I1018480,I1018511,I1018542,I1018568,I1018590,I1018662,I1090003,I1018688,I1018696,I1089994,I1018713,I1089979,I1018739,I1018747,I1018764,I1089982,I1018781,I1089991,I1018798,I1018815,I1089988,I1018654,I1018846,I1090000,I1018863,I1018880,I1018633,I1018911,I1089985,I1018928,I1018639,I1018968,I1018976,I1018648,I1019007,I1090006,I1019024,I1019041,I1019058,I1018651,I1019089,I1018630,I1019120,I1089997,I1019146,I1018645,I1019168,I1018642,I1018636,I1019240,I1019266,I1019274,I1019291,I1019317,I1019325,I1019342,I1019359,I1019376,I1019393,I1019424,I1019441,I1019458,I1019489,I1019506,I1019546,I1019554,I1019585,I1019602,I1019619,I1019636,I1019667,I1019698,I1019724,I1019746,I1019818,I1019844,I1019852,I1019869,I1019895,I1019903,I1019920,I1019937,I1019954,I1019971,I1020002,I1020019,I1020036,I1020067,I1020084,I1020124,I1020132,I1020163,I1020180,I1020197,I1020214,I1020245,I1020276,I1020302,I1020324,I1020396,I1020422,I1020430,I1020447,I1020473,I1020481,I1020498,I1020515,I1020532,I1020549,I1020580,I1020597,I1020614,I1020645,I1020662,I1020702,I1020710,I1020741,I1020758,I1020775,I1020792,I1020823,I1020854,I1020880,I1020902,I1020977,I1021003,I1021011,I1021028,I1021054,I1021062,I1021079,I1021096,I1021127,I1021158,I1021175,I1021192,I1021209,I1021226,I1021257,I1021316,I1021333,I1021359,I1021381,I1021407,I1021415,I1021432,I1021463,I1021538,I1021564,I1021572,I1021589,I1021615,I1021623,I1021640,I1021657,I1021688,I1021719,I1021736,I1021753,I1021770,I1021787,I1021818,I1021877,I1021894,I1021920,I1021942,I1021968,I1021976,I1021993,I1022024,I1022099,I1022125,I1022133,I1022150,I1022176,I1022184,I1022201,I1022218,I1022249,I1022280,I1022297,I1022314,I1022331,I1022348,I1022379,I1022438,I1022455,I1022481,I1022503,I1022529,I1022537,I1022554,I1022585,I1022660,I1022686,I1022694,I1022711,I1022737,I1022745,I1022762,I1022779,I1022810,I1022841,I1022858,I1022875,I1022892,I1022909,I1022940,I1022999,I1023016,I1023042,I1023064,I1023090,I1023098,I1023115,I1023146,I1023221,I1023247,I1023255,I1023272,I1023298,I1023306,I1023323,I1023340,I1023371,I1023402,I1023419,I1023436,I1023453,I1023470,I1023501,I1023560,I1023577,I1023603,I1023625,I1023651,I1023659,I1023676,I1023707,I1023782,I1023808,I1023816,I1023833,I1023859,I1023867,I1023884,I1023901,I1023932,I1023963,I1023980,I1023997,I1024014,I1024031,I1024062,I1024121,I1024138,I1024164,I1024186,I1024212,I1024220,I1024237,I1024268,I1024343,I1024369,I1024377,I1024394,I1024420,I1024428,I1024445,I1024462,I1024493,I1024524,I1024541,I1024558,I1024575,I1024592,I1024623,I1024682,I1024699,I1024725,I1024747,I1024773,I1024781,I1024798,I1024829,I1024904,I1024930,I1024938,I1024955,I1024981,I1024989,I1025006,I1025023,I1025054,I1025085,I1025102,I1025119,I1025136,I1025153,I1025184,I1025243,I1025260,I1025286,I1025308,I1025334,I1025342,I1025359,I1025390,I1025465,I1025491,I1025499,I1025516,I1025542,I1025550,I1025567,I1025584,I1025615,I1025646,I1025663,I1025680,I1025697,I1025714,I1025745,I1025804,I1025821,I1025847,I1025869,I1025895,I1025903,I1025920,I1025951,I1026026,I1026052,I1026060,I1026077,I1026103,I1026111,I1026128,I1026145,I1026176,I1026207,I1026224,I1026241,I1026258,I1026275,I1026306,I1026365,I1026382,I1026408,I1026430,I1026456,I1026464,I1026481,I1026512,I1026587,I1026613,I1026621,I1026638,I1026664,I1026672,I1026689,I1026706,I1026737,I1026768,I1026785,I1026802,I1026819,I1026836,I1026867,I1026926,I1026943,I1026969,I1026991,I1027017,I1027025,I1027042,I1027073,I1027148,I1027174,I1027182,I1027199,I1027225,I1027233,I1027250,I1027267,I1027298,I1027329,I1027346,I1027363,I1027380,I1027397,I1027428,I1027487,I1027504,I1027530,I1027552,I1027578,I1027586,I1027603,I1027634,I1027709,I1027735,I1027743,I1027760,I1027786,I1027794,I1027811,I1027828,I1027859,I1027890,I1027907,I1027924,I1027941,I1027958,I1027989,I1028048,I1028065,I1028091,I1028113,I1028139,I1028147,I1028164,I1028195,I1028270,I1028296,I1028304,I1028321,I1028347,I1028355,I1028372,I1028389,I1028420,I1028451,I1028468,I1028485,I1028502,I1028519,I1028550,I1028609,I1028626,I1028652,I1028674,I1028700,I1028708,I1028725,I1028756,I1028831,I1028857,I1028865,I1028882,I1028908,I1028916,I1028933,I1028950,I1028981,I1029012,I1029029,I1029046,I1029063,I1029080,I1029111,I1029170,I1029187,I1029213,I1029235,I1029261,I1029269,I1029286,I1029317,I1029392,I1029418,I1029426,I1029443,I1029469,I1029477,I1029494,I1029511,I1029542,I1029573,I1029590,I1029607,I1029624,I1029641,I1029672,I1029731,I1029748,I1029774,I1029796,I1029822,I1029830,I1029847,I1029878,I1029953,I1029979,I1029987,I1030004,I1030030,I1030038,I1030055,I1030072,I1030103,I1030134,I1030151,I1030168,I1030185,I1030202,I1030233,I1030292,I1030309,I1030335,I1030357,I1030383,I1030391,I1030408,I1030439,I1030514,I1030540,I1030557,I1030565,I1030610,I1030627,I1030644,I1030661,I1030678,I1030695,I1030712,I1030743,I1030760,I1030805,I1030822,I1030839,I1030870,I1030896,I1030904,I1030935,I1030952,I1030969,I1030995,I1031003,I1031020,I1031109,I1031135,I1031152,I1031160,I1031205,I1031222,I1031239,I1031256,I1031273,I1031290,I1031307,I1031338,I1031355,I1031400,I1031417,I1031434,I1031465,I1031491,I1031499,I1031530,I1031547,I1031564,I1031590,I1031598,I1031615,I1031704,I1031730,I1031747,I1031755,I1031800,I1031817,I1031834,I1031851,I1031868,I1031885,I1031902,I1031933,I1031950,I1031995,I1032012,I1032029,I1032060,I1032086,I1032094,I1032125,I1032142,I1032159,I1032185,I1032193,I1032210,I1032299,I1032325,I1032342,I1032350,I1032395,I1032412,I1032429,I1032446,I1032463,I1032480,I1032497,I1032528,I1032545,I1032590,I1032607,I1032624,I1032655,I1032681,I1032689,I1032720,I1032737,I1032754,I1032780,I1032788,I1032805,I1032894,I1032920,I1032937,I1032945,I1032990,I1033007,I1033024,I1033041,I1033058,I1033075,I1033092,I1033123,I1033140,I1033185,I1033202,I1033219,I1033250,I1033276,I1033284,I1033315,I1033332,I1033349,I1033375,I1033383,I1033400,I1033489,I1033515,I1033532,I1033540,I1033585,I1033602,I1033619,I1033636,I1033653,I1033670,I1033687,I1033718,I1033735,I1033780,I1033797,I1033814,I1033845,I1033871,I1033879,I1033910,I1033927,I1033944,I1033970,I1033978,I1033995,I1034084,I1034110,I1034127,I1034135,I1034180,I1034197,I1034214,I1034231,I1034248,I1034265,I1034282,I1034313,I1034330,I1034375,I1034392,I1034409,I1034440,I1034466,I1034474,I1034505,I1034522,I1034539,I1034565,I1034573,I1034590,I1034679,I1034705,I1034722,I1034730,I1034775,I1034792,I1034809,I1034826,I1034843,I1034860,I1034877,I1034908,I1034925,I1034970,I1034987,I1035004,I1035035,I1035061,I1035069,I1035100,I1035117,I1035134,I1035160,I1035168,I1035185,I1035274,I1035300,I1035317,I1035325,I1035370,I1035387,I1035404,I1035421,I1035438,I1035455,I1035472,I1035503,I1035520,I1035565,I1035582,I1035599,I1035630,I1035656,I1035664,I1035695,I1035712,I1035729,I1035755,I1035763,I1035780,I1035869,I1035895,I1035912,I1035920,I1035965,I1035982,I1035999,I1036016,I1036033,I1036050,I1036067,I1036098,I1036115,I1036160,I1036177,I1036194,I1036225,I1036251,I1036259,I1036290,I1036307,I1036324,I1036350,I1036358,I1036375,I1036464,I1036490,I1036507,I1036515,I1036560,I1036577,I1036594,I1036611,I1036628,I1036645,I1036662,I1036693,I1036710,I1036755,I1036772,I1036789,I1036820,I1036846,I1036854,I1036885,I1036902,I1036919,I1036945,I1036953,I1036970,I1037059,I1037085,I1037102,I1037110,I1037155,I1037172,I1037189,I1037206,I1037223,I1037240,I1037257,I1037288,I1037305,I1037350,I1037367,I1037384,I1037415,I1037441,I1037449,I1037480,I1037497,I1037514,I1037540,I1037548,I1037565,I1037654,I1037680,I1037697,I1037705,I1037750,I1037767,I1037784,I1037801,I1037818,I1037835,I1037852,I1037883,I1037900,I1037945,I1037962,I1037979,I1038010,I1038036,I1038044,I1038075,I1038092,I1038109,I1038135,I1038143,I1038160,I1038249,I1038275,I1038292,I1038300,I1038345,I1038362,I1038379,I1038396,I1038413,I1038430,I1038447,I1038478,I1038495,I1038540,I1038557,I1038574,I1038605,I1038631,I1038639,I1038670,I1038687,I1038704,I1038730,I1038738,I1038755,I1038844,I1038870,I1038887,I1038895,I1038940,I1038957,I1038974,I1038991,I1039008,I1039025,I1039042,I1039073,I1039090,I1039135,I1039152,I1039169,I1039200,I1039226,I1039234,I1039265,I1039282,I1039299,I1039325,I1039333,I1039350,I1039439,I1039465,I1039482,I1039490,I1039535,I1039552,I1039569,I1039586,I1039603,I1039620,I1039637,I1039668,I1039685,I1039730,I1039747,I1039764,I1039795,I1039821,I1039829,I1039860,I1039877,I1039894,I1039920,I1039928,I1039945,I1040034,I1040060,I1040077,I1040085,I1040130,I1040147,I1040164,I1040181,I1040198,I1040215,I1040232,I1040263,I1040280,I1040325,I1040342,I1040359,I1040390,I1040416,I1040424,I1040455,I1040472,I1040489,I1040515,I1040523,I1040540,I1040629,I1040655,I1040672,I1040680,I1040725,I1040742,I1040759,I1040776,I1040793,I1040810,I1040827,I1040858,I1040875,I1040920,I1040937,I1040954,I1040985,I1041011,I1041019,I1041050,I1041067,I1041084,I1041110,I1041118,I1041135,I1041224,I1041250,I1041267,I1041275,I1041320,I1041337,I1041354,I1041371,I1041388,I1041405,I1041422,I1041453,I1041470,I1041515,I1041532,I1041549,I1041580,I1041606,I1041614,I1041645,I1041662,I1041679,I1041705,I1041713,I1041730,I1041819,I1041845,I1041862,I1041870,I1041915,I1041932,I1041949,I1041966,I1041983,I1042000,I1042017,I1042048,I1042065,I1042110,I1042127,I1042144,I1042175,I1042201,I1042209,I1042240,I1042257,I1042274,I1042300,I1042308,I1042325,I1042414,I1042440,I1042457,I1042465,I1042510,I1042527,I1042544,I1042561,I1042578,I1042595,I1042612,I1042643,I1042660,I1042705,I1042722,I1042739,I1042770,I1042796,I1042804,I1042835,I1042852,I1042869,I1042895,I1042903,I1042920,I1043009,I1043035,I1043052,I1043060,I1043105,I1043122,I1043139,I1043156,I1043173,I1043190,I1043207,I1043238,I1043255,I1043300,I1043317,I1043334,I1043365,I1043391,I1043399,I1043430,I1043447,I1043464,I1043490,I1043498,I1043515,I1043604,I1043630,I1043647,I1043655,I1043700,I1043717,I1043734,I1043751,I1043768,I1043785,I1043802,I1043833,I1043850,I1043895,I1043912,I1043929,I1043960,I1043986,I1043994,I1044025,I1044042,I1044059,I1044085,I1044093,I1044110,I1044199,I1044225,I1044242,I1044250,I1044295,I1044312,I1044329,I1044346,I1044363,I1044380,I1044397,I1044428,I1044445,I1044490,I1044507,I1044524,I1044555,I1044581,I1044589,I1044620,I1044637,I1044654,I1044680,I1044688,I1044705,I1044794,I1044820,I1044837,I1044845,I1044890,I1044907,I1044924,I1044941,I1044958,I1044975,I1044992,I1045023,I1045040,I1045085,I1045102,I1045119,I1045150,I1045176,I1045184,I1045215,I1045232,I1045249,I1045275,I1045283,I1045300,I1045389,I1045415,I1045432,I1045440,I1045485,I1045502,I1045519,I1045536,I1045553,I1045570,I1045587,I1045618,I1045635,I1045680,I1045697,I1045714,I1045745,I1045771,I1045779,I1045810,I1045827,I1045844,I1045870,I1045878,I1045895,I1045984,I1046010,I1046027,I1046035,I1046080,I1046097,I1046114,I1046131,I1046148,I1046165,I1046182,I1046213,I1046230,I1046275,I1046292,I1046309,I1046340,I1046366,I1046374,I1046405,I1046422,I1046439,I1046465,I1046473,I1046490,I1046579,I1046605,I1046622,I1046630,I1046675,I1046692,I1046709,I1046726,I1046743,I1046760,I1046777,I1046808,I1046825,I1046870,I1046887,I1046904,I1046935,I1046961,I1046969,I1047000,I1047017,I1047034,I1047060,I1047068,I1047085,I1047174,I1047200,I1047217,I1047225,I1047270,I1047287,I1047304,I1047321,I1047338,I1047355,I1047372,I1047403,I1047420,I1047465,I1047482,I1047499,I1047530,I1047556,I1047564,I1047595,I1047612,I1047629,I1047655,I1047663,I1047680,I1047769,I1047795,I1047812,I1047820,I1047865,I1047882,I1047899,I1047916,I1047933,I1047950,I1047967,I1047998,I1048015,I1048060,I1048077,I1048094,I1048125,I1048151,I1048159,I1048190,I1048207,I1048224,I1048250,I1048258,I1048275,I1048364,I1048390,I1048407,I1048415,I1048460,I1048477,I1048494,I1048511,I1048528,I1048545,I1048562,I1048593,I1048610,I1048655,I1048672,I1048689,I1048720,I1048746,I1048754,I1048785,I1048802,I1048819,I1048845,I1048853,I1048870,I1048959,I1048985,I1049002,I1049010,I1049055,I1049072,I1049089,I1049106,I1049123,I1049140,I1049157,I1049188,I1049205,I1049250,I1049267,I1049284,I1049315,I1049341,I1049349,I1049380,I1049397,I1049414,I1049440,I1049448,I1049465,I1049554,I1049580,I1049597,I1049605,I1049650,I1049667,I1049684,I1049701,I1049718,I1049735,I1049752,I1049783,I1049800,I1049845,I1049862,I1049879,I1049910,I1049936,I1049944,I1049975,I1049992,I1050009,I1050035,I1050043,I1050060,I1050149,I1050175,I1050192,I1050200,I1050245,I1050262,I1050279,I1050296,I1050313,I1050330,I1050347,I1050378,I1050395,I1050440,I1050457,I1050474,I1050505,I1050531,I1050539,I1050570,I1050587,I1050604,I1050630,I1050638,I1050655,I1050744,I1050770,I1050787,I1050795,I1050840,I1050857,I1050874,I1050891,I1050908,I1050925,I1050942,I1050973,I1050990,I1051035,I1051052,I1051069,I1051100,I1051126,I1051134,I1051165,I1051182,I1051199,I1051225,I1051233,I1051250,I1051339,I1051365,I1051382,I1051390,I1051435,I1051452,I1051469,I1051486,I1051503,I1051520,I1051537,I1051568,I1051585,I1051630,I1051647,I1051664,I1051695,I1051721,I1051729,I1051760,I1051777,I1051794,I1051820,I1051828,I1051845,I1051934,I1051960,I1051977,I1051985,I1052030,I1052047,I1052064,I1052081,I1052098,I1052115,I1052132,I1052163,I1052180,I1052225,I1052242,I1052259,I1052290,I1052316,I1052324,I1052355,I1052372,I1052389,I1052415,I1052423,I1052440,I1052529,I1052555,I1052572,I1052580,I1052625,I1052642,I1052659,I1052676,I1052693,I1052710,I1052727,I1052758,I1052775,I1052820,I1052837,I1052854,I1052885,I1052911,I1052919,I1052950,I1052967,I1052984,I1053010,I1053018,I1053035,I1053124,I1053150,I1053167,I1053175,I1053220,I1053237,I1053254,I1053271,I1053288,I1053305,I1053322,I1053353,I1053370,I1053415,I1053432,I1053449,I1053480,I1053506,I1053514,I1053545,I1053562,I1053579,I1053605,I1053613,I1053630,I1053719,I1053745,I1053762,I1053770,I1053815,I1053832,I1053849,I1053866,I1053883,I1053900,I1053917,I1053948,I1053965,I1054010,I1054027,I1054044,I1054075,I1054101,I1054109,I1054140,I1054157,I1054174,I1054200,I1054208,I1054225,I1054314,I1054340,I1054357,I1054365,I1054410,I1054427,I1054444,I1054461,I1054478,I1054495,I1054512,I1054543,I1054560,I1054605,I1054622,I1054639,I1054670,I1054696,I1054704,I1054735,I1054752,I1054769,I1054795,I1054803,I1054820,I1054909,I1054935,I1054952,I1054960,I1055005,I1055022,I1055039,I1055056,I1055073,I1055090,I1055107,I1055138,I1055155,I1055200,I1055217,I1055234,I1055265,I1055291,I1055299,I1055330,I1055347,I1055364,I1055390,I1055398,I1055415,I1055504,I1055530,I1055547,I1055555,I1055600,I1055617,I1055634,I1055651,I1055668,I1055685,I1055702,I1055733,I1055750,I1055795,I1055812,I1055829,I1055860,I1055886,I1055894,I1055925,I1055942,I1055959,I1055985,I1055993,I1056010,I1056099,I1056125,I1056142,I1056150,I1056195,I1056212,I1056229,I1056246,I1056263,I1056280,I1056297,I1056328,I1056345,I1056390,I1056407,I1056424,I1056455,I1056481,I1056489,I1056520,I1056537,I1056554,I1056580,I1056588,I1056605,I1056694,I1056720,I1056737,I1056745,I1056790,I1056807,I1056824,I1056841,I1056858,I1056875,I1056892,I1056923,I1056940,I1056985,I1057002,I1057019,I1057050,I1057076,I1057084,I1057115,I1057132,I1057149,I1057175,I1057183,I1057200,I1057289,I1057315,I1057332,I1057340,I1057385,I1057402,I1057419,I1057436,I1057453,I1057470,I1057487,I1057518,I1057535,I1057580,I1057597,I1057614,I1057645,I1057671,I1057679,I1057710,I1057727,I1057744,I1057770,I1057778,I1057795,I1057884,I1057910,I1057927,I1057935,I1057980,I1057997,I1058014,I1058031,I1058048,I1058065,I1058082,I1058113,I1058130,I1058175,I1058192,I1058209,I1058240,I1058266,I1058274,I1058305,I1058322,I1058339,I1058365,I1058373,I1058390,I1058479,I1058505,I1058522,I1058530,I1058575,I1058592,I1058609,I1058626,I1058643,I1058660,I1058677,I1058708,I1058725,I1058770,I1058787,I1058804,I1058835,I1058861,I1058869,I1058900,I1058917,I1058934,I1058960,I1058968,I1058985,I1059074,I1059100,I1059117,I1059125,I1059170,I1059187,I1059204,I1059221,I1059238,I1059255,I1059272,I1059303,I1059320,I1059365,I1059382,I1059399,I1059430,I1059456,I1059464,I1059495,I1059512,I1059529,I1059555,I1059563,I1059580,I1059669,I1059695,I1059712,I1059720,I1059765,I1059782,I1059799,I1059816,I1059833,I1059850,I1059867,I1059898,I1059915,I1059960,I1059977,I1059994,I1060025,I1060051,I1060059,I1060090,I1060107,I1060124,I1060150,I1060158,I1060175,I1060264,I1060290,I1060307,I1060315,I1060360,I1060377,I1060394,I1060411,I1060428,I1060445,I1060462,I1060493,I1060510,I1060555,I1060572,I1060589,I1060620,I1060646,I1060654,I1060685,I1060702,I1060719,I1060745,I1060753,I1060770,I1060859,I1060885,I1060902,I1060910,I1060955,I1060972,I1060989,I1061006,I1061023,I1061040,I1061057,I1061088,I1061105,I1061150,I1061167,I1061184,I1061215,I1061241,I1061249,I1061280,I1061297,I1061314,I1061340,I1061348,I1061365,I1061454,I1061480,I1061497,I1061505,I1061550,I1061567,I1061584,I1061601,I1061618,I1061635,I1061652,I1061683,I1061700,I1061745,I1061762,I1061779,I1061810,I1061836,I1061844,I1061875,I1061892,I1061909,I1061935,I1061943,I1061960,I1062049,I1062075,I1062092,I1062100,I1062145,I1062162,I1062179,I1062196,I1062213,I1062230,I1062247,I1062278,I1062295,I1062340,I1062357,I1062374,I1062405,I1062431,I1062439,I1062470,I1062487,I1062504,I1062530,I1062538,I1062555,I1062644,I1062670,I1062687,I1062695,I1062740,I1062757,I1062774,I1062791,I1062808,I1062825,I1062842,I1062873,I1062890,I1062935,I1062952,I1062969,I1063000,I1063026,I1063034,I1063065,I1063082,I1063099,I1063125,I1063133,I1063150,I1063239,I1063265,I1063282,I1063290,I1063335,I1063352,I1063369,I1063386,I1063403,I1063420,I1063437,I1063468,I1063485,I1063530,I1063547,I1063564,I1063595,I1063621,I1063629,I1063660,I1063677,I1063694,I1063720,I1063728,I1063745,I1063834,I1063860,I1063877,I1063885,I1063930,I1063947,I1063964,I1063981,I1063998,I1064015,I1064032,I1064063,I1064080,I1064125,I1064142,I1064159,I1064190,I1064216,I1064224,I1064255,I1064272,I1064289,I1064315,I1064323,I1064340,I1064429,I1064455,I1064472,I1064480,I1064525,I1064542,I1064559,I1064576,I1064593,I1064610,I1064627,I1064658,I1064675,I1064720,I1064737,I1064754,I1064785,I1064811,I1064819,I1064850,I1064867,I1064884,I1064910,I1064918,I1064935,I1065024,I1065050,I1065067,I1065075,I1065120,I1065137,I1065154,I1065171,I1065188,I1065205,I1065222,I1065253,I1065270,I1065315,I1065332,I1065349,I1065380,I1065406,I1065414,I1065445,I1065462,I1065479,I1065505,I1065513,I1065530,I1065619,I1065645,I1065662,I1065670,I1065715,I1065732,I1065749,I1065766,I1065783,I1065800,I1065817,I1065848,I1065865,I1065910,I1065927,I1065944,I1065975,I1066001,I1066009,I1066040,I1066057,I1066074,I1066100,I1066108,I1066125,I1066214,I1066240,I1066257,I1066265,I1066310,I1066327,I1066344,I1066361,I1066378,I1066395,I1066412,I1066443,I1066460,I1066505,I1066522,I1066539,I1066570,I1066596,I1066604,I1066635,I1066652,I1066669,I1066695,I1066703,I1066720,I1066809,I1066835,I1066852,I1066860,I1066905,I1066922,I1066939,I1066956,I1066973,I1066990,I1067007,I1067038,I1067055,I1067100,I1067117,I1067134,I1067165,I1067191,I1067199,I1067230,I1067247,I1067264,I1067290,I1067298,I1067315,I1067404,I1067430,I1067447,I1067455,I1067500,I1067517,I1067534,I1067551,I1067568,I1067585,I1067602,I1067633,I1067650,I1067695,I1067712,I1067729,I1067760,I1067786,I1067794,I1067825,I1067842,I1067859,I1067885,I1067893,I1067910,I1067999,I1068025,I1068042,I1068050,I1068095,I1068112,I1068129,I1068146,I1068163,I1068180,I1068197,I1068228,I1068245,I1068290,I1068307,I1068324,I1068355,I1068381,I1068389,I1068420,I1068437,I1068454,I1068480,I1068488,I1068505,I1068594,I1068620,I1068637,I1068645,I1068690,I1068707,I1068724,I1068741,I1068758,I1068775,I1068792,I1068823,I1068840,I1068885,I1068902,I1068919,I1068950,I1068976,I1068984,I1069015,I1069032,I1069049,I1069075,I1069083,I1069100,I1069189,I1069215,I1069232,I1069240,I1069285,I1069302,I1069319,I1069336,I1069353,I1069370,I1069387,I1069418,I1069435,I1069480,I1069497,I1069514,I1069545,I1069571,I1069579,I1069610,I1069627,I1069644,I1069670,I1069678,I1069695,I1069784,I1069810,I1069827,I1069835,I1069880,I1069897,I1069914,I1069931,I1069948,I1069965,I1069982,I1070013,I1070030,I1070075,I1070092,I1070109,I1070140,I1070166,I1070174,I1070205,I1070222,I1070239,I1070265,I1070273,I1070290,I1070379,I1070405,I1070422,I1070430,I1070475,I1070492,I1070509,I1070526,I1070543,I1070560,I1070577,I1070608,I1070625,I1070670,I1070687,I1070704,I1070735,I1070761,I1070769,I1070800,I1070817,I1070834,I1070860,I1070868,I1070885,I1070974,I1071000,I1071017,I1071025,I1071070,I1071087,I1071104,I1071121,I1071138,I1071155,I1071172,I1071203,I1071220,I1071265,I1071282,I1071299,I1071330,I1071356,I1071364,I1071395,I1071412,I1071429,I1071455,I1071463,I1071480,I1071569,I1071595,I1071612,I1071620,I1071665,I1071682,I1071699,I1071716,I1071733,I1071750,I1071767,I1071798,I1071815,I1071860,I1071877,I1071894,I1071925,I1071951,I1071959,I1071990,I1072007,I1072024,I1072050,I1072058,I1072075,I1072164,I1072190,I1072207,I1072215,I1072260,I1072277,I1072294,I1072311,I1072328,I1072345,I1072362,I1072393,I1072410,I1072455,I1072472,I1072489,I1072520,I1072546,I1072554,I1072585,I1072602,I1072619,I1072645,I1072653,I1072670,I1072759,I1072785,I1072802,I1072810,I1072855,I1072872,I1072889,I1072906,I1072923,I1072940,I1072957,I1072988,I1073005,I1073050,I1073067,I1073084,I1073115,I1073141,I1073149,I1073180,I1073197,I1073214,I1073240,I1073248,I1073265,I1073354,I1073380,I1073397,I1073405,I1073450,I1073467,I1073484,I1073501,I1073518,I1073535,I1073552,I1073583,I1073600,I1073645,I1073662,I1073679,I1073710,I1073736,I1073744,I1073775,I1073792,I1073809,I1073835,I1073843,I1073860,I1073949,I1073975,I1073992,I1074000,I1074045,I1074062,I1074079,I1074096,I1074113,I1074130,I1074147,I1074178,I1074195,I1074240,I1074257,I1074274,I1074305,I1074331,I1074339,I1074370,I1074387,I1074404,I1074430,I1074438,I1074455,I1074544,I1074570,I1074587,I1074595,I1074640,I1074657,I1074674,I1074691,I1074708,I1074725,I1074742,I1074773,I1074790,I1074835,I1074852,I1074869,I1074900,I1074926,I1074934,I1074965,I1074982,I1074999,I1075025,I1075033,I1075050,I1075139,I1075165,I1075182,I1075190,I1075235,I1075252,I1075269,I1075286,I1075303,I1075320,I1075337,I1075368,I1075385,I1075430,I1075447,I1075464,I1075495,I1075521,I1075529,I1075560,I1075577,I1075594,I1075620,I1075628,I1075645,I1075734,I1075760,I1075777,I1075785,I1075830,I1075847,I1075864,I1075881,I1075898,I1075915,I1075932,I1075963,I1075980,I1076025,I1076042,I1076059,I1076090,I1076116,I1076124,I1076155,I1076172,I1076189,I1076215,I1076223,I1076240,I1076329,I1076355,I1076372,I1076380,I1076425,I1076442,I1076459,I1076476,I1076493,I1076510,I1076527,I1076558,I1076575,I1076620,I1076637,I1076654,I1076685,I1076711,I1076719,I1076750,I1076767,I1076784,I1076810,I1076818,I1076835,I1076924,I1076950,I1076967,I1076975,I1077020,I1077037,I1077054,I1077071,I1077088,I1077105,I1077122,I1077153,I1077170,I1077215,I1077232,I1077249,I1077280,I1077306,I1077314,I1077345,I1077362,I1077379,I1077405,I1077413,I1077430,I1077519,I1077545,I1077562,I1077570,I1077615,I1077632,I1077649,I1077666,I1077683,I1077700,I1077717,I1077748,I1077765,I1077810,I1077827,I1077844,I1077875,I1077901,I1077909,I1077940,I1077957,I1077974,I1078000,I1078008,I1078025,I1078114,I1078140,I1078157,I1078165,I1078210,I1078227,I1078244,I1078261,I1078278,I1078295,I1078312,I1078343,I1078360,I1078405,I1078422,I1078439,I1078470,I1078496,I1078504,I1078535,I1078552,I1078569,I1078595,I1078603,I1078620,I1078709,I1078735,I1078752,I1078760,I1078805,I1078822,I1078839,I1078856,I1078873,I1078890,I1078907,I1078938,I1078955,I1079000,I1079017,I1079034,I1079065,I1079091,I1079099,I1079130,I1079147,I1079164,I1079190,I1079198,I1079215,I1079304,I1079330,I1079347,I1079355,I1079400,I1079417,I1079434,I1079451,I1079468,I1079485,I1079502,I1079533,I1079550,I1079595,I1079612,I1079629,I1079660,I1079686,I1079694,I1079725,I1079742,I1079759,I1079785,I1079793,I1079810,I1079899,I1079925,I1079942,I1079950,I1079995,I1080012,I1080029,I1080046,I1080063,I1080080,I1080097,I1080128,I1080145,I1080190,I1080207,I1080224,I1080255,I1080281,I1080289,I1080320,I1080337,I1080354,I1080380,I1080388,I1080405,I1080494,I1080520,I1080537,I1080545,I1080590,I1080607,I1080624,I1080641,I1080658,I1080675,I1080692,I1080723,I1080740,I1080785,I1080802,I1080819,I1080850,I1080876,I1080884,I1080915,I1080932,I1080949,I1080975,I1080983,I1081000,I1081089,I1081115,I1081132,I1081140,I1081185,I1081202,I1081219,I1081236,I1081253,I1081270,I1081287,I1081318,I1081335,I1081380,I1081397,I1081414,I1081445,I1081471,I1081479,I1081510,I1081527,I1081544,I1081570,I1081578,I1081595,I1081684,I1081710,I1081727,I1081735,I1081780,I1081797,I1081814,I1081831,I1081848,I1081865,I1081882,I1081913,I1081930,I1081975,I1081992,I1082009,I1082040,I1082066,I1082074,I1082105,I1082122,I1082139,I1082165,I1082173,I1082190,I1082279,I1082305,I1082322,I1082330,I1082375,I1082392,I1082409,I1082426,I1082443,I1082460,I1082477,I1082508,I1082525,I1082570,I1082587,I1082604,I1082635,I1082661,I1082669,I1082700,I1082717,I1082734,I1082760,I1082768,I1082785,I1082874,I1082900,I1082917,I1082925,I1082970,I1082987,I1083004,I1083021,I1083038,I1083055,I1083072,I1083103,I1083120,I1083165,I1083182,I1083199,I1083230,I1083256,I1083264,I1083295,I1083312,I1083329,I1083355,I1083363,I1083380,I1083469,I1083495,I1083512,I1083520,I1083565,I1083582,I1083599,I1083616,I1083633,I1083650,I1083667,I1083698,I1083715,I1083760,I1083777,I1083794,I1083825,I1083851,I1083859,I1083890,I1083907,I1083924,I1083950,I1083958,I1083975,I1084064,I1084090,I1084107,I1084115,I1084160,I1084177,I1084194,I1084211,I1084228,I1084245,I1084262,I1084293,I1084310,I1084355,I1084372,I1084389,I1084420,I1084446,I1084454,I1084485,I1084502,I1084519,I1084545,I1084553,I1084570,I1084659,I1084685,I1084702,I1084710,I1084755,I1084772,I1084789,I1084806,I1084823,I1084840,I1084857,I1084888,I1084905,I1084950,I1084967,I1084984,I1085015,I1085041,I1085049,I1085080,I1085097,I1085114,I1085140,I1085148,I1085165,I1085254,I1085280,I1085297,I1085305,I1085350,I1085367,I1085384,I1085401,I1085418,I1085435,I1085452,I1085483,I1085500,I1085545,I1085562,I1085579,I1085610,I1085636,I1085644,I1085675,I1085692,I1085709,I1085735,I1085743,I1085760,I1085849,I1085875,I1085892,I1085900,I1085945,I1085962,I1085979,I1085996,I1086013,I1086030,I1086047,I1086078,I1086095,I1086140,I1086157,I1086174,I1086205,I1086231,I1086239,I1086270,I1086287,I1086304,I1086330,I1086338,I1086355,I1086444,I1086470,I1086487,I1086495,I1086540,I1086557,I1086574,I1086591,I1086608,I1086625,I1086642,I1086673,I1086690,I1086735,I1086752,I1086769,I1086800,I1086826,I1086834,I1086865,I1086882,I1086899,I1086925,I1086933,I1086950,I1087039,I1087065,I1087082,I1087090,I1087135,I1087152,I1087169,I1087186,I1087203,I1087220,I1087237,I1087268,I1087285,I1087330,I1087347,I1087364,I1087395,I1087421,I1087429,I1087460,I1087477,I1087494,I1087520,I1087528,I1087545,I1087634,I1087660,I1087677,I1087685,I1087730,I1087747,I1087764,I1087781,I1087798,I1087815,I1087832,I1087863,I1087880,I1087925,I1087942,I1087959,I1087990,I1088016,I1088024,I1088055,I1088072,I1088089,I1088115,I1088123,I1088140,I1088229,I1088255,I1088272,I1088280,I1088325,I1088342,I1088359,I1088376,I1088393,I1088410,I1088427,I1088458,I1088475,I1088520,I1088537,I1088554,I1088585,I1088611,I1088619,I1088650,I1088667,I1088684,I1088710,I1088718,I1088735,I1088824,I1088850,I1088867,I1088875,I1088920,I1088937,I1088954,I1088971,I1088988,I1089005,I1089022,I1089053,I1089070,I1089115,I1089132,I1089149,I1089180,I1089206,I1089214,I1089245,I1089262,I1089279,I1089305,I1089313,I1089330,I1089419,I1089445,I1089462,I1089470,I1089515,I1089532,I1089549,I1089566,I1089583,I1089600,I1089617,I1089648,I1089665,I1089710,I1089727,I1089744,I1089775,I1089801,I1089809,I1089840,I1089857,I1089874,I1089900,I1089908,I1089925,I1090014,I1090040,I1090057,I1090065,I1090110,I1090127,I1090144,I1090161,I1090178,I1090195,I1090212,I1090243,I1090260,I1090305,I1090322,I1090339,I1090370,I1090396,I1090404,I1090435,I1090452,I1090469,I1090495,I1090503,I1090520,I1090609,I1090635,I1090652,I1090660,I1090705,I1090722,I1090739,I1090756,I1090773,I1090790,I1090807,I1090838,I1090855,I1090900,I1090917,I1090934,I1090965,I1090991,I1090999,I1091030,I1091047,I1091064,I1091090,I1091098,I1091115,I1091204,I1091230,I1091247,I1091255,I1091300,I1091317,I1091334,I1091351,I1091368,I1091385,I1091402,I1091433,I1091450,I1091495,I1091512,I1091529,I1091560,I1091586,I1091594,I1091625,I1091642,I1091659,I1091685,I1091693,I1091710,I1091799,I1091825,I1091842,I1091850,I1091895,I1091912,I1091929,I1091946,I1091963,I1091980,I1091997,I1092028,I1092045,I1092090,I1092107,I1092124,I1092155,I1092181,I1092189,I1092220,I1092237,I1092254,I1092280,I1092288,I1092305,I1092394,I1092420,I1092437,I1092445,I1092490,I1092507,I1092524,I1092541,I1092558,I1092575,I1092592,I1092623,I1092640,I1092685,I1092702,I1092719,I1092750,I1092776,I1092784,I1092815,I1092832,I1092849,I1092875,I1092883,I1092900,I1092989,I1093015,I1093032,I1093040,I1093085,I1093102,I1093119,I1093136,I1093153,I1093170,I1093187,I1093218,I1093235,I1093280,I1093297,I1093314,I1093345,I1093371,I1093379,I1093410,I1093427,I1093444,I1093470,I1093478,I1093495,I1093584,I1093610,I1093627,I1093635,I1093680,I1093697,I1093714,I1093731,I1093748,I1093765,I1093782,I1093813,I1093830,I1093875,I1093892,I1093909,I1093940,I1093966,I1093974,I1094005,I1094022,I1094039,I1094065,I1094073,I1094090,I1094179,I1094205,I1094222,I1094230,I1094275,I1094292,I1094309,I1094326,I1094343,I1094360,I1094377,I1094408,I1094425,I1094470,I1094487,I1094504,I1094535,I1094561,I1094569,I1094600,I1094617,I1094634,I1094660,I1094668,I1094685,I1094774,I1094800,I1094817,I1094825,I1094870,I1094887,I1094904,I1094921,I1094938,I1094955,I1094972,I1095003,I1095020,I1095065,I1095082,I1095099,I1095130,I1095156,I1095164,I1095195,I1095212,I1095229,I1095255,I1095263,I1095280,I1095369,I1095395,I1095412,I1095420,I1095465,I1095482,I1095499,I1095516,I1095533,I1095550,I1095567,I1095598,I1095615,I1095660,I1095677,I1095694,I1095725,I1095751,I1095759,I1095790,I1095807,I1095824,I1095850,I1095858,I1095875,I1095964,I1095990,I1096007,I1096015,I1096060,I1096077,I1096094,I1096111,I1096128,I1096145,I1096162,I1096193,I1096210,I1096255,I1096272,I1096289,I1096320,I1096346,I1096354,I1096385,I1096402,I1096419,I1096445,I1096453,I1096470,I1096559,I1096585,I1096602,I1096610,I1096655,I1096672,I1096689,I1096706,I1096723,I1096740,I1096757,I1096788,I1096805,I1096850,I1096867,I1096884,I1096915,I1096941,I1096949,I1096980,I1096997,I1097014,I1097040,I1097048,I1097065,I1097154,I1097180,I1097197,I1097205,I1097250,I1097267,I1097284,I1097301,I1097318,I1097335,I1097352,I1097383,I1097400,I1097445,I1097462,I1097479,I1097510,I1097536,I1097544,I1097575,I1097592,I1097609,I1097635,I1097643,I1097660,I1097749,I1097775,I1097792,I1097800,I1097845,I1097862,I1097879,I1097896,I1097913,I1097930,I1097947,I1097978,I1097995,I1098040,I1098057,I1098074,I1098105,I1098131,I1098139,I1098170,I1098187,I1098204,I1098230,I1098238,I1098255,I1098344,I1098370,I1098387,I1098395,I1098440,I1098457,I1098474,I1098491,I1098508,I1098525,I1098542,I1098573,I1098590,I1098635,I1098652,I1098669,I1098700,I1098726,I1098734,I1098765,I1098782,I1098799,I1098825,I1098833,I1098850,I1098939,I1098965,I1098982,I1098990,I1099035,I1099052,I1099069,I1099086,I1099103,I1099120,I1099137,I1099168,I1099185,I1099230,I1099247,I1099264,I1099295,I1099321,I1099329,I1099360,I1099377,I1099394,I1099420,I1099428,I1099445,I1099534,I1099560,I1099577,I1099585,I1099630,I1099647,I1099664,I1099681,I1099698,I1099715,I1099732,I1099763,I1099780,I1099825,I1099842,I1099859,I1099890,I1099916,I1099924,I1099955,I1099972,I1099989,I1100015,I1100023,I1100040,I1100129,I1100155,I1100172,I1100180,I1100225,I1100242,I1100259,I1100276,I1100293,I1100310,I1100327,I1100358,I1100375,I1100420,I1100437,I1100454,I1100485,I1100511,I1100519,I1100550,I1100567,I1100584,I1100610,I1100618,I1100635,I1100724,I1100750,I1100767,I1100775,I1100820,I1100837,I1100854,I1100871,I1100888,I1100905,I1100922,I1100953,I1100970,I1101015,I1101032,I1101049,I1101080,I1101106,I1101114,I1101145,I1101162,I1101179,I1101205,I1101213,I1101230,I1101319,I1101345,I1101362,I1101370,I1101415,I1101432,I1101449,I1101466,I1101483,I1101500,I1101517,I1101548,I1101565,I1101610,I1101627,I1101644,I1101675,I1101701,I1101709,I1101740,I1101757,I1101774,I1101800,I1101808,I1101825;
not I_0 (I2722,I2690);
DFFARX1 I_1 (I630172,I2683,I2722,I2748,);
nand I_2 (I2756,I2748,I630163);
not I_3 (I2773,I2756);
DFFARX1 I_4 (I2773,I2683,I2722,I2714,);
DFFARX1 I_5 (I630169,I2683,I2722,I2813,);
not I_6 (I2821,I2813);
not I_7 (I2838,I630163);
not I_8 (I2855,I630175);
nand I_9 (I2872,I2821,I2855);
nor I_10 (I2889,I2872,I630163);
DFFARX1 I_11 (I2889,I2683,I2722,I2693,);
nor I_12 (I2920,I630175,I630163);
nand I_13 (I2937,I2813,I2920);
nor I_14 (I2954,I630184,I630181);
nor I_15 (I2696,I2872,I630184);
not I_16 (I2985,I630184);
not I_17 (I3002,I630169);
nand I_18 (I3019,I3002,I630166);
nand I_19 (I3036,I2838,I3019);
not I_20 (I3053,I3036);
nor I_21 (I3070,I630169,I630181);
nor I_22 (I2705,I3053,I3070);
nor I_23 (I3101,I630166,I630169);
and I_24 (I3118,I3101,I2954);
nor I_25 (I3135,I3036,I3118);
DFFARX1 I_26 (I3135,I2683,I2722,I2711,);
nor I_27 (I3166,I2756,I3118);
DFFARX1 I_28 (I3166,I2683,I2722,I2708,);
nor I_29 (I3197,I630166,I630178);
DFFARX1 I_30 (I3197,I2683,I2722,I3223,);
nor I_31 (I3231,I3223,I630175);
nand I_32 (I3248,I3231,I2838);
nand I_33 (I2702,I3248,I2937);
nand I_34 (I2699,I3231,I2985);
not I_35 (I3317,I2690);
DFFARX1 I_36 (I600046,I2683,I3317,I3343,);
nand I_37 (I3351,I3343,I600025);
not I_38 (I3368,I3351);
DFFARX1 I_39 (I3368,I2683,I3317,I3309,);
DFFARX1 I_40 (I600034,I2683,I3317,I3408,);
not I_41 (I3416,I3408);
not I_42 (I3433,I600040);
not I_43 (I3450,I600037);
nand I_44 (I3467,I3416,I3450);
nor I_45 (I3484,I3467,I600040);
DFFARX1 I_46 (I3484,I2683,I3317,I3288,);
nor I_47 (I3515,I600037,I600040);
nand I_48 (I3532,I3408,I3515);
nor I_49 (I3549,I600028,I600022);
nor I_50 (I3291,I3467,I600028);
not I_51 (I3580,I600028);
not I_52 (I3597,I600043);
nand I_53 (I3614,I3597,I600025);
nand I_54 (I3631,I3433,I3614);
not I_55 (I3648,I3631);
nor I_56 (I3665,I600043,I600022);
nor I_57 (I3300,I3648,I3665);
nor I_58 (I3696,I600031,I600043);
and I_59 (I3713,I3696,I3549);
nor I_60 (I3730,I3631,I3713);
DFFARX1 I_61 (I3730,I2683,I3317,I3306,);
nor I_62 (I3761,I3351,I3713);
DFFARX1 I_63 (I3761,I2683,I3317,I3303,);
nor I_64 (I3792,I600031,I600022);
DFFARX1 I_65 (I3792,I2683,I3317,I3818,);
nor I_66 (I3826,I3818,I600037);
nand I_67 (I3843,I3826,I3433);
nand I_68 (I3297,I3843,I3532);
nand I_69 (I3294,I3826,I3580);
not I_70 (I3912,I2690);
DFFARX1 I_71 (I1025430,I2683,I3912,I3938,);
nand I_72 (I3946,I3938,I1025439);
not I_73 (I3963,I3946);
DFFARX1 I_74 (I3963,I2683,I3912,I3904,);
DFFARX1 I_75 (I1025445,I2683,I3912,I4003,);
not I_76 (I4011,I4003);
not I_77 (I4028,I1025433);
not I_78 (I4045,I1025442);
nand I_79 (I4062,I4011,I4045);
nor I_80 (I4079,I4062,I1025433);
DFFARX1 I_81 (I4079,I2683,I3912,I3883,);
nor I_82 (I4110,I1025442,I1025433);
nand I_83 (I4127,I4003,I4110);
nor I_84 (I4144,I1025451,I1025448);
nor I_85 (I3886,I4062,I1025451);
not I_86 (I4175,I1025451);
not I_87 (I4192,I1025436);
nand I_88 (I4209,I4192,I1025454);
nand I_89 (I4226,I4028,I4209);
not I_90 (I4243,I4226);
nor I_91 (I4260,I1025436,I1025448);
nor I_92 (I3895,I4243,I4260);
nor I_93 (I4291,I1025430,I1025436);
and I_94 (I4308,I4291,I4144);
nor I_95 (I4325,I4226,I4308);
DFFARX1 I_96 (I4325,I2683,I3912,I3901,);
nor I_97 (I4356,I3946,I4308);
DFFARX1 I_98 (I4356,I2683,I3912,I3898,);
nor I_99 (I4387,I1025430,I1025457);
DFFARX1 I_100 (I4387,I2683,I3912,I4413,);
nor I_101 (I4421,I4413,I1025442);
nand I_102 (I4438,I4421,I4028);
nand I_103 (I3892,I4438,I4127);
nand I_104 (I3889,I4421,I4175);
not I_105 (I4507,I2690);
DFFARX1 I_106 (I482691,I2683,I4507,I4533,);
nand I_107 (I4541,I4533,I482709);
not I_108 (I4558,I4541);
DFFARX1 I_109 (I4558,I2683,I4507,I4499,);
DFFARX1 I_110 (I482703,I2683,I4507,I4598,);
not I_111 (I4606,I4598);
not I_112 (I4623,I482694);
not I_113 (I4640,I482691);
nand I_114 (I4657,I4606,I4640);
nor I_115 (I4674,I4657,I482694);
DFFARX1 I_116 (I4674,I2683,I4507,I4478,);
nor I_117 (I4705,I482691,I482694);
nand I_118 (I4722,I4598,I4705);
nor I_119 (I4739,I482700,I482688);
nor I_120 (I4481,I4657,I482700);
not I_121 (I4770,I482700);
not I_122 (I4787,I482706);
nand I_123 (I4804,I4787,I482712);
nand I_124 (I4821,I4623,I4804);
not I_125 (I4838,I4821);
nor I_126 (I4855,I482706,I482688);
nor I_127 (I4490,I4838,I4855);
nor I_128 (I4886,I482688,I482706);
and I_129 (I4903,I4886,I4739);
nor I_130 (I4920,I4821,I4903);
DFFARX1 I_131 (I4920,I2683,I4507,I4496,);
nor I_132 (I4951,I4541,I4903);
DFFARX1 I_133 (I4951,I2683,I4507,I4493,);
nor I_134 (I4982,I482688,I482697);
DFFARX1 I_135 (I4982,I2683,I4507,I5008,);
nor I_136 (I5016,I5008,I482691);
nand I_137 (I5033,I5016,I4623);
nand I_138 (I4487,I5033,I4722);
nand I_139 (I4484,I5016,I4770);
not I_140 (I5102,I2690);
DFFARX1 I_141 (I527218,I2683,I5102,I5128,);
nand I_142 (I5136,I5128,I527197);
not I_143 (I5153,I5136);
DFFARX1 I_144 (I5153,I2683,I5102,I5094,);
DFFARX1 I_145 (I527206,I2683,I5102,I5193,);
not I_146 (I5201,I5193);
not I_147 (I5218,I527212);
not I_148 (I5235,I527209);
nand I_149 (I5252,I5201,I5235);
nor I_150 (I5269,I5252,I527212);
DFFARX1 I_151 (I5269,I2683,I5102,I5073,);
nor I_152 (I5300,I527209,I527212);
nand I_153 (I5317,I5193,I5300);
nor I_154 (I5334,I527200,I527194);
nor I_155 (I5076,I5252,I527200);
not I_156 (I5365,I527200);
not I_157 (I5382,I527215);
nand I_158 (I5399,I5382,I527197);
nand I_159 (I5416,I5218,I5399);
not I_160 (I5433,I5416);
nor I_161 (I5450,I527215,I527194);
nor I_162 (I5085,I5433,I5450);
nor I_163 (I5481,I527203,I527215);
and I_164 (I5498,I5481,I5334);
nor I_165 (I5515,I5416,I5498);
DFFARX1 I_166 (I5515,I2683,I5102,I5091,);
nor I_167 (I5546,I5136,I5498);
DFFARX1 I_168 (I5546,I2683,I5102,I5088,);
nor I_169 (I5577,I527203,I527194);
DFFARX1 I_170 (I5577,I2683,I5102,I5603,);
nor I_171 (I5611,I5603,I527209);
nand I_172 (I5628,I5611,I5218);
nand I_173 (I5082,I5628,I5317);
nand I_174 (I5079,I5611,I5365);
not I_175 (I5697,I2690);
DFFARX1 I_176 (I388359,I2683,I5697,I5723,);
nand I_177 (I5731,I5723,I388341);
not I_178 (I5748,I5731);
DFFARX1 I_179 (I5748,I2683,I5697,I5689,);
DFFARX1 I_180 (I388353,I2683,I5697,I5788,);
not I_181 (I5796,I5788);
not I_182 (I5813,I388338);
not I_183 (I5830,I388347);
nand I_184 (I5847,I5796,I5830);
nor I_185 (I5864,I5847,I388338);
DFFARX1 I_186 (I5864,I2683,I5697,I5668,);
nor I_187 (I5895,I388347,I388338);
nand I_188 (I5912,I5788,I5895);
nor I_189 (I5929,I388344,I388365);
nor I_190 (I5671,I5847,I388344);
not I_191 (I5960,I388344);
not I_192 (I5977,I388356);
nand I_193 (I5994,I5977,I388362);
nand I_194 (I6011,I5813,I5994);
not I_195 (I6028,I6011);
nor I_196 (I6045,I388356,I388365);
nor I_197 (I5680,I6028,I6045);
nor I_198 (I6076,I388338,I388356);
and I_199 (I6093,I6076,I5929);
nor I_200 (I6110,I6011,I6093);
DFFARX1 I_201 (I6110,I2683,I5697,I5686,);
nor I_202 (I6141,I5731,I6093);
DFFARX1 I_203 (I6141,I2683,I5697,I5683,);
nor I_204 (I6172,I388338,I388350);
DFFARX1 I_205 (I6172,I2683,I5697,I6198,);
nor I_206 (I6206,I6198,I388347);
nand I_207 (I6223,I6206,I5813);
nand I_208 (I5677,I6223,I5912);
nand I_209 (I5674,I6206,I5960);
not I_210 (I6292,I2690);
DFFARX1 I_211 (I74343,I2683,I6292,I6318,);
nand I_212 (I6326,I6318,I74334);
not I_213 (I6343,I6326);
DFFARX1 I_214 (I6343,I2683,I6292,I6284,);
DFFARX1 I_215 (I74355,I2683,I6292,I6383,);
not I_216 (I6391,I6383);
not I_217 (I6408,I74331);
not I_218 (I6425,I74331);
nand I_219 (I6442,I6391,I6425);
nor I_220 (I6459,I6442,I74331);
DFFARX1 I_221 (I6459,I2683,I6292,I6263,);
nor I_222 (I6490,I74331,I74331);
nand I_223 (I6507,I6383,I6490);
nor I_224 (I6524,I74340,I74334);
nor I_225 (I6266,I6442,I74340);
not I_226 (I6555,I74340);
not I_227 (I6572,I74352);
nand I_228 (I6589,I6572,I74349);
nand I_229 (I6606,I6408,I6589);
not I_230 (I6623,I6606);
nor I_231 (I6640,I74352,I74334);
nor I_232 (I6275,I6623,I6640);
nor I_233 (I6671,I74346,I74352);
and I_234 (I6688,I6671,I6524);
nor I_235 (I6705,I6606,I6688);
DFFARX1 I_236 (I6705,I2683,I6292,I6281,);
nor I_237 (I6736,I6326,I6688);
DFFARX1 I_238 (I6736,I2683,I6292,I6278,);
nor I_239 (I6767,I74346,I74337);
DFFARX1 I_240 (I6767,I2683,I6292,I6793,);
nor I_241 (I6801,I6793,I74331);
nand I_242 (I6818,I6801,I6408);
nand I_243 (I6272,I6818,I6507);
nand I_244 (I6269,I6801,I6555);
not I_245 (I6887,I2690);
DFFARX1 I_246 (I287016,I2683,I6887,I6913,);
nand I_247 (I6921,I6913,I287007);
not I_248 (I6938,I6921);
DFFARX1 I_249 (I6938,I2683,I6887,I6879,);
DFFARX1 I_250 (I287010,I2683,I6887,I6978,);
not I_251 (I6986,I6978);
not I_252 (I7003,I287004);
not I_253 (I7020,I287013);
nand I_254 (I7037,I6986,I7020);
nor I_255 (I7054,I7037,I287004);
DFFARX1 I_256 (I7054,I2683,I6887,I6858,);
nor I_257 (I7085,I287013,I287004);
nand I_258 (I7102,I6978,I7085);
nor I_259 (I7119,I287001,I287019);
nor I_260 (I6861,I7037,I287001);
not I_261 (I7150,I287001);
not I_262 (I7167,I287001);
nand I_263 (I7184,I7167,I287025);
nand I_264 (I7201,I7003,I7184);
not I_265 (I7218,I7201);
nor I_266 (I7235,I287001,I287019);
nor I_267 (I6870,I7218,I7235);
nor I_268 (I7266,I287022,I287001);
and I_269 (I7283,I7266,I7119);
nor I_270 (I7300,I7201,I7283);
DFFARX1 I_271 (I7300,I2683,I6887,I6876,);
nor I_272 (I7331,I6921,I7283);
DFFARX1 I_273 (I7331,I2683,I6887,I6873,);
nor I_274 (I7362,I287022,I287028);
DFFARX1 I_275 (I7362,I2683,I6887,I7388,);
nor I_276 (I7396,I7388,I287013);
nand I_277 (I7413,I7396,I7003);
nand I_278 (I6867,I7413,I7102);
nand I_279 (I6864,I7396,I7150);
not I_280 (I7482,I2690);
DFFARX1 I_281 (I364967,I2683,I7482,I7508,);
nand I_282 (I7516,I7508,I364949);
not I_283 (I7533,I7516);
DFFARX1 I_284 (I7533,I2683,I7482,I7474,);
DFFARX1 I_285 (I364961,I2683,I7482,I7573,);
not I_286 (I7581,I7573);
not I_287 (I7598,I364946);
not I_288 (I7615,I364955);
nand I_289 (I7632,I7581,I7615);
nor I_290 (I7649,I7632,I364946);
DFFARX1 I_291 (I7649,I2683,I7482,I7453,);
nor I_292 (I7680,I364955,I364946);
nand I_293 (I7697,I7573,I7680);
nor I_294 (I7714,I364952,I364973);
nor I_295 (I7456,I7632,I364952);
not I_296 (I7745,I364952);
not I_297 (I7762,I364964);
nand I_298 (I7779,I7762,I364970);
nand I_299 (I7796,I7598,I7779);
not I_300 (I7813,I7796);
nor I_301 (I7830,I364964,I364973);
nor I_302 (I7465,I7813,I7830);
nor I_303 (I7861,I364946,I364964);
and I_304 (I7878,I7861,I7714);
nor I_305 (I7895,I7796,I7878);
DFFARX1 I_306 (I7895,I2683,I7482,I7471,);
nor I_307 (I7926,I7516,I7878);
DFFARX1 I_308 (I7926,I2683,I7482,I7468,);
nor I_309 (I7957,I364946,I364958);
DFFARX1 I_310 (I7957,I2683,I7482,I7983,);
nor I_311 (I7991,I7983,I364955);
nand I_312 (I8008,I7991,I7598);
nand I_313 (I7462,I8008,I7697);
nand I_314 (I7459,I7991,I7745);
not I_315 (I8077,I2690);
DFFARX1 I_316 (I1038229,I2683,I8077,I8103,);
nand I_317 (I8111,I8103,I1038220);
not I_318 (I8128,I8111);
DFFARX1 I_319 (I8128,I2683,I8077,I8069,);
DFFARX1 I_320 (I1038223,I2683,I8077,I8168,);
not I_321 (I8176,I8168);
not I_322 (I8193,I1038235);
not I_323 (I8210,I1038226);
nand I_324 (I8227,I8176,I8210);
nor I_325 (I8244,I8227,I1038235);
DFFARX1 I_326 (I8244,I2683,I8077,I8048,);
nor I_327 (I8275,I1038226,I1038235);
nand I_328 (I8292,I8168,I8275);
nor I_329 (I8309,I1038214,I1038214);
nor I_330 (I8051,I8227,I1038214);
not I_331 (I8340,I1038214);
not I_332 (I8357,I1038238);
nand I_333 (I8374,I8357,I1038217);
nand I_334 (I8391,I8193,I8374);
not I_335 (I8408,I8391);
nor I_336 (I8425,I1038238,I1038214);
nor I_337 (I8060,I8408,I8425);
nor I_338 (I8456,I1038232,I1038238);
and I_339 (I8473,I8456,I8309);
nor I_340 (I8490,I8391,I8473);
DFFARX1 I_341 (I8490,I2683,I8077,I8066,);
nor I_342 (I8521,I8111,I8473);
DFFARX1 I_343 (I8521,I2683,I8077,I8063,);
nor I_344 (I8552,I1038232,I1038241);
DFFARX1 I_345 (I8552,I2683,I8077,I8578,);
nor I_346 (I8586,I8578,I1038226);
nand I_347 (I8603,I8586,I8193);
nand I_348 (I8057,I8603,I8292);
nand I_349 (I8054,I8586,I8340);
not I_350 (I8672,I2690);
DFFARX1 I_351 (I858255,I2683,I8672,I8698,);
nand I_352 (I8706,I8698,I858255);
not I_353 (I8723,I8706);
DFFARX1 I_354 (I8723,I2683,I8672,I8664,);
DFFARX1 I_355 (I858270,I2683,I8672,I8763,);
not I_356 (I8771,I8763);
not I_357 (I8788,I858267);
not I_358 (I8805,I858276);
nand I_359 (I8822,I8771,I8805);
nor I_360 (I8839,I8822,I858267);
DFFARX1 I_361 (I8839,I2683,I8672,I8643,);
nor I_362 (I8870,I858276,I858267);
nand I_363 (I8887,I8763,I8870);
nor I_364 (I8904,I858264,I858273);
nor I_365 (I8646,I8822,I858264);
not I_366 (I8935,I858264);
not I_367 (I8952,I858261);
nand I_368 (I8969,I8952,I858252);
nand I_369 (I8986,I8788,I8969);
not I_370 (I9003,I8986);
nor I_371 (I9020,I858261,I858273);
nor I_372 (I8655,I9003,I9020);
nor I_373 (I9051,I858258,I858261);
and I_374 (I9068,I9051,I8904);
nor I_375 (I9085,I8986,I9068);
DFFARX1 I_376 (I9085,I2683,I8672,I8661,);
nor I_377 (I9116,I8706,I9068);
DFFARX1 I_378 (I9116,I2683,I8672,I8658,);
nor I_379 (I9147,I858258,I858252);
DFFARX1 I_380 (I9147,I2683,I8672,I9173,);
nor I_381 (I9181,I9173,I858276);
nand I_382 (I9198,I9181,I8788);
nand I_383 (I8652,I9198,I8887);
nand I_384 (I8649,I9181,I8935);
not I_385 (I9267,I2690);
DFFARX1 I_386 (I444543,I2683,I9267,I9293,);
nand I_387 (I9301,I9293,I444561);
not I_388 (I9318,I9301);
DFFARX1 I_389 (I9318,I2683,I9267,I9259,);
DFFARX1 I_390 (I444555,I2683,I9267,I9358,);
not I_391 (I9366,I9358);
not I_392 (I9383,I444546);
not I_393 (I9400,I444543);
nand I_394 (I9417,I9366,I9400);
nor I_395 (I9434,I9417,I444546);
DFFARX1 I_396 (I9434,I2683,I9267,I9238,);
nor I_397 (I9465,I444543,I444546);
nand I_398 (I9482,I9358,I9465);
nor I_399 (I9499,I444552,I444540);
nor I_400 (I9241,I9417,I444552);
not I_401 (I9530,I444552);
not I_402 (I9547,I444558);
nand I_403 (I9564,I9547,I444564);
nand I_404 (I9581,I9383,I9564);
not I_405 (I9598,I9581);
nor I_406 (I9615,I444558,I444540);
nor I_407 (I9250,I9598,I9615);
nor I_408 (I9646,I444540,I444558);
and I_409 (I9663,I9646,I9499);
nor I_410 (I9680,I9581,I9663);
DFFARX1 I_411 (I9680,I2683,I9267,I9256,);
nor I_412 (I9711,I9301,I9663);
DFFARX1 I_413 (I9711,I2683,I9267,I9253,);
nor I_414 (I9742,I444540,I444549);
DFFARX1 I_415 (I9742,I2683,I9267,I9768,);
nor I_416 (I9776,I9768,I444543);
nand I_417 (I9793,I9776,I9383);
nand I_418 (I9247,I9793,I9482);
nand I_419 (I9244,I9776,I9530);
not I_420 (I9862,I2690);
DFFARX1 I_421 (I699340,I2683,I9862,I9888,);
nand I_422 (I9896,I9888,I699331);
not I_423 (I9913,I9896);
DFFARX1 I_424 (I9913,I2683,I9862,I9854,);
DFFARX1 I_425 (I699334,I2683,I9862,I9953,);
not I_426 (I9961,I9953);
not I_427 (I9978,I699346);
not I_428 (I9995,I699325);
nand I_429 (I10012,I9961,I9995);
nor I_430 (I10029,I10012,I699346);
DFFARX1 I_431 (I10029,I2683,I9862,I9833,);
nor I_432 (I10060,I699325,I699346);
nand I_433 (I10077,I9953,I10060);
nor I_434 (I10094,I699337,I699343);
nor I_435 (I9836,I10012,I699337);
not I_436 (I10125,I699337);
not I_437 (I10142,I699328);
nand I_438 (I10159,I10142,I699319);
nand I_439 (I10176,I9978,I10159);
not I_440 (I10193,I10176);
nor I_441 (I10210,I699328,I699343);
nor I_442 (I9845,I10193,I10210);
nor I_443 (I10241,I699319,I699328);
and I_444 (I10258,I10241,I10094);
nor I_445 (I10275,I10176,I10258);
DFFARX1 I_446 (I10275,I2683,I9862,I9851,);
nor I_447 (I10306,I9896,I10258);
DFFARX1 I_448 (I10306,I2683,I9862,I9848,);
nor I_449 (I10337,I699319,I699322);
DFFARX1 I_450 (I10337,I2683,I9862,I10363,);
nor I_451 (I10371,I10363,I699325);
nand I_452 (I10388,I10371,I9978);
nand I_453 (I9842,I10388,I10077);
nand I_454 (I9839,I10371,I10125);
not I_455 (I10457,I2690);
DFFARX1 I_456 (I912009,I2683,I10457,I10483,);
nand I_457 (I10491,I10483,I912009);
not I_458 (I10508,I10491);
DFFARX1 I_459 (I10508,I2683,I10457,I10449,);
DFFARX1 I_460 (I912024,I2683,I10457,I10548,);
not I_461 (I10556,I10548);
not I_462 (I10573,I912021);
not I_463 (I10590,I912030);
nand I_464 (I10607,I10556,I10590);
nor I_465 (I10624,I10607,I912021);
DFFARX1 I_466 (I10624,I2683,I10457,I10428,);
nor I_467 (I10655,I912030,I912021);
nand I_468 (I10672,I10548,I10655);
nor I_469 (I10689,I912018,I912027);
nor I_470 (I10431,I10607,I912018);
not I_471 (I10720,I912018);
not I_472 (I10737,I912015);
nand I_473 (I10754,I10737,I912006);
nand I_474 (I10771,I10573,I10754);
not I_475 (I10788,I10771);
nor I_476 (I10805,I912015,I912027);
nor I_477 (I10440,I10788,I10805);
nor I_478 (I10836,I912012,I912015);
and I_479 (I10853,I10836,I10689);
nor I_480 (I10870,I10771,I10853);
DFFARX1 I_481 (I10870,I2683,I10457,I10446,);
nor I_482 (I10901,I10491,I10853);
DFFARX1 I_483 (I10901,I2683,I10457,I10443,);
nor I_484 (I10932,I912012,I912006);
DFFARX1 I_485 (I10932,I2683,I10457,I10958,);
nor I_486 (I10966,I10958,I912030);
nand I_487 (I10983,I10966,I10573);
nand I_488 (I10437,I10983,I10672);
nand I_489 (I10434,I10966,I10720);
not I_490 (I11052,I2690);
DFFARX1 I_491 (I851319,I2683,I11052,I11078,);
nand I_492 (I11086,I11078,I851319);
not I_493 (I11103,I11086);
DFFARX1 I_494 (I11103,I2683,I11052,I11044,);
DFFARX1 I_495 (I851334,I2683,I11052,I11143,);
not I_496 (I11151,I11143);
not I_497 (I11168,I851331);
not I_498 (I11185,I851340);
nand I_499 (I11202,I11151,I11185);
nor I_500 (I11219,I11202,I851331);
DFFARX1 I_501 (I11219,I2683,I11052,I11023,);
nor I_502 (I11250,I851340,I851331);
nand I_503 (I11267,I11143,I11250);
nor I_504 (I11284,I851328,I851337);
nor I_505 (I11026,I11202,I851328);
not I_506 (I11315,I851328);
not I_507 (I11332,I851325);
nand I_508 (I11349,I11332,I851316);
nand I_509 (I11366,I11168,I11349);
not I_510 (I11383,I11366);
nor I_511 (I11400,I851325,I851337);
nor I_512 (I11035,I11383,I11400);
nor I_513 (I11431,I851322,I851325);
and I_514 (I11448,I11431,I11284);
nor I_515 (I11465,I11366,I11448);
DFFARX1 I_516 (I11465,I2683,I11052,I11041,);
nor I_517 (I11496,I11086,I11448);
DFFARX1 I_518 (I11496,I2683,I11052,I11038,);
nor I_519 (I11527,I851322,I851316);
DFFARX1 I_520 (I11527,I2683,I11052,I11553,);
nor I_521 (I11561,I11553,I851340);
nand I_522 (I11578,I11561,I11168);
nand I_523 (I11032,I11578,I11267);
nand I_524 (I11029,I11561,I11315);
not I_525 (I11650,I2690);
DFFARX1 I_526 (I93306,I2683,I11650,I11676,);
DFFARX1 I_527 (I11676,I2683,I11650,I11693,);
not I_528 (I11701,I11693);
nand I_529 (I11718,I93306,I93321);
and I_530 (I11735,I11718,I93324);
DFFARX1 I_531 (I11735,I2683,I11650,I11761,);
DFFARX1 I_532 (I11761,I2683,I11650,I11642,);
DFFARX1 I_533 (I11761,I2683,I11650,I11633,);
DFFARX1 I_534 (I93318,I2683,I11650,I11806,);
nand I_535 (I11814,I11806,I93327);
not I_536 (I11831,I11814);
nor I_537 (I11630,I11676,I11831);
DFFARX1 I_538 (I93303,I2683,I11650,I11871,);
not I_539 (I11879,I11871);
nor I_540 (I11636,I11879,I11701);
nand I_541 (I11624,I11879,I11814);
nand I_542 (I11924,I93303,I93309);
and I_543 (I11941,I11924,I93312);
DFFARX1 I_544 (I11941,I2683,I11650,I11967,);
nor I_545 (I11975,I11967,I11676);
DFFARX1 I_546 (I11975,I2683,I11650,I11618,);
not I_547 (I12006,I11967);
nor I_548 (I12023,I93315,I93309);
not I_549 (I12040,I12023);
nor I_550 (I12057,I11814,I12040);
nor I_551 (I12074,I12006,I12057);
DFFARX1 I_552 (I12074,I2683,I11650,I11639,);
nor I_553 (I12105,I11967,I12040);
nor I_554 (I11627,I11831,I12105);
nor I_555 (I11621,I11967,I12023);
not I_556 (I12177,I2690);
DFFARX1 I_557 (I1003617,I2683,I12177,I12203,);
DFFARX1 I_558 (I12203,I2683,I12177,I12220,);
not I_559 (I12228,I12220);
nand I_560 (I12245,I1003620,I1003614);
and I_561 (I12262,I12245,I1003623);
DFFARX1 I_562 (I12262,I2683,I12177,I12288,);
DFFARX1 I_563 (I12288,I2683,I12177,I12169,);
DFFARX1 I_564 (I12288,I2683,I12177,I12160,);
DFFARX1 I_565 (I1003611,I2683,I12177,I12333,);
nand I_566 (I12341,I12333,I1003626);
not I_567 (I12358,I12341);
nor I_568 (I12157,I12203,I12358);
DFFARX1 I_569 (I1003602,I2683,I12177,I12398,);
not I_570 (I12406,I12398);
nor I_571 (I12163,I12406,I12228);
nand I_572 (I12151,I12406,I12341);
nand I_573 (I12451,I1003605,I1003605);
and I_574 (I12468,I12451,I1003602);
DFFARX1 I_575 (I12468,I2683,I12177,I12494,);
nor I_576 (I12502,I12494,I12203);
DFFARX1 I_577 (I12502,I2683,I12177,I12145,);
not I_578 (I12533,I12494);
nor I_579 (I12550,I1003608,I1003605);
not I_580 (I12567,I12550);
nor I_581 (I12584,I12341,I12567);
nor I_582 (I12601,I12533,I12584);
DFFARX1 I_583 (I12601,I2683,I12177,I12166,);
nor I_584 (I12632,I12494,I12567);
nor I_585 (I12154,I12358,I12632);
nor I_586 (I12148,I12494,I12550);
not I_587 (I12704,I2690);
DFFARX1 I_588 (I619632,I2683,I12704,I12730,);
DFFARX1 I_589 (I12730,I2683,I12704,I12747,);
not I_590 (I12755,I12747);
nand I_591 (I12772,I619623,I619644);
and I_592 (I12789,I12772,I619626);
DFFARX1 I_593 (I12789,I2683,I12704,I12815,);
DFFARX1 I_594 (I12815,I2683,I12704,I12696,);
DFFARX1 I_595 (I12815,I2683,I12704,I12687,);
DFFARX1 I_596 (I619626,I2683,I12704,I12860,);
nand I_597 (I12868,I12860,I619641);
not I_598 (I12885,I12868);
nor I_599 (I12684,I12730,I12885);
DFFARX1 I_600 (I619635,I2683,I12704,I12925,);
not I_601 (I12933,I12925);
nor I_602 (I12690,I12933,I12755);
nand I_603 (I12678,I12933,I12868);
nand I_604 (I12978,I619629,I619638);
and I_605 (I12995,I12978,I619623);
DFFARX1 I_606 (I12995,I2683,I12704,I13021,);
nor I_607 (I13029,I13021,I12730);
DFFARX1 I_608 (I13029,I2683,I12704,I12672,);
not I_609 (I13060,I13021);
nor I_610 (I13077,I619629,I619638);
not I_611 (I13094,I13077);
nor I_612 (I13111,I12868,I13094);
nor I_613 (I13128,I13060,I13111);
DFFARX1 I_614 (I13128,I2683,I12704,I12693,);
nor I_615 (I13159,I13021,I13094);
nor I_616 (I12681,I12885,I13159);
nor I_617 (I12675,I13021,I13077);
not I_618 (I13231,I2690);
DFFARX1 I_619 (I752315,I2683,I13231,I13257,);
DFFARX1 I_620 (I13257,I2683,I13231,I13274,);
not I_621 (I13282,I13274);
nand I_622 (I13299,I752291,I752318);
and I_623 (I13316,I13299,I752303);
DFFARX1 I_624 (I13316,I2683,I13231,I13342,);
DFFARX1 I_625 (I13342,I2683,I13231,I13223,);
DFFARX1 I_626 (I13342,I2683,I13231,I13214,);
DFFARX1 I_627 (I752309,I2683,I13231,I13387,);
nand I_628 (I13395,I13387,I752294);
not I_629 (I13412,I13395);
nor I_630 (I13211,I13257,I13412);
DFFARX1 I_631 (I752312,I2683,I13231,I13452,);
not I_632 (I13460,I13452);
nor I_633 (I13217,I13460,I13282);
nand I_634 (I13205,I13460,I13395);
nand I_635 (I13505,I752297,I752300);
and I_636 (I13522,I13505,I752291);
DFFARX1 I_637 (I13522,I2683,I13231,I13548,);
nor I_638 (I13556,I13548,I13257);
DFFARX1 I_639 (I13556,I2683,I13231,I13199,);
not I_640 (I13587,I13548);
nor I_641 (I13604,I752306,I752300);
not I_642 (I13621,I13604);
nor I_643 (I13638,I13395,I13621);
nor I_644 (I13655,I13587,I13638);
DFFARX1 I_645 (I13655,I2683,I13231,I13220,);
nor I_646 (I13686,I13548,I13621);
nor I_647 (I13208,I13412,I13686);
nor I_648 (I13202,I13548,I13604);
not I_649 (I13758,I2690);
DFFARX1 I_650 (I541072,I2683,I13758,I13784,);
DFFARX1 I_651 (I13784,I2683,I13758,I13801,);
not I_652 (I13809,I13801);
nand I_653 (I13826,I541087,I541090);
and I_654 (I13843,I13826,I541069);
DFFARX1 I_655 (I13843,I2683,I13758,I13869,);
DFFARX1 I_656 (I13869,I2683,I13758,I13750,);
DFFARX1 I_657 (I13869,I2683,I13758,I13741,);
DFFARX1 I_658 (I541075,I2683,I13758,I13914,);
nand I_659 (I13922,I13914,I541081);
not I_660 (I13939,I13922);
nor I_661 (I13738,I13784,I13939);
DFFARX1 I_662 (I541069,I2683,I13758,I13979,);
not I_663 (I13987,I13979);
nor I_664 (I13744,I13987,I13809);
nand I_665 (I13732,I13987,I13922);
nand I_666 (I14032,I541084,I541066);
and I_667 (I14049,I14032,I541078);
DFFARX1 I_668 (I14049,I2683,I13758,I14075,);
nor I_669 (I14083,I14075,I13784);
DFFARX1 I_670 (I14083,I2683,I13758,I13726,);
not I_671 (I14114,I14075);
nor I_672 (I14131,I541066,I541066);
not I_673 (I14148,I14131);
nor I_674 (I14165,I13922,I14148);
nor I_675 (I14182,I14114,I14165);
DFFARX1 I_676 (I14182,I2683,I13758,I13747,);
nor I_677 (I14213,I14075,I14148);
nor I_678 (I13735,I13939,I14213);
nor I_679 (I13729,I14075,I14131);
not I_680 (I14285,I2690);
DFFARX1 I_681 (I676021,I2683,I14285,I14311,);
DFFARX1 I_682 (I14311,I2683,I14285,I14328,);
not I_683 (I14336,I14328);
nand I_684 (I14353,I676012,I676033);
and I_685 (I14370,I14353,I676015);
DFFARX1 I_686 (I14370,I2683,I14285,I14396,);
DFFARX1 I_687 (I14396,I2683,I14285,I14277,);
DFFARX1 I_688 (I14396,I2683,I14285,I14268,);
DFFARX1 I_689 (I676015,I2683,I14285,I14441,);
nand I_690 (I14449,I14441,I676030);
not I_691 (I14466,I14449);
nor I_692 (I14265,I14311,I14466);
DFFARX1 I_693 (I676024,I2683,I14285,I14506,);
not I_694 (I14514,I14506);
nor I_695 (I14271,I14514,I14336);
nand I_696 (I14259,I14514,I14449);
nand I_697 (I14559,I676018,I676027);
and I_698 (I14576,I14559,I676012);
DFFARX1 I_699 (I14576,I2683,I14285,I14602,);
nor I_700 (I14610,I14602,I14311);
DFFARX1 I_701 (I14610,I2683,I14285,I14253,);
not I_702 (I14641,I14602);
nor I_703 (I14658,I676018,I676027);
not I_704 (I14675,I14658);
nor I_705 (I14692,I14449,I14675);
nor I_706 (I14709,I14641,I14692);
DFFARX1 I_707 (I14709,I2683,I14285,I14274,);
nor I_708 (I14740,I14602,I14675);
nor I_709 (I14262,I14466,I14740);
nor I_710 (I14256,I14602,I14658);
not I_711 (I14812,I2690);
DFFARX1 I_712 (I191416,I2683,I14812,I14838,);
DFFARX1 I_713 (I14838,I2683,I14812,I14855,);
not I_714 (I14863,I14855);
nand I_715 (I14880,I191434,I191419);
and I_716 (I14897,I14880,I191422);
DFFARX1 I_717 (I14897,I2683,I14812,I14923,);
DFFARX1 I_718 (I14923,I2683,I14812,I14804,);
DFFARX1 I_719 (I14923,I2683,I14812,I14795,);
DFFARX1 I_720 (I191410,I2683,I14812,I14968,);
nand I_721 (I14976,I14968,I191413);
not I_722 (I14993,I14976);
nor I_723 (I14792,I14838,I14993);
DFFARX1 I_724 (I191425,I2683,I14812,I15033,);
not I_725 (I15041,I15033);
nor I_726 (I14798,I15041,I14863);
nand I_727 (I14786,I15041,I14976);
nand I_728 (I15086,I191431,I191428);
and I_729 (I15103,I15086,I191413);
DFFARX1 I_730 (I15103,I2683,I14812,I15129,);
nor I_731 (I15137,I15129,I14838);
DFFARX1 I_732 (I15137,I2683,I14812,I14780,);
not I_733 (I15168,I15129);
nor I_734 (I15185,I191410,I191428);
not I_735 (I15202,I15185);
nor I_736 (I15219,I14976,I15202);
nor I_737 (I15236,I15168,I15219);
DFFARX1 I_738 (I15236,I2683,I14812,I14801,);
nor I_739 (I15267,I15129,I15202);
nor I_740 (I14789,I14993,I15267);
nor I_741 (I14783,I15129,I15185);
not I_742 (I15339,I2690);
DFFARX1 I_743 (I456115,I2683,I15339,I15365,);
DFFARX1 I_744 (I15365,I2683,I15339,I15382,);
not I_745 (I15390,I15382);
nand I_746 (I15407,I456100,I456118);
and I_747 (I15424,I15407,I456112);
DFFARX1 I_748 (I15424,I2683,I15339,I15450,);
DFFARX1 I_749 (I15450,I2683,I15339,I15331,);
DFFARX1 I_750 (I15450,I2683,I15339,I15322,);
DFFARX1 I_751 (I456109,I2683,I15339,I15495,);
nand I_752 (I15503,I15495,I456100);
not I_753 (I15520,I15503);
nor I_754 (I15319,I15365,I15520);
DFFARX1 I_755 (I456103,I2683,I15339,I15560,);
not I_756 (I15568,I15560);
nor I_757 (I15325,I15568,I15390);
nand I_758 (I15313,I15568,I15503);
nand I_759 (I15613,I456124,I456106);
and I_760 (I15630,I15613,I456121);
DFFARX1 I_761 (I15630,I2683,I15339,I15656,);
nor I_762 (I15664,I15656,I15365);
DFFARX1 I_763 (I15664,I2683,I15339,I15307,);
not I_764 (I15695,I15656);
nor I_765 (I15712,I456103,I456106);
not I_766 (I15729,I15712);
nor I_767 (I15746,I15503,I15729);
nor I_768 (I15763,I15695,I15746);
DFFARX1 I_769 (I15763,I2683,I15339,I15328,);
nor I_770 (I15794,I15656,I15729);
nor I_771 (I15316,I15520,I15794);
nor I_772 (I15310,I15656,I15712);
not I_773 (I15866,I2690);
DFFARX1 I_774 (I356786,I2683,I15866,I15892,);
DFFARX1 I_775 (I15892,I2683,I15866,I15909,);
not I_776 (I15917,I15909);
nand I_777 (I15934,I356786,I356789);
and I_778 (I15951,I15934,I356810);
DFFARX1 I_779 (I15951,I2683,I15866,I15977,);
DFFARX1 I_780 (I15977,I2683,I15866,I15858,);
DFFARX1 I_781 (I15977,I2683,I15866,I15849,);
DFFARX1 I_782 (I356798,I2683,I15866,I16022,);
nand I_783 (I16030,I16022,I356801);
not I_784 (I16047,I16030);
nor I_785 (I15846,I15892,I16047);
DFFARX1 I_786 (I356807,I2683,I15866,I16087,);
not I_787 (I16095,I16087);
nor I_788 (I15852,I16095,I15917);
nand I_789 (I15840,I16095,I16030);
nand I_790 (I16140,I356804,I356792);
and I_791 (I16157,I16140,I356795);
DFFARX1 I_792 (I16157,I2683,I15866,I16183,);
nor I_793 (I16191,I16183,I15892);
DFFARX1 I_794 (I16191,I2683,I15866,I15834,);
not I_795 (I16222,I16183);
nor I_796 (I16239,I356813,I356792);
not I_797 (I16256,I16239);
nor I_798 (I16273,I16030,I16256);
nor I_799 (I16290,I16222,I16273);
DFFARX1 I_800 (I16290,I2683,I15866,I15855,);
nor I_801 (I16321,I16183,I16256);
nor I_802 (I15843,I16047,I16321);
nor I_803 (I15837,I16183,I16239);
not I_804 (I16393,I2690);
DFFARX1 I_805 (I236963,I2683,I16393,I16419,);
DFFARX1 I_806 (I16419,I2683,I16393,I16436,);
not I_807 (I16444,I16436);
nand I_808 (I16461,I236960,I236954);
and I_809 (I16478,I16461,I236948);
DFFARX1 I_810 (I16478,I2683,I16393,I16504,);
DFFARX1 I_811 (I16504,I2683,I16393,I16385,);
DFFARX1 I_812 (I16504,I2683,I16393,I16376,);
DFFARX1 I_813 (I236936,I2683,I16393,I16549,);
nand I_814 (I16557,I16549,I236945);
not I_815 (I16574,I16557);
nor I_816 (I16373,I16419,I16574);
DFFARX1 I_817 (I236942,I2683,I16393,I16614,);
not I_818 (I16622,I16614);
nor I_819 (I16379,I16622,I16444);
nand I_820 (I16367,I16622,I16557);
nand I_821 (I16667,I236939,I236957);
and I_822 (I16684,I16667,I236936);
DFFARX1 I_823 (I16684,I2683,I16393,I16710,);
nor I_824 (I16718,I16710,I16419);
DFFARX1 I_825 (I16718,I2683,I16393,I16361,);
not I_826 (I16749,I16710);
nor I_827 (I16766,I236951,I236957);
not I_828 (I16783,I16766);
nor I_829 (I16800,I16557,I16783);
nor I_830 (I16817,I16749,I16800);
DFFARX1 I_831 (I16817,I2683,I16393,I16382,);
nor I_832 (I16848,I16710,I16783);
nor I_833 (I16370,I16574,I16848);
nor I_834 (I16364,I16710,I16766);
not I_835 (I16920,I2690);
DFFARX1 I_836 (I258043,I2683,I16920,I16946,);
DFFARX1 I_837 (I16946,I2683,I16920,I16963,);
not I_838 (I16971,I16963);
nand I_839 (I16988,I258040,I258034);
and I_840 (I17005,I16988,I258028);
DFFARX1 I_841 (I17005,I2683,I16920,I17031,);
DFFARX1 I_842 (I17031,I2683,I16920,I16912,);
DFFARX1 I_843 (I17031,I2683,I16920,I16903,);
DFFARX1 I_844 (I258016,I2683,I16920,I17076,);
nand I_845 (I17084,I17076,I258025);
not I_846 (I17101,I17084);
nor I_847 (I16900,I16946,I17101);
DFFARX1 I_848 (I258022,I2683,I16920,I17141,);
not I_849 (I17149,I17141);
nor I_850 (I16906,I17149,I16971);
nand I_851 (I16894,I17149,I17084);
nand I_852 (I17194,I258019,I258037);
and I_853 (I17211,I17194,I258016);
DFFARX1 I_854 (I17211,I2683,I16920,I17237,);
nor I_855 (I17245,I17237,I16946);
DFFARX1 I_856 (I17245,I2683,I16920,I16888,);
not I_857 (I17276,I17237);
nor I_858 (I17293,I258031,I258037);
not I_859 (I17310,I17293);
nor I_860 (I17327,I17084,I17310);
nor I_861 (I17344,I17276,I17327);
DFFARX1 I_862 (I17344,I2683,I16920,I16909,);
nor I_863 (I17375,I17237,I17310);
nor I_864 (I16897,I17101,I17375);
nor I_865 (I16891,I17237,I17293);
not I_866 (I17447,I2690);
DFFARX1 I_867 (I1452,I2683,I17447,I17473,);
DFFARX1 I_868 (I17473,I2683,I17447,I17490,);
not I_869 (I17498,I17490);
nand I_870 (I17515,I2156,I1396);
and I_871 (I17532,I17515,I2116);
DFFARX1 I_872 (I17532,I2683,I17447,I17558,);
DFFARX1 I_873 (I17558,I2683,I17447,I17439,);
DFFARX1 I_874 (I17558,I2683,I17447,I17430,);
DFFARX1 I_875 (I1940,I2683,I17447,I17603,);
nand I_876 (I17611,I17603,I2132);
not I_877 (I17628,I17611);
nor I_878 (I17427,I17473,I17628);
DFFARX1 I_879 (I1692,I2683,I17447,I17668,);
not I_880 (I17676,I17668);
nor I_881 (I17433,I17676,I17498);
nand I_882 (I17421,I17676,I17611);
nand I_883 (I17721,I1676,I2628);
and I_884 (I17738,I17721,I2204);
DFFARX1 I_885 (I17738,I2683,I17447,I17764,);
nor I_886 (I17772,I17764,I17473);
DFFARX1 I_887 (I17772,I2683,I17447,I17415,);
not I_888 (I17803,I17764);
nor I_889 (I17820,I2236,I2628);
not I_890 (I17837,I17820);
nor I_891 (I17854,I17611,I17837);
nor I_892 (I17871,I17803,I17854);
DFFARX1 I_893 (I17871,I2683,I17447,I17436,);
nor I_894 (I17902,I17764,I17837);
nor I_895 (I17424,I17628,I17902);
nor I_896 (I17418,I17764,I17820);
not I_897 (I17974,I2690);
DFFARX1 I_898 (I159286,I2683,I17974,I18000,);
DFFARX1 I_899 (I18000,I2683,I17974,I18017,);
not I_900 (I18025,I18017);
nand I_901 (I18042,I159304,I159289);
and I_902 (I18059,I18042,I159292);
DFFARX1 I_903 (I18059,I2683,I17974,I18085,);
DFFARX1 I_904 (I18085,I2683,I17974,I17966,);
DFFARX1 I_905 (I18085,I2683,I17974,I17957,);
DFFARX1 I_906 (I159280,I2683,I17974,I18130,);
nand I_907 (I18138,I18130,I159283);
not I_908 (I18155,I18138);
nor I_909 (I17954,I18000,I18155);
DFFARX1 I_910 (I159295,I2683,I17974,I18195,);
not I_911 (I18203,I18195);
nor I_912 (I17960,I18203,I18025);
nand I_913 (I17948,I18203,I18138);
nand I_914 (I18248,I159301,I159298);
and I_915 (I18265,I18248,I159283);
DFFARX1 I_916 (I18265,I2683,I17974,I18291,);
nor I_917 (I18299,I18291,I18000);
DFFARX1 I_918 (I18299,I2683,I17974,I17942,);
not I_919 (I18330,I18291);
nor I_920 (I18347,I159280,I159298);
not I_921 (I18364,I18347);
nor I_922 (I18381,I18138,I18364);
nor I_923 (I18398,I18330,I18381);
DFFARX1 I_924 (I18398,I2683,I17974,I17963,);
nor I_925 (I18429,I18291,I18364);
nor I_926 (I17951,I18155,I18429);
nor I_927 (I17945,I18291,I18347);
not I_928 (I18501,I2690);
DFFARX1 I_929 (I1045354,I2683,I18501,I18527,);
DFFARX1 I_930 (I18527,I2683,I18501,I18544,);
not I_931 (I18552,I18544);
nand I_932 (I18569,I1045357,I1045363);
and I_933 (I18586,I18569,I1045372);
DFFARX1 I_934 (I18586,I2683,I18501,I18612,);
DFFARX1 I_935 (I18612,I2683,I18501,I18493,);
DFFARX1 I_936 (I18612,I2683,I18501,I18484,);
DFFARX1 I_937 (I1045375,I2683,I18501,I18657,);
nand I_938 (I18665,I18657,I1045366);
not I_939 (I18682,I18665);
nor I_940 (I18481,I18527,I18682);
DFFARX1 I_941 (I1045354,I2683,I18501,I18722,);
not I_942 (I18730,I18722);
nor I_943 (I18487,I18730,I18552);
nand I_944 (I18475,I18730,I18665);
nand I_945 (I18775,I1045381,I1045360);
and I_946 (I18792,I18775,I1045369);
DFFARX1 I_947 (I18792,I2683,I18501,I18818,);
nor I_948 (I18826,I18818,I18527);
DFFARX1 I_949 (I18826,I2683,I18501,I18469,);
not I_950 (I18857,I18818);
nor I_951 (I18874,I1045378,I1045360);
not I_952 (I18891,I18874);
nor I_953 (I18908,I18665,I18891);
nor I_954 (I18925,I18857,I18908);
DFFARX1 I_955 (I18925,I2683,I18501,I18490,);
nor I_956 (I18956,I18818,I18891);
nor I_957 (I18478,I18682,I18956);
nor I_958 (I18472,I18818,I18874);
not I_959 (I19028,I2690);
DFFARX1 I_960 (I487327,I2683,I19028,I19054,);
DFFARX1 I_961 (I19054,I2683,I19028,I19071,);
not I_962 (I19079,I19071);
nand I_963 (I19096,I487312,I487330);
and I_964 (I19113,I19096,I487324);
DFFARX1 I_965 (I19113,I2683,I19028,I19139,);
DFFARX1 I_966 (I19139,I2683,I19028,I19020,);
DFFARX1 I_967 (I19139,I2683,I19028,I19011,);
DFFARX1 I_968 (I487321,I2683,I19028,I19184,);
nand I_969 (I19192,I19184,I487312);
not I_970 (I19209,I19192);
nor I_971 (I19008,I19054,I19209);
DFFARX1 I_972 (I487315,I2683,I19028,I19249,);
not I_973 (I19257,I19249);
nor I_974 (I19014,I19257,I19079);
nand I_975 (I19002,I19257,I19192);
nand I_976 (I19302,I487336,I487318);
and I_977 (I19319,I19302,I487333);
DFFARX1 I_978 (I19319,I2683,I19028,I19345,);
nor I_979 (I19353,I19345,I19054);
DFFARX1 I_980 (I19353,I2683,I19028,I18996,);
not I_981 (I19384,I19345);
nor I_982 (I19401,I487315,I487318);
not I_983 (I19418,I19401);
nor I_984 (I19435,I19192,I19418);
nor I_985 (I19452,I19384,I19435);
DFFARX1 I_986 (I19452,I2683,I19028,I19017,);
nor I_987 (I19483,I19345,I19418);
nor I_988 (I19005,I19209,I19483);
nor I_989 (I18999,I19345,I19401);
not I_990 (I19555,I2690);
DFFARX1 I_991 (I606386,I2683,I19555,I19581,);
DFFARX1 I_992 (I19581,I2683,I19555,I19598,);
not I_993 (I19606,I19598);
nand I_994 (I19623,I606401,I606404);
and I_995 (I19640,I19623,I606383);
DFFARX1 I_996 (I19640,I2683,I19555,I19666,);
DFFARX1 I_997 (I19666,I2683,I19555,I19547,);
DFFARX1 I_998 (I19666,I2683,I19555,I19538,);
DFFARX1 I_999 (I606389,I2683,I19555,I19711,);
nand I_1000 (I19719,I19711,I606395);
not I_1001 (I19736,I19719);
nor I_1002 (I19535,I19581,I19736);
DFFARX1 I_1003 (I606383,I2683,I19555,I19776,);
not I_1004 (I19784,I19776);
nor I_1005 (I19541,I19784,I19606);
nand I_1006 (I19529,I19784,I19719);
nand I_1007 (I19829,I606398,I606380);
and I_1008 (I19846,I19829,I606392);
DFFARX1 I_1009 (I19846,I2683,I19555,I19872,);
nor I_1010 (I19880,I19872,I19581);
DFFARX1 I_1011 (I19880,I2683,I19555,I19523,);
not I_1012 (I19911,I19872);
nor I_1013 (I19928,I606380,I606380);
not I_1014 (I19945,I19928);
nor I_1015 (I19962,I19719,I19945);
nor I_1016 (I19979,I19911,I19962);
DFFARX1 I_1017 (I19979,I2683,I19555,I19544,);
nor I_1018 (I20010,I19872,I19945);
nor I_1019 (I19532,I19736,I20010);
nor I_1020 (I19526,I19872,I19928);
not I_1021 (I20082,I2690);
DFFARX1 I_1022 (I542228,I2683,I20082,I20108,);
DFFARX1 I_1023 (I20108,I2683,I20082,I20125,);
not I_1024 (I20133,I20125);
nand I_1025 (I20150,I542243,I542246);
and I_1026 (I20167,I20150,I542225);
DFFARX1 I_1027 (I20167,I2683,I20082,I20193,);
DFFARX1 I_1028 (I20193,I2683,I20082,I20074,);
DFFARX1 I_1029 (I20193,I2683,I20082,I20065,);
DFFARX1 I_1030 (I542231,I2683,I20082,I20238,);
nand I_1031 (I20246,I20238,I542237);
not I_1032 (I20263,I20246);
nor I_1033 (I20062,I20108,I20263);
DFFARX1 I_1034 (I542225,I2683,I20082,I20303,);
not I_1035 (I20311,I20303);
nor I_1036 (I20068,I20311,I20133);
nand I_1037 (I20056,I20311,I20246);
nand I_1038 (I20356,I542240,I542222);
and I_1039 (I20373,I20356,I542234);
DFFARX1 I_1040 (I20373,I2683,I20082,I20399,);
nor I_1041 (I20407,I20399,I20108);
DFFARX1 I_1042 (I20407,I2683,I20082,I20050,);
not I_1043 (I20438,I20399);
nor I_1044 (I20455,I542222,I542222);
not I_1045 (I20472,I20455);
nor I_1046 (I20489,I20246,I20472);
nor I_1047 (I20506,I20438,I20489);
DFFARX1 I_1048 (I20506,I2683,I20082,I20071,);
nor I_1049 (I20537,I20399,I20472);
nor I_1050 (I20059,I20263,I20537);
nor I_1051 (I20053,I20399,I20455);
not I_1052 (I20609,I2690);
DFFARX1 I_1053 (I729705,I2683,I20609,I20635,);
DFFARX1 I_1054 (I20635,I2683,I20609,I20652,);
not I_1055 (I20660,I20652);
nand I_1056 (I20677,I729681,I729708);
and I_1057 (I20694,I20677,I729693);
DFFARX1 I_1058 (I20694,I2683,I20609,I20720,);
DFFARX1 I_1059 (I20720,I2683,I20609,I20601,);
DFFARX1 I_1060 (I20720,I2683,I20609,I20592,);
DFFARX1 I_1061 (I729699,I2683,I20609,I20765,);
nand I_1062 (I20773,I20765,I729684);
not I_1063 (I20790,I20773);
nor I_1064 (I20589,I20635,I20790);
DFFARX1 I_1065 (I729702,I2683,I20609,I20830,);
not I_1066 (I20838,I20830);
nor I_1067 (I20595,I20838,I20660);
nand I_1068 (I20583,I20838,I20773);
nand I_1069 (I20883,I729687,I729690);
and I_1070 (I20900,I20883,I729681);
DFFARX1 I_1071 (I20900,I2683,I20609,I20926,);
nor I_1072 (I20934,I20926,I20635);
DFFARX1 I_1073 (I20934,I2683,I20609,I20577,);
not I_1074 (I20965,I20926);
nor I_1075 (I20982,I729696,I729690);
not I_1076 (I20999,I20982);
nor I_1077 (I21016,I20773,I20999);
nor I_1078 (I21033,I20965,I21016);
DFFARX1 I_1079 (I21033,I2683,I20609,I20598,);
nor I_1080 (I21064,I20926,I20999);
nor I_1081 (I20586,I20790,I21064);
nor I_1082 (I20580,I20926,I20982);
not I_1083 (I21136,I2690);
DFFARX1 I_1084 (I520842,I2683,I21136,I21162,);
DFFARX1 I_1085 (I21162,I2683,I21136,I21179,);
not I_1086 (I21187,I21179);
nand I_1087 (I21204,I520857,I520860);
and I_1088 (I21221,I21204,I520839);
DFFARX1 I_1089 (I21221,I2683,I21136,I21247,);
DFFARX1 I_1090 (I21247,I2683,I21136,I21128,);
DFFARX1 I_1091 (I21247,I2683,I21136,I21119,);
DFFARX1 I_1092 (I520845,I2683,I21136,I21292,);
nand I_1093 (I21300,I21292,I520851);
not I_1094 (I21317,I21300);
nor I_1095 (I21116,I21162,I21317);
DFFARX1 I_1096 (I520839,I2683,I21136,I21357,);
not I_1097 (I21365,I21357);
nor I_1098 (I21122,I21365,I21187);
nand I_1099 (I21110,I21365,I21300);
nand I_1100 (I21410,I520854,I520836);
and I_1101 (I21427,I21410,I520848);
DFFARX1 I_1102 (I21427,I2683,I21136,I21453,);
nor I_1103 (I21461,I21453,I21162);
DFFARX1 I_1104 (I21461,I2683,I21136,I21104,);
not I_1105 (I21492,I21453);
nor I_1106 (I21509,I520836,I520836);
not I_1107 (I21526,I21509);
nor I_1108 (I21543,I21300,I21526);
nor I_1109 (I21560,I21492,I21543);
DFFARX1 I_1110 (I21560,I2683,I21136,I21125,);
nor I_1111 (I21591,I21453,I21526);
nor I_1112 (I21113,I21317,I21591);
nor I_1113 (I21107,I21453,I21509);
not I_1114 (I21663,I2690);
DFFARX1 I_1115 (I730997,I2683,I21663,I21689,);
DFFARX1 I_1116 (I21689,I2683,I21663,I21706,);
not I_1117 (I21714,I21706);
nand I_1118 (I21731,I730973,I731000);
and I_1119 (I21748,I21731,I730985);
DFFARX1 I_1120 (I21748,I2683,I21663,I21774,);
DFFARX1 I_1121 (I21774,I2683,I21663,I21655,);
DFFARX1 I_1122 (I21774,I2683,I21663,I21646,);
DFFARX1 I_1123 (I730991,I2683,I21663,I21819,);
nand I_1124 (I21827,I21819,I730976);
not I_1125 (I21844,I21827);
nor I_1126 (I21643,I21689,I21844);
DFFARX1 I_1127 (I730994,I2683,I21663,I21884,);
not I_1128 (I21892,I21884);
nor I_1129 (I21649,I21892,I21714);
nand I_1130 (I21637,I21892,I21827);
nand I_1131 (I21937,I730979,I730982);
and I_1132 (I21954,I21937,I730973);
DFFARX1 I_1133 (I21954,I2683,I21663,I21980,);
nor I_1134 (I21988,I21980,I21689);
DFFARX1 I_1135 (I21988,I2683,I21663,I21631,);
not I_1136 (I22019,I21980);
nor I_1137 (I22036,I730988,I730982);
not I_1138 (I22053,I22036);
nor I_1139 (I22070,I21827,I22053);
nor I_1140 (I22087,I22019,I22070);
DFFARX1 I_1141 (I22087,I2683,I21663,I21652,);
nor I_1142 (I22118,I21980,I22053);
nor I_1143 (I21640,I21844,I22118);
nor I_1144 (I21634,I21980,I22036);
not I_1145 (I22190,I2690);
DFFARX1 I_1146 (I284920,I2683,I22190,I22216,);
DFFARX1 I_1147 (I22216,I2683,I22190,I22233,);
not I_1148 (I22241,I22233);
nand I_1149 (I22258,I284917,I284911);
and I_1150 (I22275,I22258,I284905);
DFFARX1 I_1151 (I22275,I2683,I22190,I22301,);
DFFARX1 I_1152 (I22301,I2683,I22190,I22182,);
DFFARX1 I_1153 (I22301,I2683,I22190,I22173,);
DFFARX1 I_1154 (I284893,I2683,I22190,I22346,);
nand I_1155 (I22354,I22346,I284902);
not I_1156 (I22371,I22354);
nor I_1157 (I22170,I22216,I22371);
DFFARX1 I_1158 (I284899,I2683,I22190,I22411,);
not I_1159 (I22419,I22411);
nor I_1160 (I22176,I22419,I22241);
nand I_1161 (I22164,I22419,I22354);
nand I_1162 (I22464,I284896,I284914);
and I_1163 (I22481,I22464,I284893);
DFFARX1 I_1164 (I22481,I2683,I22190,I22507,);
nor I_1165 (I22515,I22507,I22216);
DFFARX1 I_1166 (I22515,I2683,I22190,I22158,);
not I_1167 (I22546,I22507);
nor I_1168 (I22563,I284908,I284914);
not I_1169 (I22580,I22563);
nor I_1170 (I22597,I22354,I22580);
nor I_1171 (I22614,I22546,I22597);
DFFARX1 I_1172 (I22614,I2683,I22190,I22179,);
nor I_1173 (I22645,I22507,I22580);
nor I_1174 (I22167,I22371,I22645);
nor I_1175 (I22161,I22507,I22563);
not I_1176 (I22717,I2690);
DFFARX1 I_1177 (I969534,I2683,I22717,I22743,);
DFFARX1 I_1178 (I22743,I2683,I22717,I22760,);
not I_1179 (I22768,I22760);
nand I_1180 (I22785,I969552,I969546);
and I_1181 (I22802,I22785,I969555);
DFFARX1 I_1182 (I22802,I2683,I22717,I22828,);
DFFARX1 I_1183 (I22828,I2683,I22717,I22709,);
DFFARX1 I_1184 (I22828,I2683,I22717,I22700,);
DFFARX1 I_1185 (I969540,I2683,I22717,I22873,);
nand I_1186 (I22881,I22873,I969549);
not I_1187 (I22898,I22881);
nor I_1188 (I22697,I22743,I22898);
DFFARX1 I_1189 (I969537,I2683,I22717,I22938,);
not I_1190 (I22946,I22938);
nor I_1191 (I22703,I22946,I22768);
nand I_1192 (I22691,I22946,I22881);
nand I_1193 (I22991,I969558,I969543);
and I_1194 (I23008,I22991,I969537);
DFFARX1 I_1195 (I23008,I2683,I22717,I23034,);
nor I_1196 (I23042,I23034,I22743);
DFFARX1 I_1197 (I23042,I2683,I22717,I22685,);
not I_1198 (I23073,I23034);
nor I_1199 (I23090,I969534,I969543);
not I_1200 (I23107,I23090);
nor I_1201 (I23124,I22881,I23107);
nor I_1202 (I23141,I23073,I23124);
DFFARX1 I_1203 (I23141,I2683,I22717,I22706,);
nor I_1204 (I23172,I23034,I23107);
nor I_1205 (I22694,I22898,I23172);
nor I_1206 (I22688,I23034,I23090);
not I_1207 (I23244,I2690);
DFFARX1 I_1208 (I216937,I2683,I23244,I23270,);
DFFARX1 I_1209 (I23270,I2683,I23244,I23287,);
not I_1210 (I23295,I23287);
nand I_1211 (I23312,I216934,I216928);
and I_1212 (I23329,I23312,I216922);
DFFARX1 I_1213 (I23329,I2683,I23244,I23355,);
DFFARX1 I_1214 (I23355,I2683,I23244,I23236,);
DFFARX1 I_1215 (I23355,I2683,I23244,I23227,);
DFFARX1 I_1216 (I216910,I2683,I23244,I23400,);
nand I_1217 (I23408,I23400,I216919);
not I_1218 (I23425,I23408);
nor I_1219 (I23224,I23270,I23425);
DFFARX1 I_1220 (I216916,I2683,I23244,I23465,);
not I_1221 (I23473,I23465);
nor I_1222 (I23230,I23473,I23295);
nand I_1223 (I23218,I23473,I23408);
nand I_1224 (I23518,I216913,I216931);
and I_1225 (I23535,I23518,I216910);
DFFARX1 I_1226 (I23535,I2683,I23244,I23561,);
nor I_1227 (I23569,I23561,I23270);
DFFARX1 I_1228 (I23569,I2683,I23244,I23212,);
not I_1229 (I23600,I23561);
nor I_1230 (I23617,I216925,I216931);
not I_1231 (I23634,I23617);
nor I_1232 (I23651,I23408,I23634);
nor I_1233 (I23668,I23600,I23651);
DFFARX1 I_1234 (I23668,I2683,I23244,I23233,);
nor I_1235 (I23699,I23561,I23634);
nor I_1236 (I23221,I23425,I23699);
nor I_1237 (I23215,I23561,I23617);
not I_1238 (I23771,I2690);
DFFARX1 I_1239 (I228531,I2683,I23771,I23797,);
DFFARX1 I_1240 (I23797,I2683,I23771,I23814,);
not I_1241 (I23822,I23814);
nand I_1242 (I23839,I228528,I228522);
and I_1243 (I23856,I23839,I228516);
DFFARX1 I_1244 (I23856,I2683,I23771,I23882,);
DFFARX1 I_1245 (I23882,I2683,I23771,I23763,);
DFFARX1 I_1246 (I23882,I2683,I23771,I23754,);
DFFARX1 I_1247 (I228504,I2683,I23771,I23927,);
nand I_1248 (I23935,I23927,I228513);
not I_1249 (I23952,I23935);
nor I_1250 (I23751,I23797,I23952);
DFFARX1 I_1251 (I228510,I2683,I23771,I23992,);
not I_1252 (I24000,I23992);
nor I_1253 (I23757,I24000,I23822);
nand I_1254 (I23745,I24000,I23935);
nand I_1255 (I24045,I228507,I228525);
and I_1256 (I24062,I24045,I228504);
DFFARX1 I_1257 (I24062,I2683,I23771,I24088,);
nor I_1258 (I24096,I24088,I23797);
DFFARX1 I_1259 (I24096,I2683,I23771,I23739,);
not I_1260 (I24127,I24088);
nor I_1261 (I24144,I228519,I228525);
not I_1262 (I24161,I24144);
nor I_1263 (I24178,I23935,I24161);
nor I_1264 (I24195,I24127,I24178);
DFFARX1 I_1265 (I24195,I2683,I23771,I23760,);
nor I_1266 (I24226,I24088,I24161);
nor I_1267 (I23748,I23952,I24226);
nor I_1268 (I23742,I24088,I24144);
not I_1269 (I24298,I2690);
DFFARX1 I_1270 (I1020379,I2683,I24298,I24324,);
DFFARX1 I_1271 (I24324,I2683,I24298,I24341,);
not I_1272 (I24349,I24341);
nand I_1273 (I24366,I1020382,I1020376);
and I_1274 (I24383,I24366,I1020385);
DFFARX1 I_1275 (I24383,I2683,I24298,I24409,);
DFFARX1 I_1276 (I24409,I2683,I24298,I24290,);
DFFARX1 I_1277 (I24409,I2683,I24298,I24281,);
DFFARX1 I_1278 (I1020373,I2683,I24298,I24454,);
nand I_1279 (I24462,I24454,I1020388);
not I_1280 (I24479,I24462);
nor I_1281 (I24278,I24324,I24479);
DFFARX1 I_1282 (I1020364,I2683,I24298,I24519,);
not I_1283 (I24527,I24519);
nor I_1284 (I24284,I24527,I24349);
nand I_1285 (I24272,I24527,I24462);
nand I_1286 (I24572,I1020367,I1020367);
and I_1287 (I24589,I24572,I1020364);
DFFARX1 I_1288 (I24589,I2683,I24298,I24615,);
nor I_1289 (I24623,I24615,I24324);
DFFARX1 I_1290 (I24623,I2683,I24298,I24266,);
not I_1291 (I24654,I24615);
nor I_1292 (I24671,I1020370,I1020367);
not I_1293 (I24688,I24671);
nor I_1294 (I24705,I24462,I24688);
nor I_1295 (I24722,I24654,I24705);
DFFARX1 I_1296 (I24722,I2683,I24298,I24287,);
nor I_1297 (I24753,I24615,I24688);
nor I_1298 (I24275,I24479,I24753);
nor I_1299 (I24269,I24615,I24671);
not I_1300 (I24825,I2690);
DFFARX1 I_1301 (I744563,I2683,I24825,I24851,);
DFFARX1 I_1302 (I24851,I2683,I24825,I24868,);
not I_1303 (I24876,I24868);
nand I_1304 (I24893,I744539,I744566);
and I_1305 (I24910,I24893,I744551);
DFFARX1 I_1306 (I24910,I2683,I24825,I24936,);
DFFARX1 I_1307 (I24936,I2683,I24825,I24817,);
DFFARX1 I_1308 (I24936,I2683,I24825,I24808,);
DFFARX1 I_1309 (I744557,I2683,I24825,I24981,);
nand I_1310 (I24989,I24981,I744542);
not I_1311 (I25006,I24989);
nor I_1312 (I24805,I24851,I25006);
DFFARX1 I_1313 (I744560,I2683,I24825,I25046,);
not I_1314 (I25054,I25046);
nor I_1315 (I24811,I25054,I24876);
nand I_1316 (I24799,I25054,I24989);
nand I_1317 (I25099,I744545,I744548);
and I_1318 (I25116,I25099,I744539);
DFFARX1 I_1319 (I25116,I2683,I24825,I25142,);
nor I_1320 (I25150,I25142,I24851);
DFFARX1 I_1321 (I25150,I2683,I24825,I24793,);
not I_1322 (I25181,I25142);
nor I_1323 (I25198,I744554,I744548);
not I_1324 (I25215,I25198);
nor I_1325 (I25232,I24989,I25215);
nor I_1326 (I25249,I25181,I25232);
DFFARX1 I_1327 (I25249,I2683,I24825,I24814,);
nor I_1328 (I25280,I25142,I25215);
nor I_1329 (I24802,I25006,I25280);
nor I_1330 (I24796,I25142,I25198);
not I_1331 (I25352,I2690);
DFFARX1 I_1332 (I79077,I2683,I25352,I25378,);
DFFARX1 I_1333 (I25378,I2683,I25352,I25395,);
not I_1334 (I25403,I25395);
nand I_1335 (I25420,I79077,I79092);
and I_1336 (I25437,I25420,I79095);
DFFARX1 I_1337 (I25437,I2683,I25352,I25463,);
DFFARX1 I_1338 (I25463,I2683,I25352,I25344,);
DFFARX1 I_1339 (I25463,I2683,I25352,I25335,);
DFFARX1 I_1340 (I79089,I2683,I25352,I25508,);
nand I_1341 (I25516,I25508,I79098);
not I_1342 (I25533,I25516);
nor I_1343 (I25332,I25378,I25533);
DFFARX1 I_1344 (I79074,I2683,I25352,I25573,);
not I_1345 (I25581,I25573);
nor I_1346 (I25338,I25581,I25403);
nand I_1347 (I25326,I25581,I25516);
nand I_1348 (I25626,I79074,I79080);
and I_1349 (I25643,I25626,I79083);
DFFARX1 I_1350 (I25643,I2683,I25352,I25669,);
nor I_1351 (I25677,I25669,I25378);
DFFARX1 I_1352 (I25677,I2683,I25352,I25320,);
not I_1353 (I25708,I25669);
nor I_1354 (I25725,I79086,I79080);
not I_1355 (I25742,I25725);
nor I_1356 (I25759,I25516,I25742);
nor I_1357 (I25776,I25708,I25759);
DFFARX1 I_1358 (I25776,I2683,I25352,I25341,);
nor I_1359 (I25807,I25669,I25742);
nor I_1360 (I25329,I25533,I25807);
nor I_1361 (I25323,I25669,I25725);
not I_1362 (I25879,I2690);
DFFARX1 I_1363 (I808006,I2683,I25879,I25905,);
DFFARX1 I_1364 (I25905,I2683,I25879,I25922,);
not I_1365 (I25930,I25922);
nand I_1366 (I25947,I808000,I808021);
and I_1367 (I25964,I25947,I808006);
DFFARX1 I_1368 (I25964,I2683,I25879,I25990,);
DFFARX1 I_1369 (I25990,I2683,I25879,I25871,);
DFFARX1 I_1370 (I25990,I2683,I25879,I25862,);
DFFARX1 I_1371 (I808003,I2683,I25879,I26035,);
nand I_1372 (I26043,I26035,I808012);
not I_1373 (I26060,I26043);
nor I_1374 (I25859,I25905,I26060);
DFFARX1 I_1375 (I808000,I2683,I25879,I26100,);
not I_1376 (I26108,I26100);
nor I_1377 (I25865,I26108,I25930);
nand I_1378 (I25853,I26108,I26043);
nand I_1379 (I26153,I808003,I808018);
and I_1380 (I26170,I26153,I808009);
DFFARX1 I_1381 (I26170,I2683,I25879,I26196,);
nor I_1382 (I26204,I26196,I25905);
DFFARX1 I_1383 (I26204,I2683,I25879,I25847,);
not I_1384 (I26235,I26196);
nor I_1385 (I26252,I808015,I808018);
not I_1386 (I26269,I26252);
nor I_1387 (I26286,I26043,I26269);
nor I_1388 (I26303,I26235,I26286);
DFFARX1 I_1389 (I26303,I2683,I25879,I25868,);
nor I_1390 (I26334,I26196,I26269);
nor I_1391 (I25856,I26060,I26334);
nor I_1392 (I25850,I26196,I26252);
not I_1393 (I26406,I2690);
DFFARX1 I_1394 (I471721,I2683,I26406,I26432,);
DFFARX1 I_1395 (I26432,I2683,I26406,I26449,);
not I_1396 (I26457,I26449);
nand I_1397 (I26474,I471706,I471724);
and I_1398 (I26491,I26474,I471718);
DFFARX1 I_1399 (I26491,I2683,I26406,I26517,);
DFFARX1 I_1400 (I26517,I2683,I26406,I26398,);
DFFARX1 I_1401 (I26517,I2683,I26406,I26389,);
DFFARX1 I_1402 (I471715,I2683,I26406,I26562,);
nand I_1403 (I26570,I26562,I471706);
not I_1404 (I26587,I26570);
nor I_1405 (I26386,I26432,I26587);
DFFARX1 I_1406 (I471709,I2683,I26406,I26627,);
not I_1407 (I26635,I26627);
nor I_1408 (I26392,I26635,I26457);
nand I_1409 (I26380,I26635,I26570);
nand I_1410 (I26680,I471730,I471712);
and I_1411 (I26697,I26680,I471727);
DFFARX1 I_1412 (I26697,I2683,I26406,I26723,);
nor I_1413 (I26731,I26723,I26432);
DFFARX1 I_1414 (I26731,I2683,I26406,I26374,);
not I_1415 (I26762,I26723);
nor I_1416 (I26779,I471709,I471712);
not I_1417 (I26796,I26779);
nor I_1418 (I26813,I26570,I26796);
nor I_1419 (I26830,I26762,I26813);
DFFARX1 I_1420 (I26830,I2683,I26406,I26395,);
nor I_1421 (I26861,I26723,I26796);
nor I_1422 (I26383,I26587,I26861);
nor I_1423 (I26377,I26723,I26779);
not I_1424 (I26933,I2690);
DFFARX1 I_1425 (I114670,I2683,I26933,I26959,);
DFFARX1 I_1426 (I26959,I2683,I26933,I26976,);
not I_1427 (I26984,I26976);
nand I_1428 (I27001,I114673,I114655);
and I_1429 (I27018,I27001,I114661);
DFFARX1 I_1430 (I27018,I2683,I26933,I27044,);
DFFARX1 I_1431 (I27044,I2683,I26933,I26925,);
DFFARX1 I_1432 (I27044,I2683,I26933,I26916,);
DFFARX1 I_1433 (I114664,I2683,I26933,I27089,);
nand I_1434 (I27097,I27089,I114655);
not I_1435 (I27114,I27097);
nor I_1436 (I26913,I26959,I27114);
DFFARX1 I_1437 (I114676,I2683,I26933,I27154,);
not I_1438 (I27162,I27154);
nor I_1439 (I26919,I27162,I26984);
nand I_1440 (I26907,I27162,I27097);
nand I_1441 (I27207,I114679,I114667);
and I_1442 (I27224,I27207,I114658);
DFFARX1 I_1443 (I27224,I2683,I26933,I27250,);
nor I_1444 (I27258,I27250,I26959);
DFFARX1 I_1445 (I27258,I2683,I26933,I26901,);
not I_1446 (I27289,I27250);
nor I_1447 (I27306,I114682,I114667);
not I_1448 (I27323,I27306);
nor I_1449 (I27340,I27097,I27323);
nor I_1450 (I27357,I27289,I27340);
DFFARX1 I_1451 (I27357,I2683,I26933,I26922,);
nor I_1452 (I27388,I27250,I27323);
nor I_1453 (I26910,I27114,I27388);
nor I_1454 (I26904,I27250,I27306);
not I_1455 (I27460,I2690);
DFFARX1 I_1456 (I69064,I2683,I27460,I27486,);
DFFARX1 I_1457 (I27486,I2683,I27460,I27503,);
not I_1458 (I27511,I27503);
nand I_1459 (I27528,I69064,I69079);
and I_1460 (I27545,I27528,I69082);
DFFARX1 I_1461 (I27545,I2683,I27460,I27571,);
DFFARX1 I_1462 (I27571,I2683,I27460,I27452,);
DFFARX1 I_1463 (I27571,I2683,I27460,I27443,);
DFFARX1 I_1464 (I69076,I2683,I27460,I27616,);
nand I_1465 (I27624,I27616,I69085);
not I_1466 (I27641,I27624);
nor I_1467 (I27440,I27486,I27641);
DFFARX1 I_1468 (I69061,I2683,I27460,I27681,);
not I_1469 (I27689,I27681);
nor I_1470 (I27446,I27689,I27511);
nand I_1471 (I27434,I27689,I27624);
nand I_1472 (I27734,I69061,I69067);
and I_1473 (I27751,I27734,I69070);
DFFARX1 I_1474 (I27751,I2683,I27460,I27777,);
nor I_1475 (I27785,I27777,I27486);
DFFARX1 I_1476 (I27785,I2683,I27460,I27428,);
not I_1477 (I27816,I27777);
nor I_1478 (I27833,I69073,I69067);
not I_1479 (I27850,I27833);
nor I_1480 (I27867,I27624,I27850);
nor I_1481 (I27884,I27816,I27867);
DFFARX1 I_1482 (I27884,I2683,I27460,I27449,);
nor I_1483 (I27915,I27777,I27850);
nor I_1484 (I27437,I27641,I27915);
nor I_1485 (I27431,I27777,I27833);
not I_1486 (I27987,I2690);
DFFARX1 I_1487 (I500034,I2683,I27987,I28013,);
DFFARX1 I_1488 (I28013,I2683,I27987,I28030,);
not I_1489 (I28038,I28030);
nand I_1490 (I28055,I500049,I500052);
and I_1491 (I28072,I28055,I500031);
DFFARX1 I_1492 (I28072,I2683,I27987,I28098,);
DFFARX1 I_1493 (I28098,I2683,I27987,I27979,);
DFFARX1 I_1494 (I28098,I2683,I27987,I27970,);
DFFARX1 I_1495 (I500037,I2683,I27987,I28143,);
nand I_1496 (I28151,I28143,I500043);
not I_1497 (I28168,I28151);
nor I_1498 (I27967,I28013,I28168);
DFFARX1 I_1499 (I500031,I2683,I27987,I28208,);
not I_1500 (I28216,I28208);
nor I_1501 (I27973,I28216,I28038);
nand I_1502 (I27961,I28216,I28151);
nand I_1503 (I28261,I500046,I500028);
and I_1504 (I28278,I28261,I500040);
DFFARX1 I_1505 (I28278,I2683,I27987,I28304,);
nor I_1506 (I28312,I28304,I28013);
DFFARX1 I_1507 (I28312,I2683,I27987,I27955,);
not I_1508 (I28343,I28304);
nor I_1509 (I28360,I500028,I500028);
not I_1510 (I28377,I28360);
nor I_1511 (I28394,I28151,I28377);
nor I_1512 (I28411,I28343,I28394);
DFFARX1 I_1513 (I28411,I2683,I27987,I27976,);
nor I_1514 (I28442,I28304,I28377);
nor I_1515 (I27964,I28168,I28442);
nor I_1516 (I27958,I28304,I28360);
not I_1517 (I28514,I2690);
DFFARX1 I_1518 (I598872,I2683,I28514,I28540,);
DFFARX1 I_1519 (I28540,I2683,I28514,I28557,);
not I_1520 (I28565,I28557);
nand I_1521 (I28582,I598887,I598890);
and I_1522 (I28599,I28582,I598869);
DFFARX1 I_1523 (I28599,I2683,I28514,I28625,);
DFFARX1 I_1524 (I28625,I2683,I28514,I28506,);
DFFARX1 I_1525 (I28625,I2683,I28514,I28497,);
DFFARX1 I_1526 (I598875,I2683,I28514,I28670,);
nand I_1527 (I28678,I28670,I598881);
not I_1528 (I28695,I28678);
nor I_1529 (I28494,I28540,I28695);
DFFARX1 I_1530 (I598869,I2683,I28514,I28735,);
not I_1531 (I28743,I28735);
nor I_1532 (I28500,I28743,I28565);
nand I_1533 (I28488,I28743,I28678);
nand I_1534 (I28788,I598884,I598866);
and I_1535 (I28805,I28788,I598878);
DFFARX1 I_1536 (I28805,I2683,I28514,I28831,);
nor I_1537 (I28839,I28831,I28540);
DFFARX1 I_1538 (I28839,I2683,I28514,I28482,);
not I_1539 (I28870,I28831);
nor I_1540 (I28887,I598866,I598866);
not I_1541 (I28904,I28887);
nor I_1542 (I28921,I28678,I28904);
nor I_1543 (I28938,I28870,I28921);
DFFARX1 I_1544 (I28938,I2683,I28514,I28503,);
nor I_1545 (I28969,I28831,I28904);
nor I_1546 (I28491,I28695,I28969);
nor I_1547 (I28485,I28831,I28887);
not I_1548 (I29041,I2690);
DFFARX1 I_1549 (I1037024,I2683,I29041,I29067,);
DFFARX1 I_1550 (I29067,I2683,I29041,I29084,);
not I_1551 (I29092,I29084);
nand I_1552 (I29109,I1037027,I1037033);
and I_1553 (I29126,I29109,I1037042);
DFFARX1 I_1554 (I29126,I2683,I29041,I29152,);
DFFARX1 I_1555 (I29152,I2683,I29041,I29033,);
DFFARX1 I_1556 (I29152,I2683,I29041,I29024,);
DFFARX1 I_1557 (I1037045,I2683,I29041,I29197,);
nand I_1558 (I29205,I29197,I1037036);
not I_1559 (I29222,I29205);
nor I_1560 (I29021,I29067,I29222);
DFFARX1 I_1561 (I1037024,I2683,I29041,I29262,);
not I_1562 (I29270,I29262);
nor I_1563 (I29027,I29270,I29092);
nand I_1564 (I29015,I29270,I29205);
nand I_1565 (I29315,I1037051,I1037030);
and I_1566 (I29332,I29315,I1037039);
DFFARX1 I_1567 (I29332,I2683,I29041,I29358,);
nor I_1568 (I29366,I29358,I29067);
DFFARX1 I_1569 (I29366,I2683,I29041,I29009,);
not I_1570 (I29397,I29358);
nor I_1571 (I29414,I1037048,I1037030);
not I_1572 (I29431,I29414);
nor I_1573 (I29448,I29205,I29431);
nor I_1574 (I29465,I29397,I29448);
DFFARX1 I_1575 (I29465,I2683,I29041,I29030,);
nor I_1576 (I29496,I29358,I29431);
nor I_1577 (I29018,I29222,I29496);
nor I_1578 (I29012,I29358,I29414);
not I_1579 (I29568,I2690);
DFFARX1 I_1580 (I1063799,I2683,I29568,I29594,);
DFFARX1 I_1581 (I29594,I2683,I29568,I29611,);
not I_1582 (I29619,I29611);
nand I_1583 (I29636,I1063802,I1063808);
and I_1584 (I29653,I29636,I1063817);
DFFARX1 I_1585 (I29653,I2683,I29568,I29679,);
DFFARX1 I_1586 (I29679,I2683,I29568,I29560,);
DFFARX1 I_1587 (I29679,I2683,I29568,I29551,);
DFFARX1 I_1588 (I1063820,I2683,I29568,I29724,);
nand I_1589 (I29732,I29724,I1063811);
not I_1590 (I29749,I29732);
nor I_1591 (I29548,I29594,I29749);
DFFARX1 I_1592 (I1063799,I2683,I29568,I29789,);
not I_1593 (I29797,I29789);
nor I_1594 (I29554,I29797,I29619);
nand I_1595 (I29542,I29797,I29732);
nand I_1596 (I29842,I1063826,I1063805);
and I_1597 (I29859,I29842,I1063814);
DFFARX1 I_1598 (I29859,I2683,I29568,I29885,);
nor I_1599 (I29893,I29885,I29594);
DFFARX1 I_1600 (I29893,I2683,I29568,I29536,);
not I_1601 (I29924,I29885);
nor I_1602 (I29941,I1063823,I1063805);
not I_1603 (I29958,I29941);
nor I_1604 (I29975,I29732,I29958);
nor I_1605 (I29992,I29924,I29975);
DFFARX1 I_1606 (I29992,I2683,I29568,I29557,);
nor I_1607 (I30023,I29885,I29958);
nor I_1608 (I29545,I29749,I30023);
nor I_1609 (I29539,I29885,I29941);
not I_1610 (I30095,I2690);
DFFARX1 I_1611 (I335570,I2683,I30095,I30121,);
DFFARX1 I_1612 (I30121,I2683,I30095,I30138,);
not I_1613 (I30146,I30138);
nand I_1614 (I30163,I335570,I335573);
and I_1615 (I30180,I30163,I335594);
DFFARX1 I_1616 (I30180,I2683,I30095,I30206,);
DFFARX1 I_1617 (I30206,I2683,I30095,I30087,);
DFFARX1 I_1618 (I30206,I2683,I30095,I30078,);
DFFARX1 I_1619 (I335582,I2683,I30095,I30251,);
nand I_1620 (I30259,I30251,I335585);
not I_1621 (I30276,I30259);
nor I_1622 (I30075,I30121,I30276);
DFFARX1 I_1623 (I335591,I2683,I30095,I30316,);
not I_1624 (I30324,I30316);
nor I_1625 (I30081,I30324,I30146);
nand I_1626 (I30069,I30324,I30259);
nand I_1627 (I30369,I335588,I335576);
and I_1628 (I30386,I30369,I335579);
DFFARX1 I_1629 (I30386,I2683,I30095,I30412,);
nor I_1630 (I30420,I30412,I30121);
DFFARX1 I_1631 (I30420,I2683,I30095,I30063,);
not I_1632 (I30451,I30412);
nor I_1633 (I30468,I335597,I335576);
not I_1634 (I30485,I30468);
nor I_1635 (I30502,I30259,I30485);
nor I_1636 (I30519,I30451,I30502);
DFFARX1 I_1637 (I30519,I2683,I30095,I30084,);
nor I_1638 (I30550,I30412,I30485);
nor I_1639 (I30072,I30276,I30550);
nor I_1640 (I30066,I30412,I30468);
not I_1641 (I30622,I2690);
DFFARX1 I_1642 (I115860,I2683,I30622,I30648,);
DFFARX1 I_1643 (I30648,I2683,I30622,I30665,);
not I_1644 (I30673,I30665);
nand I_1645 (I30690,I115863,I115845);
and I_1646 (I30707,I30690,I115851);
DFFARX1 I_1647 (I30707,I2683,I30622,I30733,);
DFFARX1 I_1648 (I30733,I2683,I30622,I30614,);
DFFARX1 I_1649 (I30733,I2683,I30622,I30605,);
DFFARX1 I_1650 (I115854,I2683,I30622,I30778,);
nand I_1651 (I30786,I30778,I115845);
not I_1652 (I30803,I30786);
nor I_1653 (I30602,I30648,I30803);
DFFARX1 I_1654 (I115866,I2683,I30622,I30843,);
not I_1655 (I30851,I30843);
nor I_1656 (I30608,I30851,I30673);
nand I_1657 (I30596,I30851,I30786);
nand I_1658 (I30896,I115869,I115857);
and I_1659 (I30913,I30896,I115848);
DFFARX1 I_1660 (I30913,I2683,I30622,I30939,);
nor I_1661 (I30947,I30939,I30648);
DFFARX1 I_1662 (I30947,I2683,I30622,I30590,);
not I_1663 (I30978,I30939);
nor I_1664 (I30995,I115872,I115857);
not I_1665 (I31012,I30995);
nor I_1666 (I31029,I30786,I31012);
nor I_1667 (I31046,I30978,I31029);
DFFARX1 I_1668 (I31046,I2683,I30622,I30611,);
nor I_1669 (I31077,I30939,I31012);
nor I_1670 (I30599,I30803,I31077);
nor I_1671 (I30593,I30939,I30995);
not I_1672 (I31149,I2690);
DFFARX1 I_1673 (I960830,I2683,I31149,I31175,);
DFFARX1 I_1674 (I31175,I2683,I31149,I31192,);
not I_1675 (I31200,I31192);
nand I_1676 (I31217,I960848,I960842);
and I_1677 (I31234,I31217,I960851);
DFFARX1 I_1678 (I31234,I2683,I31149,I31260,);
DFFARX1 I_1679 (I31260,I2683,I31149,I31141,);
DFFARX1 I_1680 (I31260,I2683,I31149,I31132,);
DFFARX1 I_1681 (I960836,I2683,I31149,I31305,);
nand I_1682 (I31313,I31305,I960845);
not I_1683 (I31330,I31313);
nor I_1684 (I31129,I31175,I31330);
DFFARX1 I_1685 (I960833,I2683,I31149,I31370,);
not I_1686 (I31378,I31370);
nor I_1687 (I31135,I31378,I31200);
nand I_1688 (I31123,I31378,I31313);
nand I_1689 (I31423,I960854,I960839);
and I_1690 (I31440,I31423,I960833);
DFFARX1 I_1691 (I31440,I2683,I31149,I31466,);
nor I_1692 (I31474,I31466,I31175);
DFFARX1 I_1693 (I31474,I2683,I31149,I31117,);
not I_1694 (I31505,I31466);
nor I_1695 (I31522,I960830,I960839);
not I_1696 (I31539,I31522);
nor I_1697 (I31556,I31313,I31539);
nor I_1698 (I31573,I31505,I31556);
DFFARX1 I_1699 (I31573,I2683,I31149,I31138,);
nor I_1700 (I31604,I31466,I31539);
nor I_1701 (I31126,I31330,I31604);
nor I_1702 (I31120,I31466,I31522);
not I_1703 (I31676,I2690);
DFFARX1 I_1704 (I537026,I2683,I31676,I31702,);
DFFARX1 I_1705 (I31702,I2683,I31676,I31719,);
not I_1706 (I31727,I31719);
nand I_1707 (I31744,I537041,I537044);
and I_1708 (I31761,I31744,I537023);
DFFARX1 I_1709 (I31761,I2683,I31676,I31787,);
DFFARX1 I_1710 (I31787,I2683,I31676,I31668,);
DFFARX1 I_1711 (I31787,I2683,I31676,I31659,);
DFFARX1 I_1712 (I537029,I2683,I31676,I31832,);
nand I_1713 (I31840,I31832,I537035);
not I_1714 (I31857,I31840);
nor I_1715 (I31656,I31702,I31857);
DFFARX1 I_1716 (I537023,I2683,I31676,I31897,);
not I_1717 (I31905,I31897);
nor I_1718 (I31662,I31905,I31727);
nand I_1719 (I31650,I31905,I31840);
nand I_1720 (I31950,I537038,I537020);
and I_1721 (I31967,I31950,I537032);
DFFARX1 I_1722 (I31967,I2683,I31676,I31993,);
nor I_1723 (I32001,I31993,I31702);
DFFARX1 I_1724 (I32001,I2683,I31676,I31644,);
not I_1725 (I32032,I31993);
nor I_1726 (I32049,I537020,I537020);
not I_1727 (I32066,I32049);
nor I_1728 (I32083,I31840,I32066);
nor I_1729 (I32100,I32032,I32083);
DFFARX1 I_1730 (I32100,I2683,I31676,I31665,);
nor I_1731 (I32131,I31993,I32066);
nor I_1732 (I31653,I31857,I32131);
nor I_1733 (I31647,I31993,I32049);
not I_1734 (I32203,I2690);
DFFARX1 I_1735 (I990901,I2683,I32203,I32229,);
DFFARX1 I_1736 (I32229,I2683,I32203,I32246,);
not I_1737 (I32254,I32246);
nand I_1738 (I32271,I990904,I990898);
and I_1739 (I32288,I32271,I990907);
DFFARX1 I_1740 (I32288,I2683,I32203,I32314,);
DFFARX1 I_1741 (I32314,I2683,I32203,I32195,);
DFFARX1 I_1742 (I32314,I2683,I32203,I32186,);
DFFARX1 I_1743 (I990895,I2683,I32203,I32359,);
nand I_1744 (I32367,I32359,I990910);
not I_1745 (I32384,I32367);
nor I_1746 (I32183,I32229,I32384);
DFFARX1 I_1747 (I990886,I2683,I32203,I32424,);
not I_1748 (I32432,I32424);
nor I_1749 (I32189,I32432,I32254);
nand I_1750 (I32177,I32432,I32367);
nand I_1751 (I32477,I990889,I990889);
and I_1752 (I32494,I32477,I990886);
DFFARX1 I_1753 (I32494,I2683,I32203,I32520,);
nor I_1754 (I32528,I32520,I32229);
DFFARX1 I_1755 (I32528,I2683,I32203,I32171,);
not I_1756 (I32559,I32520);
nor I_1757 (I32576,I990892,I990889);
not I_1758 (I32593,I32576);
nor I_1759 (I32610,I32367,I32593);
nor I_1760 (I32627,I32559,I32610);
DFFARX1 I_1761 (I32627,I2683,I32203,I32192,);
nor I_1762 (I32658,I32520,I32593);
nor I_1763 (I32180,I32384,I32658);
nor I_1764 (I32174,I32520,I32576);
not I_1765 (I32730,I2690);
DFFARX1 I_1766 (I489061,I2683,I32730,I32756,);
DFFARX1 I_1767 (I32756,I2683,I32730,I32773,);
not I_1768 (I32781,I32773);
nand I_1769 (I32798,I489046,I489064);
and I_1770 (I32815,I32798,I489058);
DFFARX1 I_1771 (I32815,I2683,I32730,I32841,);
DFFARX1 I_1772 (I32841,I2683,I32730,I32722,);
DFFARX1 I_1773 (I32841,I2683,I32730,I32713,);
DFFARX1 I_1774 (I489055,I2683,I32730,I32886,);
nand I_1775 (I32894,I32886,I489046);
not I_1776 (I32911,I32894);
nor I_1777 (I32710,I32756,I32911);
DFFARX1 I_1778 (I489049,I2683,I32730,I32951,);
not I_1779 (I32959,I32951);
nor I_1780 (I32716,I32959,I32781);
nand I_1781 (I32704,I32959,I32894);
nand I_1782 (I33004,I489070,I489052);
and I_1783 (I33021,I33004,I489067);
DFFARX1 I_1784 (I33021,I2683,I32730,I33047,);
nor I_1785 (I33055,I33047,I32756);
DFFARX1 I_1786 (I33055,I2683,I32730,I32698,);
not I_1787 (I33086,I33047);
nor I_1788 (I33103,I489049,I489052);
not I_1789 (I33120,I33103);
nor I_1790 (I33137,I32894,I33120);
nor I_1791 (I33154,I33086,I33137);
DFFARX1 I_1792 (I33154,I2683,I32730,I32719,);
nor I_1793 (I33185,I33047,I33120);
nor I_1794 (I32707,I32911,I33185);
nor I_1795 (I32701,I33047,I33103);
not I_1796 (I33257,I2690);
DFFARX1 I_1797 (I307581,I2683,I33257,I33283,);
DFFARX1 I_1798 (I33283,I2683,I33257,I33300,);
not I_1799 (I33308,I33300);
nand I_1800 (I33325,I307578,I307572);
and I_1801 (I33342,I33325,I307566);
DFFARX1 I_1802 (I33342,I2683,I33257,I33368,);
DFFARX1 I_1803 (I33368,I2683,I33257,I33249,);
DFFARX1 I_1804 (I33368,I2683,I33257,I33240,);
DFFARX1 I_1805 (I307554,I2683,I33257,I33413,);
nand I_1806 (I33421,I33413,I307563);
not I_1807 (I33438,I33421);
nor I_1808 (I33237,I33283,I33438);
DFFARX1 I_1809 (I307560,I2683,I33257,I33478,);
not I_1810 (I33486,I33478);
nor I_1811 (I33243,I33486,I33308);
nand I_1812 (I33231,I33486,I33421);
nand I_1813 (I33531,I307557,I307575);
and I_1814 (I33548,I33531,I307554);
DFFARX1 I_1815 (I33548,I2683,I33257,I33574,);
nor I_1816 (I33582,I33574,I33283);
DFFARX1 I_1817 (I33582,I2683,I33257,I33225,);
not I_1818 (I33613,I33574);
nor I_1819 (I33630,I307569,I307575);
not I_1820 (I33647,I33630);
nor I_1821 (I33664,I33421,I33647);
nor I_1822 (I33681,I33613,I33664);
DFFARX1 I_1823 (I33681,I2683,I33257,I33246,);
nor I_1824 (I33712,I33574,I33647);
nor I_1825 (I33234,I33438,I33712);
nor I_1826 (I33228,I33574,I33630);
not I_1827 (I33784,I2690);
DFFARX1 I_1828 (I561880,I2683,I33784,I33810,);
DFFARX1 I_1829 (I33810,I2683,I33784,I33827,);
not I_1830 (I33835,I33827);
nand I_1831 (I33852,I561895,I561898);
and I_1832 (I33869,I33852,I561877);
DFFARX1 I_1833 (I33869,I2683,I33784,I33895,);
DFFARX1 I_1834 (I33895,I2683,I33784,I33776,);
DFFARX1 I_1835 (I33895,I2683,I33784,I33767,);
DFFARX1 I_1836 (I561883,I2683,I33784,I33940,);
nand I_1837 (I33948,I33940,I561889);
not I_1838 (I33965,I33948);
nor I_1839 (I33764,I33810,I33965);
DFFARX1 I_1840 (I561877,I2683,I33784,I34005,);
not I_1841 (I34013,I34005);
nor I_1842 (I33770,I34013,I33835);
nand I_1843 (I33758,I34013,I33948);
nand I_1844 (I34058,I561892,I561874);
and I_1845 (I34075,I34058,I561886);
DFFARX1 I_1846 (I34075,I2683,I33784,I34101,);
nor I_1847 (I34109,I34101,I33810);
DFFARX1 I_1848 (I34109,I2683,I33784,I33752,);
not I_1849 (I34140,I34101);
nor I_1850 (I34157,I561874,I561874);
not I_1851 (I34174,I34157);
nor I_1852 (I34191,I33948,I34174);
nor I_1853 (I34208,I34140,I34191);
DFFARX1 I_1854 (I34208,I2683,I33784,I33773,);
nor I_1855 (I34239,I34101,I34174);
nor I_1856 (I33761,I33965,I34239);
nor I_1857 (I33755,I34101,I34157);
not I_1858 (I34311,I2690);
DFFARX1 I_1859 (I951334,I2683,I34311,I34337,);
DFFARX1 I_1860 (I34337,I2683,I34311,I34354,);
not I_1861 (I34362,I34354);
nand I_1862 (I34379,I951322,I951313);
and I_1863 (I34396,I34379,I951310);
DFFARX1 I_1864 (I34396,I2683,I34311,I34422,);
DFFARX1 I_1865 (I34422,I2683,I34311,I34303,);
DFFARX1 I_1866 (I34422,I2683,I34311,I34294,);
DFFARX1 I_1867 (I951316,I2683,I34311,I34467,);
nand I_1868 (I34475,I34467,I951328);
not I_1869 (I34492,I34475);
nor I_1870 (I34291,I34337,I34492);
DFFARX1 I_1871 (I951325,I2683,I34311,I34532,);
not I_1872 (I34540,I34532);
nor I_1873 (I34297,I34540,I34362);
nand I_1874 (I34285,I34540,I34475);
nand I_1875 (I34585,I951319,I951313);
and I_1876 (I34602,I34585,I951331);
DFFARX1 I_1877 (I34602,I2683,I34311,I34628,);
nor I_1878 (I34636,I34628,I34337);
DFFARX1 I_1879 (I34636,I2683,I34311,I34279,);
not I_1880 (I34667,I34628);
nor I_1881 (I34684,I951310,I951313);
not I_1882 (I34701,I34684);
nor I_1883 (I34718,I34475,I34701);
nor I_1884 (I34735,I34667,I34718);
DFFARX1 I_1885 (I34735,I2683,I34311,I34300,);
nor I_1886 (I34766,I34628,I34701);
nor I_1887 (I34288,I34492,I34766);
nor I_1888 (I34282,I34628,I34684);
not I_1889 (I34838,I2690);
DFFARX1 I_1890 (I649144,I2683,I34838,I34864,);
DFFARX1 I_1891 (I34864,I2683,I34838,I34881,);
not I_1892 (I34889,I34881);
nand I_1893 (I34906,I649135,I649156);
and I_1894 (I34923,I34906,I649138);
DFFARX1 I_1895 (I34923,I2683,I34838,I34949,);
DFFARX1 I_1896 (I34949,I2683,I34838,I34830,);
DFFARX1 I_1897 (I34949,I2683,I34838,I34821,);
DFFARX1 I_1898 (I649138,I2683,I34838,I34994,);
nand I_1899 (I35002,I34994,I649153);
not I_1900 (I35019,I35002);
nor I_1901 (I34818,I34864,I35019);
DFFARX1 I_1902 (I649147,I2683,I34838,I35059,);
not I_1903 (I35067,I35059);
nor I_1904 (I34824,I35067,I34889);
nand I_1905 (I34812,I35067,I35002);
nand I_1906 (I35112,I649141,I649150);
and I_1907 (I35129,I35112,I649135);
DFFARX1 I_1908 (I35129,I2683,I34838,I35155,);
nor I_1909 (I35163,I35155,I34864);
DFFARX1 I_1910 (I35163,I2683,I34838,I34806,);
not I_1911 (I35194,I35155);
nor I_1912 (I35211,I649141,I649150);
not I_1913 (I35228,I35211);
nor I_1914 (I35245,I35002,I35228);
nor I_1915 (I35262,I35194,I35245);
DFFARX1 I_1916 (I35262,I2683,I34838,I34827,);
nor I_1917 (I35293,I35155,I35228);
nor I_1918 (I34815,I35019,I35293);
nor I_1919 (I34809,I35155,I35211);
not I_1920 (I35365,I2690);
DFFARX1 I_1921 (I521420,I2683,I35365,I35391,);
DFFARX1 I_1922 (I35391,I2683,I35365,I35408,);
not I_1923 (I35416,I35408);
nand I_1924 (I35433,I521435,I521438);
and I_1925 (I35450,I35433,I521417);
DFFARX1 I_1926 (I35450,I2683,I35365,I35476,);
DFFARX1 I_1927 (I35476,I2683,I35365,I35357,);
DFFARX1 I_1928 (I35476,I2683,I35365,I35348,);
DFFARX1 I_1929 (I521423,I2683,I35365,I35521,);
nand I_1930 (I35529,I35521,I521429);
not I_1931 (I35546,I35529);
nor I_1932 (I35345,I35391,I35546);
DFFARX1 I_1933 (I521417,I2683,I35365,I35586,);
not I_1934 (I35594,I35586);
nor I_1935 (I35351,I35594,I35416);
nand I_1936 (I35339,I35594,I35529);
nand I_1937 (I35639,I521432,I521414);
and I_1938 (I35656,I35639,I521426);
DFFARX1 I_1939 (I35656,I2683,I35365,I35682,);
nor I_1940 (I35690,I35682,I35391);
DFFARX1 I_1941 (I35690,I2683,I35365,I35333,);
not I_1942 (I35721,I35682);
nor I_1943 (I35738,I521414,I521414);
not I_1944 (I35755,I35738);
nor I_1945 (I35772,I35529,I35755);
nor I_1946 (I35789,I35721,I35772);
DFFARX1 I_1947 (I35789,I2683,I35365,I35354,);
nor I_1948 (I35820,I35682,I35755);
nor I_1949 (I35342,I35546,I35820);
nor I_1950 (I35336,I35682,I35738);
not I_1951 (I35892,I2690);
DFFARX1 I_1952 (I342098,I2683,I35892,I35918,);
DFFARX1 I_1953 (I35918,I2683,I35892,I35935,);
not I_1954 (I35943,I35935);
nand I_1955 (I35960,I342098,I342101);
and I_1956 (I35977,I35960,I342122);
DFFARX1 I_1957 (I35977,I2683,I35892,I36003,);
DFFARX1 I_1958 (I36003,I2683,I35892,I35884,);
DFFARX1 I_1959 (I36003,I2683,I35892,I35875,);
DFFARX1 I_1960 (I342110,I2683,I35892,I36048,);
nand I_1961 (I36056,I36048,I342113);
not I_1962 (I36073,I36056);
nor I_1963 (I35872,I35918,I36073);
DFFARX1 I_1964 (I342119,I2683,I35892,I36113,);
not I_1965 (I36121,I36113);
nor I_1966 (I35878,I36121,I35943);
nand I_1967 (I35866,I36121,I36056);
nand I_1968 (I36166,I342116,I342104);
and I_1969 (I36183,I36166,I342107);
DFFARX1 I_1970 (I36183,I2683,I35892,I36209,);
nor I_1971 (I36217,I36209,I35918);
DFFARX1 I_1972 (I36217,I2683,I35892,I35860,);
not I_1973 (I36248,I36209);
nor I_1974 (I36265,I342125,I342104);
not I_1975 (I36282,I36265);
nor I_1976 (I36299,I36056,I36282);
nor I_1977 (I36316,I36248,I36299);
DFFARX1 I_1978 (I36316,I2683,I35892,I35881,);
nor I_1979 (I36347,I36209,I36282);
nor I_1980 (I35869,I36073,I36347);
nor I_1981 (I35863,I36209,I36265);
not I_1982 (I36419,I2690);
DFFARX1 I_1983 (I293879,I2683,I36419,I36445,);
DFFARX1 I_1984 (I36445,I2683,I36419,I36462,);
not I_1985 (I36470,I36462);
nand I_1986 (I36487,I293876,I293870);
and I_1987 (I36504,I36487,I293864);
DFFARX1 I_1988 (I36504,I2683,I36419,I36530,);
DFFARX1 I_1989 (I36530,I2683,I36419,I36411,);
DFFARX1 I_1990 (I36530,I2683,I36419,I36402,);
DFFARX1 I_1991 (I293852,I2683,I36419,I36575,);
nand I_1992 (I36583,I36575,I293861);
not I_1993 (I36600,I36583);
nor I_1994 (I36399,I36445,I36600);
DFFARX1 I_1995 (I293858,I2683,I36419,I36640,);
not I_1996 (I36648,I36640);
nor I_1997 (I36405,I36648,I36470);
nand I_1998 (I36393,I36648,I36583);
nand I_1999 (I36693,I293855,I293873);
and I_2000 (I36710,I36693,I293852);
DFFARX1 I_2001 (I36710,I2683,I36419,I36736,);
nor I_2002 (I36744,I36736,I36445);
DFFARX1 I_2003 (I36744,I2683,I36419,I36387,);
not I_2004 (I36775,I36736);
nor I_2005 (I36792,I293867,I293873);
not I_2006 (I36809,I36792);
nor I_2007 (I36826,I36583,I36809);
nor I_2008 (I36843,I36775,I36826);
DFFARX1 I_2009 (I36843,I2683,I36419,I36408,);
nor I_2010 (I36874,I36736,I36809);
nor I_2011 (I36396,I36600,I36874);
nor I_2012 (I36390,I36736,I36792);
not I_2013 (I36946,I2690);
DFFARX1 I_2014 (I914342,I2683,I36946,I36972,);
DFFARX1 I_2015 (I36972,I2683,I36946,I36989,);
not I_2016 (I36997,I36989);
nand I_2017 (I37014,I914330,I914321);
and I_2018 (I37031,I37014,I914318);
DFFARX1 I_2019 (I37031,I2683,I36946,I37057,);
DFFARX1 I_2020 (I37057,I2683,I36946,I36938,);
DFFARX1 I_2021 (I37057,I2683,I36946,I36929,);
DFFARX1 I_2022 (I914324,I2683,I36946,I37102,);
nand I_2023 (I37110,I37102,I914336);
not I_2024 (I37127,I37110);
nor I_2025 (I36926,I36972,I37127);
DFFARX1 I_2026 (I914333,I2683,I36946,I37167,);
not I_2027 (I37175,I37167);
nor I_2028 (I36932,I37175,I36997);
nand I_2029 (I36920,I37175,I37110);
nand I_2030 (I37220,I914327,I914321);
and I_2031 (I37237,I37220,I914339);
DFFARX1 I_2032 (I37237,I2683,I36946,I37263,);
nor I_2033 (I37271,I37263,I36972);
DFFARX1 I_2034 (I37271,I2683,I36946,I36914,);
not I_2035 (I37302,I37263);
nor I_2036 (I37319,I914318,I914321);
not I_2037 (I37336,I37319);
nor I_2038 (I37353,I37110,I37336);
nor I_2039 (I37370,I37302,I37353);
DFFARX1 I_2040 (I37370,I2683,I36946,I36935,);
nor I_2041 (I37401,I37263,I37336);
nor I_2042 (I36923,I37127,I37401);
nor I_2043 (I36917,I37263,I37319);
not I_2044 (I37473,I2690);
DFFARX1 I_2045 (I935728,I2683,I37473,I37499,);
DFFARX1 I_2046 (I37499,I2683,I37473,I37516,);
not I_2047 (I37524,I37516);
nand I_2048 (I37541,I935716,I935707);
and I_2049 (I37558,I37541,I935704);
DFFARX1 I_2050 (I37558,I2683,I37473,I37584,);
DFFARX1 I_2051 (I37584,I2683,I37473,I37465,);
DFFARX1 I_2052 (I37584,I2683,I37473,I37456,);
DFFARX1 I_2053 (I935710,I2683,I37473,I37629,);
nand I_2054 (I37637,I37629,I935722);
not I_2055 (I37654,I37637);
nor I_2056 (I37453,I37499,I37654);
DFFARX1 I_2057 (I935719,I2683,I37473,I37694,);
not I_2058 (I37702,I37694);
nor I_2059 (I37459,I37702,I37524);
nand I_2060 (I37447,I37702,I37637);
nand I_2061 (I37747,I935713,I935707);
and I_2062 (I37764,I37747,I935725);
DFFARX1 I_2063 (I37764,I2683,I37473,I37790,);
nor I_2064 (I37798,I37790,I37499);
DFFARX1 I_2065 (I37798,I2683,I37473,I37441,);
not I_2066 (I37829,I37790);
nor I_2067 (I37846,I935704,I935707);
not I_2068 (I37863,I37846);
nor I_2069 (I37880,I37637,I37863);
nor I_2070 (I37897,I37829,I37880);
DFFARX1 I_2071 (I37897,I2683,I37473,I37462,);
nor I_2072 (I37928,I37790,I37863);
nor I_2073 (I37450,I37654,I37928);
nor I_2074 (I37444,I37790,I37846);
not I_2075 (I38000,I2690);
DFFARX1 I_2076 (I117050,I2683,I38000,I38026,);
DFFARX1 I_2077 (I38026,I2683,I38000,I38043,);
not I_2078 (I38051,I38043);
nand I_2079 (I38068,I117053,I117035);
and I_2080 (I38085,I38068,I117041);
DFFARX1 I_2081 (I38085,I2683,I38000,I38111,);
DFFARX1 I_2082 (I38111,I2683,I38000,I37992,);
DFFARX1 I_2083 (I38111,I2683,I38000,I37983,);
DFFARX1 I_2084 (I117044,I2683,I38000,I38156,);
nand I_2085 (I38164,I38156,I117035);
not I_2086 (I38181,I38164);
nor I_2087 (I37980,I38026,I38181);
DFFARX1 I_2088 (I117056,I2683,I38000,I38221,);
not I_2089 (I38229,I38221);
nor I_2090 (I37986,I38229,I38051);
nand I_2091 (I37974,I38229,I38164);
nand I_2092 (I38274,I117059,I117047);
and I_2093 (I38291,I38274,I117038);
DFFARX1 I_2094 (I38291,I2683,I38000,I38317,);
nor I_2095 (I38325,I38317,I38026);
DFFARX1 I_2096 (I38325,I2683,I38000,I37968,);
not I_2097 (I38356,I38317);
nor I_2098 (I38373,I117062,I117047);
not I_2099 (I38390,I38373);
nor I_2100 (I38407,I38164,I38390);
nor I_2101 (I38424,I38356,I38407);
DFFARX1 I_2102 (I38424,I2683,I38000,I37989,);
nor I_2103 (I38455,I38317,I38390);
nor I_2104 (I37977,I38181,I38455);
nor I_2105 (I37971,I38317,I38373);
not I_2106 (I38527,I2690);
DFFARX1 I_2107 (I729059,I2683,I38527,I38553,);
DFFARX1 I_2108 (I38553,I2683,I38527,I38570,);
not I_2109 (I38578,I38570);
nand I_2110 (I38595,I729035,I729062);
and I_2111 (I38612,I38595,I729047);
DFFARX1 I_2112 (I38612,I2683,I38527,I38638,);
DFFARX1 I_2113 (I38638,I2683,I38527,I38519,);
DFFARX1 I_2114 (I38638,I2683,I38527,I38510,);
DFFARX1 I_2115 (I729053,I2683,I38527,I38683,);
nand I_2116 (I38691,I38683,I729038);
not I_2117 (I38708,I38691);
nor I_2118 (I38507,I38553,I38708);
DFFARX1 I_2119 (I729056,I2683,I38527,I38748,);
not I_2120 (I38756,I38748);
nor I_2121 (I38513,I38756,I38578);
nand I_2122 (I38501,I38756,I38691);
nand I_2123 (I38801,I729041,I729044);
and I_2124 (I38818,I38801,I729035);
DFFARX1 I_2125 (I38818,I2683,I38527,I38844,);
nor I_2126 (I38852,I38844,I38553);
DFFARX1 I_2127 (I38852,I2683,I38527,I38495,);
not I_2128 (I38883,I38844);
nor I_2129 (I38900,I729050,I729044);
not I_2130 (I38917,I38900);
nor I_2131 (I38934,I38691,I38917);
nor I_2132 (I38951,I38883,I38934);
DFFARX1 I_2133 (I38951,I2683,I38527,I38516,);
nor I_2134 (I38982,I38844,I38917);
nor I_2135 (I38504,I38708,I38982);
nor I_2136 (I38498,I38844,I38900);
not I_2137 (I39054,I2690);
DFFARX1 I_2138 (I251192,I2683,I39054,I39080,);
DFFARX1 I_2139 (I39080,I2683,I39054,I39097,);
not I_2140 (I39105,I39097);
nand I_2141 (I39122,I251189,I251183);
and I_2142 (I39139,I39122,I251177);
DFFARX1 I_2143 (I39139,I2683,I39054,I39165,);
DFFARX1 I_2144 (I39165,I2683,I39054,I39046,);
DFFARX1 I_2145 (I39165,I2683,I39054,I39037,);
DFFARX1 I_2146 (I251165,I2683,I39054,I39210,);
nand I_2147 (I39218,I39210,I251174);
not I_2148 (I39235,I39218);
nor I_2149 (I39034,I39080,I39235);
DFFARX1 I_2150 (I251171,I2683,I39054,I39275,);
not I_2151 (I39283,I39275);
nor I_2152 (I39040,I39283,I39105);
nand I_2153 (I39028,I39283,I39218);
nand I_2154 (I39328,I251168,I251186);
and I_2155 (I39345,I39328,I251165);
DFFARX1 I_2156 (I39345,I2683,I39054,I39371,);
nor I_2157 (I39379,I39371,I39080);
DFFARX1 I_2158 (I39379,I2683,I39054,I39022,);
not I_2159 (I39410,I39371);
nor I_2160 (I39427,I251180,I251186);
not I_2161 (I39444,I39427);
nor I_2162 (I39461,I39218,I39444);
nor I_2163 (I39478,I39410,I39461);
DFFARX1 I_2164 (I39478,I2683,I39054,I39043,);
nor I_2165 (I39509,I39371,I39444);
nor I_2166 (I39031,I39235,I39509);
nor I_2167 (I39025,I39371,I39427);
not I_2168 (I39581,I2690);
DFFARX1 I_2169 (I595404,I2683,I39581,I39607,);
DFFARX1 I_2170 (I39607,I2683,I39581,I39624,);
not I_2171 (I39632,I39624);
nand I_2172 (I39649,I595419,I595422);
and I_2173 (I39666,I39649,I595401);
DFFARX1 I_2174 (I39666,I2683,I39581,I39692,);
DFFARX1 I_2175 (I39692,I2683,I39581,I39573,);
DFFARX1 I_2176 (I39692,I2683,I39581,I39564,);
DFFARX1 I_2177 (I595407,I2683,I39581,I39737,);
nand I_2178 (I39745,I39737,I595413);
not I_2179 (I39762,I39745);
nor I_2180 (I39561,I39607,I39762);
DFFARX1 I_2181 (I595401,I2683,I39581,I39802,);
not I_2182 (I39810,I39802);
nor I_2183 (I39567,I39810,I39632);
nand I_2184 (I39555,I39810,I39745);
nand I_2185 (I39855,I595416,I595398);
and I_2186 (I39872,I39855,I595410);
DFFARX1 I_2187 (I39872,I2683,I39581,I39898,);
nor I_2188 (I39906,I39898,I39607);
DFFARX1 I_2189 (I39906,I2683,I39581,I39549,);
not I_2190 (I39937,I39898);
nor I_2191 (I39954,I595398,I595398);
not I_2192 (I39971,I39954);
nor I_2193 (I39988,I39745,I39971);
nor I_2194 (I40005,I39937,I39988);
DFFARX1 I_2195 (I40005,I2683,I39581,I39570,);
nor I_2196 (I40036,I39898,I39971);
nor I_2197 (I39558,I39762,I40036);
nor I_2198 (I39552,I39898,I39954);
not I_2199 (I40108,I2690);
DFFARX1 I_2200 (I925902,I2683,I40108,I40134,);
DFFARX1 I_2201 (I40134,I2683,I40108,I40151,);
not I_2202 (I40159,I40151);
nand I_2203 (I40176,I925890,I925881);
and I_2204 (I40193,I40176,I925878);
DFFARX1 I_2205 (I40193,I2683,I40108,I40219,);
DFFARX1 I_2206 (I40219,I2683,I40108,I40100,);
DFFARX1 I_2207 (I40219,I2683,I40108,I40091,);
DFFARX1 I_2208 (I925884,I2683,I40108,I40264,);
nand I_2209 (I40272,I40264,I925896);
not I_2210 (I40289,I40272);
nor I_2211 (I40088,I40134,I40289);
DFFARX1 I_2212 (I925893,I2683,I40108,I40329,);
not I_2213 (I40337,I40329);
nor I_2214 (I40094,I40337,I40159);
nand I_2215 (I40082,I40337,I40272);
nand I_2216 (I40382,I925887,I925881);
and I_2217 (I40399,I40382,I925899);
DFFARX1 I_2218 (I40399,I2683,I40108,I40425,);
nor I_2219 (I40433,I40425,I40134);
DFFARX1 I_2220 (I40433,I2683,I40108,I40076,);
not I_2221 (I40464,I40425);
nor I_2222 (I40481,I925878,I925881);
not I_2223 (I40498,I40481);
nor I_2224 (I40515,I40272,I40498);
nor I_2225 (I40532,I40464,I40515);
DFFARX1 I_2226 (I40532,I2683,I40108,I40097,);
nor I_2227 (I40563,I40425,I40498);
nor I_2228 (I40085,I40289,I40563);
nor I_2229 (I40079,I40425,I40481);
not I_2230 (I40635,I2690);
DFFARX1 I_2231 (I736165,I2683,I40635,I40661,);
DFFARX1 I_2232 (I40661,I2683,I40635,I40678,);
not I_2233 (I40686,I40678);
nand I_2234 (I40703,I736141,I736168);
and I_2235 (I40720,I40703,I736153);
DFFARX1 I_2236 (I40720,I2683,I40635,I40746,);
DFFARX1 I_2237 (I40746,I2683,I40635,I40627,);
DFFARX1 I_2238 (I40746,I2683,I40635,I40618,);
DFFARX1 I_2239 (I736159,I2683,I40635,I40791,);
nand I_2240 (I40799,I40791,I736144);
not I_2241 (I40816,I40799);
nor I_2242 (I40615,I40661,I40816);
DFFARX1 I_2243 (I736162,I2683,I40635,I40856,);
not I_2244 (I40864,I40856);
nor I_2245 (I40621,I40864,I40686);
nand I_2246 (I40609,I40864,I40799);
nand I_2247 (I40909,I736147,I736150);
and I_2248 (I40926,I40909,I736141);
DFFARX1 I_2249 (I40926,I2683,I40635,I40952,);
nor I_2250 (I40960,I40952,I40661);
DFFARX1 I_2251 (I40960,I2683,I40635,I40603,);
not I_2252 (I40991,I40952);
nor I_2253 (I41008,I736156,I736150);
not I_2254 (I41025,I41008);
nor I_2255 (I41042,I40799,I41025);
nor I_2256 (I41059,I40991,I41042);
DFFARX1 I_2257 (I41059,I2683,I40635,I40624,);
nor I_2258 (I41090,I40952,I41025);
nor I_2259 (I40612,I40816,I41090);
nor I_2260 (I40606,I40952,I41008);
not I_2261 (I41162,I2690);
DFFARX1 I_2262 (I690777,I2683,I41162,I41188,);
DFFARX1 I_2263 (I41188,I2683,I41162,I41205,);
not I_2264 (I41213,I41205);
nand I_2265 (I41230,I690768,I690789);
and I_2266 (I41247,I41230,I690771);
DFFARX1 I_2267 (I41247,I2683,I41162,I41273,);
DFFARX1 I_2268 (I41273,I2683,I41162,I41154,);
DFFARX1 I_2269 (I41273,I2683,I41162,I41145,);
DFFARX1 I_2270 (I690771,I2683,I41162,I41318,);
nand I_2271 (I41326,I41318,I690786);
not I_2272 (I41343,I41326);
nor I_2273 (I41142,I41188,I41343);
DFFARX1 I_2274 (I690780,I2683,I41162,I41383,);
not I_2275 (I41391,I41383);
nor I_2276 (I41148,I41391,I41213);
nand I_2277 (I41136,I41391,I41326);
nand I_2278 (I41436,I690774,I690783);
and I_2279 (I41453,I41436,I690768);
DFFARX1 I_2280 (I41453,I2683,I41162,I41479,);
nor I_2281 (I41487,I41479,I41188);
DFFARX1 I_2282 (I41487,I2683,I41162,I41130,);
not I_2283 (I41518,I41479);
nor I_2284 (I41535,I690774,I690783);
not I_2285 (I41552,I41535);
nor I_2286 (I41569,I41326,I41552);
nor I_2287 (I41586,I41518,I41569);
DFFARX1 I_2288 (I41586,I2683,I41162,I41151,);
nor I_2289 (I41617,I41479,I41552);
nor I_2290 (I41139,I41343,I41617);
nor I_2291 (I41133,I41479,I41535);
not I_2292 (I41689,I2690);
DFFARX1 I_2293 (I695520,I2683,I41689,I41715,);
DFFARX1 I_2294 (I41715,I2683,I41689,I41732,);
not I_2295 (I41740,I41732);
nand I_2296 (I41757,I695511,I695532);
and I_2297 (I41774,I41757,I695514);
DFFARX1 I_2298 (I41774,I2683,I41689,I41800,);
DFFARX1 I_2299 (I41800,I2683,I41689,I41681,);
DFFARX1 I_2300 (I41800,I2683,I41689,I41672,);
DFFARX1 I_2301 (I695514,I2683,I41689,I41845,);
nand I_2302 (I41853,I41845,I695529);
not I_2303 (I41870,I41853);
nor I_2304 (I41669,I41715,I41870);
DFFARX1 I_2305 (I695523,I2683,I41689,I41910,);
not I_2306 (I41918,I41910);
nor I_2307 (I41675,I41918,I41740);
nand I_2308 (I41663,I41918,I41853);
nand I_2309 (I41963,I695517,I695526);
and I_2310 (I41980,I41963,I695511);
DFFARX1 I_2311 (I41980,I2683,I41689,I42006,);
nor I_2312 (I42014,I42006,I41715);
DFFARX1 I_2313 (I42014,I2683,I41689,I41657,);
not I_2314 (I42045,I42006);
nor I_2315 (I42062,I695517,I695526);
not I_2316 (I42079,I42062);
nor I_2317 (I42096,I41853,I42079);
nor I_2318 (I42113,I42045,I42096);
DFFARX1 I_2319 (I42113,I2683,I41689,I41678,);
nor I_2320 (I42144,I42006,I42079);
nor I_2321 (I41666,I41870,I42144);
nor I_2322 (I41660,I42006,I42062);
not I_2323 (I42216,I2690);
DFFARX1 I_2324 (I399686,I2683,I42216,I42242,);
DFFARX1 I_2325 (I42242,I2683,I42216,I42259,);
not I_2326 (I42267,I42259);
nand I_2327 (I42284,I399692,I399680);
and I_2328 (I42301,I42284,I399677);
DFFARX1 I_2329 (I42301,I2683,I42216,I42327,);
DFFARX1 I_2330 (I42327,I2683,I42216,I42208,);
DFFARX1 I_2331 (I42327,I2683,I42216,I42199,);
DFFARX1 I_2332 (I399689,I2683,I42216,I42372,);
nand I_2333 (I42380,I42372,I399683);
not I_2334 (I42397,I42380);
nor I_2335 (I42196,I42242,I42397);
DFFARX1 I_2336 (I399701,I2683,I42216,I42437,);
not I_2337 (I42445,I42437);
nor I_2338 (I42202,I42445,I42267);
nand I_2339 (I42190,I42445,I42380);
nand I_2340 (I42490,I399695,I399698);
and I_2341 (I42507,I42490,I399680);
DFFARX1 I_2342 (I42507,I2683,I42216,I42533,);
nor I_2343 (I42541,I42533,I42242);
DFFARX1 I_2344 (I42541,I2683,I42216,I42184,);
not I_2345 (I42572,I42533);
nor I_2346 (I42589,I399677,I399698);
not I_2347 (I42606,I42589);
nor I_2348 (I42623,I42380,I42606);
nor I_2349 (I42640,I42572,I42623);
DFFARX1 I_2350 (I42640,I2683,I42216,I42205,);
nor I_2351 (I42671,I42533,I42606);
nor I_2352 (I42193,I42397,I42671);
nor I_2353 (I42187,I42533,I42589);
not I_2354 (I42743,I2690);
DFFARX1 I_2355 (I871570,I2683,I42743,I42769,);
DFFARX1 I_2356 (I42769,I2683,I42743,I42786,);
not I_2357 (I42794,I42786);
nand I_2358 (I42811,I871558,I871549);
and I_2359 (I42828,I42811,I871546);
DFFARX1 I_2360 (I42828,I2683,I42743,I42854,);
DFFARX1 I_2361 (I42854,I2683,I42743,I42735,);
DFFARX1 I_2362 (I42854,I2683,I42743,I42726,);
DFFARX1 I_2363 (I871552,I2683,I42743,I42899,);
nand I_2364 (I42907,I42899,I871564);
not I_2365 (I42924,I42907);
nor I_2366 (I42723,I42769,I42924);
DFFARX1 I_2367 (I871561,I2683,I42743,I42964,);
not I_2368 (I42972,I42964);
nor I_2369 (I42729,I42972,I42794);
nand I_2370 (I42717,I42972,I42907);
nand I_2371 (I43017,I871555,I871549);
and I_2372 (I43034,I43017,I871567);
DFFARX1 I_2373 (I43034,I2683,I42743,I43060,);
nor I_2374 (I43068,I43060,I42769);
DFFARX1 I_2375 (I43068,I2683,I42743,I42711,);
not I_2376 (I43099,I43060);
nor I_2377 (I43116,I871546,I871549);
not I_2378 (I43133,I43116);
nor I_2379 (I43150,I42907,I43133);
nor I_2380 (I43167,I43099,I43150);
DFFARX1 I_2381 (I43167,I2683,I42743,I42732,);
nor I_2382 (I43198,I43060,I43133);
nor I_2383 (I42720,I42924,I43198);
nor I_2384 (I42714,I43060,I43116);
not I_2385 (I43270,I2690);
DFFARX1 I_2386 (I895846,I2683,I43270,I43296,);
DFFARX1 I_2387 (I43296,I2683,I43270,I43313,);
not I_2388 (I43321,I43313);
nand I_2389 (I43338,I895834,I895825);
and I_2390 (I43355,I43338,I895822);
DFFARX1 I_2391 (I43355,I2683,I43270,I43381,);
DFFARX1 I_2392 (I43381,I2683,I43270,I43262,);
DFFARX1 I_2393 (I43381,I2683,I43270,I43253,);
DFFARX1 I_2394 (I895828,I2683,I43270,I43426,);
nand I_2395 (I43434,I43426,I895840);
not I_2396 (I43451,I43434);
nor I_2397 (I43250,I43296,I43451);
DFFARX1 I_2398 (I895837,I2683,I43270,I43491,);
not I_2399 (I43499,I43491);
nor I_2400 (I43256,I43499,I43321);
nand I_2401 (I43244,I43499,I43434);
nand I_2402 (I43544,I895831,I895825);
and I_2403 (I43561,I43544,I895843);
DFFARX1 I_2404 (I43561,I2683,I43270,I43587,);
nor I_2405 (I43595,I43587,I43296);
DFFARX1 I_2406 (I43595,I2683,I43270,I43238,);
not I_2407 (I43626,I43587);
nor I_2408 (I43643,I895822,I895825);
not I_2409 (I43660,I43643);
nor I_2410 (I43677,I43434,I43660);
nor I_2411 (I43694,I43626,I43677);
DFFARX1 I_2412 (I43694,I2683,I43270,I43259,);
nor I_2413 (I43725,I43587,I43660);
nor I_2414 (I43247,I43451,I43725);
nor I_2415 (I43241,I43587,I43643);
not I_2416 (I43797,I2690);
DFFARX1 I_2417 (I814177,I2683,I43797,I43823,);
DFFARX1 I_2418 (I43823,I2683,I43797,I43840,);
not I_2419 (I43848,I43840);
nand I_2420 (I43865,I814171,I814192);
and I_2421 (I43882,I43865,I814177);
DFFARX1 I_2422 (I43882,I2683,I43797,I43908,);
DFFARX1 I_2423 (I43908,I2683,I43797,I43789,);
DFFARX1 I_2424 (I43908,I2683,I43797,I43780,);
DFFARX1 I_2425 (I814174,I2683,I43797,I43953,);
nand I_2426 (I43961,I43953,I814183);
not I_2427 (I43978,I43961);
nor I_2428 (I43777,I43823,I43978);
DFFARX1 I_2429 (I814171,I2683,I43797,I44018,);
not I_2430 (I44026,I44018);
nor I_2431 (I43783,I44026,I43848);
nand I_2432 (I43771,I44026,I43961);
nand I_2433 (I44071,I814174,I814189);
and I_2434 (I44088,I44071,I814180);
DFFARX1 I_2435 (I44088,I2683,I43797,I44114,);
nor I_2436 (I44122,I44114,I43823);
DFFARX1 I_2437 (I44122,I2683,I43797,I43765,);
not I_2438 (I44153,I44114);
nor I_2439 (I44170,I814186,I814189);
not I_2440 (I44187,I44170);
nor I_2441 (I44204,I43961,I44187);
nor I_2442 (I44221,I44153,I44204);
DFFARX1 I_2443 (I44221,I2683,I43797,I43786,);
nor I_2444 (I44252,I44114,I44187);
nor I_2445 (I43774,I43978,I44252);
nor I_2446 (I43768,I44114,I44170);
not I_2447 (I44324,I2690);
DFFARX1 I_2448 (I397901,I2683,I44324,I44350,);
DFFARX1 I_2449 (I44350,I2683,I44324,I44367,);
not I_2450 (I44375,I44367);
nand I_2451 (I44392,I397907,I397895);
and I_2452 (I44409,I44392,I397892);
DFFARX1 I_2453 (I44409,I2683,I44324,I44435,);
DFFARX1 I_2454 (I44435,I2683,I44324,I44316,);
DFFARX1 I_2455 (I44435,I2683,I44324,I44307,);
DFFARX1 I_2456 (I397904,I2683,I44324,I44480,);
nand I_2457 (I44488,I44480,I397898);
not I_2458 (I44505,I44488);
nor I_2459 (I44304,I44350,I44505);
DFFARX1 I_2460 (I397916,I2683,I44324,I44545,);
not I_2461 (I44553,I44545);
nor I_2462 (I44310,I44553,I44375);
nand I_2463 (I44298,I44553,I44488);
nand I_2464 (I44598,I397910,I397913);
and I_2465 (I44615,I44598,I397895);
DFFARX1 I_2466 (I44615,I2683,I44324,I44641,);
nor I_2467 (I44649,I44641,I44350);
DFFARX1 I_2468 (I44649,I2683,I44324,I44292,);
not I_2469 (I44680,I44641);
nor I_2470 (I44697,I397892,I397913);
not I_2471 (I44714,I44697);
nor I_2472 (I44731,I44488,I44714);
nor I_2473 (I44748,I44680,I44731);
DFFARX1 I_2474 (I44748,I2683,I44324,I44313,);
nor I_2475 (I44779,I44641,I44714);
nor I_2476 (I44301,I44505,I44779);
nor I_2477 (I44295,I44641,I44697);
not I_2478 (I44851,I2690);
DFFARX1 I_2479 (I62740,I2683,I44851,I44877,);
DFFARX1 I_2480 (I44877,I2683,I44851,I44894,);
not I_2481 (I44902,I44894);
nand I_2482 (I44919,I62740,I62755);
and I_2483 (I44936,I44919,I62758);
DFFARX1 I_2484 (I44936,I2683,I44851,I44962,);
DFFARX1 I_2485 (I44962,I2683,I44851,I44843,);
DFFARX1 I_2486 (I44962,I2683,I44851,I44834,);
DFFARX1 I_2487 (I62752,I2683,I44851,I45007,);
nand I_2488 (I45015,I45007,I62761);
not I_2489 (I45032,I45015);
nor I_2490 (I44831,I44877,I45032);
DFFARX1 I_2491 (I62737,I2683,I44851,I45072,);
not I_2492 (I45080,I45072);
nor I_2493 (I44837,I45080,I44902);
nand I_2494 (I44825,I45080,I45015);
nand I_2495 (I45125,I62737,I62743);
and I_2496 (I45142,I45125,I62746);
DFFARX1 I_2497 (I45142,I2683,I44851,I45168,);
nor I_2498 (I45176,I45168,I44877);
DFFARX1 I_2499 (I45176,I2683,I44851,I44819,);
not I_2500 (I45207,I45168);
nor I_2501 (I45224,I62749,I62743);
not I_2502 (I45241,I45224);
nor I_2503 (I45258,I45015,I45241);
nor I_2504 (I45275,I45207,I45258);
DFFARX1 I_2505 (I45275,I2683,I44851,I44840,);
nor I_2506 (I45306,I45168,I45241);
nor I_2507 (I44828,I45032,I45306);
nor I_2508 (I44822,I45168,I45224);
not I_2509 (I45378,I2690);
DFFARX1 I_2510 (I583266,I2683,I45378,I45404,);
DFFARX1 I_2511 (I45404,I2683,I45378,I45421,);
not I_2512 (I45429,I45421);
nand I_2513 (I45446,I583281,I583284);
and I_2514 (I45463,I45446,I583263);
DFFARX1 I_2515 (I45463,I2683,I45378,I45489,);
DFFARX1 I_2516 (I45489,I2683,I45378,I45370,);
DFFARX1 I_2517 (I45489,I2683,I45378,I45361,);
DFFARX1 I_2518 (I583269,I2683,I45378,I45534,);
nand I_2519 (I45542,I45534,I583275);
not I_2520 (I45559,I45542);
nor I_2521 (I45358,I45404,I45559);
DFFARX1 I_2522 (I583263,I2683,I45378,I45599,);
not I_2523 (I45607,I45599);
nor I_2524 (I45364,I45607,I45429);
nand I_2525 (I45352,I45607,I45542);
nand I_2526 (I45652,I583278,I583260);
and I_2527 (I45669,I45652,I583272);
DFFARX1 I_2528 (I45669,I2683,I45378,I45695,);
nor I_2529 (I45703,I45695,I45404);
DFFARX1 I_2530 (I45703,I2683,I45378,I45346,);
not I_2531 (I45734,I45695);
nor I_2532 (I45751,I583260,I583260);
not I_2533 (I45768,I45751);
nor I_2534 (I45785,I45542,I45768);
nor I_2535 (I45802,I45734,I45785);
DFFARX1 I_2536 (I45802,I2683,I45378,I45367,);
nor I_2537 (I45833,I45695,I45768);
nor I_2538 (I45355,I45559,I45833);
nor I_2539 (I45349,I45695,I45751);
not I_2540 (I45905,I2690);
DFFARX1 I_2541 (I738749,I2683,I45905,I45931,);
DFFARX1 I_2542 (I45931,I2683,I45905,I45948,);
not I_2543 (I45956,I45948);
nand I_2544 (I45973,I738725,I738752);
and I_2545 (I45990,I45973,I738737);
DFFARX1 I_2546 (I45990,I2683,I45905,I46016,);
DFFARX1 I_2547 (I46016,I2683,I45905,I45897,);
DFFARX1 I_2548 (I46016,I2683,I45905,I45888,);
DFFARX1 I_2549 (I738743,I2683,I45905,I46061,);
nand I_2550 (I46069,I46061,I738728);
not I_2551 (I46086,I46069);
nor I_2552 (I45885,I45931,I46086);
DFFARX1 I_2553 (I738746,I2683,I45905,I46126,);
not I_2554 (I46134,I46126);
nor I_2555 (I45891,I46134,I45956);
nand I_2556 (I45879,I46134,I46069);
nand I_2557 (I46179,I738731,I738734);
and I_2558 (I46196,I46179,I738725);
DFFARX1 I_2559 (I46196,I2683,I45905,I46222,);
nor I_2560 (I46230,I46222,I45931);
DFFARX1 I_2561 (I46230,I2683,I45905,I45873,);
not I_2562 (I46261,I46222);
nor I_2563 (I46278,I738740,I738734);
not I_2564 (I46295,I46278);
nor I_2565 (I46312,I46069,I46295);
nor I_2566 (I46329,I46261,I46312);
DFFARX1 I_2567 (I46329,I2683,I45905,I45894,);
nor I_2568 (I46360,I46222,I46295);
nor I_2569 (I45882,I46086,I46360);
nor I_2570 (I45876,I46222,I46278);
not I_2571 (I46432,I2690);
DFFARX1 I_2572 (I176547,I2683,I46432,I46458,);
not I_2573 (I46466,I46458);
nand I_2574 (I46483,I176541,I176535);
and I_2575 (I46500,I46483,I176556);
DFFARX1 I_2576 (I46500,I2683,I46432,I46526,);
DFFARX1 I_2577 (I176553,I2683,I46432,I46543,);
and I_2578 (I46551,I46543,I176550);
nor I_2579 (I46568,I46526,I46551);
DFFARX1 I_2580 (I46568,I2683,I46432,I46400,);
nand I_2581 (I46599,I46543,I176550);
nand I_2582 (I46616,I46466,I46599);
not I_2583 (I46412,I46616);
DFFARX1 I_2584 (I176535,I2683,I46432,I46656,);
DFFARX1 I_2585 (I46656,I2683,I46432,I46421,);
nand I_2586 (I46678,I176538,I176538);
and I_2587 (I46695,I46678,I176559);
DFFARX1 I_2588 (I46695,I2683,I46432,I46721,);
DFFARX1 I_2589 (I46721,I2683,I46432,I46738,);
not I_2590 (I46424,I46738);
not I_2591 (I46760,I46721);
nand I_2592 (I46409,I46760,I46599);
nor I_2593 (I46791,I176544,I176538);
not I_2594 (I46808,I46791);
nor I_2595 (I46825,I46760,I46808);
nor I_2596 (I46842,I46466,I46825);
DFFARX1 I_2597 (I46842,I2683,I46432,I46418,);
nor I_2598 (I46873,I46526,I46808);
nor I_2599 (I46406,I46721,I46873);
nor I_2600 (I46415,I46656,I46791);
nor I_2601 (I46403,I46526,I46791);
not I_2602 (I46959,I2690);
DFFARX1 I_2603 (I1588,I2683,I46959,I46985,);
not I_2604 (I46993,I46985);
nand I_2605 (I47010,I2036,I1724);
and I_2606 (I47027,I47010,I1540);
DFFARX1 I_2607 (I47027,I2683,I46959,I47053,);
DFFARX1 I_2608 (I1740,I2683,I46959,I47070,);
and I_2609 (I47078,I47070,I2252);
nor I_2610 (I47095,I47053,I47078);
DFFARX1 I_2611 (I47095,I2683,I46959,I46927,);
nand I_2612 (I47126,I47070,I2252);
nand I_2613 (I47143,I46993,I47126);
not I_2614 (I46939,I47143);
DFFARX1 I_2615 (I2148,I2683,I46959,I47183,);
DFFARX1 I_2616 (I47183,I2683,I46959,I46948,);
nand I_2617 (I47205,I1900,I1684);
and I_2618 (I47222,I47205,I1844);
DFFARX1 I_2619 (I47222,I2683,I46959,I47248,);
DFFARX1 I_2620 (I47248,I2683,I46959,I47265,);
not I_2621 (I46951,I47265);
not I_2622 (I47287,I47248);
nand I_2623 (I46936,I47287,I47126);
nor I_2624 (I47318,I2468,I1684);
not I_2625 (I47335,I47318);
nor I_2626 (I47352,I47287,I47335);
nor I_2627 (I47369,I46993,I47352);
DFFARX1 I_2628 (I47369,I2683,I46959,I46945,);
nor I_2629 (I47400,I47053,I47335);
nor I_2630 (I46933,I47248,I47400);
nor I_2631 (I46942,I47183,I47318);
nor I_2632 (I46930,I47053,I47318);
not I_2633 (I47486,I2690);
DFFARX1 I_2634 (I689723,I2683,I47486,I47512,);
not I_2635 (I47520,I47512);
nand I_2636 (I47537,I689720,I689735);
and I_2637 (I47554,I47537,I689717);
DFFARX1 I_2638 (I47554,I2683,I47486,I47580,);
DFFARX1 I_2639 (I689714,I2683,I47486,I47597,);
and I_2640 (I47605,I47597,I689714);
nor I_2641 (I47622,I47580,I47605);
DFFARX1 I_2642 (I47622,I2683,I47486,I47454,);
nand I_2643 (I47653,I47597,I689714);
nand I_2644 (I47670,I47520,I47653);
not I_2645 (I47466,I47670);
DFFARX1 I_2646 (I689717,I2683,I47486,I47710,);
DFFARX1 I_2647 (I47710,I2683,I47486,I47475,);
nand I_2648 (I47732,I689729,I689720);
and I_2649 (I47749,I47732,I689732);
DFFARX1 I_2650 (I47749,I2683,I47486,I47775,);
DFFARX1 I_2651 (I47775,I2683,I47486,I47792,);
not I_2652 (I47478,I47792);
not I_2653 (I47814,I47775);
nand I_2654 (I47463,I47814,I47653);
nor I_2655 (I47845,I689726,I689720);
not I_2656 (I47862,I47845);
nor I_2657 (I47879,I47814,I47862);
nor I_2658 (I47896,I47520,I47879);
DFFARX1 I_2659 (I47896,I2683,I47486,I47472,);
nor I_2660 (I47927,I47580,I47862);
nor I_2661 (I47460,I47775,I47927);
nor I_2662 (I47469,I47710,I47845);
nor I_2663 (I47457,I47580,I47845);
not I_2664 (I48013,I2690);
DFFARX1 I_2665 (I960292,I2683,I48013,I48039,);
not I_2666 (I48047,I48039);
nand I_2667 (I48064,I960286,I960307);
and I_2668 (I48081,I48064,I960298);
DFFARX1 I_2669 (I48081,I2683,I48013,I48107,);
DFFARX1 I_2670 (I960289,I2683,I48013,I48124,);
and I_2671 (I48132,I48124,I960301);
nor I_2672 (I48149,I48107,I48132);
DFFARX1 I_2673 (I48149,I2683,I48013,I47981,);
nand I_2674 (I48180,I48124,I960301);
nand I_2675 (I48197,I48047,I48180);
not I_2676 (I47993,I48197);
DFFARX1 I_2677 (I960289,I2683,I48013,I48237,);
DFFARX1 I_2678 (I48237,I2683,I48013,I48002,);
nand I_2679 (I48259,I960310,I960295);
and I_2680 (I48276,I48259,I960286);
DFFARX1 I_2681 (I48276,I2683,I48013,I48302,);
DFFARX1 I_2682 (I48302,I2683,I48013,I48319,);
not I_2683 (I48005,I48319);
not I_2684 (I48341,I48302);
nand I_2685 (I47990,I48341,I48180);
nor I_2686 (I48372,I960304,I960295);
not I_2687 (I48389,I48372);
nor I_2688 (I48406,I48341,I48389);
nor I_2689 (I48423,I48047,I48406);
DFFARX1 I_2690 (I48423,I2683,I48013,I47999,);
nor I_2691 (I48454,I48107,I48389);
nor I_2692 (I47987,I48302,I48454);
nor I_2693 (I47996,I48237,I48372);
nor I_2694 (I47984,I48107,I48372);
not I_2695 (I48540,I2690);
DFFARX1 I_2696 (I594832,I2683,I48540,I48566,);
not I_2697 (I48574,I48566);
nand I_2698 (I48591,I594823,I594841);
and I_2699 (I48608,I48591,I594820);
DFFARX1 I_2700 (I48608,I2683,I48540,I48634,);
DFFARX1 I_2701 (I594823,I2683,I48540,I48651,);
and I_2702 (I48659,I48651,I594826);
nor I_2703 (I48676,I48634,I48659);
DFFARX1 I_2704 (I48676,I2683,I48540,I48508,);
nand I_2705 (I48707,I48651,I594826);
nand I_2706 (I48724,I48574,I48707);
not I_2707 (I48520,I48724);
DFFARX1 I_2708 (I594820,I2683,I48540,I48764,);
DFFARX1 I_2709 (I48764,I2683,I48540,I48529,);
nand I_2710 (I48786,I594838,I594829);
and I_2711 (I48803,I48786,I594844);
DFFARX1 I_2712 (I48803,I2683,I48540,I48829,);
DFFARX1 I_2713 (I48829,I2683,I48540,I48846,);
not I_2714 (I48532,I48846);
not I_2715 (I48868,I48829);
nand I_2716 (I48517,I48868,I48707);
nor I_2717 (I48899,I594835,I594829);
not I_2718 (I48916,I48899);
nor I_2719 (I48933,I48868,I48916);
nor I_2720 (I48950,I48574,I48933);
DFFARX1 I_2721 (I48950,I2683,I48540,I48526,);
nor I_2722 (I48981,I48634,I48916);
nor I_2723 (I48514,I48829,I48981);
nor I_2724 (I48523,I48764,I48899);
nor I_2725 (I48511,I48634,I48899);
not I_2726 (I49067,I2690);
DFFARX1 I_2727 (I114081,I2683,I49067,I49093,);
not I_2728 (I49101,I49093);
nand I_2729 (I49118,I114078,I114060);
and I_2730 (I49135,I49118,I114066);
DFFARX1 I_2731 (I49135,I2683,I49067,I49161,);
DFFARX1 I_2732 (I114075,I2683,I49067,I49178,);
and I_2733 (I49186,I49178,I114069);
nor I_2734 (I49203,I49161,I49186);
DFFARX1 I_2735 (I49203,I2683,I49067,I49035,);
nand I_2736 (I49234,I49178,I114069);
nand I_2737 (I49251,I49101,I49234);
not I_2738 (I49047,I49251);
DFFARX1 I_2739 (I114084,I2683,I49067,I49291,);
DFFARX1 I_2740 (I49291,I2683,I49067,I49056,);
nand I_2741 (I49313,I114072,I114063);
and I_2742 (I49330,I49313,I114060);
DFFARX1 I_2743 (I49330,I2683,I49067,I49356,);
DFFARX1 I_2744 (I49356,I2683,I49067,I49373,);
not I_2745 (I49059,I49373);
not I_2746 (I49395,I49356);
nand I_2747 (I49044,I49395,I49234);
nor I_2748 (I49426,I114087,I114063);
not I_2749 (I49443,I49426);
nor I_2750 (I49460,I49395,I49443);
nor I_2751 (I49477,I49101,I49460);
DFFARX1 I_2752 (I49477,I2683,I49067,I49053,);
nor I_2753 (I49508,I49161,I49443);
nor I_2754 (I49041,I49356,I49508);
nor I_2755 (I49050,I49291,I49426);
nor I_2756 (I49038,I49161,I49426);
not I_2757 (I49594,I2690);
DFFARX1 I_2758 (I421100,I2683,I49594,I49620,);
not I_2759 (I49628,I49620);
nand I_2760 (I49645,I421121,I421115);
and I_2761 (I49662,I49645,I421097);
DFFARX1 I_2762 (I49662,I2683,I49594,I49688,);
DFFARX1 I_2763 (I421100,I2683,I49594,I49705,);
and I_2764 (I49713,I49705,I421109);
nor I_2765 (I49730,I49688,I49713);
DFFARX1 I_2766 (I49730,I2683,I49594,I49562,);
nand I_2767 (I49761,I49705,I421109);
nand I_2768 (I49778,I49628,I49761);
not I_2769 (I49574,I49778);
DFFARX1 I_2770 (I421106,I2683,I49594,I49818,);
DFFARX1 I_2771 (I49818,I2683,I49594,I49583,);
nand I_2772 (I49840,I421112,I421103);
and I_2773 (I49857,I49840,I421097);
DFFARX1 I_2774 (I49857,I2683,I49594,I49883,);
DFFARX1 I_2775 (I49883,I2683,I49594,I49900,);
not I_2776 (I49586,I49900);
not I_2777 (I49922,I49883);
nand I_2778 (I49571,I49922,I49761);
nor I_2779 (I49953,I421118,I421103);
not I_2780 (I49970,I49953);
nor I_2781 (I49987,I49922,I49970);
nor I_2782 (I50004,I49628,I49987);
DFFARX1 I_2783 (I50004,I2683,I49594,I49580,);
nor I_2784 (I50035,I49688,I49970);
nor I_2785 (I49568,I49883,I50035);
nor I_2786 (I49577,I49818,I49953);
nor I_2787 (I49565,I49688,I49953);
not I_2788 (I50121,I2690);
DFFARX1 I_2789 (I634388,I2683,I50121,I50147,);
not I_2790 (I50155,I50147);
nand I_2791 (I50172,I634385,I634400);
and I_2792 (I50189,I50172,I634382);
DFFARX1 I_2793 (I50189,I2683,I50121,I50215,);
DFFARX1 I_2794 (I634379,I2683,I50121,I50232,);
and I_2795 (I50240,I50232,I634379);
nor I_2796 (I50257,I50215,I50240);
DFFARX1 I_2797 (I50257,I2683,I50121,I50089,);
nand I_2798 (I50288,I50232,I634379);
nand I_2799 (I50305,I50155,I50288);
not I_2800 (I50101,I50305);
DFFARX1 I_2801 (I634382,I2683,I50121,I50345,);
DFFARX1 I_2802 (I50345,I2683,I50121,I50110,);
nand I_2803 (I50367,I634394,I634385);
and I_2804 (I50384,I50367,I634397);
DFFARX1 I_2805 (I50384,I2683,I50121,I50410,);
DFFARX1 I_2806 (I50410,I2683,I50121,I50427,);
not I_2807 (I50113,I50427);
not I_2808 (I50449,I50410);
nand I_2809 (I50098,I50449,I50288);
nor I_2810 (I50480,I634391,I634385);
not I_2811 (I50497,I50480);
nor I_2812 (I50514,I50449,I50497);
nor I_2813 (I50531,I50155,I50514);
DFFARX1 I_2814 (I50531,I2683,I50121,I50107,);
nor I_2815 (I50562,I50215,I50497);
nor I_2816 (I50095,I50410,I50562);
nor I_2817 (I50104,I50345,I50480);
nor I_2818 (I50092,I50215,I50480);
not I_2819 (I50648,I2690);
DFFARX1 I_2820 (I680764,I2683,I50648,I50674,);
not I_2821 (I50682,I50674);
nand I_2822 (I50699,I680761,I680776);
and I_2823 (I50716,I50699,I680758);
DFFARX1 I_2824 (I50716,I2683,I50648,I50742,);
DFFARX1 I_2825 (I680755,I2683,I50648,I50759,);
and I_2826 (I50767,I50759,I680755);
nor I_2827 (I50784,I50742,I50767);
DFFARX1 I_2828 (I50784,I2683,I50648,I50616,);
nand I_2829 (I50815,I50759,I680755);
nand I_2830 (I50832,I50682,I50815);
not I_2831 (I50628,I50832);
DFFARX1 I_2832 (I680758,I2683,I50648,I50872,);
DFFARX1 I_2833 (I50872,I2683,I50648,I50637,);
nand I_2834 (I50894,I680770,I680761);
and I_2835 (I50911,I50894,I680773);
DFFARX1 I_2836 (I50911,I2683,I50648,I50937,);
DFFARX1 I_2837 (I50937,I2683,I50648,I50954,);
not I_2838 (I50640,I50954);
not I_2839 (I50976,I50937);
nand I_2840 (I50625,I50976,I50815);
nor I_2841 (I51007,I680767,I680761);
not I_2842 (I51024,I51007);
nor I_2843 (I51041,I50976,I51024);
nor I_2844 (I51058,I50682,I51041);
DFFARX1 I_2845 (I51058,I2683,I50648,I50634,);
nor I_2846 (I51089,I50742,I51024);
nor I_2847 (I50622,I50937,I51089);
nor I_2848 (I50631,I50872,I51007);
nor I_2849 (I50619,I50742,I51007);
not I_2850 (I51175,I2690);
DFFARX1 I_2851 (I225896,I2683,I51175,I51201,);
not I_2852 (I51209,I51201);
nand I_2853 (I51226,I225878,I225893);
and I_2854 (I51243,I51226,I225869);
DFFARX1 I_2855 (I51243,I2683,I51175,I51269,);
DFFARX1 I_2856 (I225872,I2683,I51175,I51286,);
and I_2857 (I51294,I51286,I225887);
nor I_2858 (I51311,I51269,I51294);
DFFARX1 I_2859 (I51311,I2683,I51175,I51143,);
nand I_2860 (I51342,I51286,I225887);
nand I_2861 (I51359,I51209,I51342);
not I_2862 (I51155,I51359);
DFFARX1 I_2863 (I225890,I2683,I51175,I51399,);
DFFARX1 I_2864 (I51399,I2683,I51175,I51164,);
nand I_2865 (I51421,I225869,I225881);
and I_2866 (I51438,I51421,I225875);
DFFARX1 I_2867 (I51438,I2683,I51175,I51464,);
DFFARX1 I_2868 (I51464,I2683,I51175,I51481,);
not I_2869 (I51167,I51481);
not I_2870 (I51503,I51464);
nand I_2871 (I51152,I51503,I51342);
nor I_2872 (I51534,I225884,I225881);
not I_2873 (I51551,I51534);
nor I_2874 (I51568,I51503,I51551);
nor I_2875 (I51585,I51209,I51568);
DFFARX1 I_2876 (I51585,I2683,I51175,I51161,);
nor I_2877 (I51616,I51269,I51551);
nor I_2878 (I51149,I51464,I51616);
nor I_2879 (I51158,I51399,I51534);
nor I_2880 (I51146,I51269,I51534);
not I_2881 (I51702,I2690);
DFFARX1 I_2882 (I330148,I2683,I51702,I51728,);
not I_2883 (I51736,I51728);
nand I_2884 (I51753,I330142,I330133);
and I_2885 (I51770,I51753,I330154);
DFFARX1 I_2886 (I51770,I2683,I51702,I51796,);
DFFARX1 I_2887 (I330136,I2683,I51702,I51813,);
and I_2888 (I51821,I51813,I330130);
nor I_2889 (I51838,I51796,I51821);
DFFARX1 I_2890 (I51838,I2683,I51702,I51670,);
nand I_2891 (I51869,I51813,I330130);
nand I_2892 (I51886,I51736,I51869);
not I_2893 (I51682,I51886);
DFFARX1 I_2894 (I330130,I2683,I51702,I51926,);
DFFARX1 I_2895 (I51926,I2683,I51702,I51691,);
nand I_2896 (I51948,I330157,I330139);
and I_2897 (I51965,I51948,I330145);
DFFARX1 I_2898 (I51965,I2683,I51702,I51991,);
DFFARX1 I_2899 (I51991,I2683,I51702,I52008,);
not I_2900 (I51694,I52008);
not I_2901 (I52030,I51991);
nand I_2902 (I51679,I52030,I51869);
nor I_2903 (I52061,I330151,I330139);
not I_2904 (I52078,I52061);
nor I_2905 (I52095,I52030,I52078);
nor I_2906 (I52112,I51736,I52095);
DFFARX1 I_2907 (I52112,I2683,I51702,I51688,);
nor I_2908 (I52143,I51796,I52078);
nor I_2909 (I51676,I51991,I52143);
nor I_2910 (I51685,I51926,I52061);
nor I_2911 (I51673,I51796,I52061);
not I_2912 (I52229,I2690);
DFFARX1 I_2913 (I15858,I2683,I52229,I52255,);
not I_2914 (I52263,I52255);
nand I_2915 (I52280,I15846,I15852);
and I_2916 (I52297,I52280,I15855);
DFFARX1 I_2917 (I52297,I2683,I52229,I52323,);
DFFARX1 I_2918 (I15837,I2683,I52229,I52340,);
and I_2919 (I52348,I52340,I15843);
nor I_2920 (I52365,I52323,I52348);
DFFARX1 I_2921 (I52365,I2683,I52229,I52197,);
nand I_2922 (I52396,I52340,I15843);
nand I_2923 (I52413,I52263,I52396);
not I_2924 (I52209,I52413);
DFFARX1 I_2925 (I15837,I2683,I52229,I52453,);
DFFARX1 I_2926 (I52453,I2683,I52229,I52218,);
nand I_2927 (I52475,I15840,I15834);
and I_2928 (I52492,I52475,I15849);
DFFARX1 I_2929 (I52492,I2683,I52229,I52518,);
DFFARX1 I_2930 (I52518,I2683,I52229,I52535,);
not I_2931 (I52221,I52535);
not I_2932 (I52557,I52518);
nand I_2933 (I52206,I52557,I52396);
nor I_2934 (I52588,I15834,I15834);
not I_2935 (I52605,I52588);
nor I_2936 (I52622,I52557,I52605);
nor I_2937 (I52639,I52263,I52622);
DFFARX1 I_2938 (I52639,I2683,I52229,I52215,);
nor I_2939 (I52670,I52323,I52605);
nor I_2940 (I52203,I52518,I52670);
nor I_2941 (I52212,I52453,I52588);
nor I_2942 (I52200,I52323,I52588);
not I_2943 (I52756,I2690);
DFFARX1 I_2944 (I300730,I2683,I52756,I52782,);
not I_2945 (I52790,I52782);
nand I_2946 (I52807,I300712,I300727);
and I_2947 (I52824,I52807,I300703);
DFFARX1 I_2948 (I52824,I2683,I52756,I52850,);
DFFARX1 I_2949 (I300706,I2683,I52756,I52867,);
and I_2950 (I52875,I52867,I300721);
nor I_2951 (I52892,I52850,I52875);
DFFARX1 I_2952 (I52892,I2683,I52756,I52724,);
nand I_2953 (I52923,I52867,I300721);
nand I_2954 (I52940,I52790,I52923);
not I_2955 (I52736,I52940);
DFFARX1 I_2956 (I300724,I2683,I52756,I52980,);
DFFARX1 I_2957 (I52980,I2683,I52756,I52745,);
nand I_2958 (I53002,I300703,I300715);
and I_2959 (I53019,I53002,I300709);
DFFARX1 I_2960 (I53019,I2683,I52756,I53045,);
DFFARX1 I_2961 (I53045,I2683,I52756,I53062,);
not I_2962 (I52748,I53062);
not I_2963 (I53084,I53045);
nand I_2964 (I52733,I53084,I52923);
nor I_2965 (I53115,I300718,I300715);
not I_2966 (I53132,I53115);
nor I_2967 (I53149,I53084,I53132);
nor I_2968 (I53166,I52790,I53149);
DFFARX1 I_2969 (I53166,I2683,I52756,I52742,);
nor I_2970 (I53197,I52850,I53132);
nor I_2971 (I52730,I53045,I53197);
nor I_2972 (I52739,I52980,I53115);
nor I_2973 (I52727,I52850,I53115);
not I_2974 (I53283,I2690);
DFFARX1 I_2975 (I544546,I2683,I53283,I53309,);
not I_2976 (I53317,I53309);
nand I_2977 (I53334,I544537,I544555);
and I_2978 (I53351,I53334,I544534);
DFFARX1 I_2979 (I53351,I2683,I53283,I53377,);
DFFARX1 I_2980 (I544537,I2683,I53283,I53394,);
and I_2981 (I53402,I53394,I544540);
nor I_2982 (I53419,I53377,I53402);
DFFARX1 I_2983 (I53419,I2683,I53283,I53251,);
nand I_2984 (I53450,I53394,I544540);
nand I_2985 (I53467,I53317,I53450);
not I_2986 (I53263,I53467);
DFFARX1 I_2987 (I544534,I2683,I53283,I53507,);
DFFARX1 I_2988 (I53507,I2683,I53283,I53272,);
nand I_2989 (I53529,I544552,I544543);
and I_2990 (I53546,I53529,I544558);
DFFARX1 I_2991 (I53546,I2683,I53283,I53572,);
DFFARX1 I_2992 (I53572,I2683,I53283,I53589,);
not I_2993 (I53275,I53589);
not I_2994 (I53611,I53572);
nand I_2995 (I53260,I53611,I53450);
nor I_2996 (I53642,I544549,I544543);
not I_2997 (I53659,I53642);
nor I_2998 (I53676,I53611,I53659);
nor I_2999 (I53693,I53317,I53676);
DFFARX1 I_3000 (I53693,I2683,I53283,I53269,);
nor I_3001 (I53724,I53377,I53659);
nor I_3002 (I53257,I53572,I53724);
nor I_3003 (I53266,I53507,I53642);
nor I_3004 (I53254,I53377,I53642);
not I_3005 (I53810,I2690);
DFFARX1 I_3006 (I464779,I2683,I53810,I53836,);
not I_3007 (I53844,I53836);
nand I_3008 (I53861,I464791,I464776);
and I_3009 (I53878,I53861,I464770);
DFFARX1 I_3010 (I53878,I2683,I53810,I53904,);
DFFARX1 I_3011 (I464785,I2683,I53810,I53921,);
and I_3012 (I53929,I53921,I464773);
nor I_3013 (I53946,I53904,I53929);
DFFARX1 I_3014 (I53946,I2683,I53810,I53778,);
nand I_3015 (I53977,I53921,I464773);
nand I_3016 (I53994,I53844,I53977);
not I_3017 (I53790,I53994);
DFFARX1 I_3018 (I464782,I2683,I53810,I54034,);
DFFARX1 I_3019 (I54034,I2683,I53810,I53799,);
nand I_3020 (I54056,I464788,I464794);
and I_3021 (I54073,I54056,I464770);
DFFARX1 I_3022 (I54073,I2683,I53810,I54099,);
DFFARX1 I_3023 (I54099,I2683,I53810,I54116,);
not I_3024 (I53802,I54116);
not I_3025 (I54138,I54099);
nand I_3026 (I53787,I54138,I53977);
nor I_3027 (I54169,I464773,I464794);
not I_3028 (I54186,I54169);
nor I_3029 (I54203,I54138,I54186);
nor I_3030 (I54220,I53844,I54203);
DFFARX1 I_3031 (I54220,I2683,I53810,I53796,);
nor I_3032 (I54251,I53904,I54186);
nor I_3033 (I53784,I54099,I54251);
nor I_3034 (I53793,I54034,I54169);
nor I_3035 (I53781,I53904,I54169);
not I_3036 (I54337,I2690);
DFFARX1 I_3037 (I268056,I2683,I54337,I54363,);
not I_3038 (I54371,I54363);
nand I_3039 (I54388,I268038,I268053);
and I_3040 (I54405,I54388,I268029);
DFFARX1 I_3041 (I54405,I2683,I54337,I54431,);
DFFARX1 I_3042 (I268032,I2683,I54337,I54448,);
and I_3043 (I54456,I54448,I268047);
nor I_3044 (I54473,I54431,I54456);
DFFARX1 I_3045 (I54473,I2683,I54337,I54305,);
nand I_3046 (I54504,I54448,I268047);
nand I_3047 (I54521,I54371,I54504);
not I_3048 (I54317,I54521);
DFFARX1 I_3049 (I268050,I2683,I54337,I54561,);
DFFARX1 I_3050 (I54561,I2683,I54337,I54326,);
nand I_3051 (I54583,I268029,I268041);
and I_3052 (I54600,I54583,I268035);
DFFARX1 I_3053 (I54600,I2683,I54337,I54626,);
DFFARX1 I_3054 (I54626,I2683,I54337,I54643,);
not I_3055 (I54329,I54643);
not I_3056 (I54665,I54626);
nand I_3057 (I54314,I54665,I54504);
nor I_3058 (I54696,I268044,I268041);
not I_3059 (I54713,I54696);
nor I_3060 (I54730,I54665,I54713);
nor I_3061 (I54747,I54371,I54730);
DFFARX1 I_3062 (I54747,I2683,I54337,I54323,);
nor I_3063 (I54778,I54431,I54713);
nor I_3064 (I54311,I54626,I54778);
nor I_3065 (I54320,I54561,I54696);
nor I_3066 (I54308,I54431,I54696);
not I_3067 (I54864,I2690);
DFFARX1 I_3068 (I526050,I2683,I54864,I54890,);
not I_3069 (I54898,I54890);
nand I_3070 (I54915,I526041,I526059);
and I_3071 (I54932,I54915,I526038);
DFFARX1 I_3072 (I54932,I2683,I54864,I54958,);
DFFARX1 I_3073 (I526041,I2683,I54864,I54975,);
and I_3074 (I54983,I54975,I526044);
nor I_3075 (I55000,I54958,I54983);
DFFARX1 I_3076 (I55000,I2683,I54864,I54832,);
nand I_3077 (I55031,I54975,I526044);
nand I_3078 (I55048,I54898,I55031);
not I_3079 (I54844,I55048);
DFFARX1 I_3080 (I526038,I2683,I54864,I55088,);
DFFARX1 I_3081 (I55088,I2683,I54864,I54853,);
nand I_3082 (I55110,I526056,I526047);
and I_3083 (I55127,I55110,I526062);
DFFARX1 I_3084 (I55127,I2683,I54864,I55153,);
DFFARX1 I_3085 (I55153,I2683,I54864,I55170,);
not I_3086 (I54856,I55170);
not I_3087 (I55192,I55153);
nand I_3088 (I54841,I55192,I55031);
nor I_3089 (I55223,I526053,I526047);
not I_3090 (I55240,I55223);
nor I_3091 (I55257,I55192,I55240);
nor I_3092 (I55274,I54898,I55257);
DFFARX1 I_3093 (I55274,I2683,I54864,I54850,);
nor I_3094 (I55305,I54958,I55240);
nor I_3095 (I54838,I55153,I55305);
nor I_3096 (I54847,I55088,I55223);
nor I_3097 (I54835,I54958,I55223);
not I_3098 (I55391,I2690);
DFFARX1 I_3099 (I1079876,I2683,I55391,I55417,);
not I_3100 (I55425,I55417);
nand I_3101 (I55442,I1079870,I1079891);
and I_3102 (I55459,I55442,I1079867);
DFFARX1 I_3103 (I55459,I2683,I55391,I55485,);
DFFARX1 I_3104 (I1079888,I2683,I55391,I55502,);
and I_3105 (I55510,I55502,I1079885);
nor I_3106 (I55527,I55485,I55510);
DFFARX1 I_3107 (I55527,I2683,I55391,I55359,);
nand I_3108 (I55558,I55502,I1079885);
nand I_3109 (I55575,I55425,I55558);
not I_3110 (I55371,I55575);
DFFARX1 I_3111 (I1079873,I2683,I55391,I55615,);
DFFARX1 I_3112 (I55615,I2683,I55391,I55380,);
nand I_3113 (I55637,I1079882,I1079879);
and I_3114 (I55654,I55637,I1079864);
DFFARX1 I_3115 (I55654,I2683,I55391,I55680,);
DFFARX1 I_3116 (I55680,I2683,I55391,I55697,);
not I_3117 (I55383,I55697);
not I_3118 (I55719,I55680);
nand I_3119 (I55368,I55719,I55558);
nor I_3120 (I55750,I1079864,I1079879);
not I_3121 (I55767,I55750);
nor I_3122 (I55784,I55719,I55767);
nor I_3123 (I55801,I55425,I55784);
DFFARX1 I_3124 (I55801,I2683,I55391,I55377,);
nor I_3125 (I55832,I55485,I55767);
nor I_3126 (I55365,I55680,I55832);
nor I_3127 (I55374,I55615,I55750);
nor I_3128 (I55362,I55485,I55750);
not I_3129 (I55918,I2690);
DFFARX1 I_3130 (I774910,I2683,I55918,I55944,);
not I_3131 (I55952,I55944);
nand I_3132 (I55969,I774928,I774922);
and I_3133 (I55986,I55969,I774901);
DFFARX1 I_3134 (I55986,I2683,I55918,I56012,);
DFFARX1 I_3135 (I774919,I2683,I55918,I56029,);
and I_3136 (I56037,I56029,I774904);
nor I_3137 (I56054,I56012,I56037);
DFFARX1 I_3138 (I56054,I2683,I55918,I55886,);
nand I_3139 (I56085,I56029,I774904);
nand I_3140 (I56102,I55952,I56085);
not I_3141 (I55898,I56102);
DFFARX1 I_3142 (I774916,I2683,I55918,I56142,);
DFFARX1 I_3143 (I56142,I2683,I55918,I55907,);
nand I_3144 (I56164,I774925,I774913);
and I_3145 (I56181,I56164,I774907);
DFFARX1 I_3146 (I56181,I2683,I55918,I56207,);
DFFARX1 I_3147 (I56207,I2683,I55918,I56224,);
not I_3148 (I55910,I56224);
not I_3149 (I56246,I56207);
nand I_3150 (I55895,I56246,I56085);
nor I_3151 (I56277,I774901,I774913);
not I_3152 (I56294,I56277);
nor I_3153 (I56311,I56246,I56294);
nor I_3154 (I56328,I55952,I56311);
DFFARX1 I_3155 (I56328,I2683,I55918,I55904,);
nor I_3156 (I56359,I56012,I56294);
nor I_3157 (I55892,I56207,I56359);
nor I_3158 (I55901,I56142,I56277);
nor I_3159 (I55889,I56012,I56277);
not I_3160 (I56445,I2690);
DFFARX1 I_3161 (I855368,I2683,I56445,I56471,);
not I_3162 (I56479,I56471);
nand I_3163 (I56496,I855383,I855362);
and I_3164 (I56513,I56496,I855365);
DFFARX1 I_3165 (I56513,I2683,I56445,I56539,);
DFFARX1 I_3166 (I855386,I2683,I56445,I56556,);
and I_3167 (I56564,I56556,I855365);
nor I_3168 (I56581,I56539,I56564);
DFFARX1 I_3169 (I56581,I2683,I56445,I56413,);
nand I_3170 (I56612,I56556,I855365);
nand I_3171 (I56629,I56479,I56612);
not I_3172 (I56425,I56629);
DFFARX1 I_3173 (I855362,I2683,I56445,I56669,);
DFFARX1 I_3174 (I56669,I2683,I56445,I56434,);
nand I_3175 (I56691,I855374,I855371);
and I_3176 (I56708,I56691,I855377);
DFFARX1 I_3177 (I56708,I2683,I56445,I56734,);
DFFARX1 I_3178 (I56734,I2683,I56445,I56751,);
not I_3179 (I56437,I56751);
not I_3180 (I56773,I56734);
nand I_3181 (I56422,I56773,I56612);
nor I_3182 (I56804,I855380,I855371);
not I_3183 (I56821,I56804);
nor I_3184 (I56838,I56773,I56821);
nor I_3185 (I56855,I56479,I56838);
DFFARX1 I_3186 (I56855,I2683,I56445,I56431,);
nor I_3187 (I56886,I56539,I56821);
nor I_3188 (I56419,I56734,I56886);
nor I_3189 (I56428,I56669,I56804);
nor I_3190 (I56416,I56539,I56804);
not I_3191 (I56972,I2690);
DFFARX1 I_3192 (I486743,I2683,I56972,I56998,);
not I_3193 (I57006,I56998);
nand I_3194 (I57023,I486755,I486740);
and I_3195 (I57040,I57023,I486734);
DFFARX1 I_3196 (I57040,I2683,I56972,I57066,);
DFFARX1 I_3197 (I486749,I2683,I56972,I57083,);
and I_3198 (I57091,I57083,I486737);
nor I_3199 (I57108,I57066,I57091);
DFFARX1 I_3200 (I57108,I2683,I56972,I56940,);
nand I_3201 (I57139,I57083,I486737);
nand I_3202 (I57156,I57006,I57139);
not I_3203 (I56952,I57156);
DFFARX1 I_3204 (I486746,I2683,I56972,I57196,);
DFFARX1 I_3205 (I57196,I2683,I56972,I56961,);
nand I_3206 (I57218,I486752,I486758);
and I_3207 (I57235,I57218,I486734);
DFFARX1 I_3208 (I57235,I2683,I56972,I57261,);
DFFARX1 I_3209 (I57261,I2683,I56972,I57278,);
not I_3210 (I56964,I57278);
not I_3211 (I57300,I57261);
nand I_3212 (I56949,I57300,I57139);
nor I_3213 (I57331,I486737,I486758);
not I_3214 (I57348,I57331);
nor I_3215 (I57365,I57300,I57348);
nor I_3216 (I57382,I57006,I57365);
DFFARX1 I_3217 (I57382,I2683,I56972,I56958,);
nor I_3218 (I57413,I57066,I57348);
nor I_3219 (I56946,I57261,I57413);
nor I_3220 (I56955,I57196,I57331);
nor I_3221 (I56943,I57066,I57331);
not I_3222 (I57499,I2690);
DFFARX1 I_3223 (I524316,I2683,I57499,I57525,);
not I_3224 (I57533,I57525);
nand I_3225 (I57550,I524307,I524325);
and I_3226 (I57567,I57550,I524304);
DFFARX1 I_3227 (I57567,I2683,I57499,I57593,);
DFFARX1 I_3228 (I524307,I2683,I57499,I57610,);
and I_3229 (I57618,I57610,I524310);
nor I_3230 (I57635,I57593,I57618);
DFFARX1 I_3231 (I57635,I2683,I57499,I57467,);
nand I_3232 (I57666,I57610,I524310);
nand I_3233 (I57683,I57533,I57666);
not I_3234 (I57479,I57683);
DFFARX1 I_3235 (I524304,I2683,I57499,I57723,);
DFFARX1 I_3236 (I57723,I2683,I57499,I57488,);
nand I_3237 (I57745,I524322,I524313);
and I_3238 (I57762,I57745,I524328);
DFFARX1 I_3239 (I57762,I2683,I57499,I57788,);
DFFARX1 I_3240 (I57788,I2683,I57499,I57805,);
not I_3241 (I57491,I57805);
not I_3242 (I57827,I57788);
nand I_3243 (I57476,I57827,I57666);
nor I_3244 (I57858,I524319,I524313);
not I_3245 (I57875,I57858);
nor I_3246 (I57892,I57827,I57875);
nor I_3247 (I57909,I57533,I57892);
DFFARX1 I_3248 (I57909,I2683,I57499,I57485,);
nor I_3249 (I57940,I57593,I57875);
nor I_3250 (I57473,I57788,I57940);
nor I_3251 (I57482,I57723,I57858);
nor I_3252 (I57470,I57593,I57858);
not I_3253 (I58026,I2690);
DFFARX1 I_3254 (I518536,I2683,I58026,I58052,);
not I_3255 (I58060,I58052);
nand I_3256 (I58077,I518527,I518545);
and I_3257 (I58094,I58077,I518524);
DFFARX1 I_3258 (I58094,I2683,I58026,I58120,);
DFFARX1 I_3259 (I518527,I2683,I58026,I58137,);
and I_3260 (I58145,I58137,I518530);
nor I_3261 (I58162,I58120,I58145);
DFFARX1 I_3262 (I58162,I2683,I58026,I57994,);
nand I_3263 (I58193,I58137,I518530);
nand I_3264 (I58210,I58060,I58193);
not I_3265 (I58006,I58210);
DFFARX1 I_3266 (I518524,I2683,I58026,I58250,);
DFFARX1 I_3267 (I58250,I2683,I58026,I58015,);
nand I_3268 (I58272,I518542,I518533);
and I_3269 (I58289,I58272,I518548);
DFFARX1 I_3270 (I58289,I2683,I58026,I58315,);
DFFARX1 I_3271 (I58315,I2683,I58026,I58332,);
not I_3272 (I58018,I58332);
not I_3273 (I58354,I58315);
nand I_3274 (I58003,I58354,I58193);
nor I_3275 (I58385,I518539,I518533);
not I_3276 (I58402,I58385);
nor I_3277 (I58419,I58354,I58402);
nor I_3278 (I58436,I58060,I58419);
DFFARX1 I_3279 (I58436,I2683,I58026,I58012,);
nor I_3280 (I58467,I58120,I58402);
nor I_3281 (I58000,I58315,I58467);
nor I_3282 (I58009,I58250,I58385);
nor I_3283 (I57997,I58120,I58385);
not I_3284 (I58553,I2690);
DFFARX1 I_3285 (I240652,I2683,I58553,I58579,);
not I_3286 (I58587,I58579);
nand I_3287 (I58604,I240634,I240649);
and I_3288 (I58621,I58604,I240625);
DFFARX1 I_3289 (I58621,I2683,I58553,I58647,);
DFFARX1 I_3290 (I240628,I2683,I58553,I58664,);
and I_3291 (I58672,I58664,I240643);
nor I_3292 (I58689,I58647,I58672);
DFFARX1 I_3293 (I58689,I2683,I58553,I58521,);
nand I_3294 (I58720,I58664,I240643);
nand I_3295 (I58737,I58587,I58720);
not I_3296 (I58533,I58737);
DFFARX1 I_3297 (I240646,I2683,I58553,I58777,);
DFFARX1 I_3298 (I58777,I2683,I58553,I58542,);
nand I_3299 (I58799,I240625,I240637);
and I_3300 (I58816,I58799,I240631);
DFFARX1 I_3301 (I58816,I2683,I58553,I58842,);
DFFARX1 I_3302 (I58842,I2683,I58553,I58859,);
not I_3303 (I58545,I58859);
not I_3304 (I58881,I58842);
nand I_3305 (I58530,I58881,I58720);
nor I_3306 (I58912,I240640,I240637);
not I_3307 (I58929,I58912);
nor I_3308 (I58946,I58881,I58929);
nor I_3309 (I58963,I58587,I58946);
DFFARX1 I_3310 (I58963,I2683,I58553,I58539,);
nor I_3311 (I58994,I58647,I58929);
nor I_3312 (I58527,I58842,I58994);
nor I_3313 (I58536,I58777,I58912);
nor I_3314 (I58524,I58647,I58912);
not I_3315 (I59080,I2690);
DFFARX1 I_3316 (I3898,I2683,I59080,I59106,);
not I_3317 (I59114,I59106);
nand I_3318 (I59131,I3883,I3883);
and I_3319 (I59148,I59131,I3904);
DFFARX1 I_3320 (I59148,I2683,I59080,I59174,);
DFFARX1 I_3321 (I3886,I2683,I59080,I59191,);
and I_3322 (I59199,I59191,I3895);
nor I_3323 (I59216,I59174,I59199);
DFFARX1 I_3324 (I59216,I2683,I59080,I59048,);
nand I_3325 (I59247,I59191,I3895);
nand I_3326 (I59264,I59114,I59247);
not I_3327 (I59060,I59264);
DFFARX1 I_3328 (I3889,I2683,I59080,I59304,);
DFFARX1 I_3329 (I59304,I2683,I59080,I59069,);
nand I_3330 (I59326,I3892,I3901);
and I_3331 (I59343,I59326,I3886);
DFFARX1 I_3332 (I59343,I2683,I59080,I59369,);
DFFARX1 I_3333 (I59369,I2683,I59080,I59386,);
not I_3334 (I59072,I59386);
not I_3335 (I59408,I59369);
nand I_3336 (I59057,I59408,I59247);
nor I_3337 (I59439,I3889,I3901);
not I_3338 (I59456,I59439);
nor I_3339 (I59473,I59408,I59456);
nor I_3340 (I59490,I59114,I59473);
DFFARX1 I_3341 (I59490,I2683,I59080,I59066,);
nor I_3342 (I59521,I59174,I59456);
nor I_3343 (I59054,I59369,I59521);
nor I_3344 (I59063,I59304,I59439);
nor I_3345 (I59051,I59174,I59439);
not I_3346 (I59607,I2690);
DFFARX1 I_3347 (I602924,I2683,I59607,I59633,);
not I_3348 (I59641,I59633);
nand I_3349 (I59658,I602915,I602933);
and I_3350 (I59675,I59658,I602912);
DFFARX1 I_3351 (I59675,I2683,I59607,I59701,);
DFFARX1 I_3352 (I602915,I2683,I59607,I59718,);
and I_3353 (I59726,I59718,I602918);
nor I_3354 (I59743,I59701,I59726);
DFFARX1 I_3355 (I59743,I2683,I59607,I59575,);
nand I_3356 (I59774,I59718,I602918);
nand I_3357 (I59791,I59641,I59774);
not I_3358 (I59587,I59791);
DFFARX1 I_3359 (I602912,I2683,I59607,I59831,);
DFFARX1 I_3360 (I59831,I2683,I59607,I59596,);
nand I_3361 (I59853,I602930,I602921);
and I_3362 (I59870,I59853,I602936);
DFFARX1 I_3363 (I59870,I2683,I59607,I59896,);
DFFARX1 I_3364 (I59896,I2683,I59607,I59913,);
not I_3365 (I59599,I59913);
not I_3366 (I59935,I59896);
nand I_3367 (I59584,I59935,I59774);
nor I_3368 (I59966,I602927,I602921);
not I_3369 (I59983,I59966);
nor I_3370 (I60000,I59935,I59983);
nor I_3371 (I60017,I59641,I60000);
DFFARX1 I_3372 (I60017,I2683,I59607,I59593,);
nor I_3373 (I60048,I59701,I59983);
nor I_3374 (I59581,I59896,I60048);
nor I_3375 (I59590,I59831,I59966);
nor I_3376 (I59578,I59701,I59966);
not I_3377 (I60134,I2690);
DFFARX1 I_3378 (I368772,I2683,I60134,I60160,);
not I_3379 (I60168,I60160);
nand I_3380 (I60185,I368766,I368757);
and I_3381 (I60202,I60185,I368778);
DFFARX1 I_3382 (I60202,I2683,I60134,I60228,);
DFFARX1 I_3383 (I368760,I2683,I60134,I60245,);
and I_3384 (I60253,I60245,I368754);
nor I_3385 (I60270,I60228,I60253);
DFFARX1 I_3386 (I60270,I2683,I60134,I60102,);
nand I_3387 (I60301,I60245,I368754);
nand I_3388 (I60318,I60168,I60301);
not I_3389 (I60114,I60318);
DFFARX1 I_3390 (I368754,I2683,I60134,I60358,);
DFFARX1 I_3391 (I60358,I2683,I60134,I60123,);
nand I_3392 (I60380,I368781,I368763);
and I_3393 (I60397,I60380,I368769);
DFFARX1 I_3394 (I60397,I2683,I60134,I60423,);
DFFARX1 I_3395 (I60423,I2683,I60134,I60440,);
not I_3396 (I60126,I60440);
not I_3397 (I60462,I60423);
nand I_3398 (I60111,I60462,I60301);
nor I_3399 (I60493,I368775,I368763);
not I_3400 (I60510,I60493);
nor I_3401 (I60527,I60462,I60510);
nor I_3402 (I60544,I60168,I60527);
DFFARX1 I_3403 (I60544,I2683,I60134,I60120,);
nor I_3404 (I60575,I60228,I60510);
nor I_3405 (I60108,I60423,I60575);
nor I_3406 (I60117,I60358,I60493);
nor I_3407 (I60105,I60228,I60493);
not I_3408 (I60661,I2690);
DFFARX1 I_3409 (I829936,I2683,I60661,I60687,);
not I_3410 (I60695,I60687);
nand I_3411 (I60712,I829951,I829930);
and I_3412 (I60729,I60712,I829933);
DFFARX1 I_3413 (I60729,I2683,I60661,I60755,);
DFFARX1 I_3414 (I829954,I2683,I60661,I60772,);
and I_3415 (I60780,I60772,I829933);
nor I_3416 (I60797,I60755,I60780);
DFFARX1 I_3417 (I60797,I2683,I60661,I60629,);
nand I_3418 (I60828,I60772,I829933);
nand I_3419 (I60845,I60695,I60828);
not I_3420 (I60641,I60845);
DFFARX1 I_3421 (I829930,I2683,I60661,I60885,);
DFFARX1 I_3422 (I60885,I2683,I60661,I60650,);
nand I_3423 (I60907,I829942,I829939);
and I_3424 (I60924,I60907,I829945);
DFFARX1 I_3425 (I60924,I2683,I60661,I60950,);
DFFARX1 I_3426 (I60950,I2683,I60661,I60967,);
not I_3427 (I60653,I60967);
not I_3428 (I60989,I60950);
nand I_3429 (I60638,I60989,I60828);
nor I_3430 (I61020,I829948,I829939);
not I_3431 (I61037,I61020);
nor I_3432 (I61054,I60989,I61037);
nor I_3433 (I61071,I60695,I61054);
DFFARX1 I_3434 (I61071,I2683,I60661,I60647,);
nor I_3435 (I61102,I60755,I61037);
nor I_3436 (I60635,I60950,I61102);
nor I_3437 (I60644,I60885,I61020);
nor I_3438 (I60632,I60755,I61020);
not I_3439 (I61188,I2690);
DFFARX1 I_3440 (I355172,I2683,I61188,I61214,);
not I_3441 (I61222,I61214);
nand I_3442 (I61239,I355166,I355157);
and I_3443 (I61256,I61239,I355178);
DFFARX1 I_3444 (I61256,I2683,I61188,I61282,);
DFFARX1 I_3445 (I355160,I2683,I61188,I61299,);
and I_3446 (I61307,I61299,I355154);
nor I_3447 (I61324,I61282,I61307);
DFFARX1 I_3448 (I61324,I2683,I61188,I61156,);
nand I_3449 (I61355,I61299,I355154);
nand I_3450 (I61372,I61222,I61355);
not I_3451 (I61168,I61372);
DFFARX1 I_3452 (I355154,I2683,I61188,I61412,);
DFFARX1 I_3453 (I61412,I2683,I61188,I61177,);
nand I_3454 (I61434,I355181,I355163);
and I_3455 (I61451,I61434,I355169);
DFFARX1 I_3456 (I61451,I2683,I61188,I61477,);
DFFARX1 I_3457 (I61477,I2683,I61188,I61494,);
not I_3458 (I61180,I61494);
not I_3459 (I61516,I61477);
nand I_3460 (I61165,I61516,I61355);
nor I_3461 (I61547,I355175,I355163);
not I_3462 (I61564,I61547);
nor I_3463 (I61581,I61516,I61564);
nor I_3464 (I61598,I61222,I61581);
DFFARX1 I_3465 (I61598,I2683,I61188,I61174,);
nor I_3466 (I61629,I61282,I61564);
nor I_3467 (I61162,I61477,I61629);
nor I_3468 (I61171,I61412,I61547);
nor I_3469 (I61159,I61282,I61547);
not I_3470 (I61715,I2690);
DFFARX1 I_3471 (I1964,I2683,I61715,I61741,);
not I_3472 (I61749,I61741);
nand I_3473 (I61766,I2284,I2340);
and I_3474 (I61783,I61766,I2212);
DFFARX1 I_3475 (I61783,I2683,I61715,I61809,);
DFFARX1 I_3476 (I1660,I2683,I61715,I61826,);
and I_3477 (I61834,I61826,I2388);
nor I_3478 (I61851,I61809,I61834);
DFFARX1 I_3479 (I61851,I2683,I61715,I61683,);
nand I_3480 (I61882,I61826,I2388);
nand I_3481 (I61899,I61749,I61882);
not I_3482 (I61695,I61899);
DFFARX1 I_3483 (I2516,I2683,I61715,I61939,);
DFFARX1 I_3484 (I61939,I2683,I61715,I61704,);
nand I_3485 (I61961,I2660,I2588);
and I_3486 (I61978,I61961,I2108);
DFFARX1 I_3487 (I61978,I2683,I61715,I62004,);
DFFARX1 I_3488 (I62004,I2683,I61715,I62021,);
not I_3489 (I61707,I62021);
not I_3490 (I62043,I62004);
nand I_3491 (I61692,I62043,I61882);
nor I_3492 (I62074,I2532,I2588);
not I_3493 (I62091,I62074);
nor I_3494 (I62108,I62043,I62091);
nor I_3495 (I62125,I61749,I62108);
DFFARX1 I_3496 (I62125,I2683,I61715,I61701,);
nor I_3497 (I62156,I61809,I62091);
nor I_3498 (I61689,I62004,I62156);
nor I_3499 (I61698,I61939,I62074);
nor I_3500 (I61686,I61809,I62074);
not I_3501 (I62242,I2690);
DFFARX1 I_3502 (I847276,I2683,I62242,I62268,);
not I_3503 (I62276,I62268);
nand I_3504 (I62293,I847291,I847270);
and I_3505 (I62310,I62293,I847273);
DFFARX1 I_3506 (I62310,I2683,I62242,I62336,);
DFFARX1 I_3507 (I847294,I2683,I62242,I62353,);
and I_3508 (I62361,I62353,I847273);
nor I_3509 (I62378,I62336,I62361);
DFFARX1 I_3510 (I62378,I2683,I62242,I62210,);
nand I_3511 (I62409,I62353,I847273);
nand I_3512 (I62426,I62276,I62409);
not I_3513 (I62222,I62426);
DFFARX1 I_3514 (I847270,I2683,I62242,I62466,);
DFFARX1 I_3515 (I62466,I2683,I62242,I62231,);
nand I_3516 (I62488,I847282,I847279);
and I_3517 (I62505,I62488,I847285);
DFFARX1 I_3518 (I62505,I2683,I62242,I62531,);
DFFARX1 I_3519 (I62531,I2683,I62242,I62548,);
not I_3520 (I62234,I62548);
not I_3521 (I62570,I62531);
nand I_3522 (I62219,I62570,I62409);
nor I_3523 (I62601,I847288,I847279);
not I_3524 (I62618,I62601);
nor I_3525 (I62635,I62570,I62618);
nor I_3526 (I62652,I62276,I62635);
DFFARX1 I_3527 (I62652,I2683,I62242,I62228,);
nor I_3528 (I62683,I62336,I62618);
nor I_3529 (I62216,I62531,I62683);
nor I_3530 (I62225,I62466,I62601);
nor I_3531 (I62213,I62336,I62601);
not I_3532 (I62769,I2690);
DFFARX1 I_3533 (I844964,I2683,I62769,I62795,);
not I_3534 (I62803,I62795);
nand I_3535 (I62820,I844979,I844958);
and I_3536 (I62837,I62820,I844961);
DFFARX1 I_3537 (I62837,I2683,I62769,I62863,);
DFFARX1 I_3538 (I844982,I2683,I62769,I62880,);
and I_3539 (I62888,I62880,I844961);
nor I_3540 (I62905,I62863,I62888);
DFFARX1 I_3541 (I62905,I2683,I62769,I62737,);
nand I_3542 (I62936,I62880,I844961);
nand I_3543 (I62953,I62803,I62936);
not I_3544 (I62749,I62953);
DFFARX1 I_3545 (I844958,I2683,I62769,I62993,);
DFFARX1 I_3546 (I62993,I2683,I62769,I62758,);
nand I_3547 (I63015,I844970,I844967);
and I_3548 (I63032,I63015,I844973);
DFFARX1 I_3549 (I63032,I2683,I62769,I63058,);
DFFARX1 I_3550 (I63058,I2683,I62769,I63075,);
not I_3551 (I62761,I63075);
not I_3552 (I63097,I63058);
nand I_3553 (I62746,I63097,I62936);
nor I_3554 (I63128,I844976,I844967);
not I_3555 (I63145,I63128);
nor I_3556 (I63162,I63097,I63145);
nor I_3557 (I63179,I62803,I63162);
DFFARX1 I_3558 (I63179,I2683,I62769,I62755,);
nor I_3559 (I63210,I62863,I63145);
nor I_3560 (I62743,I63058,I63210);
nor I_3561 (I62752,I62993,I63128);
nor I_3562 (I62740,I62863,I63128);
not I_3563 (I63296,I2690);
DFFARX1 I_3564 (I31141,I2683,I63296,I63322,);
not I_3565 (I63330,I63322);
nand I_3566 (I63347,I31129,I31135);
and I_3567 (I63364,I63347,I31138);
DFFARX1 I_3568 (I63364,I2683,I63296,I63390,);
DFFARX1 I_3569 (I31120,I2683,I63296,I63407,);
and I_3570 (I63415,I63407,I31126);
nor I_3571 (I63432,I63390,I63415);
DFFARX1 I_3572 (I63432,I2683,I63296,I63264,);
nand I_3573 (I63463,I63407,I31126);
nand I_3574 (I63480,I63330,I63463);
not I_3575 (I63276,I63480);
DFFARX1 I_3576 (I31120,I2683,I63296,I63520,);
DFFARX1 I_3577 (I63520,I2683,I63296,I63285,);
nand I_3578 (I63542,I31123,I31117);
and I_3579 (I63559,I63542,I31132);
DFFARX1 I_3580 (I63559,I2683,I63296,I63585,);
DFFARX1 I_3581 (I63585,I2683,I63296,I63602,);
not I_3582 (I63288,I63602);
not I_3583 (I63624,I63585);
nand I_3584 (I63273,I63624,I63463);
nor I_3585 (I63655,I31117,I31117);
not I_3586 (I63672,I63655);
nor I_3587 (I63689,I63624,I63672);
nor I_3588 (I63706,I63330,I63689);
DFFARX1 I_3589 (I63706,I2683,I63296,I63282,);
nor I_3590 (I63737,I63390,I63672);
nor I_3591 (I63270,I63585,I63737);
nor I_3592 (I63279,I63520,I63655);
nor I_3593 (I63267,I63390,I63655);
not I_3594 (I63823,I2690);
DFFARX1 I_3595 (I465935,I2683,I63823,I63849,);
not I_3596 (I63857,I63849);
nand I_3597 (I63874,I465947,I465932);
and I_3598 (I63891,I63874,I465926);
DFFARX1 I_3599 (I63891,I2683,I63823,I63917,);
DFFARX1 I_3600 (I465941,I2683,I63823,I63934,);
and I_3601 (I63942,I63934,I465929);
nor I_3602 (I63959,I63917,I63942);
DFFARX1 I_3603 (I63959,I2683,I63823,I63791,);
nand I_3604 (I63990,I63934,I465929);
nand I_3605 (I64007,I63857,I63990);
not I_3606 (I63803,I64007);
DFFARX1 I_3607 (I465938,I2683,I63823,I64047,);
DFFARX1 I_3608 (I64047,I2683,I63823,I63812,);
nand I_3609 (I64069,I465944,I465950);
and I_3610 (I64086,I64069,I465926);
DFFARX1 I_3611 (I64086,I2683,I63823,I64112,);
DFFARX1 I_3612 (I64112,I2683,I63823,I64129,);
not I_3613 (I63815,I64129);
not I_3614 (I64151,I64112);
nand I_3615 (I63800,I64151,I63990);
nor I_3616 (I64182,I465929,I465950);
not I_3617 (I64199,I64182);
nor I_3618 (I64216,I64151,I64199);
nor I_3619 (I64233,I63857,I64216);
DFFARX1 I_3620 (I64233,I2683,I63823,I63809,);
nor I_3621 (I64264,I63917,I64199);
nor I_3622 (I63797,I64112,I64264);
nor I_3623 (I63806,I64047,I64182);
nor I_3624 (I63794,I63917,I64182);
not I_3625 (I64350,I2690);
DFFARX1 I_3626 (I244341,I2683,I64350,I64376,);
not I_3627 (I64384,I64376);
nand I_3628 (I64401,I244323,I244338);
and I_3629 (I64418,I64401,I244314);
DFFARX1 I_3630 (I64418,I2683,I64350,I64444,);
DFFARX1 I_3631 (I244317,I2683,I64350,I64461,);
and I_3632 (I64469,I64461,I244332);
nor I_3633 (I64486,I64444,I64469);
DFFARX1 I_3634 (I64486,I2683,I64350,I64318,);
nand I_3635 (I64517,I64461,I244332);
nand I_3636 (I64534,I64384,I64517);
not I_3637 (I64330,I64534);
DFFARX1 I_3638 (I244335,I2683,I64350,I64574,);
DFFARX1 I_3639 (I64574,I2683,I64350,I64339,);
nand I_3640 (I64596,I244314,I244326);
and I_3641 (I64613,I64596,I244320);
DFFARX1 I_3642 (I64613,I2683,I64350,I64639,);
DFFARX1 I_3643 (I64639,I2683,I64350,I64656,);
not I_3644 (I64342,I64656);
not I_3645 (I64678,I64639);
nand I_3646 (I64327,I64678,I64517);
nor I_3647 (I64709,I244329,I244326);
not I_3648 (I64726,I64709);
nor I_3649 (I64743,I64678,I64726);
nor I_3650 (I64760,I64384,I64743);
DFFARX1 I_3651 (I64760,I2683,I64350,I64336,);
nor I_3652 (I64791,I64444,I64726);
nor I_3653 (I64324,I64639,I64791);
nor I_3654 (I64333,I64574,I64709);
nor I_3655 (I64321,I64444,I64709);
not I_3656 (I64877,I2690);
DFFARX1 I_3657 (I605236,I2683,I64877,I64903,);
not I_3658 (I64911,I64903);
nand I_3659 (I64928,I605227,I605245);
and I_3660 (I64945,I64928,I605224);
DFFARX1 I_3661 (I64945,I2683,I64877,I64971,);
DFFARX1 I_3662 (I605227,I2683,I64877,I64988,);
and I_3663 (I64996,I64988,I605230);
nor I_3664 (I65013,I64971,I64996);
DFFARX1 I_3665 (I65013,I2683,I64877,I64845,);
nand I_3666 (I65044,I64988,I605230);
nand I_3667 (I65061,I64911,I65044);
not I_3668 (I64857,I65061);
DFFARX1 I_3669 (I605224,I2683,I64877,I65101,);
DFFARX1 I_3670 (I65101,I2683,I64877,I64866,);
nand I_3671 (I65123,I605242,I605233);
and I_3672 (I65140,I65123,I605248);
DFFARX1 I_3673 (I65140,I2683,I64877,I65166,);
DFFARX1 I_3674 (I65166,I2683,I64877,I65183,);
not I_3675 (I64869,I65183);
not I_3676 (I65205,I65166);
nand I_3677 (I64854,I65205,I65044);
nor I_3678 (I65236,I605239,I605233);
not I_3679 (I65253,I65236);
nor I_3680 (I65270,I65205,I65253);
nor I_3681 (I65287,I64911,I65270);
DFFARX1 I_3682 (I65287,I2683,I64877,I64863,);
nor I_3683 (I65318,I64971,I65253);
nor I_3684 (I64851,I65166,I65318);
nor I_3685 (I64860,I65101,I65236);
nor I_3686 (I64848,I64971,I65236);
not I_3687 (I65404,I2690);
DFFARX1 I_3688 (I438191,I2683,I65404,I65430,);
not I_3689 (I65438,I65430);
nand I_3690 (I65455,I438203,I438188);
and I_3691 (I65472,I65455,I438182);
DFFARX1 I_3692 (I65472,I2683,I65404,I65498,);
DFFARX1 I_3693 (I438197,I2683,I65404,I65515,);
and I_3694 (I65523,I65515,I438185);
nor I_3695 (I65540,I65498,I65523);
DFFARX1 I_3696 (I65540,I2683,I65404,I65372,);
nand I_3697 (I65571,I65515,I438185);
nand I_3698 (I65588,I65438,I65571);
not I_3699 (I65384,I65588);
DFFARX1 I_3700 (I438194,I2683,I65404,I65628,);
DFFARX1 I_3701 (I65628,I2683,I65404,I65393,);
nand I_3702 (I65650,I438200,I438206);
and I_3703 (I65667,I65650,I438182);
DFFARX1 I_3704 (I65667,I2683,I65404,I65693,);
DFFARX1 I_3705 (I65693,I2683,I65404,I65710,);
not I_3706 (I65396,I65710);
not I_3707 (I65732,I65693);
nand I_3708 (I65381,I65732,I65571);
nor I_3709 (I65763,I438185,I438206);
not I_3710 (I65780,I65763);
nor I_3711 (I65797,I65732,I65780);
nor I_3712 (I65814,I65438,I65797);
DFFARX1 I_3713 (I65814,I2683,I65404,I65390,);
nor I_3714 (I65845,I65498,I65780);
nor I_3715 (I65378,I65693,I65845);
nor I_3716 (I65387,I65628,I65763);
nor I_3717 (I65375,I65498,I65763);
not I_3718 (I65931,I2690);
DFFARX1 I_3719 (I394920,I2683,I65931,I65957,);
not I_3720 (I65965,I65957);
nand I_3721 (I65982,I394941,I394935);
and I_3722 (I65999,I65982,I394917);
DFFARX1 I_3723 (I65999,I2683,I65931,I66025,);
DFFARX1 I_3724 (I394920,I2683,I65931,I66042,);
and I_3725 (I66050,I66042,I394929);
nor I_3726 (I66067,I66025,I66050);
DFFARX1 I_3727 (I66067,I2683,I65931,I65899,);
nand I_3728 (I66098,I66042,I394929);
nand I_3729 (I66115,I65965,I66098);
not I_3730 (I65911,I66115);
DFFARX1 I_3731 (I394926,I2683,I65931,I66155,);
DFFARX1 I_3732 (I66155,I2683,I65931,I65920,);
nand I_3733 (I66177,I394932,I394923);
and I_3734 (I66194,I66177,I394917);
DFFARX1 I_3735 (I66194,I2683,I65931,I66220,);
DFFARX1 I_3736 (I66220,I2683,I65931,I66237,);
not I_3737 (I65923,I66237);
not I_3738 (I66259,I66220);
nand I_3739 (I65908,I66259,I66098);
nor I_3740 (I66290,I394938,I394923);
not I_3741 (I66307,I66290);
nor I_3742 (I66324,I66259,I66307);
nor I_3743 (I66341,I65965,I66324);
DFFARX1 I_3744 (I66341,I2683,I65931,I65917,);
nor I_3745 (I66372,I66025,I66307);
nor I_3746 (I65905,I66220,I66372);
nor I_3747 (I65914,I66155,I66290);
nor I_3748 (I65902,I66025,I66290);
not I_3749 (I66458,I2690);
DFFARX1 I_3750 (I586162,I2683,I66458,I66484,);
not I_3751 (I66492,I66484);
nand I_3752 (I66509,I586153,I586171);
and I_3753 (I66526,I66509,I586150);
DFFARX1 I_3754 (I66526,I2683,I66458,I66552,);
DFFARX1 I_3755 (I586153,I2683,I66458,I66569,);
and I_3756 (I66577,I66569,I586156);
nor I_3757 (I66594,I66552,I66577);
DFFARX1 I_3758 (I66594,I2683,I66458,I66426,);
nand I_3759 (I66625,I66569,I586156);
nand I_3760 (I66642,I66492,I66625);
not I_3761 (I66438,I66642);
DFFARX1 I_3762 (I586150,I2683,I66458,I66682,);
DFFARX1 I_3763 (I66682,I2683,I66458,I66447,);
nand I_3764 (I66704,I586168,I586159);
and I_3765 (I66721,I66704,I586174);
DFFARX1 I_3766 (I66721,I2683,I66458,I66747,);
DFFARX1 I_3767 (I66747,I2683,I66458,I66764,);
not I_3768 (I66450,I66764);
not I_3769 (I66786,I66747);
nand I_3770 (I66435,I66786,I66625);
nor I_3771 (I66817,I586165,I586159);
not I_3772 (I66834,I66817);
nor I_3773 (I66851,I66786,I66834);
nor I_3774 (I66868,I66492,I66851);
DFFARX1 I_3775 (I66868,I2683,I66458,I66444,);
nor I_3776 (I66899,I66552,I66834);
nor I_3777 (I66432,I66747,I66899);
nor I_3778 (I66441,I66682,I66817);
nor I_3779 (I66429,I66552,I66817);
not I_3780 (I66985,I2690);
DFFARX1 I_3781 (I1043581,I2683,I66985,I67011,);
not I_3782 (I67019,I67011);
nand I_3783 (I67036,I1043575,I1043596);
and I_3784 (I67053,I67036,I1043572);
DFFARX1 I_3785 (I67053,I2683,I66985,I67079,);
DFFARX1 I_3786 (I1043593,I2683,I66985,I67096,);
and I_3787 (I67104,I67096,I1043590);
nor I_3788 (I67121,I67079,I67104);
DFFARX1 I_3789 (I67121,I2683,I66985,I66953,);
nand I_3790 (I67152,I67096,I1043590);
nand I_3791 (I67169,I67019,I67152);
not I_3792 (I66965,I67169);
DFFARX1 I_3793 (I1043578,I2683,I66985,I67209,);
DFFARX1 I_3794 (I67209,I2683,I66985,I66974,);
nand I_3795 (I67231,I1043587,I1043584);
and I_3796 (I67248,I67231,I1043569);
DFFARX1 I_3797 (I67248,I2683,I66985,I67274,);
DFFARX1 I_3798 (I67274,I2683,I66985,I67291,);
not I_3799 (I66977,I67291);
not I_3800 (I67313,I67274);
nand I_3801 (I66962,I67313,I67152);
nor I_3802 (I67344,I1043569,I1043584);
not I_3803 (I67361,I67344);
nor I_3804 (I67378,I67313,I67361);
nor I_3805 (I67395,I67019,I67378);
DFFARX1 I_3806 (I67395,I2683,I66985,I66971,);
nor I_3807 (I67426,I67079,I67361);
nor I_3808 (I66959,I67274,I67426);
nor I_3809 (I66968,I67209,I67344);
nor I_3810 (I66956,I67079,I67344);
not I_3811 (I67512,I2690);
DFFARX1 I_3812 (I406225,I2683,I67512,I67538,);
not I_3813 (I67546,I67538);
nand I_3814 (I67563,I406246,I406240);
and I_3815 (I67580,I67563,I406222);
DFFARX1 I_3816 (I67580,I2683,I67512,I67606,);
DFFARX1 I_3817 (I406225,I2683,I67512,I67623,);
and I_3818 (I67631,I67623,I406234);
nor I_3819 (I67648,I67606,I67631);
DFFARX1 I_3820 (I67648,I2683,I67512,I67480,);
nand I_3821 (I67679,I67623,I406234);
nand I_3822 (I67696,I67546,I67679);
not I_3823 (I67492,I67696);
DFFARX1 I_3824 (I406231,I2683,I67512,I67736,);
DFFARX1 I_3825 (I67736,I2683,I67512,I67501,);
nand I_3826 (I67758,I406237,I406228);
and I_3827 (I67775,I67758,I406222);
DFFARX1 I_3828 (I67775,I2683,I67512,I67801,);
DFFARX1 I_3829 (I67801,I2683,I67512,I67818,);
not I_3830 (I67504,I67818);
not I_3831 (I67840,I67801);
nand I_3832 (I67489,I67840,I67679);
nor I_3833 (I67871,I406243,I406228);
not I_3834 (I67888,I67871);
nor I_3835 (I67905,I67840,I67888);
nor I_3836 (I67922,I67546,I67905);
DFFARX1 I_3837 (I67922,I2683,I67512,I67498,);
nor I_3838 (I67953,I67606,I67888);
nor I_3839 (I67486,I67801,I67953);
nor I_3840 (I67495,I67736,I67871);
nor I_3841 (I67483,I67606,I67871);
not I_3842 (I68039,I2690);
DFFARX1 I_3843 (I919526,I2683,I68039,I68065,);
not I_3844 (I68073,I68065);
nand I_3845 (I68090,I919541,I919520);
and I_3846 (I68107,I68090,I919523);
DFFARX1 I_3847 (I68107,I2683,I68039,I68133,);
DFFARX1 I_3848 (I919544,I2683,I68039,I68150,);
and I_3849 (I68158,I68150,I919523);
nor I_3850 (I68175,I68133,I68158);
DFFARX1 I_3851 (I68175,I2683,I68039,I68007,);
nand I_3852 (I68206,I68150,I919523);
nand I_3853 (I68223,I68073,I68206);
not I_3854 (I68019,I68223);
DFFARX1 I_3855 (I919520,I2683,I68039,I68263,);
DFFARX1 I_3856 (I68263,I2683,I68039,I68028,);
nand I_3857 (I68285,I919532,I919529);
and I_3858 (I68302,I68285,I919535);
DFFARX1 I_3859 (I68302,I2683,I68039,I68328,);
DFFARX1 I_3860 (I68328,I2683,I68039,I68345,);
not I_3861 (I68031,I68345);
not I_3862 (I68367,I68328);
nand I_3863 (I68016,I68367,I68206);
nor I_3864 (I68398,I919538,I919529);
not I_3865 (I68415,I68398);
nor I_3866 (I68432,I68367,I68415);
nor I_3867 (I68449,I68073,I68432);
DFFARX1 I_3868 (I68449,I2683,I68039,I68025,);
nor I_3869 (I68480,I68133,I68415);
nor I_3870 (I68013,I68328,I68480);
nor I_3871 (I68022,I68263,I68398);
nor I_3872 (I68010,I68133,I68398);
not I_3873 (I68566,I2690);
DFFARX1 I_3874 (I958660,I2683,I68566,I68592,);
not I_3875 (I68600,I68592);
nand I_3876 (I68617,I958654,I958675);
and I_3877 (I68634,I68617,I958666);
DFFARX1 I_3878 (I68634,I2683,I68566,I68660,);
DFFARX1 I_3879 (I958657,I2683,I68566,I68677,);
and I_3880 (I68685,I68677,I958669);
nor I_3881 (I68702,I68660,I68685);
DFFARX1 I_3882 (I68702,I2683,I68566,I68534,);
nand I_3883 (I68733,I68677,I958669);
nand I_3884 (I68750,I68600,I68733);
not I_3885 (I68546,I68750);
DFFARX1 I_3886 (I958657,I2683,I68566,I68790,);
DFFARX1 I_3887 (I68790,I2683,I68566,I68555,);
nand I_3888 (I68812,I958678,I958663);
and I_3889 (I68829,I68812,I958654);
DFFARX1 I_3890 (I68829,I2683,I68566,I68855,);
DFFARX1 I_3891 (I68855,I2683,I68566,I68872,);
not I_3892 (I68558,I68872);
not I_3893 (I68894,I68855);
nand I_3894 (I68543,I68894,I68733);
nor I_3895 (I68925,I958672,I958663);
not I_3896 (I68942,I68925);
nor I_3897 (I68959,I68894,I68942);
nor I_3898 (I68976,I68600,I68959);
DFFARX1 I_3899 (I68976,I2683,I68566,I68552,);
nor I_3900 (I69007,I68660,I68942);
nor I_3901 (I68540,I68855,I69007);
nor I_3902 (I68549,I68790,I68925);
nor I_3903 (I68537,I68660,I68925);
not I_3904 (I69093,I2690);
DFFARX1 I_3905 (I797905,I2683,I69093,I69119,);
not I_3906 (I69127,I69119);
nand I_3907 (I69144,I797902,I797908);
and I_3908 (I69161,I69144,I797905);
DFFARX1 I_3909 (I69161,I2683,I69093,I69187,);
DFFARX1 I_3910 (I797908,I2683,I69093,I69204,);
and I_3911 (I69212,I69204,I797902);
nor I_3912 (I69229,I69187,I69212);
DFFARX1 I_3913 (I69229,I2683,I69093,I69061,);
nand I_3914 (I69260,I69204,I797902);
nand I_3915 (I69277,I69127,I69260);
not I_3916 (I69073,I69277);
DFFARX1 I_3917 (I797911,I2683,I69093,I69317,);
DFFARX1 I_3918 (I69317,I2683,I69093,I69082,);
nand I_3919 (I69339,I797914,I797923);
and I_3920 (I69356,I69339,I797917);
DFFARX1 I_3921 (I69356,I2683,I69093,I69382,);
DFFARX1 I_3922 (I69382,I2683,I69093,I69399,);
not I_3923 (I69085,I69399);
not I_3924 (I69421,I69382);
nand I_3925 (I69070,I69421,I69260);
nor I_3926 (I69452,I797920,I797923);
not I_3927 (I69469,I69452);
nor I_3928 (I69486,I69421,I69469);
nor I_3929 (I69503,I69127,I69486);
DFFARX1 I_3930 (I69503,I2683,I69093,I69079,);
nor I_3931 (I69534,I69187,I69469);
nor I_3932 (I69067,I69382,I69534);
nor I_3933 (I69076,I69317,I69452);
nor I_3934 (I69064,I69187,I69452);
not I_3935 (I69620,I2690);
DFFARX1 I_3936 (I1032871,I2683,I69620,I69646,);
not I_3937 (I69654,I69646);
nand I_3938 (I69671,I1032865,I1032886);
and I_3939 (I69688,I69671,I1032862);
DFFARX1 I_3940 (I69688,I2683,I69620,I69714,);
DFFARX1 I_3941 (I1032883,I2683,I69620,I69731,);
and I_3942 (I69739,I69731,I1032880);
nor I_3943 (I69756,I69714,I69739);
DFFARX1 I_3944 (I69756,I2683,I69620,I69588,);
nand I_3945 (I69787,I69731,I1032880);
nand I_3946 (I69804,I69654,I69787);
not I_3947 (I69600,I69804);
DFFARX1 I_3948 (I1032868,I2683,I69620,I69844,);
DFFARX1 I_3949 (I69844,I2683,I69620,I69609,);
nand I_3950 (I69866,I1032877,I1032874);
and I_3951 (I69883,I69866,I1032859);
DFFARX1 I_3952 (I69883,I2683,I69620,I69909,);
DFFARX1 I_3953 (I69909,I2683,I69620,I69926,);
not I_3954 (I69612,I69926);
not I_3955 (I69948,I69909);
nand I_3956 (I69597,I69948,I69787);
nor I_3957 (I69979,I1032859,I1032874);
not I_3958 (I69996,I69979);
nor I_3959 (I70013,I69948,I69996);
nor I_3960 (I70030,I69654,I70013);
DFFARX1 I_3961 (I70030,I2683,I69620,I69606,);
nor I_3962 (I70061,I69714,I69996);
nor I_3963 (I69594,I69909,I70061);
nor I_3964 (I69603,I69844,I69979);
nor I_3965 (I69591,I69714,I69979);
not I_3966 (I70147,I2690);
DFFARX1 I_3967 (I1000155,I2683,I70147,I70173,);
not I_3968 (I70181,I70173);
nand I_3969 (I70198,I1000158,I1000152);
and I_3970 (I70215,I70198,I1000149);
DFFARX1 I_3971 (I70215,I2683,I70147,I70241,);
DFFARX1 I_3972 (I1000134,I2683,I70147,I70258,);
and I_3973 (I70266,I70258,I1000143);
nor I_3974 (I70283,I70241,I70266);
DFFARX1 I_3975 (I70283,I2683,I70147,I70115,);
nand I_3976 (I70314,I70258,I1000143);
nand I_3977 (I70331,I70181,I70314);
not I_3978 (I70127,I70331);
DFFARX1 I_3979 (I1000134,I2683,I70147,I70371,);
DFFARX1 I_3980 (I70371,I2683,I70147,I70136,);
nand I_3981 (I70393,I1000137,I1000140);
and I_3982 (I70410,I70393,I1000146);
DFFARX1 I_3983 (I70410,I2683,I70147,I70436,);
DFFARX1 I_3984 (I70436,I2683,I70147,I70453,);
not I_3985 (I70139,I70453);
not I_3986 (I70475,I70436);
nand I_3987 (I70124,I70475,I70314);
nor I_3988 (I70506,I1000137,I1000140);
not I_3989 (I70523,I70506);
nor I_3990 (I70540,I70475,I70523);
nor I_3991 (I70557,I70181,I70540);
DFFARX1 I_3992 (I70557,I2683,I70147,I70133,);
nor I_3993 (I70588,I70241,I70523);
nor I_3994 (I70121,I70436,I70588);
nor I_3995 (I70130,I70371,I70506);
nor I_3996 (I70118,I70241,I70506);
not I_3997 (I70674,I2690);
DFFARX1 I_3998 (I348644,I2683,I70674,I70700,);
not I_3999 (I70708,I70700);
nand I_4000 (I70725,I348638,I348629);
and I_4001 (I70742,I70725,I348650);
DFFARX1 I_4002 (I70742,I2683,I70674,I70768,);
DFFARX1 I_4003 (I348632,I2683,I70674,I70785,);
and I_4004 (I70793,I70785,I348626);
nor I_4005 (I70810,I70768,I70793);
DFFARX1 I_4006 (I70810,I2683,I70674,I70642,);
nand I_4007 (I70841,I70785,I348626);
nand I_4008 (I70858,I70708,I70841);
not I_4009 (I70654,I70858);
DFFARX1 I_4010 (I348626,I2683,I70674,I70898,);
DFFARX1 I_4011 (I70898,I2683,I70674,I70663,);
nand I_4012 (I70920,I348653,I348635);
and I_4013 (I70937,I70920,I348641);
DFFARX1 I_4014 (I70937,I2683,I70674,I70963,);
DFFARX1 I_4015 (I70963,I2683,I70674,I70980,);
not I_4016 (I70666,I70980);
not I_4017 (I71002,I70963);
nand I_4018 (I70651,I71002,I70841);
nor I_4019 (I71033,I348647,I348635);
not I_4020 (I71050,I71033);
nor I_4021 (I71067,I71002,I71050);
nor I_4022 (I71084,I70708,I71067);
DFFARX1 I_4023 (I71084,I2683,I70674,I70660,);
nor I_4024 (I71115,I70768,I71050);
nor I_4025 (I70648,I70963,I71115);
nor I_4026 (I70657,I70898,I71033);
nor I_4027 (I70645,I70768,I71033);
not I_4028 (I71201,I2690);
DFFARX1 I_4029 (I809125,I2683,I71201,I71227,);
not I_4030 (I71235,I71227);
nand I_4031 (I71252,I809122,I809128);
and I_4032 (I71269,I71252,I809125);
DFFARX1 I_4033 (I71269,I2683,I71201,I71295,);
DFFARX1 I_4034 (I809128,I2683,I71201,I71312,);
and I_4035 (I71320,I71312,I809122);
nor I_4036 (I71337,I71295,I71320);
DFFARX1 I_4037 (I71337,I2683,I71201,I71169,);
nand I_4038 (I71368,I71312,I809122);
nand I_4039 (I71385,I71235,I71368);
not I_4040 (I71181,I71385);
DFFARX1 I_4041 (I809131,I2683,I71201,I71425,);
DFFARX1 I_4042 (I71425,I2683,I71201,I71190,);
nand I_4043 (I71447,I809134,I809143);
and I_4044 (I71464,I71447,I809137);
DFFARX1 I_4045 (I71464,I2683,I71201,I71490,);
DFFARX1 I_4046 (I71490,I2683,I71201,I71507,);
not I_4047 (I71193,I71507);
not I_4048 (I71529,I71490);
nand I_4049 (I71178,I71529,I71368);
nor I_4050 (I71560,I809140,I809143);
not I_4051 (I71577,I71560);
nor I_4052 (I71594,I71529,I71577);
nor I_4053 (I71611,I71235,I71594);
DFFARX1 I_4054 (I71611,I2683,I71201,I71187,);
nor I_4055 (I71642,I71295,I71577);
nor I_4056 (I71175,I71490,I71642);
nor I_4057 (I71184,I71425,I71560);
nor I_4058 (I71172,I71295,I71560);
not I_4059 (I71728,I2690);
DFFARX1 I_4060 (I139062,I2683,I71728,I71754,);
not I_4061 (I71762,I71754);
nand I_4062 (I71779,I139056,I139050);
and I_4063 (I71796,I71779,I139071);
DFFARX1 I_4064 (I71796,I2683,I71728,I71822,);
DFFARX1 I_4065 (I139068,I2683,I71728,I71839,);
and I_4066 (I71847,I71839,I139065);
nor I_4067 (I71864,I71822,I71847);
DFFARX1 I_4068 (I71864,I2683,I71728,I71696,);
nand I_4069 (I71895,I71839,I139065);
nand I_4070 (I71912,I71762,I71895);
not I_4071 (I71708,I71912);
DFFARX1 I_4072 (I139050,I2683,I71728,I71952,);
DFFARX1 I_4073 (I71952,I2683,I71728,I71717,);
nand I_4074 (I71974,I139053,I139053);
and I_4075 (I71991,I71974,I139074);
DFFARX1 I_4076 (I71991,I2683,I71728,I72017,);
DFFARX1 I_4077 (I72017,I2683,I71728,I72034,);
not I_4078 (I71720,I72034);
not I_4079 (I72056,I72017);
nand I_4080 (I71705,I72056,I71895);
nor I_4081 (I72087,I139059,I139053);
not I_4082 (I72104,I72087);
nor I_4083 (I72121,I72056,I72104);
nor I_4084 (I72138,I71762,I72121);
DFFARX1 I_4085 (I72138,I2683,I71728,I71714,);
nor I_4086 (I72169,I71822,I72104);
nor I_4087 (I71702,I72017,I72169);
nor I_4088 (I71711,I71952,I72087);
nor I_4089 (I71699,I71822,I72087);
not I_4090 (I72255,I2690);
DFFARX1 I_4091 (I1001889,I2683,I72255,I72281,);
not I_4092 (I72289,I72281);
nand I_4093 (I72306,I1001892,I1001886);
and I_4094 (I72323,I72306,I1001883);
DFFARX1 I_4095 (I72323,I2683,I72255,I72349,);
DFFARX1 I_4096 (I1001868,I2683,I72255,I72366,);
and I_4097 (I72374,I72366,I1001877);
nor I_4098 (I72391,I72349,I72374);
DFFARX1 I_4099 (I72391,I2683,I72255,I72223,);
nand I_4100 (I72422,I72366,I1001877);
nand I_4101 (I72439,I72289,I72422);
not I_4102 (I72235,I72439);
DFFARX1 I_4103 (I1001868,I2683,I72255,I72479,);
DFFARX1 I_4104 (I72479,I2683,I72255,I72244,);
nand I_4105 (I72501,I1001871,I1001874);
and I_4106 (I72518,I72501,I1001880);
DFFARX1 I_4107 (I72518,I2683,I72255,I72544,);
DFFARX1 I_4108 (I72544,I2683,I72255,I72561,);
not I_4109 (I72247,I72561);
not I_4110 (I72583,I72544);
nand I_4111 (I72232,I72583,I72422);
nor I_4112 (I72614,I1001871,I1001874);
not I_4113 (I72631,I72614);
nor I_4114 (I72648,I72583,I72631);
nor I_4115 (I72665,I72289,I72648);
DFFARX1 I_4116 (I72665,I2683,I72255,I72241,);
nor I_4117 (I72696,I72349,I72631);
nor I_4118 (I72229,I72544,I72696);
nor I_4119 (I72238,I72479,I72614);
nor I_4120 (I72226,I72349,I72614);
not I_4121 (I72782,I2690);
DFFARX1 I_4122 (I283866,I2683,I72782,I72808,);
not I_4123 (I72816,I72808);
nand I_4124 (I72833,I283848,I283863);
and I_4125 (I72850,I72833,I283839);
DFFARX1 I_4126 (I72850,I2683,I72782,I72876,);
DFFARX1 I_4127 (I283842,I2683,I72782,I72893,);
and I_4128 (I72901,I72893,I283857);
nor I_4129 (I72918,I72876,I72901);
DFFARX1 I_4130 (I72918,I2683,I72782,I72750,);
nand I_4131 (I72949,I72893,I283857);
nand I_4132 (I72966,I72816,I72949);
not I_4133 (I72762,I72966);
DFFARX1 I_4134 (I283860,I2683,I72782,I73006,);
DFFARX1 I_4135 (I73006,I2683,I72782,I72771,);
nand I_4136 (I73028,I283839,I283851);
and I_4137 (I73045,I73028,I283845);
DFFARX1 I_4138 (I73045,I2683,I72782,I73071,);
DFFARX1 I_4139 (I73071,I2683,I72782,I73088,);
not I_4140 (I72774,I73088);
not I_4141 (I73110,I73071);
nand I_4142 (I72759,I73110,I72949);
nor I_4143 (I73141,I283854,I283851);
not I_4144 (I73158,I73141);
nor I_4145 (I73175,I73110,I73158);
nor I_4146 (I73192,I72816,I73175);
DFFARX1 I_4147 (I73192,I2683,I72782,I72768,);
nor I_4148 (I73223,I72876,I73158);
nor I_4149 (I72756,I73071,I73223);
nor I_4150 (I72765,I73006,I73141);
nor I_4151 (I72753,I72876,I73141);
not I_4152 (I73309,I2690);
DFFARX1 I_4153 (I703204,I2683,I73309,I73335,);
not I_4154 (I73343,I73335);
nand I_4155 (I73360,I703222,I703216);
and I_4156 (I73377,I73360,I703195);
DFFARX1 I_4157 (I73377,I2683,I73309,I73403,);
DFFARX1 I_4158 (I703213,I2683,I73309,I73420,);
and I_4159 (I73428,I73420,I703198);
nor I_4160 (I73445,I73403,I73428);
DFFARX1 I_4161 (I73445,I2683,I73309,I73277,);
nand I_4162 (I73476,I73420,I703198);
nand I_4163 (I73493,I73343,I73476);
not I_4164 (I73289,I73493);
DFFARX1 I_4165 (I703210,I2683,I73309,I73533,);
DFFARX1 I_4166 (I73533,I2683,I73309,I73298,);
nand I_4167 (I73555,I703219,I703207);
and I_4168 (I73572,I73555,I703201);
DFFARX1 I_4169 (I73572,I2683,I73309,I73598,);
DFFARX1 I_4170 (I73598,I2683,I73309,I73615,);
not I_4171 (I73301,I73615);
not I_4172 (I73637,I73598);
nand I_4173 (I73286,I73637,I73476);
nor I_4174 (I73668,I703195,I703207);
not I_4175 (I73685,I73668);
nor I_4176 (I73702,I73637,I73685);
nor I_4177 (I73719,I73343,I73702);
DFFARX1 I_4178 (I73719,I2683,I73309,I73295,);
nor I_4179 (I73750,I73403,I73685);
nor I_4180 (I73283,I73598,I73750);
nor I_4181 (I73292,I73533,I73668);
nor I_4182 (I73280,I73403,I73668);
not I_4183 (I73836,I2690);
DFFARX1 I_4184 (I1027674,I2683,I73836,I73862,);
not I_4185 (I73870,I73862);
nand I_4186 (I73887,I1027680,I1027698);
and I_4187 (I73904,I73887,I1027695);
DFFARX1 I_4188 (I73904,I2683,I73836,I73930,);
DFFARX1 I_4189 (I1027692,I2683,I73836,I73947,);
and I_4190 (I73955,I73947,I1027686);
nor I_4191 (I73972,I73930,I73955);
DFFARX1 I_4192 (I73972,I2683,I73836,I73804,);
nand I_4193 (I74003,I73947,I1027686);
nand I_4194 (I74020,I73870,I74003);
not I_4195 (I73816,I74020);
DFFARX1 I_4196 (I1027674,I2683,I73836,I74060,);
DFFARX1 I_4197 (I74060,I2683,I73836,I73825,);
nand I_4198 (I74082,I1027689,I1027677);
and I_4199 (I74099,I74082,I1027701);
DFFARX1 I_4200 (I74099,I2683,I73836,I74125,);
DFFARX1 I_4201 (I74125,I2683,I73836,I74142,);
not I_4202 (I73828,I74142);
not I_4203 (I74164,I74125);
nand I_4204 (I73813,I74164,I74003);
nor I_4205 (I74195,I1027683,I1027677);
not I_4206 (I74212,I74195);
nor I_4207 (I74229,I74164,I74212);
nor I_4208 (I74246,I73870,I74229);
DFFARX1 I_4209 (I74246,I2683,I73836,I73822,);
nor I_4210 (I74277,I73930,I74212);
nor I_4211 (I73810,I74125,I74277);
nor I_4212 (I73819,I74060,I74195);
nor I_4213 (I73807,I73930,I74195);
not I_4214 (I74363,I2690);
DFFARX1 I_4215 (I865772,I2683,I74363,I74389,);
not I_4216 (I74397,I74389);
nand I_4217 (I74414,I865787,I865766);
and I_4218 (I74431,I74414,I865769);
DFFARX1 I_4219 (I74431,I2683,I74363,I74457,);
DFFARX1 I_4220 (I865790,I2683,I74363,I74474,);
and I_4221 (I74482,I74474,I865769);
nor I_4222 (I74499,I74457,I74482);
DFFARX1 I_4223 (I74499,I2683,I74363,I74331,);
nand I_4224 (I74530,I74474,I865769);
nand I_4225 (I74547,I74397,I74530);
not I_4226 (I74343,I74547);
DFFARX1 I_4227 (I865766,I2683,I74363,I74587,);
DFFARX1 I_4228 (I74587,I2683,I74363,I74352,);
nand I_4229 (I74609,I865778,I865775);
and I_4230 (I74626,I74609,I865781);
DFFARX1 I_4231 (I74626,I2683,I74363,I74652,);
DFFARX1 I_4232 (I74652,I2683,I74363,I74669,);
not I_4233 (I74355,I74669);
not I_4234 (I74691,I74652);
nand I_4235 (I74340,I74691,I74530);
nor I_4236 (I74722,I865784,I865775);
not I_4237 (I74739,I74722);
nor I_4238 (I74756,I74691,I74739);
nor I_4239 (I74773,I74397,I74756);
DFFARX1 I_4240 (I74773,I2683,I74363,I74349,);
nor I_4241 (I74804,I74457,I74739);
nor I_4242 (I74337,I74652,I74804);
nor I_4243 (I74346,I74587,I74722);
nor I_4244 (I74334,I74457,I74722);
not I_4245 (I74890,I2690);
DFFARX1 I_4246 (I402655,I2683,I74890,I74916,);
not I_4247 (I74924,I74916);
nand I_4248 (I74941,I402676,I402670);
and I_4249 (I74958,I74941,I402652);
DFFARX1 I_4250 (I74958,I2683,I74890,I74984,);
DFFARX1 I_4251 (I402655,I2683,I74890,I75001,);
and I_4252 (I75009,I75001,I402664);
nor I_4253 (I75026,I74984,I75009);
DFFARX1 I_4254 (I75026,I2683,I74890,I74858,);
nand I_4255 (I75057,I75001,I402664);
nand I_4256 (I75074,I74924,I75057);
not I_4257 (I74870,I75074);
DFFARX1 I_4258 (I402661,I2683,I74890,I75114,);
DFFARX1 I_4259 (I75114,I2683,I74890,I74879,);
nand I_4260 (I75136,I402667,I402658);
and I_4261 (I75153,I75136,I402652);
DFFARX1 I_4262 (I75153,I2683,I74890,I75179,);
DFFARX1 I_4263 (I75179,I2683,I74890,I75196,);
not I_4264 (I74882,I75196);
not I_4265 (I75218,I75179);
nand I_4266 (I74867,I75218,I75057);
nor I_4267 (I75249,I402673,I402658);
not I_4268 (I75266,I75249);
nor I_4269 (I75283,I75218,I75266);
nor I_4270 (I75300,I74924,I75283);
DFFARX1 I_4271 (I75300,I2683,I74890,I74876,);
nor I_4272 (I75331,I74984,I75266);
nor I_4273 (I74864,I75179,I75331);
nor I_4274 (I74873,I75114,I75249);
nor I_4275 (I74861,I74984,I75249);
not I_4276 (I75417,I2690);
DFFARX1 I_4277 (I758114,I2683,I75417,I75443,);
not I_4278 (I75451,I75443);
nand I_4279 (I75468,I758132,I758126);
and I_4280 (I75485,I75468,I758105);
DFFARX1 I_4281 (I75485,I2683,I75417,I75511,);
DFFARX1 I_4282 (I758123,I2683,I75417,I75528,);
and I_4283 (I75536,I75528,I758108);
nor I_4284 (I75553,I75511,I75536);
DFFARX1 I_4285 (I75553,I2683,I75417,I75385,);
nand I_4286 (I75584,I75528,I758108);
nand I_4287 (I75601,I75451,I75584);
not I_4288 (I75397,I75601);
DFFARX1 I_4289 (I758120,I2683,I75417,I75641,);
DFFARX1 I_4290 (I75641,I2683,I75417,I75406,);
nand I_4291 (I75663,I758129,I758117);
and I_4292 (I75680,I75663,I758111);
DFFARX1 I_4293 (I75680,I2683,I75417,I75706,);
DFFARX1 I_4294 (I75706,I2683,I75417,I75723,);
not I_4295 (I75409,I75723);
not I_4296 (I75745,I75706);
nand I_4297 (I75394,I75745,I75584);
nor I_4298 (I75776,I758105,I758117);
not I_4299 (I75793,I75776);
nor I_4300 (I75810,I75745,I75793);
nor I_4301 (I75827,I75451,I75810);
DFFARX1 I_4302 (I75827,I2683,I75417,I75403,);
nor I_4303 (I75858,I75511,I75793);
nor I_4304 (I75391,I75706,I75858);
nor I_4305 (I75400,I75641,I75776);
nor I_4306 (I75388,I75511,I75776);
not I_4307 (I75944,I2690);
DFFARX1 I_4308 (I29033,I2683,I75944,I75970,);
not I_4309 (I75978,I75970);
nand I_4310 (I75995,I29021,I29027);
and I_4311 (I76012,I75995,I29030);
DFFARX1 I_4312 (I76012,I2683,I75944,I76038,);
DFFARX1 I_4313 (I29012,I2683,I75944,I76055,);
and I_4314 (I76063,I76055,I29018);
nor I_4315 (I76080,I76038,I76063);
DFFARX1 I_4316 (I76080,I2683,I75944,I75912,);
nand I_4317 (I76111,I76055,I29018);
nand I_4318 (I76128,I75978,I76111);
not I_4319 (I75924,I76128);
DFFARX1 I_4320 (I29012,I2683,I75944,I76168,);
DFFARX1 I_4321 (I76168,I2683,I75944,I75933,);
nand I_4322 (I76190,I29015,I29009);
and I_4323 (I76207,I76190,I29024);
DFFARX1 I_4324 (I76207,I2683,I75944,I76233,);
DFFARX1 I_4325 (I76233,I2683,I75944,I76250,);
not I_4326 (I75936,I76250);
not I_4327 (I76272,I76233);
nand I_4328 (I75921,I76272,I76111);
nor I_4329 (I76303,I29009,I29009);
not I_4330 (I76320,I76303);
nor I_4331 (I76337,I76272,I76320);
nor I_4332 (I76354,I75978,I76337);
DFFARX1 I_4333 (I76354,I2683,I75944,I75930,);
nor I_4334 (I76385,I76038,I76320);
nor I_4335 (I75918,I76233,I76385);
nor I_4336 (I75927,I76168,I76303);
nor I_4337 (I75915,I76038,I76303);
not I_4338 (I76471,I2690);
DFFARX1 I_4339 (I806881,I2683,I76471,I76497,);
not I_4340 (I76505,I76497);
nand I_4341 (I76522,I806878,I806884);
and I_4342 (I76539,I76522,I806881);
DFFARX1 I_4343 (I76539,I2683,I76471,I76565,);
DFFARX1 I_4344 (I806884,I2683,I76471,I76582,);
and I_4345 (I76590,I76582,I806878);
nor I_4346 (I76607,I76565,I76590);
DFFARX1 I_4347 (I76607,I2683,I76471,I76439,);
nand I_4348 (I76638,I76582,I806878);
nand I_4349 (I76655,I76505,I76638);
not I_4350 (I76451,I76655);
DFFARX1 I_4351 (I806887,I2683,I76471,I76695,);
DFFARX1 I_4352 (I76695,I2683,I76471,I76460,);
nand I_4353 (I76717,I806890,I806899);
and I_4354 (I76734,I76717,I806893);
DFFARX1 I_4355 (I76734,I2683,I76471,I76760,);
DFFARX1 I_4356 (I76760,I2683,I76471,I76777,);
not I_4357 (I76463,I76777);
not I_4358 (I76799,I76760);
nand I_4359 (I76448,I76799,I76638);
nor I_4360 (I76830,I806896,I806899);
not I_4361 (I76847,I76830);
nor I_4362 (I76864,I76799,I76847);
nor I_4363 (I76881,I76505,I76864);
DFFARX1 I_4364 (I76881,I2683,I76471,I76457,);
nor I_4365 (I76912,I76565,I76847);
nor I_4366 (I76445,I76760,I76912);
nor I_4367 (I76454,I76695,I76830);
nor I_4368 (I76442,I76565,I76830);
not I_4369 (I76998,I2690);
DFFARX1 I_4370 (I379108,I2683,I76998,I77024,);
not I_4371 (I77032,I77024);
nand I_4372 (I77049,I379102,I379093);
and I_4373 (I77066,I77049,I379114);
DFFARX1 I_4374 (I77066,I2683,I76998,I77092,);
DFFARX1 I_4375 (I379096,I2683,I76998,I77109,);
and I_4376 (I77117,I77109,I379090);
nor I_4377 (I77134,I77092,I77117);
DFFARX1 I_4378 (I77134,I2683,I76998,I76966,);
nand I_4379 (I77165,I77109,I379090);
nand I_4380 (I77182,I77032,I77165);
not I_4381 (I76978,I77182);
DFFARX1 I_4382 (I379090,I2683,I76998,I77222,);
DFFARX1 I_4383 (I77222,I2683,I76998,I76987,);
nand I_4384 (I77244,I379117,I379099);
and I_4385 (I77261,I77244,I379105);
DFFARX1 I_4386 (I77261,I2683,I76998,I77287,);
DFFARX1 I_4387 (I77287,I2683,I76998,I77304,);
not I_4388 (I76990,I77304);
not I_4389 (I77326,I77287);
nand I_4390 (I76975,I77326,I77165);
nor I_4391 (I77357,I379111,I379099);
not I_4392 (I77374,I77357);
nor I_4393 (I77391,I77326,I77374);
nor I_4394 (I77408,I77032,I77391);
DFFARX1 I_4395 (I77408,I2683,I76998,I76984,);
nor I_4396 (I77439,I77092,I77374);
nor I_4397 (I76972,I77287,I77439);
nor I_4398 (I76981,I77222,I77357);
nor I_4399 (I76969,I77092,I77357);
not I_4400 (I77525,I2690);
DFFARX1 I_4401 (I600612,I2683,I77525,I77551,);
not I_4402 (I77559,I77551);
nand I_4403 (I77576,I600603,I600621);
and I_4404 (I77593,I77576,I600600);
DFFARX1 I_4405 (I77593,I2683,I77525,I77619,);
DFFARX1 I_4406 (I600603,I2683,I77525,I77636,);
and I_4407 (I77644,I77636,I600606);
nor I_4408 (I77661,I77619,I77644);
DFFARX1 I_4409 (I77661,I2683,I77525,I77493,);
nand I_4410 (I77692,I77636,I600606);
nand I_4411 (I77709,I77559,I77692);
not I_4412 (I77505,I77709);
DFFARX1 I_4413 (I600600,I2683,I77525,I77749,);
DFFARX1 I_4414 (I77749,I2683,I77525,I77514,);
nand I_4415 (I77771,I600618,I600609);
and I_4416 (I77788,I77771,I600624);
DFFARX1 I_4417 (I77788,I2683,I77525,I77814,);
DFFARX1 I_4418 (I77814,I2683,I77525,I77831,);
not I_4419 (I77517,I77831);
not I_4420 (I77853,I77814);
nand I_4421 (I77502,I77853,I77692);
nor I_4422 (I77884,I600615,I600609);
not I_4423 (I77901,I77884);
nor I_4424 (I77918,I77853,I77901);
nor I_4425 (I77935,I77559,I77918);
DFFARX1 I_4426 (I77935,I2683,I77525,I77511,);
nor I_4427 (I77966,I77619,I77901);
nor I_4428 (I77499,I77814,I77966);
nor I_4429 (I77508,I77749,I77884);
nor I_4430 (I77496,I77619,I77884);
not I_4431 (I78052,I2690);
DFFARX1 I_4432 (I657049,I2683,I78052,I78078,);
not I_4433 (I78086,I78078);
nand I_4434 (I78103,I657046,I657061);
and I_4435 (I78120,I78103,I657043);
DFFARX1 I_4436 (I78120,I2683,I78052,I78146,);
DFFARX1 I_4437 (I657040,I2683,I78052,I78163,);
and I_4438 (I78171,I78163,I657040);
nor I_4439 (I78188,I78146,I78171);
DFFARX1 I_4440 (I78188,I2683,I78052,I78020,);
nand I_4441 (I78219,I78163,I657040);
nand I_4442 (I78236,I78086,I78219);
not I_4443 (I78032,I78236);
DFFARX1 I_4444 (I657043,I2683,I78052,I78276,);
DFFARX1 I_4445 (I78276,I2683,I78052,I78041,);
nand I_4446 (I78298,I657055,I657046);
and I_4447 (I78315,I78298,I657058);
DFFARX1 I_4448 (I78315,I2683,I78052,I78341,);
DFFARX1 I_4449 (I78341,I2683,I78052,I78358,);
not I_4450 (I78044,I78358);
not I_4451 (I78380,I78341);
nand I_4452 (I78029,I78380,I78219);
nor I_4453 (I78411,I657052,I657046);
not I_4454 (I78428,I78411);
nor I_4455 (I78445,I78380,I78428);
nor I_4456 (I78462,I78086,I78445);
DFFARX1 I_4457 (I78462,I2683,I78052,I78038,);
nor I_4458 (I78493,I78146,I78428);
nor I_4459 (I78026,I78341,I78493);
nor I_4460 (I78035,I78276,I78411);
nor I_4461 (I78023,I78146,I78411);
not I_4462 (I78579,I2690);
DFFARX1 I_4463 (I502930,I2683,I78579,I78605,);
not I_4464 (I78613,I78605);
nand I_4465 (I78630,I502921,I502939);
and I_4466 (I78647,I78630,I502918);
DFFARX1 I_4467 (I78647,I2683,I78579,I78673,);
DFFARX1 I_4468 (I502921,I2683,I78579,I78690,);
and I_4469 (I78698,I78690,I502924);
nor I_4470 (I78715,I78673,I78698);
DFFARX1 I_4471 (I78715,I2683,I78579,I78547,);
nand I_4472 (I78746,I78690,I502924);
nand I_4473 (I78763,I78613,I78746);
not I_4474 (I78559,I78763);
DFFARX1 I_4475 (I502918,I2683,I78579,I78803,);
DFFARX1 I_4476 (I78803,I2683,I78579,I78568,);
nand I_4477 (I78825,I502936,I502927);
and I_4478 (I78842,I78825,I502942);
DFFARX1 I_4479 (I78842,I2683,I78579,I78868,);
DFFARX1 I_4480 (I78868,I2683,I78579,I78885,);
not I_4481 (I78571,I78885);
not I_4482 (I78907,I78868);
nand I_4483 (I78556,I78907,I78746);
nor I_4484 (I78938,I502933,I502927);
not I_4485 (I78955,I78938);
nor I_4486 (I78972,I78907,I78955);
nor I_4487 (I78989,I78613,I78972);
DFFARX1 I_4488 (I78989,I2683,I78579,I78565,);
nor I_4489 (I79020,I78673,I78955);
nor I_4490 (I78553,I78868,I79020);
nor I_4491 (I78562,I78803,I78938);
nor I_4492 (I78550,I78673,I78938);
not I_4493 (I79106,I2690);
DFFARX1 I_4494 (I563620,I2683,I79106,I79132,);
not I_4495 (I79140,I79132);
nand I_4496 (I79157,I563611,I563629);
and I_4497 (I79174,I79157,I563608);
DFFARX1 I_4498 (I79174,I2683,I79106,I79200,);
DFFARX1 I_4499 (I563611,I2683,I79106,I79217,);
and I_4500 (I79225,I79217,I563614);
nor I_4501 (I79242,I79200,I79225);
DFFARX1 I_4502 (I79242,I2683,I79106,I79074,);
nand I_4503 (I79273,I79217,I563614);
nand I_4504 (I79290,I79140,I79273);
not I_4505 (I79086,I79290);
DFFARX1 I_4506 (I563608,I2683,I79106,I79330,);
DFFARX1 I_4507 (I79330,I2683,I79106,I79095,);
nand I_4508 (I79352,I563626,I563617);
and I_4509 (I79369,I79352,I563632);
DFFARX1 I_4510 (I79369,I2683,I79106,I79395,);
DFFARX1 I_4511 (I79395,I2683,I79106,I79412,);
not I_4512 (I79098,I79412);
not I_4513 (I79434,I79395);
nand I_4514 (I79083,I79434,I79273);
nor I_4515 (I79465,I563623,I563617);
not I_4516 (I79482,I79465);
nor I_4517 (I79499,I79434,I79482);
nor I_4518 (I79516,I79140,I79499);
DFFARX1 I_4519 (I79516,I2683,I79106,I79092,);
nor I_4520 (I79547,I79200,I79482);
nor I_4521 (I79080,I79395,I79547);
nor I_4522 (I79089,I79330,I79465);
nor I_4523 (I79077,I79200,I79465);
not I_4524 (I79633,I2690);
DFFARX1 I_4525 (I262786,I2683,I79633,I79659,);
not I_4526 (I79667,I79659);
nand I_4527 (I79684,I262768,I262783);
and I_4528 (I79701,I79684,I262759);
DFFARX1 I_4529 (I79701,I2683,I79633,I79727,);
DFFARX1 I_4530 (I262762,I2683,I79633,I79744,);
and I_4531 (I79752,I79744,I262777);
nor I_4532 (I79769,I79727,I79752);
DFFARX1 I_4533 (I79769,I2683,I79633,I79601,);
nand I_4534 (I79800,I79744,I262777);
nand I_4535 (I79817,I79667,I79800);
not I_4536 (I79613,I79817);
DFFARX1 I_4537 (I262780,I2683,I79633,I79857,);
DFFARX1 I_4538 (I79857,I2683,I79633,I79622,);
nand I_4539 (I79879,I262759,I262771);
and I_4540 (I79896,I79879,I262765);
DFFARX1 I_4541 (I79896,I2683,I79633,I79922,);
DFFARX1 I_4542 (I79922,I2683,I79633,I79939,);
not I_4543 (I79625,I79939);
not I_4544 (I79961,I79922);
nand I_4545 (I79610,I79961,I79800);
nor I_4546 (I79992,I262774,I262771);
not I_4547 (I80009,I79992);
nor I_4548 (I80026,I79961,I80009);
nor I_4549 (I80043,I79667,I80026);
DFFARX1 I_4550 (I80043,I2683,I79633,I79619,);
nor I_4551 (I80074,I79727,I80009);
nor I_4552 (I79607,I79922,I80074);
nor I_4553 (I79616,I79857,I79992);
nor I_4554 (I79604,I79727,I79992);
not I_4555 (I80160,I2690);
DFFARX1 I_4556 (I321444,I2683,I80160,I80186,);
not I_4557 (I80194,I80186);
nand I_4558 (I80211,I321438,I321429);
and I_4559 (I80228,I80211,I321450);
DFFARX1 I_4560 (I80228,I2683,I80160,I80254,);
DFFARX1 I_4561 (I321432,I2683,I80160,I80271,);
and I_4562 (I80279,I80271,I321426);
nor I_4563 (I80296,I80254,I80279);
DFFARX1 I_4564 (I80296,I2683,I80160,I80128,);
nand I_4565 (I80327,I80271,I321426);
nand I_4566 (I80344,I80194,I80327);
not I_4567 (I80140,I80344);
DFFARX1 I_4568 (I321426,I2683,I80160,I80384,);
DFFARX1 I_4569 (I80384,I2683,I80160,I80149,);
nand I_4570 (I80406,I321453,I321435);
and I_4571 (I80423,I80406,I321441);
DFFARX1 I_4572 (I80423,I2683,I80160,I80449,);
DFFARX1 I_4573 (I80449,I2683,I80160,I80466,);
not I_4574 (I80152,I80466);
not I_4575 (I80488,I80449);
nand I_4576 (I80137,I80488,I80327);
nor I_4577 (I80519,I321447,I321435);
not I_4578 (I80536,I80519);
nor I_4579 (I80553,I80488,I80536);
nor I_4580 (I80570,I80194,I80553);
DFFARX1 I_4581 (I80570,I2683,I80160,I80146,);
nor I_4582 (I80601,I80254,I80536);
nor I_4583 (I80134,I80449,I80601);
nor I_4584 (I80143,I80384,I80519);
nor I_4585 (I80131,I80254,I80519);
not I_4586 (I80687,I2690);
DFFARX1 I_4587 (I144417,I2683,I80687,I80713,);
not I_4588 (I80721,I80713);
nand I_4589 (I80738,I144411,I144405);
and I_4590 (I80755,I80738,I144426);
DFFARX1 I_4591 (I80755,I2683,I80687,I80781,);
DFFARX1 I_4592 (I144423,I2683,I80687,I80798,);
and I_4593 (I80806,I80798,I144420);
nor I_4594 (I80823,I80781,I80806);
DFFARX1 I_4595 (I80823,I2683,I80687,I80655,);
nand I_4596 (I80854,I80798,I144420);
nand I_4597 (I80871,I80721,I80854);
not I_4598 (I80667,I80871);
DFFARX1 I_4599 (I144405,I2683,I80687,I80911,);
DFFARX1 I_4600 (I80911,I2683,I80687,I80676,);
nand I_4601 (I80933,I144408,I144408);
and I_4602 (I80950,I80933,I144429);
DFFARX1 I_4603 (I80950,I2683,I80687,I80976,);
DFFARX1 I_4604 (I80976,I2683,I80687,I80993,);
not I_4605 (I80679,I80993);
not I_4606 (I81015,I80976);
nand I_4607 (I80664,I81015,I80854);
nor I_4608 (I81046,I144414,I144408);
not I_4609 (I81063,I81046);
nor I_4610 (I81080,I81015,I81063);
nor I_4611 (I81097,I80721,I81080);
DFFARX1 I_4612 (I81097,I2683,I80687,I80673,);
nor I_4613 (I81128,I80781,I81063);
nor I_4614 (I80661,I80976,I81128);
nor I_4615 (I80670,I80911,I81046);
nor I_4616 (I80658,I80781,I81046);
not I_4617 (I81214,I2690);
DFFARX1 I_4618 (I400275,I2683,I81214,I81240,);
not I_4619 (I81248,I81240);
nand I_4620 (I81265,I400296,I400290);
and I_4621 (I81282,I81265,I400272);
DFFARX1 I_4622 (I81282,I2683,I81214,I81308,);
DFFARX1 I_4623 (I400275,I2683,I81214,I81325,);
and I_4624 (I81333,I81325,I400284);
nor I_4625 (I81350,I81308,I81333);
DFFARX1 I_4626 (I81350,I2683,I81214,I81182,);
nand I_4627 (I81381,I81325,I400284);
nand I_4628 (I81398,I81248,I81381);
not I_4629 (I81194,I81398);
DFFARX1 I_4630 (I400281,I2683,I81214,I81438,);
DFFARX1 I_4631 (I81438,I2683,I81214,I81203,);
nand I_4632 (I81460,I400287,I400278);
and I_4633 (I81477,I81460,I400272);
DFFARX1 I_4634 (I81477,I2683,I81214,I81503,);
DFFARX1 I_4635 (I81503,I2683,I81214,I81520,);
not I_4636 (I81206,I81520);
not I_4637 (I81542,I81503);
nand I_4638 (I81191,I81542,I81381);
nor I_4639 (I81573,I400293,I400278);
not I_4640 (I81590,I81573);
nor I_4641 (I81607,I81542,I81590);
nor I_4642 (I81624,I81248,I81607);
DFFARX1 I_4643 (I81624,I2683,I81214,I81200,);
nor I_4644 (I81655,I81308,I81590);
nor I_4645 (I81188,I81503,I81655);
nor I_4646 (I81197,I81438,I81573);
nor I_4647 (I81185,I81308,I81573);
not I_4648 (I81741,I2690);
DFFARX1 I_4649 (I745840,I2683,I81741,I81767,);
not I_4650 (I81775,I81767);
nand I_4651 (I81792,I745858,I745852);
and I_4652 (I81809,I81792,I745831);
DFFARX1 I_4653 (I81809,I2683,I81741,I81835,);
DFFARX1 I_4654 (I745849,I2683,I81741,I81852,);
and I_4655 (I81860,I81852,I745834);
nor I_4656 (I81877,I81835,I81860);
DFFARX1 I_4657 (I81877,I2683,I81741,I81709,);
nand I_4658 (I81908,I81852,I745834);
nand I_4659 (I81925,I81775,I81908);
not I_4660 (I81721,I81925);
DFFARX1 I_4661 (I745846,I2683,I81741,I81965,);
DFFARX1 I_4662 (I81965,I2683,I81741,I81730,);
nand I_4663 (I81987,I745855,I745843);
and I_4664 (I82004,I81987,I745837);
DFFARX1 I_4665 (I82004,I2683,I81741,I82030,);
DFFARX1 I_4666 (I82030,I2683,I81741,I82047,);
not I_4667 (I81733,I82047);
not I_4668 (I82069,I82030);
nand I_4669 (I81718,I82069,I81908);
nor I_4670 (I82100,I745831,I745843);
not I_4671 (I82117,I82100);
nor I_4672 (I82134,I82069,I82117);
nor I_4673 (I82151,I81775,I82134);
DFFARX1 I_4674 (I82151,I2683,I81741,I81727,);
nor I_4675 (I82182,I81835,I82117);
nor I_4676 (I81715,I82030,I82182);
nor I_4677 (I81724,I81965,I82100);
nor I_4678 (I81712,I81835,I82100);
not I_4679 (I82268,I2690);
DFFARX1 I_4680 (I237490,I2683,I82268,I82294,);
not I_4681 (I82302,I82294);
nand I_4682 (I82319,I237472,I237487);
and I_4683 (I82336,I82319,I237463);
DFFARX1 I_4684 (I82336,I2683,I82268,I82362,);
DFFARX1 I_4685 (I237466,I2683,I82268,I82379,);
and I_4686 (I82387,I82379,I237481);
nor I_4687 (I82404,I82362,I82387);
DFFARX1 I_4688 (I82404,I2683,I82268,I82236,);
nand I_4689 (I82435,I82379,I237481);
nand I_4690 (I82452,I82302,I82435);
not I_4691 (I82248,I82452);
DFFARX1 I_4692 (I237484,I2683,I82268,I82492,);
DFFARX1 I_4693 (I82492,I2683,I82268,I82257,);
nand I_4694 (I82514,I237463,I237475);
and I_4695 (I82531,I82514,I237469);
DFFARX1 I_4696 (I82531,I2683,I82268,I82557,);
DFFARX1 I_4697 (I82557,I2683,I82268,I82574,);
not I_4698 (I82260,I82574);
not I_4699 (I82596,I82557);
nand I_4700 (I82245,I82596,I82435);
nor I_4701 (I82627,I237478,I237475);
not I_4702 (I82644,I82627);
nor I_4703 (I82661,I82596,I82644);
nor I_4704 (I82678,I82302,I82661);
DFFARX1 I_4705 (I82678,I2683,I82268,I82254,);
nor I_4706 (I82709,I82362,I82644);
nor I_4707 (I82242,I82557,I82709);
nor I_4708 (I82251,I82492,I82627);
nor I_4709 (I82239,I82362,I82627);
not I_4710 (I82795,I2690);
DFFARX1 I_4711 (I903920,I2683,I82795,I82821,);
not I_4712 (I82829,I82821);
nand I_4713 (I82846,I903935,I903914);
and I_4714 (I82863,I82846,I903917);
DFFARX1 I_4715 (I82863,I2683,I82795,I82889,);
DFFARX1 I_4716 (I903938,I2683,I82795,I82906,);
and I_4717 (I82914,I82906,I903917);
nor I_4718 (I82931,I82889,I82914);
DFFARX1 I_4719 (I82931,I2683,I82795,I82763,);
nand I_4720 (I82962,I82906,I903917);
nand I_4721 (I82979,I82829,I82962);
not I_4722 (I82775,I82979);
DFFARX1 I_4723 (I903914,I2683,I82795,I83019,);
DFFARX1 I_4724 (I83019,I2683,I82795,I82784,);
nand I_4725 (I83041,I903926,I903923);
and I_4726 (I83058,I83041,I903929);
DFFARX1 I_4727 (I83058,I2683,I82795,I83084,);
DFFARX1 I_4728 (I83084,I2683,I82795,I83101,);
not I_4729 (I82787,I83101);
not I_4730 (I83123,I83084);
nand I_4731 (I82772,I83123,I82962);
nor I_4732 (I83154,I903932,I903923);
not I_4733 (I83171,I83154);
nor I_4734 (I83188,I83123,I83171);
nor I_4735 (I83205,I82829,I83188);
DFFARX1 I_4736 (I83205,I2683,I82795,I82781,);
nor I_4737 (I83236,I82889,I83171);
nor I_4738 (I82769,I83084,I83236);
nor I_4739 (I82778,I83019,I83154);
nor I_4740 (I82766,I82889,I83154);
not I_4741 (I83322,I2690);
DFFARX1 I_4742 (I500618,I2683,I83322,I83348,);
not I_4743 (I83356,I83348);
nand I_4744 (I83373,I500609,I500627);
and I_4745 (I83390,I83373,I500606);
DFFARX1 I_4746 (I83390,I2683,I83322,I83416,);
DFFARX1 I_4747 (I500609,I2683,I83322,I83433,);
and I_4748 (I83441,I83433,I500612);
nor I_4749 (I83458,I83416,I83441);
DFFARX1 I_4750 (I83458,I2683,I83322,I83290,);
nand I_4751 (I83489,I83433,I500612);
nand I_4752 (I83506,I83356,I83489);
not I_4753 (I83302,I83506);
DFFARX1 I_4754 (I500606,I2683,I83322,I83546,);
DFFARX1 I_4755 (I83546,I2683,I83322,I83311,);
nand I_4756 (I83568,I500624,I500615);
and I_4757 (I83585,I83568,I500630);
DFFARX1 I_4758 (I83585,I2683,I83322,I83611,);
DFFARX1 I_4759 (I83611,I2683,I83322,I83628,);
not I_4760 (I83314,I83628);
not I_4761 (I83650,I83611);
nand I_4762 (I83299,I83650,I83489);
nor I_4763 (I83681,I500621,I500615);
not I_4764 (I83698,I83681);
nor I_4765 (I83715,I83650,I83698);
nor I_4766 (I83732,I83356,I83715);
DFFARX1 I_4767 (I83732,I2683,I83322,I83308,);
nor I_4768 (I83763,I83416,I83698);
nor I_4769 (I83296,I83611,I83763);
nor I_4770 (I83305,I83546,I83681);
nor I_4771 (I83293,I83416,I83681);
not I_4772 (I83849,I2690);
DFFARX1 I_4773 (I822028,I2683,I83849,I83875,);
not I_4774 (I83883,I83875);
nand I_4775 (I83900,I822025,I822031);
and I_4776 (I83917,I83900,I822028);
DFFARX1 I_4777 (I83917,I2683,I83849,I83943,);
DFFARX1 I_4778 (I822031,I2683,I83849,I83960,);
and I_4779 (I83968,I83960,I822025);
nor I_4780 (I83985,I83943,I83968);
DFFARX1 I_4781 (I83985,I2683,I83849,I83817,);
nand I_4782 (I84016,I83960,I822025);
nand I_4783 (I84033,I83883,I84016);
not I_4784 (I83829,I84033);
DFFARX1 I_4785 (I822034,I2683,I83849,I84073,);
DFFARX1 I_4786 (I84073,I2683,I83849,I83838,);
nand I_4787 (I84095,I822037,I822046);
and I_4788 (I84112,I84095,I822040);
DFFARX1 I_4789 (I84112,I2683,I83849,I84138,);
DFFARX1 I_4790 (I84138,I2683,I83849,I84155,);
not I_4791 (I83841,I84155);
not I_4792 (I84177,I84138);
nand I_4793 (I83826,I84177,I84016);
nor I_4794 (I84208,I822043,I822046);
not I_4795 (I84225,I84208);
nor I_4796 (I84242,I84177,I84225);
nor I_4797 (I84259,I83883,I84242);
DFFARX1 I_4798 (I84259,I2683,I83849,I83835,);
nor I_4799 (I84290,I83943,I84225);
nor I_4800 (I83823,I84138,I84290);
nor I_4801 (I83832,I84073,I84208);
nor I_4802 (I83820,I83943,I84208);
not I_4803 (I84376,I2690);
DFFARX1 I_4804 (I172977,I2683,I84376,I84402,);
not I_4805 (I84410,I84402);
nand I_4806 (I84427,I172971,I172965);
and I_4807 (I84444,I84427,I172986);
DFFARX1 I_4808 (I84444,I2683,I84376,I84470,);
DFFARX1 I_4809 (I172983,I2683,I84376,I84487,);
and I_4810 (I84495,I84487,I172980);
nor I_4811 (I84512,I84470,I84495);
DFFARX1 I_4812 (I84512,I2683,I84376,I84344,);
nand I_4813 (I84543,I84487,I172980);
nand I_4814 (I84560,I84410,I84543);
not I_4815 (I84356,I84560);
DFFARX1 I_4816 (I172965,I2683,I84376,I84600,);
DFFARX1 I_4817 (I84600,I2683,I84376,I84365,);
nand I_4818 (I84622,I172968,I172968);
and I_4819 (I84639,I84622,I172989);
DFFARX1 I_4820 (I84639,I2683,I84376,I84665,);
DFFARX1 I_4821 (I84665,I2683,I84376,I84682,);
not I_4822 (I84368,I84682);
not I_4823 (I84704,I84665);
nand I_4824 (I84353,I84704,I84543);
nor I_4825 (I84735,I172974,I172968);
not I_4826 (I84752,I84735);
nor I_4827 (I84769,I84704,I84752);
nor I_4828 (I84786,I84410,I84769);
DFFARX1 I_4829 (I84786,I2683,I84376,I84362,);
nor I_4830 (I84817,I84470,I84752);
nor I_4831 (I84350,I84665,I84817);
nor I_4832 (I84359,I84600,I84735);
nor I_4833 (I84347,I84470,I84735);
not I_4834 (I84903,I2690);
DFFARX1 I_4835 (I1023747,I2683,I84903,I84929,);
not I_4836 (I84937,I84929);
nand I_4837 (I84954,I1023753,I1023771);
and I_4838 (I84971,I84954,I1023768);
DFFARX1 I_4839 (I84971,I2683,I84903,I84997,);
DFFARX1 I_4840 (I1023765,I2683,I84903,I85014,);
and I_4841 (I85022,I85014,I1023759);
nor I_4842 (I85039,I84997,I85022);
DFFARX1 I_4843 (I85039,I2683,I84903,I84871,);
nand I_4844 (I85070,I85014,I1023759);
nand I_4845 (I85087,I84937,I85070);
not I_4846 (I84883,I85087);
DFFARX1 I_4847 (I1023747,I2683,I84903,I85127,);
DFFARX1 I_4848 (I85127,I2683,I84903,I84892,);
nand I_4849 (I85149,I1023762,I1023750);
and I_4850 (I85166,I85149,I1023774);
DFFARX1 I_4851 (I85166,I2683,I84903,I85192,);
DFFARX1 I_4852 (I85192,I2683,I84903,I85209,);
not I_4853 (I84895,I85209);
not I_4854 (I85231,I85192);
nand I_4855 (I84880,I85231,I85070);
nor I_4856 (I85262,I1023756,I1023750);
not I_4857 (I85279,I85262);
nor I_4858 (I85296,I85231,I85279);
nor I_4859 (I85313,I84937,I85296);
DFFARX1 I_4860 (I85313,I2683,I84903,I84889,);
nor I_4861 (I85344,I84997,I85279);
nor I_4862 (I84877,I85192,I85344);
nor I_4863 (I84886,I85127,I85262);
nor I_4864 (I84874,I84997,I85262);
not I_4865 (I85430,I2690);
DFFARX1 I_4866 (I797344,I2683,I85430,I85456,);
not I_4867 (I85464,I85456);
nand I_4868 (I85481,I797341,I797347);
and I_4869 (I85498,I85481,I797344);
DFFARX1 I_4870 (I85498,I2683,I85430,I85524,);
DFFARX1 I_4871 (I797347,I2683,I85430,I85541,);
and I_4872 (I85549,I85541,I797341);
nor I_4873 (I85566,I85524,I85549);
DFFARX1 I_4874 (I85566,I2683,I85430,I85398,);
nand I_4875 (I85597,I85541,I797341);
nand I_4876 (I85614,I85464,I85597);
not I_4877 (I85410,I85614);
DFFARX1 I_4878 (I797350,I2683,I85430,I85654,);
DFFARX1 I_4879 (I85654,I2683,I85430,I85419,);
nand I_4880 (I85676,I797353,I797362);
and I_4881 (I85693,I85676,I797356);
DFFARX1 I_4882 (I85693,I2683,I85430,I85719,);
DFFARX1 I_4883 (I85719,I2683,I85430,I85736,);
not I_4884 (I85422,I85736);
not I_4885 (I85758,I85719);
nand I_4886 (I85407,I85758,I85597);
nor I_4887 (I85789,I797359,I797362);
not I_4888 (I85806,I85789);
nor I_4889 (I85823,I85758,I85806);
nor I_4890 (I85840,I85464,I85823);
DFFARX1 I_4891 (I85840,I2683,I85430,I85416,);
nor I_4892 (I85871,I85524,I85806);
nor I_4893 (I85404,I85719,I85871);
nor I_4894 (I85413,I85654,I85789);
nor I_4895 (I85401,I85524,I85789);
not I_4896 (I85957,I2690);
DFFARX1 I_4897 (I617374,I2683,I85957,I85983,);
not I_4898 (I85991,I85983);
nand I_4899 (I86008,I617365,I617383);
and I_4900 (I86025,I86008,I617362);
DFFARX1 I_4901 (I86025,I2683,I85957,I86051,);
DFFARX1 I_4902 (I617365,I2683,I85957,I86068,);
and I_4903 (I86076,I86068,I617368);
nor I_4904 (I86093,I86051,I86076);
DFFARX1 I_4905 (I86093,I2683,I85957,I85925,);
nand I_4906 (I86124,I86068,I617368);
nand I_4907 (I86141,I85991,I86124);
not I_4908 (I85937,I86141);
DFFARX1 I_4909 (I617362,I2683,I85957,I86181,);
DFFARX1 I_4910 (I86181,I2683,I85957,I85946,);
nand I_4911 (I86203,I617380,I617371);
and I_4912 (I86220,I86203,I617386);
DFFARX1 I_4913 (I86220,I2683,I85957,I86246,);
DFFARX1 I_4914 (I86246,I2683,I85957,I86263,);
not I_4915 (I85949,I86263);
not I_4916 (I86285,I86246);
nand I_4917 (I85934,I86285,I86124);
nor I_4918 (I86316,I617377,I617371);
not I_4919 (I86333,I86316);
nor I_4920 (I86350,I86285,I86333);
nor I_4921 (I86367,I85991,I86350);
DFFARX1 I_4922 (I86367,I2683,I85957,I85943,);
nor I_4923 (I86398,I86051,I86333);
nor I_4924 (I85931,I86246,I86398);
nor I_4925 (I85940,I86181,I86316);
nor I_4926 (I85928,I86051,I86316);
not I_4927 (I86484,I2690);
DFFARX1 I_4928 (I966820,I2683,I86484,I86510,);
not I_4929 (I86518,I86510);
nand I_4930 (I86535,I966814,I966835);
and I_4931 (I86552,I86535,I966826);
DFFARX1 I_4932 (I86552,I2683,I86484,I86578,);
DFFARX1 I_4933 (I966817,I2683,I86484,I86595,);
and I_4934 (I86603,I86595,I966829);
nor I_4935 (I86620,I86578,I86603);
DFFARX1 I_4936 (I86620,I2683,I86484,I86452,);
nand I_4937 (I86651,I86595,I966829);
nand I_4938 (I86668,I86518,I86651);
not I_4939 (I86464,I86668);
DFFARX1 I_4940 (I966817,I2683,I86484,I86708,);
DFFARX1 I_4941 (I86708,I2683,I86484,I86473,);
nand I_4942 (I86730,I966838,I966823);
and I_4943 (I86747,I86730,I966814);
DFFARX1 I_4944 (I86747,I2683,I86484,I86773,);
DFFARX1 I_4945 (I86773,I2683,I86484,I86790,);
not I_4946 (I86476,I86790);
not I_4947 (I86812,I86773);
nand I_4948 (I86461,I86812,I86651);
nor I_4949 (I86843,I966832,I966823);
not I_4950 (I86860,I86843);
nor I_4951 (I86877,I86812,I86860);
nor I_4952 (I86894,I86518,I86877);
DFFARX1 I_4953 (I86894,I2683,I86484,I86470,);
nor I_4954 (I86925,I86578,I86860);
nor I_4955 (I86458,I86773,I86925);
nor I_4956 (I86467,I86708,I86843);
nor I_4957 (I86455,I86578,I86843);
not I_4958 (I87011,I2690);
DFFARX1 I_4959 (I243287,I2683,I87011,I87037,);
not I_4960 (I87045,I87037);
nand I_4961 (I87062,I243269,I243284);
and I_4962 (I87079,I87062,I243260);
DFFARX1 I_4963 (I87079,I2683,I87011,I87105,);
DFFARX1 I_4964 (I243263,I2683,I87011,I87122,);
and I_4965 (I87130,I87122,I243278);
nor I_4966 (I87147,I87105,I87130);
DFFARX1 I_4967 (I87147,I2683,I87011,I86979,);
nand I_4968 (I87178,I87122,I243278);
nand I_4969 (I87195,I87045,I87178);
not I_4970 (I86991,I87195);
DFFARX1 I_4971 (I243281,I2683,I87011,I87235,);
DFFARX1 I_4972 (I87235,I2683,I87011,I87000,);
nand I_4973 (I87257,I243260,I243272);
and I_4974 (I87274,I87257,I243266);
DFFARX1 I_4975 (I87274,I2683,I87011,I87300,);
DFFARX1 I_4976 (I87300,I2683,I87011,I87317,);
not I_4977 (I87003,I87317);
not I_4978 (I87339,I87300);
nand I_4979 (I86988,I87339,I87178);
nor I_4980 (I87370,I243275,I243272);
not I_4981 (I87387,I87370);
nor I_4982 (I87404,I87339,I87387);
nor I_4983 (I87421,I87045,I87404);
DFFARX1 I_4984 (I87421,I2683,I87011,I86997,);
nor I_4985 (I87452,I87105,I87387);
nor I_4986 (I86985,I87300,I87452);
nor I_4987 (I86994,I87235,I87370);
nor I_4988 (I86982,I87105,I87370);
not I_4989 (I87538,I2690);
DFFARX1 I_4990 (I367684,I2683,I87538,I87564,);
not I_4991 (I87572,I87564);
nand I_4992 (I87589,I367678,I367669);
and I_4993 (I87606,I87589,I367690);
DFFARX1 I_4994 (I87606,I2683,I87538,I87632,);
DFFARX1 I_4995 (I367672,I2683,I87538,I87649,);
and I_4996 (I87657,I87649,I367666);
nor I_4997 (I87674,I87632,I87657);
DFFARX1 I_4998 (I87674,I2683,I87538,I87506,);
nand I_4999 (I87705,I87649,I367666);
nand I_5000 (I87722,I87572,I87705);
not I_5001 (I87518,I87722);
DFFARX1 I_5002 (I367666,I2683,I87538,I87762,);
DFFARX1 I_5003 (I87762,I2683,I87538,I87527,);
nand I_5004 (I87784,I367693,I367675);
and I_5005 (I87801,I87784,I367681);
DFFARX1 I_5006 (I87801,I2683,I87538,I87827,);
DFFARX1 I_5007 (I87827,I2683,I87538,I87844,);
not I_5008 (I87530,I87844);
not I_5009 (I87866,I87827);
nand I_5010 (I87515,I87866,I87705);
nor I_5011 (I87897,I367687,I367675);
not I_5012 (I87914,I87897);
nor I_5013 (I87931,I87866,I87914);
nor I_5014 (I87948,I87572,I87931);
DFFARX1 I_5015 (I87948,I2683,I87538,I87524,);
nor I_5016 (I87979,I87632,I87914);
nor I_5017 (I87512,I87827,I87979);
nor I_5018 (I87521,I87762,I87897);
nor I_5019 (I87509,I87632,I87897);
not I_5020 (I88065,I2690);
DFFARX1 I_5021 (I608126,I2683,I88065,I88091,);
not I_5022 (I88099,I88091);
nand I_5023 (I88116,I608117,I608135);
and I_5024 (I88133,I88116,I608114);
DFFARX1 I_5025 (I88133,I2683,I88065,I88159,);
DFFARX1 I_5026 (I608117,I2683,I88065,I88176,);
and I_5027 (I88184,I88176,I608120);
nor I_5028 (I88201,I88159,I88184);
DFFARX1 I_5029 (I88201,I2683,I88065,I88033,);
nand I_5030 (I88232,I88176,I608120);
nand I_5031 (I88249,I88099,I88232);
not I_5032 (I88045,I88249);
DFFARX1 I_5033 (I608114,I2683,I88065,I88289,);
DFFARX1 I_5034 (I88289,I2683,I88065,I88054,);
nand I_5035 (I88311,I608132,I608123);
and I_5036 (I88328,I88311,I608138);
DFFARX1 I_5037 (I88328,I2683,I88065,I88354,);
DFFARX1 I_5038 (I88354,I2683,I88065,I88371,);
not I_5039 (I88057,I88371);
not I_5040 (I88393,I88354);
nand I_5041 (I88042,I88393,I88232);
nor I_5042 (I88424,I608129,I608123);
not I_5043 (I88441,I88424);
nor I_5044 (I88458,I88393,I88441);
nor I_5045 (I88475,I88099,I88458);
DFFARX1 I_5046 (I88475,I2683,I88065,I88051,);
nor I_5047 (I88506,I88159,I88441);
nor I_5048 (I88039,I88354,I88506);
nor I_5049 (I88048,I88289,I88424);
nor I_5050 (I88036,I88159,I88424);
not I_5051 (I88592,I2690);
DFFARX1 I_5052 (I860570,I2683,I88592,I88618,);
not I_5053 (I88626,I88618);
nand I_5054 (I88643,I860585,I860564);
and I_5055 (I88660,I88643,I860567);
DFFARX1 I_5056 (I88660,I2683,I88592,I88686,);
DFFARX1 I_5057 (I860588,I2683,I88592,I88703,);
and I_5058 (I88711,I88703,I860567);
nor I_5059 (I88728,I88686,I88711);
DFFARX1 I_5060 (I88728,I2683,I88592,I88560,);
nand I_5061 (I88759,I88703,I860567);
nand I_5062 (I88776,I88626,I88759);
not I_5063 (I88572,I88776);
DFFARX1 I_5064 (I860564,I2683,I88592,I88816,);
DFFARX1 I_5065 (I88816,I2683,I88592,I88581,);
nand I_5066 (I88838,I860576,I860573);
and I_5067 (I88855,I88838,I860579);
DFFARX1 I_5068 (I88855,I2683,I88592,I88881,);
DFFARX1 I_5069 (I88881,I2683,I88592,I88898,);
not I_5070 (I88584,I88898);
not I_5071 (I88920,I88881);
nand I_5072 (I88569,I88920,I88759);
nor I_5073 (I88951,I860582,I860573);
not I_5074 (I88968,I88951);
nor I_5075 (I88985,I88920,I88968);
nor I_5076 (I89002,I88626,I88985);
DFFARX1 I_5077 (I89002,I2683,I88592,I88578,);
nor I_5078 (I89033,I88686,I88968);
nor I_5079 (I88566,I88881,I89033);
nor I_5080 (I88575,I88816,I88951);
nor I_5081 (I88563,I88686,I88951);
not I_5082 (I89119,I2690);
DFFARX1 I_5083 (I658103,I2683,I89119,I89145,);
not I_5084 (I89153,I89145);
nand I_5085 (I89170,I658100,I658115);
and I_5086 (I89187,I89170,I658097);
DFFARX1 I_5087 (I89187,I2683,I89119,I89213,);
DFFARX1 I_5088 (I658094,I2683,I89119,I89230,);
and I_5089 (I89238,I89230,I658094);
nor I_5090 (I89255,I89213,I89238);
DFFARX1 I_5091 (I89255,I2683,I89119,I89087,);
nand I_5092 (I89286,I89230,I658094);
nand I_5093 (I89303,I89153,I89286);
not I_5094 (I89099,I89303);
DFFARX1 I_5095 (I658097,I2683,I89119,I89343,);
DFFARX1 I_5096 (I89343,I2683,I89119,I89108,);
nand I_5097 (I89365,I658109,I658100);
and I_5098 (I89382,I89365,I658112);
DFFARX1 I_5099 (I89382,I2683,I89119,I89408,);
DFFARX1 I_5100 (I89408,I2683,I89119,I89425,);
not I_5101 (I89111,I89425);
not I_5102 (I89447,I89408);
nand I_5103 (I89096,I89447,I89286);
nor I_5104 (I89478,I658106,I658100);
not I_5105 (I89495,I89478);
nor I_5106 (I89512,I89447,I89495);
nor I_5107 (I89529,I89153,I89512);
DFFARX1 I_5108 (I89529,I2683,I89119,I89105,);
nor I_5109 (I89560,I89213,I89495);
nor I_5110 (I89093,I89408,I89560);
nor I_5111 (I89102,I89343,I89478);
nor I_5112 (I89090,I89213,I89478);
not I_5113 (I89646,I2690);
DFFARX1 I_5114 (I809686,I2683,I89646,I89672,);
not I_5115 (I89680,I89672);
nand I_5116 (I89697,I809683,I809689);
and I_5117 (I89714,I89697,I809686);
DFFARX1 I_5118 (I89714,I2683,I89646,I89740,);
DFFARX1 I_5119 (I809689,I2683,I89646,I89757,);
and I_5120 (I89765,I89757,I809683);
nor I_5121 (I89782,I89740,I89765);
DFFARX1 I_5122 (I89782,I2683,I89646,I89614,);
nand I_5123 (I89813,I89757,I809683);
nand I_5124 (I89830,I89680,I89813);
not I_5125 (I89626,I89830);
DFFARX1 I_5126 (I809692,I2683,I89646,I89870,);
DFFARX1 I_5127 (I89870,I2683,I89646,I89635,);
nand I_5128 (I89892,I809695,I809704);
and I_5129 (I89909,I89892,I809698);
DFFARX1 I_5130 (I89909,I2683,I89646,I89935,);
DFFARX1 I_5131 (I89935,I2683,I89646,I89952,);
not I_5132 (I89638,I89952);
not I_5133 (I89974,I89935);
nand I_5134 (I89623,I89974,I89813);
nor I_5135 (I90005,I809701,I809704);
not I_5136 (I90022,I90005);
nor I_5137 (I90039,I89974,I90022);
nor I_5138 (I90056,I89680,I90039);
DFFARX1 I_5139 (I90056,I2683,I89646,I89632,);
nor I_5140 (I90087,I89740,I90022);
nor I_5141 (I89620,I89935,I90087);
nor I_5142 (I89629,I89870,I90005);
nor I_5143 (I89617,I89740,I90005);
not I_5144 (I90173,I2690);
DFFARX1 I_5145 (I167027,I2683,I90173,I90199,);
not I_5146 (I90207,I90199);
nand I_5147 (I90224,I167021,I167015);
and I_5148 (I90241,I90224,I167036);
DFFARX1 I_5149 (I90241,I2683,I90173,I90267,);
DFFARX1 I_5150 (I167033,I2683,I90173,I90284,);
and I_5151 (I90292,I90284,I167030);
nor I_5152 (I90309,I90267,I90292);
DFFARX1 I_5153 (I90309,I2683,I90173,I90141,);
nand I_5154 (I90340,I90284,I167030);
nand I_5155 (I90357,I90207,I90340);
not I_5156 (I90153,I90357);
DFFARX1 I_5157 (I167015,I2683,I90173,I90397,);
DFFARX1 I_5158 (I90397,I2683,I90173,I90162,);
nand I_5159 (I90419,I167018,I167018);
and I_5160 (I90436,I90419,I167039);
DFFARX1 I_5161 (I90436,I2683,I90173,I90462,);
DFFARX1 I_5162 (I90462,I2683,I90173,I90479,);
not I_5163 (I90165,I90479);
not I_5164 (I90501,I90462);
nand I_5165 (I90150,I90501,I90340);
nor I_5166 (I90532,I167024,I167018);
not I_5167 (I90549,I90532);
nor I_5168 (I90566,I90501,I90549);
nor I_5169 (I90583,I90207,I90566);
DFFARX1 I_5170 (I90583,I2683,I90173,I90159,);
nor I_5171 (I90614,I90267,I90549);
nor I_5172 (I90147,I90462,I90614);
nor I_5173 (I90156,I90397,I90532);
nor I_5174 (I90144,I90267,I90532);
not I_5175 (I90700,I2690);
DFFARX1 I_5176 (I325252,I2683,I90700,I90726,);
not I_5177 (I90734,I90726);
nand I_5178 (I90751,I325246,I325237);
and I_5179 (I90768,I90751,I325258);
DFFARX1 I_5180 (I90768,I2683,I90700,I90794,);
DFFARX1 I_5181 (I325240,I2683,I90700,I90811,);
and I_5182 (I90819,I90811,I325234);
nor I_5183 (I90836,I90794,I90819);
DFFARX1 I_5184 (I90836,I2683,I90700,I90668,);
nand I_5185 (I90867,I90811,I325234);
nand I_5186 (I90884,I90734,I90867);
not I_5187 (I90680,I90884);
DFFARX1 I_5188 (I325234,I2683,I90700,I90924,);
DFFARX1 I_5189 (I90924,I2683,I90700,I90689,);
nand I_5190 (I90946,I325261,I325243);
and I_5191 (I90963,I90946,I325249);
DFFARX1 I_5192 (I90963,I2683,I90700,I90989,);
DFFARX1 I_5193 (I90989,I2683,I90700,I91006,);
not I_5194 (I90692,I91006);
not I_5195 (I91028,I90989);
nand I_5196 (I90677,I91028,I90867);
nor I_5197 (I91059,I325255,I325243);
not I_5198 (I91076,I91059);
nor I_5199 (I91093,I91028,I91076);
nor I_5200 (I91110,I90734,I91093);
DFFARX1 I_5201 (I91110,I2683,I90700,I90686,);
nor I_5202 (I91141,I90794,I91076);
nor I_5203 (I90674,I90989,I91141);
nor I_5204 (I90683,I90924,I91059);
nor I_5205 (I90671,I90794,I91059);
not I_5206 (I91227,I2690);
DFFARX1 I_5207 (I258570,I2683,I91227,I91253,);
not I_5208 (I91261,I91253);
nand I_5209 (I91278,I258552,I258567);
and I_5210 (I91295,I91278,I258543);
DFFARX1 I_5211 (I91295,I2683,I91227,I91321,);
DFFARX1 I_5212 (I258546,I2683,I91227,I91338,);
and I_5213 (I91346,I91338,I258561);
nor I_5214 (I91363,I91321,I91346);
DFFARX1 I_5215 (I91363,I2683,I91227,I91195,);
nand I_5216 (I91394,I91338,I258561);
nand I_5217 (I91411,I91261,I91394);
not I_5218 (I91207,I91411);
DFFARX1 I_5219 (I258564,I2683,I91227,I91451,);
DFFARX1 I_5220 (I91451,I2683,I91227,I91216,);
nand I_5221 (I91473,I258543,I258555);
and I_5222 (I91490,I91473,I258549);
DFFARX1 I_5223 (I91490,I2683,I91227,I91516,);
DFFARX1 I_5224 (I91516,I2683,I91227,I91533,);
not I_5225 (I91219,I91533);
not I_5226 (I91555,I91516);
nand I_5227 (I91204,I91555,I91394);
nor I_5228 (I91586,I258558,I258555);
not I_5229 (I91603,I91586);
nor I_5230 (I91620,I91555,I91603);
nor I_5231 (I91637,I91261,I91620);
DFFARX1 I_5232 (I91637,I2683,I91227,I91213,);
nor I_5233 (I91668,I91321,I91603);
nor I_5234 (I91201,I91516,I91668);
nor I_5235 (I91210,I91451,I91586);
nor I_5236 (I91198,I91321,I91586);
not I_5237 (I91754,I2690);
DFFARX1 I_5238 (I725814,I2683,I91754,I91780,);
not I_5239 (I91788,I91780);
nand I_5240 (I91805,I725832,I725826);
and I_5241 (I91822,I91805,I725805);
DFFARX1 I_5242 (I91822,I2683,I91754,I91848,);
DFFARX1 I_5243 (I725823,I2683,I91754,I91865,);
and I_5244 (I91873,I91865,I725808);
nor I_5245 (I91890,I91848,I91873);
DFFARX1 I_5246 (I91890,I2683,I91754,I91722,);
nand I_5247 (I91921,I91865,I725808);
nand I_5248 (I91938,I91788,I91921);
not I_5249 (I91734,I91938);
DFFARX1 I_5250 (I725820,I2683,I91754,I91978,);
DFFARX1 I_5251 (I91978,I2683,I91754,I91743,);
nand I_5252 (I92000,I725829,I725817);
and I_5253 (I92017,I92000,I725811);
DFFARX1 I_5254 (I92017,I2683,I91754,I92043,);
DFFARX1 I_5255 (I92043,I2683,I91754,I92060,);
not I_5256 (I91746,I92060);
not I_5257 (I92082,I92043);
nand I_5258 (I91731,I92082,I91921);
nor I_5259 (I92113,I725805,I725817);
not I_5260 (I92130,I92113);
nor I_5261 (I92147,I92082,I92130);
nor I_5262 (I92164,I91788,I92147);
DFFARX1 I_5263 (I92164,I2683,I91754,I91740,);
nor I_5264 (I92195,I91848,I92130);
nor I_5265 (I91728,I92043,I92195);
nor I_5266 (I91737,I91978,I92113);
nor I_5267 (I91725,I91848,I92113);
not I_5268 (I92281,I2690);
DFFARX1 I_5269 (I149772,I2683,I92281,I92307,);
not I_5270 (I92315,I92307);
nand I_5271 (I92332,I149766,I149760);
and I_5272 (I92349,I92332,I149781);
DFFARX1 I_5273 (I92349,I2683,I92281,I92375,);
DFFARX1 I_5274 (I149778,I2683,I92281,I92392,);
and I_5275 (I92400,I92392,I149775);
nor I_5276 (I92417,I92375,I92400);
DFFARX1 I_5277 (I92417,I2683,I92281,I92249,);
nand I_5278 (I92448,I92392,I149775);
nand I_5279 (I92465,I92315,I92448);
not I_5280 (I92261,I92465);
DFFARX1 I_5281 (I149760,I2683,I92281,I92505,);
DFFARX1 I_5282 (I92505,I2683,I92281,I92270,);
nand I_5283 (I92527,I149763,I149763);
and I_5284 (I92544,I92527,I149784);
DFFARX1 I_5285 (I92544,I2683,I92281,I92570,);
DFFARX1 I_5286 (I92570,I2683,I92281,I92587,);
not I_5287 (I92273,I92587);
not I_5288 (I92609,I92570);
nand I_5289 (I92258,I92609,I92448);
nor I_5290 (I92640,I149769,I149763);
not I_5291 (I92657,I92640);
nor I_5292 (I92674,I92609,I92657);
nor I_5293 (I92691,I92315,I92674);
DFFARX1 I_5294 (I92691,I2683,I92281,I92267,);
nor I_5295 (I92722,I92375,I92657);
nor I_5296 (I92255,I92570,I92722);
nor I_5297 (I92264,I92505,I92640);
nor I_5298 (I92252,I92375,I92640);
not I_5299 (I92808,I2690);
DFFARX1 I_5300 (I1082256,I2683,I92808,I92834,);
not I_5301 (I92842,I92834);
nand I_5302 (I92859,I1082250,I1082271);
and I_5303 (I92876,I92859,I1082247);
DFFARX1 I_5304 (I92876,I2683,I92808,I92902,);
DFFARX1 I_5305 (I1082268,I2683,I92808,I92919,);
and I_5306 (I92927,I92919,I1082265);
nor I_5307 (I92944,I92902,I92927);
DFFARX1 I_5308 (I92944,I2683,I92808,I92776,);
nand I_5309 (I92975,I92919,I1082265);
nand I_5310 (I92992,I92842,I92975);
not I_5311 (I92788,I92992);
DFFARX1 I_5312 (I1082253,I2683,I92808,I93032,);
DFFARX1 I_5313 (I93032,I2683,I92808,I92797,);
nand I_5314 (I93054,I1082262,I1082259);
and I_5315 (I93071,I93054,I1082244);
DFFARX1 I_5316 (I93071,I2683,I92808,I93097,);
DFFARX1 I_5317 (I93097,I2683,I92808,I93114,);
not I_5318 (I92800,I93114);
not I_5319 (I93136,I93097);
nand I_5320 (I92785,I93136,I92975);
nor I_5321 (I93167,I1082244,I1082259);
not I_5322 (I93184,I93167);
nor I_5323 (I93201,I93136,I93184);
nor I_5324 (I93218,I92842,I93201);
DFFARX1 I_5325 (I93218,I2683,I92808,I92794,);
nor I_5326 (I93249,I92902,I93184);
nor I_5327 (I92782,I93097,I93249);
nor I_5328 (I92791,I93032,I93167);
nor I_5329 (I92779,I92902,I93167);
not I_5330 (I93335,I2690);
DFFARX1 I_5331 (I621213,I2683,I93335,I93361,);
not I_5332 (I93369,I93361);
nand I_5333 (I93386,I621210,I621225);
and I_5334 (I93403,I93386,I621207);
DFFARX1 I_5335 (I93403,I2683,I93335,I93429,);
DFFARX1 I_5336 (I621204,I2683,I93335,I93446,);
and I_5337 (I93454,I93446,I621204);
nor I_5338 (I93471,I93429,I93454);
DFFARX1 I_5339 (I93471,I2683,I93335,I93303,);
nand I_5340 (I93502,I93446,I621204);
nand I_5341 (I93519,I93369,I93502);
not I_5342 (I93315,I93519);
DFFARX1 I_5343 (I621207,I2683,I93335,I93559,);
DFFARX1 I_5344 (I93559,I2683,I93335,I93324,);
nand I_5345 (I93581,I621219,I621210);
and I_5346 (I93598,I93581,I621222);
DFFARX1 I_5347 (I93598,I2683,I93335,I93624,);
DFFARX1 I_5348 (I93624,I2683,I93335,I93641,);
not I_5349 (I93327,I93641);
not I_5350 (I93663,I93624);
nand I_5351 (I93312,I93663,I93502);
nor I_5352 (I93694,I621216,I621210);
not I_5353 (I93711,I93694);
nor I_5354 (I93728,I93663,I93711);
nor I_5355 (I93745,I93369,I93728);
DFFARX1 I_5356 (I93745,I2683,I93335,I93321,);
nor I_5357 (I93776,I93429,I93711);
nor I_5358 (I93309,I93624,I93776);
nor I_5359 (I93318,I93559,I93694);
nor I_5360 (I93306,I93429,I93694);
not I_5361 (I93862,I2690);
DFFARX1 I_5362 (I1051911,I2683,I93862,I93888,);
not I_5363 (I93896,I93888);
nand I_5364 (I93913,I1051905,I1051926);
and I_5365 (I93930,I93913,I1051902);
DFFARX1 I_5366 (I93930,I2683,I93862,I93956,);
DFFARX1 I_5367 (I1051923,I2683,I93862,I93973,);
and I_5368 (I93981,I93973,I1051920);
nor I_5369 (I93998,I93956,I93981);
DFFARX1 I_5370 (I93998,I2683,I93862,I93830,);
nand I_5371 (I94029,I93973,I1051920);
nand I_5372 (I94046,I93896,I94029);
not I_5373 (I93842,I94046);
DFFARX1 I_5374 (I1051908,I2683,I93862,I94086,);
DFFARX1 I_5375 (I94086,I2683,I93862,I93851,);
nand I_5376 (I94108,I1051917,I1051914);
and I_5377 (I94125,I94108,I1051899);
DFFARX1 I_5378 (I94125,I2683,I93862,I94151,);
DFFARX1 I_5379 (I94151,I2683,I93862,I94168,);
not I_5380 (I93854,I94168);
not I_5381 (I94190,I94151);
nand I_5382 (I93839,I94190,I94029);
nor I_5383 (I94221,I1051899,I1051914);
not I_5384 (I94238,I94221);
nor I_5385 (I94255,I94190,I94238);
nor I_5386 (I94272,I93896,I94255);
DFFARX1 I_5387 (I94272,I2683,I93862,I93848,);
nor I_5388 (I94303,I93956,I94238);
nor I_5389 (I93836,I94151,I94303);
nor I_5390 (I93845,I94086,I94221);
nor I_5391 (I93833,I93956,I94221);
not I_5392 (I94389,I2690);
DFFARX1 I_5393 (I219045,I2683,I94389,I94415,);
not I_5394 (I94423,I94415);
nand I_5395 (I94440,I219027,I219042);
and I_5396 (I94457,I94440,I219018);
DFFARX1 I_5397 (I94457,I2683,I94389,I94483,);
DFFARX1 I_5398 (I219021,I2683,I94389,I94500,);
and I_5399 (I94508,I94500,I219036);
nor I_5400 (I94525,I94483,I94508);
DFFARX1 I_5401 (I94525,I2683,I94389,I94357,);
nand I_5402 (I94556,I94500,I219036);
nand I_5403 (I94573,I94423,I94556);
not I_5404 (I94369,I94573);
DFFARX1 I_5405 (I219039,I2683,I94389,I94613,);
DFFARX1 I_5406 (I94613,I2683,I94389,I94378,);
nand I_5407 (I94635,I219018,I219030);
and I_5408 (I94652,I94635,I219024);
DFFARX1 I_5409 (I94652,I2683,I94389,I94678,);
DFFARX1 I_5410 (I94678,I2683,I94389,I94695,);
not I_5411 (I94381,I94695);
not I_5412 (I94717,I94678);
nand I_5413 (I94366,I94717,I94556);
nor I_5414 (I94748,I219033,I219030);
not I_5415 (I94765,I94748);
nor I_5416 (I94782,I94717,I94765);
nor I_5417 (I94799,I94423,I94782);
DFFARX1 I_5418 (I94799,I2683,I94389,I94375,);
nor I_5419 (I94830,I94483,I94765);
nor I_5420 (I94363,I94678,I94830);
nor I_5421 (I94372,I94613,I94748);
nor I_5422 (I94360,I94483,I94748);
not I_5423 (I94916,I2690);
DFFARX1 I_5424 (I215883,I2683,I94916,I94942,);
not I_5425 (I94950,I94942);
nand I_5426 (I94967,I215865,I215880);
and I_5427 (I94984,I94967,I215856);
DFFARX1 I_5428 (I94984,I2683,I94916,I95010,);
DFFARX1 I_5429 (I215859,I2683,I94916,I95027,);
and I_5430 (I95035,I95027,I215874);
nor I_5431 (I95052,I95010,I95035);
DFFARX1 I_5432 (I95052,I2683,I94916,I94884,);
nand I_5433 (I95083,I95027,I215874);
nand I_5434 (I95100,I94950,I95083);
not I_5435 (I94896,I95100);
DFFARX1 I_5436 (I215877,I2683,I94916,I95140,);
DFFARX1 I_5437 (I95140,I2683,I94916,I94905,);
nand I_5438 (I95162,I215856,I215868);
and I_5439 (I95179,I95162,I215862);
DFFARX1 I_5440 (I95179,I2683,I94916,I95205,);
DFFARX1 I_5441 (I95205,I2683,I94916,I95222,);
not I_5442 (I94908,I95222);
not I_5443 (I95244,I95205);
nand I_5444 (I94893,I95244,I95083);
nor I_5445 (I95275,I215871,I215868);
not I_5446 (I95292,I95275);
nor I_5447 (I95309,I95244,I95292);
nor I_5448 (I95326,I94950,I95309);
DFFARX1 I_5449 (I95326,I2683,I94916,I94902,);
nor I_5450 (I95357,I95010,I95292);
nor I_5451 (I94890,I95205,I95357);
nor I_5452 (I94899,I95140,I95275);
nor I_5453 (I94887,I95010,I95275);
not I_5454 (I95443,I2690);
DFFARX1 I_5455 (I407415,I2683,I95443,I95469,);
not I_5456 (I95477,I95469);
nand I_5457 (I95494,I407436,I407430);
and I_5458 (I95511,I95494,I407412);
DFFARX1 I_5459 (I95511,I2683,I95443,I95537,);
DFFARX1 I_5460 (I407415,I2683,I95443,I95554,);
and I_5461 (I95562,I95554,I407424);
nor I_5462 (I95579,I95537,I95562);
DFFARX1 I_5463 (I95579,I2683,I95443,I95411,);
nand I_5464 (I95610,I95554,I407424);
nand I_5465 (I95627,I95477,I95610);
not I_5466 (I95423,I95627);
DFFARX1 I_5467 (I407421,I2683,I95443,I95667,);
DFFARX1 I_5468 (I95667,I2683,I95443,I95432,);
nand I_5469 (I95689,I407427,I407418);
and I_5470 (I95706,I95689,I407412);
DFFARX1 I_5471 (I95706,I2683,I95443,I95732,);
DFFARX1 I_5472 (I95732,I2683,I95443,I95749,);
not I_5473 (I95435,I95749);
not I_5474 (I95771,I95732);
nand I_5475 (I95420,I95771,I95610);
nor I_5476 (I95802,I407433,I407418);
not I_5477 (I95819,I95802);
nor I_5478 (I95836,I95771,I95819);
nor I_5479 (I95853,I95477,I95836);
DFFARX1 I_5480 (I95853,I2683,I95443,I95429,);
nor I_5481 (I95884,I95537,I95819);
nor I_5482 (I95417,I95732,I95884);
nor I_5483 (I95426,I95667,I95802);
nor I_5484 (I95414,I95537,I95802);
not I_5485 (I95970,I2690);
DFFARX1 I_5486 (I938600,I2683,I95970,I95996,);
not I_5487 (I96004,I95996);
nand I_5488 (I96021,I938615,I938594);
and I_5489 (I96038,I96021,I938597);
DFFARX1 I_5490 (I96038,I2683,I95970,I96064,);
DFFARX1 I_5491 (I938618,I2683,I95970,I96081,);
and I_5492 (I96089,I96081,I938597);
nor I_5493 (I96106,I96064,I96089);
DFFARX1 I_5494 (I96106,I2683,I95970,I95938,);
nand I_5495 (I96137,I96081,I938597);
nand I_5496 (I96154,I96004,I96137);
not I_5497 (I95950,I96154);
DFFARX1 I_5498 (I938594,I2683,I95970,I96194,);
DFFARX1 I_5499 (I96194,I2683,I95970,I95959,);
nand I_5500 (I96216,I938606,I938603);
and I_5501 (I96233,I96216,I938609);
DFFARX1 I_5502 (I96233,I2683,I95970,I96259,);
DFFARX1 I_5503 (I96259,I2683,I95970,I96276,);
not I_5504 (I95962,I96276);
not I_5505 (I96298,I96259);
nand I_5506 (I95947,I96298,I96137);
nor I_5507 (I96329,I938612,I938603);
not I_5508 (I96346,I96329);
nor I_5509 (I96363,I96298,I96346);
nor I_5510 (I96380,I96004,I96363);
DFFARX1 I_5511 (I96380,I2683,I95970,I95956,);
nor I_5512 (I96411,I96064,I96346);
nor I_5513 (I95944,I96259,I96411);
nor I_5514 (I95953,I96194,I96329);
nor I_5515 (I95941,I96064,I96329);
not I_5516 (I96497,I2690);
DFFARX1 I_5517 (I193207,I2683,I96497,I96523,);
not I_5518 (I96531,I96523);
nand I_5519 (I96548,I193201,I193195);
and I_5520 (I96565,I96548,I193216);
DFFARX1 I_5521 (I96565,I2683,I96497,I96591,);
DFFARX1 I_5522 (I193213,I2683,I96497,I96608,);
and I_5523 (I96616,I96608,I193210);
nor I_5524 (I96633,I96591,I96616);
DFFARX1 I_5525 (I96633,I2683,I96497,I96465,);
nand I_5526 (I96664,I96608,I193210);
nand I_5527 (I96681,I96531,I96664);
not I_5528 (I96477,I96681);
DFFARX1 I_5529 (I193195,I2683,I96497,I96721,);
DFFARX1 I_5530 (I96721,I2683,I96497,I96486,);
nand I_5531 (I96743,I193198,I193198);
and I_5532 (I96760,I96743,I193219);
DFFARX1 I_5533 (I96760,I2683,I96497,I96786,);
DFFARX1 I_5534 (I96786,I2683,I96497,I96803,);
not I_5535 (I96489,I96803);
not I_5536 (I96825,I96786);
nand I_5537 (I96474,I96825,I96664);
nor I_5538 (I96856,I193204,I193198);
not I_5539 (I96873,I96856);
nor I_5540 (I96890,I96825,I96873);
nor I_5541 (I96907,I96531,I96890);
DFFARX1 I_5542 (I96907,I2683,I96497,I96483,);
nor I_5543 (I96938,I96591,I96873);
nor I_5544 (I96471,I96786,I96938);
nor I_5545 (I96480,I96721,I96856);
nor I_5546 (I96468,I96591,I96856);
not I_5547 (I97024,I2690);
DFFARX1 I_5548 (I983684,I2683,I97024,I97050,);
not I_5549 (I97058,I97050);
nand I_5550 (I97075,I983678,I983699);
and I_5551 (I97092,I97075,I983690);
DFFARX1 I_5552 (I97092,I2683,I97024,I97118,);
DFFARX1 I_5553 (I983681,I2683,I97024,I97135,);
and I_5554 (I97143,I97135,I983693);
nor I_5555 (I97160,I97118,I97143);
DFFARX1 I_5556 (I97160,I2683,I97024,I96992,);
nand I_5557 (I97191,I97135,I983693);
nand I_5558 (I97208,I97058,I97191);
not I_5559 (I97004,I97208);
DFFARX1 I_5560 (I983681,I2683,I97024,I97248,);
DFFARX1 I_5561 (I97248,I2683,I97024,I97013,);
nand I_5562 (I97270,I983702,I983687);
and I_5563 (I97287,I97270,I983678);
DFFARX1 I_5564 (I97287,I2683,I97024,I97313,);
DFFARX1 I_5565 (I97313,I2683,I97024,I97330,);
not I_5566 (I97016,I97330);
not I_5567 (I97352,I97313);
nand I_5568 (I97001,I97352,I97191);
nor I_5569 (I97383,I983696,I983687);
not I_5570 (I97400,I97383);
nor I_5571 (I97417,I97352,I97400);
nor I_5572 (I97434,I97058,I97417);
DFFARX1 I_5573 (I97434,I2683,I97024,I97010,);
nor I_5574 (I97465,I97118,I97400);
nor I_5575 (I96998,I97313,I97465);
nor I_5576 (I97007,I97248,I97383);
nor I_5577 (I96995,I97118,I97383);
not I_5578 (I97551,I2690);
DFFARX1 I_5579 (I515646,I2683,I97551,I97577,);
not I_5580 (I97585,I97577);
nand I_5581 (I97602,I515637,I515655);
and I_5582 (I97619,I97602,I515634);
DFFARX1 I_5583 (I97619,I2683,I97551,I97645,);
DFFARX1 I_5584 (I515637,I2683,I97551,I97662,);
and I_5585 (I97670,I97662,I515640);
nor I_5586 (I97687,I97645,I97670);
DFFARX1 I_5587 (I97687,I2683,I97551,I97519,);
nand I_5588 (I97718,I97662,I515640);
nand I_5589 (I97735,I97585,I97718);
not I_5590 (I97531,I97735);
DFFARX1 I_5591 (I515634,I2683,I97551,I97775,);
DFFARX1 I_5592 (I97775,I2683,I97551,I97540,);
nand I_5593 (I97797,I515652,I515643);
and I_5594 (I97814,I97797,I515658);
DFFARX1 I_5595 (I97814,I2683,I97551,I97840,);
DFFARX1 I_5596 (I97840,I2683,I97551,I97857,);
not I_5597 (I97543,I97857);
not I_5598 (I97879,I97840);
nand I_5599 (I97528,I97879,I97718);
nor I_5600 (I97910,I515649,I515643);
not I_5601 (I97927,I97910);
nor I_5602 (I97944,I97879,I97927);
nor I_5603 (I97961,I97585,I97944);
DFFARX1 I_5604 (I97961,I2683,I97551,I97537,);
nor I_5605 (I97992,I97645,I97927);
nor I_5606 (I97525,I97840,I97992);
nor I_5607 (I97534,I97775,I97910);
nor I_5608 (I97522,I97645,I97910);
not I_5609 (I98078,I2690);
DFFARX1 I_5610 (I863460,I2683,I98078,I98104,);
not I_5611 (I98112,I98104);
nand I_5612 (I98129,I863475,I863454);
and I_5613 (I98146,I98129,I863457);
DFFARX1 I_5614 (I98146,I2683,I98078,I98172,);
DFFARX1 I_5615 (I863478,I2683,I98078,I98189,);
and I_5616 (I98197,I98189,I863457);
nor I_5617 (I98214,I98172,I98197);
DFFARX1 I_5618 (I98214,I2683,I98078,I98046,);
nand I_5619 (I98245,I98189,I863457);
nand I_5620 (I98262,I98112,I98245);
not I_5621 (I98058,I98262);
DFFARX1 I_5622 (I863454,I2683,I98078,I98302,);
DFFARX1 I_5623 (I98302,I2683,I98078,I98067,);
nand I_5624 (I98324,I863466,I863463);
and I_5625 (I98341,I98324,I863469);
DFFARX1 I_5626 (I98341,I2683,I98078,I98367,);
DFFARX1 I_5627 (I98367,I2683,I98078,I98384,);
not I_5628 (I98070,I98384);
not I_5629 (I98406,I98367);
nand I_5630 (I98055,I98406,I98245);
nor I_5631 (I98437,I863472,I863463);
not I_5632 (I98454,I98437);
nor I_5633 (I98471,I98406,I98454);
nor I_5634 (I98488,I98112,I98471);
DFFARX1 I_5635 (I98488,I2683,I98078,I98064,);
nor I_5636 (I98519,I98172,I98454);
nor I_5637 (I98052,I98367,I98519);
nor I_5638 (I98061,I98302,I98437);
nor I_5639 (I98049,I98172,I98437);
not I_5640 (I98605,I2690);
DFFARX1 I_5641 (I421695,I2683,I98605,I98631,);
not I_5642 (I98639,I98631);
nand I_5643 (I98656,I421716,I421710);
and I_5644 (I98673,I98656,I421692);
DFFARX1 I_5645 (I98673,I2683,I98605,I98699,);
DFFARX1 I_5646 (I421695,I2683,I98605,I98716,);
and I_5647 (I98724,I98716,I421704);
nor I_5648 (I98741,I98699,I98724);
DFFARX1 I_5649 (I98741,I2683,I98605,I98573,);
nand I_5650 (I98772,I98716,I421704);
nand I_5651 (I98789,I98639,I98772);
not I_5652 (I98585,I98789);
DFFARX1 I_5653 (I421701,I2683,I98605,I98829,);
DFFARX1 I_5654 (I98829,I2683,I98605,I98594,);
nand I_5655 (I98851,I421707,I421698);
and I_5656 (I98868,I98851,I421692);
DFFARX1 I_5657 (I98868,I2683,I98605,I98894,);
DFFARX1 I_5658 (I98894,I2683,I98605,I98911,);
not I_5659 (I98597,I98911);
not I_5660 (I98933,I98894);
nand I_5661 (I98582,I98933,I98772);
nor I_5662 (I98964,I421713,I421698);
not I_5663 (I98981,I98964);
nor I_5664 (I98998,I98933,I98981);
nor I_5665 (I99015,I98639,I98998);
DFFARX1 I_5666 (I99015,I2683,I98605,I98591,);
nor I_5667 (I99046,I98699,I98981);
nor I_5668 (I98579,I98894,I99046);
nor I_5669 (I98588,I98829,I98964);
nor I_5670 (I98576,I98699,I98964);
not I_5671 (I99132,I2690);
DFFARX1 I_5672 (I549748,I2683,I99132,I99158,);
not I_5673 (I99166,I99158);
nand I_5674 (I99183,I549739,I549757);
and I_5675 (I99200,I99183,I549736);
DFFARX1 I_5676 (I99200,I2683,I99132,I99226,);
DFFARX1 I_5677 (I549739,I2683,I99132,I99243,);
and I_5678 (I99251,I99243,I549742);
nor I_5679 (I99268,I99226,I99251);
DFFARX1 I_5680 (I99268,I2683,I99132,I99100,);
nand I_5681 (I99299,I99243,I549742);
nand I_5682 (I99316,I99166,I99299);
not I_5683 (I99112,I99316);
DFFARX1 I_5684 (I549736,I2683,I99132,I99356,);
DFFARX1 I_5685 (I99356,I2683,I99132,I99121,);
nand I_5686 (I99378,I549754,I549745);
and I_5687 (I99395,I99378,I549760);
DFFARX1 I_5688 (I99395,I2683,I99132,I99421,);
DFFARX1 I_5689 (I99421,I2683,I99132,I99438,);
not I_5690 (I99124,I99438);
not I_5691 (I99460,I99421);
nand I_5692 (I99109,I99460,I99299);
nor I_5693 (I99491,I549751,I549745);
not I_5694 (I99508,I99491);
nor I_5695 (I99525,I99460,I99508);
nor I_5696 (I99542,I99166,I99525);
DFFARX1 I_5697 (I99542,I2683,I99132,I99118,);
nor I_5698 (I99573,I99226,I99508);
nor I_5699 (I99106,I99421,I99573);
nor I_5700 (I99115,I99356,I99491);
nor I_5701 (I99103,I99226,I99491);
not I_5702 (I99659,I2690);
DFFARX1 I_5703 (I32195,I2683,I99659,I99685,);
not I_5704 (I99693,I99685);
nand I_5705 (I99710,I32183,I32189);
and I_5706 (I99727,I99710,I32192);
DFFARX1 I_5707 (I99727,I2683,I99659,I99753,);
DFFARX1 I_5708 (I32174,I2683,I99659,I99770,);
and I_5709 (I99778,I99770,I32180);
nor I_5710 (I99795,I99753,I99778);
DFFARX1 I_5711 (I99795,I2683,I99659,I99627,);
nand I_5712 (I99826,I99770,I32180);
nand I_5713 (I99843,I99693,I99826);
not I_5714 (I99639,I99843);
DFFARX1 I_5715 (I32174,I2683,I99659,I99883,);
DFFARX1 I_5716 (I99883,I2683,I99659,I99648,);
nand I_5717 (I99905,I32177,I32171);
and I_5718 (I99922,I99905,I32186);
DFFARX1 I_5719 (I99922,I2683,I99659,I99948,);
DFFARX1 I_5720 (I99948,I2683,I99659,I99965,);
not I_5721 (I99651,I99965);
not I_5722 (I99987,I99948);
nand I_5723 (I99636,I99987,I99826);
nor I_5724 (I100018,I32171,I32171);
not I_5725 (I100035,I100018);
nor I_5726 (I100052,I99987,I100035);
nor I_5727 (I100069,I99693,I100052);
DFFARX1 I_5728 (I100069,I2683,I99659,I99645,);
nor I_5729 (I100100,I99753,I100035);
nor I_5730 (I99633,I99948,I100100);
nor I_5731 (I99642,I99883,I100018);
nor I_5732 (I99630,I99753,I100018);
not I_5733 (I100186,I2690);
DFFARX1 I_5734 (I599456,I2683,I100186,I100212,);
not I_5735 (I100220,I100212);
nand I_5736 (I100237,I599447,I599465);
and I_5737 (I100254,I100237,I599444);
DFFARX1 I_5738 (I100254,I2683,I100186,I100280,);
DFFARX1 I_5739 (I599447,I2683,I100186,I100297,);
and I_5740 (I100305,I100297,I599450);
nor I_5741 (I100322,I100280,I100305);
DFFARX1 I_5742 (I100322,I2683,I100186,I100154,);
nand I_5743 (I100353,I100297,I599450);
nand I_5744 (I100370,I100220,I100353);
not I_5745 (I100166,I100370);
DFFARX1 I_5746 (I599444,I2683,I100186,I100410,);
DFFARX1 I_5747 (I100410,I2683,I100186,I100175,);
nand I_5748 (I100432,I599462,I599453);
and I_5749 (I100449,I100432,I599468);
DFFARX1 I_5750 (I100449,I2683,I100186,I100475,);
DFFARX1 I_5751 (I100475,I2683,I100186,I100492,);
not I_5752 (I100178,I100492);
not I_5753 (I100514,I100475);
nand I_5754 (I100163,I100514,I100353);
nor I_5755 (I100545,I599459,I599453);
not I_5756 (I100562,I100545);
nor I_5757 (I100579,I100514,I100562);
nor I_5758 (I100596,I100220,I100579);
DFFARX1 I_5759 (I100596,I2683,I100186,I100172,);
nor I_5760 (I100627,I100280,I100562);
nor I_5761 (I100160,I100475,I100627);
nor I_5762 (I100169,I100410,I100545);
nor I_5763 (I100157,I100280,I100545);
not I_5764 (I100713,I2690);
DFFARX1 I_5765 (I1092371,I2683,I100713,I100739,);
not I_5766 (I100747,I100739);
nand I_5767 (I100764,I1092365,I1092386);
and I_5768 (I100781,I100764,I1092362);
DFFARX1 I_5769 (I100781,I2683,I100713,I100807,);
DFFARX1 I_5770 (I1092383,I2683,I100713,I100824,);
and I_5771 (I100832,I100824,I1092380);
nor I_5772 (I100849,I100807,I100832);
DFFARX1 I_5773 (I100849,I2683,I100713,I100681,);
nand I_5774 (I100880,I100824,I1092380);
nand I_5775 (I100897,I100747,I100880);
not I_5776 (I100693,I100897);
DFFARX1 I_5777 (I1092368,I2683,I100713,I100937,);
DFFARX1 I_5778 (I100937,I2683,I100713,I100702,);
nand I_5779 (I100959,I1092377,I1092374);
and I_5780 (I100976,I100959,I1092359);
DFFARX1 I_5781 (I100976,I2683,I100713,I101002,);
DFFARX1 I_5782 (I101002,I2683,I100713,I101019,);
not I_5783 (I100705,I101019);
not I_5784 (I101041,I101002);
nand I_5785 (I100690,I101041,I100880);
nor I_5786 (I101072,I1092359,I1092374);
not I_5787 (I101089,I101072);
nor I_5788 (I101106,I101041,I101089);
nor I_5789 (I101123,I100747,I101106);
DFFARX1 I_5790 (I101123,I2683,I100713,I100699,);
nor I_5791 (I101154,I100807,I101089);
nor I_5792 (I100687,I101002,I101154);
nor I_5793 (I100696,I100937,I101072);
nor I_5794 (I100684,I100807,I101072);
not I_5795 (I101240,I2690);
DFFARX1 I_5796 (I903342,I2683,I101240,I101266,);
not I_5797 (I101274,I101266);
nand I_5798 (I101291,I903357,I903336);
and I_5799 (I101308,I101291,I903339);
DFFARX1 I_5800 (I101308,I2683,I101240,I101334,);
DFFARX1 I_5801 (I903360,I2683,I101240,I101351,);
and I_5802 (I101359,I101351,I903339);
nor I_5803 (I101376,I101334,I101359);
DFFARX1 I_5804 (I101376,I2683,I101240,I101208,);
nand I_5805 (I101407,I101351,I903339);
nand I_5806 (I101424,I101274,I101407);
not I_5807 (I101220,I101424);
DFFARX1 I_5808 (I903336,I2683,I101240,I101464,);
DFFARX1 I_5809 (I101464,I2683,I101240,I101229,);
nand I_5810 (I101486,I903348,I903345);
and I_5811 (I101503,I101486,I903351);
DFFARX1 I_5812 (I101503,I2683,I101240,I101529,);
DFFARX1 I_5813 (I101529,I2683,I101240,I101546,);
not I_5814 (I101232,I101546);
not I_5815 (I101568,I101529);
nand I_5816 (I101217,I101568,I101407);
nor I_5817 (I101599,I903354,I903345);
not I_5818 (I101616,I101599);
nor I_5819 (I101633,I101568,I101616);
nor I_5820 (I101650,I101274,I101633);
DFFARX1 I_5821 (I101650,I2683,I101240,I101226,);
nor I_5822 (I101681,I101334,I101616);
nor I_5823 (I101214,I101529,I101681);
nor I_5824 (I101223,I101464,I101599);
nor I_5825 (I101211,I101334,I101599);
not I_5826 (I101767,I2690);
DFFARX1 I_5827 (I1086421,I2683,I101767,I101793,);
not I_5828 (I101801,I101793);
nand I_5829 (I101818,I1086415,I1086436);
and I_5830 (I101835,I101818,I1086412);
DFFARX1 I_5831 (I101835,I2683,I101767,I101861,);
DFFARX1 I_5832 (I1086433,I2683,I101767,I101878,);
and I_5833 (I101886,I101878,I1086430);
nor I_5834 (I101903,I101861,I101886);
DFFARX1 I_5835 (I101903,I2683,I101767,I101735,);
nand I_5836 (I101934,I101878,I1086430);
nand I_5837 (I101951,I101801,I101934);
not I_5838 (I101747,I101951);
DFFARX1 I_5839 (I1086418,I2683,I101767,I101991,);
DFFARX1 I_5840 (I101991,I2683,I101767,I101756,);
nand I_5841 (I102013,I1086427,I1086424);
and I_5842 (I102030,I102013,I1086409);
DFFARX1 I_5843 (I102030,I2683,I101767,I102056,);
DFFARX1 I_5844 (I102056,I2683,I101767,I102073,);
not I_5845 (I101759,I102073);
not I_5846 (I102095,I102056);
nand I_5847 (I101744,I102095,I101934);
nor I_5848 (I102126,I1086409,I1086424);
not I_5849 (I102143,I102126);
nor I_5850 (I102160,I102095,I102143);
nor I_5851 (I102177,I101801,I102160);
DFFARX1 I_5852 (I102177,I2683,I101767,I101753,);
nor I_5853 (I102208,I101861,I102143);
nor I_5854 (I101741,I102056,I102208);
nor I_5855 (I101750,I101991,I102126);
nor I_5856 (I101738,I101861,I102126);
not I_5857 (I102294,I2690);
DFFARX1 I_5858 (I1045961,I2683,I102294,I102320,);
not I_5859 (I102328,I102320);
nand I_5860 (I102345,I1045955,I1045976);
and I_5861 (I102362,I102345,I1045952);
DFFARX1 I_5862 (I102362,I2683,I102294,I102388,);
DFFARX1 I_5863 (I1045973,I2683,I102294,I102405,);
and I_5864 (I102413,I102405,I1045970);
nor I_5865 (I102430,I102388,I102413);
DFFARX1 I_5866 (I102430,I2683,I102294,I102262,);
nand I_5867 (I102461,I102405,I1045970);
nand I_5868 (I102478,I102328,I102461);
not I_5869 (I102274,I102478);
DFFARX1 I_5870 (I1045958,I2683,I102294,I102518,);
DFFARX1 I_5871 (I102518,I2683,I102294,I102283,);
nand I_5872 (I102540,I1045967,I1045964);
and I_5873 (I102557,I102540,I1045949);
DFFARX1 I_5874 (I102557,I2683,I102294,I102583,);
DFFARX1 I_5875 (I102583,I2683,I102294,I102600,);
not I_5876 (I102286,I102600);
not I_5877 (I102622,I102583);
nand I_5878 (I102271,I102622,I102461);
nor I_5879 (I102653,I1045949,I1045964);
not I_5880 (I102670,I102653);
nor I_5881 (I102687,I102622,I102670);
nor I_5882 (I102704,I102328,I102687);
DFFARX1 I_5883 (I102704,I2683,I102294,I102280,);
nor I_5884 (I102735,I102388,I102670);
nor I_5885 (I102268,I102583,I102735);
nor I_5886 (I102277,I102518,I102653);
nor I_5887 (I102265,I102388,I102653);
not I_5888 (I102821,I2690);
DFFARX1 I_5889 (I467091,I2683,I102821,I102847,);
not I_5890 (I102855,I102847);
nand I_5891 (I102872,I467103,I467088);
and I_5892 (I102889,I102872,I467082);
DFFARX1 I_5893 (I102889,I2683,I102821,I102915,);
DFFARX1 I_5894 (I467097,I2683,I102821,I102932,);
and I_5895 (I102940,I102932,I467085);
nor I_5896 (I102957,I102915,I102940);
DFFARX1 I_5897 (I102957,I2683,I102821,I102789,);
nand I_5898 (I102988,I102932,I467085);
nand I_5899 (I103005,I102855,I102988);
not I_5900 (I102801,I103005);
DFFARX1 I_5901 (I467094,I2683,I102821,I103045,);
DFFARX1 I_5902 (I103045,I2683,I102821,I102810,);
nand I_5903 (I103067,I467100,I467106);
and I_5904 (I103084,I103067,I467082);
DFFARX1 I_5905 (I103084,I2683,I102821,I103110,);
DFFARX1 I_5906 (I103110,I2683,I102821,I103127,);
not I_5907 (I102813,I103127);
not I_5908 (I103149,I103110);
nand I_5909 (I102798,I103149,I102988);
nor I_5910 (I103180,I467085,I467106);
not I_5911 (I103197,I103180);
nor I_5912 (I103214,I103149,I103197);
nor I_5913 (I103231,I102855,I103214);
DFFARX1 I_5914 (I103231,I2683,I102821,I102807,);
nor I_5915 (I103262,I102915,I103197);
nor I_5916 (I102795,I103110,I103262);
nor I_5917 (I102804,I103045,I103180);
nor I_5918 (I102792,I102915,I103180);
not I_5919 (I103348,I2690);
DFFARX1 I_5920 (I178927,I2683,I103348,I103374,);
not I_5921 (I103382,I103374);
nand I_5922 (I103399,I178921,I178915);
and I_5923 (I103416,I103399,I178936);
DFFARX1 I_5924 (I103416,I2683,I103348,I103442,);
DFFARX1 I_5925 (I178933,I2683,I103348,I103459,);
and I_5926 (I103467,I103459,I178930);
nor I_5927 (I103484,I103442,I103467);
DFFARX1 I_5928 (I103484,I2683,I103348,I103316,);
nand I_5929 (I103515,I103459,I178930);
nand I_5930 (I103532,I103382,I103515);
not I_5931 (I103328,I103532);
DFFARX1 I_5932 (I178915,I2683,I103348,I103572,);
DFFARX1 I_5933 (I103572,I2683,I103348,I103337,);
nand I_5934 (I103594,I178918,I178918);
and I_5935 (I103611,I103594,I178939);
DFFARX1 I_5936 (I103611,I2683,I103348,I103637,);
DFFARX1 I_5937 (I103637,I2683,I103348,I103654,);
not I_5938 (I103340,I103654);
not I_5939 (I103676,I103637);
nand I_5940 (I103325,I103676,I103515);
nor I_5941 (I103707,I178924,I178918);
not I_5942 (I103724,I103707);
nor I_5943 (I103741,I103676,I103724);
nor I_5944 (I103758,I103382,I103741);
DFFARX1 I_5945 (I103758,I2683,I103348,I103334,);
nor I_5946 (I103789,I103442,I103724);
nor I_5947 (I103322,I103637,I103789);
nor I_5948 (I103331,I103572,I103707);
nor I_5949 (I103319,I103442,I103707);
not I_5950 (I103875,I2690);
DFFARX1 I_5951 (I696574,I2683,I103875,I103901,);
not I_5952 (I103909,I103901);
nand I_5953 (I103926,I696571,I696586);
and I_5954 (I103943,I103926,I696568);
DFFARX1 I_5955 (I103943,I2683,I103875,I103969,);
DFFARX1 I_5956 (I696565,I2683,I103875,I103986,);
and I_5957 (I103994,I103986,I696565);
nor I_5958 (I104011,I103969,I103994);
DFFARX1 I_5959 (I104011,I2683,I103875,I103843,);
nand I_5960 (I104042,I103986,I696565);
nand I_5961 (I104059,I103909,I104042);
not I_5962 (I103855,I104059);
DFFARX1 I_5963 (I696568,I2683,I103875,I104099,);
DFFARX1 I_5964 (I104099,I2683,I103875,I103864,);
nand I_5965 (I104121,I696580,I696571);
and I_5966 (I104138,I104121,I696583);
DFFARX1 I_5967 (I104138,I2683,I103875,I104164,);
DFFARX1 I_5968 (I104164,I2683,I103875,I104181,);
not I_5969 (I103867,I104181);
not I_5970 (I104203,I104164);
nand I_5971 (I103852,I104203,I104042);
nor I_5972 (I104234,I696577,I696571);
not I_5973 (I104251,I104234);
nor I_5974 (I104268,I104203,I104251);
nor I_5975 (I104285,I103909,I104268);
DFFARX1 I_5976 (I104285,I2683,I103875,I103861,);
nor I_5977 (I104316,I103969,I104251);
nor I_5978 (I103849,I104164,I104316);
nor I_5979 (I103858,I104099,I104234);
nor I_5980 (I103846,I103969,I104234);
not I_5981 (I104402,I2690);
DFFARX1 I_5982 (I18493,I2683,I104402,I104428,);
not I_5983 (I104436,I104428);
nand I_5984 (I104453,I18481,I18487);
and I_5985 (I104470,I104453,I18490);
DFFARX1 I_5986 (I104470,I2683,I104402,I104496,);
DFFARX1 I_5987 (I18472,I2683,I104402,I104513,);
and I_5988 (I104521,I104513,I18478);
nor I_5989 (I104538,I104496,I104521);
DFFARX1 I_5990 (I104538,I2683,I104402,I104370,);
nand I_5991 (I104569,I104513,I18478);
nand I_5992 (I104586,I104436,I104569);
not I_5993 (I104382,I104586);
DFFARX1 I_5994 (I18472,I2683,I104402,I104626,);
DFFARX1 I_5995 (I104626,I2683,I104402,I104391,);
nand I_5996 (I104648,I18475,I18469);
and I_5997 (I104665,I104648,I18484);
DFFARX1 I_5998 (I104665,I2683,I104402,I104691,);
DFFARX1 I_5999 (I104691,I2683,I104402,I104708,);
not I_6000 (I104394,I104708);
not I_6001 (I104730,I104691);
nand I_6002 (I104379,I104730,I104569);
nor I_6003 (I104761,I18469,I18469);
not I_6004 (I104778,I104761);
nor I_6005 (I104795,I104730,I104778);
nor I_6006 (I104812,I104436,I104795);
DFFARX1 I_6007 (I104812,I2683,I104402,I104388,);
nor I_6008 (I104843,I104496,I104778);
nor I_6009 (I104376,I104691,I104843);
nor I_6010 (I104385,I104626,I104761);
nor I_6011 (I104373,I104496,I104761);
not I_6012 (I104929,I2690);
DFFARX1 I_6013 (I1026552,I2683,I104929,I104955,);
not I_6014 (I104963,I104955);
nand I_6015 (I104980,I1026558,I1026576);
and I_6016 (I104997,I104980,I1026573);
DFFARX1 I_6017 (I104997,I2683,I104929,I105023,);
DFFARX1 I_6018 (I1026570,I2683,I104929,I105040,);
and I_6019 (I105048,I105040,I1026564);
nor I_6020 (I105065,I105023,I105048);
DFFARX1 I_6021 (I105065,I2683,I104929,I104897,);
nand I_6022 (I105096,I105040,I1026564);
nand I_6023 (I105113,I104963,I105096);
not I_6024 (I104909,I105113);
DFFARX1 I_6025 (I1026552,I2683,I104929,I105153,);
DFFARX1 I_6026 (I105153,I2683,I104929,I104918,);
nand I_6027 (I105175,I1026567,I1026555);
and I_6028 (I105192,I105175,I1026579);
DFFARX1 I_6029 (I105192,I2683,I104929,I105218,);
DFFARX1 I_6030 (I105218,I2683,I104929,I105235,);
not I_6031 (I104921,I105235);
not I_6032 (I105257,I105218);
nand I_6033 (I104906,I105257,I105096);
nor I_6034 (I105288,I1026561,I1026555);
not I_6035 (I105305,I105288);
nor I_6036 (I105322,I105257,I105305);
nor I_6037 (I105339,I104963,I105322);
DFFARX1 I_6038 (I105339,I2683,I104929,I104915,);
nor I_6039 (I105370,I105023,I105305);
nor I_6040 (I104903,I105218,I105370);
nor I_6041 (I104912,I105153,I105288);
nor I_6042 (I104900,I105023,I105288);
not I_6043 (I105456,I2690);
DFFARX1 I_6044 (I785246,I2683,I105456,I105482,);
not I_6045 (I105490,I105482);
nand I_6046 (I105507,I785264,I785258);
and I_6047 (I105524,I105507,I785237);
DFFARX1 I_6048 (I105524,I2683,I105456,I105550,);
DFFARX1 I_6049 (I785255,I2683,I105456,I105567,);
and I_6050 (I105575,I105567,I785240);
nor I_6051 (I105592,I105550,I105575);
DFFARX1 I_6052 (I105592,I2683,I105456,I105424,);
nand I_6053 (I105623,I105567,I785240);
nand I_6054 (I105640,I105490,I105623);
not I_6055 (I105436,I105640);
DFFARX1 I_6056 (I785252,I2683,I105456,I105680,);
DFFARX1 I_6057 (I105680,I2683,I105456,I105445,);
nand I_6058 (I105702,I785261,I785249);
and I_6059 (I105719,I105702,I785243);
DFFARX1 I_6060 (I105719,I2683,I105456,I105745,);
DFFARX1 I_6061 (I105745,I2683,I105456,I105762,);
not I_6062 (I105448,I105762);
not I_6063 (I105784,I105745);
nand I_6064 (I105433,I105784,I105623);
nor I_6065 (I105815,I785237,I785249);
not I_6066 (I105832,I105815);
nor I_6067 (I105849,I105784,I105832);
nor I_6068 (I105866,I105490,I105849);
DFFARX1 I_6069 (I105866,I2683,I105456,I105442,);
nor I_6070 (I105897,I105550,I105832);
nor I_6071 (I105430,I105745,I105897);
nor I_6072 (I105439,I105680,I105815);
nor I_6073 (I105427,I105550,I105815);
not I_6074 (I105983,I2690);
DFFARX1 I_6075 (I285974,I2683,I105983,I106009,);
not I_6076 (I106017,I106009);
nand I_6077 (I106034,I285956,I285971);
and I_6078 (I106051,I106034,I285947);
DFFARX1 I_6079 (I106051,I2683,I105983,I106077,);
DFFARX1 I_6080 (I285950,I2683,I105983,I106094,);
and I_6081 (I106102,I106094,I285965);
nor I_6082 (I106119,I106077,I106102);
DFFARX1 I_6083 (I106119,I2683,I105983,I105951,);
nand I_6084 (I106150,I106094,I285965);
nand I_6085 (I106167,I106017,I106150);
not I_6086 (I105963,I106167);
DFFARX1 I_6087 (I285968,I2683,I105983,I106207,);
DFFARX1 I_6088 (I106207,I2683,I105983,I105972,);
nand I_6089 (I106229,I285947,I285959);
and I_6090 (I106246,I106229,I285953);
DFFARX1 I_6091 (I106246,I2683,I105983,I106272,);
DFFARX1 I_6092 (I106272,I2683,I105983,I106289,);
not I_6093 (I105975,I106289);
not I_6094 (I106311,I106272);
nand I_6095 (I105960,I106311,I106150);
nor I_6096 (I106342,I285962,I285959);
not I_6097 (I106359,I106342);
nor I_6098 (I106376,I106311,I106359);
nor I_6099 (I106393,I106017,I106376);
DFFARX1 I_6100 (I106393,I2683,I105983,I105969,);
nor I_6101 (I106424,I106077,I106359);
nor I_6102 (I105957,I106272,I106424);
nor I_6103 (I105966,I106207,I106342);
nor I_6104 (I105954,I106077,I106342);
not I_6105 (I106510,I2690);
DFFARX1 I_6106 (I149177,I2683,I106510,I106536,);
not I_6107 (I106544,I106536);
nand I_6108 (I106561,I149171,I149165);
and I_6109 (I106578,I106561,I149186);
DFFARX1 I_6110 (I106578,I2683,I106510,I106604,);
DFFARX1 I_6111 (I149183,I2683,I106510,I106621,);
and I_6112 (I106629,I106621,I149180);
nor I_6113 (I106646,I106604,I106629);
DFFARX1 I_6114 (I106646,I2683,I106510,I106478,);
nand I_6115 (I106677,I106621,I149180);
nand I_6116 (I106694,I106544,I106677);
not I_6117 (I106490,I106694);
DFFARX1 I_6118 (I149165,I2683,I106510,I106734,);
DFFARX1 I_6119 (I106734,I2683,I106510,I106499,);
nand I_6120 (I106756,I149168,I149168);
and I_6121 (I106773,I106756,I149189);
DFFARX1 I_6122 (I106773,I2683,I106510,I106799,);
DFFARX1 I_6123 (I106799,I2683,I106510,I106816,);
not I_6124 (I106502,I106816);
not I_6125 (I106838,I106799);
nand I_6126 (I106487,I106838,I106677);
nor I_6127 (I106869,I149174,I149168);
not I_6128 (I106886,I106869);
nor I_6129 (I106903,I106838,I106886);
nor I_6130 (I106920,I106544,I106903);
DFFARX1 I_6131 (I106920,I2683,I106510,I106496,);
nor I_6132 (I106951,I106604,I106886);
nor I_6133 (I106484,I106799,I106951);
nor I_6134 (I106493,I106734,I106869);
nor I_6135 (I106481,I106604,I106869);
not I_6136 (I107037,I2690);
DFFARX1 I_6137 (I902764,I2683,I107037,I107063,);
not I_6138 (I107071,I107063);
nand I_6139 (I107088,I902779,I902758);
and I_6140 (I107105,I107088,I902761);
DFFARX1 I_6141 (I107105,I2683,I107037,I107131,);
DFFARX1 I_6142 (I902782,I2683,I107037,I107148,);
and I_6143 (I107156,I107148,I902761);
nor I_6144 (I107173,I107131,I107156);
DFFARX1 I_6145 (I107173,I2683,I107037,I107005,);
nand I_6146 (I107204,I107148,I902761);
nand I_6147 (I107221,I107071,I107204);
not I_6148 (I107017,I107221);
DFFARX1 I_6149 (I902758,I2683,I107037,I107261,);
DFFARX1 I_6150 (I107261,I2683,I107037,I107026,);
nand I_6151 (I107283,I902770,I902767);
and I_6152 (I107300,I107283,I902773);
DFFARX1 I_6153 (I107300,I2683,I107037,I107326,);
DFFARX1 I_6154 (I107326,I2683,I107037,I107343,);
not I_6155 (I107029,I107343);
not I_6156 (I107365,I107326);
nand I_6157 (I107014,I107365,I107204);
nor I_6158 (I107396,I902776,I902767);
not I_6159 (I107413,I107396);
nor I_6160 (I107430,I107365,I107413);
nor I_6161 (I107447,I107071,I107430);
DFFARX1 I_6162 (I107447,I2683,I107037,I107023,);
nor I_6163 (I107478,I107131,I107413);
nor I_6164 (I107011,I107326,I107478);
nor I_6165 (I107020,I107261,I107396);
nor I_6166 (I107008,I107131,I107396);
not I_6167 (I107564,I2690);
DFFARX1 I_6168 (I408010,I2683,I107564,I107590,);
not I_6169 (I107598,I107590);
nand I_6170 (I107615,I408031,I408025);
and I_6171 (I107632,I107615,I408007);
DFFARX1 I_6172 (I107632,I2683,I107564,I107658,);
DFFARX1 I_6173 (I408010,I2683,I107564,I107675,);
and I_6174 (I107683,I107675,I408019);
nor I_6175 (I107700,I107658,I107683);
DFFARX1 I_6176 (I107700,I2683,I107564,I107532,);
nand I_6177 (I107731,I107675,I408019);
nand I_6178 (I107748,I107598,I107731);
not I_6179 (I107544,I107748);
DFFARX1 I_6180 (I408016,I2683,I107564,I107788,);
DFFARX1 I_6181 (I107788,I2683,I107564,I107553,);
nand I_6182 (I107810,I408022,I408013);
and I_6183 (I107827,I107810,I408007);
DFFARX1 I_6184 (I107827,I2683,I107564,I107853,);
DFFARX1 I_6185 (I107853,I2683,I107564,I107870,);
not I_6186 (I107556,I107870);
not I_6187 (I107892,I107853);
nand I_6188 (I107541,I107892,I107731);
nor I_6189 (I107923,I408028,I408013);
not I_6190 (I107940,I107923);
nor I_6191 (I107957,I107892,I107940);
nor I_6192 (I107974,I107598,I107957);
DFFARX1 I_6193 (I107974,I2683,I107564,I107550,);
nor I_6194 (I108005,I107658,I107940);
nor I_6195 (I107538,I107853,I108005);
nor I_6196 (I107547,I107788,I107923);
nor I_6197 (I107535,I107658,I107923);
not I_6198 (I108091,I2690);
DFFARX1 I_6199 (I584428,I2683,I108091,I108117,);
not I_6200 (I108125,I108117);
nand I_6201 (I108142,I584419,I584437);
and I_6202 (I108159,I108142,I584416);
DFFARX1 I_6203 (I108159,I2683,I108091,I108185,);
DFFARX1 I_6204 (I584419,I2683,I108091,I108202,);
and I_6205 (I108210,I108202,I584422);
nor I_6206 (I108227,I108185,I108210);
DFFARX1 I_6207 (I108227,I2683,I108091,I108059,);
nand I_6208 (I108258,I108202,I584422);
nand I_6209 (I108275,I108125,I108258);
not I_6210 (I108071,I108275);
DFFARX1 I_6211 (I584416,I2683,I108091,I108315,);
DFFARX1 I_6212 (I108315,I2683,I108091,I108080,);
nand I_6213 (I108337,I584434,I584425);
and I_6214 (I108354,I108337,I584440);
DFFARX1 I_6215 (I108354,I2683,I108091,I108380,);
DFFARX1 I_6216 (I108380,I2683,I108091,I108397,);
not I_6217 (I108083,I108397);
not I_6218 (I108419,I108380);
nand I_6219 (I108068,I108419,I108258);
nor I_6220 (I108450,I584431,I584425);
not I_6221 (I108467,I108450);
nor I_6222 (I108484,I108419,I108467);
nor I_6223 (I108501,I108125,I108484);
DFFARX1 I_6224 (I108501,I2683,I108091,I108077,);
nor I_6225 (I108532,I108185,I108467);
nor I_6226 (I108065,I108380,I108532);
nor I_6227 (I108074,I108315,I108450);
nor I_6228 (I108062,I108185,I108450);
not I_6229 (I108618,I2690);
DFFARX1 I_6230 (I820906,I2683,I108618,I108644,);
not I_6231 (I108652,I108644);
nand I_6232 (I108669,I820903,I820909);
and I_6233 (I108686,I108669,I820906);
DFFARX1 I_6234 (I108686,I2683,I108618,I108712,);
DFFARX1 I_6235 (I820909,I2683,I108618,I108729,);
and I_6236 (I108737,I108729,I820903);
nor I_6237 (I108754,I108712,I108737);
DFFARX1 I_6238 (I108754,I2683,I108618,I108586,);
nand I_6239 (I108785,I108729,I820903);
nand I_6240 (I108802,I108652,I108785);
not I_6241 (I108598,I108802);
DFFARX1 I_6242 (I820912,I2683,I108618,I108842,);
DFFARX1 I_6243 (I108842,I2683,I108618,I108607,);
nand I_6244 (I108864,I820915,I820924);
and I_6245 (I108881,I108864,I820918);
DFFARX1 I_6246 (I108881,I2683,I108618,I108907,);
DFFARX1 I_6247 (I108907,I2683,I108618,I108924,);
not I_6248 (I108610,I108924);
not I_6249 (I108946,I108907);
nand I_6250 (I108595,I108946,I108785);
nor I_6251 (I108977,I820921,I820924);
not I_6252 (I108994,I108977);
nor I_6253 (I109011,I108946,I108994);
nor I_6254 (I109028,I108652,I109011);
DFFARX1 I_6255 (I109028,I2683,I108618,I108604,);
nor I_6256 (I109059,I108712,I108994);
nor I_6257 (I108592,I108907,I109059);
nor I_6258 (I108601,I108842,I108977);
nor I_6259 (I108589,I108712,I108977);
not I_6260 (I109145,I2690);
DFFARX1 I_6261 (I515068,I2683,I109145,I109171,);
not I_6262 (I109179,I109171);
nand I_6263 (I109196,I515059,I515077);
and I_6264 (I109213,I109196,I515056);
DFFARX1 I_6265 (I109213,I2683,I109145,I109239,);
DFFARX1 I_6266 (I515059,I2683,I109145,I109256,);
and I_6267 (I109264,I109256,I515062);
nor I_6268 (I109281,I109239,I109264);
DFFARX1 I_6269 (I109281,I2683,I109145,I109113,);
nand I_6270 (I109312,I109256,I515062);
nand I_6271 (I109329,I109179,I109312);
not I_6272 (I109125,I109329);
DFFARX1 I_6273 (I515056,I2683,I109145,I109369,);
DFFARX1 I_6274 (I109369,I2683,I109145,I109134,);
nand I_6275 (I109391,I515074,I515065);
and I_6276 (I109408,I109391,I515080);
DFFARX1 I_6277 (I109408,I2683,I109145,I109434,);
DFFARX1 I_6278 (I109434,I2683,I109145,I109451,);
not I_6279 (I109137,I109451);
not I_6280 (I109473,I109434);
nand I_6281 (I109122,I109473,I109312);
nor I_6282 (I109504,I515071,I515065);
not I_6283 (I109521,I109504);
nor I_6284 (I109538,I109473,I109521);
nor I_6285 (I109555,I109179,I109538);
DFFARX1 I_6286 (I109555,I2683,I109145,I109131,);
nor I_6287 (I109586,I109239,I109521);
nor I_6288 (I109119,I109434,I109586);
nor I_6289 (I109128,I109369,I109504);
nor I_6290 (I109116,I109239,I109504);
not I_6291 (I109672,I2690);
DFFARX1 I_6292 (I411580,I2683,I109672,I109698,);
not I_6293 (I109706,I109698);
nand I_6294 (I109723,I411601,I411595);
and I_6295 (I109740,I109723,I411577);
DFFARX1 I_6296 (I109740,I2683,I109672,I109766,);
DFFARX1 I_6297 (I411580,I2683,I109672,I109783,);
and I_6298 (I109791,I109783,I411589);
nor I_6299 (I109808,I109766,I109791);
DFFARX1 I_6300 (I109808,I2683,I109672,I109640,);
nand I_6301 (I109839,I109783,I411589);
nand I_6302 (I109856,I109706,I109839);
not I_6303 (I109652,I109856);
DFFARX1 I_6304 (I411586,I2683,I109672,I109896,);
DFFARX1 I_6305 (I109896,I2683,I109672,I109661,);
nand I_6306 (I109918,I411592,I411583);
and I_6307 (I109935,I109918,I411577);
DFFARX1 I_6308 (I109935,I2683,I109672,I109961,);
DFFARX1 I_6309 (I109961,I2683,I109672,I109978,);
not I_6310 (I109664,I109978);
not I_6311 (I110000,I109961);
nand I_6312 (I109649,I110000,I109839);
nor I_6313 (I110031,I411598,I411583);
not I_6314 (I110048,I110031);
nor I_6315 (I110065,I110000,I110048);
nor I_6316 (I110082,I109706,I110065);
DFFARX1 I_6317 (I110082,I2683,I109672,I109658,);
nor I_6318 (I110113,I109766,I110048);
nor I_6319 (I109646,I109961,I110113);
nor I_6320 (I109655,I109896,I110031);
nor I_6321 (I109643,I109766,I110031);
not I_6322 (I110199,I2690);
DFFARX1 I_6323 (I613906,I2683,I110199,I110225,);
not I_6324 (I110233,I110225);
nand I_6325 (I110250,I613897,I613915);
and I_6326 (I110267,I110250,I613894);
DFFARX1 I_6327 (I110267,I2683,I110199,I110293,);
DFFARX1 I_6328 (I613897,I2683,I110199,I110310,);
and I_6329 (I110318,I110310,I613900);
nor I_6330 (I110335,I110293,I110318);
DFFARX1 I_6331 (I110335,I2683,I110199,I110167,);
nand I_6332 (I110366,I110310,I613900);
nand I_6333 (I110383,I110233,I110366);
not I_6334 (I110179,I110383);
DFFARX1 I_6335 (I613894,I2683,I110199,I110423,);
DFFARX1 I_6336 (I110423,I2683,I110199,I110188,);
nand I_6337 (I110445,I613912,I613903);
and I_6338 (I110462,I110445,I613918);
DFFARX1 I_6339 (I110462,I2683,I110199,I110488,);
DFFARX1 I_6340 (I110488,I2683,I110199,I110505,);
not I_6341 (I110191,I110505);
not I_6342 (I110527,I110488);
nand I_6343 (I110176,I110527,I110366);
nor I_6344 (I110558,I613909,I613903);
not I_6345 (I110575,I110558);
nor I_6346 (I110592,I110527,I110575);
nor I_6347 (I110609,I110233,I110592);
DFFARX1 I_6348 (I110609,I2683,I110199,I110185,);
nor I_6349 (I110640,I110293,I110575);
nor I_6350 (I110173,I110488,I110640);
nor I_6351 (I110182,I110423,I110558);
nor I_6352 (I110170,I110293,I110558);
not I_6353 (I110726,I2690);
DFFARX1 I_6354 (I897562,I2683,I110726,I110752,);
not I_6355 (I110760,I110752);
nand I_6356 (I110777,I897577,I897556);
and I_6357 (I110794,I110777,I897559);
DFFARX1 I_6358 (I110794,I2683,I110726,I110820,);
DFFARX1 I_6359 (I897580,I2683,I110726,I110837,);
and I_6360 (I110845,I110837,I897559);
nor I_6361 (I110862,I110820,I110845);
DFFARX1 I_6362 (I110862,I2683,I110726,I110694,);
nand I_6363 (I110893,I110837,I897559);
nand I_6364 (I110910,I110760,I110893);
not I_6365 (I110706,I110910);
DFFARX1 I_6366 (I897556,I2683,I110726,I110950,);
DFFARX1 I_6367 (I110950,I2683,I110726,I110715,);
nand I_6368 (I110972,I897568,I897565);
and I_6369 (I110989,I110972,I897571);
DFFARX1 I_6370 (I110989,I2683,I110726,I111015,);
DFFARX1 I_6371 (I111015,I2683,I110726,I111032,);
not I_6372 (I110718,I111032);
not I_6373 (I111054,I111015);
nand I_6374 (I110703,I111054,I110893);
nor I_6375 (I111085,I897574,I897565);
not I_6376 (I111102,I111085);
nor I_6377 (I111119,I111054,I111102);
nor I_6378 (I111136,I110760,I111119);
DFFARX1 I_6379 (I111136,I2683,I110726,I110712,);
nor I_6380 (I111167,I110820,I111102);
nor I_6381 (I110700,I111015,I111167);
nor I_6382 (I110709,I110950,I111085);
nor I_6383 (I110697,I110820,I111085);
not I_6384 (I111253,I2690);
DFFARX1 I_6385 (I931086,I2683,I111253,I111279,);
not I_6386 (I111287,I111279);
nand I_6387 (I111304,I931101,I931080);
and I_6388 (I111321,I111304,I931083);
DFFARX1 I_6389 (I111321,I2683,I111253,I111347,);
DFFARX1 I_6390 (I931104,I2683,I111253,I111364,);
and I_6391 (I111372,I111364,I931083);
nor I_6392 (I111389,I111347,I111372);
DFFARX1 I_6393 (I111389,I2683,I111253,I111221,);
nand I_6394 (I111420,I111364,I931083);
nand I_6395 (I111437,I111287,I111420);
not I_6396 (I111233,I111437);
DFFARX1 I_6397 (I931080,I2683,I111253,I111477,);
DFFARX1 I_6398 (I111477,I2683,I111253,I111242,);
nand I_6399 (I111499,I931092,I931089);
and I_6400 (I111516,I111499,I931095);
DFFARX1 I_6401 (I111516,I2683,I111253,I111542,);
DFFARX1 I_6402 (I111542,I2683,I111253,I111559,);
not I_6403 (I111245,I111559);
not I_6404 (I111581,I111542);
nand I_6405 (I111230,I111581,I111420);
nor I_6406 (I111612,I931098,I931089);
not I_6407 (I111629,I111612);
nor I_6408 (I111646,I111581,I111629);
nor I_6409 (I111663,I111287,I111646);
DFFARX1 I_6410 (I111663,I2683,I111253,I111239,);
nor I_6411 (I111694,I111347,I111629);
nor I_6412 (I111227,I111542,I111694);
nor I_6413 (I111236,I111477,I111612);
nor I_6414 (I111224,I111347,I111612);
not I_6415 (I111780,I2690);
DFFARX1 I_6416 (I263313,I2683,I111780,I111806,);
not I_6417 (I111814,I111806);
nand I_6418 (I111831,I263295,I263310);
and I_6419 (I111848,I111831,I263286);
DFFARX1 I_6420 (I111848,I2683,I111780,I111874,);
DFFARX1 I_6421 (I263289,I2683,I111780,I111891,);
and I_6422 (I111899,I111891,I263304);
nor I_6423 (I111916,I111874,I111899);
DFFARX1 I_6424 (I111916,I2683,I111780,I111748,);
nand I_6425 (I111947,I111891,I263304);
nand I_6426 (I111964,I111814,I111947);
not I_6427 (I111760,I111964);
DFFARX1 I_6428 (I263307,I2683,I111780,I112004,);
DFFARX1 I_6429 (I112004,I2683,I111780,I111769,);
nand I_6430 (I112026,I263286,I263298);
and I_6431 (I112043,I112026,I263292);
DFFARX1 I_6432 (I112043,I2683,I111780,I112069,);
DFFARX1 I_6433 (I112069,I2683,I111780,I112086,);
not I_6434 (I111772,I112086);
not I_6435 (I112108,I112069);
nand I_6436 (I111757,I112108,I111947);
nor I_6437 (I112139,I263301,I263298);
not I_6438 (I112156,I112139);
nor I_6439 (I112173,I112108,I112156);
nor I_6440 (I112190,I111814,I112173);
DFFARX1 I_6441 (I112190,I2683,I111780,I111766,);
nor I_6442 (I112221,I111874,I112156);
nor I_6443 (I111754,I112069,I112221);
nor I_6444 (I111763,I112004,I112139);
nor I_6445 (I111751,I111874,I112139);
not I_6446 (I112310,I2690);
DFFARX1 I_6447 (I286483,I2683,I112310,I112336,);
not I_6448 (I112344,I112336);
DFFARX1 I_6449 (I286480,I2683,I112310,I112370,);
not I_6450 (I112378,I286477);
or I_6451 (I112395,I286489,I286477);
nor I_6452 (I112412,I112370,I286489);
nand I_6453 (I112287,I112378,I112412);
nor I_6454 (I112443,I286498,I286489);
nand I_6455 (I112281,I112443,I112378);
not I_6456 (I112474,I286495);
nand I_6457 (I112491,I112378,I112474);
nor I_6458 (I112508,I286474,I286474);
not I_6459 (I112525,I112508);
nor I_6460 (I112542,I112525,I112491);
nor I_6461 (I112559,I112443,I112542);
DFFARX1 I_6462 (I112559,I2683,I112310,I112296,);
nor I_6463 (I112293,I112508,I112395);
DFFARX1 I_6464 (I112508,I2683,I112310,I112299,);
nor I_6465 (I112618,I112474,I286474);
nor I_6466 (I112635,I112618,I286477);
nor I_6467 (I112652,I286486,I286501);
DFFARX1 I_6468 (I112652,I2683,I112310,I112678,);
nor I_6469 (I112278,I112678,I112635);
DFFARX1 I_6470 (I112678,I2683,I112310,I112709,);
nand I_6471 (I112717,I112709,I286492);
nor I_6472 (I112302,I112344,I112717);
not I_6473 (I112748,I112678);
nand I_6474 (I112765,I112748,I286492);
nor I_6475 (I112782,I112344,I112765);
nor I_6476 (I112284,I112370,I112782);
nor I_6477 (I112813,I286486,I286498);
nor I_6478 (I112830,I112370,I112813);
DFFARX1 I_6479 (I112830,I2683,I112310,I112275,);
and I_6480 (I112290,I112443,I286486);
not I_6481 (I112905,I2690);
DFFARX1 I_6482 (I434151,I2683,I112905,I112931,);
not I_6483 (I112939,I112931);
DFFARX1 I_6484 (I434136,I2683,I112905,I112965,);
not I_6485 (I112973,I434160);
or I_6486 (I112990,I434139,I434160);
nor I_6487 (I113007,I112965,I434139);
nand I_6488 (I112882,I112973,I113007);
nor I_6489 (I113038,I434142,I434139);
nand I_6490 (I112876,I113038,I112973);
not I_6491 (I113069,I434145);
nand I_6492 (I113086,I112973,I113069);
nor I_6493 (I113103,I434148,I434154);
not I_6494 (I113120,I113103);
nor I_6495 (I113137,I113120,I113086);
nor I_6496 (I113154,I113038,I113137);
DFFARX1 I_6497 (I113154,I2683,I112905,I112891,);
nor I_6498 (I112888,I113103,I112990);
DFFARX1 I_6499 (I113103,I2683,I112905,I112894,);
nor I_6500 (I113213,I113069,I434148);
nor I_6501 (I113230,I113213,I434160);
nor I_6502 (I113247,I434157,I434139);
DFFARX1 I_6503 (I113247,I2683,I112905,I113273,);
nor I_6504 (I112873,I113273,I113230);
DFFARX1 I_6505 (I113273,I2683,I112905,I113304,);
nand I_6506 (I113312,I113304,I434136);
nor I_6507 (I112897,I112939,I113312);
not I_6508 (I113343,I113273);
nand I_6509 (I113360,I113343,I434136);
nor I_6510 (I113377,I112939,I113360);
nor I_6511 (I112879,I112965,I113377);
nor I_6512 (I113408,I434157,I434142);
nor I_6513 (I113425,I112965,I113408);
DFFARX1 I_6514 (I113425,I2683,I112905,I112870,);
and I_6515 (I112885,I113038,I434157);
not I_6516 (I113500,I2690);
DFFARX1 I_6517 (I945533,I2683,I113500,I113526,);
not I_6518 (I113534,I113526);
DFFARX1 I_6519 (I945530,I2683,I113500,I113560,);
not I_6520 (I113568,I945539);
or I_6521 (I113585,I945530,I945539);
nor I_6522 (I113602,I113560,I945530);
nand I_6523 (I113477,I113568,I113602);
nor I_6524 (I113633,I945542,I945530);
nand I_6525 (I113471,I113633,I113568);
not I_6526 (I113664,I945536);
nand I_6527 (I113681,I113568,I113664);
nor I_6528 (I113698,I945533,I945551);
not I_6529 (I113715,I113698);
nor I_6530 (I113732,I113715,I113681);
nor I_6531 (I113749,I113633,I113732);
DFFARX1 I_6532 (I113749,I2683,I113500,I113486,);
nor I_6533 (I113483,I113698,I113585);
DFFARX1 I_6534 (I113698,I2683,I113500,I113489,);
nor I_6535 (I113808,I113664,I945533);
nor I_6536 (I113825,I113808,I945539);
nor I_6537 (I113842,I945554,I945548);
DFFARX1 I_6538 (I113842,I2683,I113500,I113868,);
nor I_6539 (I113468,I113868,I113825);
DFFARX1 I_6540 (I113868,I2683,I113500,I113899,);
nand I_6541 (I113907,I113899,I945545);
nor I_6542 (I113492,I113534,I113907);
not I_6543 (I113938,I113868);
nand I_6544 (I113955,I113938,I945545);
nor I_6545 (I113972,I113534,I113955);
nor I_6546 (I113474,I113560,I113972);
nor I_6547 (I114003,I945554,I945542);
nor I_6548 (I114020,I113560,I114003);
DFFARX1 I_6549 (I114020,I2683,I113500,I113465,);
and I_6550 (I113480,I113633,I945554);
not I_6551 (I114095,I2690);
DFFARX1 I_6552 (I491373,I2683,I114095,I114121,);
not I_6553 (I114129,I114121);
DFFARX1 I_6554 (I491358,I2683,I114095,I114155,);
not I_6555 (I114163,I491382);
or I_6556 (I114180,I491361,I491382);
nor I_6557 (I114197,I114155,I491361);
nand I_6558 (I114072,I114163,I114197);
nor I_6559 (I114228,I491364,I491361);
nand I_6560 (I114066,I114228,I114163);
not I_6561 (I114259,I491367);
nand I_6562 (I114276,I114163,I114259);
nor I_6563 (I114293,I491370,I491376);
not I_6564 (I114310,I114293);
nor I_6565 (I114327,I114310,I114276);
nor I_6566 (I114344,I114228,I114327);
DFFARX1 I_6567 (I114344,I2683,I114095,I114081,);
nor I_6568 (I114078,I114293,I114180);
DFFARX1 I_6569 (I114293,I2683,I114095,I114084,);
nor I_6570 (I114403,I114259,I491370);
nor I_6571 (I114420,I114403,I491382);
nor I_6572 (I114437,I491379,I491361);
DFFARX1 I_6573 (I114437,I2683,I114095,I114463,);
nor I_6574 (I114063,I114463,I114420);
DFFARX1 I_6575 (I114463,I2683,I114095,I114494,);
nand I_6576 (I114502,I114494,I491358);
nor I_6577 (I114087,I114129,I114502);
not I_6578 (I114533,I114463);
nand I_6579 (I114550,I114533,I491358);
nor I_6580 (I114567,I114129,I114550);
nor I_6581 (I114069,I114155,I114567);
nor I_6582 (I114598,I491379,I491364);
nor I_6583 (I114615,I114155,I114598);
DFFARX1 I_6584 (I114615,I2683,I114095,I114060,);
and I_6585 (I114075,I114228,I491379);
not I_6586 (I114690,I2690);
DFFARX1 I_6587 (I875595,I2683,I114690,I114716,);
not I_6588 (I114724,I114716);
DFFARX1 I_6589 (I875592,I2683,I114690,I114750,);
not I_6590 (I114758,I875601);
or I_6591 (I114775,I875592,I875601);
nor I_6592 (I114792,I114750,I875592);
nand I_6593 (I114667,I114758,I114792);
nor I_6594 (I114823,I875604,I875592);
nand I_6595 (I114661,I114823,I114758);
not I_6596 (I114854,I875598);
nand I_6597 (I114871,I114758,I114854);
nor I_6598 (I114888,I875595,I875613);
not I_6599 (I114905,I114888);
nor I_6600 (I114922,I114905,I114871);
nor I_6601 (I114939,I114823,I114922);
DFFARX1 I_6602 (I114939,I2683,I114690,I114676,);
nor I_6603 (I114673,I114888,I114775);
DFFARX1 I_6604 (I114888,I2683,I114690,I114679,);
nor I_6605 (I114998,I114854,I875595);
nor I_6606 (I115015,I114998,I875601);
nor I_6607 (I115032,I875616,I875610);
DFFARX1 I_6608 (I115032,I2683,I114690,I115058,);
nor I_6609 (I114658,I115058,I115015);
DFFARX1 I_6610 (I115058,I2683,I114690,I115089,);
nand I_6611 (I115097,I115089,I875607);
nor I_6612 (I114682,I114724,I115097);
not I_6613 (I115128,I115058);
nand I_6614 (I115145,I115128,I875607);
nor I_6615 (I115162,I114724,I115145);
nor I_6616 (I114664,I114750,I115162);
nor I_6617 (I115193,I875616,I875604);
nor I_6618 (I115210,I114750,I115193);
DFFARX1 I_6619 (I115210,I2683,I114690,I114655,);
and I_6620 (I114670,I114823,I875616);
not I_6621 (I115285,I2690);
DFFARX1 I_6622 (I259079,I2683,I115285,I115311,);
not I_6623 (I115319,I115311);
DFFARX1 I_6624 (I259076,I2683,I115285,I115345,);
not I_6625 (I115353,I259073);
or I_6626 (I115370,I259085,I259073);
nor I_6627 (I115387,I115345,I259085);
nand I_6628 (I115262,I115353,I115387);
nor I_6629 (I115418,I259094,I259085);
nand I_6630 (I115256,I115418,I115353);
not I_6631 (I115449,I259091);
nand I_6632 (I115466,I115353,I115449);
nor I_6633 (I115483,I259070,I259070);
not I_6634 (I115500,I115483);
nor I_6635 (I115517,I115500,I115466);
nor I_6636 (I115534,I115418,I115517);
DFFARX1 I_6637 (I115534,I2683,I115285,I115271,);
nor I_6638 (I115268,I115483,I115370);
DFFARX1 I_6639 (I115483,I2683,I115285,I115274,);
nor I_6640 (I115593,I115449,I259070);
nor I_6641 (I115610,I115593,I259073);
nor I_6642 (I115627,I259082,I259097);
DFFARX1 I_6643 (I115627,I2683,I115285,I115653,);
nor I_6644 (I115253,I115653,I115610);
DFFARX1 I_6645 (I115653,I2683,I115285,I115684,);
nand I_6646 (I115692,I115684,I259088);
nor I_6647 (I115277,I115319,I115692);
not I_6648 (I115723,I115653);
nand I_6649 (I115740,I115723,I259088);
nor I_6650 (I115757,I115319,I115740);
nor I_6651 (I115259,I115345,I115757);
nor I_6652 (I115788,I259082,I259094);
nor I_6653 (I115805,I115345,I115788);
DFFARX1 I_6654 (I115805,I2683,I115285,I115250,);
and I_6655 (I115265,I115418,I259082);
not I_6656 (I115880,I2690);
DFFARX1 I_6657 (I678126,I2683,I115880,I115906,);
not I_6658 (I115914,I115906);
DFFARX1 I_6659 (I678126,I2683,I115880,I115940,);
not I_6660 (I115948,I678123);
or I_6661 (I115965,I678135,I678123);
nor I_6662 (I115982,I115940,I678135);
nand I_6663 (I115857,I115948,I115982);
nor I_6664 (I116013,I678129,I678135);
nand I_6665 (I115851,I116013,I115948);
not I_6666 (I116044,I678141);
nand I_6667 (I116061,I115948,I116044);
nor I_6668 (I116078,I678132,I678120);
not I_6669 (I116095,I116078);
nor I_6670 (I116112,I116095,I116061);
nor I_6671 (I116129,I116013,I116112);
DFFARX1 I_6672 (I116129,I2683,I115880,I115866,);
nor I_6673 (I115863,I116078,I115965);
DFFARX1 I_6674 (I116078,I2683,I115880,I115869,);
nor I_6675 (I116188,I116044,I678132);
nor I_6676 (I116205,I116188,I678123);
nor I_6677 (I116222,I678123,I678120);
DFFARX1 I_6678 (I116222,I2683,I115880,I116248,);
nor I_6679 (I115848,I116248,I116205);
DFFARX1 I_6680 (I116248,I2683,I115880,I116279,);
nand I_6681 (I116287,I116279,I678138);
nor I_6682 (I115872,I115914,I116287);
not I_6683 (I116318,I116248);
nand I_6684 (I116335,I116318,I678138);
nor I_6685 (I116352,I115914,I116335);
nor I_6686 (I115854,I115940,I116352);
nor I_6687 (I116383,I678123,I678129);
nor I_6688 (I116400,I115940,I116383);
DFFARX1 I_6689 (I116400,I2683,I115880,I115845,);
and I_6690 (I115860,I116013,I678123);
not I_6691 (I116475,I2690);
DFFARX1 I_6692 (I973889,I2683,I116475,I116501,);
not I_6693 (I116509,I116501);
DFFARX1 I_6694 (I973901,I2683,I116475,I116535,);
not I_6695 (I116543,I973907);
or I_6696 (I116560,I973886,I973907);
nor I_6697 (I116577,I116535,I973886);
nand I_6698 (I116452,I116543,I116577);
nor I_6699 (I116608,I973904,I973886);
nand I_6700 (I116446,I116608,I116543);
not I_6701 (I116639,I973889);
nand I_6702 (I116656,I116543,I116639);
nor I_6703 (I116673,I973892,I973886);
not I_6704 (I116690,I116673);
nor I_6705 (I116707,I116690,I116656);
nor I_6706 (I116724,I116608,I116707);
DFFARX1 I_6707 (I116724,I2683,I116475,I116461,);
nor I_6708 (I116458,I116673,I116560);
DFFARX1 I_6709 (I116673,I2683,I116475,I116464,);
nor I_6710 (I116783,I116639,I973892);
nor I_6711 (I116800,I116783,I973907);
nor I_6712 (I116817,I973910,I973898);
DFFARX1 I_6713 (I116817,I2683,I116475,I116843,);
nor I_6714 (I116443,I116843,I116800);
DFFARX1 I_6715 (I116843,I2683,I116475,I116874,);
nand I_6716 (I116882,I116874,I973895);
nor I_6717 (I116467,I116509,I116882);
not I_6718 (I116913,I116843);
nand I_6719 (I116930,I116913,I973895);
nor I_6720 (I116947,I116509,I116930);
nor I_6721 (I116449,I116535,I116947);
nor I_6722 (I116978,I973910,I973904);
nor I_6723 (I116995,I116535,I116978);
DFFARX1 I_6724 (I116995,I2683,I116475,I116440,);
and I_6725 (I116455,I116608,I973910);
not I_6726 (I117070,I2690);
DFFARX1 I_6727 (I298077,I2683,I117070,I117096,);
not I_6728 (I117104,I117096);
DFFARX1 I_6729 (I298074,I2683,I117070,I117130,);
not I_6730 (I117138,I298071);
or I_6731 (I117155,I298083,I298071);
nor I_6732 (I117172,I117130,I298083);
nand I_6733 (I117047,I117138,I117172);
nor I_6734 (I117203,I298092,I298083);
nand I_6735 (I117041,I117203,I117138);
not I_6736 (I117234,I298089);
nand I_6737 (I117251,I117138,I117234);
nor I_6738 (I117268,I298068,I298068);
not I_6739 (I117285,I117268);
nor I_6740 (I117302,I117285,I117251);
nor I_6741 (I117319,I117203,I117302);
DFFARX1 I_6742 (I117319,I2683,I117070,I117056,);
nor I_6743 (I117053,I117268,I117155);
DFFARX1 I_6744 (I117268,I2683,I117070,I117059,);
nor I_6745 (I117378,I117234,I298068);
nor I_6746 (I117395,I117378,I298071);
nor I_6747 (I117412,I298080,I298095);
DFFARX1 I_6748 (I117412,I2683,I117070,I117438,);
nor I_6749 (I117038,I117438,I117395);
DFFARX1 I_6750 (I117438,I2683,I117070,I117469,);
nand I_6751 (I117477,I117469,I298086);
nor I_6752 (I117062,I117104,I117477);
not I_6753 (I117508,I117438);
nand I_6754 (I117525,I117508,I298086);
nor I_6755 (I117542,I117104,I117525);
nor I_6756 (I117044,I117130,I117542);
nor I_6757 (I117573,I298080,I298092);
nor I_6758 (I117590,I117130,I117573);
DFFARX1 I_6759 (I117590,I2683,I117070,I117035,);
and I_6760 (I117050,I117203,I298080);
not I_6761 (I117665,I2690);
DFFARX1 I_6762 (I976065,I2683,I117665,I117691,);
not I_6763 (I117699,I117691);
DFFARX1 I_6764 (I976077,I2683,I117665,I117725,);
not I_6765 (I117733,I976083);
or I_6766 (I117750,I976062,I976083);
nor I_6767 (I117767,I117725,I976062);
nand I_6768 (I117642,I117733,I117767);
nor I_6769 (I117798,I976080,I976062);
nand I_6770 (I117636,I117798,I117733);
not I_6771 (I117829,I976065);
nand I_6772 (I117846,I117733,I117829);
nor I_6773 (I117863,I976068,I976062);
not I_6774 (I117880,I117863);
nor I_6775 (I117897,I117880,I117846);
nor I_6776 (I117914,I117798,I117897);
DFFARX1 I_6777 (I117914,I2683,I117665,I117651,);
nor I_6778 (I117648,I117863,I117750);
DFFARX1 I_6779 (I117863,I2683,I117665,I117654,);
nor I_6780 (I117973,I117829,I976068);
nor I_6781 (I117990,I117973,I976083);
nor I_6782 (I118007,I976086,I976074);
DFFARX1 I_6783 (I118007,I2683,I117665,I118033,);
nor I_6784 (I117633,I118033,I117990);
DFFARX1 I_6785 (I118033,I2683,I117665,I118064,);
nand I_6786 (I118072,I118064,I976071);
nor I_6787 (I117657,I117699,I118072);
not I_6788 (I118103,I118033);
nand I_6789 (I118120,I118103,I976071);
nor I_6790 (I118137,I117699,I118120);
nor I_6791 (I117639,I117725,I118137);
nor I_6792 (I118168,I976086,I976080);
nor I_6793 (I118185,I117725,I118168);
DFFARX1 I_6794 (I118185,I2683,I117665,I117630,);
and I_6795 (I117645,I117798,I976086);
not I_6796 (I118260,I2690);
DFFARX1 I_6797 (I662843,I2683,I118260,I118286,);
not I_6798 (I118294,I118286);
DFFARX1 I_6799 (I662843,I2683,I118260,I118320,);
not I_6800 (I118328,I662840);
or I_6801 (I118345,I662852,I662840);
nor I_6802 (I118362,I118320,I662852);
nand I_6803 (I118237,I118328,I118362);
nor I_6804 (I118393,I662846,I662852);
nand I_6805 (I118231,I118393,I118328);
not I_6806 (I118424,I662858);
nand I_6807 (I118441,I118328,I118424);
nor I_6808 (I118458,I662849,I662837);
not I_6809 (I118475,I118458);
nor I_6810 (I118492,I118475,I118441);
nor I_6811 (I118509,I118393,I118492);
DFFARX1 I_6812 (I118509,I2683,I118260,I118246,);
nor I_6813 (I118243,I118458,I118345);
DFFARX1 I_6814 (I118458,I2683,I118260,I118249,);
nor I_6815 (I118568,I118424,I662849);
nor I_6816 (I118585,I118568,I662840);
nor I_6817 (I118602,I662840,I662837);
DFFARX1 I_6818 (I118602,I2683,I118260,I118628,);
nor I_6819 (I118228,I118628,I118585);
DFFARX1 I_6820 (I118628,I2683,I118260,I118659,);
nand I_6821 (I118667,I118659,I662855);
nor I_6822 (I118252,I118294,I118667);
not I_6823 (I118698,I118628);
nand I_6824 (I118715,I118698,I662855);
nor I_6825 (I118732,I118294,I118715);
nor I_6826 (I118234,I118320,I118732);
nor I_6827 (I118763,I662840,I662846);
nor I_6828 (I118780,I118320,I118763);
DFFARX1 I_6829 (I118780,I2683,I118260,I118225,);
and I_6830 (I118240,I118393,I662840);
not I_6831 (I118855,I2690);
DFFARX1 I_6832 (I212176,I2683,I118855,I118881,);
not I_6833 (I118889,I118881);
DFFARX1 I_6834 (I212173,I2683,I118855,I118915,);
not I_6835 (I118923,I212170);
or I_6836 (I118940,I212182,I212170);
nor I_6837 (I118957,I118915,I212182);
nand I_6838 (I118832,I118923,I118957);
nor I_6839 (I118988,I212191,I212182);
nand I_6840 (I118826,I118988,I118923);
not I_6841 (I119019,I212188);
nand I_6842 (I119036,I118923,I119019);
nor I_6843 (I119053,I212167,I212167);
not I_6844 (I119070,I119053);
nor I_6845 (I119087,I119070,I119036);
nor I_6846 (I119104,I118988,I119087);
DFFARX1 I_6847 (I119104,I2683,I118855,I118841,);
nor I_6848 (I118838,I119053,I118940);
DFFARX1 I_6849 (I119053,I2683,I118855,I118844,);
nor I_6850 (I119163,I119019,I212167);
nor I_6851 (I119180,I119163,I212170);
nor I_6852 (I119197,I212179,I212194);
DFFARX1 I_6853 (I119197,I2683,I118855,I119223,);
nor I_6854 (I118823,I119223,I119180);
DFFARX1 I_6855 (I119223,I2683,I118855,I119254,);
nand I_6856 (I119262,I119254,I212185);
nor I_6857 (I118847,I118889,I119262);
not I_6858 (I119293,I119223);
nand I_6859 (I119310,I119293,I212185);
nor I_6860 (I119327,I118889,I119310);
nor I_6861 (I118829,I118915,I119327);
nor I_6862 (I119358,I212179,I212191);
nor I_6863 (I119375,I118915,I119358);
DFFARX1 I_6864 (I119375,I2683,I118855,I118820,);
and I_6865 (I118835,I118988,I212179);
not I_6866 (I119450,I2690);
DFFARX1 I_6867 (I360618,I2683,I119450,I119476,);
not I_6868 (I119484,I119476);
DFFARX1 I_6869 (I360612,I2683,I119450,I119510,);
not I_6870 (I119518,I360609);
or I_6871 (I119535,I360600,I360609);
nor I_6872 (I119552,I119510,I360600);
nand I_6873 (I119427,I119518,I119552);
nor I_6874 (I119583,I360603,I360600);
nand I_6875 (I119421,I119583,I119518);
not I_6876 (I119614,I360606);
nand I_6877 (I119631,I119518,I119614);
nor I_6878 (I119648,I360594,I360621);
not I_6879 (I119665,I119648);
nor I_6880 (I119682,I119665,I119631);
nor I_6881 (I119699,I119583,I119682);
DFFARX1 I_6882 (I119699,I2683,I119450,I119436,);
nor I_6883 (I119433,I119648,I119535);
DFFARX1 I_6884 (I119648,I2683,I119450,I119439,);
nor I_6885 (I119758,I119614,I360594);
nor I_6886 (I119775,I119758,I360609);
nor I_6887 (I119792,I360597,I360594);
DFFARX1 I_6888 (I119792,I2683,I119450,I119818,);
nor I_6889 (I119418,I119818,I119775);
DFFARX1 I_6890 (I119818,I2683,I119450,I119849,);
nand I_6891 (I119857,I119849,I360615);
nor I_6892 (I119442,I119484,I119857);
not I_6893 (I119888,I119818);
nand I_6894 (I119905,I119888,I360615);
nor I_6895 (I119922,I119484,I119905);
nor I_6896 (I119424,I119510,I119922);
nor I_6897 (I119953,I360597,I360603);
nor I_6898 (I119970,I119510,I119953);
DFFARX1 I_6899 (I119970,I2683,I119450,I119415,);
and I_6900 (I119430,I119583,I360597);
not I_6901 (I120045,I2690);
DFFARX1 I_6902 (I701909,I2683,I120045,I120071,);
not I_6903 (I120079,I120071);
DFFARX1 I_6904 (I701930,I2683,I120045,I120105,);
not I_6905 (I120113,I701912);
or I_6906 (I120130,I701903,I701912);
nor I_6907 (I120147,I120105,I701903);
nand I_6908 (I120022,I120113,I120147);
nor I_6909 (I120178,I701915,I701903);
nand I_6910 (I120016,I120178,I120113);
not I_6911 (I120209,I701906);
nand I_6912 (I120226,I120113,I120209);
nor I_6913 (I120243,I701924,I701927);
not I_6914 (I120260,I120243);
nor I_6915 (I120277,I120260,I120226);
nor I_6916 (I120294,I120178,I120277);
DFFARX1 I_6917 (I120294,I2683,I120045,I120031,);
nor I_6918 (I120028,I120243,I120130);
DFFARX1 I_6919 (I120243,I2683,I120045,I120034,);
nor I_6920 (I120353,I120209,I701924);
nor I_6921 (I120370,I120353,I701912);
nor I_6922 (I120387,I701918,I701921);
DFFARX1 I_6923 (I120387,I2683,I120045,I120413,);
nor I_6924 (I120013,I120413,I120370);
DFFARX1 I_6925 (I120413,I2683,I120045,I120444,);
nand I_6926 (I120452,I120444,I701903);
nor I_6927 (I120037,I120079,I120452);
not I_6928 (I120483,I120413);
nand I_6929 (I120500,I120483,I701903);
nor I_6930 (I120517,I120079,I120500);
nor I_6931 (I120019,I120105,I120517);
nor I_6932 (I120548,I701918,I701915);
nor I_6933 (I120565,I120105,I120548);
DFFARX1 I_6934 (I120565,I2683,I120045,I120010,);
and I_6935 (I120025,I120178,I701918);
not I_6936 (I120640,I2690);
DFFARX1 I_6937 (I767801,I2683,I120640,I120666,);
not I_6938 (I120674,I120666);
DFFARX1 I_6939 (I767822,I2683,I120640,I120700,);
not I_6940 (I120708,I767804);
or I_6941 (I120725,I767795,I767804);
nor I_6942 (I120742,I120700,I767795);
nand I_6943 (I120617,I120708,I120742);
nor I_6944 (I120773,I767807,I767795);
nand I_6945 (I120611,I120773,I120708);
not I_6946 (I120804,I767798);
nand I_6947 (I120821,I120708,I120804);
nor I_6948 (I120838,I767816,I767819);
not I_6949 (I120855,I120838);
nor I_6950 (I120872,I120855,I120821);
nor I_6951 (I120889,I120773,I120872);
DFFARX1 I_6952 (I120889,I2683,I120640,I120626,);
nor I_6953 (I120623,I120838,I120725);
DFFARX1 I_6954 (I120838,I2683,I120640,I120629,);
nor I_6955 (I120948,I120804,I767816);
nor I_6956 (I120965,I120948,I767804);
nor I_6957 (I120982,I767810,I767813);
DFFARX1 I_6958 (I120982,I2683,I120640,I121008,);
nor I_6959 (I120608,I121008,I120965);
DFFARX1 I_6960 (I121008,I2683,I120640,I121039,);
nand I_6961 (I121047,I121039,I767795);
nor I_6962 (I120632,I120674,I121047);
not I_6963 (I121078,I121008);
nand I_6964 (I121095,I121078,I767795);
nor I_6965 (I121112,I120674,I121095);
nor I_6966 (I120614,I120700,I121112);
nor I_6967 (I121143,I767810,I767807);
nor I_6968 (I121160,I120700,I121143);
DFFARX1 I_6969 (I121160,I2683,I120640,I120605,);
and I_6970 (I120620,I120773,I767810);
not I_6971 (I121235,I2690);
DFFARX1 I_6972 (I888311,I2683,I121235,I121261,);
not I_6973 (I121269,I121261);
DFFARX1 I_6974 (I888308,I2683,I121235,I121295,);
not I_6975 (I121303,I888317);
or I_6976 (I121320,I888308,I888317);
nor I_6977 (I121337,I121295,I888308);
nand I_6978 (I121212,I121303,I121337);
nor I_6979 (I121368,I888320,I888308);
nand I_6980 (I121206,I121368,I121303);
not I_6981 (I121399,I888314);
nand I_6982 (I121416,I121303,I121399);
nor I_6983 (I121433,I888311,I888329);
not I_6984 (I121450,I121433);
nor I_6985 (I121467,I121450,I121416);
nor I_6986 (I121484,I121368,I121467);
DFFARX1 I_6987 (I121484,I2683,I121235,I121221,);
nor I_6988 (I121218,I121433,I121320);
DFFARX1 I_6989 (I121433,I2683,I121235,I121224,);
nor I_6990 (I121543,I121399,I888311);
nor I_6991 (I121560,I121543,I888317);
nor I_6992 (I121577,I888332,I888326);
DFFARX1 I_6993 (I121577,I2683,I121235,I121603,);
nor I_6994 (I121203,I121603,I121560);
DFFARX1 I_6995 (I121603,I2683,I121235,I121634,);
nand I_6996 (I121642,I121634,I888323);
nor I_6997 (I121227,I121269,I121642);
not I_6998 (I121673,I121603);
nand I_6999 (I121690,I121673,I888323);
nor I_7000 (I121707,I121269,I121690);
nor I_7001 (I121209,I121295,I121707);
nor I_7002 (I121738,I888332,I888320);
nor I_7003 (I121755,I121295,I121738);
DFFARX1 I_7004 (I121755,I2683,I121235,I121200,);
and I_7005 (I121215,I121368,I888332);
not I_7006 (I121827,I2690);
DFFARX1 I_7007 (I760058,I2683,I121827,I121853,);
DFFARX1 I_7008 (I121853,I2683,I121827,I121870,);
not I_7009 (I121819,I121870);
not I_7010 (I121892,I121853);
DFFARX1 I_7011 (I760067,I2683,I121827,I121918,);
not I_7012 (I121926,I121918);
and I_7013 (I121943,I121892,I760055);
not I_7014 (I121960,I760046);
nand I_7015 (I121977,I121960,I760055);
not I_7016 (I121994,I760052);
nor I_7017 (I122011,I121994,I760070);
nand I_7018 (I122028,I122011,I760043);
nor I_7019 (I122045,I122028,I121977);
DFFARX1 I_7020 (I122045,I2683,I121827,I121795,);
not I_7021 (I122076,I122028);
not I_7022 (I122093,I760070);
nand I_7023 (I122110,I122093,I760055);
nor I_7024 (I122127,I760070,I760046);
nand I_7025 (I121807,I121943,I122127);
nand I_7026 (I121801,I121892,I760070);
nand I_7027 (I122172,I121994,I760049);
DFFARX1 I_7028 (I122172,I2683,I121827,I121816,);
DFFARX1 I_7029 (I122172,I2683,I121827,I121810,);
not I_7030 (I122217,I760049);
nor I_7031 (I122234,I122217,I760061);
and I_7032 (I122251,I122234,I760043);
or I_7033 (I122268,I122251,I760064);
DFFARX1 I_7034 (I122268,I2683,I121827,I122294,);
nand I_7035 (I122302,I122294,I121960);
nor I_7036 (I121804,I122302,I122110);
nor I_7037 (I121798,I122294,I121926);
DFFARX1 I_7038 (I122294,I2683,I121827,I122356,);
not I_7039 (I122364,I122356);
nor I_7040 (I121813,I122364,I122076);
not I_7041 (I122422,I2690);
DFFARX1 I_7042 (I276461,I2683,I122422,I122448,);
DFFARX1 I_7043 (I122448,I2683,I122422,I122465,);
not I_7044 (I122414,I122465);
not I_7045 (I122487,I122448);
DFFARX1 I_7046 (I276476,I2683,I122422,I122513,);
not I_7047 (I122521,I122513);
and I_7048 (I122538,I122487,I276473);
not I_7049 (I122555,I276461);
nand I_7050 (I122572,I122555,I276473);
not I_7051 (I122589,I276470);
nor I_7052 (I122606,I122589,I276485);
nand I_7053 (I122623,I122606,I276482);
nor I_7054 (I122640,I122623,I122572);
DFFARX1 I_7055 (I122640,I2683,I122422,I122390,);
not I_7056 (I122671,I122623);
not I_7057 (I122688,I276485);
nand I_7058 (I122705,I122688,I276473);
nor I_7059 (I122722,I276485,I276461);
nand I_7060 (I122402,I122538,I122722);
nand I_7061 (I122396,I122487,I276485);
nand I_7062 (I122767,I122589,I276479);
DFFARX1 I_7063 (I122767,I2683,I122422,I122411,);
DFFARX1 I_7064 (I122767,I2683,I122422,I122405,);
not I_7065 (I122812,I276479);
nor I_7066 (I122829,I122812,I276467);
and I_7067 (I122846,I122829,I276488);
or I_7068 (I122863,I122846,I276464);
DFFARX1 I_7069 (I122863,I2683,I122422,I122889,);
nand I_7070 (I122897,I122889,I122555);
nor I_7071 (I122399,I122897,I122705);
nor I_7072 (I122393,I122889,I122521);
DFFARX1 I_7073 (I122889,I2683,I122422,I122951,);
not I_7074 (I122959,I122951);
nor I_7075 (I122408,I122959,I122671);
not I_7076 (I123017,I2690);
DFFARX1 I_7077 (I952466,I2683,I123017,I123043,);
DFFARX1 I_7078 (I123043,I2683,I123017,I123060,);
not I_7079 (I123009,I123060);
not I_7080 (I123082,I123043);
DFFARX1 I_7081 (I952466,I2683,I123017,I123108,);
not I_7082 (I123116,I123108);
and I_7083 (I123133,I123082,I952469);
not I_7084 (I123150,I952481);
nand I_7085 (I123167,I123150,I952469);
not I_7086 (I123184,I952487);
nor I_7087 (I123201,I123184,I952478);
nand I_7088 (I123218,I123201,I952484);
nor I_7089 (I123235,I123218,I123167);
DFFARX1 I_7090 (I123235,I2683,I123017,I122985,);
not I_7091 (I123266,I123218);
not I_7092 (I123283,I952478);
nand I_7093 (I123300,I123283,I952469);
nor I_7094 (I123317,I952478,I952481);
nand I_7095 (I122997,I123133,I123317);
nand I_7096 (I122991,I123082,I952478);
nand I_7097 (I123362,I123184,I952475);
DFFARX1 I_7098 (I123362,I2683,I123017,I123006,);
DFFARX1 I_7099 (I123362,I2683,I123017,I123000,);
not I_7100 (I123407,I952475);
nor I_7101 (I123424,I123407,I952472);
and I_7102 (I123441,I123424,I952490);
or I_7103 (I123458,I123441,I952469);
DFFARX1 I_7104 (I123458,I2683,I123017,I123484,);
nand I_7105 (I123492,I123484,I123150);
nor I_7106 (I122994,I123492,I123300);
nor I_7107 (I122988,I123484,I123116);
DFFARX1 I_7108 (I123484,I2683,I123017,I123546,);
not I_7109 (I123554,I123546);
nor I_7110 (I123003,I123554,I123266);
not I_7111 (I123612,I2690);
DFFARX1 I_7112 (I25871,I2683,I123612,I123638,);
DFFARX1 I_7113 (I123638,I2683,I123612,I123655,);
not I_7114 (I123604,I123655);
not I_7115 (I123677,I123638);
DFFARX1 I_7116 (I25847,I2683,I123612,I123703,);
not I_7117 (I123711,I123703);
and I_7118 (I123728,I123677,I25862);
not I_7119 (I123745,I25850);
nand I_7120 (I123762,I123745,I25862);
not I_7121 (I123779,I25853);
nor I_7122 (I123796,I123779,I25865);
nand I_7123 (I123813,I123796,I25856);
nor I_7124 (I123830,I123813,I123762);
DFFARX1 I_7125 (I123830,I2683,I123612,I123580,);
not I_7126 (I123861,I123813);
not I_7127 (I123878,I25865);
nand I_7128 (I123895,I123878,I25862);
nor I_7129 (I123912,I25865,I25850);
nand I_7130 (I123592,I123728,I123912);
nand I_7131 (I123586,I123677,I25865);
nand I_7132 (I123957,I123779,I25859);
DFFARX1 I_7133 (I123957,I2683,I123612,I123601,);
DFFARX1 I_7134 (I123957,I2683,I123612,I123595,);
not I_7135 (I124002,I25859);
nor I_7136 (I124019,I124002,I25850);
and I_7137 (I124036,I124019,I25847);
or I_7138 (I124053,I124036,I25868);
DFFARX1 I_7139 (I124053,I2683,I123612,I124079,);
nand I_7140 (I124087,I124079,I123745);
nor I_7141 (I123589,I124087,I123895);
nor I_7142 (I123583,I124079,I123711);
DFFARX1 I_7143 (I124079,I2683,I123612,I124141,);
not I_7144 (I124149,I124141);
nor I_7145 (I123598,I124149,I123861);
not I_7146 (I124207,I2690);
DFFARX1 I_7147 (I490217,I2683,I124207,I124233,);
DFFARX1 I_7148 (I124233,I2683,I124207,I124250,);
not I_7149 (I124199,I124250);
not I_7150 (I124272,I124233);
DFFARX1 I_7151 (I490208,I2683,I124207,I124298,);
not I_7152 (I124306,I124298);
and I_7153 (I124323,I124272,I490226);
not I_7154 (I124340,I490223);
nand I_7155 (I124357,I124340,I490226);
not I_7156 (I124374,I490202);
nor I_7157 (I124391,I124374,I490205);
nand I_7158 (I124408,I124391,I490214);
nor I_7159 (I124425,I124408,I124357);
DFFARX1 I_7160 (I124425,I2683,I124207,I124175,);
not I_7161 (I124456,I124408);
not I_7162 (I124473,I490205);
nand I_7163 (I124490,I124473,I490226);
nor I_7164 (I124507,I490205,I490223);
nand I_7165 (I124187,I124323,I124507);
nand I_7166 (I124181,I124272,I490205);
nand I_7167 (I124552,I124374,I490220);
DFFARX1 I_7168 (I124552,I2683,I124207,I124196,);
DFFARX1 I_7169 (I124552,I2683,I124207,I124190,);
not I_7170 (I124597,I490220);
nor I_7171 (I124614,I124597,I490202);
and I_7172 (I124631,I124614,I490211);
or I_7173 (I124648,I124631,I490205);
DFFARX1 I_7174 (I124648,I2683,I124207,I124674,);
nand I_7175 (I124682,I124674,I124340);
nor I_7176 (I124184,I124682,I124490);
nor I_7177 (I124178,I124674,I124306);
DFFARX1 I_7178 (I124674,I2683,I124207,I124736,);
not I_7179 (I124744,I124736);
nor I_7180 (I124193,I124744,I124456);
not I_7181 (I124802,I2690);
DFFARX1 I_7182 (I922410,I2683,I124802,I124828,);
DFFARX1 I_7183 (I124828,I2683,I124802,I124845,);
not I_7184 (I124794,I124845);
not I_7185 (I124867,I124828);
DFFARX1 I_7186 (I922410,I2683,I124802,I124893,);
not I_7187 (I124901,I124893);
and I_7188 (I124918,I124867,I922413);
not I_7189 (I124935,I922425);
nand I_7190 (I124952,I124935,I922413);
not I_7191 (I124969,I922431);
nor I_7192 (I124986,I124969,I922422);
nand I_7193 (I125003,I124986,I922428);
nor I_7194 (I125020,I125003,I124952);
DFFARX1 I_7195 (I125020,I2683,I124802,I124770,);
not I_7196 (I125051,I125003);
not I_7197 (I125068,I922422);
nand I_7198 (I125085,I125068,I922413);
nor I_7199 (I125102,I922422,I922425);
nand I_7200 (I124782,I124918,I125102);
nand I_7201 (I124776,I124867,I922422);
nand I_7202 (I125147,I124969,I922419);
DFFARX1 I_7203 (I125147,I2683,I124802,I124791,);
DFFARX1 I_7204 (I125147,I2683,I124802,I124785,);
not I_7205 (I125192,I922419);
nor I_7206 (I125209,I125192,I922416);
and I_7207 (I125226,I125209,I922434);
or I_7208 (I125243,I125226,I922413);
DFFARX1 I_7209 (I125243,I2683,I124802,I125269,);
nand I_7210 (I125277,I125269,I124935);
nor I_7211 (I124779,I125277,I125085);
nor I_7212 (I124773,I125269,I124901);
DFFARX1 I_7213 (I125269,I2683,I124802,I125331,);
not I_7214 (I125339,I125331);
nor I_7215 (I124788,I125339,I125051);
not I_7216 (I125397,I2690);
DFFARX1 I_7217 (I535876,I2683,I125397,I125423,);
DFFARX1 I_7218 (I125423,I2683,I125397,I125440,);
not I_7219 (I125389,I125440);
not I_7220 (I125462,I125423);
DFFARX1 I_7221 (I535873,I2683,I125397,I125488,);
not I_7222 (I125496,I125488);
and I_7223 (I125513,I125462,I535879);
not I_7224 (I125530,I535864);
nand I_7225 (I125547,I125530,I535879);
not I_7226 (I125564,I535867);
nor I_7227 (I125581,I125564,I535888);
nand I_7228 (I125598,I125581,I535885);
nor I_7229 (I125615,I125598,I125547);
DFFARX1 I_7230 (I125615,I2683,I125397,I125365,);
not I_7231 (I125646,I125598);
not I_7232 (I125663,I535888);
nand I_7233 (I125680,I125663,I535879);
nor I_7234 (I125697,I535888,I535864);
nand I_7235 (I125377,I125513,I125697);
nand I_7236 (I125371,I125462,I535888);
nand I_7237 (I125742,I125564,I535864);
DFFARX1 I_7238 (I125742,I2683,I125397,I125386,);
DFFARX1 I_7239 (I125742,I2683,I125397,I125380,);
not I_7240 (I125787,I535864);
nor I_7241 (I125804,I125787,I535870);
and I_7242 (I125821,I125804,I535882);
or I_7243 (I125838,I125821,I535867);
DFFARX1 I_7244 (I125838,I2683,I125397,I125864,);
nand I_7245 (I125872,I125864,I125530);
nor I_7246 (I125374,I125872,I125680);
nor I_7247 (I125368,I125864,I125496);
DFFARX1 I_7248 (I125864,I2683,I125397,I125926,);
not I_7249 (I125934,I125926);
nor I_7250 (I125383,I125934,I125646);
not I_7251 (I125992,I2690);
DFFARX1 I_7252 (I629115,I2683,I125992,I126018,);
DFFARX1 I_7253 (I126018,I2683,I125992,I126035,);
not I_7254 (I125984,I126035);
not I_7255 (I126057,I126018);
DFFARX1 I_7256 (I629109,I2683,I125992,I126083,);
not I_7257 (I126091,I126083);
and I_7258 (I126108,I126057,I629127);
not I_7259 (I126125,I629115);
nand I_7260 (I126142,I126125,I629127);
not I_7261 (I126159,I629109);
nor I_7262 (I126176,I126159,I629121);
nand I_7263 (I126193,I126176,I629112);
nor I_7264 (I126210,I126193,I126142);
DFFARX1 I_7265 (I126210,I2683,I125992,I125960,);
not I_7266 (I126241,I126193);
not I_7267 (I126258,I629121);
nand I_7268 (I126275,I126258,I629127);
nor I_7269 (I126292,I629121,I629115);
nand I_7270 (I125972,I126108,I126292);
nand I_7271 (I125966,I126057,I629121);
nand I_7272 (I126337,I126159,I629124);
DFFARX1 I_7273 (I126337,I2683,I125992,I125981,);
DFFARX1 I_7274 (I126337,I2683,I125992,I125975,);
not I_7275 (I126382,I629124);
nor I_7276 (I126399,I126382,I629130);
and I_7277 (I126416,I126399,I629112);
or I_7278 (I126433,I126416,I629118);
DFFARX1 I_7279 (I126433,I2683,I125992,I126459,);
nand I_7280 (I126467,I126459,I126125);
nor I_7281 (I125969,I126467,I126275);
nor I_7282 (I125963,I126459,I126091);
DFFARX1 I_7283 (I126459,I2683,I125992,I126521,);
not I_7284 (I126529,I126521);
nor I_7285 (I125978,I126529,I126241);
not I_7286 (I126587,I2690);
DFFARX1 I_7287 (I509288,I2683,I126587,I126613,);
DFFARX1 I_7288 (I126613,I2683,I126587,I126630,);
not I_7289 (I126579,I126630);
not I_7290 (I126652,I126613);
DFFARX1 I_7291 (I509285,I2683,I126587,I126678,);
not I_7292 (I126686,I126678);
and I_7293 (I126703,I126652,I509291);
not I_7294 (I126720,I509276);
nand I_7295 (I126737,I126720,I509291);
not I_7296 (I126754,I509279);
nor I_7297 (I126771,I126754,I509300);
nand I_7298 (I126788,I126771,I509297);
nor I_7299 (I126805,I126788,I126737);
DFFARX1 I_7300 (I126805,I2683,I126587,I126555,);
not I_7301 (I126836,I126788);
not I_7302 (I126853,I509300);
nand I_7303 (I126870,I126853,I509291);
nor I_7304 (I126887,I509300,I509276);
nand I_7305 (I126567,I126703,I126887);
nand I_7306 (I126561,I126652,I509300);
nand I_7307 (I126932,I126754,I509276);
DFFARX1 I_7308 (I126932,I2683,I126587,I126576,);
DFFARX1 I_7309 (I126932,I2683,I126587,I126570,);
not I_7310 (I126977,I509276);
nor I_7311 (I126994,I126977,I509282);
and I_7312 (I127011,I126994,I509294);
or I_7313 (I127028,I127011,I509279);
DFFARX1 I_7314 (I127028,I2683,I126587,I127054,);
nand I_7315 (I127062,I127054,I126720);
nor I_7316 (I126564,I127062,I126870);
nor I_7317 (I126558,I127054,I126686);
DFFARX1 I_7318 (I127054,I2683,I126587,I127116,);
not I_7319 (I127124,I127116);
nor I_7320 (I126573,I127124,I126836);
not I_7321 (I127182,I2690);
DFFARX1 I_7322 (I234301,I2683,I127182,I127208,);
DFFARX1 I_7323 (I127208,I2683,I127182,I127225,);
not I_7324 (I127174,I127225);
not I_7325 (I127247,I127208);
DFFARX1 I_7326 (I234316,I2683,I127182,I127273,);
not I_7327 (I127281,I127273);
and I_7328 (I127298,I127247,I234313);
not I_7329 (I127315,I234301);
nand I_7330 (I127332,I127315,I234313);
not I_7331 (I127349,I234310);
nor I_7332 (I127366,I127349,I234325);
nand I_7333 (I127383,I127366,I234322);
nor I_7334 (I127400,I127383,I127332);
DFFARX1 I_7335 (I127400,I2683,I127182,I127150,);
not I_7336 (I127431,I127383);
not I_7337 (I127448,I234325);
nand I_7338 (I127465,I127448,I234313);
nor I_7339 (I127482,I234325,I234301);
nand I_7340 (I127162,I127298,I127482);
nand I_7341 (I127156,I127247,I234325);
nand I_7342 (I127527,I127349,I234319);
DFFARX1 I_7343 (I127527,I2683,I127182,I127171,);
DFFARX1 I_7344 (I127527,I2683,I127182,I127165,);
not I_7345 (I127572,I234319);
nor I_7346 (I127589,I127572,I234307);
and I_7347 (I127606,I127589,I234328);
or I_7348 (I127623,I127606,I234304);
DFFARX1 I_7349 (I127623,I2683,I127182,I127649,);
nand I_7350 (I127657,I127649,I127315);
nor I_7351 (I127159,I127657,I127465);
nor I_7352 (I127153,I127649,I127281);
DFFARX1 I_7353 (I127649,I2683,I127182,I127711,);
not I_7354 (I127719,I127711);
nor I_7355 (I127168,I127719,I127431);
not I_7356 (I127777,I2690);
DFFARX1 I_7357 (I21128,I2683,I127777,I127803,);
DFFARX1 I_7358 (I127803,I2683,I127777,I127820,);
not I_7359 (I127769,I127820);
not I_7360 (I127842,I127803);
DFFARX1 I_7361 (I21104,I2683,I127777,I127868,);
not I_7362 (I127876,I127868);
and I_7363 (I127893,I127842,I21119);
not I_7364 (I127910,I21107);
nand I_7365 (I127927,I127910,I21119);
not I_7366 (I127944,I21110);
nor I_7367 (I127961,I127944,I21122);
nand I_7368 (I127978,I127961,I21113);
nor I_7369 (I127995,I127978,I127927);
DFFARX1 I_7370 (I127995,I2683,I127777,I127745,);
not I_7371 (I128026,I127978);
not I_7372 (I128043,I21122);
nand I_7373 (I128060,I128043,I21119);
nor I_7374 (I128077,I21122,I21107);
nand I_7375 (I127757,I127893,I128077);
nand I_7376 (I127751,I127842,I21122);
nand I_7377 (I128122,I127944,I21116);
DFFARX1 I_7378 (I128122,I2683,I127777,I127766,);
DFFARX1 I_7379 (I128122,I2683,I127777,I127760,);
not I_7380 (I128167,I21116);
nor I_7381 (I128184,I128167,I21107);
and I_7382 (I128201,I128184,I21104);
or I_7383 (I128218,I128201,I21125);
DFFARX1 I_7384 (I128218,I2683,I127777,I128244,);
nand I_7385 (I128252,I128244,I127910);
nor I_7386 (I127754,I128252,I128060);
nor I_7387 (I127748,I128244,I127876);
DFFARX1 I_7388 (I128244,I2683,I127777,I128306,);
not I_7389 (I128314,I128306);
nor I_7390 (I127763,I128314,I128026);
not I_7391 (I128372,I2690);
DFFARX1 I_7392 (I601190,I2683,I128372,I128398,);
DFFARX1 I_7393 (I128398,I2683,I128372,I128415,);
not I_7394 (I128364,I128415);
not I_7395 (I128437,I128398);
DFFARX1 I_7396 (I601187,I2683,I128372,I128463,);
not I_7397 (I128471,I128463);
and I_7398 (I128488,I128437,I601193);
not I_7399 (I128505,I601178);
nand I_7400 (I128522,I128505,I601193);
not I_7401 (I128539,I601181);
nor I_7402 (I128556,I128539,I601202);
nand I_7403 (I128573,I128556,I601199);
nor I_7404 (I128590,I128573,I128522);
DFFARX1 I_7405 (I128590,I2683,I128372,I128340,);
not I_7406 (I128621,I128573);
not I_7407 (I128638,I601202);
nand I_7408 (I128655,I128638,I601193);
nor I_7409 (I128672,I601202,I601178);
nand I_7410 (I128352,I128488,I128672);
nand I_7411 (I128346,I128437,I601202);
nand I_7412 (I128717,I128539,I601178);
DFFARX1 I_7413 (I128717,I2683,I128372,I128361,);
DFFARX1 I_7414 (I128717,I2683,I128372,I128355,);
not I_7415 (I128762,I601178);
nor I_7416 (I128779,I128762,I601184);
and I_7417 (I128796,I128779,I601196);
or I_7418 (I128813,I128796,I601181);
DFFARX1 I_7419 (I128813,I2683,I128372,I128839,);
nand I_7420 (I128847,I128839,I128505);
nor I_7421 (I128349,I128847,I128655);
nor I_7422 (I128343,I128839,I128471);
DFFARX1 I_7423 (I128839,I2683,I128372,I128901,);
not I_7424 (I128909,I128901);
nor I_7425 (I128358,I128909,I128621);
not I_7426 (I128967,I2690);
DFFARX1 I_7427 (I1005339,I2683,I128967,I128993,);
DFFARX1 I_7428 (I128993,I2683,I128967,I129010,);
not I_7429 (I128959,I129010);
not I_7430 (I129032,I128993);
DFFARX1 I_7431 (I1005351,I2683,I128967,I129058,);
not I_7432 (I129066,I129058);
and I_7433 (I129083,I129032,I1005345);
not I_7434 (I129100,I1005357);
nand I_7435 (I129117,I129100,I1005345);
not I_7436 (I129134,I1005342);
nor I_7437 (I129151,I129134,I1005354);
nand I_7438 (I129168,I129151,I1005336);
nor I_7439 (I129185,I129168,I129117);
DFFARX1 I_7440 (I129185,I2683,I128967,I128935,);
not I_7441 (I129216,I129168);
not I_7442 (I129233,I1005354);
nand I_7443 (I129250,I129233,I1005345);
nor I_7444 (I129267,I1005354,I1005357);
nand I_7445 (I128947,I129083,I129267);
nand I_7446 (I128941,I129032,I1005354);
nand I_7447 (I129312,I129134,I1005348);
DFFARX1 I_7448 (I129312,I2683,I128967,I128956,);
DFFARX1 I_7449 (I129312,I2683,I128967,I128950,);
not I_7450 (I129357,I1005348);
nor I_7451 (I129374,I129357,I1005339);
and I_7452 (I129391,I129374,I1005336);
or I_7453 (I129408,I129391,I1005360);
DFFARX1 I_7454 (I129408,I2683,I128967,I129434,);
nand I_7455 (I129442,I129434,I129100);
nor I_7456 (I128944,I129442,I129250);
nor I_7457 (I128938,I129434,I129066);
DFFARX1 I_7458 (I129434,I2683,I128967,I129496,);
not I_7459 (I129504,I129496);
nor I_7460 (I128953,I129504,I129216);
not I_7461 (I129562,I2690);
DFFARX1 I_7462 (I388906,I2683,I129562,I129588,);
DFFARX1 I_7463 (I129588,I2683,I129562,I129605,);
not I_7464 (I129554,I129605);
not I_7465 (I129627,I129588);
DFFARX1 I_7466 (I388894,I2683,I129562,I129653,);
not I_7467 (I129661,I129653);
and I_7468 (I129678,I129627,I388903);
not I_7469 (I129695,I388900);
nand I_7470 (I129712,I129695,I388903);
not I_7471 (I129729,I388891);
nor I_7472 (I129746,I129729,I388897);
nand I_7473 (I129763,I129746,I388882);
nor I_7474 (I129780,I129763,I129712);
DFFARX1 I_7475 (I129780,I2683,I129562,I129530,);
not I_7476 (I129811,I129763);
not I_7477 (I129828,I388897);
nand I_7478 (I129845,I129828,I388903);
nor I_7479 (I129862,I388897,I388900);
nand I_7480 (I129542,I129678,I129862);
nand I_7481 (I129536,I129627,I388897);
nand I_7482 (I129907,I129729,I388882);
DFFARX1 I_7483 (I129907,I2683,I129562,I129551,);
DFFARX1 I_7484 (I129907,I2683,I129562,I129545,);
not I_7485 (I129952,I388882);
nor I_7486 (I129969,I129952,I388888);
and I_7487 (I129986,I129969,I388885);
or I_7488 (I130003,I129986,I388909);
DFFARX1 I_7489 (I130003,I2683,I129562,I130029,);
nand I_7490 (I130037,I130029,I129695);
nor I_7491 (I129539,I130037,I129845);
nor I_7492 (I129533,I130029,I129661);
DFFARX1 I_7493 (I130029,I2683,I129562,I130091,);
not I_7494 (I130099,I130091);
nor I_7495 (I129548,I130099,I129811);
not I_7496 (I130157,I2690);
DFFARX1 I_7497 (I926456,I2683,I130157,I130183,);
DFFARX1 I_7498 (I130183,I2683,I130157,I130200,);
not I_7499 (I130149,I130200);
not I_7500 (I130222,I130183);
DFFARX1 I_7501 (I926456,I2683,I130157,I130248,);
not I_7502 (I130256,I130248);
and I_7503 (I130273,I130222,I926459);
not I_7504 (I130290,I926471);
nand I_7505 (I130307,I130290,I926459);
not I_7506 (I130324,I926477);
nor I_7507 (I130341,I130324,I926468);
nand I_7508 (I130358,I130341,I926474);
nor I_7509 (I130375,I130358,I130307);
DFFARX1 I_7510 (I130375,I2683,I130157,I130125,);
not I_7511 (I130406,I130358);
not I_7512 (I130423,I926468);
nand I_7513 (I130440,I130423,I926459);
nor I_7514 (I130457,I926468,I926471);
nand I_7515 (I130137,I130273,I130457);
nand I_7516 (I130131,I130222,I926468);
nand I_7517 (I130502,I130324,I926465);
DFFARX1 I_7518 (I130502,I2683,I130157,I130146,);
DFFARX1 I_7519 (I130502,I2683,I130157,I130140,);
not I_7520 (I130547,I926465);
nor I_7521 (I130564,I130547,I926462);
and I_7522 (I130581,I130564,I926480);
or I_7523 (I130598,I130581,I926459);
DFFARX1 I_7524 (I130598,I2683,I130157,I130624,);
nand I_7525 (I130632,I130624,I130290);
nor I_7526 (I130134,I130632,I130440);
nor I_7527 (I130128,I130624,I130256);
DFFARX1 I_7528 (I130624,I2683,I130157,I130686,);
not I_7529 (I130694,I130686);
nor I_7530 (I130143,I130694,I130406);
not I_7531 (I130752,I2690);
DFFARX1 I_7532 (I691828,I2683,I130752,I130778,);
DFFARX1 I_7533 (I130778,I2683,I130752,I130795,);
not I_7534 (I130744,I130795);
not I_7535 (I130817,I130778);
DFFARX1 I_7536 (I691822,I2683,I130752,I130843,);
not I_7537 (I130851,I130843);
and I_7538 (I130868,I130817,I691840);
not I_7539 (I130885,I691828);
nand I_7540 (I130902,I130885,I691840);
not I_7541 (I130919,I691822);
nor I_7542 (I130936,I130919,I691834);
nand I_7543 (I130953,I130936,I691825);
nor I_7544 (I130970,I130953,I130902);
DFFARX1 I_7545 (I130970,I2683,I130752,I130720,);
not I_7546 (I131001,I130953);
not I_7547 (I131018,I691834);
nand I_7548 (I131035,I131018,I691840);
nor I_7549 (I131052,I691834,I691828);
nand I_7550 (I130732,I130868,I131052);
nand I_7551 (I130726,I130817,I691834);
nand I_7552 (I131097,I130919,I691837);
DFFARX1 I_7553 (I131097,I2683,I130752,I130741,);
DFFARX1 I_7554 (I131097,I2683,I130752,I130735,);
not I_7555 (I131142,I691837);
nor I_7556 (I131159,I131142,I691843);
and I_7557 (I131176,I131159,I691825);
or I_7558 (I131193,I131176,I691831);
DFFARX1 I_7559 (I131193,I2683,I130752,I131219,);
nand I_7560 (I131227,I131219,I130885);
nor I_7561 (I130729,I131227,I131035);
nor I_7562 (I130723,I131219,I130851);
DFFARX1 I_7563 (I131219,I2683,I130752,I131281,);
not I_7564 (I131289,I131281);
nor I_7565 (I130738,I131289,I131001);
not I_7566 (I131347,I2690);
DFFARX1 I_7567 (I86988,I2683,I131347,I131373,);
DFFARX1 I_7568 (I131373,I2683,I131347,I131390,);
not I_7569 (I131339,I131390);
not I_7570 (I131412,I131373);
DFFARX1 I_7571 (I86982,I2683,I131347,I131438,);
not I_7572 (I131446,I131438);
and I_7573 (I131463,I131412,I86979);
not I_7574 (I131480,I87000);
nand I_7575 (I131497,I131480,I86979);
not I_7576 (I131514,I86994);
nor I_7577 (I131531,I131514,I86985);
nand I_7578 (I131548,I131531,I86991);
nor I_7579 (I131565,I131548,I131497);
DFFARX1 I_7580 (I131565,I2683,I131347,I131315,);
not I_7581 (I131596,I131548);
not I_7582 (I131613,I86985);
nand I_7583 (I131630,I131613,I86979);
nor I_7584 (I131647,I86985,I87000);
nand I_7585 (I131327,I131463,I131647);
nand I_7586 (I131321,I131412,I86985);
nand I_7587 (I131692,I131514,I86979);
DFFARX1 I_7588 (I131692,I2683,I131347,I131336,);
DFFARX1 I_7589 (I131692,I2683,I131347,I131330,);
not I_7590 (I131737,I86979);
nor I_7591 (I131754,I131737,I86997);
and I_7592 (I131771,I131754,I87003);
or I_7593 (I131788,I131771,I86982);
DFFARX1 I_7594 (I131788,I2683,I131347,I131814,);
nand I_7595 (I131822,I131814,I131480);
nor I_7596 (I131324,I131822,I131630);
nor I_7597 (I131318,I131814,I131446);
DFFARX1 I_7598 (I131814,I2683,I131347,I131876,);
not I_7599 (I131884,I131876);
nor I_7600 (I131333,I131884,I131596);
not I_7601 (I131942,I2690);
DFFARX1 I_7602 (I827638,I2683,I131942,I131968,);
DFFARX1 I_7603 (I131968,I2683,I131942,I131985,);
not I_7604 (I131934,I131985);
not I_7605 (I132007,I131968);
DFFARX1 I_7606 (I827647,I2683,I131942,I132033,);
not I_7607 (I132041,I132033);
and I_7608 (I132058,I132007,I827641);
not I_7609 (I132075,I827635);
nand I_7610 (I132092,I132075,I827641);
not I_7611 (I132109,I827650);
nor I_7612 (I132126,I132109,I827638);
nand I_7613 (I132143,I132126,I827644);
nor I_7614 (I132160,I132143,I132092);
DFFARX1 I_7615 (I132160,I2683,I131942,I131910,);
not I_7616 (I132191,I132143);
not I_7617 (I132208,I827638);
nand I_7618 (I132225,I132208,I827641);
nor I_7619 (I132242,I827638,I827635);
nand I_7620 (I131922,I132058,I132242);
nand I_7621 (I131916,I132007,I827638);
nand I_7622 (I132287,I132109,I827641);
DFFARX1 I_7623 (I132287,I2683,I131942,I131931,);
DFFARX1 I_7624 (I132287,I2683,I131942,I131925,);
not I_7625 (I132332,I827641);
nor I_7626 (I132349,I132332,I827656);
and I_7627 (I132366,I132349,I827653);
or I_7628 (I132383,I132366,I827635);
DFFARX1 I_7629 (I132383,I2683,I131942,I132409,);
nand I_7630 (I132417,I132409,I132075);
nor I_7631 (I131919,I132417,I132225);
nor I_7632 (I131913,I132409,I132041);
DFFARX1 I_7633 (I132409,I2683,I131942,I132471,);
not I_7634 (I132479,I132471);
nor I_7635 (I131928,I132479,I132191);
not I_7636 (I132537,I2690);
DFFARX1 I_7637 (I508132,I2683,I132537,I132563,);
DFFARX1 I_7638 (I132563,I2683,I132537,I132580,);
not I_7639 (I132529,I132580);
not I_7640 (I132602,I132563);
DFFARX1 I_7641 (I508129,I2683,I132537,I132628,);
not I_7642 (I132636,I132628);
and I_7643 (I132653,I132602,I508135);
not I_7644 (I132670,I508120);
nand I_7645 (I132687,I132670,I508135);
not I_7646 (I132704,I508123);
nor I_7647 (I132721,I132704,I508144);
nand I_7648 (I132738,I132721,I508141);
nor I_7649 (I132755,I132738,I132687);
DFFARX1 I_7650 (I132755,I2683,I132537,I132505,);
not I_7651 (I132786,I132738);
not I_7652 (I132803,I508144);
nand I_7653 (I132820,I132803,I508135);
nor I_7654 (I132837,I508144,I508120);
nand I_7655 (I132517,I132653,I132837);
nand I_7656 (I132511,I132602,I508144);
nand I_7657 (I132882,I132704,I508120);
DFFARX1 I_7658 (I132882,I2683,I132537,I132526,);
DFFARX1 I_7659 (I132882,I2683,I132537,I132520,);
not I_7660 (I132927,I508120);
nor I_7661 (I132944,I132927,I508126);
and I_7662 (I132961,I132944,I508138);
or I_7663 (I132978,I132961,I508123);
DFFARX1 I_7664 (I132978,I2683,I132537,I133004,);
nand I_7665 (I133012,I133004,I132670);
nor I_7666 (I132514,I133012,I132820);
nor I_7667 (I132508,I133004,I132636);
DFFARX1 I_7668 (I133004,I2683,I132537,I133066,);
not I_7669 (I133074,I133066);
nor I_7670 (I132523,I133074,I132786);
not I_7671 (I133132,I2690);
DFFARX1 I_7672 (I536454,I2683,I133132,I133158,);
DFFARX1 I_7673 (I133158,I2683,I133132,I133175,);
not I_7674 (I133124,I133175);
not I_7675 (I133197,I133158);
DFFARX1 I_7676 (I536451,I2683,I133132,I133223,);
not I_7677 (I133231,I133223);
and I_7678 (I133248,I133197,I536457);
not I_7679 (I133265,I536442);
nand I_7680 (I133282,I133265,I536457);
not I_7681 (I133299,I536445);
nor I_7682 (I133316,I133299,I536466);
nand I_7683 (I133333,I133316,I536463);
nor I_7684 (I133350,I133333,I133282);
DFFARX1 I_7685 (I133350,I2683,I133132,I133100,);
not I_7686 (I133381,I133333);
not I_7687 (I133398,I536466);
nand I_7688 (I133415,I133398,I536457);
nor I_7689 (I133432,I536466,I536442);
nand I_7690 (I133112,I133248,I133432);
nand I_7691 (I133106,I133197,I536466);
nand I_7692 (I133477,I133299,I536442);
DFFARX1 I_7693 (I133477,I2683,I133132,I133121,);
DFFARX1 I_7694 (I133477,I2683,I133132,I133115,);
not I_7695 (I133522,I536442);
nor I_7696 (I133539,I133522,I536448);
and I_7697 (I133556,I133539,I536460);
or I_7698 (I133573,I133556,I536445);
DFFARX1 I_7699 (I133573,I2683,I133132,I133599,);
nand I_7700 (I133607,I133599,I133265);
nor I_7701 (I133109,I133607,I133415);
nor I_7702 (I133103,I133599,I133231);
DFFARX1 I_7703 (I133599,I2683,I133132,I133661,);
not I_7704 (I133669,I133661);
nor I_7705 (I133118,I133669,I133381);
not I_7706 (I133727,I2690);
DFFARX1 I_7707 (I533564,I2683,I133727,I133753,);
DFFARX1 I_7708 (I133753,I2683,I133727,I133770,);
not I_7709 (I133719,I133770);
not I_7710 (I133792,I133753);
DFFARX1 I_7711 (I533561,I2683,I133727,I133818,);
not I_7712 (I133826,I133818);
and I_7713 (I133843,I133792,I533567);
not I_7714 (I133860,I533552);
nand I_7715 (I133877,I133860,I533567);
not I_7716 (I133894,I533555);
nor I_7717 (I133911,I133894,I533576);
nand I_7718 (I133928,I133911,I533573);
nor I_7719 (I133945,I133928,I133877);
DFFARX1 I_7720 (I133945,I2683,I133727,I133695,);
not I_7721 (I133976,I133928);
not I_7722 (I133993,I533576);
nand I_7723 (I134010,I133993,I533567);
nor I_7724 (I134027,I533576,I533552);
nand I_7725 (I133707,I133843,I134027);
nand I_7726 (I133701,I133792,I533576);
nand I_7727 (I134072,I133894,I533552);
DFFARX1 I_7728 (I134072,I2683,I133727,I133716,);
DFFARX1 I_7729 (I134072,I2683,I133727,I133710,);
not I_7730 (I134117,I533552);
nor I_7731 (I134134,I134117,I533558);
and I_7732 (I134151,I134134,I533570);
or I_7733 (I134168,I134151,I533555);
DFFARX1 I_7734 (I134168,I2683,I133727,I134194,);
nand I_7735 (I134202,I134194,I133860);
nor I_7736 (I133704,I134202,I134010);
nor I_7737 (I133698,I134194,I133826);
DFFARX1 I_7738 (I134194,I2683,I133727,I134256,);
not I_7739 (I134264,I134256);
nor I_7740 (I133713,I134264,I133976);
not I_7741 (I134322,I2690);
DFFARX1 I_7742 (I604658,I2683,I134322,I134348,);
DFFARX1 I_7743 (I134348,I2683,I134322,I134365,);
not I_7744 (I134314,I134365);
not I_7745 (I134387,I134348);
DFFARX1 I_7746 (I604655,I2683,I134322,I134413,);
not I_7747 (I134421,I134413);
and I_7748 (I134438,I134387,I604661);
not I_7749 (I134455,I604646);
nand I_7750 (I134472,I134455,I604661);
not I_7751 (I134489,I604649);
nor I_7752 (I134506,I134489,I604670);
nand I_7753 (I134523,I134506,I604667);
nor I_7754 (I134540,I134523,I134472);
DFFARX1 I_7755 (I134540,I2683,I134322,I134290,);
not I_7756 (I134571,I134523);
not I_7757 (I134588,I604670);
nand I_7758 (I134605,I134588,I604661);
nor I_7759 (I134622,I604670,I604646);
nand I_7760 (I134302,I134438,I134622);
nand I_7761 (I134296,I134387,I604670);
nand I_7762 (I134667,I134489,I604646);
DFFARX1 I_7763 (I134667,I2683,I134322,I134311,);
DFFARX1 I_7764 (I134667,I2683,I134322,I134305,);
not I_7765 (I134712,I604646);
nor I_7766 (I134729,I134712,I604652);
and I_7767 (I134746,I134729,I604664);
or I_7768 (I134763,I134746,I604649);
DFFARX1 I_7769 (I134763,I2683,I134322,I134789,);
nand I_7770 (I134797,I134789,I134455);
nor I_7771 (I134299,I134797,I134605);
nor I_7772 (I134293,I134789,I134421);
DFFARX1 I_7773 (I134789,I2683,I134322,I134851,);
not I_7774 (I134859,I134851);
nor I_7775 (I134308,I134859,I134571);
not I_7776 (I134917,I2690);
DFFARX1 I_7777 (I366602,I2683,I134917,I134943,);
DFFARX1 I_7778 (I134943,I2683,I134917,I134960,);
not I_7779 (I134909,I134960);
not I_7780 (I134982,I134943);
DFFARX1 I_7781 (I366590,I2683,I134917,I135008,);
not I_7782 (I135016,I135008);
and I_7783 (I135033,I134982,I366599);
not I_7784 (I135050,I366596);
nand I_7785 (I135067,I135050,I366599);
not I_7786 (I135084,I366587);
nor I_7787 (I135101,I135084,I366593);
nand I_7788 (I135118,I135101,I366578);
nor I_7789 (I135135,I135118,I135067);
DFFARX1 I_7790 (I135135,I2683,I134917,I134885,);
not I_7791 (I135166,I135118);
not I_7792 (I135183,I366593);
nand I_7793 (I135200,I135183,I366599);
nor I_7794 (I135217,I366593,I366596);
nand I_7795 (I134897,I135033,I135217);
nand I_7796 (I134891,I134982,I366593);
nand I_7797 (I135262,I135084,I366578);
DFFARX1 I_7798 (I135262,I2683,I134917,I134906,);
DFFARX1 I_7799 (I135262,I2683,I134917,I134900,);
not I_7800 (I135307,I366578);
nor I_7801 (I135324,I135307,I366584);
and I_7802 (I135341,I135324,I366581);
or I_7803 (I135358,I135341,I366605);
DFFARX1 I_7804 (I135358,I2683,I134917,I135384,);
nand I_7805 (I135392,I135384,I135050);
nor I_7806 (I134894,I135392,I135200);
nor I_7807 (I134888,I135384,I135016);
DFFARX1 I_7808 (I135384,I2683,I134917,I135446,);
not I_7809 (I135454,I135446);
nor I_7810 (I134903,I135454,I135166);
not I_7811 (I135512,I2690);
DFFARX1 I_7812 (I637020,I2683,I135512,I135538,);
DFFARX1 I_7813 (I135538,I2683,I135512,I135555,);
not I_7814 (I135504,I135555);
not I_7815 (I135577,I135538);
DFFARX1 I_7816 (I637014,I2683,I135512,I135603,);
not I_7817 (I135611,I135603);
and I_7818 (I135628,I135577,I637032);
not I_7819 (I135645,I637020);
nand I_7820 (I135662,I135645,I637032);
not I_7821 (I135679,I637014);
nor I_7822 (I135696,I135679,I637026);
nand I_7823 (I135713,I135696,I637017);
nor I_7824 (I135730,I135713,I135662);
DFFARX1 I_7825 (I135730,I2683,I135512,I135480,);
not I_7826 (I135761,I135713);
not I_7827 (I135778,I637026);
nand I_7828 (I135795,I135778,I637032);
nor I_7829 (I135812,I637026,I637020);
nand I_7830 (I135492,I135628,I135812);
nand I_7831 (I135486,I135577,I637026);
nand I_7832 (I135857,I135679,I637029);
DFFARX1 I_7833 (I135857,I2683,I135512,I135501,);
DFFARX1 I_7834 (I135857,I2683,I135512,I135495,);
not I_7835 (I135902,I637029);
nor I_7836 (I135919,I135902,I637035);
and I_7837 (I135936,I135919,I637017);
or I_7838 (I135953,I135936,I637023);
DFFARX1 I_7839 (I135953,I2683,I135512,I135979,);
nand I_7840 (I135987,I135979,I135645);
nor I_7841 (I135489,I135987,I135795);
nor I_7842 (I135483,I135979,I135611);
DFFARX1 I_7843 (I135979,I2683,I135512,I136041,);
not I_7844 (I136049,I136041);
nor I_7845 (I135498,I136049,I135761);
not I_7846 (I136107,I2690);
DFFARX1 I_7847 (I787836,I2683,I136107,I136133,);
DFFARX1 I_7848 (I136133,I2683,I136107,I136150,);
not I_7849 (I136099,I136150);
not I_7850 (I136172,I136133);
DFFARX1 I_7851 (I787845,I2683,I136107,I136198,);
not I_7852 (I136206,I136198);
and I_7853 (I136223,I136172,I787833);
not I_7854 (I136240,I787824);
nand I_7855 (I136257,I136240,I787833);
not I_7856 (I136274,I787830);
nor I_7857 (I136291,I136274,I787848);
nand I_7858 (I136308,I136291,I787821);
nor I_7859 (I136325,I136308,I136257);
DFFARX1 I_7860 (I136325,I2683,I136107,I136075,);
not I_7861 (I136356,I136308);
not I_7862 (I136373,I787848);
nand I_7863 (I136390,I136373,I787833);
nor I_7864 (I136407,I787848,I787824);
nand I_7865 (I136087,I136223,I136407);
nand I_7866 (I136081,I136172,I787848);
nand I_7867 (I136452,I136274,I787827);
DFFARX1 I_7868 (I136452,I2683,I136107,I136096,);
DFFARX1 I_7869 (I136452,I2683,I136107,I136090,);
not I_7870 (I136497,I787827);
nor I_7871 (I136514,I136497,I787839);
and I_7872 (I136531,I136514,I787821);
or I_7873 (I136548,I136531,I787842);
DFFARX1 I_7874 (I136548,I2683,I136107,I136574,);
nand I_7875 (I136582,I136574,I136240);
nor I_7876 (I136084,I136582,I136390);
nor I_7877 (I136078,I136574,I136206);
DFFARX1 I_7878 (I136574,I2683,I136107,I136636,);
not I_7879 (I136644,I136636);
nor I_7880 (I136093,I136644,I136356);
not I_7881 (I136702,I2690);
DFFARX1 I_7882 (I635439,I2683,I136702,I136728,);
DFFARX1 I_7883 (I136728,I2683,I136702,I136745,);
not I_7884 (I136694,I136745);
not I_7885 (I136767,I136728);
DFFARX1 I_7886 (I635433,I2683,I136702,I136793,);
not I_7887 (I136801,I136793);
and I_7888 (I136818,I136767,I635451);
not I_7889 (I136835,I635439);
nand I_7890 (I136852,I136835,I635451);
not I_7891 (I136869,I635433);
nor I_7892 (I136886,I136869,I635445);
nand I_7893 (I136903,I136886,I635436);
nor I_7894 (I136920,I136903,I136852);
DFFARX1 I_7895 (I136920,I2683,I136702,I136670,);
not I_7896 (I136951,I136903);
not I_7897 (I136968,I635445);
nand I_7898 (I136985,I136968,I635451);
nor I_7899 (I137002,I635445,I635439);
nand I_7900 (I136682,I136818,I137002);
nand I_7901 (I136676,I136767,I635445);
nand I_7902 (I137047,I136869,I635448);
DFFARX1 I_7903 (I137047,I2683,I136702,I136691,);
DFFARX1 I_7904 (I137047,I2683,I136702,I136685,);
not I_7905 (I137092,I635448);
nor I_7906 (I137109,I137092,I635454);
and I_7907 (I137126,I137109,I635436);
or I_7908 (I137143,I137126,I635442);
DFFARX1 I_7909 (I137143,I2683,I136702,I137169,);
nand I_7910 (I137177,I137169,I136835);
nor I_7911 (I136679,I137177,I136985);
nor I_7912 (I136673,I137169,I136801);
DFFARX1 I_7913 (I137169,I2683,I136702,I137231,);
not I_7914 (I137239,I137231);
nor I_7915 (I136688,I137239,I136951);
not I_7916 (I137297,I2690);
DFFARX1 I_7917 (I858830,I2683,I137297,I137323,);
DFFARX1 I_7918 (I137323,I2683,I137297,I137340,);
not I_7919 (I137289,I137340);
not I_7920 (I137362,I137323);
DFFARX1 I_7921 (I858830,I2683,I137297,I137388,);
not I_7922 (I137396,I137388);
and I_7923 (I137413,I137362,I858833);
not I_7924 (I137430,I858845);
nand I_7925 (I137447,I137430,I858833);
not I_7926 (I137464,I858851);
nor I_7927 (I137481,I137464,I858842);
nand I_7928 (I137498,I137481,I858848);
nor I_7929 (I137515,I137498,I137447);
DFFARX1 I_7930 (I137515,I2683,I137297,I137265,);
not I_7931 (I137546,I137498);
not I_7932 (I137563,I858842);
nand I_7933 (I137580,I137563,I858833);
nor I_7934 (I137597,I858842,I858845);
nand I_7935 (I137277,I137413,I137597);
nand I_7936 (I137271,I137362,I858842);
nand I_7937 (I137642,I137464,I858839);
DFFARX1 I_7938 (I137642,I2683,I137297,I137286,);
DFFARX1 I_7939 (I137642,I2683,I137297,I137280,);
not I_7940 (I137687,I858839);
nor I_7941 (I137704,I137687,I858836);
and I_7942 (I137721,I137704,I858854);
or I_7943 (I137738,I137721,I858833);
DFFARX1 I_7944 (I137738,I2683,I137297,I137764,);
nand I_7945 (I137772,I137764,I137430);
nor I_7946 (I137274,I137772,I137580);
nor I_7947 (I137268,I137764,I137396);
DFFARX1 I_7948 (I137764,I2683,I137297,I137826,);
not I_7949 (I137834,I137826);
nor I_7950 (I137283,I137834,I137546);
not I_7951 (I137892,I2690);
DFFARX1 I_7952 (I47463,I2683,I137892,I137918,);
DFFARX1 I_7953 (I137918,I2683,I137892,I137935,);
not I_7954 (I137884,I137935);
not I_7955 (I137957,I137918);
DFFARX1 I_7956 (I47457,I2683,I137892,I137983,);
not I_7957 (I137991,I137983);
and I_7958 (I138008,I137957,I47454);
not I_7959 (I138025,I47475);
nand I_7960 (I138042,I138025,I47454);
not I_7961 (I138059,I47469);
nor I_7962 (I138076,I138059,I47460);
nand I_7963 (I138093,I138076,I47466);
nor I_7964 (I138110,I138093,I138042);
DFFARX1 I_7965 (I138110,I2683,I137892,I137860,);
not I_7966 (I138141,I138093);
not I_7967 (I138158,I47460);
nand I_7968 (I138175,I138158,I47454);
nor I_7969 (I138192,I47460,I47475);
nand I_7970 (I137872,I138008,I138192);
nand I_7971 (I137866,I137957,I47460);
nand I_7972 (I138237,I138059,I47454);
DFFARX1 I_7973 (I138237,I2683,I137892,I137881,);
DFFARX1 I_7974 (I138237,I2683,I137892,I137875,);
not I_7975 (I138282,I47454);
nor I_7976 (I138299,I138282,I47472);
and I_7977 (I138316,I138299,I47478);
or I_7978 (I138333,I138316,I47457);
DFFARX1 I_7979 (I138333,I2683,I137892,I138359,);
nand I_7980 (I138367,I138359,I138025);
nor I_7981 (I137869,I138367,I138175);
nor I_7982 (I137863,I138359,I137991);
DFFARX1 I_7983 (I138359,I2683,I137892,I138421,);
not I_7984 (I138429,I138421);
nor I_7985 (I137878,I138429,I138141);
not I_7986 (I138487,I2690);
DFFARX1 I_7987 (I885996,I2683,I138487,I138513,);
DFFARX1 I_7988 (I138513,I2683,I138487,I138530,);
not I_7989 (I138479,I138530);
not I_7990 (I138552,I138513);
DFFARX1 I_7991 (I885996,I2683,I138487,I138578,);
not I_7992 (I138586,I138578);
and I_7993 (I138603,I138552,I885999);
not I_7994 (I138620,I886011);
nand I_7995 (I138637,I138620,I885999);
not I_7996 (I138654,I886017);
nor I_7997 (I138671,I138654,I886008);
nand I_7998 (I138688,I138671,I886014);
nor I_7999 (I138705,I138688,I138637);
DFFARX1 I_8000 (I138705,I2683,I138487,I138455,);
not I_8001 (I138736,I138688);
not I_8002 (I138753,I886008);
nand I_8003 (I138770,I138753,I885999);
nor I_8004 (I138787,I886008,I886011);
nand I_8005 (I138467,I138603,I138787);
nand I_8006 (I138461,I138552,I886008);
nand I_8007 (I138832,I138654,I886005);
DFFARX1 I_8008 (I138832,I2683,I138487,I138476,);
DFFARX1 I_8009 (I138832,I2683,I138487,I138470,);
not I_8010 (I138877,I886005);
nor I_8011 (I138894,I138877,I886002);
and I_8012 (I138911,I138894,I886020);
or I_8013 (I138928,I138911,I885999);
DFFARX1 I_8014 (I138928,I2683,I138487,I138954,);
nand I_8015 (I138962,I138954,I138620);
nor I_8016 (I138464,I138962,I138770);
nor I_8017 (I138458,I138954,I138586);
DFFARX1 I_8018 (I138954,I2683,I138487,I139016,);
not I_8019 (I139024,I139016);
nor I_8020 (I138473,I139024,I138736);
not I_8021 (I139082,I2690);
DFFARX1 I_8022 (I438775,I2683,I139082,I139108,);
DFFARX1 I_8023 (I139108,I2683,I139082,I139125,);
not I_8024 (I139074,I139125);
not I_8025 (I139147,I139108);
DFFARX1 I_8026 (I438766,I2683,I139082,I139173,);
not I_8027 (I139181,I139173);
and I_8028 (I139198,I139147,I438784);
not I_8029 (I139215,I438781);
nand I_8030 (I139232,I139215,I438784);
not I_8031 (I139249,I438760);
nor I_8032 (I139266,I139249,I438763);
nand I_8033 (I139283,I139266,I438772);
nor I_8034 (I139300,I139283,I139232);
DFFARX1 I_8035 (I139300,I2683,I139082,I139050,);
not I_8036 (I139331,I139283);
not I_8037 (I139348,I438763);
nand I_8038 (I139365,I139348,I438784);
nor I_8039 (I139382,I438763,I438781);
nand I_8040 (I139062,I139198,I139382);
nand I_8041 (I139056,I139147,I438763);
nand I_8042 (I139427,I139249,I438778);
DFFARX1 I_8043 (I139427,I2683,I139082,I139071,);
DFFARX1 I_8044 (I139427,I2683,I139082,I139065,);
not I_8045 (I139472,I438778);
nor I_8046 (I139489,I139472,I438760);
and I_8047 (I139506,I139489,I438769);
or I_8048 (I139523,I139506,I438763);
DFFARX1 I_8049 (I139523,I2683,I139082,I139549,);
nand I_8050 (I139557,I139549,I139215);
nor I_8051 (I139059,I139557,I139365);
nor I_8052 (I139053,I139549,I139181);
DFFARX1 I_8053 (I139549,I2683,I139082,I139611,);
not I_8054 (I139619,I139611);
nor I_8055 (I139068,I139619,I139331);
not I_8056 (I139677,I2690);
DFFARX1 I_8057 (I293325,I2683,I139677,I139703,);
DFFARX1 I_8058 (I139703,I2683,I139677,I139720,);
not I_8059 (I139669,I139720);
not I_8060 (I139742,I139703);
DFFARX1 I_8061 (I293340,I2683,I139677,I139768,);
not I_8062 (I139776,I139768);
and I_8063 (I139793,I139742,I293337);
not I_8064 (I139810,I293325);
nand I_8065 (I139827,I139810,I293337);
not I_8066 (I139844,I293334);
nor I_8067 (I139861,I139844,I293349);
nand I_8068 (I139878,I139861,I293346);
nor I_8069 (I139895,I139878,I139827);
DFFARX1 I_8070 (I139895,I2683,I139677,I139645,);
not I_8071 (I139926,I139878);
not I_8072 (I139943,I293349);
nand I_8073 (I139960,I139943,I293337);
nor I_8074 (I139977,I293349,I293325);
nand I_8075 (I139657,I139793,I139977);
nand I_8076 (I139651,I139742,I293349);
nand I_8077 (I140022,I139844,I293343);
DFFARX1 I_8078 (I140022,I2683,I139677,I139666,);
DFFARX1 I_8079 (I140022,I2683,I139677,I139660,);
not I_8080 (I140067,I293343);
nor I_8081 (I140084,I140067,I293331);
and I_8082 (I140101,I140084,I293352);
or I_8083 (I140118,I140101,I293328);
DFFARX1 I_8084 (I140118,I2683,I139677,I140144,);
nand I_8085 (I140152,I140144,I139810);
nor I_8086 (I139654,I140152,I139960);
nor I_8087 (I139648,I140144,I139776);
DFFARX1 I_8088 (I140144,I2683,I139677,I140206,);
not I_8089 (I140214,I140206);
nor I_8090 (I139663,I140214,I139926);
not I_8091 (I140272,I2690);
DFFARX1 I_8092 (I867500,I2683,I140272,I140298,);
DFFARX1 I_8093 (I140298,I2683,I140272,I140315,);
not I_8094 (I140264,I140315);
not I_8095 (I140337,I140298);
DFFARX1 I_8096 (I867500,I2683,I140272,I140363,);
not I_8097 (I140371,I140363);
and I_8098 (I140388,I140337,I867503);
not I_8099 (I140405,I867515);
nand I_8100 (I140422,I140405,I867503);
not I_8101 (I140439,I867521);
nor I_8102 (I140456,I140439,I867512);
nand I_8103 (I140473,I140456,I867518);
nor I_8104 (I140490,I140473,I140422);
DFFARX1 I_8105 (I140490,I2683,I140272,I140240,);
not I_8106 (I140521,I140473);
not I_8107 (I140538,I867512);
nand I_8108 (I140555,I140538,I867503);
nor I_8109 (I140572,I867512,I867515);
nand I_8110 (I140252,I140388,I140572);
nand I_8111 (I140246,I140337,I867512);
nand I_8112 (I140617,I140439,I867509);
DFFARX1 I_8113 (I140617,I2683,I140272,I140261,);
DFFARX1 I_8114 (I140617,I2683,I140272,I140255,);
not I_8115 (I140662,I867509);
nor I_8116 (I140679,I140662,I867506);
and I_8117 (I140696,I140679,I867524);
or I_8118 (I140713,I140696,I867503);
DFFARX1 I_8119 (I140713,I2683,I140272,I140739,);
nand I_8120 (I140747,I140739,I140405);
nor I_8121 (I140249,I140747,I140555);
nor I_8122 (I140243,I140739,I140371);
DFFARX1 I_8123 (I140739,I2683,I140272,I140801,);
not I_8124 (I140809,I140801);
nor I_8125 (I140258,I140809,I140521);
not I_8126 (I140867,I2690);
DFFARX1 I_8127 (I736802,I2683,I140867,I140893,);
DFFARX1 I_8128 (I140893,I2683,I140867,I140910,);
not I_8129 (I140859,I140910);
not I_8130 (I140932,I140893);
DFFARX1 I_8131 (I736811,I2683,I140867,I140958,);
not I_8132 (I140966,I140958);
and I_8133 (I140983,I140932,I736799);
not I_8134 (I141000,I736790);
nand I_8135 (I141017,I141000,I736799);
not I_8136 (I141034,I736796);
nor I_8137 (I141051,I141034,I736814);
nand I_8138 (I141068,I141051,I736787);
nor I_8139 (I141085,I141068,I141017);
DFFARX1 I_8140 (I141085,I2683,I140867,I140835,);
not I_8141 (I141116,I141068);
not I_8142 (I141133,I736814);
nand I_8143 (I141150,I141133,I736799);
nor I_8144 (I141167,I736814,I736790);
nand I_8145 (I140847,I140983,I141167);
nand I_8146 (I140841,I140932,I736814);
nand I_8147 (I141212,I141034,I736793);
DFFARX1 I_8148 (I141212,I2683,I140867,I140856,);
DFFARX1 I_8149 (I141212,I2683,I140867,I140850,);
not I_8150 (I141257,I736793);
nor I_8151 (I141274,I141257,I736805);
and I_8152 (I141291,I141274,I736787);
or I_8153 (I141308,I141291,I736808);
DFFARX1 I_8154 (I141308,I2683,I140867,I141334,);
nand I_8155 (I141342,I141334,I141000);
nor I_8156 (I140844,I141342,I141150);
nor I_8157 (I140838,I141334,I140966);
DFFARX1 I_8158 (I141334,I2683,I140867,I141396,);
not I_8159 (I141404,I141396);
nor I_8160 (I140853,I141404,I141116);
not I_8161 (I141462,I2690);
DFFARX1 I_8162 (I23763,I2683,I141462,I141488,);
DFFARX1 I_8163 (I141488,I2683,I141462,I141505,);
not I_8164 (I141454,I141505);
not I_8165 (I141527,I141488);
DFFARX1 I_8166 (I23739,I2683,I141462,I141553,);
not I_8167 (I141561,I141553);
and I_8168 (I141578,I141527,I23754);
not I_8169 (I141595,I23742);
nand I_8170 (I141612,I141595,I23754);
not I_8171 (I141629,I23745);
nor I_8172 (I141646,I141629,I23757);
nand I_8173 (I141663,I141646,I23748);
nor I_8174 (I141680,I141663,I141612);
DFFARX1 I_8175 (I141680,I2683,I141462,I141430,);
not I_8176 (I141711,I141663);
not I_8177 (I141728,I23757);
nand I_8178 (I141745,I141728,I23754);
nor I_8179 (I141762,I23757,I23742);
nand I_8180 (I141442,I141578,I141762);
nand I_8181 (I141436,I141527,I23757);
nand I_8182 (I141807,I141629,I23751);
DFFARX1 I_8183 (I141807,I2683,I141462,I141451,);
DFFARX1 I_8184 (I141807,I2683,I141462,I141445,);
not I_8185 (I141852,I23751);
nor I_8186 (I141869,I141852,I23742);
and I_8187 (I141886,I141869,I23739);
or I_8188 (I141903,I141886,I23760);
DFFARX1 I_8189 (I141903,I2683,I141462,I141929,);
nand I_8190 (I141937,I141929,I141595);
nor I_8191 (I141439,I141937,I141745);
nor I_8192 (I141433,I141929,I141561);
DFFARX1 I_8193 (I141929,I2683,I141462,I141991,);
not I_8194 (I141999,I141991);
nor I_8195 (I141448,I141999,I141711);
not I_8196 (I142057,I2690);
DFFARX1 I_8197 (I626480,I2683,I142057,I142083,);
DFFARX1 I_8198 (I142083,I2683,I142057,I142100,);
not I_8199 (I142049,I142100);
not I_8200 (I142122,I142083);
DFFARX1 I_8201 (I626474,I2683,I142057,I142148,);
not I_8202 (I142156,I142148);
and I_8203 (I142173,I142122,I626492);
not I_8204 (I142190,I626480);
nand I_8205 (I142207,I142190,I626492);
not I_8206 (I142224,I626474);
nor I_8207 (I142241,I142224,I626486);
nand I_8208 (I142258,I142241,I626477);
nor I_8209 (I142275,I142258,I142207);
DFFARX1 I_8210 (I142275,I2683,I142057,I142025,);
not I_8211 (I142306,I142258);
not I_8212 (I142323,I626486);
nand I_8213 (I142340,I142323,I626492);
nor I_8214 (I142357,I626486,I626480);
nand I_8215 (I142037,I142173,I142357);
nand I_8216 (I142031,I142122,I626486);
nand I_8217 (I142402,I142224,I626489);
DFFARX1 I_8218 (I142402,I2683,I142057,I142046,);
DFFARX1 I_8219 (I142402,I2683,I142057,I142040,);
not I_8220 (I142447,I626489);
nor I_8221 (I142464,I142447,I626495);
and I_8222 (I142481,I142464,I626477);
or I_8223 (I142498,I142481,I626483);
DFFARX1 I_8224 (I142498,I2683,I142057,I142524,);
nand I_8225 (I142532,I142524,I142190);
nor I_8226 (I142034,I142532,I142340);
nor I_8227 (I142028,I142524,I142156);
DFFARX1 I_8228 (I142524,I2683,I142057,I142586,);
not I_8229 (I142594,I142586);
nor I_8230 (I142043,I142594,I142306);
not I_8231 (I142652,I2690);
DFFARX1 I_8232 (I763934,I2683,I142652,I142678,);
DFFARX1 I_8233 (I142678,I2683,I142652,I142695,);
not I_8234 (I142644,I142695);
not I_8235 (I142717,I142678);
DFFARX1 I_8236 (I763943,I2683,I142652,I142743,);
not I_8237 (I142751,I142743);
and I_8238 (I142768,I142717,I763931);
not I_8239 (I142785,I763922);
nand I_8240 (I142802,I142785,I763931);
not I_8241 (I142819,I763928);
nor I_8242 (I142836,I142819,I763946);
nand I_8243 (I142853,I142836,I763919);
nor I_8244 (I142870,I142853,I142802);
DFFARX1 I_8245 (I142870,I2683,I142652,I142620,);
not I_8246 (I142901,I142853);
not I_8247 (I142918,I763946);
nand I_8248 (I142935,I142918,I763931);
nor I_8249 (I142952,I763946,I763922);
nand I_8250 (I142632,I142768,I142952);
nand I_8251 (I142626,I142717,I763946);
nand I_8252 (I142997,I142819,I763925);
DFFARX1 I_8253 (I142997,I2683,I142652,I142641,);
DFFARX1 I_8254 (I142997,I2683,I142652,I142635,);
not I_8255 (I143042,I763925);
nor I_8256 (I143059,I143042,I763937);
and I_8257 (I143076,I143059,I763919);
or I_8258 (I143093,I143076,I763940);
DFFARX1 I_8259 (I143093,I2683,I142652,I143119,);
nand I_8260 (I143127,I143119,I142785);
nor I_8261 (I142629,I143127,I142935);
nor I_8262 (I142623,I143119,I142751);
DFFARX1 I_8263 (I143119,I2683,I142652,I143181,);
not I_8264 (I143189,I143181);
nor I_8265 (I142638,I143189,I142901);
not I_8266 (I143247,I2690);
DFFARX1 I_8267 (I890042,I2683,I143247,I143273,);
DFFARX1 I_8268 (I143273,I2683,I143247,I143290,);
not I_8269 (I143239,I143290);
not I_8270 (I143312,I143273);
DFFARX1 I_8271 (I890042,I2683,I143247,I143338,);
not I_8272 (I143346,I143338);
and I_8273 (I143363,I143312,I890045);
not I_8274 (I143380,I890057);
nand I_8275 (I143397,I143380,I890045);
not I_8276 (I143414,I890063);
nor I_8277 (I143431,I143414,I890054);
nand I_8278 (I143448,I143431,I890060);
nor I_8279 (I143465,I143448,I143397);
DFFARX1 I_8280 (I143465,I2683,I143247,I143215,);
not I_8281 (I143496,I143448);
not I_8282 (I143513,I890054);
nand I_8283 (I143530,I143513,I890045);
nor I_8284 (I143547,I890054,I890057);
nand I_8285 (I143227,I143363,I143547);
nand I_8286 (I143221,I143312,I890054);
nand I_8287 (I143592,I143414,I890051);
DFFARX1 I_8288 (I143592,I2683,I143247,I143236,);
DFFARX1 I_8289 (I143592,I2683,I143247,I143230,);
not I_8290 (I143637,I890051);
nor I_8291 (I143654,I143637,I890048);
and I_8292 (I143671,I143654,I890066);
or I_8293 (I143688,I143671,I890045);
DFFARX1 I_8294 (I143688,I2683,I143247,I143714,);
nand I_8295 (I143722,I143714,I143380);
nor I_8296 (I143224,I143722,I143530);
nor I_8297 (I143218,I143714,I143346);
DFFARX1 I_8298 (I143714,I2683,I143247,I143776,);
not I_8299 (I143784,I143776);
nor I_8300 (I143233,I143784,I143496);
not I_8301 (I143842,I2690);
DFFARX1 I_8302 (I292798,I2683,I143842,I143868,);
DFFARX1 I_8303 (I143868,I2683,I143842,I143885,);
not I_8304 (I143834,I143885);
not I_8305 (I143907,I143868);
DFFARX1 I_8306 (I292813,I2683,I143842,I143933,);
not I_8307 (I143941,I143933);
and I_8308 (I143958,I143907,I292810);
not I_8309 (I143975,I292798);
nand I_8310 (I143992,I143975,I292810);
not I_8311 (I144009,I292807);
nor I_8312 (I144026,I144009,I292822);
nand I_8313 (I144043,I144026,I292819);
nor I_8314 (I144060,I144043,I143992);
DFFARX1 I_8315 (I144060,I2683,I143842,I143810,);
not I_8316 (I144091,I144043);
not I_8317 (I144108,I292822);
nand I_8318 (I144125,I144108,I292810);
nor I_8319 (I144142,I292822,I292798);
nand I_8320 (I143822,I143958,I144142);
nand I_8321 (I143816,I143907,I292822);
nand I_8322 (I144187,I144009,I292816);
DFFARX1 I_8323 (I144187,I2683,I143842,I143831,);
DFFARX1 I_8324 (I144187,I2683,I143842,I143825,);
not I_8325 (I144232,I292816);
nor I_8326 (I144249,I144232,I292804);
and I_8327 (I144266,I144249,I292825);
or I_8328 (I144283,I144266,I292801);
DFFARX1 I_8329 (I144283,I2683,I143842,I144309,);
nand I_8330 (I144317,I144309,I143975);
nor I_8331 (I143819,I144317,I144125);
nor I_8332 (I143813,I144309,I143941);
DFFARX1 I_8333 (I144309,I2683,I143842,I144371,);
not I_8334 (I144379,I144371);
nor I_8335 (I143828,I144379,I144091);
not I_8336 (I144437,I2690);
DFFARX1 I_8337 (I19020,I2683,I144437,I144463,);
DFFARX1 I_8338 (I144463,I2683,I144437,I144480,);
not I_8339 (I144429,I144480);
not I_8340 (I144502,I144463);
DFFARX1 I_8341 (I18996,I2683,I144437,I144528,);
not I_8342 (I144536,I144528);
and I_8343 (I144553,I144502,I19011);
not I_8344 (I144570,I18999);
nand I_8345 (I144587,I144570,I19011);
not I_8346 (I144604,I19002);
nor I_8347 (I144621,I144604,I19014);
nand I_8348 (I144638,I144621,I19005);
nor I_8349 (I144655,I144638,I144587);
DFFARX1 I_8350 (I144655,I2683,I144437,I144405,);
not I_8351 (I144686,I144638);
not I_8352 (I144703,I19014);
nand I_8353 (I144720,I144703,I19011);
nor I_8354 (I144737,I19014,I18999);
nand I_8355 (I144417,I144553,I144737);
nand I_8356 (I144411,I144502,I19014);
nand I_8357 (I144782,I144604,I19008);
DFFARX1 I_8358 (I144782,I2683,I144437,I144426,);
DFFARX1 I_8359 (I144782,I2683,I144437,I144420,);
not I_8360 (I144827,I19008);
nor I_8361 (I144844,I144827,I18999);
and I_8362 (I144861,I144844,I18996);
or I_8363 (I144878,I144861,I19017);
DFFARX1 I_8364 (I144878,I2683,I144437,I144904,);
nand I_8365 (I144912,I144904,I144570);
nor I_8366 (I144414,I144912,I144720);
nor I_8367 (I144408,I144904,I144536);
DFFARX1 I_8368 (I144904,I2683,I144437,I144966,);
not I_8369 (I144974,I144966);
nor I_8370 (I144423,I144974,I144686);
not I_8371 (I145032,I2690);
DFFARX1 I_8372 (I496572,I2683,I145032,I145058,);
DFFARX1 I_8373 (I145058,I2683,I145032,I145075,);
not I_8374 (I145024,I145075);
not I_8375 (I145097,I145058);
DFFARX1 I_8376 (I496569,I2683,I145032,I145123,);
not I_8377 (I145131,I145123);
and I_8378 (I145148,I145097,I496575);
not I_8379 (I145165,I496560);
nand I_8380 (I145182,I145165,I496575);
not I_8381 (I145199,I496563);
nor I_8382 (I145216,I145199,I496584);
nand I_8383 (I145233,I145216,I496581);
nor I_8384 (I145250,I145233,I145182);
DFFARX1 I_8385 (I145250,I2683,I145032,I145000,);
not I_8386 (I145281,I145233);
not I_8387 (I145298,I496584);
nand I_8388 (I145315,I145298,I496575);
nor I_8389 (I145332,I496584,I496560);
nand I_8390 (I145012,I145148,I145332);
nand I_8391 (I145006,I145097,I496584);
nand I_8392 (I145377,I145199,I496560);
DFFARX1 I_8393 (I145377,I2683,I145032,I145021,);
DFFARX1 I_8394 (I145377,I2683,I145032,I145015,);
not I_8395 (I145422,I496560);
nor I_8396 (I145439,I145422,I496566);
and I_8397 (I145456,I145439,I496578);
or I_8398 (I145473,I145456,I496563);
DFFARX1 I_8399 (I145473,I2683,I145032,I145499,);
nand I_8400 (I145507,I145499,I145165);
nor I_8401 (I145009,I145507,I145315);
nor I_8402 (I145003,I145499,I145131);
DFFARX1 I_8403 (I145499,I2683,I145032,I145561,);
not I_8404 (I145569,I145561);
nor I_8405 (I145018,I145569,I145281);
not I_8406 (I145627,I2690);
DFFARX1 I_8407 (I778792,I2683,I145627,I145653,);
DFFARX1 I_8408 (I145653,I2683,I145627,I145670,);
not I_8409 (I145619,I145670);
not I_8410 (I145692,I145653);
DFFARX1 I_8411 (I778801,I2683,I145627,I145718,);
not I_8412 (I145726,I145718);
and I_8413 (I145743,I145692,I778789);
not I_8414 (I145760,I778780);
nand I_8415 (I145777,I145760,I778789);
not I_8416 (I145794,I778786);
nor I_8417 (I145811,I145794,I778804);
nand I_8418 (I145828,I145811,I778777);
nor I_8419 (I145845,I145828,I145777);
DFFARX1 I_8420 (I145845,I2683,I145627,I145595,);
not I_8421 (I145876,I145828);
not I_8422 (I145893,I778804);
nand I_8423 (I145910,I145893,I778789);
nor I_8424 (I145927,I778804,I778780);
nand I_8425 (I145607,I145743,I145927);
nand I_8426 (I145601,I145692,I778804);
nand I_8427 (I145972,I145794,I778783);
DFFARX1 I_8428 (I145972,I2683,I145627,I145616,);
DFFARX1 I_8429 (I145972,I2683,I145627,I145610,);
not I_8430 (I146017,I778783);
nor I_8431 (I146034,I146017,I778795);
and I_8432 (I146051,I146034,I778777);
or I_8433 (I146068,I146051,I778798);
DFFARX1 I_8434 (I146068,I2683,I145627,I146094,);
nand I_8435 (I146102,I146094,I145760);
nor I_8436 (I145604,I146102,I145910);
nor I_8437 (I145598,I146094,I145726);
DFFARX1 I_8438 (I146094,I2683,I145627,I146156,);
not I_8439 (I146164,I146156);
nor I_8440 (I145613,I146164,I145876);
not I_8441 (I146222,I2690);
DFFARX1 I_8442 (I834554,I2683,I146222,I146248,);
DFFARX1 I_8443 (I146248,I2683,I146222,I146265,);
not I_8444 (I146214,I146265);
not I_8445 (I146287,I146248);
DFFARX1 I_8446 (I834554,I2683,I146222,I146313,);
not I_8447 (I146321,I146313);
and I_8448 (I146338,I146287,I834557);
not I_8449 (I146355,I834569);
nand I_8450 (I146372,I146355,I834557);
not I_8451 (I146389,I834575);
nor I_8452 (I146406,I146389,I834566);
nand I_8453 (I146423,I146406,I834572);
nor I_8454 (I146440,I146423,I146372);
DFFARX1 I_8455 (I146440,I2683,I146222,I146190,);
not I_8456 (I146471,I146423);
not I_8457 (I146488,I834566);
nand I_8458 (I146505,I146488,I834557);
nor I_8459 (I146522,I834566,I834569);
nand I_8460 (I146202,I146338,I146522);
nand I_8461 (I146196,I146287,I834566);
nand I_8462 (I146567,I146389,I834563);
DFFARX1 I_8463 (I146567,I2683,I146222,I146211,);
DFFARX1 I_8464 (I146567,I2683,I146222,I146205,);
not I_8465 (I146612,I834563);
nor I_8466 (I146629,I146612,I834560);
and I_8467 (I146646,I146629,I834578);
or I_8468 (I146663,I146646,I834557);
DFFARX1 I_8469 (I146663,I2683,I146222,I146689,);
nand I_8470 (I146697,I146689,I146355);
nor I_8471 (I146199,I146697,I146505);
nor I_8472 (I146193,I146689,I146321);
DFFARX1 I_8473 (I146689,I2683,I146222,I146751,);
not I_8474 (I146759,I146751);
nor I_8475 (I146208,I146759,I146471);
not I_8476 (I146817,I2690);
DFFARX1 I_8477 (I461317,I2683,I146817,I146843,);
DFFARX1 I_8478 (I146843,I2683,I146817,I146860,);
not I_8479 (I146809,I146860);
not I_8480 (I146882,I146843);
DFFARX1 I_8481 (I461308,I2683,I146817,I146908,);
not I_8482 (I146916,I146908);
and I_8483 (I146933,I146882,I461326);
not I_8484 (I146950,I461323);
nand I_8485 (I146967,I146950,I461326);
not I_8486 (I146984,I461302);
nor I_8487 (I147001,I146984,I461305);
nand I_8488 (I147018,I147001,I461314);
nor I_8489 (I147035,I147018,I146967);
DFFARX1 I_8490 (I147035,I2683,I146817,I146785,);
not I_8491 (I147066,I147018);
not I_8492 (I147083,I461305);
nand I_8493 (I147100,I147083,I461326);
nor I_8494 (I147117,I461305,I461323);
nand I_8495 (I146797,I146933,I147117);
nand I_8496 (I146791,I146882,I461305);
nand I_8497 (I147162,I146984,I461320);
DFFARX1 I_8498 (I147162,I2683,I146817,I146806,);
DFFARX1 I_8499 (I147162,I2683,I146817,I146800,);
not I_8500 (I147207,I461320);
nor I_8501 (I147224,I147207,I461302);
and I_8502 (I147241,I147224,I461311);
or I_8503 (I147258,I147241,I461305);
DFFARX1 I_8504 (I147258,I2683,I146817,I147284,);
nand I_8505 (I147292,I147284,I146950);
nor I_8506 (I146794,I147292,I147100);
nor I_8507 (I146788,I147284,I146916);
DFFARX1 I_8508 (I147284,I2683,I146817,I147346,);
not I_8509 (I147354,I147346);
nor I_8510 (I146803,I147354,I147066);
not I_8511 (I147412,I2690);
DFFARX1 I_8512 (I319818,I2683,I147412,I147438,);
DFFARX1 I_8513 (I147438,I2683,I147412,I147455,);
not I_8514 (I147404,I147455);
not I_8515 (I147477,I147438);
DFFARX1 I_8516 (I319806,I2683,I147412,I147503,);
not I_8517 (I147511,I147503);
and I_8518 (I147528,I147477,I319815);
not I_8519 (I147545,I319812);
nand I_8520 (I147562,I147545,I319815);
not I_8521 (I147579,I319803);
nor I_8522 (I147596,I147579,I319809);
nand I_8523 (I147613,I147596,I319794);
nor I_8524 (I147630,I147613,I147562);
DFFARX1 I_8525 (I147630,I2683,I147412,I147380,);
not I_8526 (I147661,I147613);
not I_8527 (I147678,I319809);
nand I_8528 (I147695,I147678,I319815);
nor I_8529 (I147712,I319809,I319812);
nand I_8530 (I147392,I147528,I147712);
nand I_8531 (I147386,I147477,I319809);
nand I_8532 (I147757,I147579,I319794);
DFFARX1 I_8533 (I147757,I2683,I147412,I147401,);
DFFARX1 I_8534 (I147757,I2683,I147412,I147395,);
not I_8535 (I147802,I319794);
nor I_8536 (I147819,I147802,I319800);
and I_8537 (I147836,I147819,I319797);
or I_8538 (I147853,I147836,I319821);
DFFARX1 I_8539 (I147853,I2683,I147412,I147879,);
nand I_8540 (I147887,I147879,I147545);
nor I_8541 (I147389,I147887,I147695);
nor I_8542 (I147383,I147879,I147511);
DFFARX1 I_8543 (I147879,I2683,I147412,I147941,);
not I_8544 (I147949,I147941);
nor I_8545 (I147398,I147949,I147661);
not I_8546 (I148007,I2690);
DFFARX1 I_8547 (I1042400,I2683,I148007,I148033,);
DFFARX1 I_8548 (I148033,I2683,I148007,I148050,);
not I_8549 (I147999,I148050);
not I_8550 (I148072,I148033);
DFFARX1 I_8551 (I1042391,I2683,I148007,I148098,);
not I_8552 (I148106,I148098);
and I_8553 (I148123,I148072,I1042385);
not I_8554 (I148140,I1042379);
nand I_8555 (I148157,I148140,I1042385);
not I_8556 (I148174,I1042406);
nor I_8557 (I148191,I148174,I1042379);
nand I_8558 (I148208,I148191,I1042403);
nor I_8559 (I148225,I148208,I148157);
DFFARX1 I_8560 (I148225,I2683,I148007,I147975,);
not I_8561 (I148256,I148208);
not I_8562 (I148273,I1042379);
nand I_8563 (I148290,I148273,I1042385);
nor I_8564 (I148307,I1042379,I1042379);
nand I_8565 (I147987,I148123,I148307);
nand I_8566 (I147981,I148072,I1042379);
nand I_8567 (I148352,I148174,I1042388);
DFFARX1 I_8568 (I148352,I2683,I148007,I147996,);
DFFARX1 I_8569 (I148352,I2683,I148007,I147990,);
not I_8570 (I148397,I1042388);
nor I_8571 (I148414,I148397,I1042394);
and I_8572 (I148431,I148414,I1042397);
or I_8573 (I148448,I148431,I1042382);
DFFARX1 I_8574 (I148448,I2683,I148007,I148474,);
nand I_8575 (I148482,I148474,I148140);
nor I_8576 (I147984,I148482,I148290);
nor I_8577 (I147978,I148474,I148106);
DFFARX1 I_8578 (I148474,I2683,I148007,I148536,);
not I_8579 (I148544,I148536);
nor I_8580 (I147993,I148544,I148256);
not I_8581 (I148602,I2690);
DFFARX1 I_8582 (I513334,I2683,I148602,I148628,);
DFFARX1 I_8583 (I148628,I2683,I148602,I148645,);
not I_8584 (I148594,I148645);
not I_8585 (I148667,I148628);
DFFARX1 I_8586 (I513331,I2683,I148602,I148693,);
not I_8587 (I148701,I148693);
and I_8588 (I148718,I148667,I513337);
not I_8589 (I148735,I513322);
nand I_8590 (I148752,I148735,I513337);
not I_8591 (I148769,I513325);
nor I_8592 (I148786,I148769,I513346);
nand I_8593 (I148803,I148786,I513343);
nor I_8594 (I148820,I148803,I148752);
DFFARX1 I_8595 (I148820,I2683,I148602,I148570,);
not I_8596 (I148851,I148803);
not I_8597 (I148868,I513346);
nand I_8598 (I148885,I148868,I513337);
nor I_8599 (I148902,I513346,I513322);
nand I_8600 (I148582,I148718,I148902);
nand I_8601 (I148576,I148667,I513346);
nand I_8602 (I148947,I148769,I513322);
DFFARX1 I_8603 (I148947,I2683,I148602,I148591,);
DFFARX1 I_8604 (I148947,I2683,I148602,I148585,);
not I_8605 (I148992,I513322);
nor I_8606 (I149009,I148992,I513328);
and I_8607 (I149026,I149009,I513340);
or I_8608 (I149043,I149026,I513325);
DFFARX1 I_8609 (I149043,I2683,I148602,I149069,);
nand I_8610 (I149077,I149069,I148735);
nor I_8611 (I148579,I149077,I148885);
nor I_8612 (I148573,I149069,I148701);
DFFARX1 I_8613 (I149069,I2683,I148602,I149131,);
not I_8614 (I149139,I149131);
nor I_8615 (I148588,I149139,I148851);
not I_8616 (I149197,I2690);
DFFARX1 I_8617 (I93839,I2683,I149197,I149223,);
DFFARX1 I_8618 (I149223,I2683,I149197,I149240,);
not I_8619 (I149189,I149240);
not I_8620 (I149262,I149223);
DFFARX1 I_8621 (I93833,I2683,I149197,I149288,);
not I_8622 (I149296,I149288);
and I_8623 (I149313,I149262,I93830);
not I_8624 (I149330,I93851);
nand I_8625 (I149347,I149330,I93830);
not I_8626 (I149364,I93845);
nor I_8627 (I149381,I149364,I93836);
nand I_8628 (I149398,I149381,I93842);
nor I_8629 (I149415,I149398,I149347);
DFFARX1 I_8630 (I149415,I2683,I149197,I149165,);
not I_8631 (I149446,I149398);
not I_8632 (I149463,I93836);
nand I_8633 (I149480,I149463,I93830);
nor I_8634 (I149497,I93836,I93851);
nand I_8635 (I149177,I149313,I149497);
nand I_8636 (I149171,I149262,I93836);
nand I_8637 (I149542,I149364,I93830);
DFFARX1 I_8638 (I149542,I2683,I149197,I149186,);
DFFARX1 I_8639 (I149542,I2683,I149197,I149180,);
not I_8640 (I149587,I93830);
nor I_8641 (I149604,I149587,I93848);
and I_8642 (I149621,I149604,I93854);
or I_8643 (I149638,I149621,I93833);
DFFARX1 I_8644 (I149638,I2683,I149197,I149664,);
nand I_8645 (I149672,I149664,I149330);
nor I_8646 (I149174,I149672,I149480);
nor I_8647 (I149168,I149664,I149296);
DFFARX1 I_8648 (I149664,I2683,I149197,I149726,);
not I_8649 (I149734,I149726);
nor I_8650 (I149183,I149734,I149446);
not I_8651 (I149792,I2690);
DFFARX1 I_8652 (I1094760,I2683,I149792,I149818,);
DFFARX1 I_8653 (I149818,I2683,I149792,I149835,);
not I_8654 (I149784,I149835);
not I_8655 (I149857,I149818);
DFFARX1 I_8656 (I1094751,I2683,I149792,I149883,);
not I_8657 (I149891,I149883);
and I_8658 (I149908,I149857,I1094745);
not I_8659 (I149925,I1094739);
nand I_8660 (I149942,I149925,I1094745);
not I_8661 (I149959,I1094766);
nor I_8662 (I149976,I149959,I1094739);
nand I_8663 (I149993,I149976,I1094763);
nor I_8664 (I150010,I149993,I149942);
DFFARX1 I_8665 (I150010,I2683,I149792,I149760,);
not I_8666 (I150041,I149993);
not I_8667 (I150058,I1094739);
nand I_8668 (I150075,I150058,I1094745);
nor I_8669 (I150092,I1094739,I1094739);
nand I_8670 (I149772,I149908,I150092);
nand I_8671 (I149766,I149857,I1094739);
nand I_8672 (I150137,I149959,I1094748);
DFFARX1 I_8673 (I150137,I2683,I149792,I149781,);
DFFARX1 I_8674 (I150137,I2683,I149792,I149775,);
not I_8675 (I150182,I1094748);
nor I_8676 (I150199,I150182,I1094754);
and I_8677 (I150216,I150199,I1094757);
or I_8678 (I150233,I150216,I1094742);
DFFARX1 I_8679 (I150233,I2683,I149792,I150259,);
nand I_8680 (I150267,I150259,I149925);
nor I_8681 (I149769,I150267,I150075);
nor I_8682 (I149763,I150259,I149891);
DFFARX1 I_8683 (I150259,I2683,I149792,I150321,);
not I_8684 (I150329,I150321);
nor I_8685 (I149778,I150329,I150041);
not I_8686 (I150387,I2690);
DFFARX1 I_8687 (I471143,I2683,I150387,I150413,);
DFFARX1 I_8688 (I150413,I2683,I150387,I150430,);
not I_8689 (I150379,I150430);
not I_8690 (I150452,I150413);
DFFARX1 I_8691 (I471134,I2683,I150387,I150478,);
not I_8692 (I150486,I150478);
and I_8693 (I150503,I150452,I471152);
not I_8694 (I150520,I471149);
nand I_8695 (I150537,I150520,I471152);
not I_8696 (I150554,I471128);
nor I_8697 (I150571,I150554,I471131);
nand I_8698 (I150588,I150571,I471140);
nor I_8699 (I150605,I150588,I150537);
DFFARX1 I_8700 (I150605,I2683,I150387,I150355,);
not I_8701 (I150636,I150588);
not I_8702 (I150653,I471131);
nand I_8703 (I150670,I150653,I471152);
nor I_8704 (I150687,I471131,I471149);
nand I_8705 (I150367,I150503,I150687);
nand I_8706 (I150361,I150452,I471131);
nand I_8707 (I150732,I150554,I471146);
DFFARX1 I_8708 (I150732,I2683,I150387,I150376,);
DFFARX1 I_8709 (I150732,I2683,I150387,I150370,);
not I_8710 (I150777,I471146);
nor I_8711 (I150794,I150777,I471128);
and I_8712 (I150811,I150794,I471137);
or I_8713 (I150828,I150811,I471131);
DFFARX1 I_8714 (I150828,I2683,I150387,I150854,);
nand I_8715 (I150862,I150854,I150520);
nor I_8716 (I150364,I150862,I150670);
nor I_8717 (I150358,I150854,I150486);
DFFARX1 I_8718 (I150854,I2683,I150387,I150916,);
not I_8719 (I150924,I150916);
nor I_8720 (I150373,I150924,I150636);
not I_8721 (I150982,I2690);
DFFARX1 I_8722 (I772332,I2683,I150982,I151008,);
DFFARX1 I_8723 (I151008,I2683,I150982,I151025,);
not I_8724 (I150974,I151025);
not I_8725 (I151047,I151008);
DFFARX1 I_8726 (I772341,I2683,I150982,I151073,);
not I_8727 (I151081,I151073);
and I_8728 (I151098,I151047,I772329);
not I_8729 (I151115,I772320);
nand I_8730 (I151132,I151115,I772329);
not I_8731 (I151149,I772326);
nor I_8732 (I151166,I151149,I772344);
nand I_8733 (I151183,I151166,I772317);
nor I_8734 (I151200,I151183,I151132);
DFFARX1 I_8735 (I151200,I2683,I150982,I150950,);
not I_8736 (I151231,I151183);
not I_8737 (I151248,I772344);
nand I_8738 (I151265,I151248,I772329);
nor I_8739 (I151282,I772344,I772320);
nand I_8740 (I150962,I151098,I151282);
nand I_8741 (I150956,I151047,I772344);
nand I_8742 (I151327,I151149,I772323);
DFFARX1 I_8743 (I151327,I2683,I150982,I150971,);
DFFARX1 I_8744 (I151327,I2683,I150982,I150965,);
not I_8745 (I151372,I772323);
nor I_8746 (I151389,I151372,I772335);
and I_8747 (I151406,I151389,I772317);
or I_8748 (I151423,I151406,I772338);
DFFARX1 I_8749 (I151423,I2683,I150982,I151449,);
nand I_8750 (I151457,I151449,I151115);
nor I_8751 (I150959,I151457,I151265);
nor I_8752 (I150953,I151449,I151081);
DFFARX1 I_8753 (I151449,I2683,I150982,I151511,);
not I_8754 (I151519,I151511);
nor I_8755 (I150968,I151519,I151231);
not I_8756 (I151577,I2690);
DFFARX1 I_8757 (I354634,I2683,I151577,I151603,);
DFFARX1 I_8758 (I151603,I2683,I151577,I151620,);
not I_8759 (I151569,I151620);
not I_8760 (I151642,I151603);
DFFARX1 I_8761 (I354622,I2683,I151577,I151668,);
not I_8762 (I151676,I151668);
and I_8763 (I151693,I151642,I354631);
not I_8764 (I151710,I354628);
nand I_8765 (I151727,I151710,I354631);
not I_8766 (I151744,I354619);
nor I_8767 (I151761,I151744,I354625);
nand I_8768 (I151778,I151761,I354610);
nor I_8769 (I151795,I151778,I151727);
DFFARX1 I_8770 (I151795,I2683,I151577,I151545,);
not I_8771 (I151826,I151778);
not I_8772 (I151843,I354625);
nand I_8773 (I151860,I151843,I354631);
nor I_8774 (I151877,I354625,I354628);
nand I_8775 (I151557,I151693,I151877);
nand I_8776 (I151551,I151642,I354625);
nand I_8777 (I151922,I151744,I354610);
DFFARX1 I_8778 (I151922,I2683,I151577,I151566,);
DFFARX1 I_8779 (I151922,I2683,I151577,I151560,);
not I_8780 (I151967,I354610);
nor I_8781 (I151984,I151967,I354616);
and I_8782 (I152001,I151984,I354613);
or I_8783 (I152018,I152001,I354637);
DFFARX1 I_8784 (I152018,I2683,I151577,I152044,);
nand I_8785 (I152052,I152044,I151710);
nor I_8786 (I151554,I152052,I151860);
nor I_8787 (I151548,I152044,I151676);
DFFARX1 I_8788 (I152044,I2683,I151577,I152106,);
not I_8789 (I152114,I152106);
nor I_8790 (I151563,I152114,I151826);
not I_8791 (I152172,I2690);
DFFARX1 I_8792 (I254854,I2683,I152172,I152198,);
DFFARX1 I_8793 (I152198,I2683,I152172,I152215,);
not I_8794 (I152164,I152215);
not I_8795 (I152237,I152198);
DFFARX1 I_8796 (I254869,I2683,I152172,I152263,);
not I_8797 (I152271,I152263);
and I_8798 (I152288,I152237,I254866);
not I_8799 (I152305,I254854);
nand I_8800 (I152322,I152305,I254866);
not I_8801 (I152339,I254863);
nor I_8802 (I152356,I152339,I254878);
nand I_8803 (I152373,I152356,I254875);
nor I_8804 (I152390,I152373,I152322);
DFFARX1 I_8805 (I152390,I2683,I152172,I152140,);
not I_8806 (I152421,I152373);
not I_8807 (I152438,I254878);
nand I_8808 (I152455,I152438,I254866);
nor I_8809 (I152472,I254878,I254854);
nand I_8810 (I152152,I152288,I152472);
nand I_8811 (I152146,I152237,I254878);
nand I_8812 (I152517,I152339,I254872);
DFFARX1 I_8813 (I152517,I2683,I152172,I152161,);
DFFARX1 I_8814 (I152517,I2683,I152172,I152155,);
not I_8815 (I152562,I254872);
nor I_8816 (I152579,I152562,I254860);
and I_8817 (I152596,I152579,I254881);
or I_8818 (I152613,I152596,I254857);
DFFARX1 I_8819 (I152613,I2683,I152172,I152639,);
nand I_8820 (I152647,I152639,I152305);
nor I_8821 (I152149,I152647,I152455);
nor I_8822 (I152143,I152639,I152271);
DFFARX1 I_8823 (I152639,I2683,I152172,I152701,);
not I_8824 (I152709,I152701);
nor I_8825 (I152158,I152709,I152421);
not I_8826 (I152767,I2690);
DFFARX1 I_8827 (I226396,I2683,I152767,I152793,);
DFFARX1 I_8828 (I152793,I2683,I152767,I152810,);
not I_8829 (I152759,I152810);
not I_8830 (I152832,I152793);
DFFARX1 I_8831 (I226411,I2683,I152767,I152858,);
not I_8832 (I152866,I152858);
and I_8833 (I152883,I152832,I226408);
not I_8834 (I152900,I226396);
nand I_8835 (I152917,I152900,I226408);
not I_8836 (I152934,I226405);
nor I_8837 (I152951,I152934,I226420);
nand I_8838 (I152968,I152951,I226417);
nor I_8839 (I152985,I152968,I152917);
DFFARX1 I_8840 (I152985,I2683,I152767,I152735,);
not I_8841 (I153016,I152968);
not I_8842 (I153033,I226420);
nand I_8843 (I153050,I153033,I226408);
nor I_8844 (I153067,I226420,I226396);
nand I_8845 (I152747,I152883,I153067);
nand I_8846 (I152741,I152832,I226420);
nand I_8847 (I153112,I152934,I226414);
DFFARX1 I_8848 (I153112,I2683,I152767,I152756,);
DFFARX1 I_8849 (I153112,I2683,I152767,I152750,);
not I_8850 (I153157,I226414);
nor I_8851 (I153174,I153157,I226402);
and I_8852 (I153191,I153174,I226423);
or I_8853 (I153208,I153191,I226399);
DFFARX1 I_8854 (I153208,I2683,I152767,I153234,);
nand I_8855 (I153242,I153234,I152900);
nor I_8856 (I152744,I153242,I153050);
nor I_8857 (I152738,I153234,I152866);
DFFARX1 I_8858 (I153234,I2683,I152767,I153296,);
not I_8859 (I153304,I153296);
nor I_8860 (I152753,I153304,I153016);
not I_8861 (I153362,I2690);
DFFARX1 I_8862 (I418134,I2683,I153362,I153388,);
DFFARX1 I_8863 (I153388,I2683,I153362,I153405,);
not I_8864 (I153354,I153405);
not I_8865 (I153427,I153388);
DFFARX1 I_8866 (I418128,I2683,I153362,I153453,);
not I_8867 (I153461,I153453);
and I_8868 (I153478,I153427,I418143);
not I_8869 (I153495,I418140);
nand I_8870 (I153512,I153495,I418143);
not I_8871 (I153529,I418131);
nor I_8872 (I153546,I153529,I418122);
nand I_8873 (I153563,I153546,I418125);
nor I_8874 (I153580,I153563,I153512);
DFFARX1 I_8875 (I153580,I2683,I153362,I153330,);
not I_8876 (I153611,I153563);
not I_8877 (I153628,I418122);
nand I_8878 (I153645,I153628,I418143);
nor I_8879 (I153662,I418122,I418140);
nand I_8880 (I153342,I153478,I153662);
nand I_8881 (I153336,I153427,I418122);
nand I_8882 (I153707,I153529,I418146);
DFFARX1 I_8883 (I153707,I2683,I153362,I153351,);
DFFARX1 I_8884 (I153707,I2683,I153362,I153345,);
not I_8885 (I153752,I418146);
nor I_8886 (I153769,I153752,I418137);
and I_8887 (I153786,I153769,I418122);
or I_8888 (I153803,I153786,I418125);
DFFARX1 I_8889 (I153803,I2683,I153362,I153829,);
nand I_8890 (I153837,I153829,I153495);
nor I_8891 (I153339,I153837,I153645);
nor I_8892 (I153333,I153829,I153461);
DFFARX1 I_8893 (I153829,I2683,I153362,I153891,);
not I_8894 (I153899,I153891);
nor I_8895 (I153348,I153899,I153611);
not I_8896 (I153957,I2690);
DFFARX1 I_8897 (I857674,I2683,I153957,I153983,);
DFFARX1 I_8898 (I153983,I2683,I153957,I154000,);
not I_8899 (I153949,I154000);
not I_8900 (I154022,I153983);
DFFARX1 I_8901 (I857674,I2683,I153957,I154048,);
not I_8902 (I154056,I154048);
and I_8903 (I154073,I154022,I857677);
not I_8904 (I154090,I857689);
nand I_8905 (I154107,I154090,I857677);
not I_8906 (I154124,I857695);
nor I_8907 (I154141,I154124,I857686);
nand I_8908 (I154158,I154141,I857692);
nor I_8909 (I154175,I154158,I154107);
DFFARX1 I_8910 (I154175,I2683,I153957,I153925,);
not I_8911 (I154206,I154158);
not I_8912 (I154223,I857686);
nand I_8913 (I154240,I154223,I857677);
nor I_8914 (I154257,I857686,I857689);
nand I_8915 (I153937,I154073,I154257);
nand I_8916 (I153931,I154022,I857686);
nand I_8917 (I154302,I154124,I857683);
DFFARX1 I_8918 (I154302,I2683,I153957,I153946,);
DFFARX1 I_8919 (I154302,I2683,I153957,I153940,);
not I_8920 (I154347,I857683);
nor I_8921 (I154364,I154347,I857680);
and I_8922 (I154381,I154364,I857698);
or I_8923 (I154398,I154381,I857677);
DFFARX1 I_8924 (I154398,I2683,I153957,I154424,);
nand I_8925 (I154432,I154424,I154090);
nor I_8926 (I153934,I154432,I154240);
nor I_8927 (I153928,I154424,I154056);
DFFARX1 I_8928 (I154424,I2683,I153957,I154486,);
not I_8929 (I154494,I154486);
nor I_8930 (I153943,I154494,I154206);
not I_8931 (I154552,I2690);
DFFARX1 I_8932 (I678653,I2683,I154552,I154578,);
DFFARX1 I_8933 (I154578,I2683,I154552,I154595,);
not I_8934 (I154544,I154595);
not I_8935 (I154617,I154578);
DFFARX1 I_8936 (I678647,I2683,I154552,I154643,);
not I_8937 (I154651,I154643);
and I_8938 (I154668,I154617,I678665);
not I_8939 (I154685,I678653);
nand I_8940 (I154702,I154685,I678665);
not I_8941 (I154719,I678647);
nor I_8942 (I154736,I154719,I678659);
nand I_8943 (I154753,I154736,I678650);
nor I_8944 (I154770,I154753,I154702);
DFFARX1 I_8945 (I154770,I2683,I154552,I154520,);
not I_8946 (I154801,I154753);
not I_8947 (I154818,I678659);
nand I_8948 (I154835,I154818,I678665);
nor I_8949 (I154852,I678659,I678653);
nand I_8950 (I154532,I154668,I154852);
nand I_8951 (I154526,I154617,I678659);
nand I_8952 (I154897,I154719,I678662);
DFFARX1 I_8953 (I154897,I2683,I154552,I154541,);
DFFARX1 I_8954 (I154897,I2683,I154552,I154535,);
not I_8955 (I154942,I678662);
nor I_8956 (I154959,I154942,I678668);
and I_8957 (I154976,I154959,I678650);
or I_8958 (I154993,I154976,I678656);
DFFARX1 I_8959 (I154993,I2683,I154552,I155019,);
nand I_8960 (I155027,I155019,I154685);
nor I_8961 (I154529,I155027,I154835);
nor I_8962 (I154523,I155019,I154651);
DFFARX1 I_8963 (I155019,I2683,I154552,I155081,);
not I_8964 (I155089,I155081);
nor I_8965 (I154538,I155089,I154801);
not I_8966 (I155147,I2690);
DFFARX1 I_8967 (I1006495,I2683,I155147,I155173,);
DFFARX1 I_8968 (I155173,I2683,I155147,I155190,);
not I_8969 (I155139,I155190);
not I_8970 (I155212,I155173);
DFFARX1 I_8971 (I1006507,I2683,I155147,I155238,);
not I_8972 (I155246,I155238);
and I_8973 (I155263,I155212,I1006501);
not I_8974 (I155280,I1006513);
nand I_8975 (I155297,I155280,I1006501);
not I_8976 (I155314,I1006498);
nor I_8977 (I155331,I155314,I1006510);
nand I_8978 (I155348,I155331,I1006492);
nor I_8979 (I155365,I155348,I155297);
DFFARX1 I_8980 (I155365,I2683,I155147,I155115,);
not I_8981 (I155396,I155348);
not I_8982 (I155413,I1006510);
nand I_8983 (I155430,I155413,I1006501);
nor I_8984 (I155447,I1006510,I1006513);
nand I_8985 (I155127,I155263,I155447);
nand I_8986 (I155121,I155212,I1006510);
nand I_8987 (I155492,I155314,I1006504);
DFFARX1 I_8988 (I155492,I2683,I155147,I155136,);
DFFARX1 I_8989 (I155492,I2683,I155147,I155130,);
not I_8990 (I155537,I1006504);
nor I_8991 (I155554,I155537,I1006495);
and I_8992 (I155571,I155554,I1006492);
or I_8993 (I155588,I155571,I1006516);
DFFARX1 I_8994 (I155588,I2683,I155147,I155614,);
nand I_8995 (I155622,I155614,I155280);
nor I_8996 (I155124,I155622,I155430);
nor I_8997 (I155118,I155614,I155246);
DFFARX1 I_8998 (I155614,I2683,I155147,I155676,);
not I_8999 (I155684,I155676);
nor I_9000 (I155133,I155684,I155396);
not I_9001 (I155742,I2690);
DFFARX1 I_9002 (I1056085,I2683,I155742,I155768,);
DFFARX1 I_9003 (I155768,I2683,I155742,I155785,);
not I_9004 (I155734,I155785);
not I_9005 (I155807,I155768);
DFFARX1 I_9006 (I1056076,I2683,I155742,I155833,);
not I_9007 (I155841,I155833);
and I_9008 (I155858,I155807,I1056070);
not I_9009 (I155875,I1056064);
nand I_9010 (I155892,I155875,I1056070);
not I_9011 (I155909,I1056091);
nor I_9012 (I155926,I155909,I1056064);
nand I_9013 (I155943,I155926,I1056088);
nor I_9014 (I155960,I155943,I155892);
DFFARX1 I_9015 (I155960,I2683,I155742,I155710,);
not I_9016 (I155991,I155943);
not I_9017 (I156008,I1056064);
nand I_9018 (I156025,I156008,I1056070);
nor I_9019 (I156042,I1056064,I1056064);
nand I_9020 (I155722,I155858,I156042);
nand I_9021 (I155716,I155807,I1056064);
nand I_9022 (I156087,I155909,I1056073);
DFFARX1 I_9023 (I156087,I2683,I155742,I155731,);
DFFARX1 I_9024 (I156087,I2683,I155742,I155725,);
not I_9025 (I156132,I1056073);
nor I_9026 (I156149,I156132,I1056079);
and I_9027 (I156166,I156149,I1056082);
or I_9028 (I156183,I156166,I1056067);
DFFARX1 I_9029 (I156183,I2683,I155742,I156209,);
nand I_9030 (I156217,I156209,I155875);
nor I_9031 (I155719,I156217,I156025);
nor I_9032 (I155713,I156209,I155841);
DFFARX1 I_9033 (I156209,I2683,I155742,I156271,);
not I_9034 (I156279,I156271);
nor I_9035 (I155728,I156279,I155991);
not I_9036 (I156337,I2690);
DFFARX1 I_9037 (I320906,I2683,I156337,I156363,);
DFFARX1 I_9038 (I156363,I2683,I156337,I156380,);
not I_9039 (I156329,I156380);
not I_9040 (I156402,I156363);
DFFARX1 I_9041 (I320894,I2683,I156337,I156428,);
not I_9042 (I156436,I156428);
and I_9043 (I156453,I156402,I320903);
not I_9044 (I156470,I320900);
nand I_9045 (I156487,I156470,I320903);
not I_9046 (I156504,I320891);
nor I_9047 (I156521,I156504,I320897);
nand I_9048 (I156538,I156521,I320882);
nor I_9049 (I156555,I156538,I156487);
DFFARX1 I_9050 (I156555,I2683,I156337,I156305,);
not I_9051 (I156586,I156538);
not I_9052 (I156603,I320897);
nand I_9053 (I156620,I156603,I320903);
nor I_9054 (I156637,I320897,I320900);
nand I_9055 (I156317,I156453,I156637);
nand I_9056 (I156311,I156402,I320897);
nand I_9057 (I156682,I156504,I320882);
DFFARX1 I_9058 (I156682,I2683,I156337,I156326,);
DFFARX1 I_9059 (I156682,I2683,I156337,I156320,);
not I_9060 (I156727,I320882);
nor I_9061 (I156744,I156727,I320888);
and I_9062 (I156761,I156744,I320885);
or I_9063 (I156778,I156761,I320909);
DFFARX1 I_9064 (I156778,I2683,I156337,I156804,);
nand I_9065 (I156812,I156804,I156470);
nor I_9066 (I156314,I156812,I156620);
nor I_9067 (I156308,I156804,I156436);
DFFARX1 I_9068 (I156804,I2683,I156337,I156866,);
not I_9069 (I156874,I156866);
nor I_9070 (I156323,I156874,I156586);
not I_9071 (I156932,I2690);
DFFARX1 I_9072 (I967376,I2683,I156932,I156958,);
DFFARX1 I_9073 (I156958,I2683,I156932,I156975,);
not I_9074 (I156924,I156975);
not I_9075 (I156997,I156958);
DFFARX1 I_9076 (I967361,I2683,I156932,I157023,);
not I_9077 (I157031,I157023);
and I_9078 (I157048,I156997,I967379);
not I_9079 (I157065,I967361);
nand I_9080 (I157082,I157065,I967379);
not I_9081 (I157099,I967382);
nor I_9082 (I157116,I157099,I967373);
nand I_9083 (I157133,I157116,I967370);
nor I_9084 (I157150,I157133,I157082);
DFFARX1 I_9085 (I157150,I2683,I156932,I156900,);
not I_9086 (I157181,I157133);
not I_9087 (I157198,I967373);
nand I_9088 (I157215,I157198,I967379);
nor I_9089 (I157232,I967373,I967361);
nand I_9090 (I156912,I157048,I157232);
nand I_9091 (I156906,I156997,I967373);
nand I_9092 (I157277,I157099,I967367);
DFFARX1 I_9093 (I157277,I2683,I156932,I156921,);
DFFARX1 I_9094 (I157277,I2683,I156932,I156915,);
not I_9095 (I157322,I967367);
nor I_9096 (I157339,I157322,I967358);
and I_9097 (I157356,I157339,I967364);
or I_9098 (I157373,I157356,I967358);
DFFARX1 I_9099 (I157373,I2683,I156932,I157399,);
nand I_9100 (I157407,I157399,I157065);
nor I_9101 (I156909,I157407,I157215);
nor I_9102 (I156903,I157399,I157031);
DFFARX1 I_9103 (I157399,I2683,I156932,I157461,);
not I_9104 (I157469,I157461);
nor I_9105 (I156918,I157469,I157181);
not I_9106 (I157527,I2690);
DFFARX1 I_9107 (I412184,I2683,I157527,I157553,);
DFFARX1 I_9108 (I157553,I2683,I157527,I157570,);
not I_9109 (I157519,I157570);
not I_9110 (I157592,I157553);
DFFARX1 I_9111 (I412178,I2683,I157527,I157618,);
not I_9112 (I157626,I157618);
and I_9113 (I157643,I157592,I412193);
not I_9114 (I157660,I412190);
nand I_9115 (I157677,I157660,I412193);
not I_9116 (I157694,I412181);
nor I_9117 (I157711,I157694,I412172);
nand I_9118 (I157728,I157711,I412175);
nor I_9119 (I157745,I157728,I157677);
DFFARX1 I_9120 (I157745,I2683,I157527,I157495,);
not I_9121 (I157776,I157728);
not I_9122 (I157793,I412172);
nand I_9123 (I157810,I157793,I412193);
nor I_9124 (I157827,I412172,I412190);
nand I_9125 (I157507,I157643,I157827);
nand I_9126 (I157501,I157592,I412172);
nand I_9127 (I157872,I157694,I412196);
DFFARX1 I_9128 (I157872,I2683,I157527,I157516,);
DFFARX1 I_9129 (I157872,I2683,I157527,I157510,);
not I_9130 (I157917,I412196);
nor I_9131 (I157934,I157917,I412187);
and I_9132 (I157951,I157934,I412172);
or I_9133 (I157968,I157951,I412175);
DFFARX1 I_9134 (I157968,I2683,I157527,I157994,);
nand I_9135 (I158002,I157994,I157660);
nor I_9136 (I157504,I158002,I157810);
nor I_9137 (I157498,I157994,I157626);
DFFARX1 I_9138 (I157994,I2683,I157527,I158056,);
not I_9139 (I158064,I158056);
nor I_9140 (I157513,I158064,I157776);
not I_9141 (I158122,I2690);
DFFARX1 I_9142 (I708378,I2683,I158122,I158148,);
DFFARX1 I_9143 (I158148,I2683,I158122,I158165,);
not I_9144 (I158114,I158165);
not I_9145 (I158187,I158148);
DFFARX1 I_9146 (I708387,I2683,I158122,I158213,);
not I_9147 (I158221,I158213);
and I_9148 (I158238,I158187,I708375);
not I_9149 (I158255,I708366);
nand I_9150 (I158272,I158255,I708375);
not I_9151 (I158289,I708372);
nor I_9152 (I158306,I158289,I708390);
nand I_9153 (I158323,I158306,I708363);
nor I_9154 (I158340,I158323,I158272);
DFFARX1 I_9155 (I158340,I2683,I158122,I158090,);
not I_9156 (I158371,I158323);
not I_9157 (I158388,I708390);
nand I_9158 (I158405,I158388,I708375);
nor I_9159 (I158422,I708390,I708366);
nand I_9160 (I158102,I158238,I158422);
nand I_9161 (I158096,I158187,I708390);
nand I_9162 (I158467,I158289,I708369);
DFFARX1 I_9163 (I158467,I2683,I158122,I158111,);
DFFARX1 I_9164 (I158467,I2683,I158122,I158105,);
not I_9165 (I158512,I708369);
nor I_9166 (I158529,I158512,I708381);
and I_9167 (I158546,I158529,I708363);
or I_9168 (I158563,I158546,I708384);
DFFARX1 I_9169 (I158563,I2683,I158122,I158589,);
nand I_9170 (I158597,I158589,I158255);
nor I_9171 (I158099,I158597,I158405);
nor I_9172 (I158093,I158589,I158221);
DFFARX1 I_9173 (I158589,I2683,I158122,I158651,);
not I_9174 (I158659,I158651);
nor I_9175 (I158108,I158659,I158371);
not I_9176 (I158717,I2690);
DFFARX1 I_9177 (I375306,I2683,I158717,I158743,);
DFFARX1 I_9178 (I158743,I2683,I158717,I158760,);
not I_9179 (I158709,I158760);
not I_9180 (I158782,I158743);
DFFARX1 I_9181 (I375294,I2683,I158717,I158808,);
not I_9182 (I158816,I158808);
and I_9183 (I158833,I158782,I375303);
not I_9184 (I158850,I375300);
nand I_9185 (I158867,I158850,I375303);
not I_9186 (I158884,I375291);
nor I_9187 (I158901,I158884,I375297);
nand I_9188 (I158918,I158901,I375282);
nor I_9189 (I158935,I158918,I158867);
DFFARX1 I_9190 (I158935,I2683,I158717,I158685,);
not I_9191 (I158966,I158918);
not I_9192 (I158983,I375297);
nand I_9193 (I159000,I158983,I375303);
nor I_9194 (I159017,I375297,I375300);
nand I_9195 (I158697,I158833,I159017);
nand I_9196 (I158691,I158782,I375297);
nand I_9197 (I159062,I158884,I375282);
DFFARX1 I_9198 (I159062,I2683,I158717,I158706,);
DFFARX1 I_9199 (I159062,I2683,I158717,I158700,);
not I_9200 (I159107,I375282);
nor I_9201 (I159124,I159107,I375288);
and I_9202 (I159141,I159124,I375285);
or I_9203 (I159158,I159141,I375309);
DFFARX1 I_9204 (I159158,I2683,I158717,I159184,);
nand I_9205 (I159192,I159184,I158850);
nor I_9206 (I158694,I159192,I159000);
nor I_9207 (I158688,I159184,I158816);
DFFARX1 I_9208 (I159184,I2683,I158717,I159246,);
not I_9209 (I159254,I159246);
nor I_9210 (I158703,I159254,I158966);
not I_9211 (I159312,I2690);
DFFARX1 I_9212 (I994357,I2683,I159312,I159338,);
DFFARX1 I_9213 (I159338,I2683,I159312,I159355,);
not I_9214 (I159304,I159355);
not I_9215 (I159377,I159338);
DFFARX1 I_9216 (I994369,I2683,I159312,I159403,);
not I_9217 (I159411,I159403);
and I_9218 (I159428,I159377,I994363);
not I_9219 (I159445,I994375);
nand I_9220 (I159462,I159445,I994363);
not I_9221 (I159479,I994360);
nor I_9222 (I159496,I159479,I994372);
nand I_9223 (I159513,I159496,I994354);
nor I_9224 (I159530,I159513,I159462);
DFFARX1 I_9225 (I159530,I2683,I159312,I159280,);
not I_9226 (I159561,I159513);
not I_9227 (I159578,I994372);
nand I_9228 (I159595,I159578,I994363);
nor I_9229 (I159612,I994372,I994375);
nand I_9230 (I159292,I159428,I159612);
nand I_9231 (I159286,I159377,I994372);
nand I_9232 (I159657,I159479,I994366);
DFFARX1 I_9233 (I159657,I2683,I159312,I159301,);
DFFARX1 I_9234 (I159657,I2683,I159312,I159295,);
not I_9235 (I159702,I994366);
nor I_9236 (I159719,I159702,I994357);
and I_9237 (I159736,I159719,I994354);
or I_9238 (I159753,I159736,I994378);
DFFARX1 I_9239 (I159753,I2683,I159312,I159779,);
nand I_9240 (I159787,I159779,I159445);
nor I_9241 (I159289,I159787,I159595);
nor I_9242 (I159283,I159779,I159411);
DFFARX1 I_9243 (I159779,I2683,I159312,I159841,);
not I_9244 (I159849,I159841);
nor I_9245 (I159298,I159849,I159561);
not I_9246 (I159907,I2690);
DFFARX1 I_9247 (I1087620,I2683,I159907,I159933,);
DFFARX1 I_9248 (I159933,I2683,I159907,I159950,);
not I_9249 (I159899,I159950);
not I_9250 (I159972,I159933);
DFFARX1 I_9251 (I1087611,I2683,I159907,I159998,);
not I_9252 (I160006,I159998);
and I_9253 (I160023,I159972,I1087605);
not I_9254 (I160040,I1087599);
nand I_9255 (I160057,I160040,I1087605);
not I_9256 (I160074,I1087626);
nor I_9257 (I160091,I160074,I1087599);
nand I_9258 (I160108,I160091,I1087623);
nor I_9259 (I160125,I160108,I160057);
DFFARX1 I_9260 (I160125,I2683,I159907,I159875,);
not I_9261 (I160156,I160108);
not I_9262 (I160173,I1087599);
nand I_9263 (I160190,I160173,I1087605);
nor I_9264 (I160207,I1087599,I1087599);
nand I_9265 (I159887,I160023,I160207);
nand I_9266 (I159881,I159972,I1087599);
nand I_9267 (I160252,I160074,I1087608);
DFFARX1 I_9268 (I160252,I2683,I159907,I159896,);
DFFARX1 I_9269 (I160252,I2683,I159907,I159890,);
not I_9270 (I160297,I1087608);
nor I_9271 (I160314,I160297,I1087614);
and I_9272 (I160331,I160314,I1087617);
or I_9273 (I160348,I160331,I1087602);
DFFARX1 I_9274 (I160348,I2683,I159907,I160374,);
nand I_9275 (I160382,I160374,I160040);
nor I_9276 (I159884,I160382,I160190);
nor I_9277 (I159878,I160374,I160006);
DFFARX1 I_9278 (I160374,I2683,I159907,I160436,);
not I_9279 (I160444,I160436);
nor I_9280 (I159893,I160444,I160156);
not I_9281 (I160502,I2690);
DFFARX1 I_9282 (I90150,I2683,I160502,I160528,);
DFFARX1 I_9283 (I160528,I2683,I160502,I160545,);
not I_9284 (I160494,I160545);
not I_9285 (I160567,I160528);
DFFARX1 I_9286 (I90144,I2683,I160502,I160593,);
not I_9287 (I160601,I160593);
and I_9288 (I160618,I160567,I90141);
not I_9289 (I160635,I90162);
nand I_9290 (I160652,I160635,I90141);
not I_9291 (I160669,I90156);
nor I_9292 (I160686,I160669,I90147);
nand I_9293 (I160703,I160686,I90153);
nor I_9294 (I160720,I160703,I160652);
DFFARX1 I_9295 (I160720,I2683,I160502,I160470,);
not I_9296 (I160751,I160703);
not I_9297 (I160768,I90147);
nand I_9298 (I160785,I160768,I90141);
nor I_9299 (I160802,I90147,I90162);
nand I_9300 (I160482,I160618,I160802);
nand I_9301 (I160476,I160567,I90147);
nand I_9302 (I160847,I160669,I90141);
DFFARX1 I_9303 (I160847,I2683,I160502,I160491,);
DFFARX1 I_9304 (I160847,I2683,I160502,I160485,);
not I_9305 (I160892,I90141);
nor I_9306 (I160909,I160892,I90159);
and I_9307 (I160926,I160909,I90165);
or I_9308 (I160943,I160926,I90144);
DFFARX1 I_9309 (I160943,I2683,I160502,I160969,);
nand I_9310 (I160977,I160969,I160635);
nor I_9311 (I160479,I160977,I160785);
nor I_9312 (I160473,I160969,I160601);
DFFARX1 I_9313 (I160969,I2683,I160502,I161031,);
not I_9314 (I161039,I161031);
nor I_9315 (I160488,I161039,I160751);
not I_9316 (I161097,I2690);
DFFARX1 I_9317 (I465363,I2683,I161097,I161123,);
DFFARX1 I_9318 (I161123,I2683,I161097,I161140,);
not I_9319 (I161089,I161140);
not I_9320 (I161162,I161123);
DFFARX1 I_9321 (I465354,I2683,I161097,I161188,);
not I_9322 (I161196,I161188);
and I_9323 (I161213,I161162,I465372);
not I_9324 (I161230,I465369);
nand I_9325 (I161247,I161230,I465372);
not I_9326 (I161264,I465348);
nor I_9327 (I161281,I161264,I465351);
nand I_9328 (I161298,I161281,I465360);
nor I_9329 (I161315,I161298,I161247);
DFFARX1 I_9330 (I161315,I2683,I161097,I161065,);
not I_9331 (I161346,I161298);
not I_9332 (I161363,I465351);
nand I_9333 (I161380,I161363,I465372);
nor I_9334 (I161397,I465351,I465369);
nand I_9335 (I161077,I161213,I161397);
nand I_9336 (I161071,I161162,I465351);
nand I_9337 (I161442,I161264,I465366);
DFFARX1 I_9338 (I161442,I2683,I161097,I161086,);
DFFARX1 I_9339 (I161442,I2683,I161097,I161080,);
not I_9340 (I161487,I465366);
nor I_9341 (I161504,I161487,I465348);
and I_9342 (I161521,I161504,I465357);
or I_9343 (I161538,I161521,I465351);
DFFARX1 I_9344 (I161538,I2683,I161097,I161564,);
nand I_9345 (I161572,I161564,I161230);
nor I_9346 (I161074,I161572,I161380);
nor I_9347 (I161068,I161564,I161196);
DFFARX1 I_9348 (I161564,I2683,I161097,I161626,);
not I_9349 (I161634,I161626);
nor I_9350 (I161083,I161634,I161346);
not I_9351 (I161692,I2690);
DFFARX1 I_9352 (I698152,I2683,I161692,I161718,);
DFFARX1 I_9353 (I161718,I2683,I161692,I161735,);
not I_9354 (I161684,I161735);
not I_9355 (I161757,I161718);
DFFARX1 I_9356 (I698146,I2683,I161692,I161783,);
not I_9357 (I161791,I161783);
and I_9358 (I161808,I161757,I698164);
not I_9359 (I161825,I698152);
nand I_9360 (I161842,I161825,I698164);
not I_9361 (I161859,I698146);
nor I_9362 (I161876,I161859,I698158);
nand I_9363 (I161893,I161876,I698149);
nor I_9364 (I161910,I161893,I161842);
DFFARX1 I_9365 (I161910,I2683,I161692,I161660,);
not I_9366 (I161941,I161893);
not I_9367 (I161958,I698158);
nand I_9368 (I161975,I161958,I698164);
nor I_9369 (I161992,I698158,I698152);
nand I_9370 (I161672,I161808,I161992);
nand I_9371 (I161666,I161757,I698158);
nand I_9372 (I162037,I161859,I698161);
DFFARX1 I_9373 (I162037,I2683,I161692,I161681,);
DFFARX1 I_9374 (I162037,I2683,I161692,I161675,);
not I_9375 (I162082,I698161);
nor I_9376 (I162099,I162082,I698167);
and I_9377 (I162116,I162099,I698149);
or I_9378 (I162133,I162116,I698155);
DFFARX1 I_9379 (I162133,I2683,I161692,I162159,);
nand I_9380 (I162167,I162159,I161825);
nor I_9381 (I161669,I162167,I161975);
nor I_9382 (I161663,I162159,I161791);
DFFARX1 I_9383 (I162159,I2683,I161692,I162221,);
not I_9384 (I162229,I162221);
nor I_9385 (I161678,I162229,I161941);
not I_9386 (I162287,I2690);
DFFARX1 I_9387 (I931658,I2683,I162287,I162313,);
DFFARX1 I_9388 (I162313,I2683,I162287,I162330,);
not I_9389 (I162279,I162330);
not I_9390 (I162352,I162313);
DFFARX1 I_9391 (I931658,I2683,I162287,I162378,);
not I_9392 (I162386,I162378);
and I_9393 (I162403,I162352,I931661);
not I_9394 (I162420,I931673);
nand I_9395 (I162437,I162420,I931661);
not I_9396 (I162454,I931679);
nor I_9397 (I162471,I162454,I931670);
nand I_9398 (I162488,I162471,I931676);
nor I_9399 (I162505,I162488,I162437);
DFFARX1 I_9400 (I162505,I2683,I162287,I162255,);
not I_9401 (I162536,I162488);
not I_9402 (I162553,I931670);
nand I_9403 (I162570,I162553,I931661);
nor I_9404 (I162587,I931670,I931673);
nand I_9405 (I162267,I162403,I162587);
nand I_9406 (I162261,I162352,I931670);
nand I_9407 (I162632,I162454,I931667);
DFFARX1 I_9408 (I162632,I2683,I162287,I162276,);
DFFARX1 I_9409 (I162632,I2683,I162287,I162270,);
not I_9410 (I162677,I931667);
nor I_9411 (I162694,I162677,I931664);
and I_9412 (I162711,I162694,I931682);
or I_9413 (I162728,I162711,I931661);
DFFARX1 I_9414 (I162728,I2683,I162287,I162754,);
nand I_9415 (I162762,I162754,I162420);
nor I_9416 (I162264,I162762,I162570);
nor I_9417 (I162258,I162754,I162386);
DFFARX1 I_9418 (I162754,I2683,I162287,I162816,);
not I_9419 (I162824,I162816);
nor I_9420 (I162273,I162824,I162536);
not I_9421 (I162882,I2690);
DFFARX1 I_9422 (I925300,I2683,I162882,I162908,);
DFFARX1 I_9423 (I162908,I2683,I162882,I162925,);
not I_9424 (I162874,I162925);
not I_9425 (I162947,I162908);
DFFARX1 I_9426 (I925300,I2683,I162882,I162973,);
not I_9427 (I162981,I162973);
and I_9428 (I162998,I162947,I925303);
not I_9429 (I163015,I925315);
nand I_9430 (I163032,I163015,I925303);
not I_9431 (I163049,I925321);
nor I_9432 (I163066,I163049,I925312);
nand I_9433 (I163083,I163066,I925318);
nor I_9434 (I163100,I163083,I163032);
DFFARX1 I_9435 (I163100,I2683,I162882,I162850,);
not I_9436 (I163131,I163083);
not I_9437 (I163148,I925312);
nand I_9438 (I163165,I163148,I925303);
nor I_9439 (I163182,I925312,I925315);
nand I_9440 (I162862,I162998,I163182);
nand I_9441 (I162856,I162947,I925312);
nand I_9442 (I163227,I163049,I925309);
DFFARX1 I_9443 (I163227,I2683,I162882,I162871,);
DFFARX1 I_9444 (I163227,I2683,I162882,I162865,);
not I_9445 (I163272,I925309);
nor I_9446 (I163289,I163272,I925306);
and I_9447 (I163306,I163289,I925324);
or I_9448 (I163323,I163306,I925303);
DFFARX1 I_9449 (I163323,I2683,I162882,I163349,);
nand I_9450 (I163357,I163349,I163015);
nor I_9451 (I162859,I163357,I163165);
nor I_9452 (I162853,I163349,I162981);
DFFARX1 I_9453 (I163349,I2683,I162882,I163411,);
not I_9454 (I163419,I163411);
nor I_9455 (I162868,I163419,I163131);
not I_9456 (I163477,I2690);
DFFARX1 I_9457 (I294906,I2683,I163477,I163503,);
DFFARX1 I_9458 (I163503,I2683,I163477,I163520,);
not I_9459 (I163469,I163520);
not I_9460 (I163542,I163503);
DFFARX1 I_9461 (I294921,I2683,I163477,I163568,);
not I_9462 (I163576,I163568);
and I_9463 (I163593,I163542,I294918);
not I_9464 (I163610,I294906);
nand I_9465 (I163627,I163610,I294918);
not I_9466 (I163644,I294915);
nor I_9467 (I163661,I163644,I294930);
nand I_9468 (I163678,I163661,I294927);
nor I_9469 (I163695,I163678,I163627);
DFFARX1 I_9470 (I163695,I2683,I163477,I163445,);
not I_9471 (I163726,I163678);
not I_9472 (I163743,I294930);
nand I_9473 (I163760,I163743,I294918);
nor I_9474 (I163777,I294930,I294906);
nand I_9475 (I163457,I163593,I163777);
nand I_9476 (I163451,I163542,I294930);
nand I_9477 (I163822,I163644,I294924);
DFFARX1 I_9478 (I163822,I2683,I163477,I163466,);
DFFARX1 I_9479 (I163822,I2683,I163477,I163460,);
not I_9480 (I163867,I294924);
nor I_9481 (I163884,I163867,I294912);
and I_9482 (I163901,I163884,I294933);
or I_9483 (I163918,I163901,I294909);
DFFARX1 I_9484 (I163918,I2683,I163477,I163944,);
nand I_9485 (I163952,I163944,I163610);
nor I_9486 (I163454,I163952,I163760);
nor I_9487 (I163448,I163944,I163576);
DFFARX1 I_9488 (I163944,I2683,I163477,I164006,);
not I_9489 (I164014,I164006);
nor I_9490 (I163463,I164014,I163726);
not I_9491 (I164072,I2690);
DFFARX1 I_9492 (I975536,I2683,I164072,I164098,);
DFFARX1 I_9493 (I164098,I2683,I164072,I164115,);
not I_9494 (I164064,I164115);
not I_9495 (I164137,I164098);
DFFARX1 I_9496 (I975521,I2683,I164072,I164163,);
not I_9497 (I164171,I164163);
and I_9498 (I164188,I164137,I975539);
not I_9499 (I164205,I975521);
nand I_9500 (I164222,I164205,I975539);
not I_9501 (I164239,I975542);
nor I_9502 (I164256,I164239,I975533);
nand I_9503 (I164273,I164256,I975530);
nor I_9504 (I164290,I164273,I164222);
DFFARX1 I_9505 (I164290,I2683,I164072,I164040,);
not I_9506 (I164321,I164273);
not I_9507 (I164338,I975533);
nand I_9508 (I164355,I164338,I975539);
nor I_9509 (I164372,I975533,I975521);
nand I_9510 (I164052,I164188,I164372);
nand I_9511 (I164046,I164137,I975533);
nand I_9512 (I164417,I164239,I975527);
DFFARX1 I_9513 (I164417,I2683,I164072,I164061,);
DFFARX1 I_9514 (I164417,I2683,I164072,I164055,);
not I_9515 (I164462,I975527);
nor I_9516 (I164479,I164462,I975518);
and I_9517 (I164496,I164479,I975524);
or I_9518 (I164513,I164496,I975518);
DFFARX1 I_9519 (I164513,I2683,I164072,I164539,);
nand I_9520 (I164547,I164539,I164205);
nor I_9521 (I164049,I164547,I164355);
nor I_9522 (I164043,I164539,I164171);
DFFARX1 I_9523 (I164539,I2683,I164072,I164601,);
not I_9524 (I164609,I164601);
nor I_9525 (I164058,I164609,I164321);
not I_9526 (I164667,I2690);
DFFARX1 I_9527 (I526628,I2683,I164667,I164693,);
DFFARX1 I_9528 (I164693,I2683,I164667,I164710,);
not I_9529 (I164659,I164710);
not I_9530 (I164732,I164693);
DFFARX1 I_9531 (I526625,I2683,I164667,I164758,);
not I_9532 (I164766,I164758);
and I_9533 (I164783,I164732,I526631);
not I_9534 (I164800,I526616);
nand I_9535 (I164817,I164800,I526631);
not I_9536 (I164834,I526619);
nor I_9537 (I164851,I164834,I526640);
nand I_9538 (I164868,I164851,I526637);
nor I_9539 (I164885,I164868,I164817);
DFFARX1 I_9540 (I164885,I2683,I164667,I164635,);
not I_9541 (I164916,I164868);
not I_9542 (I164933,I526640);
nand I_9543 (I164950,I164933,I526631);
nor I_9544 (I164967,I526640,I526616);
nand I_9545 (I164647,I164783,I164967);
nand I_9546 (I164641,I164732,I526640);
nand I_9547 (I165012,I164834,I526616);
DFFARX1 I_9548 (I165012,I2683,I164667,I164656,);
DFFARX1 I_9549 (I165012,I2683,I164667,I164650,);
not I_9550 (I165057,I526616);
nor I_9551 (I165074,I165057,I526622);
and I_9552 (I165091,I165074,I526634);
or I_9553 (I165108,I165091,I526619);
DFFARX1 I_9554 (I165108,I2683,I164667,I165134,);
nand I_9555 (I165142,I165134,I164800);
nor I_9556 (I164644,I165142,I164950);
nor I_9557 (I164638,I165134,I164766);
DFFARX1 I_9558 (I165134,I2683,I164667,I165196,);
not I_9559 (I165204,I165196);
nor I_9560 (I164653,I165204,I164916);
not I_9561 (I165262,I2690);
DFFARX1 I_9562 (I29560,I2683,I165262,I165288,);
DFFARX1 I_9563 (I165288,I2683,I165262,I165305,);
not I_9564 (I165254,I165305);
not I_9565 (I165327,I165288);
DFFARX1 I_9566 (I29536,I2683,I165262,I165353,);
not I_9567 (I165361,I165353);
and I_9568 (I165378,I165327,I29551);
not I_9569 (I165395,I29539);
nand I_9570 (I165412,I165395,I29551);
not I_9571 (I165429,I29542);
nor I_9572 (I165446,I165429,I29554);
nand I_9573 (I165463,I165446,I29545);
nor I_9574 (I165480,I165463,I165412);
DFFARX1 I_9575 (I165480,I2683,I165262,I165230,);
not I_9576 (I165511,I165463);
not I_9577 (I165528,I29554);
nand I_9578 (I165545,I165528,I29551);
nor I_9579 (I165562,I29554,I29539);
nand I_9580 (I165242,I165378,I165562);
nand I_9581 (I165236,I165327,I29554);
nand I_9582 (I165607,I165429,I29548);
DFFARX1 I_9583 (I165607,I2683,I165262,I165251,);
DFFARX1 I_9584 (I165607,I2683,I165262,I165245,);
not I_9585 (I165652,I29548);
nor I_9586 (I165669,I165652,I29539);
and I_9587 (I165686,I165669,I29536);
or I_9588 (I165703,I165686,I29557);
DFFARX1 I_9589 (I165703,I2683,I165262,I165729,);
nand I_9590 (I165737,I165729,I165395);
nor I_9591 (I165239,I165737,I165545);
nor I_9592 (I165233,I165729,I165361);
DFFARX1 I_9593 (I165729,I2683,I165262,I165791,);
not I_9594 (I165799,I165791);
nor I_9595 (I165248,I165799,I165511);
not I_9596 (I165857,I2690);
DFFARX1 I_9597 (I881950,I2683,I165857,I165883,);
DFFARX1 I_9598 (I165883,I2683,I165857,I165900,);
not I_9599 (I165849,I165900);
not I_9600 (I165922,I165883);
DFFARX1 I_9601 (I881950,I2683,I165857,I165948,);
not I_9602 (I165956,I165948);
and I_9603 (I165973,I165922,I881953);
not I_9604 (I165990,I881965);
nand I_9605 (I166007,I165990,I881953);
not I_9606 (I166024,I881971);
nor I_9607 (I166041,I166024,I881962);
nand I_9608 (I166058,I166041,I881968);
nor I_9609 (I166075,I166058,I166007);
DFFARX1 I_9610 (I166075,I2683,I165857,I165825,);
not I_9611 (I166106,I166058);
not I_9612 (I166123,I881962);
nand I_9613 (I166140,I166123,I881953);
nor I_9614 (I166157,I881962,I881965);
nand I_9615 (I165837,I165973,I166157);
nand I_9616 (I165831,I165922,I881962);
nand I_9617 (I166202,I166024,I881959);
DFFARX1 I_9618 (I166202,I2683,I165857,I165846,);
DFFARX1 I_9619 (I166202,I2683,I165857,I165840,);
not I_9620 (I166247,I881959);
nor I_9621 (I166264,I166247,I881956);
and I_9622 (I166281,I166264,I881974);
or I_9623 (I166298,I166281,I881953);
DFFARX1 I_9624 (I166298,I2683,I165857,I166324,);
nand I_9625 (I166332,I166324,I165990);
nor I_9626 (I165834,I166332,I166140);
nor I_9627 (I165828,I166324,I165956);
DFFARX1 I_9628 (I166324,I2683,I165857,I166386,);
not I_9629 (I166394,I166386);
nor I_9630 (I165843,I166394,I166106);
not I_9631 (I166452,I2690);
DFFARX1 I_9632 (I280677,I2683,I166452,I166478,);
DFFARX1 I_9633 (I166478,I2683,I166452,I166495,);
not I_9634 (I166444,I166495);
not I_9635 (I166517,I166478);
DFFARX1 I_9636 (I280692,I2683,I166452,I166543,);
not I_9637 (I166551,I166543);
and I_9638 (I166568,I166517,I280689);
not I_9639 (I166585,I280677);
nand I_9640 (I166602,I166585,I280689);
not I_9641 (I166619,I280686);
nor I_9642 (I166636,I166619,I280701);
nand I_9643 (I166653,I166636,I280698);
nor I_9644 (I166670,I166653,I166602);
DFFARX1 I_9645 (I166670,I2683,I166452,I166420,);
not I_9646 (I166701,I166653);
not I_9647 (I166718,I280701);
nand I_9648 (I166735,I166718,I280689);
nor I_9649 (I166752,I280701,I280677);
nand I_9650 (I166432,I166568,I166752);
nand I_9651 (I166426,I166517,I280701);
nand I_9652 (I166797,I166619,I280695);
DFFARX1 I_9653 (I166797,I2683,I166452,I166441,);
DFFARX1 I_9654 (I166797,I2683,I166452,I166435,);
not I_9655 (I166842,I280695);
nor I_9656 (I166859,I166842,I280683);
and I_9657 (I166876,I166859,I280704);
or I_9658 (I166893,I166876,I280680);
DFFARX1 I_9659 (I166893,I2683,I166452,I166919,);
nand I_9660 (I166927,I166919,I166585);
nor I_9661 (I166429,I166927,I166735);
nor I_9662 (I166423,I166919,I166551);
DFFARX1 I_9663 (I166919,I2683,I166452,I166981,);
not I_9664 (I166989,I166981);
nor I_9665 (I166438,I166989,I166701);
not I_9666 (I167047,I2690);
DFFARX1 I_9667 (I611016,I2683,I167047,I167073,);
DFFARX1 I_9668 (I167073,I2683,I167047,I167090,);
not I_9669 (I167039,I167090);
not I_9670 (I167112,I167073);
DFFARX1 I_9671 (I611013,I2683,I167047,I167138,);
not I_9672 (I167146,I167138);
and I_9673 (I167163,I167112,I611019);
not I_9674 (I167180,I611004);
nand I_9675 (I167197,I167180,I611019);
not I_9676 (I167214,I611007);
nor I_9677 (I167231,I167214,I611028);
nand I_9678 (I167248,I167231,I611025);
nor I_9679 (I167265,I167248,I167197);
DFFARX1 I_9680 (I167265,I2683,I167047,I167015,);
not I_9681 (I167296,I167248);
not I_9682 (I167313,I611028);
nand I_9683 (I167330,I167313,I611019);
nor I_9684 (I167347,I611028,I611004);
nand I_9685 (I167027,I167163,I167347);
nand I_9686 (I167021,I167112,I611028);
nand I_9687 (I167392,I167214,I611004);
DFFARX1 I_9688 (I167392,I2683,I167047,I167036,);
DFFARX1 I_9689 (I167392,I2683,I167047,I167030,);
not I_9690 (I167437,I611004);
nor I_9691 (I167454,I167437,I611010);
and I_9692 (I167471,I167454,I611022);
or I_9693 (I167488,I167471,I611007);
DFFARX1 I_9694 (I167488,I2683,I167047,I167514,);
nand I_9695 (I167522,I167514,I167180);
nor I_9696 (I167024,I167522,I167330);
nor I_9697 (I167018,I167514,I167146);
DFFARX1 I_9698 (I167514,I2683,I167047,I167576,);
not I_9699 (I167584,I167576);
nor I_9700 (I167033,I167584,I167296);
not I_9701 (I167642,I2690);
DFFARX1 I_9702 (I269083,I2683,I167642,I167668,);
DFFARX1 I_9703 (I167668,I2683,I167642,I167685,);
not I_9704 (I167634,I167685);
not I_9705 (I167707,I167668);
DFFARX1 I_9706 (I269098,I2683,I167642,I167733,);
not I_9707 (I167741,I167733);
and I_9708 (I167758,I167707,I269095);
not I_9709 (I167775,I269083);
nand I_9710 (I167792,I167775,I269095);
not I_9711 (I167809,I269092);
nor I_9712 (I167826,I167809,I269107);
nand I_9713 (I167843,I167826,I269104);
nor I_9714 (I167860,I167843,I167792);
DFFARX1 I_9715 (I167860,I2683,I167642,I167610,);
not I_9716 (I167891,I167843);
not I_9717 (I167908,I269107);
nand I_9718 (I167925,I167908,I269095);
nor I_9719 (I167942,I269107,I269083);
nand I_9720 (I167622,I167758,I167942);
nand I_9721 (I167616,I167707,I269107);
nand I_9722 (I167987,I167809,I269101);
DFFARX1 I_9723 (I167987,I2683,I167642,I167631,);
DFFARX1 I_9724 (I167987,I2683,I167642,I167625,);
not I_9725 (I168032,I269101);
nor I_9726 (I168049,I168032,I269089);
and I_9727 (I168066,I168049,I269110);
or I_9728 (I168083,I168066,I269086);
DFFARX1 I_9729 (I168083,I2683,I167642,I168109,);
nand I_9730 (I168117,I168109,I167775);
nor I_9731 (I167619,I168117,I167925);
nor I_9732 (I167613,I168109,I167741);
DFFARX1 I_9733 (I168109,I2683,I167642,I168171,);
not I_9734 (I168179,I168171);
nor I_9735 (I167628,I168179,I167891);
not I_9736 (I168237,I2690);
DFFARX1 I_9737 (I957040,I2683,I168237,I168263,);
DFFARX1 I_9738 (I168263,I2683,I168237,I168280,);
not I_9739 (I168229,I168280);
not I_9740 (I168302,I168263);
DFFARX1 I_9741 (I957025,I2683,I168237,I168328,);
not I_9742 (I168336,I168328);
and I_9743 (I168353,I168302,I957043);
not I_9744 (I168370,I957025);
nand I_9745 (I168387,I168370,I957043);
not I_9746 (I168404,I957046);
nor I_9747 (I168421,I168404,I957037);
nand I_9748 (I168438,I168421,I957034);
nor I_9749 (I168455,I168438,I168387);
DFFARX1 I_9750 (I168455,I2683,I168237,I168205,);
not I_9751 (I168486,I168438);
not I_9752 (I168503,I957037);
nand I_9753 (I168520,I168503,I957043);
nor I_9754 (I168537,I957037,I957025);
nand I_9755 (I168217,I168353,I168537);
nand I_9756 (I168211,I168302,I957037);
nand I_9757 (I168582,I168404,I957031);
DFFARX1 I_9758 (I168582,I2683,I168237,I168226,);
DFFARX1 I_9759 (I168582,I2683,I168237,I168220,);
not I_9760 (I168627,I957031);
nor I_9761 (I168644,I168627,I957022);
and I_9762 (I168661,I168644,I957028);
or I_9763 (I168678,I168661,I957022);
DFFARX1 I_9764 (I168678,I2683,I168237,I168704,);
nand I_9765 (I168712,I168704,I168370);
nor I_9766 (I168214,I168712,I168520);
nor I_9767 (I168208,I168704,I168336);
DFFARX1 I_9768 (I168704,I2683,I168237,I168766,);
not I_9769 (I168774,I168766);
nor I_9770 (I168223,I168774,I168486);
not I_9771 (I168832,I2690);
DFFARX1 I_9772 (I347018,I2683,I168832,I168858,);
DFFARX1 I_9773 (I168858,I2683,I168832,I168875,);
not I_9774 (I168824,I168875);
not I_9775 (I168897,I168858);
DFFARX1 I_9776 (I347006,I2683,I168832,I168923,);
not I_9777 (I168931,I168923);
and I_9778 (I168948,I168897,I347015);
not I_9779 (I168965,I347012);
nand I_9780 (I168982,I168965,I347015);
not I_9781 (I168999,I347003);
nor I_9782 (I169016,I168999,I347009);
nand I_9783 (I169033,I169016,I346994);
nor I_9784 (I169050,I169033,I168982);
DFFARX1 I_9785 (I169050,I2683,I168832,I168800,);
not I_9786 (I169081,I169033);
not I_9787 (I169098,I347009);
nand I_9788 (I169115,I169098,I347015);
nor I_9789 (I169132,I347009,I347012);
nand I_9790 (I168812,I168948,I169132);
nand I_9791 (I168806,I168897,I347009);
nand I_9792 (I169177,I168999,I346994);
DFFARX1 I_9793 (I169177,I2683,I168832,I168821,);
DFFARX1 I_9794 (I169177,I2683,I168832,I168815,);
not I_9795 (I169222,I346994);
nor I_9796 (I169239,I169222,I347000);
and I_9797 (I169256,I169239,I346997);
or I_9798 (I169273,I169256,I347021);
DFFARX1 I_9799 (I169273,I2683,I168832,I169299,);
nand I_9800 (I169307,I169299,I168965);
nor I_9801 (I168809,I169307,I169115);
nor I_9802 (I168803,I169299,I168931);
DFFARX1 I_9803 (I169299,I2683,I168832,I169361,);
not I_9804 (I169369,I169361);
nor I_9805 (I168818,I169369,I169081);
not I_9806 (I169427,I2690);
DFFARX1 I_9807 (I632277,I2683,I169427,I169453,);
DFFARX1 I_9808 (I169453,I2683,I169427,I169470,);
not I_9809 (I169419,I169470);
not I_9810 (I169492,I169453);
DFFARX1 I_9811 (I632271,I2683,I169427,I169518,);
not I_9812 (I169526,I169518);
and I_9813 (I169543,I169492,I632289);
not I_9814 (I169560,I632277);
nand I_9815 (I169577,I169560,I632289);
not I_9816 (I169594,I632271);
nor I_9817 (I169611,I169594,I632283);
nand I_9818 (I169628,I169611,I632274);
nor I_9819 (I169645,I169628,I169577);
DFFARX1 I_9820 (I169645,I2683,I169427,I169395,);
not I_9821 (I169676,I169628);
not I_9822 (I169693,I632283);
nand I_9823 (I169710,I169693,I632289);
nor I_9824 (I169727,I632283,I632277);
nand I_9825 (I169407,I169543,I169727);
nand I_9826 (I169401,I169492,I632283);
nand I_9827 (I169772,I169594,I632286);
DFFARX1 I_9828 (I169772,I2683,I169427,I169416,);
DFFARX1 I_9829 (I169772,I2683,I169427,I169410,);
not I_9830 (I169817,I632286);
nor I_9831 (I169834,I169817,I632292);
and I_9832 (I169851,I169834,I632274);
or I_9833 (I169868,I169851,I632280);
DFFARX1 I_9834 (I169868,I2683,I169427,I169894,);
nand I_9835 (I169902,I169894,I169560);
nor I_9836 (I169404,I169902,I169710);
nor I_9837 (I169398,I169894,I169526);
DFFARX1 I_9838 (I169894,I2683,I169427,I169956,);
not I_9839 (I169964,I169956);
nor I_9840 (I169413,I169964,I169676);
not I_9841 (I170022,I2690);
DFFARX1 I_9842 (I615062,I2683,I170022,I170048,);
DFFARX1 I_9843 (I170048,I2683,I170022,I170065,);
not I_9844 (I170014,I170065);
not I_9845 (I170087,I170048);
DFFARX1 I_9846 (I615059,I2683,I170022,I170113,);
not I_9847 (I170121,I170113);
and I_9848 (I170138,I170087,I615065);
not I_9849 (I170155,I615050);
nand I_9850 (I170172,I170155,I615065);
not I_9851 (I170189,I615053);
nor I_9852 (I170206,I170189,I615074);
nand I_9853 (I170223,I170206,I615071);
nor I_9854 (I170240,I170223,I170172);
DFFARX1 I_9855 (I170240,I2683,I170022,I169990,);
not I_9856 (I170271,I170223);
not I_9857 (I170288,I615074);
nand I_9858 (I170305,I170288,I615065);
nor I_9859 (I170322,I615074,I615050);
nand I_9860 (I170002,I170138,I170322);
nand I_9861 (I169996,I170087,I615074);
nand I_9862 (I170367,I170189,I615050);
DFFARX1 I_9863 (I170367,I2683,I170022,I170011,);
DFFARX1 I_9864 (I170367,I2683,I170022,I170005,);
not I_9865 (I170412,I615050);
nor I_9866 (I170429,I170412,I615056);
and I_9867 (I170446,I170429,I615068);
or I_9868 (I170463,I170446,I615053);
DFFARX1 I_9869 (I170463,I2683,I170022,I170489,);
nand I_9870 (I170497,I170489,I170155);
nor I_9871 (I169999,I170497,I170305);
nor I_9872 (I169993,I170489,I170121);
DFFARX1 I_9873 (I170489,I2683,I170022,I170551,);
not I_9874 (I170559,I170551);
nor I_9875 (I170008,I170559,I170271);
not I_9876 (I170617,I2690);
DFFARX1 I_9877 (I47990,I2683,I170617,I170643,);
DFFARX1 I_9878 (I170643,I2683,I170617,I170660,);
not I_9879 (I170609,I170660);
not I_9880 (I170682,I170643);
DFFARX1 I_9881 (I47984,I2683,I170617,I170708,);
not I_9882 (I170716,I170708);
and I_9883 (I170733,I170682,I47981);
not I_9884 (I170750,I48002);
nand I_9885 (I170767,I170750,I47981);
not I_9886 (I170784,I47996);
nor I_9887 (I170801,I170784,I47987);
nand I_9888 (I170818,I170801,I47993);
nor I_9889 (I170835,I170818,I170767);
DFFARX1 I_9890 (I170835,I2683,I170617,I170585,);
not I_9891 (I170866,I170818);
not I_9892 (I170883,I47987);
nand I_9893 (I170900,I170883,I47981);
nor I_9894 (I170917,I47987,I48002);
nand I_9895 (I170597,I170733,I170917);
nand I_9896 (I170591,I170682,I47987);
nand I_9897 (I170962,I170784,I47981);
DFFARX1 I_9898 (I170962,I2683,I170617,I170606,);
DFFARX1 I_9899 (I170962,I2683,I170617,I170600,);
not I_9900 (I171007,I47981);
nor I_9901 (I171024,I171007,I47999);
and I_9902 (I171041,I171024,I48005);
or I_9903 (I171058,I171041,I47984);
DFFARX1 I_9904 (I171058,I2683,I170617,I171084,);
nand I_9905 (I171092,I171084,I170750);
nor I_9906 (I170594,I171092,I170900);
nor I_9907 (I170588,I171084,I170716);
DFFARX1 I_9908 (I171084,I2683,I170617,I171146,);
not I_9909 (I171154,I171146);
nor I_9910 (I170603,I171154,I170866);
not I_9911 (I171212,I2690);
DFFARX1 I_9912 (I1812,I2683,I171212,I171238,);
DFFARX1 I_9913 (I171238,I2683,I171212,I171255,);
not I_9914 (I171204,I171255);
not I_9915 (I171277,I171238);
DFFARX1 I_9916 (I2372,I2683,I171212,I171303,);
not I_9917 (I171311,I171303);
and I_9918 (I171328,I171277,I2668);
not I_9919 (I171345,I2020);
nand I_9920 (I171362,I171345,I2668);
not I_9921 (I171379,I1772);
nor I_9922 (I171396,I171379,I2028);
nand I_9923 (I171413,I171396,I1876);
nor I_9924 (I171430,I171413,I171362);
DFFARX1 I_9925 (I171430,I2683,I171212,I171180,);
not I_9926 (I171461,I171413);
not I_9927 (I171478,I2028);
nand I_9928 (I171495,I171478,I2668);
nor I_9929 (I171512,I2028,I2020);
nand I_9930 (I171192,I171328,I171512);
nand I_9931 (I171186,I171277,I2028);
nand I_9932 (I171557,I171379,I1668);
DFFARX1 I_9933 (I171557,I2683,I171212,I171201,);
DFFARX1 I_9934 (I171557,I2683,I171212,I171195,);
not I_9935 (I171602,I1668);
nor I_9936 (I171619,I171602,I2196);
and I_9937 (I171636,I171619,I1756);
or I_9938 (I171653,I171636,I1980);
DFFARX1 I_9939 (I171653,I2683,I171212,I171679,);
nand I_9940 (I171687,I171679,I171345);
nor I_9941 (I171189,I171687,I171495);
nor I_9942 (I171183,I171679,I171311);
DFFARX1 I_9943 (I171679,I2683,I171212,I171741,);
not I_9944 (I171749,I171741);
nor I_9945 (I171198,I171749,I171461);
not I_9946 (I171807,I2690);
DFFARX1 I_9947 (I485015,I2683,I171807,I171833,);
DFFARX1 I_9948 (I171833,I2683,I171807,I171850,);
not I_9949 (I171799,I171850);
not I_9950 (I171872,I171833);
DFFARX1 I_9951 (I485006,I2683,I171807,I171898,);
not I_9952 (I171906,I171898);
and I_9953 (I171923,I171872,I485024);
not I_9954 (I171940,I485021);
nand I_9955 (I171957,I171940,I485024);
not I_9956 (I171974,I485000);
nor I_9957 (I171991,I171974,I485003);
nand I_9958 (I172008,I171991,I485012);
nor I_9959 (I172025,I172008,I171957);
DFFARX1 I_9960 (I172025,I2683,I171807,I171775,);
not I_9961 (I172056,I172008);
not I_9962 (I172073,I485003);
nand I_9963 (I172090,I172073,I485024);
nor I_9964 (I172107,I485003,I485021);
nand I_9965 (I171787,I171923,I172107);
nand I_9966 (I171781,I171872,I485003);
nand I_9967 (I172152,I171974,I485018);
DFFARX1 I_9968 (I172152,I2683,I171807,I171796,);
DFFARX1 I_9969 (I172152,I2683,I171807,I171790,);
not I_9970 (I172197,I485018);
nor I_9971 (I172214,I172197,I485000);
and I_9972 (I172231,I172214,I485009);
or I_9973 (I172248,I172231,I485003);
DFFARX1 I_9974 (I172248,I2683,I171807,I172274,);
nand I_9975 (I172282,I172274,I171940);
nor I_9976 (I171784,I172282,I172090);
nor I_9977 (I171778,I172274,I171906);
DFFARX1 I_9978 (I172274,I2683,I171807,I172336,);
not I_9979 (I172344,I172336);
nor I_9980 (I171793,I172344,I172056);
not I_9981 (I172402,I2690);
DFFARX1 I_9982 (I652303,I2683,I172402,I172428,);
DFFARX1 I_9983 (I172428,I2683,I172402,I172445,);
not I_9984 (I172394,I172445);
not I_9985 (I172467,I172428);
DFFARX1 I_9986 (I652297,I2683,I172402,I172493,);
not I_9987 (I172501,I172493);
and I_9988 (I172518,I172467,I652315);
not I_9989 (I172535,I652303);
nand I_9990 (I172552,I172535,I652315);
not I_9991 (I172569,I652297);
nor I_9992 (I172586,I172569,I652309);
nand I_9993 (I172603,I172586,I652300);
nor I_9994 (I172620,I172603,I172552);
DFFARX1 I_9995 (I172620,I2683,I172402,I172370,);
not I_9996 (I172651,I172603);
not I_9997 (I172668,I652309);
nand I_9998 (I172685,I172668,I652315);
nor I_9999 (I172702,I652309,I652303);
nand I_10000 (I172382,I172518,I172702);
nand I_10001 (I172376,I172467,I652309);
nand I_10002 (I172747,I172569,I652312);
DFFARX1 I_10003 (I172747,I2683,I172402,I172391,);
DFFARX1 I_10004 (I172747,I2683,I172402,I172385,);
not I_10005 (I172792,I652312);
nor I_10006 (I172809,I172792,I652318);
and I_10007 (I172826,I172809,I652300);
or I_10008 (I172843,I172826,I652306);
DFFARX1 I_10009 (I172843,I2683,I172402,I172869,);
nand I_10010 (I172877,I172869,I172535);
nor I_10011 (I172379,I172877,I172685);
nor I_10012 (I172373,I172869,I172501);
DFFARX1 I_10013 (I172869,I2683,I172402,I172931,);
not I_10014 (I172939,I172931);
nor I_10015 (I172388,I172939,I172651);
not I_10016 (I172997,I2690);
DFFARX1 I_10017 (I69597,I2683,I172997,I173023,);
DFFARX1 I_10018 (I173023,I2683,I172997,I173040,);
not I_10019 (I172989,I173040);
not I_10020 (I173062,I173023);
DFFARX1 I_10021 (I69591,I2683,I172997,I173088,);
not I_10022 (I173096,I173088);
and I_10023 (I173113,I173062,I69588);
not I_10024 (I173130,I69609);
nand I_10025 (I173147,I173130,I69588);
not I_10026 (I173164,I69603);
nor I_10027 (I173181,I173164,I69594);
nand I_10028 (I173198,I173181,I69600);
nor I_10029 (I173215,I173198,I173147);
DFFARX1 I_10030 (I173215,I2683,I172997,I172965,);
not I_10031 (I173246,I173198);
not I_10032 (I173263,I69594);
nand I_10033 (I173280,I173263,I69588);
nor I_10034 (I173297,I69594,I69609);
nand I_10035 (I172977,I173113,I173297);
nand I_10036 (I172971,I173062,I69594);
nand I_10037 (I173342,I173164,I69588);
DFFARX1 I_10038 (I173342,I2683,I172997,I172986,);
DFFARX1 I_10039 (I173342,I2683,I172997,I172980,);
not I_10040 (I173387,I69588);
nor I_10041 (I173404,I173387,I69606);
and I_10042 (I173421,I173404,I69612);
or I_10043 (I173438,I173421,I69591);
DFFARX1 I_10044 (I173438,I2683,I172997,I173464,);
nand I_10045 (I173472,I173464,I173130);
nor I_10046 (I172974,I173472,I173280);
nor I_10047 (I172968,I173464,I173096);
DFFARX1 I_10048 (I173464,I2683,I172997,I173526,);
not I_10049 (I173534,I173526);
nor I_10050 (I172983,I173534,I173246);
not I_10051 (I173592,I2690);
DFFARX1 I_10052 (I92258,I2683,I173592,I173618,);
DFFARX1 I_10053 (I173618,I2683,I173592,I173635,);
not I_10054 (I173584,I173635);
not I_10055 (I173657,I173618);
DFFARX1 I_10056 (I92252,I2683,I173592,I173683,);
not I_10057 (I173691,I173683);
and I_10058 (I173708,I173657,I92249);
not I_10059 (I173725,I92270);
nand I_10060 (I173742,I173725,I92249);
not I_10061 (I173759,I92264);
nor I_10062 (I173776,I173759,I92255);
nand I_10063 (I173793,I173776,I92261);
nor I_10064 (I173810,I173793,I173742);
DFFARX1 I_10065 (I173810,I2683,I173592,I173560,);
not I_10066 (I173841,I173793);
not I_10067 (I173858,I92255);
nand I_10068 (I173875,I173858,I92249);
nor I_10069 (I173892,I92255,I92270);
nand I_10070 (I173572,I173708,I173892);
nand I_10071 (I173566,I173657,I92255);
nand I_10072 (I173937,I173759,I92249);
DFFARX1 I_10073 (I173937,I2683,I173592,I173581,);
DFFARX1 I_10074 (I173937,I2683,I173592,I173575,);
not I_10075 (I173982,I92249);
nor I_10076 (I173999,I173982,I92267);
and I_10077 (I174016,I173999,I92273);
or I_10078 (I174033,I174016,I92252);
DFFARX1 I_10079 (I174033,I2683,I173592,I174059,);
nand I_10080 (I174067,I174059,I173725);
nor I_10081 (I173569,I174067,I173875);
nor I_10082 (I173563,I174059,I173691);
DFFARX1 I_10083 (I174059,I2683,I173592,I174121,);
not I_10084 (I174129,I174121);
nor I_10085 (I173578,I174129,I173841);
not I_10086 (I174187,I2690);
DFFARX1 I_10087 (I802393,I2683,I174187,I174213,);
DFFARX1 I_10088 (I174213,I2683,I174187,I174230,);
not I_10089 (I174179,I174230);
not I_10090 (I174252,I174213);
DFFARX1 I_10091 (I802402,I2683,I174187,I174278,);
not I_10092 (I174286,I174278);
and I_10093 (I174303,I174252,I802396);
not I_10094 (I174320,I802390);
nand I_10095 (I174337,I174320,I802396);
not I_10096 (I174354,I802405);
nor I_10097 (I174371,I174354,I802393);
nand I_10098 (I174388,I174371,I802399);
nor I_10099 (I174405,I174388,I174337);
DFFARX1 I_10100 (I174405,I2683,I174187,I174155,);
not I_10101 (I174436,I174388);
not I_10102 (I174453,I802393);
nand I_10103 (I174470,I174453,I802396);
nor I_10104 (I174487,I802393,I802390);
nand I_10105 (I174167,I174303,I174487);
nand I_10106 (I174161,I174252,I802393);
nand I_10107 (I174532,I174354,I802396);
DFFARX1 I_10108 (I174532,I2683,I174187,I174176,);
DFFARX1 I_10109 (I174532,I2683,I174187,I174170,);
not I_10110 (I174577,I802396);
nor I_10111 (I174594,I174577,I802411);
and I_10112 (I174611,I174594,I802408);
or I_10113 (I174628,I174611,I802390);
DFFARX1 I_10114 (I174628,I2683,I174187,I174654,);
nand I_10115 (I174662,I174654,I174320);
nor I_10116 (I174164,I174662,I174470);
nor I_10117 (I174158,I174654,I174286);
DFFARX1 I_10118 (I174654,I2683,I174187,I174716,);
not I_10119 (I174724,I174716);
nor I_10120 (I174173,I174724,I174436);
not I_10121 (I174782,I2690);
DFFARX1 I_10122 (I663370,I2683,I174782,I174808,);
DFFARX1 I_10123 (I174808,I2683,I174782,I174825,);
not I_10124 (I174774,I174825);
not I_10125 (I174847,I174808);
DFFARX1 I_10126 (I663364,I2683,I174782,I174873,);
not I_10127 (I174881,I174873);
and I_10128 (I174898,I174847,I663382);
not I_10129 (I174915,I663370);
nand I_10130 (I174932,I174915,I663382);
not I_10131 (I174949,I663364);
nor I_10132 (I174966,I174949,I663376);
nand I_10133 (I174983,I174966,I663367);
nor I_10134 (I175000,I174983,I174932);
DFFARX1 I_10135 (I175000,I2683,I174782,I174750,);
not I_10136 (I175031,I174983);
not I_10137 (I175048,I663376);
nand I_10138 (I175065,I175048,I663382);
nor I_10139 (I175082,I663376,I663370);
nand I_10140 (I174762,I174898,I175082);
nand I_10141 (I174756,I174847,I663376);
nand I_10142 (I175127,I174949,I663379);
DFFARX1 I_10143 (I175127,I2683,I174782,I174771,);
DFFARX1 I_10144 (I175127,I2683,I174782,I174765,);
not I_10145 (I175172,I663379);
nor I_10146 (I175189,I175172,I663385);
and I_10147 (I175206,I175189,I663367);
or I_10148 (I175223,I175206,I663373);
DFFARX1 I_10149 (I175223,I2683,I174782,I175249,);
nand I_10150 (I175257,I175249,I174915);
nor I_10151 (I174759,I175257,I175065);
nor I_10152 (I174753,I175249,I174881);
DFFARX1 I_10153 (I175249,I2683,I174782,I175311,);
not I_10154 (I175319,I175311);
nor I_10155 (I174768,I175319,I175031);
not I_10156 (I175377,I2690);
DFFARX1 I_10157 (I105960,I2683,I175377,I175403,);
DFFARX1 I_10158 (I175403,I2683,I175377,I175420,);
not I_10159 (I175369,I175420);
not I_10160 (I175442,I175403);
DFFARX1 I_10161 (I105954,I2683,I175377,I175468,);
not I_10162 (I175476,I175468);
and I_10163 (I175493,I175442,I105951);
not I_10164 (I175510,I105972);
nand I_10165 (I175527,I175510,I105951);
not I_10166 (I175544,I105966);
nor I_10167 (I175561,I175544,I105957);
nand I_10168 (I175578,I175561,I105963);
nor I_10169 (I175595,I175578,I175527);
DFFARX1 I_10170 (I175595,I2683,I175377,I175345,);
not I_10171 (I175626,I175578);
not I_10172 (I175643,I105957);
nand I_10173 (I175660,I175643,I105951);
nor I_10174 (I175677,I105957,I105972);
nand I_10175 (I175357,I175493,I175677);
nand I_10176 (I175351,I175442,I105957);
nand I_10177 (I175722,I175544,I105951);
DFFARX1 I_10178 (I175722,I2683,I175377,I175366,);
DFFARX1 I_10179 (I175722,I2683,I175377,I175360,);
not I_10180 (I175767,I105951);
nor I_10181 (I175784,I175767,I105969);
and I_10182 (I175801,I175784,I105975);
or I_10183 (I175818,I175801,I105954);
DFFARX1 I_10184 (I175818,I2683,I175377,I175844,);
nand I_10185 (I175852,I175844,I175510);
nor I_10186 (I175354,I175852,I175660);
nor I_10187 (I175348,I175844,I175476);
DFFARX1 I_10188 (I175844,I2683,I175377,I175906,);
not I_10189 (I175914,I175906);
nor I_10190 (I175363,I175914,I175626);
not I_10191 (I175972,I2690);
DFFARX1 I_10192 (I859986,I2683,I175972,I175998,);
DFFARX1 I_10193 (I175998,I2683,I175972,I176015,);
not I_10194 (I175964,I176015);
not I_10195 (I176037,I175998);
DFFARX1 I_10196 (I859986,I2683,I175972,I176063,);
not I_10197 (I176071,I176063);
and I_10198 (I176088,I176037,I859989);
not I_10199 (I176105,I860001);
nand I_10200 (I176122,I176105,I859989);
not I_10201 (I176139,I860007);
nor I_10202 (I176156,I176139,I859998);
nand I_10203 (I176173,I176156,I860004);
nor I_10204 (I176190,I176173,I176122);
DFFARX1 I_10205 (I176190,I2683,I175972,I175940,);
not I_10206 (I176221,I176173);
not I_10207 (I176238,I859998);
nand I_10208 (I176255,I176238,I859989);
nor I_10209 (I176272,I859998,I860001);
nand I_10210 (I175952,I176088,I176272);
nand I_10211 (I175946,I176037,I859998);
nand I_10212 (I176317,I176139,I859995);
DFFARX1 I_10213 (I176317,I2683,I175972,I175961,);
DFFARX1 I_10214 (I176317,I2683,I175972,I175955,);
not I_10215 (I176362,I859995);
nor I_10216 (I176379,I176362,I859992);
and I_10217 (I176396,I176379,I860010);
or I_10218 (I176413,I176396,I859989);
DFFARX1 I_10219 (I176413,I2683,I175972,I176439,);
nand I_10220 (I176447,I176439,I176105);
nor I_10221 (I175949,I176447,I176255);
nor I_10222 (I175943,I176439,I176071);
DFFARX1 I_10223 (I176439,I2683,I175972,I176501,);
not I_10224 (I176509,I176501);
nor I_10225 (I175958,I176509,I176221);
not I_10226 (I176567,I2690);
DFFARX1 I_10227 (I909694,I2683,I176567,I176593,);
DFFARX1 I_10228 (I176593,I2683,I176567,I176610,);
not I_10229 (I176559,I176610);
not I_10230 (I176632,I176593);
DFFARX1 I_10231 (I909694,I2683,I176567,I176658,);
not I_10232 (I176666,I176658);
and I_10233 (I176683,I176632,I909697);
not I_10234 (I176700,I909709);
nand I_10235 (I176717,I176700,I909697);
not I_10236 (I176734,I909715);
nor I_10237 (I176751,I176734,I909706);
nand I_10238 (I176768,I176751,I909712);
nor I_10239 (I176785,I176768,I176717);
DFFARX1 I_10240 (I176785,I2683,I176567,I176535,);
not I_10241 (I176816,I176768);
not I_10242 (I176833,I909706);
nand I_10243 (I176850,I176833,I909697);
nor I_10244 (I176867,I909706,I909709);
nand I_10245 (I176547,I176683,I176867);
nand I_10246 (I176541,I176632,I909706);
nand I_10247 (I176912,I176734,I909703);
DFFARX1 I_10248 (I176912,I2683,I176567,I176556,);
DFFARX1 I_10249 (I176912,I2683,I176567,I176550,);
not I_10250 (I176957,I909703);
nor I_10251 (I176974,I176957,I909700);
and I_10252 (I176991,I176974,I909718);
or I_10253 (I177008,I176991,I909697);
DFFARX1 I_10254 (I177008,I2683,I176567,I177034,);
nand I_10255 (I177042,I177034,I176700);
nor I_10256 (I176544,I177042,I176850);
nor I_10257 (I176538,I177034,I176666);
DFFARX1 I_10258 (I177034,I2683,I176567,I177096,);
not I_10259 (I177104,I177096);
nor I_10260 (I176553,I177104,I176816);
not I_10261 (I177162,I2690);
DFFARX1 I_10262 (I751660,I2683,I177162,I177188,);
DFFARX1 I_10263 (I177188,I2683,I177162,I177205,);
not I_10264 (I177154,I177205);
not I_10265 (I177227,I177188);
DFFARX1 I_10266 (I751669,I2683,I177162,I177253,);
not I_10267 (I177261,I177253);
and I_10268 (I177278,I177227,I751657);
not I_10269 (I177295,I751648);
nand I_10270 (I177312,I177295,I751657);
not I_10271 (I177329,I751654);
nor I_10272 (I177346,I177329,I751672);
nand I_10273 (I177363,I177346,I751645);
nor I_10274 (I177380,I177363,I177312);
DFFARX1 I_10275 (I177380,I2683,I177162,I177130,);
not I_10276 (I177411,I177363);
not I_10277 (I177428,I751672);
nand I_10278 (I177445,I177428,I751657);
nor I_10279 (I177462,I751672,I751648);
nand I_10280 (I177142,I177278,I177462);
nand I_10281 (I177136,I177227,I751672);
nand I_10282 (I177507,I177329,I751651);
DFFARX1 I_10283 (I177507,I2683,I177162,I177151,);
DFFARX1 I_10284 (I177507,I2683,I177162,I177145,);
not I_10285 (I177552,I751651);
nor I_10286 (I177569,I177552,I751663);
and I_10287 (I177586,I177569,I751645);
or I_10288 (I177603,I177586,I751666);
DFFARX1 I_10289 (I177603,I2683,I177162,I177629,);
nand I_10290 (I177637,I177629,I177295);
nor I_10291 (I177139,I177637,I177445);
nor I_10292 (I177133,I177629,I177261);
DFFARX1 I_10293 (I177629,I2683,I177162,I177691,);
not I_10294 (I177699,I177691);
nor I_10295 (I177148,I177699,I177411);
not I_10296 (I177757,I2690);
DFFARX1 I_10297 (I628588,I2683,I177757,I177783,);
DFFARX1 I_10298 (I177783,I2683,I177757,I177800,);
not I_10299 (I177749,I177800);
not I_10300 (I177822,I177783);
DFFARX1 I_10301 (I628582,I2683,I177757,I177848,);
not I_10302 (I177856,I177848);
and I_10303 (I177873,I177822,I628600);
not I_10304 (I177890,I628588);
nand I_10305 (I177907,I177890,I628600);
not I_10306 (I177924,I628582);
nor I_10307 (I177941,I177924,I628594);
nand I_10308 (I177958,I177941,I628585);
nor I_10309 (I177975,I177958,I177907);
DFFARX1 I_10310 (I177975,I2683,I177757,I177725,);
not I_10311 (I178006,I177958);
not I_10312 (I178023,I628594);
nand I_10313 (I178040,I178023,I628600);
nor I_10314 (I178057,I628594,I628588);
nand I_10315 (I177737,I177873,I178057);
nand I_10316 (I177731,I177822,I628594);
nand I_10317 (I178102,I177924,I628597);
DFFARX1 I_10318 (I178102,I2683,I177757,I177746,);
DFFARX1 I_10319 (I178102,I2683,I177757,I177740,);
not I_10320 (I178147,I628597);
nor I_10321 (I178164,I178147,I628603);
and I_10322 (I178181,I178164,I628585);
or I_10323 (I178198,I178181,I628591);
DFFARX1 I_10324 (I178198,I2683,I177757,I178224,);
nand I_10325 (I178232,I178224,I177890);
nor I_10326 (I177734,I178232,I178040);
nor I_10327 (I177728,I178224,I177856);
DFFARX1 I_10328 (I178224,I2683,I177757,I178286,);
not I_10329 (I178294,I178286);
nor I_10330 (I177743,I178294,I178006);
not I_10331 (I178352,I2690);
DFFARX1 I_10332 (I732280,I2683,I178352,I178378,);
DFFARX1 I_10333 (I178378,I2683,I178352,I178395,);
not I_10334 (I178344,I178395);
not I_10335 (I178417,I178378);
DFFARX1 I_10336 (I732289,I2683,I178352,I178443,);
not I_10337 (I178451,I178443);
and I_10338 (I178468,I178417,I732277);
not I_10339 (I178485,I732268);
nand I_10340 (I178502,I178485,I732277);
not I_10341 (I178519,I732274);
nor I_10342 (I178536,I178519,I732292);
nand I_10343 (I178553,I178536,I732265);
nor I_10344 (I178570,I178553,I178502);
DFFARX1 I_10345 (I178570,I2683,I178352,I178320,);
not I_10346 (I178601,I178553);
not I_10347 (I178618,I732292);
nand I_10348 (I178635,I178618,I732277);
nor I_10349 (I178652,I732292,I732268);
nand I_10350 (I178332,I178468,I178652);
nand I_10351 (I178326,I178417,I732292);
nand I_10352 (I178697,I178519,I732271);
DFFARX1 I_10353 (I178697,I2683,I178352,I178341,);
DFFARX1 I_10354 (I178697,I2683,I178352,I178335,);
not I_10355 (I178742,I732271);
nor I_10356 (I178759,I178742,I732283);
and I_10357 (I178776,I178759,I732265);
or I_10358 (I178793,I178776,I732286);
DFFARX1 I_10359 (I178793,I2683,I178352,I178819,);
nand I_10360 (I178827,I178819,I178485);
nor I_10361 (I178329,I178827,I178635);
nor I_10362 (I178323,I178819,I178451);
DFFARX1 I_10363 (I178819,I2683,I178352,I178881,);
not I_10364 (I178889,I178881);
nor I_10365 (I178338,I178889,I178601);
not I_10366 (I178947,I2690);
DFFARX1 I_10367 (I531830,I2683,I178947,I178973,);
DFFARX1 I_10368 (I178973,I2683,I178947,I178990,);
not I_10369 (I178939,I178990);
not I_10370 (I179012,I178973);
DFFARX1 I_10371 (I531827,I2683,I178947,I179038,);
not I_10372 (I179046,I179038);
and I_10373 (I179063,I179012,I531833);
not I_10374 (I179080,I531818);
nand I_10375 (I179097,I179080,I531833);
not I_10376 (I179114,I531821);
nor I_10377 (I179131,I179114,I531842);
nand I_10378 (I179148,I179131,I531839);
nor I_10379 (I179165,I179148,I179097);
DFFARX1 I_10380 (I179165,I2683,I178947,I178915,);
not I_10381 (I179196,I179148);
not I_10382 (I179213,I531842);
nand I_10383 (I179230,I179213,I531833);
nor I_10384 (I179247,I531842,I531818);
nand I_10385 (I178927,I179063,I179247);
nand I_10386 (I178921,I179012,I531842);
nand I_10387 (I179292,I179114,I531818);
DFFARX1 I_10388 (I179292,I2683,I178947,I178936,);
DFFARX1 I_10389 (I179292,I2683,I178947,I178930,);
not I_10390 (I179337,I531818);
nor I_10391 (I179354,I179337,I531824);
and I_10392 (I179371,I179354,I531836);
or I_10393 (I179388,I179371,I531821);
DFFARX1 I_10394 (I179388,I2683,I178947,I179414,);
nand I_10395 (I179422,I179414,I179080);
nor I_10396 (I178924,I179422,I179230);
nor I_10397 (I178918,I179414,I179046);
DFFARX1 I_10398 (I179414,I2683,I178947,I179476,);
not I_10399 (I179484,I179476);
nor I_10400 (I178933,I179484,I179196);
not I_10401 (I179542,I2690);
DFFARX1 I_10402 (I938016,I2683,I179542,I179568,);
DFFARX1 I_10403 (I179568,I2683,I179542,I179585,);
not I_10404 (I179534,I179585);
not I_10405 (I179607,I179568);
DFFARX1 I_10406 (I938016,I2683,I179542,I179633,);
not I_10407 (I179641,I179633);
and I_10408 (I179658,I179607,I938019);
not I_10409 (I179675,I938031);
nand I_10410 (I179692,I179675,I938019);
not I_10411 (I179709,I938037);
nor I_10412 (I179726,I179709,I938028);
nand I_10413 (I179743,I179726,I938034);
nor I_10414 (I179760,I179743,I179692);
DFFARX1 I_10415 (I179760,I2683,I179542,I179510,);
not I_10416 (I179791,I179743);
not I_10417 (I179808,I938028);
nand I_10418 (I179825,I179808,I938019);
nor I_10419 (I179842,I938028,I938031);
nand I_10420 (I179522,I179658,I179842);
nand I_10421 (I179516,I179607,I938028);
nand I_10422 (I179887,I179709,I938025);
DFFARX1 I_10423 (I179887,I2683,I179542,I179531,);
DFFARX1 I_10424 (I179887,I2683,I179542,I179525,);
not I_10425 (I179932,I938025);
nor I_10426 (I179949,I179932,I938022);
and I_10427 (I179966,I179949,I938040);
or I_10428 (I179983,I179966,I938019);
DFFARX1 I_10429 (I179983,I2683,I179542,I180009,);
nand I_10430 (I180017,I180009,I179675);
nor I_10431 (I179519,I180017,I179825);
nor I_10432 (I179513,I180009,I179641);
DFFARX1 I_10433 (I180009,I2683,I179542,I180071,);
not I_10434 (I180079,I180071);
nor I_10435 (I179528,I180079,I179791);
not I_10436 (I180137,I2690);
DFFARX1 I_10437 (I650195,I2683,I180137,I180163,);
DFFARX1 I_10438 (I180163,I2683,I180137,I180180,);
not I_10439 (I180129,I180180);
not I_10440 (I180202,I180163);
DFFARX1 I_10441 (I650189,I2683,I180137,I180228,);
not I_10442 (I180236,I180228);
and I_10443 (I180253,I180202,I650207);
not I_10444 (I180270,I650195);
nand I_10445 (I180287,I180270,I650207);
not I_10446 (I180304,I650189);
nor I_10447 (I180321,I180304,I650201);
nand I_10448 (I180338,I180321,I650192);
nor I_10449 (I180355,I180338,I180287);
DFFARX1 I_10450 (I180355,I2683,I180137,I180105,);
not I_10451 (I180386,I180338);
not I_10452 (I180403,I650201);
nand I_10453 (I180420,I180403,I650207);
nor I_10454 (I180437,I650201,I650195);
nand I_10455 (I180117,I180253,I180437);
nand I_10456 (I180111,I180202,I650201);
nand I_10457 (I180482,I180304,I650204);
DFFARX1 I_10458 (I180482,I2683,I180137,I180126,);
DFFARX1 I_10459 (I180482,I2683,I180137,I180120,);
not I_10460 (I180527,I650204);
nor I_10461 (I180544,I180527,I650210);
and I_10462 (I180561,I180544,I650192);
or I_10463 (I180578,I180561,I650198);
DFFARX1 I_10464 (I180578,I2683,I180137,I180604,);
nand I_10465 (I180612,I180604,I180270);
nor I_10466 (I180114,I180612,I180420);
nor I_10467 (I180108,I180604,I180236);
DFFARX1 I_10468 (I180604,I2683,I180137,I180666,);
not I_10469 (I180674,I180666);
nor I_10470 (I180123,I180674,I180386);
not I_10471 (I180732,I2690);
DFFARX1 I_10472 (I313351,I2683,I180732,I180758,);
DFFARX1 I_10473 (I180758,I2683,I180732,I180775,);
not I_10474 (I180724,I180775);
not I_10475 (I180797,I180758);
DFFARX1 I_10476 (I313366,I2683,I180732,I180823,);
not I_10477 (I180831,I180823);
and I_10478 (I180848,I180797,I313363);
not I_10479 (I180865,I313351);
nand I_10480 (I180882,I180865,I313363);
not I_10481 (I180899,I313360);
nor I_10482 (I180916,I180899,I313375);
nand I_10483 (I180933,I180916,I313372);
nor I_10484 (I180950,I180933,I180882);
DFFARX1 I_10485 (I180950,I2683,I180732,I180700,);
not I_10486 (I180981,I180933);
not I_10487 (I180998,I313375);
nand I_10488 (I181015,I180998,I313363);
nor I_10489 (I181032,I313375,I313351);
nand I_10490 (I180712,I180848,I181032);
nand I_10491 (I180706,I180797,I313375);
nand I_10492 (I181077,I180899,I313369);
DFFARX1 I_10493 (I181077,I2683,I180732,I180721,);
DFFARX1 I_10494 (I181077,I2683,I180732,I180715,);
not I_10495 (I181122,I313369);
nor I_10496 (I181139,I181122,I313357);
and I_10497 (I181156,I181139,I313378);
or I_10498 (I181173,I181156,I313354);
DFFARX1 I_10499 (I181173,I2683,I180732,I181199,);
nand I_10500 (I181207,I181199,I180865);
nor I_10501 (I180709,I181207,I181015);
nor I_10502 (I180703,I181199,I180831);
DFFARX1 I_10503 (I181199,I2683,I180732,I181261,);
not I_10504 (I181269,I181261);
nor I_10505 (I180718,I181269,I180981);
not I_10506 (I181327,I2690);
DFFARX1 I_10507 (I901024,I2683,I181327,I181353,);
DFFARX1 I_10508 (I181353,I2683,I181327,I181370,);
not I_10509 (I181319,I181370);
not I_10510 (I181392,I181353);
DFFARX1 I_10511 (I901024,I2683,I181327,I181418,);
not I_10512 (I181426,I181418);
and I_10513 (I181443,I181392,I901027);
not I_10514 (I181460,I901039);
nand I_10515 (I181477,I181460,I901027);
not I_10516 (I181494,I901045);
nor I_10517 (I181511,I181494,I901036);
nand I_10518 (I181528,I181511,I901042);
nor I_10519 (I181545,I181528,I181477);
DFFARX1 I_10520 (I181545,I2683,I181327,I181295,);
not I_10521 (I181576,I181528);
not I_10522 (I181593,I901036);
nand I_10523 (I181610,I181593,I901027);
nor I_10524 (I181627,I901036,I901039);
nand I_10525 (I181307,I181443,I181627);
nand I_10526 (I181301,I181392,I901036);
nand I_10527 (I181672,I181494,I901033);
DFFARX1 I_10528 (I181672,I2683,I181327,I181316,);
DFFARX1 I_10529 (I181672,I2683,I181327,I181310,);
not I_10530 (I181717,I901033);
nor I_10531 (I181734,I181717,I901030);
and I_10532 (I181751,I181734,I901048);
or I_10533 (I181768,I181751,I901027);
DFFARX1 I_10534 (I181768,I2683,I181327,I181794,);
nand I_10535 (I181802,I181794,I181460);
nor I_10536 (I181304,I181802,I181610);
nor I_10537 (I181298,I181794,I181426);
DFFARX1 I_10538 (I181794,I2683,I181327,I181856,);
not I_10539 (I181864,I181856);
nor I_10540 (I181313,I181864,I181576);
not I_10541 (I181922,I2690);
DFFARX1 I_10542 (I785898,I2683,I181922,I181948,);
DFFARX1 I_10543 (I181948,I2683,I181922,I181965,);
not I_10544 (I181914,I181965);
not I_10545 (I181987,I181948);
DFFARX1 I_10546 (I785907,I2683,I181922,I182013,);
not I_10547 (I182021,I182013);
and I_10548 (I182038,I181987,I785895);
not I_10549 (I182055,I785886);
nand I_10550 (I182072,I182055,I785895);
not I_10551 (I182089,I785892);
nor I_10552 (I182106,I182089,I785910);
nand I_10553 (I182123,I182106,I785883);
nor I_10554 (I182140,I182123,I182072);
DFFARX1 I_10555 (I182140,I2683,I181922,I181890,);
not I_10556 (I182171,I182123);
not I_10557 (I182188,I785910);
nand I_10558 (I182205,I182188,I785895);
nor I_10559 (I182222,I785910,I785886);
nand I_10560 (I181902,I182038,I182222);
nand I_10561 (I181896,I181987,I785910);
nand I_10562 (I182267,I182089,I785889);
DFFARX1 I_10563 (I182267,I2683,I181922,I181911,);
DFFARX1 I_10564 (I182267,I2683,I181922,I181905,);
not I_10565 (I182312,I785889);
nor I_10566 (I182329,I182312,I785901);
and I_10567 (I182346,I182329,I785883);
or I_10568 (I182363,I182346,I785904);
DFFARX1 I_10569 (I182363,I2683,I181922,I182389,);
nand I_10570 (I182397,I182389,I182055);
nor I_10571 (I181899,I182397,I182205);
nor I_10572 (I181893,I182389,I182021);
DFFARX1 I_10573 (I182389,I2683,I181922,I182451,);
not I_10574 (I182459,I182451);
nor I_10575 (I181908,I182459,I182171);
not I_10576 (I182517,I2690);
DFFARX1 I_10577 (I430034,I2683,I182517,I182543,);
DFFARX1 I_10578 (I182543,I2683,I182517,I182560,);
not I_10579 (I182509,I182560);
not I_10580 (I182582,I182543);
DFFARX1 I_10581 (I430028,I2683,I182517,I182608,);
not I_10582 (I182616,I182608);
and I_10583 (I182633,I182582,I430043);
not I_10584 (I182650,I430040);
nand I_10585 (I182667,I182650,I430043);
not I_10586 (I182684,I430031);
nor I_10587 (I182701,I182684,I430022);
nand I_10588 (I182718,I182701,I430025);
nor I_10589 (I182735,I182718,I182667);
DFFARX1 I_10590 (I182735,I2683,I182517,I182485,);
not I_10591 (I182766,I182718);
not I_10592 (I182783,I430022);
nand I_10593 (I182800,I182783,I430043);
nor I_10594 (I182817,I430022,I430040);
nand I_10595 (I182497,I182633,I182817);
nand I_10596 (I182491,I182582,I430022);
nand I_10597 (I182862,I182684,I430046);
DFFARX1 I_10598 (I182862,I2683,I182517,I182506,);
DFFARX1 I_10599 (I182862,I2683,I182517,I182500,);
not I_10600 (I182907,I430046);
nor I_10601 (I182924,I182907,I430037);
and I_10602 (I182941,I182924,I430022);
or I_10603 (I182958,I182941,I430025);
DFFARX1 I_10604 (I182958,I2683,I182517,I182984,);
nand I_10605 (I182992,I182984,I182650);
nor I_10606 (I182494,I182992,I182800);
nor I_10607 (I182488,I182984,I182616);
DFFARX1 I_10608 (I182984,I2683,I182517,I183046,);
not I_10609 (I183054,I183046);
nor I_10610 (I182503,I183054,I182766);
not I_10611 (I183112,I2690);
DFFARX1 I_10612 (I30614,I2683,I183112,I183138,);
DFFARX1 I_10613 (I183138,I2683,I183112,I183155,);
not I_10614 (I183104,I183155);
not I_10615 (I183177,I183138);
DFFARX1 I_10616 (I30590,I2683,I183112,I183203,);
not I_10617 (I183211,I183203);
and I_10618 (I183228,I183177,I30605);
not I_10619 (I183245,I30593);
nand I_10620 (I183262,I183245,I30605);
not I_10621 (I183279,I30596);
nor I_10622 (I183296,I183279,I30608);
nand I_10623 (I183313,I183296,I30599);
nor I_10624 (I183330,I183313,I183262);
DFFARX1 I_10625 (I183330,I2683,I183112,I183080,);
not I_10626 (I183361,I183313);
not I_10627 (I183378,I30608);
nand I_10628 (I183395,I183378,I30605);
nor I_10629 (I183412,I30608,I30593);
nand I_10630 (I183092,I183228,I183412);
nand I_10631 (I183086,I183177,I30608);
nand I_10632 (I183457,I183279,I30602);
DFFARX1 I_10633 (I183457,I2683,I183112,I183101,);
DFFARX1 I_10634 (I183457,I2683,I183112,I183095,);
not I_10635 (I183502,I30602);
nor I_10636 (I183519,I183502,I30593);
and I_10637 (I183536,I183519,I30590);
or I_10638 (I183553,I183536,I30611);
DFFARX1 I_10639 (I183553,I2683,I183112,I183579,);
nand I_10640 (I183587,I183579,I183245);
nor I_10641 (I183089,I183587,I183395);
nor I_10642 (I183083,I183579,I183211);
DFFARX1 I_10643 (I183579,I2683,I183112,I183641,);
not I_10644 (I183649,I183641);
nor I_10645 (I183098,I183649,I183361);
not I_10646 (I183707,I2690);
DFFARX1 I_10647 (I898712,I2683,I183707,I183733,);
DFFARX1 I_10648 (I183733,I2683,I183707,I183750,);
not I_10649 (I183699,I183750);
not I_10650 (I183772,I183733);
DFFARX1 I_10651 (I898712,I2683,I183707,I183798,);
not I_10652 (I183806,I183798);
and I_10653 (I183823,I183772,I898715);
not I_10654 (I183840,I898727);
nand I_10655 (I183857,I183840,I898715);
not I_10656 (I183874,I898733);
nor I_10657 (I183891,I183874,I898724);
nand I_10658 (I183908,I183891,I898730);
nor I_10659 (I183925,I183908,I183857);
DFFARX1 I_10660 (I183925,I2683,I183707,I183675,);
not I_10661 (I183956,I183908);
not I_10662 (I183973,I898724);
nand I_10663 (I183990,I183973,I898715);
nor I_10664 (I184007,I898724,I898727);
nand I_10665 (I183687,I183823,I184007);
nand I_10666 (I183681,I183772,I898724);
nand I_10667 (I184052,I183874,I898721);
DFFARX1 I_10668 (I184052,I2683,I183707,I183696,);
DFFARX1 I_10669 (I184052,I2683,I183707,I183690,);
not I_10670 (I184097,I898721);
nor I_10671 (I184114,I184097,I898718);
and I_10672 (I184131,I184114,I898736);
or I_10673 (I184148,I184131,I898715);
DFFARX1 I_10674 (I184148,I2683,I183707,I184174,);
nand I_10675 (I184182,I184174,I183840);
nor I_10676 (I183684,I184182,I183990);
nor I_10677 (I183678,I184174,I183806);
DFFARX1 I_10678 (I184174,I2683,I183707,I184236,);
not I_10679 (I184244,I184236);
nor I_10680 (I183693,I184244,I183956);
not I_10681 (I184302,I2690);
DFFARX1 I_10682 (I944952,I2683,I184302,I184328,);
DFFARX1 I_10683 (I184328,I2683,I184302,I184345,);
not I_10684 (I184294,I184345);
not I_10685 (I184367,I184328);
DFFARX1 I_10686 (I944952,I2683,I184302,I184393,);
not I_10687 (I184401,I184393);
and I_10688 (I184418,I184367,I944955);
not I_10689 (I184435,I944967);
nand I_10690 (I184452,I184435,I944955);
not I_10691 (I184469,I944973);
nor I_10692 (I184486,I184469,I944964);
nand I_10693 (I184503,I184486,I944970);
nor I_10694 (I184520,I184503,I184452);
DFFARX1 I_10695 (I184520,I2683,I184302,I184270,);
not I_10696 (I184551,I184503);
not I_10697 (I184568,I944964);
nand I_10698 (I184585,I184568,I944955);
nor I_10699 (I184602,I944964,I944967);
nand I_10700 (I184282,I184418,I184602);
nand I_10701 (I184276,I184367,I944964);
nand I_10702 (I184647,I184469,I944961);
DFFARX1 I_10703 (I184647,I2683,I184302,I184291,);
DFFARX1 I_10704 (I184647,I2683,I184302,I184285,);
not I_10705 (I184692,I944961);
nor I_10706 (I184709,I184692,I944958);
and I_10707 (I184726,I184709,I944976);
or I_10708 (I184743,I184726,I944955);
DFFARX1 I_10709 (I184743,I2683,I184302,I184769,);
nand I_10710 (I184777,I184769,I184435);
nor I_10711 (I184279,I184777,I184585);
nor I_10712 (I184273,I184769,I184401);
DFFARX1 I_10713 (I184769,I2683,I184302,I184831,);
not I_10714 (I184839,I184831);
nor I_10715 (I184288,I184839,I184551);
not I_10716 (I184897,I2690);
DFFARX1 I_10717 (I548592,I2683,I184897,I184923,);
DFFARX1 I_10718 (I184923,I2683,I184897,I184940,);
not I_10719 (I184889,I184940);
not I_10720 (I184962,I184923);
DFFARX1 I_10721 (I548589,I2683,I184897,I184988,);
not I_10722 (I184996,I184988);
and I_10723 (I185013,I184962,I548595);
not I_10724 (I185030,I548580);
nand I_10725 (I185047,I185030,I548595);
not I_10726 (I185064,I548583);
nor I_10727 (I185081,I185064,I548604);
nand I_10728 (I185098,I185081,I548601);
nor I_10729 (I185115,I185098,I185047);
DFFARX1 I_10730 (I185115,I2683,I184897,I184865,);
not I_10731 (I185146,I185098);
not I_10732 (I185163,I548604);
nand I_10733 (I185180,I185163,I548595);
nor I_10734 (I185197,I548604,I548580);
nand I_10735 (I184877,I185013,I185197);
nand I_10736 (I184871,I184962,I548604);
nand I_10737 (I185242,I185064,I548580);
DFFARX1 I_10738 (I185242,I2683,I184897,I184886,);
DFFARX1 I_10739 (I185242,I2683,I184897,I184880,);
not I_10740 (I185287,I548580);
nor I_10741 (I185304,I185287,I548586);
and I_10742 (I185321,I185304,I548598);
or I_10743 (I185338,I185321,I548583);
DFFARX1 I_10744 (I185338,I2683,I184897,I185364,);
nand I_10745 (I185372,I185364,I185030);
nor I_10746 (I184874,I185372,I185180);
nor I_10747 (I184868,I185364,I184996);
DFFARX1 I_10748 (I185364,I2683,I184897,I185426,);
not I_10749 (I185434,I185426);
nor I_10750 (I184883,I185434,I185146);
not I_10751 (I185492,I2690);
DFFARX1 I_10752 (I586740,I2683,I185492,I185518,);
DFFARX1 I_10753 (I185518,I2683,I185492,I185535,);
not I_10754 (I185484,I185535);
not I_10755 (I185557,I185518);
DFFARX1 I_10756 (I586737,I2683,I185492,I185583,);
not I_10757 (I185591,I185583);
and I_10758 (I185608,I185557,I586743);
not I_10759 (I185625,I586728);
nand I_10760 (I185642,I185625,I586743);
not I_10761 (I185659,I586731);
nor I_10762 (I185676,I185659,I586752);
nand I_10763 (I185693,I185676,I586749);
nor I_10764 (I185710,I185693,I185642);
DFFARX1 I_10765 (I185710,I2683,I185492,I185460,);
not I_10766 (I185741,I185693);
not I_10767 (I185758,I586752);
nand I_10768 (I185775,I185758,I586743);
nor I_10769 (I185792,I586752,I586728);
nand I_10770 (I185472,I185608,I185792);
nand I_10771 (I185466,I185557,I586752);
nand I_10772 (I185837,I185659,I586728);
DFFARX1 I_10773 (I185837,I2683,I185492,I185481,);
DFFARX1 I_10774 (I185837,I2683,I185492,I185475,);
not I_10775 (I185882,I586728);
nor I_10776 (I185899,I185882,I586734);
and I_10777 (I185916,I185899,I586746);
or I_10778 (I185933,I185916,I586731);
DFFARX1 I_10779 (I185933,I2683,I185492,I185959,);
nand I_10780 (I185967,I185959,I185625);
nor I_10781 (I185469,I185967,I185775);
nor I_10782 (I185463,I185959,I185591);
DFFARX1 I_10783 (I185959,I2683,I185492,I186021,);
not I_10784 (I186029,I186021);
nor I_10785 (I185478,I186029,I185741);
not I_10786 (I186087,I2690);
DFFARX1 I_10787 (I462473,I2683,I186087,I186113,);
DFFARX1 I_10788 (I186113,I2683,I186087,I186130,);
not I_10789 (I186079,I186130);
not I_10790 (I186152,I186113);
DFFARX1 I_10791 (I462464,I2683,I186087,I186178,);
not I_10792 (I186186,I186178);
and I_10793 (I186203,I186152,I462482);
not I_10794 (I186220,I462479);
nand I_10795 (I186237,I186220,I462482);
not I_10796 (I186254,I462458);
nor I_10797 (I186271,I186254,I462461);
nand I_10798 (I186288,I186271,I462470);
nor I_10799 (I186305,I186288,I186237);
DFFARX1 I_10800 (I186305,I2683,I186087,I186055,);
not I_10801 (I186336,I186288);
not I_10802 (I186353,I462461);
nand I_10803 (I186370,I186353,I462482);
nor I_10804 (I186387,I462461,I462479);
nand I_10805 (I186067,I186203,I186387);
nand I_10806 (I186061,I186152,I462461);
nand I_10807 (I186432,I186254,I462476);
DFFARX1 I_10808 (I186432,I2683,I186087,I186076,);
DFFARX1 I_10809 (I186432,I2683,I186087,I186070,);
not I_10810 (I186477,I462476);
nor I_10811 (I186494,I186477,I462458);
and I_10812 (I186511,I186494,I462467);
or I_10813 (I186528,I186511,I462461);
DFFARX1 I_10814 (I186528,I2683,I186087,I186554,);
nand I_10815 (I186562,I186554,I186220);
nor I_10816 (I186064,I186562,I186370);
nor I_10817 (I186058,I186554,I186186);
DFFARX1 I_10818 (I186554,I2683,I186087,I186616,);
not I_10819 (I186624,I186616);
nor I_10820 (I186073,I186624,I186336);
not I_10821 (I186682,I2690);
DFFARX1 I_10822 (I1088810,I2683,I186682,I186708,);
DFFARX1 I_10823 (I186708,I2683,I186682,I186725,);
not I_10824 (I186674,I186725);
not I_10825 (I186747,I186708);
DFFARX1 I_10826 (I1088801,I2683,I186682,I186773,);
not I_10827 (I186781,I186773);
and I_10828 (I186798,I186747,I1088795);
not I_10829 (I186815,I1088789);
nand I_10830 (I186832,I186815,I1088795);
not I_10831 (I186849,I1088816);
nor I_10832 (I186866,I186849,I1088789);
nand I_10833 (I186883,I186866,I1088813);
nor I_10834 (I186900,I186883,I186832);
DFFARX1 I_10835 (I186900,I2683,I186682,I186650,);
not I_10836 (I186931,I186883);
not I_10837 (I186948,I1088789);
nand I_10838 (I186965,I186948,I1088795);
nor I_10839 (I186982,I1088789,I1088789);
nand I_10840 (I186662,I186798,I186982);
nand I_10841 (I186656,I186747,I1088789);
nand I_10842 (I187027,I186849,I1088798);
DFFARX1 I_10843 (I187027,I2683,I186682,I186671,);
DFFARX1 I_10844 (I187027,I2683,I186682,I186665,);
not I_10845 (I187072,I1088798);
nor I_10846 (I187089,I187072,I1088804);
and I_10847 (I187106,I187089,I1088807);
or I_10848 (I187123,I187106,I1088792);
DFFARX1 I_10849 (I187123,I2683,I186682,I187149,);
nand I_10850 (I187157,I187149,I186815);
nor I_10851 (I186659,I187157,I186965);
nor I_10852 (I186653,I187149,I186781);
DFFARX1 I_10853 (I187149,I2683,I186682,I187211,);
not I_10854 (I187219,I187211);
nor I_10855 (I186668,I187219,I186931);
not I_10856 (I187277,I2690);
DFFARX1 I_10857 (I964112,I2683,I187277,I187303,);
DFFARX1 I_10858 (I187303,I2683,I187277,I187320,);
not I_10859 (I187269,I187320);
not I_10860 (I187342,I187303);
DFFARX1 I_10861 (I964097,I2683,I187277,I187368,);
not I_10862 (I187376,I187368);
and I_10863 (I187393,I187342,I964115);
not I_10864 (I187410,I964097);
nand I_10865 (I187427,I187410,I964115);
not I_10866 (I187444,I964118);
nor I_10867 (I187461,I187444,I964109);
nand I_10868 (I187478,I187461,I964106);
nor I_10869 (I187495,I187478,I187427);
DFFARX1 I_10870 (I187495,I2683,I187277,I187245,);
not I_10871 (I187526,I187478);
not I_10872 (I187543,I964109);
nand I_10873 (I187560,I187543,I964115);
nor I_10874 (I187577,I964109,I964097);
nand I_10875 (I187257,I187393,I187577);
nand I_10876 (I187251,I187342,I964109);
nand I_10877 (I187622,I187444,I964103);
DFFARX1 I_10878 (I187622,I2683,I187277,I187266,);
DFFARX1 I_10879 (I187622,I2683,I187277,I187260,);
not I_10880 (I187667,I964103);
nor I_10881 (I187684,I187667,I964094);
and I_10882 (I187701,I187684,I964100);
or I_10883 (I187718,I187701,I964094);
DFFARX1 I_10884 (I187718,I2683,I187277,I187744,);
nand I_10885 (I187752,I187744,I187410);
nor I_10886 (I187254,I187752,I187560);
nor I_10887 (I187248,I187744,I187376);
DFFARX1 I_10888 (I187744,I2683,I187277,I187806,);
not I_10889 (I187814,I187806);
nor I_10890 (I187263,I187814,I187526);
not I_10891 (I187872,I2690);
DFFARX1 I_10892 (I737448,I2683,I187872,I187898,);
DFFARX1 I_10893 (I187898,I2683,I187872,I187915,);
not I_10894 (I187864,I187915);
not I_10895 (I187937,I187898);
DFFARX1 I_10896 (I737457,I2683,I187872,I187963,);
not I_10897 (I187971,I187963);
and I_10898 (I187988,I187937,I737445);
not I_10899 (I188005,I737436);
nand I_10900 (I188022,I188005,I737445);
not I_10901 (I188039,I737442);
nor I_10902 (I188056,I188039,I737460);
nand I_10903 (I188073,I188056,I737433);
nor I_10904 (I188090,I188073,I188022);
DFFARX1 I_10905 (I188090,I2683,I187872,I187840,);
not I_10906 (I188121,I188073);
not I_10907 (I188138,I737460);
nand I_10908 (I188155,I188138,I737445);
nor I_10909 (I188172,I737460,I737436);
nand I_10910 (I187852,I187988,I188172);
nand I_10911 (I187846,I187937,I737460);
nand I_10912 (I188217,I188039,I737439);
DFFARX1 I_10913 (I188217,I2683,I187872,I187861,);
DFFARX1 I_10914 (I188217,I2683,I187872,I187855,);
not I_10915 (I188262,I737439);
nor I_10916 (I188279,I188262,I737451);
and I_10917 (I188296,I188279,I737433);
or I_10918 (I188313,I188296,I737454);
DFFARX1 I_10919 (I188313,I2683,I187872,I188339,);
nand I_10920 (I188347,I188339,I188005);
nor I_10921 (I187849,I188347,I188155);
nor I_10922 (I187843,I188339,I187971);
DFFARX1 I_10923 (I188339,I2683,I187872,I188401,);
not I_10924 (I188409,I188401);
nor I_10925 (I187858,I188409,I188121);
not I_10926 (I188467,I2690);
DFFARX1 I_10927 (I771040,I2683,I188467,I188493,);
DFFARX1 I_10928 (I188493,I2683,I188467,I188510,);
not I_10929 (I188459,I188510);
not I_10930 (I188532,I188493);
DFFARX1 I_10931 (I771049,I2683,I188467,I188558,);
not I_10932 (I188566,I188558);
and I_10933 (I188583,I188532,I771037);
not I_10934 (I188600,I771028);
nand I_10935 (I188617,I188600,I771037);
not I_10936 (I188634,I771034);
nor I_10937 (I188651,I188634,I771052);
nand I_10938 (I188668,I188651,I771025);
nor I_10939 (I188685,I188668,I188617);
DFFARX1 I_10940 (I188685,I2683,I188467,I188435,);
not I_10941 (I188716,I188668);
not I_10942 (I188733,I771052);
nand I_10943 (I188750,I188733,I771037);
nor I_10944 (I188767,I771052,I771028);
nand I_10945 (I188447,I188583,I188767);
nand I_10946 (I188441,I188532,I771052);
nand I_10947 (I188812,I188634,I771031);
DFFARX1 I_10948 (I188812,I2683,I188467,I188456,);
DFFARX1 I_10949 (I188812,I2683,I188467,I188450,);
not I_10950 (I188857,I771031);
nor I_10951 (I188874,I188857,I771043);
and I_10952 (I188891,I188874,I771025);
or I_10953 (I188908,I188891,I771046);
DFFARX1 I_10954 (I188908,I2683,I188467,I188934,);
nand I_10955 (I188942,I188934,I188600);
nor I_10956 (I188444,I188942,I188750);
nor I_10957 (I188438,I188934,I188566);
DFFARX1 I_10958 (I188934,I2683,I188467,I188996,);
not I_10959 (I189004,I188996);
nor I_10960 (I188453,I189004,I188716);
not I_10961 (I189062,I2690);
DFFARX1 I_10962 (I529518,I2683,I189062,I189088,);
DFFARX1 I_10963 (I189088,I2683,I189062,I189105,);
not I_10964 (I189054,I189105);
not I_10965 (I189127,I189088);
DFFARX1 I_10966 (I529515,I2683,I189062,I189153,);
not I_10967 (I189161,I189153);
and I_10968 (I189178,I189127,I529521);
not I_10969 (I189195,I529506);
nand I_10970 (I189212,I189195,I529521);
not I_10971 (I189229,I529509);
nor I_10972 (I189246,I189229,I529530);
nand I_10973 (I189263,I189246,I529527);
nor I_10974 (I189280,I189263,I189212);
DFFARX1 I_10975 (I189280,I2683,I189062,I189030,);
not I_10976 (I189311,I189263);
not I_10977 (I189328,I529530);
nand I_10978 (I189345,I189328,I529521);
nor I_10979 (I189362,I529530,I529506);
nand I_10980 (I189042,I189178,I189362);
nand I_10981 (I189036,I189127,I529530);
nand I_10982 (I189407,I189229,I529506);
DFFARX1 I_10983 (I189407,I2683,I189062,I189051,);
DFFARX1 I_10984 (I189407,I2683,I189062,I189045,);
not I_10985 (I189452,I529506);
nor I_10986 (I189469,I189452,I529512);
and I_10987 (I189486,I189469,I529524);
or I_10988 (I189503,I189486,I529509);
DFFARX1 I_10989 (I189503,I2683,I189062,I189529,);
nand I_10990 (I189537,I189529,I189195);
nor I_10991 (I189039,I189537,I189345);
nor I_10992 (I189033,I189529,I189161);
DFFARX1 I_10993 (I189529,I2683,I189062,I189591,);
not I_10994 (I189599,I189591);
nor I_10995 (I189048,I189599,I189311);
not I_10996 (I189657,I2690);
DFFARX1 I_10997 (I354090,I2683,I189657,I189683,);
DFFARX1 I_10998 (I189683,I2683,I189657,I189700,);
not I_10999 (I189649,I189700);
not I_11000 (I189722,I189683);
DFFARX1 I_11001 (I354078,I2683,I189657,I189748,);
not I_11002 (I189756,I189748);
and I_11003 (I189773,I189722,I354087);
not I_11004 (I189790,I354084);
nand I_11005 (I189807,I189790,I354087);
not I_11006 (I189824,I354075);
nor I_11007 (I189841,I189824,I354081);
nand I_11008 (I189858,I189841,I354066);
nor I_11009 (I189875,I189858,I189807);
DFFARX1 I_11010 (I189875,I2683,I189657,I189625,);
not I_11011 (I189906,I189858);
not I_11012 (I189923,I354081);
nand I_11013 (I189940,I189923,I354087);
nor I_11014 (I189957,I354081,I354084);
nand I_11015 (I189637,I189773,I189957);
nand I_11016 (I189631,I189722,I354081);
nand I_11017 (I190002,I189824,I354066);
DFFARX1 I_11018 (I190002,I2683,I189657,I189646,);
DFFARX1 I_11019 (I190002,I2683,I189657,I189640,);
not I_11020 (I190047,I354066);
nor I_11021 (I190064,I190047,I354072);
and I_11022 (I190081,I190064,I354069);
or I_11023 (I190098,I190081,I354093);
DFFARX1 I_11024 (I190098,I2683,I189657,I190124,);
nand I_11025 (I190132,I190124,I189790);
nor I_11026 (I189634,I190132,I189940);
nor I_11027 (I189628,I190124,I189756);
DFFARX1 I_11028 (I190124,I2683,I189657,I190186,);
not I_11029 (I190194,I190186);
nor I_11030 (I189643,I190194,I189906);
not I_11031 (I190252,I2690);
DFFARX1 I_11032 (I435307,I2683,I190252,I190278,);
DFFARX1 I_11033 (I190278,I2683,I190252,I190295,);
not I_11034 (I190244,I190295);
not I_11035 (I190317,I190278);
DFFARX1 I_11036 (I435298,I2683,I190252,I190343,);
not I_11037 (I190351,I190343);
and I_11038 (I190368,I190317,I435316);
not I_11039 (I190385,I435313);
nand I_11040 (I190402,I190385,I435316);
not I_11041 (I190419,I435292);
nor I_11042 (I190436,I190419,I435295);
nand I_11043 (I190453,I190436,I435304);
nor I_11044 (I190470,I190453,I190402);
DFFARX1 I_11045 (I190470,I2683,I190252,I190220,);
not I_11046 (I190501,I190453);
not I_11047 (I190518,I435295);
nand I_11048 (I190535,I190518,I435316);
nor I_11049 (I190552,I435295,I435313);
nand I_11050 (I190232,I190368,I190552);
nand I_11051 (I190226,I190317,I435295);
nand I_11052 (I190597,I190419,I435310);
DFFARX1 I_11053 (I190597,I2683,I190252,I190241,);
DFFARX1 I_11054 (I190597,I2683,I190252,I190235,);
not I_11055 (I190642,I435310);
nor I_11056 (I190659,I190642,I435292);
and I_11057 (I190676,I190659,I435301);
or I_11058 (I190693,I190676,I435295);
DFFARX1 I_11059 (I190693,I2683,I190252,I190719,);
nand I_11060 (I190727,I190719,I190385);
nor I_11061 (I190229,I190727,I190535);
nor I_11062 (I190223,I190719,I190351);
DFFARX1 I_11063 (I190719,I2683,I190252,I190781,);
not I_11064 (I190789,I190781);
nor I_11065 (I190238,I190789,I190501);
not I_11066 (I190847,I2690);
DFFARX1 I_11067 (I877326,I2683,I190847,I190873,);
DFFARX1 I_11068 (I190873,I2683,I190847,I190890,);
not I_11069 (I190839,I190890);
not I_11070 (I190912,I190873);
DFFARX1 I_11071 (I877326,I2683,I190847,I190938,);
not I_11072 (I190946,I190938);
and I_11073 (I190963,I190912,I877329);
not I_11074 (I190980,I877341);
nand I_11075 (I190997,I190980,I877329);
not I_11076 (I191014,I877347);
nor I_11077 (I191031,I191014,I877338);
nand I_11078 (I191048,I191031,I877344);
nor I_11079 (I191065,I191048,I190997);
DFFARX1 I_11080 (I191065,I2683,I190847,I190815,);
not I_11081 (I191096,I191048);
not I_11082 (I191113,I877338);
nand I_11083 (I191130,I191113,I877329);
nor I_11084 (I191147,I877338,I877341);
nand I_11085 (I190827,I190963,I191147);
nand I_11086 (I190821,I190912,I877338);
nand I_11087 (I191192,I191014,I877335);
DFFARX1 I_11088 (I191192,I2683,I190847,I190836,);
DFFARX1 I_11089 (I191192,I2683,I190847,I190830,);
not I_11090 (I191237,I877335);
nor I_11091 (I191254,I191237,I877332);
and I_11092 (I191271,I191254,I877350);
or I_11093 (I191288,I191271,I877329);
DFFARX1 I_11094 (I191288,I2683,I190847,I191314,);
nand I_11095 (I191322,I191314,I190980);
nor I_11096 (I190824,I191322,I191130);
nor I_11097 (I190818,I191314,I190946);
DFFARX1 I_11098 (I191314,I2683,I190847,I191376,);
not I_11099 (I191384,I191376);
nor I_11100 (I190833,I191384,I191096);
not I_11101 (I191442,I2690);
DFFARX1 I_11102 (I289636,I2683,I191442,I191468,);
DFFARX1 I_11103 (I191468,I2683,I191442,I191485,);
not I_11104 (I191434,I191485);
not I_11105 (I191507,I191468);
DFFARX1 I_11106 (I289651,I2683,I191442,I191533,);
not I_11107 (I191541,I191533);
and I_11108 (I191558,I191507,I289648);
not I_11109 (I191575,I289636);
nand I_11110 (I191592,I191575,I289648);
not I_11111 (I191609,I289645);
nor I_11112 (I191626,I191609,I289660);
nand I_11113 (I191643,I191626,I289657);
nor I_11114 (I191660,I191643,I191592);
DFFARX1 I_11115 (I191660,I2683,I191442,I191410,);
not I_11116 (I191691,I191643);
not I_11117 (I191708,I289660);
nand I_11118 (I191725,I191708,I289648);
nor I_11119 (I191742,I289660,I289636);
nand I_11120 (I191422,I191558,I191742);
nand I_11121 (I191416,I191507,I289660);
nand I_11122 (I191787,I191609,I289654);
DFFARX1 I_11123 (I191787,I2683,I191442,I191431,);
DFFARX1 I_11124 (I191787,I2683,I191442,I191425,);
not I_11125 (I191832,I289654);
nor I_11126 (I191849,I191832,I289642);
and I_11127 (I191866,I191849,I289663);
or I_11128 (I191883,I191866,I289639);
DFFARX1 I_11129 (I191883,I2683,I191442,I191909,);
nand I_11130 (I191917,I191909,I191575);
nor I_11131 (I191419,I191917,I191725);
nor I_11132 (I191413,I191909,I191541);
DFFARX1 I_11133 (I191909,I2683,I191442,I191971,);
not I_11134 (I191979,I191971);
nor I_11135 (I191428,I191979,I191691);
not I_11136 (I192037,I2690);
DFFARX1 I_11137 (I791712,I2683,I192037,I192063,);
DFFARX1 I_11138 (I192063,I2683,I192037,I192080,);
not I_11139 (I192029,I192080);
not I_11140 (I192102,I192063);
DFFARX1 I_11141 (I791721,I2683,I192037,I192128,);
not I_11142 (I192136,I192128);
and I_11143 (I192153,I192102,I791709);
not I_11144 (I192170,I791700);
nand I_11145 (I192187,I192170,I791709);
not I_11146 (I192204,I791706);
nor I_11147 (I192221,I192204,I791724);
nand I_11148 (I192238,I192221,I791697);
nor I_11149 (I192255,I192238,I192187);
DFFARX1 I_11150 (I192255,I2683,I192037,I192005,);
not I_11151 (I192286,I192238);
not I_11152 (I192303,I791724);
nand I_11153 (I192320,I192303,I791709);
nor I_11154 (I192337,I791724,I791700);
nand I_11155 (I192017,I192153,I192337);
nand I_11156 (I192011,I192102,I791724);
nand I_11157 (I192382,I192204,I791703);
DFFARX1 I_11158 (I192382,I2683,I192037,I192026,);
DFFARX1 I_11159 (I192382,I2683,I192037,I192020,);
not I_11160 (I192427,I791703);
nor I_11161 (I192444,I192427,I791715);
and I_11162 (I192461,I192444,I791697);
or I_11163 (I192478,I192461,I791718);
DFFARX1 I_11164 (I192478,I2683,I192037,I192504,);
nand I_11165 (I192512,I192504,I192170);
nor I_11166 (I192014,I192512,I192320);
nor I_11167 (I192008,I192504,I192136);
DFFARX1 I_11168 (I192504,I2683,I192037,I192566,);
not I_11169 (I192574,I192566);
nor I_11170 (I192023,I192574,I192286);
not I_11171 (I192632,I2690);
DFFARX1 I_11172 (I1035855,I2683,I192632,I192658,);
DFFARX1 I_11173 (I192658,I2683,I192632,I192675,);
not I_11174 (I192624,I192675);
not I_11175 (I192697,I192658);
DFFARX1 I_11176 (I1035846,I2683,I192632,I192723,);
not I_11177 (I192731,I192723);
and I_11178 (I192748,I192697,I1035840);
not I_11179 (I192765,I1035834);
nand I_11180 (I192782,I192765,I1035840);
not I_11181 (I192799,I1035861);
nor I_11182 (I192816,I192799,I1035834);
nand I_11183 (I192833,I192816,I1035858);
nor I_11184 (I192850,I192833,I192782);
DFFARX1 I_11185 (I192850,I2683,I192632,I192600,);
not I_11186 (I192881,I192833);
not I_11187 (I192898,I1035834);
nand I_11188 (I192915,I192898,I1035840);
nor I_11189 (I192932,I1035834,I1035834);
nand I_11190 (I192612,I192748,I192932);
nand I_11191 (I192606,I192697,I1035834);
nand I_11192 (I192977,I192799,I1035843);
DFFARX1 I_11193 (I192977,I2683,I192632,I192621,);
DFFARX1 I_11194 (I192977,I2683,I192632,I192615,);
not I_11195 (I193022,I1035843);
nor I_11196 (I193039,I193022,I1035849);
and I_11197 (I193056,I193039,I1035852);
or I_11198 (I193073,I193056,I1035837);
DFFARX1 I_11199 (I193073,I2683,I192632,I193099,);
nand I_11200 (I193107,I193099,I192765);
nor I_11201 (I192609,I193107,I192915);
nor I_11202 (I192603,I193099,I192731);
DFFARX1 I_11203 (I193099,I2683,I192632,I193161,);
not I_11204 (I193169,I193161);
nor I_11205 (I192618,I193169,I192881);
not I_11206 (I193227,I2690);
DFFARX1 I_11207 (I214802,I2683,I193227,I193253,);
DFFARX1 I_11208 (I193253,I2683,I193227,I193270,);
not I_11209 (I193219,I193270);
not I_11210 (I193292,I193253);
DFFARX1 I_11211 (I214817,I2683,I193227,I193318,);
not I_11212 (I193326,I193318);
and I_11213 (I193343,I193292,I214814);
not I_11214 (I193360,I214802);
nand I_11215 (I193377,I193360,I214814);
not I_11216 (I193394,I214811);
nor I_11217 (I193411,I193394,I214826);
nand I_11218 (I193428,I193411,I214823);
nor I_11219 (I193445,I193428,I193377);
DFFARX1 I_11220 (I193445,I2683,I193227,I193195,);
not I_11221 (I193476,I193428);
not I_11222 (I193493,I214826);
nand I_11223 (I193510,I193493,I214814);
nor I_11224 (I193527,I214826,I214802);
nand I_11225 (I193207,I193343,I193527);
nand I_11226 (I193201,I193292,I214826);
nand I_11227 (I193572,I193394,I214820);
DFFARX1 I_11228 (I193572,I2683,I193227,I193216,);
DFFARX1 I_11229 (I193572,I2683,I193227,I193210,);
not I_11230 (I193617,I214820);
nor I_11231 (I193634,I193617,I214808);
and I_11232 (I193651,I193634,I214829);
or I_11233 (I193668,I193651,I214805);
DFFARX1 I_11234 (I193668,I2683,I193227,I193694,);
nand I_11235 (I193702,I193694,I193360);
nor I_11236 (I193204,I193702,I193510);
nor I_11237 (I193198,I193694,I193326);
DFFARX1 I_11238 (I193694,I2683,I193227,I193756,);
not I_11239 (I193764,I193756);
nor I_11240 (I193213,I193764,I193476);
not I_11241 (I193822,I2690);
DFFARX1 I_11242 (I1020969,I2683,I193822,I193848,);
DFFARX1 I_11243 (I193848,I2683,I193822,I193865,);
not I_11244 (I193814,I193865);
not I_11245 (I193887,I193848);
DFFARX1 I_11246 (I1020942,I2683,I193822,I193913,);
not I_11247 (I193921,I193913);
and I_11248 (I193938,I193887,I1020966);
not I_11249 (I193955,I1020963);
nand I_11250 (I193972,I193955,I1020966);
not I_11251 (I193989,I1020942);
nor I_11252 (I194006,I193989,I1020960);
nand I_11253 (I194023,I194006,I1020948);
nor I_11254 (I194040,I194023,I193972);
DFFARX1 I_11255 (I194040,I2683,I193822,I193790,);
not I_11256 (I194071,I194023);
not I_11257 (I194088,I1020960);
nand I_11258 (I194105,I194088,I1020966);
nor I_11259 (I194122,I1020960,I1020963);
nand I_11260 (I193802,I193938,I194122);
nand I_11261 (I193796,I193887,I1020960);
nand I_11262 (I194167,I193989,I1020954);
DFFARX1 I_11263 (I194167,I2683,I193822,I193811,);
DFFARX1 I_11264 (I194167,I2683,I193822,I193805,);
not I_11265 (I194212,I1020954);
nor I_11266 (I194229,I194212,I1020957);
and I_11267 (I194246,I194229,I1020945);
or I_11268 (I194263,I194246,I1020951);
DFFARX1 I_11269 (I194263,I2683,I193822,I194289,);
nand I_11270 (I194297,I194289,I193955);
nor I_11271 (I193799,I194297,I194105);
nor I_11272 (I193793,I194289,I193921);
DFFARX1 I_11273 (I194289,I2683,I193822,I194351,);
not I_11274 (I194359,I194351);
nor I_11275 (I193808,I194359,I194071);
not I_11276 (I194417,I2690);
DFFARX1 I_11277 (I738094,I2683,I194417,I194443,);
DFFARX1 I_11278 (I194443,I2683,I194417,I194460,);
not I_11279 (I194409,I194460);
not I_11280 (I194482,I194443);
DFFARX1 I_11281 (I738103,I2683,I194417,I194508,);
not I_11282 (I194516,I194508);
and I_11283 (I194533,I194482,I738091);
not I_11284 (I194550,I738082);
nand I_11285 (I194567,I194550,I738091);
not I_11286 (I194584,I738088);
nor I_11287 (I194601,I194584,I738106);
nand I_11288 (I194618,I194601,I738079);
nor I_11289 (I194635,I194618,I194567);
DFFARX1 I_11290 (I194635,I2683,I194417,I194385,);
not I_11291 (I194666,I194618);
not I_11292 (I194683,I738106);
nand I_11293 (I194700,I194683,I738091);
nor I_11294 (I194717,I738106,I738082);
nand I_11295 (I194397,I194533,I194717);
nand I_11296 (I194391,I194482,I738106);
nand I_11297 (I194762,I194584,I738085);
DFFARX1 I_11298 (I194762,I2683,I194417,I194406,);
DFFARX1 I_11299 (I194762,I2683,I194417,I194400,);
not I_11300 (I194807,I738085);
nor I_11301 (I194824,I194807,I738097);
and I_11302 (I194841,I194824,I738079);
or I_11303 (I194858,I194841,I738100);
DFFARX1 I_11304 (I194858,I2683,I194417,I194884,);
nand I_11305 (I194892,I194884,I194550);
nor I_11306 (I194394,I194892,I194700);
nor I_11307 (I194388,I194884,I194516);
DFFARX1 I_11308 (I194884,I2683,I194417,I194946,);
not I_11309 (I194954,I194946);
nor I_11310 (I194403,I194954,I194666);
not I_11311 (I195012,I2690);
DFFARX1 I_11312 (I994935,I2683,I195012,I195038,);
DFFARX1 I_11313 (I195038,I2683,I195012,I195055,);
not I_11314 (I195004,I195055);
not I_11315 (I195077,I195038);
DFFARX1 I_11316 (I994947,I2683,I195012,I195103,);
not I_11317 (I195111,I195103);
and I_11318 (I195128,I195077,I994941);
not I_11319 (I195145,I994953);
nand I_11320 (I195162,I195145,I994941);
not I_11321 (I195179,I994938);
nor I_11322 (I195196,I195179,I994950);
nand I_11323 (I195213,I195196,I994932);
nor I_11324 (I195230,I195213,I195162);
DFFARX1 I_11325 (I195230,I2683,I195012,I194980,);
not I_11326 (I195261,I195213);
not I_11327 (I195278,I994950);
nand I_11328 (I195295,I195278,I994941);
nor I_11329 (I195312,I994950,I994953);
nand I_11330 (I194992,I195128,I195312);
nand I_11331 (I194986,I195077,I994950);
nand I_11332 (I195357,I195179,I994944);
DFFARX1 I_11333 (I195357,I2683,I195012,I195001,);
DFFARX1 I_11334 (I195357,I2683,I195012,I194995,);
not I_11335 (I195402,I994944);
nor I_11336 (I195419,I195402,I994935);
and I_11337 (I195436,I195419,I994932);
or I_11338 (I195453,I195436,I994956);
DFFARX1 I_11339 (I195453,I2683,I195012,I195479,);
nand I_11340 (I195487,I195479,I195145);
nor I_11341 (I194989,I195487,I195295);
nor I_11342 (I194983,I195479,I195111);
DFFARX1 I_11343 (I195479,I2683,I195012,I195541,);
not I_11344 (I195549,I195541);
nor I_11345 (I194998,I195549,I195261);
not I_11346 (I195607,I2690);
DFFARX1 I_11347 (I365514,I2683,I195607,I195633,);
DFFARX1 I_11348 (I195633,I2683,I195607,I195650,);
not I_11349 (I195599,I195650);
not I_11350 (I195672,I195633);
DFFARX1 I_11351 (I365502,I2683,I195607,I195698,);
not I_11352 (I195706,I195698);
and I_11353 (I195723,I195672,I365511);
not I_11354 (I195740,I365508);
nand I_11355 (I195757,I195740,I365511);
not I_11356 (I195774,I365499);
nor I_11357 (I195791,I195774,I365505);
nand I_11358 (I195808,I195791,I365490);
nor I_11359 (I195825,I195808,I195757);
DFFARX1 I_11360 (I195825,I2683,I195607,I195575,);
not I_11361 (I195856,I195808);
not I_11362 (I195873,I365505);
nand I_11363 (I195890,I195873,I365511);
nor I_11364 (I195907,I365505,I365508);
nand I_11365 (I195587,I195723,I195907);
nand I_11366 (I195581,I195672,I365505);
nand I_11367 (I195952,I195774,I365490);
DFFARX1 I_11368 (I195952,I2683,I195607,I195596,);
DFFARX1 I_11369 (I195952,I2683,I195607,I195590,);
not I_11370 (I195997,I365490);
nor I_11371 (I196014,I195997,I365496);
and I_11372 (I196031,I196014,I365493);
or I_11373 (I196048,I196031,I365517);
DFFARX1 I_11374 (I196048,I2683,I195607,I196074,);
nand I_11375 (I196082,I196074,I195740);
nor I_11376 (I195584,I196082,I195890);
nor I_11377 (I195578,I196074,I195706);
DFFARX1 I_11378 (I196074,I2683,I195607,I196136,);
not I_11379 (I196144,I196136);
nor I_11380 (I195593,I196144,I195856);
not I_11381 (I196202,I2690);
DFFARX1 I_11382 (I2711,I2683,I196202,I196228,);
DFFARX1 I_11383 (I196228,I2683,I196202,I196245,);
not I_11384 (I196194,I196245);
not I_11385 (I196267,I196228);
DFFARX1 I_11386 (I2708,I2683,I196202,I196293,);
not I_11387 (I196301,I196293);
and I_11388 (I196318,I196267,I2699);
not I_11389 (I196335,I2696);
nand I_11390 (I196352,I196335,I2699);
not I_11391 (I196369,I2696);
nor I_11392 (I196386,I196369,I2693);
nand I_11393 (I196403,I196386,I2705);
nor I_11394 (I196420,I196403,I196352);
DFFARX1 I_11395 (I196420,I2683,I196202,I196170,);
not I_11396 (I196451,I196403);
not I_11397 (I196468,I2693);
nand I_11398 (I196485,I196468,I2699);
nor I_11399 (I196502,I2693,I2696);
nand I_11400 (I196182,I196318,I196502);
nand I_11401 (I196176,I196267,I2693);
nand I_11402 (I196547,I196369,I2702);
DFFARX1 I_11403 (I196547,I2683,I196202,I196191,);
DFFARX1 I_11404 (I196547,I2683,I196202,I196185,);
not I_11405 (I196592,I2702);
nor I_11406 (I196609,I196592,I2714);
and I_11407 (I196626,I196609,I2699);
or I_11408 (I196643,I196626,I2693);
DFFARX1 I_11409 (I196643,I2683,I196202,I196669,);
nand I_11410 (I196677,I196669,I196335);
nor I_11411 (I196179,I196677,I196485);
nor I_11412 (I196173,I196669,I196301);
DFFARX1 I_11413 (I196669,I2683,I196202,I196731,);
not I_11414 (I196739,I196731);
nor I_11415 (I196188,I196739,I196451);
not I_11416 (I196797,I2690);
DFFARX1 I_11417 (I670221,I2683,I196797,I196823,);
DFFARX1 I_11418 (I196823,I2683,I196797,I196840,);
not I_11419 (I196789,I196840);
not I_11420 (I196862,I196823);
DFFARX1 I_11421 (I670215,I2683,I196797,I196888,);
not I_11422 (I196896,I196888);
and I_11423 (I196913,I196862,I670233);
not I_11424 (I196930,I670221);
nand I_11425 (I196947,I196930,I670233);
not I_11426 (I196964,I670215);
nor I_11427 (I196981,I196964,I670227);
nand I_11428 (I196998,I196981,I670218);
nor I_11429 (I197015,I196998,I196947);
DFFARX1 I_11430 (I197015,I2683,I196797,I196765,);
not I_11431 (I197046,I196998);
not I_11432 (I197063,I670227);
nand I_11433 (I197080,I197063,I670233);
nor I_11434 (I197097,I670227,I670221);
nand I_11435 (I196777,I196913,I197097);
nand I_11436 (I196771,I196862,I670227);
nand I_11437 (I197142,I196964,I670230);
DFFARX1 I_11438 (I197142,I2683,I196797,I196786,);
DFFARX1 I_11439 (I197142,I2683,I196797,I196780,);
not I_11440 (I197187,I670230);
nor I_11441 (I197204,I197187,I670236);
and I_11442 (I197221,I197204,I670218);
or I_11443 (I197238,I197221,I670224);
DFFARX1 I_11444 (I197238,I2683,I196797,I197264,);
nand I_11445 (I197272,I197264,I196930);
nor I_11446 (I196774,I197272,I197080);
nor I_11447 (I196768,I197264,I196896);
DFFARX1 I_11448 (I197264,I2683,I196797,I197326,);
not I_11449 (I197334,I197326);
nor I_11450 (I196783,I197334,I197046);
not I_11451 (I197392,I2690);
DFFARX1 I_11452 (I514490,I2683,I197392,I197418,);
DFFARX1 I_11453 (I197418,I2683,I197392,I197435,);
not I_11454 (I197384,I197435);
not I_11455 (I197457,I197418);
DFFARX1 I_11456 (I514487,I2683,I197392,I197483,);
not I_11457 (I197491,I197483);
and I_11458 (I197508,I197457,I514493);
not I_11459 (I197525,I514478);
nand I_11460 (I197542,I197525,I514493);
not I_11461 (I197559,I514481);
nor I_11462 (I197576,I197559,I514502);
nand I_11463 (I197593,I197576,I514499);
nor I_11464 (I197610,I197593,I197542);
DFFARX1 I_11465 (I197610,I2683,I197392,I197360,);
not I_11466 (I197641,I197593);
not I_11467 (I197658,I514502);
nand I_11468 (I197675,I197658,I514493);
nor I_11469 (I197692,I514502,I514478);
nand I_11470 (I197372,I197508,I197692);
nand I_11471 (I197366,I197457,I514502);
nand I_11472 (I197737,I197559,I514478);
DFFARX1 I_11473 (I197737,I2683,I197392,I197381,);
DFFARX1 I_11474 (I197737,I2683,I197392,I197375,);
not I_11475 (I197782,I514478);
nor I_11476 (I197799,I197782,I514484);
and I_11477 (I197816,I197799,I514496);
or I_11478 (I197833,I197816,I514481);
DFFARX1 I_11479 (I197833,I2683,I197392,I197859,);
nand I_11480 (I197867,I197859,I197525);
nor I_11481 (I197369,I197867,I197675);
nor I_11482 (I197363,I197859,I197491);
DFFARX1 I_11483 (I197859,I2683,I197392,I197921,);
not I_11484 (I197929,I197921);
nor I_11485 (I197378,I197929,I197641);
not I_11486 (I197987,I2690);
DFFARX1 I_11487 (I264340,I2683,I197987,I198013,);
DFFARX1 I_11488 (I198013,I2683,I197987,I198030,);
not I_11489 (I197979,I198030);
not I_11490 (I198052,I198013);
DFFARX1 I_11491 (I264355,I2683,I197987,I198078,);
not I_11492 (I198086,I198078);
and I_11493 (I198103,I198052,I264352);
not I_11494 (I198120,I264340);
nand I_11495 (I198137,I198120,I264352);
not I_11496 (I198154,I264349);
nor I_11497 (I198171,I198154,I264364);
nand I_11498 (I198188,I198171,I264361);
nor I_11499 (I198205,I198188,I198137);
DFFARX1 I_11500 (I198205,I2683,I197987,I197955,);
not I_11501 (I198236,I198188);
not I_11502 (I198253,I264364);
nand I_11503 (I198270,I198253,I264352);
nor I_11504 (I198287,I264364,I264340);
nand I_11505 (I197967,I198103,I198287);
nand I_11506 (I197961,I198052,I264364);
nand I_11507 (I198332,I198154,I264358);
DFFARX1 I_11508 (I198332,I2683,I197987,I197976,);
DFFARX1 I_11509 (I198332,I2683,I197987,I197970,);
not I_11510 (I198377,I264358);
nor I_11511 (I198394,I198377,I264346);
and I_11512 (I198411,I198394,I264367);
or I_11513 (I198428,I198411,I264343);
DFFARX1 I_11514 (I198428,I2683,I197987,I198454,);
nand I_11515 (I198462,I198454,I198120);
nor I_11516 (I197964,I198462,I198270);
nor I_11517 (I197958,I198454,I198086);
DFFARX1 I_11518 (I198454,I2683,I197987,I198516,);
not I_11519 (I198524,I198516);
nor I_11520 (I197973,I198524,I198236);
not I_11521 (I198582,I2690);
DFFARX1 I_11522 (I1000715,I2683,I198582,I198608,);
DFFARX1 I_11523 (I198608,I2683,I198582,I198625,);
not I_11524 (I198574,I198625);
not I_11525 (I198647,I198608);
DFFARX1 I_11526 (I1000727,I2683,I198582,I198673,);
not I_11527 (I198681,I198673);
and I_11528 (I198698,I198647,I1000721);
not I_11529 (I198715,I1000733);
nand I_11530 (I198732,I198715,I1000721);
not I_11531 (I198749,I1000718);
nor I_11532 (I198766,I198749,I1000730);
nand I_11533 (I198783,I198766,I1000712);
nor I_11534 (I198800,I198783,I198732);
DFFARX1 I_11535 (I198800,I2683,I198582,I198550,);
not I_11536 (I198831,I198783);
not I_11537 (I198848,I1000730);
nand I_11538 (I198865,I198848,I1000721);
nor I_11539 (I198882,I1000730,I1000733);
nand I_11540 (I198562,I198698,I198882);
nand I_11541 (I198556,I198647,I1000730);
nand I_11542 (I198927,I198749,I1000724);
DFFARX1 I_11543 (I198927,I2683,I198582,I198571,);
DFFARX1 I_11544 (I198927,I2683,I198582,I198565,);
not I_11545 (I198972,I1000724);
nor I_11546 (I198989,I198972,I1000715);
and I_11547 (I199006,I198989,I1000712);
or I_11548 (I199023,I199006,I1000736);
DFFARX1 I_11549 (I199023,I2683,I198582,I199049,);
nand I_11550 (I199057,I199049,I198715);
nor I_11551 (I198559,I199057,I198865);
nor I_11552 (I198553,I199049,I198681);
DFFARX1 I_11553 (I199049,I2683,I198582,I199111,);
not I_11554 (I199119,I199111);
nor I_11555 (I198568,I199119,I198831);
not I_11556 (I199177,I2690);
DFFARX1 I_11557 (I304919,I2683,I199177,I199203,);
DFFARX1 I_11558 (I199203,I2683,I199177,I199220,);
not I_11559 (I199169,I199220);
not I_11560 (I199242,I199203);
DFFARX1 I_11561 (I304934,I2683,I199177,I199268,);
not I_11562 (I199276,I199268);
and I_11563 (I199293,I199242,I304931);
not I_11564 (I199310,I304919);
nand I_11565 (I199327,I199310,I304931);
not I_11566 (I199344,I304928);
nor I_11567 (I199361,I199344,I304943);
nand I_11568 (I199378,I199361,I304940);
nor I_11569 (I199395,I199378,I199327);
DFFARX1 I_11570 (I199395,I2683,I199177,I199145,);
not I_11571 (I199426,I199378);
not I_11572 (I199443,I304943);
nand I_11573 (I199460,I199443,I304931);
nor I_11574 (I199477,I304943,I304919);
nand I_11575 (I199157,I199293,I199477);
nand I_11576 (I199151,I199242,I304943);
nand I_11577 (I199522,I199344,I304937);
DFFARX1 I_11578 (I199522,I2683,I199177,I199166,);
DFFARX1 I_11579 (I199522,I2683,I199177,I199160,);
not I_11580 (I199567,I304937);
nor I_11581 (I199584,I199567,I304925);
and I_11582 (I199601,I199584,I304946);
or I_11583 (I199618,I199601,I304922);
DFFARX1 I_11584 (I199618,I2683,I199177,I199644,);
nand I_11585 (I199652,I199644,I199310);
nor I_11586 (I199154,I199652,I199460);
nor I_11587 (I199148,I199644,I199276);
DFFARX1 I_11588 (I199644,I2683,I199177,I199706,);
not I_11589 (I199714,I199706);
nor I_11590 (I199163,I199714,I199426);
not I_11591 (I199772,I2690);
DFFARX1 I_11592 (I684450,I2683,I199772,I199798,);
DFFARX1 I_11593 (I199798,I2683,I199772,I199815,);
not I_11594 (I199764,I199815);
not I_11595 (I199837,I199798);
DFFARX1 I_11596 (I684444,I2683,I199772,I199863,);
not I_11597 (I199871,I199863);
and I_11598 (I199888,I199837,I684462);
not I_11599 (I199905,I684450);
nand I_11600 (I199922,I199905,I684462);
not I_11601 (I199939,I684444);
nor I_11602 (I199956,I199939,I684456);
nand I_11603 (I199973,I199956,I684447);
nor I_11604 (I199990,I199973,I199922);
DFFARX1 I_11605 (I199990,I2683,I199772,I199740,);
not I_11606 (I200021,I199973);
not I_11607 (I200038,I684456);
nand I_11608 (I200055,I200038,I684462);
nor I_11609 (I200072,I684456,I684450);
nand I_11610 (I199752,I199888,I200072);
nand I_11611 (I199746,I199837,I684456);
nand I_11612 (I200117,I199939,I684459);
DFFARX1 I_11613 (I200117,I2683,I199772,I199761,);
DFFARX1 I_11614 (I200117,I2683,I199772,I199755,);
not I_11615 (I200162,I684459);
nor I_11616 (I200179,I200162,I684465);
and I_11617 (I200196,I200179,I684447);
or I_11618 (I200213,I200196,I684453);
DFFARX1 I_11619 (I200213,I2683,I199772,I200239,);
nand I_11620 (I200247,I200239,I199905);
nor I_11621 (I199749,I200247,I200055);
nor I_11622 (I199743,I200239,I199871);
DFFARX1 I_11623 (I200239,I2683,I199772,I200301,);
not I_11624 (I200309,I200301);
nor I_11625 (I199758,I200309,I200021);
not I_11626 (I200367,I2690);
DFFARX1 I_11627 (I241679,I2683,I200367,I200393,);
DFFARX1 I_11628 (I200393,I2683,I200367,I200410,);
not I_11629 (I200359,I200410);
not I_11630 (I200432,I200393);
DFFARX1 I_11631 (I241694,I2683,I200367,I200458,);
not I_11632 (I200466,I200458);
and I_11633 (I200483,I200432,I241691);
not I_11634 (I200500,I241679);
nand I_11635 (I200517,I200500,I241691);
not I_11636 (I200534,I241688);
nor I_11637 (I200551,I200534,I241703);
nand I_11638 (I200568,I200551,I241700);
nor I_11639 (I200585,I200568,I200517);
DFFARX1 I_11640 (I200585,I2683,I200367,I200335,);
not I_11641 (I200616,I200568);
not I_11642 (I200633,I241703);
nand I_11643 (I200650,I200633,I241691);
nor I_11644 (I200667,I241703,I241679);
nand I_11645 (I200347,I200483,I200667);
nand I_11646 (I200341,I200432,I241703);
nand I_11647 (I200712,I200534,I241697);
DFFARX1 I_11648 (I200712,I2683,I200367,I200356,);
DFFARX1 I_11649 (I200712,I2683,I200367,I200350,);
not I_11650 (I200757,I241697);
nor I_11651 (I200774,I200757,I241685);
and I_11652 (I200791,I200774,I241706);
or I_11653 (I200808,I200791,I241682);
DFFARX1 I_11654 (I200808,I2683,I200367,I200834,);
nand I_11655 (I200842,I200834,I200500);
nor I_11656 (I200344,I200842,I200650);
nor I_11657 (I200338,I200834,I200466);
DFFARX1 I_11658 (I200834,I2683,I200367,I200896,);
not I_11659 (I200904,I200896);
nor I_11660 (I200353,I200904,I200616);
not I_11661 (I200962,I2690);
DFFARX1 I_11662 (I66435,I2683,I200962,I200988,);
DFFARX1 I_11663 (I200988,I2683,I200962,I201005,);
not I_11664 (I200954,I201005);
not I_11665 (I201027,I200988);
DFFARX1 I_11666 (I66429,I2683,I200962,I201053,);
not I_11667 (I201061,I201053);
and I_11668 (I201078,I201027,I66426);
not I_11669 (I201095,I66447);
nand I_11670 (I201112,I201095,I66426);
not I_11671 (I201129,I66441);
nor I_11672 (I201146,I201129,I66432);
nand I_11673 (I201163,I201146,I66438);
nor I_11674 (I201180,I201163,I201112);
DFFARX1 I_11675 (I201180,I2683,I200962,I200930,);
not I_11676 (I201211,I201163);
not I_11677 (I201228,I66432);
nand I_11678 (I201245,I201228,I66426);
nor I_11679 (I201262,I66432,I66447);
nand I_11680 (I200942,I201078,I201262);
nand I_11681 (I200936,I201027,I66432);
nand I_11682 (I201307,I201129,I66426);
DFFARX1 I_11683 (I201307,I2683,I200962,I200951,);
DFFARX1 I_11684 (I201307,I2683,I200962,I200945,);
not I_11685 (I201352,I66426);
nor I_11686 (I201369,I201352,I66444);
and I_11687 (I201386,I201369,I66450);
or I_11688 (I201403,I201386,I66429);
DFFARX1 I_11689 (I201403,I2683,I200962,I201429,);
nand I_11690 (I201437,I201429,I201095);
nor I_11691 (I200939,I201437,I201245);
nor I_11692 (I200933,I201429,I201061);
DFFARX1 I_11693 (I201429,I2683,I200962,I201491,);
not I_11694 (I201499,I201491);
nor I_11695 (I200948,I201499,I201211);
not I_11696 (I201557,I2690);
DFFARX1 I_11697 (I511022,I2683,I201557,I201583,);
DFFARX1 I_11698 (I201583,I2683,I201557,I201600,);
not I_11699 (I201549,I201600);
not I_11700 (I201622,I201583);
DFFARX1 I_11701 (I511019,I2683,I201557,I201648,);
not I_11702 (I201656,I201648);
and I_11703 (I201673,I201622,I511025);
not I_11704 (I201690,I511010);
nand I_11705 (I201707,I201690,I511025);
not I_11706 (I201724,I511013);
nor I_11707 (I201741,I201724,I511034);
nand I_11708 (I201758,I201741,I511031);
nor I_11709 (I201775,I201758,I201707);
DFFARX1 I_11710 (I201775,I2683,I201557,I201525,);
not I_11711 (I201806,I201758);
not I_11712 (I201823,I511034);
nand I_11713 (I201840,I201823,I511025);
nor I_11714 (I201857,I511034,I511010);
nand I_11715 (I201537,I201673,I201857);
nand I_11716 (I201531,I201622,I511034);
nand I_11717 (I201902,I201724,I511010);
DFFARX1 I_11718 (I201902,I2683,I201557,I201546,);
DFFARX1 I_11719 (I201902,I2683,I201557,I201540,);
not I_11720 (I201947,I511010);
nor I_11721 (I201964,I201947,I511016);
and I_11722 (I201981,I201964,I511028);
or I_11723 (I201998,I201981,I511013);
DFFARX1 I_11724 (I201998,I2683,I201557,I202024,);
nand I_11725 (I202032,I202024,I201690);
nor I_11726 (I201534,I202032,I201840);
nor I_11727 (I201528,I202024,I201656);
DFFARX1 I_11728 (I202024,I2683,I201557,I202086,);
not I_11729 (I202094,I202086);
nor I_11730 (I201543,I202094,I201806);
not I_11731 (I202152,I2690);
DFFARX1 I_11732 (I350282,I2683,I202152,I202178,);
DFFARX1 I_11733 (I202178,I2683,I202152,I202195,);
not I_11734 (I202144,I202195);
not I_11735 (I202217,I202178);
DFFARX1 I_11736 (I350270,I2683,I202152,I202243,);
not I_11737 (I202251,I202243);
and I_11738 (I202268,I202217,I350279);
not I_11739 (I202285,I350276);
nand I_11740 (I202302,I202285,I350279);
not I_11741 (I202319,I350267);
nor I_11742 (I202336,I202319,I350273);
nand I_11743 (I202353,I202336,I350258);
nor I_11744 (I202370,I202353,I202302);
DFFARX1 I_11745 (I202370,I2683,I202152,I202120,);
not I_11746 (I202401,I202353);
not I_11747 (I202418,I350273);
nand I_11748 (I202435,I202418,I350279);
nor I_11749 (I202452,I350273,I350276);
nand I_11750 (I202132,I202268,I202452);
nand I_11751 (I202126,I202217,I350273);
nand I_11752 (I202497,I202319,I350258);
DFFARX1 I_11753 (I202497,I2683,I202152,I202141,);
DFFARX1 I_11754 (I202497,I2683,I202152,I202135,);
not I_11755 (I202542,I350258);
nor I_11756 (I202559,I202542,I350264);
and I_11757 (I202576,I202559,I350261);
or I_11758 (I202593,I202576,I350285);
DFFARX1 I_11759 (I202593,I2683,I202152,I202619,);
nand I_11760 (I202627,I202619,I202285);
nor I_11761 (I202129,I202627,I202435);
nor I_11762 (I202123,I202619,I202251);
DFFARX1 I_11763 (I202619,I2683,I202152,I202681,);
not I_11764 (I202689,I202681);
nor I_11765 (I202138,I202689,I202401);
not I_11766 (I202747,I2690);
DFFARX1 I_11767 (I333418,I2683,I202747,I202773,);
DFFARX1 I_11768 (I202773,I2683,I202747,I202790,);
not I_11769 (I202739,I202790);
not I_11770 (I202812,I202773);
DFFARX1 I_11771 (I333406,I2683,I202747,I202838,);
not I_11772 (I202846,I202838);
and I_11773 (I202863,I202812,I333415);
not I_11774 (I202880,I333412);
nand I_11775 (I202897,I202880,I333415);
not I_11776 (I202914,I333403);
nor I_11777 (I202931,I202914,I333409);
nand I_11778 (I202948,I202931,I333394);
nor I_11779 (I202965,I202948,I202897);
DFFARX1 I_11780 (I202965,I2683,I202747,I202715,);
not I_11781 (I202996,I202948);
not I_11782 (I203013,I333409);
nand I_11783 (I203030,I203013,I333415);
nor I_11784 (I203047,I333409,I333412);
nand I_11785 (I202727,I202863,I203047);
nand I_11786 (I202721,I202812,I333409);
nand I_11787 (I203092,I202914,I333394);
DFFARX1 I_11788 (I203092,I2683,I202747,I202736,);
DFFARX1 I_11789 (I203092,I2683,I202747,I202730,);
not I_11790 (I203137,I333394);
nor I_11791 (I203154,I203137,I333400);
and I_11792 (I203171,I203154,I333397);
or I_11793 (I203188,I203171,I333421);
DFFARX1 I_11794 (I203188,I2683,I202747,I203214,);
nand I_11795 (I203222,I203214,I202880);
nor I_11796 (I202724,I203222,I203030);
nor I_11797 (I202718,I203214,I202846);
DFFARX1 I_11798 (I203214,I2683,I202747,I203276,);
not I_11799 (I203284,I203276);
nor I_11800 (I202733,I203284,I202996);
not I_11801 (I203342,I2690);
DFFARX1 I_11802 (I120028,I2683,I203342,I203368,);
DFFARX1 I_11803 (I203368,I2683,I203342,I203385,);
not I_11804 (I203334,I203385);
not I_11805 (I203407,I203368);
DFFARX1 I_11806 (I120013,I2683,I203342,I203433,);
not I_11807 (I203441,I203433);
and I_11808 (I203458,I203407,I120034);
not I_11809 (I203475,I120025);
nand I_11810 (I203492,I203475,I120034);
not I_11811 (I203509,I120010);
nor I_11812 (I203526,I203509,I120022);
nand I_11813 (I203543,I203526,I120037);
nor I_11814 (I203560,I203543,I203492);
DFFARX1 I_11815 (I203560,I2683,I203342,I203310,);
not I_11816 (I203591,I203543);
not I_11817 (I203608,I120022);
nand I_11818 (I203625,I203608,I120034);
nor I_11819 (I203642,I120022,I120025);
nand I_11820 (I203322,I203458,I203642);
nand I_11821 (I203316,I203407,I120022);
nand I_11822 (I203687,I203509,I120016);
DFFARX1 I_11823 (I203687,I2683,I203342,I203331,);
DFFARX1 I_11824 (I203687,I2683,I203342,I203325,);
not I_11825 (I203732,I120016);
nor I_11826 (I203749,I203732,I120019);
and I_11827 (I203766,I203749,I120010);
or I_11828 (I203783,I203766,I120031);
DFFARX1 I_11829 (I203783,I2683,I203342,I203809,);
nand I_11830 (I203817,I203809,I203475);
nor I_11831 (I203319,I203817,I203625);
nor I_11832 (I203313,I203809,I203441);
DFFARX1 I_11833 (I203809,I2683,I203342,I203871,);
not I_11834 (I203879,I203871);
nor I_11835 (I203328,I203879,I203591);
not I_11836 (I203937,I2690);
DFFARX1 I_11837 (I495419,I2683,I203937,I203963,);
DFFARX1 I_11838 (I203963,I2683,I203937,I203980,);
not I_11839 (I203929,I203980);
not I_11840 (I204002,I203963);
DFFARX1 I_11841 (I495410,I2683,I203937,I204028,);
not I_11842 (I204036,I204028);
and I_11843 (I204053,I204002,I495428);
not I_11844 (I204070,I495425);
nand I_11845 (I204087,I204070,I495428);
not I_11846 (I204104,I495404);
nor I_11847 (I204121,I204104,I495407);
nand I_11848 (I204138,I204121,I495416);
nor I_11849 (I204155,I204138,I204087);
DFFARX1 I_11850 (I204155,I2683,I203937,I203905,);
not I_11851 (I204186,I204138);
not I_11852 (I204203,I495407);
nand I_11853 (I204220,I204203,I495428);
nor I_11854 (I204237,I495407,I495425);
nand I_11855 (I203917,I204053,I204237);
nand I_11856 (I203911,I204002,I495407);
nand I_11857 (I204282,I204104,I495422);
DFFARX1 I_11858 (I204282,I2683,I203937,I203926,);
DFFARX1 I_11859 (I204282,I2683,I203937,I203920,);
not I_11860 (I204327,I495422);
nor I_11861 (I204344,I204327,I495404);
and I_11862 (I204361,I204344,I495413);
or I_11863 (I204378,I204361,I495407);
DFFARX1 I_11864 (I204378,I2683,I203937,I204404,);
nand I_11865 (I204412,I204404,I204070);
nor I_11866 (I203914,I204412,I204220);
nor I_11867 (I203908,I204404,I204036);
DFFARX1 I_11868 (I204404,I2683,I203937,I204466,);
not I_11869 (I204474,I204466);
nor I_11870 (I203923,I204474,I204186);
not I_11871 (I204532,I2690);
DFFARX1 I_11872 (I264867,I2683,I204532,I204558,);
DFFARX1 I_11873 (I204558,I2683,I204532,I204575,);
not I_11874 (I204524,I204575);
not I_11875 (I204597,I204558);
DFFARX1 I_11876 (I264882,I2683,I204532,I204623,);
not I_11877 (I204631,I204623);
and I_11878 (I204648,I204597,I264879);
not I_11879 (I204665,I264867);
nand I_11880 (I204682,I204665,I264879);
not I_11881 (I204699,I264876);
nor I_11882 (I204716,I204699,I264891);
nand I_11883 (I204733,I204716,I264888);
nor I_11884 (I204750,I204733,I204682);
DFFARX1 I_11885 (I204750,I2683,I204532,I204500,);
not I_11886 (I204781,I204733);
not I_11887 (I204798,I264891);
nand I_11888 (I204815,I204798,I264879);
nor I_11889 (I204832,I264891,I264867);
nand I_11890 (I204512,I204648,I204832);
nand I_11891 (I204506,I204597,I264891);
nand I_11892 (I204877,I204699,I264885);
DFFARX1 I_11893 (I204877,I2683,I204532,I204521,);
DFFARX1 I_11894 (I204877,I2683,I204532,I204515,);
not I_11895 (I204922,I264885);
nor I_11896 (I204939,I204922,I264873);
and I_11897 (I204956,I204939,I264894);
or I_11898 (I204973,I204956,I264870);
DFFARX1 I_11899 (I204973,I2683,I204532,I204999,);
nand I_11900 (I205007,I204999,I204665);
nor I_11901 (I204509,I205007,I204815);
nor I_11902 (I204503,I204999,I204631);
DFFARX1 I_11903 (I204999,I2683,I204532,I205061,);
not I_11904 (I205069,I205061);
nor I_11905 (I204518,I205069,I204781);
not I_11906 (I205127,I2690);
DFFARX1 I_11907 (I310716,I2683,I205127,I205153,);
DFFARX1 I_11908 (I205153,I2683,I205127,I205170,);
not I_11909 (I205119,I205170);
not I_11910 (I205192,I205153);
DFFARX1 I_11911 (I310731,I2683,I205127,I205218,);
not I_11912 (I205226,I205218);
and I_11913 (I205243,I205192,I310728);
not I_11914 (I205260,I310716);
nand I_11915 (I205277,I205260,I310728);
not I_11916 (I205294,I310725);
nor I_11917 (I205311,I205294,I310740);
nand I_11918 (I205328,I205311,I310737);
nor I_11919 (I205345,I205328,I205277);
DFFARX1 I_11920 (I205345,I2683,I205127,I205095,);
not I_11921 (I205376,I205328);
not I_11922 (I205393,I310740);
nand I_11923 (I205410,I205393,I310728);
nor I_11924 (I205427,I310740,I310716);
nand I_11925 (I205107,I205243,I205427);
nand I_11926 (I205101,I205192,I310740);
nand I_11927 (I205472,I205294,I310734);
DFFARX1 I_11928 (I205472,I2683,I205127,I205116,);
DFFARX1 I_11929 (I205472,I2683,I205127,I205110,);
not I_11930 (I205517,I310734);
nor I_11931 (I205534,I205517,I310722);
and I_11932 (I205551,I205534,I310743);
or I_11933 (I205568,I205551,I310719);
DFFARX1 I_11934 (I205568,I2683,I205127,I205594,);
nand I_11935 (I205602,I205594,I205260);
nor I_11936 (I205104,I205602,I205410);
nor I_11937 (I205098,I205594,I205226);
DFFARX1 I_11938 (I205594,I2683,I205127,I205656,);
not I_11939 (I205664,I205656);
nor I_11940 (I205113,I205664,I205376);
not I_11941 (I205722,I2690);
DFFARX1 I_11942 (I281204,I2683,I205722,I205748,);
DFFARX1 I_11943 (I205748,I2683,I205722,I205765,);
not I_11944 (I205714,I205765);
not I_11945 (I205787,I205748);
DFFARX1 I_11946 (I281219,I2683,I205722,I205813,);
not I_11947 (I205821,I205813);
and I_11948 (I205838,I205787,I281216);
not I_11949 (I205855,I281204);
nand I_11950 (I205872,I205855,I281216);
not I_11951 (I205889,I281213);
nor I_11952 (I205906,I205889,I281228);
nand I_11953 (I205923,I205906,I281225);
nor I_11954 (I205940,I205923,I205872);
DFFARX1 I_11955 (I205940,I2683,I205722,I205690,);
not I_11956 (I205971,I205923);
not I_11957 (I205988,I281228);
nand I_11958 (I206005,I205988,I281216);
nor I_11959 (I206022,I281228,I281204);
nand I_11960 (I205702,I205838,I206022);
nand I_11961 (I205696,I205787,I281228);
nand I_11962 (I206067,I205889,I281222);
DFFARX1 I_11963 (I206067,I2683,I205722,I205711,);
DFFARX1 I_11964 (I206067,I2683,I205722,I205705,);
not I_11965 (I206112,I281222);
nor I_11966 (I206129,I206112,I281210);
and I_11967 (I206146,I206129,I281231);
or I_11968 (I206163,I206146,I281207);
DFFARX1 I_11969 (I206163,I2683,I205722,I206189,);
nand I_11970 (I206197,I206189,I205855);
nor I_11971 (I205699,I206197,I206005);
nor I_11972 (I205693,I206189,I205821);
DFFARX1 I_11973 (I206189,I2683,I205722,I206251,);
not I_11974 (I206259,I206251);
nor I_11975 (I205708,I206259,I205971);
not I_11976 (I206317,I2690);
DFFARX1 I_11977 (I880216,I2683,I206317,I206343,);
DFFARX1 I_11978 (I206343,I2683,I206317,I206360,);
not I_11979 (I206309,I206360);
not I_11980 (I206382,I206343);
DFFARX1 I_11981 (I880216,I2683,I206317,I206408,);
not I_11982 (I206416,I206408);
and I_11983 (I206433,I206382,I880219);
not I_11984 (I206450,I880231);
nand I_11985 (I206467,I206450,I880219);
not I_11986 (I206484,I880237);
nor I_11987 (I206501,I206484,I880228);
nand I_11988 (I206518,I206501,I880234);
nor I_11989 (I206535,I206518,I206467);
DFFARX1 I_11990 (I206535,I2683,I206317,I206285,);
not I_11991 (I206566,I206518);
not I_11992 (I206583,I880228);
nand I_11993 (I206600,I206583,I880219);
nor I_11994 (I206617,I880228,I880231);
nand I_11995 (I206297,I206433,I206617);
nand I_11996 (I206291,I206382,I880228);
nand I_11997 (I206662,I206484,I880225);
DFFARX1 I_11998 (I206662,I2683,I206317,I206306,);
DFFARX1 I_11999 (I206662,I2683,I206317,I206300,);
not I_12000 (I206707,I880225);
nor I_12001 (I206724,I206707,I880222);
and I_12002 (I206741,I206724,I880240);
or I_12003 (I206758,I206741,I880219);
DFFARX1 I_12004 (I206758,I2683,I206317,I206784,);
nand I_12005 (I206792,I206784,I206450);
nor I_12006 (I206294,I206792,I206600);
nor I_12007 (I206288,I206784,I206416);
DFFARX1 I_12008 (I206784,I2683,I206317,I206846,);
not I_12009 (I206854,I206846);
nor I_12010 (I206303,I206854,I206566);
not I_12011 (I206912,I2690);
DFFARX1 I_12012 (I754890,I2683,I206912,I206938,);
DFFARX1 I_12013 (I206938,I2683,I206912,I206955,);
not I_12014 (I206904,I206955);
not I_12015 (I206977,I206938);
DFFARX1 I_12016 (I754899,I2683,I206912,I207003,);
not I_12017 (I207011,I207003);
and I_12018 (I207028,I206977,I754887);
not I_12019 (I207045,I754878);
nand I_12020 (I207062,I207045,I754887);
not I_12021 (I207079,I754884);
nor I_12022 (I207096,I207079,I754902);
nand I_12023 (I207113,I207096,I754875);
nor I_12024 (I207130,I207113,I207062);
DFFARX1 I_12025 (I207130,I2683,I206912,I206880,);
not I_12026 (I207161,I207113);
not I_12027 (I207178,I754902);
nand I_12028 (I207195,I207178,I754887);
nor I_12029 (I207212,I754902,I754878);
nand I_12030 (I206892,I207028,I207212);
nand I_12031 (I206886,I206977,I754902);
nand I_12032 (I207257,I207079,I754881);
DFFARX1 I_12033 (I207257,I2683,I206912,I206901,);
DFFARX1 I_12034 (I207257,I2683,I206912,I206895,);
not I_12035 (I207302,I754881);
nor I_12036 (I207319,I207302,I754893);
and I_12037 (I207336,I207319,I754875);
or I_12038 (I207353,I207336,I754896);
DFFARX1 I_12039 (I207353,I2683,I206912,I207379,);
nand I_12040 (I207387,I207379,I207045);
nor I_12041 (I206889,I207387,I207195);
nor I_12042 (I206883,I207379,I207011);
DFFARX1 I_12043 (I207379,I2683,I206912,I207441,);
not I_12044 (I207449,I207441);
nor I_12045 (I206898,I207449,I207161);
not I_12046 (I207507,I2690);
DFFARX1 I_12047 (I671275,I2683,I207507,I207533,);
DFFARX1 I_12048 (I207533,I2683,I207507,I207550,);
not I_12049 (I207499,I207550);
not I_12050 (I207572,I207533);
DFFARX1 I_12051 (I671269,I2683,I207507,I207598,);
not I_12052 (I207606,I207598);
and I_12053 (I207623,I207572,I671287);
not I_12054 (I207640,I671275);
nand I_12055 (I207657,I207640,I671287);
not I_12056 (I207674,I671269);
nor I_12057 (I207691,I207674,I671281);
nand I_12058 (I207708,I207691,I671272);
nor I_12059 (I207725,I207708,I207657);
DFFARX1 I_12060 (I207725,I2683,I207507,I207475,);
not I_12061 (I207756,I207708);
not I_12062 (I207773,I671281);
nand I_12063 (I207790,I207773,I671287);
nor I_12064 (I207807,I671281,I671275);
nand I_12065 (I207487,I207623,I207807);
nand I_12066 (I207481,I207572,I671281);
nand I_12067 (I207852,I207674,I671284);
DFFARX1 I_12068 (I207852,I2683,I207507,I207496,);
DFFARX1 I_12069 (I207852,I2683,I207507,I207490,);
not I_12070 (I207897,I671284);
nor I_12071 (I207914,I207897,I671290);
and I_12072 (I207931,I207914,I671272);
or I_12073 (I207948,I207931,I671278);
DFFARX1 I_12074 (I207948,I2683,I207507,I207974,);
nand I_12075 (I207982,I207974,I207640);
nor I_12076 (I207484,I207982,I207790);
nor I_12077 (I207478,I207974,I207606);
DFFARX1 I_12078 (I207974,I2683,I207507,I208036,);
not I_12079 (I208044,I208036);
nor I_12080 (I207493,I208044,I207756);
not I_12081 (I208102,I2690);
DFFARX1 I_12082 (I916630,I2683,I208102,I208128,);
DFFARX1 I_12083 (I208128,I2683,I208102,I208145,);
not I_12084 (I208094,I208145);
not I_12085 (I208167,I208128);
DFFARX1 I_12086 (I916630,I2683,I208102,I208193,);
not I_12087 (I208201,I208193);
and I_12088 (I208218,I208167,I916633);
not I_12089 (I208235,I916645);
nand I_12090 (I208252,I208235,I916633);
not I_12091 (I208269,I916651);
nor I_12092 (I208286,I208269,I916642);
nand I_12093 (I208303,I208286,I916648);
nor I_12094 (I208320,I208303,I208252);
DFFARX1 I_12095 (I208320,I2683,I208102,I208070,);
not I_12096 (I208351,I208303);
not I_12097 (I208368,I916642);
nand I_12098 (I208385,I208368,I916633);
nor I_12099 (I208402,I916642,I916645);
nand I_12100 (I208082,I208218,I208402);
nand I_12101 (I208076,I208167,I916642);
nand I_12102 (I208447,I208269,I916639);
DFFARX1 I_12103 (I208447,I2683,I208102,I208091,);
DFFARX1 I_12104 (I208447,I2683,I208102,I208085,);
not I_12105 (I208492,I916639);
nor I_12106 (I208509,I208492,I916636);
and I_12107 (I208526,I208509,I916654);
or I_12108 (I208543,I208526,I916633);
DFFARX1 I_12109 (I208543,I2683,I208102,I208569,);
nand I_12110 (I208577,I208569,I208235);
nor I_12111 (I208079,I208577,I208385);
nor I_12112 (I208073,I208569,I208201);
DFFARX1 I_12113 (I208569,I2683,I208102,I208631,);
not I_12114 (I208639,I208631);
nor I_12115 (I208088,I208639,I208351);
not I_12116 (I208697,I2690);
DFFARX1 I_12117 (I1012275,I2683,I208697,I208723,);
DFFARX1 I_12118 (I208723,I2683,I208697,I208740,);
not I_12119 (I208689,I208740);
not I_12120 (I208762,I208723);
DFFARX1 I_12121 (I1012287,I2683,I208697,I208788,);
not I_12122 (I208796,I208788);
and I_12123 (I208813,I208762,I1012281);
not I_12124 (I208830,I1012293);
nand I_12125 (I208847,I208830,I1012281);
not I_12126 (I208864,I1012278);
nor I_12127 (I208881,I208864,I1012290);
nand I_12128 (I208898,I208881,I1012272);
nor I_12129 (I208915,I208898,I208847);
DFFARX1 I_12130 (I208915,I2683,I208697,I208665,);
not I_12131 (I208946,I208898);
not I_12132 (I208963,I1012290);
nand I_12133 (I208980,I208963,I1012281);
nor I_12134 (I208997,I1012290,I1012293);
nand I_12135 (I208677,I208813,I208997);
nand I_12136 (I208671,I208762,I1012290);
nand I_12137 (I209042,I208864,I1012284);
DFFARX1 I_12138 (I209042,I2683,I208697,I208686,);
DFFARX1 I_12139 (I209042,I2683,I208697,I208680,);
not I_12140 (I209087,I1012284);
nor I_12141 (I209104,I209087,I1012275);
and I_12142 (I209121,I209104,I1012272);
or I_12143 (I209138,I209121,I1012296);
DFFARX1 I_12144 (I209138,I2683,I208697,I209164,);
nand I_12145 (I209172,I209164,I208830);
nor I_12146 (I208674,I209172,I208980);
nor I_12147 (I208668,I209164,I208796);
DFFARX1 I_12148 (I209164,I2683,I208697,I209226,);
not I_12149 (I209234,I209226);
nor I_12150 (I208683,I209234,I208946);
not I_12151 (I209292,I2690);
DFFARX1 I_12152 (I474033,I2683,I209292,I209318,);
DFFARX1 I_12153 (I209318,I2683,I209292,I209335,);
not I_12154 (I209284,I209335);
not I_12155 (I209357,I209318);
DFFARX1 I_12156 (I474024,I2683,I209292,I209383,);
not I_12157 (I209391,I209383);
and I_12158 (I209408,I209357,I474042);
not I_12159 (I209425,I474039);
nand I_12160 (I209442,I209425,I474042);
not I_12161 (I209459,I474018);
nor I_12162 (I209476,I209459,I474021);
nand I_12163 (I209493,I209476,I474030);
nor I_12164 (I209510,I209493,I209442);
DFFARX1 I_12165 (I209510,I2683,I209292,I209260,);
not I_12166 (I209541,I209493);
not I_12167 (I209558,I474021);
nand I_12168 (I209575,I209558,I474042);
nor I_12169 (I209592,I474021,I474039);
nand I_12170 (I209272,I209408,I209592);
nand I_12171 (I209266,I209357,I474021);
nand I_12172 (I209637,I209459,I474036);
DFFARX1 I_12173 (I209637,I2683,I209292,I209281,);
DFFARX1 I_12174 (I209637,I2683,I209292,I209275,);
not I_12175 (I209682,I474036);
nor I_12176 (I209699,I209682,I474018);
and I_12177 (I209716,I209699,I474027);
or I_12178 (I209733,I209716,I474021);
DFFARX1 I_12179 (I209733,I2683,I209292,I209759,);
nand I_12180 (I209767,I209759,I209425);
nor I_12181 (I209269,I209767,I209575);
nor I_12182 (I209263,I209759,I209391);
DFFARX1 I_12183 (I209759,I2683,I209292,I209821,);
not I_12184 (I209829,I209821);
nor I_12185 (I209278,I209829,I209541);
not I_12186 (I209887,I2690);
DFFARX1 I_12187 (I847848,I2683,I209887,I209913,);
DFFARX1 I_12188 (I209913,I2683,I209887,I209930,);
not I_12189 (I209879,I209930);
not I_12190 (I209952,I209913);
DFFARX1 I_12191 (I847848,I2683,I209887,I209978,);
not I_12192 (I209986,I209978);
and I_12193 (I210003,I209952,I847851);
not I_12194 (I210020,I847863);
nand I_12195 (I210037,I210020,I847851);
not I_12196 (I210054,I847869);
nor I_12197 (I210071,I210054,I847860);
nand I_12198 (I210088,I210071,I847866);
nor I_12199 (I210105,I210088,I210037);
DFFARX1 I_12200 (I210105,I2683,I209887,I209855,);
not I_12201 (I210136,I210088);
not I_12202 (I210153,I847860);
nand I_12203 (I210170,I210153,I847851);
nor I_12204 (I210187,I847860,I847863);
nand I_12205 (I209867,I210003,I210187);
nand I_12206 (I209861,I209952,I847860);
nand I_12207 (I210232,I210054,I847857);
DFFARX1 I_12208 (I210232,I2683,I209887,I209876,);
DFFARX1 I_12209 (I210232,I2683,I209887,I209870,);
not I_12210 (I210277,I847857);
nor I_12211 (I210294,I210277,I847854);
and I_12212 (I210311,I210294,I847872);
or I_12213 (I210328,I210311,I847851);
DFFARX1 I_12214 (I210328,I2683,I209887,I210354,);
nand I_12215 (I210362,I210354,I210020);
nor I_12216 (I209864,I210362,I210170);
nor I_12217 (I209858,I210354,I209986);
DFFARX1 I_12218 (I210354,I2683,I209887,I210416,);
not I_12219 (I210424,I210416);
nor I_12220 (I209873,I210424,I210136);
not I_12221 (I210482,I2690);
DFFARX1 I_12222 (I380746,I2683,I210482,I210508,);
DFFARX1 I_12223 (I210508,I2683,I210482,I210525,);
not I_12224 (I210474,I210525);
not I_12225 (I210547,I210508);
DFFARX1 I_12226 (I380734,I2683,I210482,I210573,);
not I_12227 (I210581,I210573);
and I_12228 (I210598,I210547,I380743);
not I_12229 (I210615,I380740);
nand I_12230 (I210632,I210615,I380743);
not I_12231 (I210649,I380731);
nor I_12232 (I210666,I210649,I380737);
nand I_12233 (I210683,I210666,I380722);
nor I_12234 (I210700,I210683,I210632);
DFFARX1 I_12235 (I210700,I2683,I210482,I210450,);
not I_12236 (I210731,I210683);
not I_12237 (I210748,I380737);
nand I_12238 (I210765,I210748,I380743);
nor I_12239 (I210782,I380737,I380740);
nand I_12240 (I210462,I210598,I210782);
nand I_12241 (I210456,I210547,I380737);
nand I_12242 (I210827,I210649,I380722);
DFFARX1 I_12243 (I210827,I2683,I210482,I210471,);
DFFARX1 I_12244 (I210827,I2683,I210482,I210465,);
not I_12245 (I210872,I380722);
nor I_12246 (I210889,I210872,I380728);
and I_12247 (I210906,I210889,I380725);
or I_12248 (I210923,I210906,I380749);
DFFARX1 I_12249 (I210923,I2683,I210482,I210949,);
nand I_12250 (I210957,I210949,I210615);
nor I_12251 (I210459,I210957,I210765);
nor I_12252 (I210453,I210949,I210581);
DFFARX1 I_12253 (I210949,I2683,I210482,I211011,);
not I_12254 (I211019,I211011);
nor I_12255 (I210468,I211019,I210731);
not I_12256 (I211077,I2690);
DFFARX1 I_12257 (I651249,I2683,I211077,I211103,);
DFFARX1 I_12258 (I211103,I2683,I211077,I211120,);
not I_12259 (I211069,I211120);
not I_12260 (I211142,I211103);
DFFARX1 I_12261 (I651243,I2683,I211077,I211168,);
not I_12262 (I211176,I211168);
and I_12263 (I211193,I211142,I651261);
not I_12264 (I211210,I651249);
nand I_12265 (I211227,I211210,I651261);
not I_12266 (I211244,I651243);
nor I_12267 (I211261,I211244,I651255);
nand I_12268 (I211278,I211261,I651246);
nor I_12269 (I211295,I211278,I211227);
DFFARX1 I_12270 (I211295,I2683,I211077,I211045,);
not I_12271 (I211326,I211278);
not I_12272 (I211343,I651255);
nand I_12273 (I211360,I211343,I651261);
nor I_12274 (I211377,I651255,I651249);
nand I_12275 (I211057,I211193,I211377);
nand I_12276 (I211051,I211142,I651255);
nand I_12277 (I211422,I211244,I651258);
DFFARX1 I_12278 (I211422,I2683,I211077,I211066,);
DFFARX1 I_12279 (I211422,I2683,I211077,I211060,);
not I_12280 (I211467,I651258);
nor I_12281 (I211484,I211467,I651264);
and I_12282 (I211501,I211484,I651246);
or I_12283 (I211518,I211501,I651252);
DFFARX1 I_12284 (I211518,I2683,I211077,I211544,);
nand I_12285 (I211552,I211544,I211210);
nor I_12286 (I211054,I211552,I211360);
nor I_12287 (I211048,I211544,I211176);
DFFARX1 I_12288 (I211544,I2683,I211077,I211606,);
not I_12289 (I211614,I211606);
nor I_12290 (I211063,I211614,I211326);
not I_12291 (I211675,I2690);
DFFARX1 I_12292 (I506398,I2683,I211675,I211701,);
nand I_12293 (I211709,I506389,I506404);
and I_12294 (I211726,I211709,I506410);
DFFARX1 I_12295 (I211726,I2683,I211675,I211752,);
nor I_12296 (I211643,I211752,I211701);
not I_12297 (I211774,I211752);
DFFARX1 I_12298 (I506395,I2683,I211675,I211800,);
nand I_12299 (I211808,I211800,I506389);
not I_12300 (I211825,I211808);
DFFARX1 I_12301 (I211825,I2683,I211675,I211851,);
not I_12302 (I211667,I211851);
nor I_12303 (I211873,I211701,I211808);
nor I_12304 (I211649,I211752,I211873);
DFFARX1 I_12305 (I506392,I2683,I211675,I211913,);
DFFARX1 I_12306 (I211913,I2683,I211675,I211930,);
not I_12307 (I211938,I211930);
not I_12308 (I211955,I211913);
nand I_12309 (I211652,I211955,I211774);
nand I_12310 (I211986,I506386,I506401);
and I_12311 (I212003,I211986,I506386);
DFFARX1 I_12312 (I212003,I2683,I211675,I212029,);
nor I_12313 (I212037,I212029,I211701);
DFFARX1 I_12314 (I212037,I2683,I211675,I211640,);
DFFARX1 I_12315 (I212029,I2683,I211675,I211658,);
nor I_12316 (I212082,I506407,I506401);
not I_12317 (I212099,I212082);
nor I_12318 (I211661,I211938,I212099);
nand I_12319 (I211646,I211955,I212099);
nor I_12320 (I211655,I211701,I212082);
DFFARX1 I_12321 (I212082,I2683,I211675,I211664,);
not I_12322 (I212202,I2690);
DFFARX1 I_12323 (I666002,I2683,I212202,I212228,);
nand I_12324 (I212236,I666005,I665999);
and I_12325 (I212253,I212236,I666011);
DFFARX1 I_12326 (I212253,I2683,I212202,I212279,);
nor I_12327 (I212170,I212279,I212228);
not I_12328 (I212301,I212279);
DFFARX1 I_12329 (I666014,I2683,I212202,I212327,);
nand I_12330 (I212335,I212327,I666005);
not I_12331 (I212352,I212335);
DFFARX1 I_12332 (I212352,I2683,I212202,I212378,);
not I_12333 (I212194,I212378);
nor I_12334 (I212400,I212228,I212335);
nor I_12335 (I212176,I212279,I212400);
DFFARX1 I_12336 (I666017,I2683,I212202,I212440,);
DFFARX1 I_12337 (I212440,I2683,I212202,I212457,);
not I_12338 (I212465,I212457);
not I_12339 (I212482,I212440);
nand I_12340 (I212179,I212482,I212301);
nand I_12341 (I212513,I665999,I666008);
and I_12342 (I212530,I212513,I666002);
DFFARX1 I_12343 (I212530,I2683,I212202,I212556,);
nor I_12344 (I212564,I212556,I212228);
DFFARX1 I_12345 (I212564,I2683,I212202,I212167,);
DFFARX1 I_12346 (I212556,I2683,I212202,I212185,);
nor I_12347 (I212609,I666020,I666008);
not I_12348 (I212626,I212609);
nor I_12349 (I212188,I212465,I212626);
nand I_12350 (I212173,I212482,I212626);
nor I_12351 (I212182,I212228,I212609);
DFFARX1 I_12352 (I212609,I2683,I212202,I212191,);
not I_12353 (I212729,I2690);
DFFARX1 I_12354 (I315998,I2683,I212729,I212755,);
nand I_12355 (I212763,I316010,I315989);
and I_12356 (I212780,I212763,I316013);
DFFARX1 I_12357 (I212780,I2683,I212729,I212806,);
nor I_12358 (I212697,I212806,I212755);
not I_12359 (I212828,I212806);
DFFARX1 I_12360 (I316004,I2683,I212729,I212854,);
nand I_12361 (I212862,I212854,I315986);
not I_12362 (I212879,I212862);
DFFARX1 I_12363 (I212879,I2683,I212729,I212905,);
not I_12364 (I212721,I212905);
nor I_12365 (I212927,I212755,I212862);
nor I_12366 (I212703,I212806,I212927);
DFFARX1 I_12367 (I316001,I2683,I212729,I212967,);
DFFARX1 I_12368 (I212967,I2683,I212729,I212984,);
not I_12369 (I212992,I212984);
not I_12370 (I213009,I212967);
nand I_12371 (I212706,I213009,I212828);
nand I_12372 (I213040,I315986,I315992);
and I_12373 (I213057,I213040,I315995);
DFFARX1 I_12374 (I213057,I2683,I212729,I213083,);
nor I_12375 (I213091,I213083,I212755);
DFFARX1 I_12376 (I213091,I2683,I212729,I212694,);
DFFARX1 I_12377 (I213083,I2683,I212729,I212712,);
nor I_12378 (I213136,I316007,I315992);
not I_12379 (I213153,I213136);
nor I_12380 (I212715,I212992,I213153);
nand I_12381 (I212700,I213009,I213153);
nor I_12382 (I212709,I212755,I213136);
DFFARX1 I_12383 (I213136,I2683,I212729,I212718,);
not I_12384 (I213256,I2690);
DFFARX1 I_12385 (I982608,I2683,I213256,I213282,);
nand I_12386 (I213290,I982590,I982614);
and I_12387 (I213307,I213290,I982605);
DFFARX1 I_12388 (I213307,I2683,I213256,I213333,);
nor I_12389 (I213224,I213333,I213282);
not I_12390 (I213355,I213333);
DFFARX1 I_12391 (I982611,I2683,I213256,I213381,);
nand I_12392 (I213389,I213381,I982599);
not I_12393 (I213406,I213389);
DFFARX1 I_12394 (I213406,I2683,I213256,I213432,);
not I_12395 (I213248,I213432);
nor I_12396 (I213454,I213282,I213389);
nor I_12397 (I213230,I213333,I213454);
DFFARX1 I_12398 (I982590,I2683,I213256,I213494,);
DFFARX1 I_12399 (I213494,I2683,I213256,I213511,);
not I_12400 (I213519,I213511);
not I_12401 (I213536,I213494);
nand I_12402 (I213233,I213536,I213355);
nand I_12403 (I213567,I982596,I982593);
and I_12404 (I213584,I213567,I982602);
DFFARX1 I_12405 (I213584,I2683,I213256,I213610,);
nor I_12406 (I213618,I213610,I213282);
DFFARX1 I_12407 (I213618,I2683,I213256,I213221,);
DFFARX1 I_12408 (I213610,I2683,I213256,I213239,);
nor I_12409 (I213663,I982593,I982593);
not I_12410 (I213680,I213663);
nor I_12411 (I213242,I213519,I213680);
nand I_12412 (I213227,I213536,I213680);
nor I_12413 (I213236,I213282,I213663);
DFFARX1 I_12414 (I213663,I2683,I213256,I213245,);
not I_12415 (I213783,I2690);
DFFARX1 I_12416 (I86455,I2683,I213783,I213809,);
nand I_12417 (I213817,I86467,I86476);
and I_12418 (I213834,I213817,I86455);
DFFARX1 I_12419 (I213834,I2683,I213783,I213860,);
nor I_12420 (I213751,I213860,I213809);
not I_12421 (I213882,I213860);
DFFARX1 I_12422 (I86470,I2683,I213783,I213908,);
nand I_12423 (I213916,I213908,I86458);
not I_12424 (I213933,I213916);
DFFARX1 I_12425 (I213933,I2683,I213783,I213959,);
not I_12426 (I213775,I213959);
nor I_12427 (I213981,I213809,I213916);
nor I_12428 (I213757,I213860,I213981);
DFFARX1 I_12429 (I86461,I2683,I213783,I214021,);
DFFARX1 I_12430 (I214021,I2683,I213783,I214038,);
not I_12431 (I214046,I214038);
not I_12432 (I214063,I214021);
nand I_12433 (I213760,I214063,I213882);
nand I_12434 (I214094,I86452,I86452);
and I_12435 (I214111,I214094,I86464);
DFFARX1 I_12436 (I214111,I2683,I213783,I214137,);
nor I_12437 (I214145,I214137,I213809);
DFFARX1 I_12438 (I214145,I2683,I213783,I213748,);
DFFARX1 I_12439 (I214137,I2683,I213783,I213766,);
nor I_12440 (I214190,I86473,I86452);
not I_12441 (I214207,I214190);
nor I_12442 (I213769,I214046,I214207);
nand I_12443 (I213754,I214063,I214207);
nor I_12444 (I213763,I213809,I214190);
DFFARX1 I_12445 (I214190,I2683,I213783,I213772,);
not I_12446 (I214310,I2690);
DFFARX1 I_12447 (I65375,I2683,I214310,I214336,);
nand I_12448 (I214344,I65387,I65396);
and I_12449 (I214361,I214344,I65375);
DFFARX1 I_12450 (I214361,I2683,I214310,I214387,);
nor I_12451 (I214278,I214387,I214336);
not I_12452 (I214409,I214387);
DFFARX1 I_12453 (I65390,I2683,I214310,I214435,);
nand I_12454 (I214443,I214435,I65378);
not I_12455 (I214460,I214443);
DFFARX1 I_12456 (I214460,I2683,I214310,I214486,);
not I_12457 (I214302,I214486);
nor I_12458 (I214508,I214336,I214443);
nor I_12459 (I214284,I214387,I214508);
DFFARX1 I_12460 (I65381,I2683,I214310,I214548,);
DFFARX1 I_12461 (I214548,I2683,I214310,I214565,);
not I_12462 (I214573,I214565);
not I_12463 (I214590,I214548);
nand I_12464 (I214287,I214590,I214409);
nand I_12465 (I214621,I65372,I65372);
and I_12466 (I214638,I214621,I65384);
DFFARX1 I_12467 (I214638,I2683,I214310,I214664,);
nor I_12468 (I214672,I214664,I214336);
DFFARX1 I_12469 (I214672,I2683,I214310,I214275,);
DFFARX1 I_12470 (I214664,I2683,I214310,I214293,);
nor I_12471 (I214717,I65393,I65372);
not I_12472 (I214734,I214717);
nor I_12473 (I214296,I214573,I214734);
nand I_12474 (I214281,I214590,I214734);
nor I_12475 (I214290,I214336,I214717);
DFFARX1 I_12476 (I214717,I2683,I214310,I214299,);
not I_12477 (I214837,I2690);
DFFARX1 I_12478 (I597722,I2683,I214837,I214863,);
nand I_12479 (I214871,I597713,I597728);
and I_12480 (I214888,I214871,I597734);
DFFARX1 I_12481 (I214888,I2683,I214837,I214914,);
nor I_12482 (I214805,I214914,I214863);
not I_12483 (I214936,I214914);
DFFARX1 I_12484 (I597719,I2683,I214837,I214962,);
nand I_12485 (I214970,I214962,I597713);
not I_12486 (I214987,I214970);
DFFARX1 I_12487 (I214987,I2683,I214837,I215013,);
not I_12488 (I214829,I215013);
nor I_12489 (I215035,I214863,I214970);
nor I_12490 (I214811,I214914,I215035);
DFFARX1 I_12491 (I597716,I2683,I214837,I215075,);
DFFARX1 I_12492 (I215075,I2683,I214837,I215092,);
not I_12493 (I215100,I215092);
not I_12494 (I215117,I215075);
nand I_12495 (I214814,I215117,I214936);
nand I_12496 (I215148,I597710,I597725);
and I_12497 (I215165,I215148,I597710);
DFFARX1 I_12498 (I215165,I2683,I214837,I215191,);
nor I_12499 (I215199,I215191,I214863);
DFFARX1 I_12500 (I215199,I2683,I214837,I214802,);
DFFARX1 I_12501 (I215191,I2683,I214837,I214820,);
nor I_12502 (I215244,I597731,I597725);
not I_12503 (I215261,I215244);
nor I_12504 (I214823,I215100,I215261);
nand I_12505 (I214808,I215117,I215261);
nor I_12506 (I214817,I214863,I215244);
DFFARX1 I_12507 (I215244,I2683,I214837,I214826,);
not I_12508 (I215364,I2690);
DFFARX1 I_12509 (I326878,I2683,I215364,I215390,);
nand I_12510 (I215398,I326890,I326869);
and I_12511 (I215415,I215398,I326893);
DFFARX1 I_12512 (I215415,I2683,I215364,I215441,);
nor I_12513 (I215332,I215441,I215390);
not I_12514 (I215463,I215441);
DFFARX1 I_12515 (I326884,I2683,I215364,I215489,);
nand I_12516 (I215497,I215489,I326866);
not I_12517 (I215514,I215497);
DFFARX1 I_12518 (I215514,I2683,I215364,I215540,);
not I_12519 (I215356,I215540);
nor I_12520 (I215562,I215390,I215497);
nor I_12521 (I215338,I215441,I215562);
DFFARX1 I_12522 (I326881,I2683,I215364,I215602,);
DFFARX1 I_12523 (I215602,I2683,I215364,I215619,);
not I_12524 (I215627,I215619);
not I_12525 (I215644,I215602);
nand I_12526 (I215341,I215644,I215463);
nand I_12527 (I215675,I326866,I326872);
and I_12528 (I215692,I215675,I326875);
DFFARX1 I_12529 (I215692,I2683,I215364,I215718,);
nor I_12530 (I215726,I215718,I215390);
DFFARX1 I_12531 (I215726,I2683,I215364,I215329,);
DFFARX1 I_12532 (I215718,I2683,I215364,I215347,);
nor I_12533 (I215771,I326887,I326872);
not I_12534 (I215788,I215771);
nor I_12535 (I215350,I215627,I215788);
nand I_12536 (I215335,I215644,I215788);
nor I_12537 (I215344,I215390,I215771);
DFFARX1 I_12538 (I215771,I2683,I215364,I215353,);
not I_12539 (I215891,I2690);
DFFARX1 I_12540 (I179510,I2683,I215891,I215917,);
nand I_12541 (I215925,I179510,I179516);
and I_12542 (I215942,I215925,I179534);
DFFARX1 I_12543 (I215942,I2683,I215891,I215968,);
nor I_12544 (I215859,I215968,I215917);
not I_12545 (I215990,I215968);
DFFARX1 I_12546 (I179522,I2683,I215891,I216016,);
nand I_12547 (I216024,I216016,I179519);
not I_12548 (I216041,I216024);
DFFARX1 I_12549 (I216041,I2683,I215891,I216067,);
not I_12550 (I215883,I216067);
nor I_12551 (I216089,I215917,I216024);
nor I_12552 (I215865,I215968,I216089);
DFFARX1 I_12553 (I179528,I2683,I215891,I216129,);
DFFARX1 I_12554 (I216129,I2683,I215891,I216146,);
not I_12555 (I216154,I216146);
not I_12556 (I216171,I216129);
nand I_12557 (I215868,I216171,I215990);
nand I_12558 (I216202,I179513,I179513);
and I_12559 (I216219,I216202,I179525);
DFFARX1 I_12560 (I216219,I2683,I215891,I216245,);
nor I_12561 (I216253,I216245,I215917);
DFFARX1 I_12562 (I216253,I2683,I215891,I215856,);
DFFARX1 I_12563 (I216245,I2683,I215891,I215874,);
nor I_12564 (I216298,I179531,I179513);
not I_12565 (I216315,I216298);
nor I_12566 (I215877,I216154,I216315);
nand I_12567 (I215862,I216171,I216315);
nor I_12568 (I215871,I215917,I216298);
DFFARX1 I_12569 (I216298,I2683,I215891,I215880,);
not I_12570 (I216418,I2690);
DFFARX1 I_12571 (I962480,I2683,I216418,I216444,);
nand I_12572 (I216452,I962462,I962486);
and I_12573 (I216469,I216452,I962477);
DFFARX1 I_12574 (I216469,I2683,I216418,I216495,);
nor I_12575 (I216386,I216495,I216444);
not I_12576 (I216517,I216495);
DFFARX1 I_12577 (I962483,I2683,I216418,I216543,);
nand I_12578 (I216551,I216543,I962471);
not I_12579 (I216568,I216551);
DFFARX1 I_12580 (I216568,I2683,I216418,I216594,);
not I_12581 (I216410,I216594);
nor I_12582 (I216616,I216444,I216551);
nor I_12583 (I216392,I216495,I216616);
DFFARX1 I_12584 (I962462,I2683,I216418,I216656,);
DFFARX1 I_12585 (I216656,I2683,I216418,I216673,);
not I_12586 (I216681,I216673);
not I_12587 (I216698,I216656);
nand I_12588 (I216395,I216698,I216517);
nand I_12589 (I216729,I962468,I962465);
and I_12590 (I216746,I216729,I962474);
DFFARX1 I_12591 (I216746,I2683,I216418,I216772,);
nor I_12592 (I216780,I216772,I216444);
DFFARX1 I_12593 (I216780,I2683,I216418,I216383,);
DFFARX1 I_12594 (I216772,I2683,I216418,I216401,);
nor I_12595 (I216825,I962465,I962465);
not I_12596 (I216842,I216825);
nor I_12597 (I216404,I216681,I216842);
nand I_12598 (I216389,I216698,I216842);
nor I_12599 (I216398,I216444,I216825);
DFFARX1 I_12600 (I216825,I2683,I216418,I216407,);
not I_12601 (I216945,I2690);
DFFARX1 I_12602 (I499462,I2683,I216945,I216971,);
nand I_12603 (I216979,I499453,I499468);
and I_12604 (I216996,I216979,I499474);
DFFARX1 I_12605 (I216996,I2683,I216945,I217022,);
nor I_12606 (I216913,I217022,I216971);
not I_12607 (I217044,I217022);
DFFARX1 I_12608 (I499459,I2683,I216945,I217070,);
nand I_12609 (I217078,I217070,I499453);
not I_12610 (I217095,I217078);
DFFARX1 I_12611 (I217095,I2683,I216945,I217121,);
not I_12612 (I216937,I217121);
nor I_12613 (I217143,I216971,I217078);
nor I_12614 (I216919,I217022,I217143);
DFFARX1 I_12615 (I499456,I2683,I216945,I217183,);
DFFARX1 I_12616 (I217183,I2683,I216945,I217200,);
not I_12617 (I217208,I217200);
not I_12618 (I217225,I217183);
nand I_12619 (I216922,I217225,I217044);
nand I_12620 (I217256,I499450,I499465);
and I_12621 (I217273,I217256,I499450);
DFFARX1 I_12622 (I217273,I2683,I216945,I217299,);
nor I_12623 (I217307,I217299,I216971);
DFFARX1 I_12624 (I217307,I2683,I216945,I216910,);
DFFARX1 I_12625 (I217299,I2683,I216945,I216928,);
nor I_12626 (I217352,I499471,I499465);
not I_12627 (I217369,I217352);
nor I_12628 (I216931,I217208,I217369);
nand I_12629 (I216916,I217225,I217369);
nor I_12630 (I216925,I216971,I217352);
DFFARX1 I_12631 (I217352,I2683,I216945,I216934,);
not I_12632 (I217472,I2690);
DFFARX1 I_12633 (I396705,I2683,I217472,I217498,);
nand I_12634 (I217506,I396705,I396717);
and I_12635 (I217523,I217506,I396702);
DFFARX1 I_12636 (I217523,I2683,I217472,I217549,);
nor I_12637 (I217440,I217549,I217498);
not I_12638 (I217571,I217549);
DFFARX1 I_12639 (I396726,I2683,I217472,I217597,);
nand I_12640 (I217605,I217597,I396723);
not I_12641 (I217622,I217605);
DFFARX1 I_12642 (I217622,I2683,I217472,I217648,);
not I_12643 (I217464,I217648);
nor I_12644 (I217670,I217498,I217605);
nor I_12645 (I217446,I217549,I217670);
DFFARX1 I_12646 (I396714,I2683,I217472,I217710,);
DFFARX1 I_12647 (I217710,I2683,I217472,I217727,);
not I_12648 (I217735,I217727);
not I_12649 (I217752,I217710);
nand I_12650 (I217449,I217752,I217571);
nand I_12651 (I217783,I396702,I396711);
and I_12652 (I217800,I217783,I396720);
DFFARX1 I_12653 (I217800,I2683,I217472,I217826,);
nor I_12654 (I217834,I217826,I217498);
DFFARX1 I_12655 (I217834,I2683,I217472,I217437,);
DFFARX1 I_12656 (I217826,I2683,I217472,I217455,);
nor I_12657 (I217879,I396708,I396711);
not I_12658 (I217896,I217879);
nor I_12659 (I217458,I217735,I217896);
nand I_12660 (I217443,I217752,I217896);
nor I_12661 (I217452,I217498,I217879);
DFFARX1 I_12662 (I217879,I2683,I217472,I217461,);
not I_12663 (I217999,I2690);
DFFARX1 I_12664 (I1015755,I2683,I217999,I218025,);
nand I_12665 (I218033,I1015752,I1015743);
and I_12666 (I218050,I218033,I1015740);
DFFARX1 I_12667 (I218050,I2683,I217999,I218076,);
nor I_12668 (I217967,I218076,I218025);
not I_12669 (I218098,I218076);
DFFARX1 I_12670 (I1015749,I2683,I217999,I218124,);
nand I_12671 (I218132,I218124,I1015758);
not I_12672 (I218149,I218132);
DFFARX1 I_12673 (I218149,I2683,I217999,I218175,);
not I_12674 (I217991,I218175);
nor I_12675 (I218197,I218025,I218132);
nor I_12676 (I217973,I218076,I218197);
DFFARX1 I_12677 (I1015761,I2683,I217999,I218237,);
DFFARX1 I_12678 (I218237,I2683,I217999,I218254,);
not I_12679 (I218262,I218254);
not I_12680 (I218279,I218237);
nand I_12681 (I217976,I218279,I218098);
nand I_12682 (I218310,I1015740,I1015746);
and I_12683 (I218327,I218310,I1015764);
DFFARX1 I_12684 (I218327,I2683,I217999,I218353,);
nor I_12685 (I218361,I218353,I218025);
DFFARX1 I_12686 (I218361,I2683,I217999,I217964,);
DFFARX1 I_12687 (I218353,I2683,I217999,I217982,);
nor I_12688 (I218406,I1015743,I1015746);
not I_12689 (I218423,I218406);
nor I_12690 (I217985,I218262,I218423);
nand I_12691 (I217970,I218279,I218423);
nor I_12692 (I217979,I218025,I218406);
DFFARX1 I_12693 (I218406,I2683,I217999,I217988,);
not I_12694 (I218526,I2690);
DFFARX1 I_12695 (I950154,I2683,I218526,I218552,);
nand I_12696 (I218560,I950169,I950154);
and I_12697 (I218577,I218560,I950172);
DFFARX1 I_12698 (I218577,I2683,I218526,I218603,);
nor I_12699 (I218494,I218603,I218552);
not I_12700 (I218625,I218603);
DFFARX1 I_12701 (I950178,I2683,I218526,I218651,);
nand I_12702 (I218659,I218651,I950160);
not I_12703 (I218676,I218659);
DFFARX1 I_12704 (I218676,I2683,I218526,I218702,);
not I_12705 (I218518,I218702);
nor I_12706 (I218724,I218552,I218659);
nor I_12707 (I218500,I218603,I218724);
DFFARX1 I_12708 (I950157,I2683,I218526,I218764,);
DFFARX1 I_12709 (I218764,I2683,I218526,I218781,);
not I_12710 (I218789,I218781);
not I_12711 (I218806,I218764);
nand I_12712 (I218503,I218806,I218625);
nand I_12713 (I218837,I950157,I950163);
and I_12714 (I218854,I218837,I950175);
DFFARX1 I_12715 (I218854,I2683,I218526,I218880,);
nor I_12716 (I218888,I218880,I218552);
DFFARX1 I_12717 (I218888,I2683,I218526,I218491,);
DFFARX1 I_12718 (I218880,I2683,I218526,I218509,);
nor I_12719 (I218933,I950166,I950163);
not I_12720 (I218950,I218933);
nor I_12721 (I218512,I218789,I218950);
nand I_12722 (I218497,I218806,I218950);
nor I_12723 (I218506,I218552,I218933);
DFFARX1 I_12724 (I218933,I2683,I218526,I218515,);
not I_12725 (I219053,I2690);
DFFARX1 I_12726 (I476923,I2683,I219053,I219079,);
nand I_12727 (I219087,I476908,I476911);
and I_12728 (I219104,I219087,I476926);
DFFARX1 I_12729 (I219104,I2683,I219053,I219130,);
nor I_12730 (I219021,I219130,I219079);
not I_12731 (I219152,I219130);
DFFARX1 I_12732 (I476920,I2683,I219053,I219178,);
nand I_12733 (I219186,I219178,I476911);
not I_12734 (I219203,I219186);
DFFARX1 I_12735 (I219203,I2683,I219053,I219229,);
not I_12736 (I219045,I219229);
nor I_12737 (I219251,I219079,I219186);
nor I_12738 (I219027,I219130,I219251);
DFFARX1 I_12739 (I476917,I2683,I219053,I219291,);
DFFARX1 I_12740 (I219291,I2683,I219053,I219308,);
not I_12741 (I219316,I219308);
not I_12742 (I219333,I219291);
nand I_12743 (I219030,I219333,I219152);
nand I_12744 (I219364,I476932,I476908);
and I_12745 (I219381,I219364,I476929);
DFFARX1 I_12746 (I219381,I2683,I219053,I219407,);
nor I_12747 (I219415,I219407,I219079);
DFFARX1 I_12748 (I219415,I2683,I219053,I219018,);
DFFARX1 I_12749 (I219407,I2683,I219053,I219036,);
nor I_12750 (I219460,I476914,I476908);
not I_12751 (I219477,I219460);
nor I_12752 (I219039,I219316,I219477);
nand I_12753 (I219024,I219333,I219477);
nor I_12754 (I219033,I219079,I219460);
DFFARX1 I_12755 (I219460,I2683,I219053,I219042,);
not I_12756 (I219580,I2690);
DFFARX1 I_12757 (I755524,I2683,I219580,I219606,);
nand I_12758 (I219614,I755521,I755539);
and I_12759 (I219631,I219614,I755530);
DFFARX1 I_12760 (I219631,I2683,I219580,I219657,);
nor I_12761 (I219548,I219657,I219606);
not I_12762 (I219679,I219657);
DFFARX1 I_12763 (I755545,I2683,I219580,I219705,);
nand I_12764 (I219713,I219705,I755527);
not I_12765 (I219730,I219713);
DFFARX1 I_12766 (I219730,I2683,I219580,I219756,);
not I_12767 (I219572,I219756);
nor I_12768 (I219778,I219606,I219713);
nor I_12769 (I219554,I219657,I219778);
DFFARX1 I_12770 (I755533,I2683,I219580,I219818,);
DFFARX1 I_12771 (I219818,I2683,I219580,I219835,);
not I_12772 (I219843,I219835);
not I_12773 (I219860,I219818);
nand I_12774 (I219557,I219860,I219679);
nand I_12775 (I219891,I755521,I755548);
and I_12776 (I219908,I219891,I755536);
DFFARX1 I_12777 (I219908,I2683,I219580,I219934,);
nor I_12778 (I219942,I219934,I219606);
DFFARX1 I_12779 (I219942,I2683,I219580,I219545,);
DFFARX1 I_12780 (I219934,I2683,I219580,I219563,);
nor I_12781 (I219987,I755542,I755548);
not I_12782 (I220004,I219987);
nor I_12783 (I219566,I219843,I220004);
nand I_12784 (I219551,I219860,I220004);
nor I_12785 (I219560,I219606,I219987);
DFFARX1 I_12786 (I219987,I2683,I219580,I219569,);
not I_12787 (I220107,I2690);
DFFARX1 I_12788 (I336670,I2683,I220107,I220133,);
nand I_12789 (I220141,I336682,I336661);
and I_12790 (I220158,I220141,I336685);
DFFARX1 I_12791 (I220158,I2683,I220107,I220184,);
nor I_12792 (I220075,I220184,I220133);
not I_12793 (I220206,I220184);
DFFARX1 I_12794 (I336676,I2683,I220107,I220232,);
nand I_12795 (I220240,I220232,I336658);
not I_12796 (I220257,I220240);
DFFARX1 I_12797 (I220257,I2683,I220107,I220283,);
not I_12798 (I220099,I220283);
nor I_12799 (I220305,I220133,I220240);
nor I_12800 (I220081,I220184,I220305);
DFFARX1 I_12801 (I336673,I2683,I220107,I220345,);
DFFARX1 I_12802 (I220345,I2683,I220107,I220362,);
not I_12803 (I220370,I220362);
not I_12804 (I220387,I220345);
nand I_12805 (I220084,I220387,I220206);
nand I_12806 (I220418,I336658,I336664);
and I_12807 (I220435,I220418,I336667);
DFFARX1 I_12808 (I220435,I2683,I220107,I220461,);
nor I_12809 (I220469,I220461,I220133);
DFFARX1 I_12810 (I220469,I2683,I220107,I220072,);
DFFARX1 I_12811 (I220461,I2683,I220107,I220090,);
nor I_12812 (I220514,I336679,I336664);
not I_12813 (I220531,I220514);
nor I_12814 (I220093,I220370,I220531);
nand I_12815 (I220078,I220387,I220531);
nor I_12816 (I220087,I220133,I220514);
DFFARX1 I_12817 (I220514,I2683,I220107,I220096,);
not I_12818 (I220634,I2690);
DFFARX1 I_12819 (I56943,I2683,I220634,I220660,);
nand I_12820 (I220668,I56955,I56964);
and I_12821 (I220685,I220668,I56943);
DFFARX1 I_12822 (I220685,I2683,I220634,I220711,);
nor I_12823 (I220602,I220711,I220660);
not I_12824 (I220733,I220711);
DFFARX1 I_12825 (I56958,I2683,I220634,I220759,);
nand I_12826 (I220767,I220759,I56946);
not I_12827 (I220784,I220767);
DFFARX1 I_12828 (I220784,I2683,I220634,I220810,);
not I_12829 (I220626,I220810);
nor I_12830 (I220832,I220660,I220767);
nor I_12831 (I220608,I220711,I220832);
DFFARX1 I_12832 (I56949,I2683,I220634,I220872,);
DFFARX1 I_12833 (I220872,I2683,I220634,I220889,);
not I_12834 (I220897,I220889);
not I_12835 (I220914,I220872);
nand I_12836 (I220611,I220914,I220733);
nand I_12837 (I220945,I56940,I56940);
and I_12838 (I220962,I220945,I56952);
DFFARX1 I_12839 (I220962,I2683,I220634,I220988,);
nor I_12840 (I220996,I220988,I220660);
DFFARX1 I_12841 (I220996,I2683,I220634,I220599,);
DFFARX1 I_12842 (I220988,I2683,I220634,I220617,);
nor I_12843 (I221041,I56961,I56940);
not I_12844 (I221058,I221041);
nor I_12845 (I220620,I220897,I221058);
nand I_12846 (I220605,I220914,I221058);
nor I_12847 (I220614,I220660,I221041);
DFFARX1 I_12848 (I221041,I2683,I220634,I220623,);
not I_12849 (I221161,I2690);
DFFARX1 I_12850 (I1062630,I2683,I221161,I221187,);
nand I_12851 (I221195,I1062609,I1062609);
and I_12852 (I221212,I221195,I1062636);
DFFARX1 I_12853 (I221212,I2683,I221161,I221238,);
nor I_12854 (I221129,I221238,I221187);
not I_12855 (I221260,I221238);
DFFARX1 I_12856 (I1062624,I2683,I221161,I221286,);
nand I_12857 (I221294,I221286,I1062627);
not I_12858 (I221311,I221294);
DFFARX1 I_12859 (I221311,I2683,I221161,I221337,);
not I_12860 (I221153,I221337);
nor I_12861 (I221359,I221187,I221294);
nor I_12862 (I221135,I221238,I221359);
DFFARX1 I_12863 (I1062618,I2683,I221161,I221399,);
DFFARX1 I_12864 (I221399,I2683,I221161,I221416,);
not I_12865 (I221424,I221416);
not I_12866 (I221441,I221399);
nand I_12867 (I221138,I221441,I221260);
nand I_12868 (I221472,I1062615,I1062612);
and I_12869 (I221489,I221472,I1062633);
DFFARX1 I_12870 (I221489,I2683,I221161,I221515,);
nor I_12871 (I221523,I221515,I221187);
DFFARX1 I_12872 (I221523,I2683,I221161,I221126,);
DFFARX1 I_12873 (I221515,I2683,I221161,I221144,);
nor I_12874 (I221568,I1062621,I1062612);
not I_12875 (I221585,I221568);
nor I_12876 (I221147,I221424,I221585);
nand I_12877 (I221132,I221441,I221585);
nor I_12878 (I221141,I221187,I221568);
DFFARX1 I_12879 (I221568,I2683,I221161,I221150,);
not I_12880 (I221688,I2690);
DFFARX1 I_12881 (I740666,I2683,I221688,I221714,);
nand I_12882 (I221722,I740663,I740681);
and I_12883 (I221739,I221722,I740672);
DFFARX1 I_12884 (I221739,I2683,I221688,I221765,);
nor I_12885 (I221656,I221765,I221714);
not I_12886 (I221787,I221765);
DFFARX1 I_12887 (I740687,I2683,I221688,I221813,);
nand I_12888 (I221821,I221813,I740669);
not I_12889 (I221838,I221821);
DFFARX1 I_12890 (I221838,I2683,I221688,I221864,);
not I_12891 (I221680,I221864);
nor I_12892 (I221886,I221714,I221821);
nor I_12893 (I221662,I221765,I221886);
DFFARX1 I_12894 (I740675,I2683,I221688,I221926,);
DFFARX1 I_12895 (I221926,I2683,I221688,I221943,);
not I_12896 (I221951,I221943);
not I_12897 (I221968,I221926);
nand I_12898 (I221665,I221968,I221787);
nand I_12899 (I221999,I740663,I740690);
and I_12900 (I222016,I221999,I740678);
DFFARX1 I_12901 (I222016,I2683,I221688,I222042,);
nor I_12902 (I222050,I222042,I221714);
DFFARX1 I_12903 (I222050,I2683,I221688,I221653,);
DFFARX1 I_12904 (I222042,I2683,I221688,I221671,);
nor I_12905 (I222095,I740684,I740690);
not I_12906 (I222112,I222095);
nor I_12907 (I221674,I221951,I222112);
nand I_12908 (I221659,I221968,I222112);
nor I_12909 (I221668,I221714,I222095);
DFFARX1 I_12910 (I222095,I2683,I221688,I221677,);
not I_12911 (I222215,I2690);
DFFARX1 I_12912 (I34806,I2683,I222215,I222241,);
nand I_12913 (I222249,I34830,I34809);
and I_12914 (I222266,I222249,I34806);
DFFARX1 I_12915 (I222266,I2683,I222215,I222292,);
nor I_12916 (I222183,I222292,I222241);
not I_12917 (I222314,I222292);
DFFARX1 I_12918 (I34812,I2683,I222215,I222340,);
nand I_12919 (I222348,I222340,I34821);
not I_12920 (I222365,I222348);
DFFARX1 I_12921 (I222365,I2683,I222215,I222391,);
not I_12922 (I222207,I222391);
nor I_12923 (I222413,I222241,I222348);
nor I_12924 (I222189,I222292,I222413);
DFFARX1 I_12925 (I34815,I2683,I222215,I222453,);
DFFARX1 I_12926 (I222453,I2683,I222215,I222470,);
not I_12927 (I222478,I222470);
not I_12928 (I222495,I222453);
nand I_12929 (I222192,I222495,I222314);
nand I_12930 (I222526,I34827,I34809);
and I_12931 (I222543,I222526,I34818);
DFFARX1 I_12932 (I222543,I2683,I222215,I222569,);
nor I_12933 (I222577,I222569,I222241);
DFFARX1 I_12934 (I222577,I2683,I222215,I222180,);
DFFARX1 I_12935 (I222569,I2683,I222215,I222198,);
nor I_12936 (I222622,I34824,I34809);
not I_12937 (I222639,I222622);
nor I_12938 (I222201,I222478,I222639);
nand I_12939 (I222186,I222495,I222639);
nor I_12940 (I222195,I222241,I222622);
DFFARX1 I_12941 (I222622,I2683,I222215,I222204,);
not I_12942 (I222742,I2690);
DFFARX1 I_12943 (I36914,I2683,I222742,I222768,);
nand I_12944 (I222776,I36938,I36917);
and I_12945 (I222793,I222776,I36914);
DFFARX1 I_12946 (I222793,I2683,I222742,I222819,);
nor I_12947 (I222710,I222819,I222768);
not I_12948 (I222841,I222819);
DFFARX1 I_12949 (I36920,I2683,I222742,I222867,);
nand I_12950 (I222875,I222867,I36929);
not I_12951 (I222892,I222875);
DFFARX1 I_12952 (I222892,I2683,I222742,I222918,);
not I_12953 (I222734,I222918);
nor I_12954 (I222940,I222768,I222875);
nor I_12955 (I222716,I222819,I222940);
DFFARX1 I_12956 (I36923,I2683,I222742,I222980,);
DFFARX1 I_12957 (I222980,I2683,I222742,I222997,);
not I_12958 (I223005,I222997);
not I_12959 (I223022,I222980);
nand I_12960 (I222719,I223022,I222841);
nand I_12961 (I223053,I36935,I36917);
and I_12962 (I223070,I223053,I36926);
DFFARX1 I_12963 (I223070,I2683,I222742,I223096,);
nor I_12964 (I223104,I223096,I222768);
DFFARX1 I_12965 (I223104,I2683,I222742,I222707,);
DFFARX1 I_12966 (I223096,I2683,I222742,I222725,);
nor I_12967 (I223149,I36932,I36917);
not I_12968 (I223166,I223149);
nor I_12969 (I222728,I223005,I223166);
nand I_12970 (I222713,I223022,I223166);
nor I_12971 (I222722,I222768,I223149);
DFFARX1 I_12972 (I223149,I2683,I222742,I222731,);
not I_12973 (I223269,I2690);
DFFARX1 I_12974 (I578648,I2683,I223269,I223295,);
nand I_12975 (I223303,I578639,I578654);
and I_12976 (I223320,I223303,I578660);
DFFARX1 I_12977 (I223320,I2683,I223269,I223346,);
nor I_12978 (I223237,I223346,I223295);
not I_12979 (I223368,I223346);
DFFARX1 I_12980 (I578645,I2683,I223269,I223394,);
nand I_12981 (I223402,I223394,I578639);
not I_12982 (I223419,I223402);
DFFARX1 I_12983 (I223419,I2683,I223269,I223445,);
not I_12984 (I223261,I223445);
nor I_12985 (I223467,I223295,I223402);
nor I_12986 (I223243,I223346,I223467);
DFFARX1 I_12987 (I578642,I2683,I223269,I223507,);
DFFARX1 I_12988 (I223507,I2683,I223269,I223524,);
not I_12989 (I223532,I223524);
not I_12990 (I223549,I223507);
nand I_12991 (I223246,I223549,I223368);
nand I_12992 (I223580,I578636,I578651);
and I_12993 (I223597,I223580,I578636);
DFFARX1 I_12994 (I223597,I2683,I223269,I223623,);
nor I_12995 (I223631,I223623,I223295);
DFFARX1 I_12996 (I223631,I2683,I223269,I223234,);
DFFARX1 I_12997 (I223623,I2683,I223269,I223252,);
nor I_12998 (I223676,I578657,I578651);
not I_12999 (I223693,I223676);
nor I_13000 (I223255,I223532,I223693);
nand I_13001 (I223240,I223549,I223693);
nor I_13002 (I223249,I223295,I223676);
DFFARX1 I_13003 (I223676,I2683,I223269,I223258,);
not I_13004 (I223796,I2690);
DFFARX1 I_13005 (I391070,I2683,I223796,I223822,);
nand I_13006 (I223830,I391082,I391061);
and I_13007 (I223847,I223830,I391085);
DFFARX1 I_13008 (I223847,I2683,I223796,I223873,);
nor I_13009 (I223764,I223873,I223822);
not I_13010 (I223895,I223873);
DFFARX1 I_13011 (I391076,I2683,I223796,I223921,);
nand I_13012 (I223929,I223921,I391058);
not I_13013 (I223946,I223929);
DFFARX1 I_13014 (I223946,I2683,I223796,I223972,);
not I_13015 (I223788,I223972);
nor I_13016 (I223994,I223822,I223929);
nor I_13017 (I223770,I223873,I223994);
DFFARX1 I_13018 (I391073,I2683,I223796,I224034,);
DFFARX1 I_13019 (I224034,I2683,I223796,I224051,);
not I_13020 (I224059,I224051);
not I_13021 (I224076,I224034);
nand I_13022 (I223773,I224076,I223895);
nand I_13023 (I224107,I391058,I391064);
and I_13024 (I224124,I224107,I391067);
DFFARX1 I_13025 (I224124,I2683,I223796,I224150,);
nor I_13026 (I224158,I224150,I223822);
DFFARX1 I_13027 (I224158,I2683,I223796,I223761,);
DFFARX1 I_13028 (I224150,I2683,I223796,I223779,);
nor I_13029 (I224203,I391079,I391064);
not I_13030 (I224220,I224203);
nor I_13031 (I223782,I224059,I224220);
nand I_13032 (I223767,I224076,I224220);
nor I_13033 (I223776,I223822,I224203);
DFFARX1 I_13034 (I224203,I2683,I223796,I223785,);
not I_13035 (I224323,I2690);
DFFARX1 I_13036 (I12145,I2683,I224323,I224349,);
nand I_13037 (I224357,I12169,I12148);
and I_13038 (I224374,I224357,I12145);
DFFARX1 I_13039 (I224374,I2683,I224323,I224400,);
nor I_13040 (I224291,I224400,I224349);
not I_13041 (I224422,I224400);
DFFARX1 I_13042 (I12151,I2683,I224323,I224448,);
nand I_13043 (I224456,I224448,I12160);
not I_13044 (I224473,I224456);
DFFARX1 I_13045 (I224473,I2683,I224323,I224499,);
not I_13046 (I224315,I224499);
nor I_13047 (I224521,I224349,I224456);
nor I_13048 (I224297,I224400,I224521);
DFFARX1 I_13049 (I12154,I2683,I224323,I224561,);
DFFARX1 I_13050 (I224561,I2683,I224323,I224578,);
not I_13051 (I224586,I224578);
not I_13052 (I224603,I224561);
nand I_13053 (I224300,I224603,I224422);
nand I_13054 (I224634,I12166,I12148);
and I_13055 (I224651,I224634,I12157);
DFFARX1 I_13056 (I224651,I2683,I224323,I224677,);
nor I_13057 (I224685,I224677,I224349);
DFFARX1 I_13058 (I224685,I2683,I224323,I224288,);
DFFARX1 I_13059 (I224677,I2683,I224323,I224306,);
nor I_13060 (I224730,I12163,I12148);
not I_13061 (I224747,I224730);
nor I_13062 (I224309,I224586,I224747);
nand I_13063 (I224294,I224603,I224747);
nor I_13064 (I224303,I224349,I224730);
DFFARX1 I_13065 (I224730,I2683,I224323,I224312,);
not I_13066 (I224850,I2690);
DFFARX1 I_13067 (I592520,I2683,I224850,I224876,);
nand I_13068 (I224884,I592511,I592526);
and I_13069 (I224901,I224884,I592532);
DFFARX1 I_13070 (I224901,I2683,I224850,I224927,);
nor I_13071 (I224818,I224927,I224876);
not I_13072 (I224949,I224927);
DFFARX1 I_13073 (I592517,I2683,I224850,I224975,);
nand I_13074 (I224983,I224975,I592511);
not I_13075 (I225000,I224983);
DFFARX1 I_13076 (I225000,I2683,I224850,I225026,);
not I_13077 (I224842,I225026);
nor I_13078 (I225048,I224876,I224983);
nor I_13079 (I224824,I224927,I225048);
DFFARX1 I_13080 (I592514,I2683,I224850,I225088,);
DFFARX1 I_13081 (I225088,I2683,I224850,I225105,);
not I_13082 (I225113,I225105);
not I_13083 (I225130,I225088);
nand I_13084 (I224827,I225130,I224949);
nand I_13085 (I225161,I592508,I592523);
and I_13086 (I225178,I225161,I592508);
DFFARX1 I_13087 (I225178,I2683,I224850,I225204,);
nor I_13088 (I225212,I225204,I224876);
DFFARX1 I_13089 (I225212,I2683,I224850,I224815,);
DFFARX1 I_13090 (I225204,I2683,I224850,I224833,);
nor I_13091 (I225257,I592529,I592523);
not I_13092 (I225274,I225257);
nor I_13093 (I224836,I225113,I225274);
nand I_13094 (I224821,I225130,I225274);
nor I_13095 (I224830,I224876,I225257);
DFFARX1 I_13096 (I225257,I2683,I224850,I224839,);
not I_13097 (I225377,I2690);
DFFARX1 I_13098 (I1002461,I2683,I225377,I225403,);
nand I_13099 (I225411,I1002458,I1002449);
and I_13100 (I225428,I225411,I1002446);
DFFARX1 I_13101 (I225428,I2683,I225377,I225454,);
nor I_13102 (I225345,I225454,I225403);
not I_13103 (I225476,I225454);
DFFARX1 I_13104 (I1002455,I2683,I225377,I225502,);
nand I_13105 (I225510,I225502,I1002464);
not I_13106 (I225527,I225510);
DFFARX1 I_13107 (I225527,I2683,I225377,I225553,);
not I_13108 (I225369,I225553);
nor I_13109 (I225575,I225403,I225510);
nor I_13110 (I225351,I225454,I225575);
DFFARX1 I_13111 (I1002467,I2683,I225377,I225615,);
DFFARX1 I_13112 (I225615,I2683,I225377,I225632,);
not I_13113 (I225640,I225632);
not I_13114 (I225657,I225615);
nand I_13115 (I225354,I225657,I225476);
nand I_13116 (I225688,I1002446,I1002452);
and I_13117 (I225705,I225688,I1002470);
DFFARX1 I_13118 (I225705,I2683,I225377,I225731,);
nor I_13119 (I225739,I225731,I225403);
DFFARX1 I_13120 (I225739,I2683,I225377,I225342,);
DFFARX1 I_13121 (I225731,I2683,I225377,I225360,);
nor I_13122 (I225784,I1002449,I1002452);
not I_13123 (I225801,I225784);
nor I_13124 (I225363,I225640,I225801);
nand I_13125 (I225348,I225657,I225801);
nor I_13126 (I225357,I225403,I225784);
DFFARX1 I_13127 (I225784,I2683,I225377,I225366,);
not I_13128 (I225904,I2690);
DFFARX1 I_13129 (I819223,I2683,I225904,I225930,);
nand I_13130 (I225938,I819220,I819223);
and I_13131 (I225955,I225938,I819232);
DFFARX1 I_13132 (I225955,I2683,I225904,I225981,);
nor I_13133 (I225872,I225981,I225930);
not I_13134 (I226003,I225981);
DFFARX1 I_13135 (I819220,I2683,I225904,I226029,);
nand I_13136 (I226037,I226029,I819238);
not I_13137 (I226054,I226037);
DFFARX1 I_13138 (I226054,I2683,I225904,I226080,);
not I_13139 (I225896,I226080);
nor I_13140 (I226102,I225930,I226037);
nor I_13141 (I225878,I225981,I226102);
DFFARX1 I_13142 (I819226,I2683,I225904,I226142,);
DFFARX1 I_13143 (I226142,I2683,I225904,I226159,);
not I_13144 (I226167,I226159);
not I_13145 (I226184,I226142);
nand I_13146 (I225881,I226184,I226003);
nand I_13147 (I226215,I819235,I819241);
and I_13148 (I226232,I226215,I819226);
DFFARX1 I_13149 (I226232,I2683,I225904,I226258,);
nor I_13150 (I226266,I226258,I225930);
DFFARX1 I_13151 (I226266,I2683,I225904,I225869,);
DFFARX1 I_13152 (I226258,I2683,I225904,I225887,);
nor I_13153 (I226311,I819229,I819241);
not I_13154 (I226328,I226311);
nor I_13155 (I225890,I226167,I226328);
nand I_13156 (I225875,I226184,I226328);
nor I_13157 (I225884,I225930,I226311);
DFFARX1 I_13158 (I226311,I2683,I225904,I225893,);
not I_13159 (I226431,I2690);
DFFARX1 I_13160 (I204500,I2683,I226431,I226457,);
nand I_13161 (I226465,I204500,I204506);
and I_13162 (I226482,I226465,I204524);
DFFARX1 I_13163 (I226482,I2683,I226431,I226508,);
nor I_13164 (I226399,I226508,I226457);
not I_13165 (I226530,I226508);
DFFARX1 I_13166 (I204512,I2683,I226431,I226556,);
nand I_13167 (I226564,I226556,I204509);
not I_13168 (I226581,I226564);
DFFARX1 I_13169 (I226581,I2683,I226431,I226607,);
not I_13170 (I226423,I226607);
nor I_13171 (I226629,I226457,I226564);
nor I_13172 (I226405,I226508,I226629);
DFFARX1 I_13173 (I204518,I2683,I226431,I226669,);
DFFARX1 I_13174 (I226669,I2683,I226431,I226686,);
not I_13175 (I226694,I226686);
not I_13176 (I226711,I226669);
nand I_13177 (I226408,I226711,I226530);
nand I_13178 (I226742,I204503,I204503);
and I_13179 (I226759,I226742,I204515);
DFFARX1 I_13180 (I226759,I2683,I226431,I226785,);
nor I_13181 (I226793,I226785,I226457);
DFFARX1 I_13182 (I226793,I2683,I226431,I226396,);
DFFARX1 I_13183 (I226785,I2683,I226431,I226414,);
nor I_13184 (I226838,I204521,I204503);
not I_13185 (I226855,I226838);
nor I_13186 (I226417,I226694,I226855);
nand I_13187 (I226402,I226711,I226855);
nor I_13188 (I226411,I226457,I226838);
DFFARX1 I_13189 (I226838,I2683,I226431,I226420,);
not I_13190 (I226958,I2690);
DFFARX1 I_13191 (I2396,I2683,I226958,I226984,);
nand I_13192 (I226992,I2172,I1644);
and I_13193 (I227009,I226992,I1956);
DFFARX1 I_13194 (I227009,I2683,I226958,I227035,);
nor I_13195 (I226926,I227035,I226984);
not I_13196 (I227057,I227035);
DFFARX1 I_13197 (I1532,I2683,I226958,I227083,);
nand I_13198 (I227091,I227083,I1852);
not I_13199 (I227108,I227091);
DFFARX1 I_13200 (I227108,I2683,I226958,I227134,);
not I_13201 (I226950,I227134);
nor I_13202 (I227156,I226984,I227091);
nor I_13203 (I226932,I227035,I227156);
DFFARX1 I_13204 (I2124,I2683,I226958,I227196,);
DFFARX1 I_13205 (I227196,I2683,I226958,I227213,);
not I_13206 (I227221,I227213);
not I_13207 (I227238,I227196);
nand I_13208 (I226935,I227238,I227057);
nand I_13209 (I227269,I2484,I2444);
and I_13210 (I227286,I227269,I1580);
DFFARX1 I_13211 (I227286,I2683,I226958,I227312,);
nor I_13212 (I227320,I227312,I226984);
DFFARX1 I_13213 (I227320,I2683,I226958,I226923,);
DFFARX1 I_13214 (I227312,I2683,I226958,I226941,);
nor I_13215 (I227365,I1860,I2444);
not I_13216 (I227382,I227365);
nor I_13217 (I226944,I227221,I227382);
nand I_13218 (I226929,I227238,I227382);
nor I_13219 (I226938,I226984,I227365);
DFFARX1 I_13220 (I227365,I2683,I226958,I226947,);
not I_13221 (I227485,I2690);
DFFARX1 I_13222 (I545124,I2683,I227485,I227511,);
nand I_13223 (I227519,I545115,I545130);
and I_13224 (I227536,I227519,I545136);
DFFARX1 I_13225 (I227536,I2683,I227485,I227562,);
nor I_13226 (I227453,I227562,I227511);
not I_13227 (I227584,I227562);
DFFARX1 I_13228 (I545121,I2683,I227485,I227610,);
nand I_13229 (I227618,I227610,I545115);
not I_13230 (I227635,I227618);
DFFARX1 I_13231 (I227635,I2683,I227485,I227661,);
not I_13232 (I227477,I227661);
nor I_13233 (I227683,I227511,I227618);
nor I_13234 (I227459,I227562,I227683);
DFFARX1 I_13235 (I545118,I2683,I227485,I227723,);
DFFARX1 I_13236 (I227723,I2683,I227485,I227740,);
not I_13237 (I227748,I227740);
not I_13238 (I227765,I227723);
nand I_13239 (I227462,I227765,I227584);
nand I_13240 (I227796,I545112,I545127);
and I_13241 (I227813,I227796,I545112);
DFFARX1 I_13242 (I227813,I2683,I227485,I227839,);
nor I_13243 (I227847,I227839,I227511);
DFFARX1 I_13244 (I227847,I2683,I227485,I227450,);
DFFARX1 I_13245 (I227839,I2683,I227485,I227468,);
nor I_13246 (I227892,I545133,I545127);
not I_13247 (I227909,I227892);
nor I_13248 (I227471,I227748,I227909);
nand I_13249 (I227456,I227765,I227909);
nor I_13250 (I227465,I227511,I227892);
DFFARX1 I_13251 (I227892,I2683,I227485,I227474,);
not I_13252 (I228012,I2690);
DFFARX1 I_13253 (I900446,I2683,I228012,I228038,);
nand I_13254 (I228046,I900461,I900446);
and I_13255 (I228063,I228046,I900464);
DFFARX1 I_13256 (I228063,I2683,I228012,I228089,);
nor I_13257 (I227980,I228089,I228038);
not I_13258 (I228111,I228089);
DFFARX1 I_13259 (I900470,I2683,I228012,I228137,);
nand I_13260 (I228145,I228137,I900452);
not I_13261 (I228162,I228145);
DFFARX1 I_13262 (I228162,I2683,I228012,I228188,);
not I_13263 (I228004,I228188);
nor I_13264 (I228210,I228038,I228145);
nor I_13265 (I227986,I228089,I228210);
DFFARX1 I_13266 (I900449,I2683,I228012,I228250,);
DFFARX1 I_13267 (I228250,I2683,I228012,I228267,);
not I_13268 (I228275,I228267);
not I_13269 (I228292,I228250);
nand I_13270 (I227989,I228292,I228111);
nand I_13271 (I228323,I900449,I900455);
and I_13272 (I228340,I228323,I900467);
DFFARX1 I_13273 (I228340,I2683,I228012,I228366,);
nor I_13274 (I228374,I228366,I228038);
DFFARX1 I_13275 (I228374,I2683,I228012,I227977,);
DFFARX1 I_13276 (I228366,I2683,I228012,I227995,);
nor I_13277 (I228419,I900458,I900455);
not I_13278 (I228436,I228419);
nor I_13279 (I227998,I228275,I228436);
nand I_13280 (I227983,I228292,I228436);
nor I_13281 (I227992,I228038,I228419);
DFFARX1 I_13282 (I228419,I2683,I228012,I228001,);
not I_13283 (I228539,I2690);
DFFARX1 I_13284 (I202715,I2683,I228539,I228565,);
nand I_13285 (I228573,I202715,I202721);
and I_13286 (I228590,I228573,I202739);
DFFARX1 I_13287 (I228590,I2683,I228539,I228616,);
nor I_13288 (I228507,I228616,I228565);
not I_13289 (I228638,I228616);
DFFARX1 I_13290 (I202727,I2683,I228539,I228664,);
nand I_13291 (I228672,I228664,I202724);
not I_13292 (I228689,I228672);
DFFARX1 I_13293 (I228689,I2683,I228539,I228715,);
not I_13294 (I228531,I228715);
nor I_13295 (I228737,I228565,I228672);
nor I_13296 (I228513,I228616,I228737);
DFFARX1 I_13297 (I202733,I2683,I228539,I228777,);
DFFARX1 I_13298 (I228777,I2683,I228539,I228794,);
not I_13299 (I228802,I228794);
not I_13300 (I228819,I228777);
nand I_13301 (I228516,I228819,I228638);
nand I_13302 (I228850,I202718,I202718);
and I_13303 (I228867,I228850,I202730);
DFFARX1 I_13304 (I228867,I2683,I228539,I228893,);
nor I_13305 (I228901,I228893,I228565);
DFFARX1 I_13306 (I228901,I2683,I228539,I228504,);
DFFARX1 I_13307 (I228893,I2683,I228539,I228522,);
nor I_13308 (I228946,I202736,I202718);
not I_13309 (I228963,I228946);
nor I_13310 (I228525,I228802,I228963);
nand I_13311 (I228510,I228819,I228963);
nor I_13312 (I228519,I228565,I228946);
DFFARX1 I_13313 (I228946,I2683,I228539,I228528,);
not I_13314 (I229066,I2690);
DFFARX1 I_13315 (I418720,I2683,I229066,I229092,);
nand I_13316 (I229100,I418720,I418732);
and I_13317 (I229117,I229100,I418717);
DFFARX1 I_13318 (I229117,I2683,I229066,I229143,);
nor I_13319 (I229034,I229143,I229092);
not I_13320 (I229165,I229143);
DFFARX1 I_13321 (I418741,I2683,I229066,I229191,);
nand I_13322 (I229199,I229191,I418738);
not I_13323 (I229216,I229199);
DFFARX1 I_13324 (I229216,I2683,I229066,I229242,);
not I_13325 (I229058,I229242);
nor I_13326 (I229264,I229092,I229199);
nor I_13327 (I229040,I229143,I229264);
DFFARX1 I_13328 (I418729,I2683,I229066,I229304,);
DFFARX1 I_13329 (I229304,I2683,I229066,I229321,);
not I_13330 (I229329,I229321);
not I_13331 (I229346,I229304);
nand I_13332 (I229043,I229346,I229165);
nand I_13333 (I229377,I418717,I418726);
and I_13334 (I229394,I229377,I418735);
DFFARX1 I_13335 (I229394,I2683,I229066,I229420,);
nor I_13336 (I229428,I229420,I229092);
DFFARX1 I_13337 (I229428,I2683,I229066,I229031,);
DFFARX1 I_13338 (I229420,I2683,I229066,I229049,);
nor I_13339 (I229473,I418723,I418726);
not I_13340 (I229490,I229473);
nor I_13341 (I229052,I229329,I229490);
nand I_13342 (I229037,I229346,I229490);
nor I_13343 (I229046,I229092,I229473);
DFFARX1 I_13344 (I229473,I2683,I229066,I229055,);
not I_13345 (I229593,I2690);
DFFARX1 I_13346 (I806320,I2683,I229593,I229619,);
nand I_13347 (I229627,I806317,I806320);
and I_13348 (I229644,I229627,I806329);
DFFARX1 I_13349 (I229644,I2683,I229593,I229670,);
nor I_13350 (I229561,I229670,I229619);
not I_13351 (I229692,I229670);
DFFARX1 I_13352 (I806317,I2683,I229593,I229718,);
nand I_13353 (I229726,I229718,I806335);
not I_13354 (I229743,I229726);
DFFARX1 I_13355 (I229743,I2683,I229593,I229769,);
not I_13356 (I229585,I229769);
nor I_13357 (I229791,I229619,I229726);
nor I_13358 (I229567,I229670,I229791);
DFFARX1 I_13359 (I806323,I2683,I229593,I229831,);
DFFARX1 I_13360 (I229831,I2683,I229593,I229848,);
not I_13361 (I229856,I229848);
not I_13362 (I229873,I229831);
nand I_13363 (I229570,I229873,I229692);
nand I_13364 (I229904,I806332,I806338);
and I_13365 (I229921,I229904,I806323);
DFFARX1 I_13366 (I229921,I2683,I229593,I229947,);
nor I_13367 (I229955,I229947,I229619);
DFFARX1 I_13368 (I229955,I2683,I229593,I229558,);
DFFARX1 I_13369 (I229947,I2683,I229593,I229576,);
nor I_13370 (I230000,I806326,I806338);
not I_13371 (I230017,I230000);
nor I_13372 (I229579,I229856,I230017);
nand I_13373 (I229564,I229873,I230017);
nor I_13374 (I229573,I229619,I230000);
DFFARX1 I_13375 (I230000,I2683,I229593,I229582,);
not I_13376 (I230120,I2690);
DFFARX1 I_13377 (I498884,I2683,I230120,I230146,);
nand I_13378 (I230154,I498875,I498890);
and I_13379 (I230171,I230154,I498896);
DFFARX1 I_13380 (I230171,I2683,I230120,I230197,);
nor I_13381 (I230088,I230197,I230146);
not I_13382 (I230219,I230197);
DFFARX1 I_13383 (I498881,I2683,I230120,I230245,);
nand I_13384 (I230253,I230245,I498875);
not I_13385 (I230270,I230253);
DFFARX1 I_13386 (I230270,I2683,I230120,I230296,);
not I_13387 (I230112,I230296);
nor I_13388 (I230318,I230146,I230253);
nor I_13389 (I230094,I230197,I230318);
DFFARX1 I_13390 (I498878,I2683,I230120,I230358,);
DFFARX1 I_13391 (I230358,I2683,I230120,I230375,);
not I_13392 (I230383,I230375);
not I_13393 (I230400,I230358);
nand I_13394 (I230097,I230400,I230219);
nand I_13395 (I230431,I498872,I498887);
and I_13396 (I230448,I230431,I498872);
DFFARX1 I_13397 (I230448,I2683,I230120,I230474,);
nor I_13398 (I230482,I230474,I230146);
DFFARX1 I_13399 (I230482,I2683,I230120,I230085,);
DFFARX1 I_13400 (I230474,I2683,I230120,I230103,);
nor I_13401 (I230527,I498893,I498887);
not I_13402 (I230544,I230527);
nor I_13403 (I230106,I230383,I230544);
nand I_13404 (I230091,I230400,I230544);
nor I_13405 (I230100,I230146,I230527);
DFFARX1 I_13406 (I230527,I2683,I230120,I230109,);
not I_13407 (I230647,I2690);
DFFARX1 I_13408 (I878482,I2683,I230647,I230673,);
nand I_13409 (I230681,I878497,I878482);
and I_13410 (I230698,I230681,I878500);
DFFARX1 I_13411 (I230698,I2683,I230647,I230724,);
nor I_13412 (I230615,I230724,I230673);
not I_13413 (I230746,I230724);
DFFARX1 I_13414 (I878506,I2683,I230647,I230772,);
nand I_13415 (I230780,I230772,I878488);
not I_13416 (I230797,I230780);
DFFARX1 I_13417 (I230797,I2683,I230647,I230823,);
not I_13418 (I230639,I230823);
nor I_13419 (I230845,I230673,I230780);
nor I_13420 (I230621,I230724,I230845);
DFFARX1 I_13421 (I878485,I2683,I230647,I230885,);
DFFARX1 I_13422 (I230885,I2683,I230647,I230902,);
not I_13423 (I230910,I230902);
not I_13424 (I230927,I230885);
nand I_13425 (I230624,I230927,I230746);
nand I_13426 (I230958,I878485,I878491);
and I_13427 (I230975,I230958,I878503);
DFFARX1 I_13428 (I230975,I2683,I230647,I231001,);
nor I_13429 (I231009,I231001,I230673);
DFFARX1 I_13430 (I231009,I2683,I230647,I230612,);
DFFARX1 I_13431 (I231001,I2683,I230647,I230630,);
nor I_13432 (I231054,I878494,I878491);
not I_13433 (I231071,I231054);
nor I_13434 (I230633,I230910,I231071);
nand I_13435 (I230618,I230927,I231071);
nor I_13436 (I230627,I230673,I231054);
DFFARX1 I_13437 (I231054,I2683,I230647,I230636,);
not I_13438 (I231174,I2690);
DFFARX1 I_13439 (I197955,I2683,I231174,I231200,);
nand I_13440 (I231208,I197955,I197961);
and I_13441 (I231225,I231208,I197979);
DFFARX1 I_13442 (I231225,I2683,I231174,I231251,);
nor I_13443 (I231142,I231251,I231200);
not I_13444 (I231273,I231251);
DFFARX1 I_13445 (I197967,I2683,I231174,I231299,);
nand I_13446 (I231307,I231299,I197964);
not I_13447 (I231324,I231307);
DFFARX1 I_13448 (I231324,I2683,I231174,I231350,);
not I_13449 (I231166,I231350);
nor I_13450 (I231372,I231200,I231307);
nor I_13451 (I231148,I231251,I231372);
DFFARX1 I_13452 (I197973,I2683,I231174,I231412,);
DFFARX1 I_13453 (I231412,I2683,I231174,I231429,);
not I_13454 (I231437,I231429);
not I_13455 (I231454,I231412);
nand I_13456 (I231151,I231454,I231273);
nand I_13457 (I231485,I197958,I197958);
and I_13458 (I231502,I231485,I197970);
DFFARX1 I_13459 (I231502,I2683,I231174,I231528,);
nor I_13460 (I231536,I231528,I231200);
DFFARX1 I_13461 (I231536,I2683,I231174,I231139,);
DFFARX1 I_13462 (I231528,I2683,I231174,I231157,);
nor I_13463 (I231581,I197976,I197958);
not I_13464 (I231598,I231581);
nor I_13465 (I231160,I231437,I231598);
nand I_13466 (I231145,I231454,I231598);
nor I_13467 (I231154,I231200,I231581);
DFFARX1 I_13468 (I231581,I2683,I231174,I231163,);
not I_13469 (I231701,I2690);
DFFARX1 I_13470 (I845536,I2683,I231701,I231727,);
nand I_13471 (I231735,I845551,I845536);
and I_13472 (I231752,I231735,I845554);
DFFARX1 I_13473 (I231752,I2683,I231701,I231778,);
nor I_13474 (I231669,I231778,I231727);
not I_13475 (I231800,I231778);
DFFARX1 I_13476 (I845560,I2683,I231701,I231826,);
nand I_13477 (I231834,I231826,I845542);
not I_13478 (I231851,I231834);
DFFARX1 I_13479 (I231851,I2683,I231701,I231877,);
not I_13480 (I231693,I231877);
nor I_13481 (I231899,I231727,I231834);
nor I_13482 (I231675,I231778,I231899);
DFFARX1 I_13483 (I845539,I2683,I231701,I231939,);
DFFARX1 I_13484 (I231939,I2683,I231701,I231956,);
not I_13485 (I231964,I231956);
not I_13486 (I231981,I231939);
nand I_13487 (I231678,I231981,I231800);
nand I_13488 (I232012,I845539,I845545);
and I_13489 (I232029,I232012,I845557);
DFFARX1 I_13490 (I232029,I2683,I231701,I232055,);
nor I_13491 (I232063,I232055,I231727);
DFFARX1 I_13492 (I232063,I2683,I231701,I231666,);
DFFARX1 I_13493 (I232055,I2683,I231701,I231684,);
nor I_13494 (I232108,I845548,I845545);
not I_13495 (I232125,I232108);
nor I_13496 (I231687,I231964,I232125);
nand I_13497 (I231672,I231981,I232125);
nor I_13498 (I231681,I231727,I232108);
DFFARX1 I_13499 (I232108,I2683,I231701,I231690,);
not I_13500 (I232228,I2690);
DFFARX1 I_13501 (I645449,I2683,I232228,I232254,);
nand I_13502 (I232262,I645452,I645446);
and I_13503 (I232279,I232262,I645458);
DFFARX1 I_13504 (I232279,I2683,I232228,I232305,);
nor I_13505 (I232196,I232305,I232254);
not I_13506 (I232327,I232305);
DFFARX1 I_13507 (I645461,I2683,I232228,I232353,);
nand I_13508 (I232361,I232353,I645452);
not I_13509 (I232378,I232361);
DFFARX1 I_13510 (I232378,I2683,I232228,I232404,);
not I_13511 (I232220,I232404);
nor I_13512 (I232426,I232254,I232361);
nor I_13513 (I232202,I232305,I232426);
DFFARX1 I_13514 (I645464,I2683,I232228,I232466,);
DFFARX1 I_13515 (I232466,I2683,I232228,I232483,);
not I_13516 (I232491,I232483);
not I_13517 (I232508,I232466);
nand I_13518 (I232205,I232508,I232327);
nand I_13519 (I232539,I645446,I645455);
and I_13520 (I232556,I232539,I645449);
DFFARX1 I_13521 (I232556,I2683,I232228,I232582,);
nor I_13522 (I232590,I232582,I232254);
DFFARX1 I_13523 (I232590,I2683,I232228,I232193,);
DFFARX1 I_13524 (I232582,I2683,I232228,I232211,);
nor I_13525 (I232635,I645467,I645455);
not I_13526 (I232652,I232635);
nor I_13527 (I232214,I232491,I232652);
nand I_13528 (I232199,I232508,I232652);
nor I_13529 (I232208,I232254,I232635);
DFFARX1 I_13530 (I232635,I2683,I232228,I232217,);
not I_13531 (I232755,I2690);
DFFARX1 I_13532 (I723870,I2683,I232755,I232781,);
nand I_13533 (I232789,I723867,I723885);
and I_13534 (I232806,I232789,I723876);
DFFARX1 I_13535 (I232806,I2683,I232755,I232832,);
nor I_13536 (I232723,I232832,I232781);
not I_13537 (I232854,I232832);
DFFARX1 I_13538 (I723891,I2683,I232755,I232880,);
nand I_13539 (I232888,I232880,I723873);
not I_13540 (I232905,I232888);
DFFARX1 I_13541 (I232905,I2683,I232755,I232931,);
not I_13542 (I232747,I232931);
nor I_13543 (I232953,I232781,I232888);
nor I_13544 (I232729,I232832,I232953);
DFFARX1 I_13545 (I723879,I2683,I232755,I232993,);
DFFARX1 I_13546 (I232993,I2683,I232755,I233010,);
not I_13547 (I233018,I233010);
not I_13548 (I233035,I232993);
nand I_13549 (I232732,I233035,I232854);
nand I_13550 (I233066,I723867,I723894);
and I_13551 (I233083,I233066,I723882);
DFFARX1 I_13552 (I233083,I2683,I232755,I233109,);
nor I_13553 (I233117,I233109,I232781);
DFFARX1 I_13554 (I233117,I2683,I232755,I232720,);
DFFARX1 I_13555 (I233109,I2683,I232755,I232738,);
nor I_13556 (I233162,I723888,I723894);
not I_13557 (I233179,I233162);
nor I_13558 (I232741,I233018,I233179);
nand I_13559 (I232726,I233035,I233179);
nor I_13560 (I232735,I232781,I233162);
DFFARX1 I_13561 (I233162,I2683,I232755,I232744,);
not I_13562 (I233282,I2690);
DFFARX1 I_13563 (I997837,I2683,I233282,I233308,);
nand I_13564 (I233316,I997834,I997825);
and I_13565 (I233333,I233316,I997822);
DFFARX1 I_13566 (I233333,I2683,I233282,I233359,);
nor I_13567 (I233250,I233359,I233308);
not I_13568 (I233381,I233359);
DFFARX1 I_13569 (I997831,I2683,I233282,I233407,);
nand I_13570 (I233415,I233407,I997840);
not I_13571 (I233432,I233415);
DFFARX1 I_13572 (I233432,I2683,I233282,I233458,);
not I_13573 (I233274,I233458);
nor I_13574 (I233480,I233308,I233415);
nor I_13575 (I233256,I233359,I233480);
DFFARX1 I_13576 (I997843,I2683,I233282,I233520,);
DFFARX1 I_13577 (I233520,I2683,I233282,I233537,);
not I_13578 (I233545,I233537);
not I_13579 (I233562,I233520);
nand I_13580 (I233259,I233562,I233381);
nand I_13581 (I233593,I997822,I997828);
and I_13582 (I233610,I233593,I997846);
DFFARX1 I_13583 (I233610,I2683,I233282,I233636,);
nor I_13584 (I233644,I233636,I233308);
DFFARX1 I_13585 (I233644,I2683,I233282,I233247,);
DFFARX1 I_13586 (I233636,I2683,I233282,I233265,);
nor I_13587 (I233689,I997825,I997828);
not I_13588 (I233706,I233689);
nor I_13589 (I233268,I233545,I233706);
nand I_13590 (I233253,I233562,I233706);
nor I_13591 (I233262,I233308,I233689);
DFFARX1 I_13592 (I233689,I2683,I233282,I233271,);
not I_13593 (I233809,I2690);
DFFARX1 I_13594 (I667056,I2683,I233809,I233835,);
nand I_13595 (I233843,I667059,I667053);
and I_13596 (I233860,I233843,I667065);
DFFARX1 I_13597 (I233860,I2683,I233809,I233886,);
nor I_13598 (I233777,I233886,I233835);
not I_13599 (I233908,I233886);
DFFARX1 I_13600 (I667068,I2683,I233809,I233934,);
nand I_13601 (I233942,I233934,I667059);
not I_13602 (I233959,I233942);
DFFARX1 I_13603 (I233959,I2683,I233809,I233985,);
not I_13604 (I233801,I233985);
nor I_13605 (I234007,I233835,I233942);
nor I_13606 (I233783,I233886,I234007);
DFFARX1 I_13607 (I667071,I2683,I233809,I234047,);
DFFARX1 I_13608 (I234047,I2683,I233809,I234064,);
not I_13609 (I234072,I234064);
not I_13610 (I234089,I234047);
nand I_13611 (I233786,I234089,I233908);
nand I_13612 (I234120,I667053,I667062);
and I_13613 (I234137,I234120,I667056);
DFFARX1 I_13614 (I234137,I2683,I233809,I234163,);
nor I_13615 (I234171,I234163,I233835);
DFFARX1 I_13616 (I234171,I2683,I233809,I233774,);
DFFARX1 I_13617 (I234163,I2683,I233809,I233792,);
nor I_13618 (I234216,I667074,I667062);
not I_13619 (I234233,I234216);
nor I_13620 (I233795,I234072,I234233);
nand I_13621 (I233780,I234089,I234233);
nor I_13622 (I233789,I233835,I234216);
DFFARX1 I_13623 (I234216,I2683,I233809,I233798,);
not I_13624 (I234336,I2690);
DFFARX1 I_13625 (I1044185,I2683,I234336,I234362,);
nand I_13626 (I234370,I1044164,I1044164);
and I_13627 (I234387,I234370,I1044191);
DFFARX1 I_13628 (I234387,I2683,I234336,I234413,);
nor I_13629 (I234304,I234413,I234362);
not I_13630 (I234435,I234413);
DFFARX1 I_13631 (I1044179,I2683,I234336,I234461,);
nand I_13632 (I234469,I234461,I1044182);
not I_13633 (I234486,I234469);
DFFARX1 I_13634 (I234486,I2683,I234336,I234512,);
not I_13635 (I234328,I234512);
nor I_13636 (I234534,I234362,I234469);
nor I_13637 (I234310,I234413,I234534);
DFFARX1 I_13638 (I1044173,I2683,I234336,I234574,);
DFFARX1 I_13639 (I234574,I2683,I234336,I234591,);
not I_13640 (I234599,I234591);
not I_13641 (I234616,I234574);
nand I_13642 (I234313,I234616,I234435);
nand I_13643 (I234647,I1044170,I1044167);
and I_13644 (I234664,I234647,I1044188);
DFFARX1 I_13645 (I234664,I2683,I234336,I234690,);
nor I_13646 (I234698,I234690,I234362);
DFFARX1 I_13647 (I234698,I2683,I234336,I234301,);
DFFARX1 I_13648 (I234690,I2683,I234336,I234319,);
nor I_13649 (I234743,I1044176,I1044167);
not I_13650 (I234760,I234743);
nor I_13651 (I234322,I234599,I234760);
nand I_13652 (I234307,I234616,I234760);
nor I_13653 (I234316,I234362,I234743);
DFFARX1 I_13654 (I234743,I2683,I234336,I234325,);
not I_13655 (I234863,I2690);
DFFARX1 I_13656 (I479813,I2683,I234863,I234889,);
nand I_13657 (I234897,I479798,I479801);
and I_13658 (I234914,I234897,I479816);
DFFARX1 I_13659 (I234914,I2683,I234863,I234940,);
nor I_13660 (I234831,I234940,I234889);
not I_13661 (I234962,I234940);
DFFARX1 I_13662 (I479810,I2683,I234863,I234988,);
nand I_13663 (I234996,I234988,I479801);
not I_13664 (I235013,I234996);
DFFARX1 I_13665 (I235013,I2683,I234863,I235039,);
not I_13666 (I234855,I235039);
nor I_13667 (I235061,I234889,I234996);
nor I_13668 (I234837,I234940,I235061);
DFFARX1 I_13669 (I479807,I2683,I234863,I235101,);
DFFARX1 I_13670 (I235101,I2683,I234863,I235118,);
not I_13671 (I235126,I235118);
not I_13672 (I235143,I235101);
nand I_13673 (I234840,I235143,I234962);
nand I_13674 (I235174,I479822,I479798);
and I_13675 (I235191,I235174,I479819);
DFFARX1 I_13676 (I235191,I2683,I234863,I235217,);
nor I_13677 (I235225,I235217,I234889);
DFFARX1 I_13678 (I235225,I2683,I234863,I234828,);
DFFARX1 I_13679 (I235217,I2683,I234863,I234846,);
nor I_13680 (I235270,I479804,I479798);
not I_13681 (I235287,I235270);
nor I_13682 (I234849,I235126,I235287);
nand I_13683 (I234834,I235143,I235287);
nor I_13684 (I234843,I234889,I235270);
DFFARX1 I_13685 (I235270,I2683,I234863,I234852,);
not I_13686 (I235390,I2690);
DFFARX1 I_13687 (I1078695,I2683,I235390,I235416,);
nand I_13688 (I235424,I1078674,I1078674);
and I_13689 (I235441,I235424,I1078701);
DFFARX1 I_13690 (I235441,I2683,I235390,I235467,);
nor I_13691 (I235358,I235467,I235416);
not I_13692 (I235489,I235467);
DFFARX1 I_13693 (I1078689,I2683,I235390,I235515,);
nand I_13694 (I235523,I235515,I1078692);
not I_13695 (I235540,I235523);
DFFARX1 I_13696 (I235540,I2683,I235390,I235566,);
not I_13697 (I235382,I235566);
nor I_13698 (I235588,I235416,I235523);
nor I_13699 (I235364,I235467,I235588);
DFFARX1 I_13700 (I1078683,I2683,I235390,I235628,);
DFFARX1 I_13701 (I235628,I2683,I235390,I235645,);
not I_13702 (I235653,I235645);
not I_13703 (I235670,I235628);
nand I_13704 (I235367,I235670,I235489);
nand I_13705 (I235701,I1078680,I1078677);
and I_13706 (I235718,I235701,I1078698);
DFFARX1 I_13707 (I235718,I2683,I235390,I235744,);
nor I_13708 (I235752,I235744,I235416);
DFFARX1 I_13709 (I235752,I2683,I235390,I235355,);
DFFARX1 I_13710 (I235744,I2683,I235390,I235373,);
nor I_13711 (I235797,I1078686,I1078677);
not I_13712 (I235814,I235797);
nor I_13713 (I235376,I235653,I235814);
nand I_13714 (I235361,I235670,I235814);
nor I_13715 (I235370,I235416,I235797);
DFFARX1 I_13716 (I235797,I2683,I235390,I235379,);
not I_13717 (I235917,I2690);
DFFARX1 I_13718 (I44819,I2683,I235917,I235943,);
nand I_13719 (I235951,I44843,I44822);
and I_13720 (I235968,I235951,I44819);
DFFARX1 I_13721 (I235968,I2683,I235917,I235994,);
nor I_13722 (I235885,I235994,I235943);
not I_13723 (I236016,I235994);
DFFARX1 I_13724 (I44825,I2683,I235917,I236042,);
nand I_13725 (I236050,I236042,I44834);
not I_13726 (I236067,I236050);
DFFARX1 I_13727 (I236067,I2683,I235917,I236093,);
not I_13728 (I235909,I236093);
nor I_13729 (I236115,I235943,I236050);
nor I_13730 (I235891,I235994,I236115);
DFFARX1 I_13731 (I44828,I2683,I235917,I236155,);
DFFARX1 I_13732 (I236155,I2683,I235917,I236172,);
not I_13733 (I236180,I236172);
not I_13734 (I236197,I236155);
nand I_13735 (I235894,I236197,I236016);
nand I_13736 (I236228,I44840,I44822);
and I_13737 (I236245,I236228,I44831);
DFFARX1 I_13738 (I236245,I2683,I235917,I236271,);
nor I_13739 (I236279,I236271,I235943);
DFFARX1 I_13740 (I236279,I2683,I235917,I235882,);
DFFARX1 I_13741 (I236271,I2683,I235917,I235900,);
nor I_13742 (I236324,I44837,I44822);
not I_13743 (I236341,I236324);
nor I_13744 (I235903,I236180,I236341);
nand I_13745 (I235888,I236197,I236341);
nor I_13746 (I235897,I235943,I236324);
DFFARX1 I_13747 (I236324,I2683,I235917,I235906,);
not I_13748 (I236444,I2690);
DFFARX1 I_13749 (I660732,I2683,I236444,I236470,);
nand I_13750 (I236478,I660735,I660729);
and I_13751 (I236495,I236478,I660741);
DFFARX1 I_13752 (I236495,I2683,I236444,I236521,);
nor I_13753 (I236412,I236521,I236470);
not I_13754 (I236543,I236521);
DFFARX1 I_13755 (I660744,I2683,I236444,I236569,);
nand I_13756 (I236577,I236569,I660735);
not I_13757 (I236594,I236577);
DFFARX1 I_13758 (I236594,I2683,I236444,I236620,);
not I_13759 (I236436,I236620);
nor I_13760 (I236642,I236470,I236577);
nor I_13761 (I236418,I236521,I236642);
DFFARX1 I_13762 (I660747,I2683,I236444,I236682,);
DFFARX1 I_13763 (I236682,I2683,I236444,I236699,);
not I_13764 (I236707,I236699);
not I_13765 (I236724,I236682);
nand I_13766 (I236421,I236724,I236543);
nand I_13767 (I236755,I660729,I660738);
and I_13768 (I236772,I236755,I660732);
DFFARX1 I_13769 (I236772,I2683,I236444,I236798,);
nor I_13770 (I236806,I236798,I236470);
DFFARX1 I_13771 (I236806,I2683,I236444,I236409,);
DFFARX1 I_13772 (I236798,I2683,I236444,I236427,);
nor I_13773 (I236851,I660750,I660738);
not I_13774 (I236868,I236851);
nor I_13775 (I236430,I236707,I236868);
nand I_13776 (I236415,I236724,I236868);
nor I_13777 (I236424,I236470,I236851);
DFFARX1 I_13778 (I236851,I2683,I236444,I236433,);
not I_13779 (I236971,I2690);
DFFARX1 I_13780 (I369854,I2683,I236971,I236997,);
nand I_13781 (I237005,I369866,I369845);
and I_13782 (I237022,I237005,I369869);
DFFARX1 I_13783 (I237022,I2683,I236971,I237048,);
nor I_13784 (I236939,I237048,I236997);
not I_13785 (I237070,I237048);
DFFARX1 I_13786 (I369860,I2683,I236971,I237096,);
nand I_13787 (I237104,I237096,I369842);
not I_13788 (I237121,I237104);
DFFARX1 I_13789 (I237121,I2683,I236971,I237147,);
not I_13790 (I236963,I237147);
nor I_13791 (I237169,I236997,I237104);
nor I_13792 (I236945,I237048,I237169);
DFFARX1 I_13793 (I369857,I2683,I236971,I237209,);
DFFARX1 I_13794 (I237209,I2683,I236971,I237226,);
not I_13795 (I237234,I237226);
not I_13796 (I237251,I237209);
nand I_13797 (I236948,I237251,I237070);
nand I_13798 (I237282,I369842,I369848);
and I_13799 (I237299,I237282,I369851);
DFFARX1 I_13800 (I237299,I2683,I236971,I237325,);
nor I_13801 (I237333,I237325,I236997);
DFFARX1 I_13802 (I237333,I2683,I236971,I236936,);
DFFARX1 I_13803 (I237325,I2683,I236971,I236954,);
nor I_13804 (I237378,I369863,I369848);
not I_13805 (I237395,I237378);
nor I_13806 (I236957,I237234,I237395);
nand I_13807 (I236942,I237251,I237395);
nor I_13808 (I236951,I236997,I237378);
DFFARX1 I_13809 (I237378,I2683,I236971,I236960,);
not I_13810 (I237498,I2690);
DFFARX1 I_13811 (I389982,I2683,I237498,I237524,);
nand I_13812 (I237532,I389994,I389973);
and I_13813 (I237549,I237532,I389997);
DFFARX1 I_13814 (I237549,I2683,I237498,I237575,);
nor I_13815 (I237466,I237575,I237524);
not I_13816 (I237597,I237575);
DFFARX1 I_13817 (I389988,I2683,I237498,I237623,);
nand I_13818 (I237631,I237623,I389970);
not I_13819 (I237648,I237631);
DFFARX1 I_13820 (I237648,I2683,I237498,I237674,);
not I_13821 (I237490,I237674);
nor I_13822 (I237696,I237524,I237631);
nor I_13823 (I237472,I237575,I237696);
DFFARX1 I_13824 (I389985,I2683,I237498,I237736,);
DFFARX1 I_13825 (I237736,I2683,I237498,I237753,);
not I_13826 (I237761,I237753);
not I_13827 (I237778,I237736);
nand I_13828 (I237475,I237778,I237597);
nand I_13829 (I237809,I389970,I389976);
and I_13830 (I237826,I237809,I389979);
DFFARX1 I_13831 (I237826,I2683,I237498,I237852,);
nor I_13832 (I237860,I237852,I237524);
DFFARX1 I_13833 (I237860,I2683,I237498,I237463,);
DFFARX1 I_13834 (I237852,I2683,I237498,I237481,);
nor I_13835 (I237905,I389991,I389976);
not I_13836 (I237922,I237905);
nor I_13837 (I237484,I237761,I237922);
nand I_13838 (I237469,I237778,I237922);
nor I_13839 (I237478,I237524,I237905);
DFFARX1 I_13840 (I237905,I2683,I237498,I237487,);
not I_13841 (I238025,I2690);
DFFARX1 I_13842 (I169395,I2683,I238025,I238051,);
nand I_13843 (I238059,I169395,I169401);
and I_13844 (I238076,I238059,I169419);
DFFARX1 I_13845 (I238076,I2683,I238025,I238102,);
nor I_13846 (I237993,I238102,I238051);
not I_13847 (I238124,I238102);
DFFARX1 I_13848 (I169407,I2683,I238025,I238150,);
nand I_13849 (I238158,I238150,I169404);
not I_13850 (I238175,I238158);
DFFARX1 I_13851 (I238175,I2683,I238025,I238201,);
not I_13852 (I238017,I238201);
nor I_13853 (I238223,I238051,I238158);
nor I_13854 (I237999,I238102,I238223);
DFFARX1 I_13855 (I169413,I2683,I238025,I238263,);
DFFARX1 I_13856 (I238263,I2683,I238025,I238280,);
not I_13857 (I238288,I238280);
not I_13858 (I238305,I238263);
nand I_13859 (I238002,I238305,I238124);
nand I_13860 (I238336,I169398,I169398);
and I_13861 (I238353,I238336,I169410);
DFFARX1 I_13862 (I238353,I2683,I238025,I238379,);
nor I_13863 (I238387,I238379,I238051);
DFFARX1 I_13864 (I238387,I2683,I238025,I237990,);
DFFARX1 I_13865 (I238379,I2683,I238025,I238008,);
nor I_13866 (I238432,I169416,I169398);
not I_13867 (I238449,I238432);
nor I_13868 (I238011,I238288,I238449);
nand I_13869 (I237996,I238305,I238449);
nor I_13870 (I238005,I238051,I238432);
DFFARX1 I_13871 (I238432,I2683,I238025,I238014,);
not I_13872 (I238552,I2690);
DFFARX1 I_13873 (I151545,I2683,I238552,I238578,);
nand I_13874 (I238586,I151545,I151551);
and I_13875 (I238603,I238586,I151569);
DFFARX1 I_13876 (I238603,I2683,I238552,I238629,);
nor I_13877 (I238520,I238629,I238578);
not I_13878 (I238651,I238629);
DFFARX1 I_13879 (I151557,I2683,I238552,I238677,);
nand I_13880 (I238685,I238677,I151554);
not I_13881 (I238702,I238685);
DFFARX1 I_13882 (I238702,I2683,I238552,I238728,);
not I_13883 (I238544,I238728);
nor I_13884 (I238750,I238578,I238685);
nor I_13885 (I238526,I238629,I238750);
DFFARX1 I_13886 (I151563,I2683,I238552,I238790,);
DFFARX1 I_13887 (I238790,I2683,I238552,I238807,);
not I_13888 (I238815,I238807);
not I_13889 (I238832,I238790);
nand I_13890 (I238529,I238832,I238651);
nand I_13891 (I238863,I151548,I151548);
and I_13892 (I238880,I238863,I151560);
DFFARX1 I_13893 (I238880,I2683,I238552,I238906,);
nor I_13894 (I238914,I238906,I238578);
DFFARX1 I_13895 (I238914,I2683,I238552,I238517,);
DFFARX1 I_13896 (I238906,I2683,I238552,I238535,);
nor I_13897 (I238959,I151566,I151548);
not I_13898 (I238976,I238959);
nor I_13899 (I238538,I238815,I238976);
nand I_13900 (I238523,I238832,I238976);
nor I_13901 (I238532,I238578,I238959);
DFFARX1 I_13902 (I238959,I2683,I238552,I238541,);
not I_13903 (I239079,I2690);
DFFARX1 I_13904 (I805198,I2683,I239079,I239105,);
nand I_13905 (I239113,I805195,I805198);
and I_13906 (I239130,I239113,I805207);
DFFARX1 I_13907 (I239130,I2683,I239079,I239156,);
nor I_13908 (I239047,I239156,I239105);
not I_13909 (I239178,I239156);
DFFARX1 I_13910 (I805195,I2683,I239079,I239204,);
nand I_13911 (I239212,I239204,I805213);
not I_13912 (I239229,I239212);
DFFARX1 I_13913 (I239229,I2683,I239079,I239255,);
not I_13914 (I239071,I239255);
nor I_13915 (I239277,I239105,I239212);
nor I_13916 (I239053,I239156,I239277);
DFFARX1 I_13917 (I805201,I2683,I239079,I239317,);
DFFARX1 I_13918 (I239317,I2683,I239079,I239334,);
not I_13919 (I239342,I239334);
not I_13920 (I239359,I239317);
nand I_13921 (I239056,I239359,I239178);
nand I_13922 (I239390,I805210,I805216);
and I_13923 (I239407,I239390,I805201);
DFFARX1 I_13924 (I239407,I2683,I239079,I239433,);
nor I_13925 (I239441,I239433,I239105);
DFFARX1 I_13926 (I239441,I2683,I239079,I239044,);
DFFARX1 I_13927 (I239433,I2683,I239079,I239062,);
nor I_13928 (I239486,I805204,I805216);
not I_13929 (I239503,I239486);
nor I_13930 (I239065,I239342,I239503);
nand I_13931 (I239050,I239359,I239503);
nor I_13932 (I239059,I239105,I239486);
DFFARX1 I_13933 (I239486,I2683,I239079,I239068,);
not I_13934 (I239606,I2690);
DFFARX1 I_13935 (I589630,I2683,I239606,I239632,);
nand I_13936 (I239640,I589621,I589636);
and I_13937 (I239657,I239640,I589642);
DFFARX1 I_13938 (I239657,I2683,I239606,I239683,);
nor I_13939 (I239574,I239683,I239632);
not I_13940 (I239705,I239683);
DFFARX1 I_13941 (I589627,I2683,I239606,I239731,);
nand I_13942 (I239739,I239731,I589621);
not I_13943 (I239756,I239739);
DFFARX1 I_13944 (I239756,I2683,I239606,I239782,);
not I_13945 (I239598,I239782);
nor I_13946 (I239804,I239632,I239739);
nor I_13947 (I239580,I239683,I239804);
DFFARX1 I_13948 (I589624,I2683,I239606,I239844,);
DFFARX1 I_13949 (I239844,I2683,I239606,I239861,);
not I_13950 (I239869,I239861);
not I_13951 (I239886,I239844);
nand I_13952 (I239583,I239886,I239705);
nand I_13953 (I239917,I589618,I589633);
and I_13954 (I239934,I239917,I589618);
DFFARX1 I_13955 (I239934,I2683,I239606,I239960,);
nor I_13956 (I239968,I239960,I239632);
DFFARX1 I_13957 (I239968,I2683,I239606,I239571,);
DFFARX1 I_13958 (I239960,I2683,I239606,I239589,);
nor I_13959 (I240013,I589639,I589633);
not I_13960 (I240030,I240013);
nor I_13961 (I239592,I239869,I240030);
nand I_13962 (I239577,I239886,I240030);
nor I_13963 (I239586,I239632,I240013);
DFFARX1 I_13964 (I240013,I2683,I239606,I239595,);
not I_13965 (I240133,I2690);
DFFARX1 I_13966 (I105427,I2683,I240133,I240159,);
nand I_13967 (I240167,I105439,I105448);
and I_13968 (I240184,I240167,I105427);
DFFARX1 I_13969 (I240184,I2683,I240133,I240210,);
nor I_13970 (I240101,I240210,I240159);
not I_13971 (I240232,I240210);
DFFARX1 I_13972 (I105442,I2683,I240133,I240258,);
nand I_13973 (I240266,I240258,I105430);
not I_13974 (I240283,I240266);
DFFARX1 I_13975 (I240283,I2683,I240133,I240309,);
not I_13976 (I240125,I240309);
nor I_13977 (I240331,I240159,I240266);
nor I_13978 (I240107,I240210,I240331);
DFFARX1 I_13979 (I105433,I2683,I240133,I240371,);
DFFARX1 I_13980 (I240371,I2683,I240133,I240388,);
not I_13981 (I240396,I240388);
not I_13982 (I240413,I240371);
nand I_13983 (I240110,I240413,I240232);
nand I_13984 (I240444,I105424,I105424);
and I_13985 (I240461,I240444,I105436);
DFFARX1 I_13986 (I240461,I2683,I240133,I240487,);
nor I_13987 (I240495,I240487,I240159);
DFFARX1 I_13988 (I240495,I2683,I240133,I240098,);
DFFARX1 I_13989 (I240487,I2683,I240133,I240116,);
nor I_13990 (I240540,I105445,I105424);
not I_13991 (I240557,I240540);
nor I_13992 (I240119,I240396,I240557);
nand I_13993 (I240104,I240413,I240557);
nor I_13994 (I240113,I240159,I240540);
DFFARX1 I_13995 (I240540,I2683,I240133,I240122,);
not I_13996 (I240660,I2690);
DFFARX1 I_13997 (I494841,I2683,I240660,I240686,);
nand I_13998 (I240694,I494826,I494829);
and I_13999 (I240711,I240694,I494844);
DFFARX1 I_14000 (I240711,I2683,I240660,I240737,);
nor I_14001 (I240628,I240737,I240686);
not I_14002 (I240759,I240737);
DFFARX1 I_14003 (I494838,I2683,I240660,I240785,);
nand I_14004 (I240793,I240785,I494829);
not I_14005 (I240810,I240793);
DFFARX1 I_14006 (I240810,I2683,I240660,I240836,);
not I_14007 (I240652,I240836);
nor I_14008 (I240858,I240686,I240793);
nor I_14009 (I240634,I240737,I240858);
DFFARX1 I_14010 (I494835,I2683,I240660,I240898,);
DFFARX1 I_14011 (I240898,I2683,I240660,I240915,);
not I_14012 (I240923,I240915);
not I_14013 (I240940,I240898);
nand I_14014 (I240637,I240940,I240759);
nand I_14015 (I240971,I494850,I494826);
and I_14016 (I240988,I240971,I494847);
DFFARX1 I_14017 (I240988,I2683,I240660,I241014,);
nor I_14018 (I241022,I241014,I240686);
DFFARX1 I_14019 (I241022,I2683,I240660,I240625,);
DFFARX1 I_14020 (I241014,I2683,I240660,I240643,);
nor I_14021 (I241067,I494832,I494826);
not I_14022 (I241084,I241067);
nor I_14023 (I240646,I240923,I241084);
nand I_14024 (I240631,I240940,I241084);
nor I_14025 (I240640,I240686,I241067);
DFFARX1 I_14026 (I241067,I2683,I240660,I240649,);
not I_14027 (I241187,I2690);
DFFARX1 I_14028 (I640706,I2683,I241187,I241213,);
nand I_14029 (I241221,I640709,I640703);
and I_14030 (I241238,I241221,I640715);
DFFARX1 I_14031 (I241238,I2683,I241187,I241264,);
nor I_14032 (I241155,I241264,I241213);
not I_14033 (I241286,I241264);
DFFARX1 I_14034 (I640718,I2683,I241187,I241312,);
nand I_14035 (I241320,I241312,I640709);
not I_14036 (I241337,I241320);
DFFARX1 I_14037 (I241337,I2683,I241187,I241363,);
not I_14038 (I241179,I241363);
nor I_14039 (I241385,I241213,I241320);
nor I_14040 (I241161,I241264,I241385);
DFFARX1 I_14041 (I640721,I2683,I241187,I241425,);
DFFARX1 I_14042 (I241425,I2683,I241187,I241442,);
not I_14043 (I241450,I241442);
not I_14044 (I241467,I241425);
nand I_14045 (I241164,I241467,I241286);
nand I_14046 (I241498,I640703,I640712);
and I_14047 (I241515,I241498,I640706);
DFFARX1 I_14048 (I241515,I2683,I241187,I241541,);
nor I_14049 (I241549,I241541,I241213);
DFFARX1 I_14050 (I241549,I2683,I241187,I241152,);
DFFARX1 I_14051 (I241541,I2683,I241187,I241170,);
nor I_14052 (I241594,I640724,I640712);
not I_14053 (I241611,I241594);
nor I_14054 (I241173,I241450,I241611);
nand I_14055 (I241158,I241467,I241611);
nor I_14056 (I241167,I241213,I241594);
DFFARX1 I_14057 (I241594,I2683,I241187,I241176,);
not I_14058 (I241714,I2690);
DFFARX1 I_14059 (I325790,I2683,I241714,I241740,);
nand I_14060 (I241748,I325802,I325781);
and I_14061 (I241765,I241748,I325805);
DFFARX1 I_14062 (I241765,I2683,I241714,I241791,);
nor I_14063 (I241682,I241791,I241740);
not I_14064 (I241813,I241791);
DFFARX1 I_14065 (I325796,I2683,I241714,I241839,);
nand I_14066 (I241847,I241839,I325778);
not I_14067 (I241864,I241847);
DFFARX1 I_14068 (I241864,I2683,I241714,I241890,);
not I_14069 (I241706,I241890);
nor I_14070 (I241912,I241740,I241847);
nor I_14071 (I241688,I241791,I241912);
DFFARX1 I_14072 (I325793,I2683,I241714,I241952,);
DFFARX1 I_14073 (I241952,I2683,I241714,I241969,);
not I_14074 (I241977,I241969);
not I_14075 (I241994,I241952);
nand I_14076 (I241691,I241994,I241813);
nand I_14077 (I242025,I325778,I325784);
and I_14078 (I242042,I242025,I325787);
DFFARX1 I_14079 (I242042,I2683,I241714,I242068,);
nor I_14080 (I242076,I242068,I241740);
DFFARX1 I_14081 (I242076,I2683,I241714,I241679,);
DFFARX1 I_14082 (I242068,I2683,I241714,I241697,);
nor I_14083 (I242121,I325799,I325784);
not I_14084 (I242138,I242121);
nor I_14085 (I241700,I241977,I242138);
nand I_14086 (I241685,I241994,I242138);
nor I_14087 (I241694,I241740,I242121);
DFFARX1 I_14088 (I242121,I2683,I241714,I241703,);
not I_14089 (I242241,I2690);
DFFARX1 I_14090 (I391614,I2683,I242241,I242267,);
nand I_14091 (I242275,I391626,I391605);
and I_14092 (I242292,I242275,I391629);
DFFARX1 I_14093 (I242292,I2683,I242241,I242318,);
nor I_14094 (I242209,I242318,I242267);
not I_14095 (I242340,I242318);
DFFARX1 I_14096 (I391620,I2683,I242241,I242366,);
nand I_14097 (I242374,I242366,I391602);
not I_14098 (I242391,I242374);
DFFARX1 I_14099 (I242391,I2683,I242241,I242417,);
not I_14100 (I242233,I242417);
nor I_14101 (I242439,I242267,I242374);
nor I_14102 (I242215,I242318,I242439);
DFFARX1 I_14103 (I391617,I2683,I242241,I242479,);
DFFARX1 I_14104 (I242479,I2683,I242241,I242496,);
not I_14105 (I242504,I242496);
not I_14106 (I242521,I242479);
nand I_14107 (I242218,I242521,I242340);
nand I_14108 (I242552,I391602,I391608);
and I_14109 (I242569,I242552,I391611);
DFFARX1 I_14110 (I242569,I2683,I242241,I242595,);
nor I_14111 (I242603,I242595,I242267);
DFFARX1 I_14112 (I242603,I2683,I242241,I242206,);
DFFARX1 I_14113 (I242595,I2683,I242241,I242224,);
nor I_14114 (I242648,I391623,I391608);
not I_14115 (I242665,I242648);
nor I_14116 (I242227,I242504,I242665);
nand I_14117 (I242212,I242521,I242665);
nor I_14118 (I242221,I242267,I242648);
DFFARX1 I_14119 (I242648,I2683,I242241,I242230,);
not I_14120 (I242768,I2690);
DFFARX1 I_14121 (I696041,I2683,I242768,I242794,);
nand I_14122 (I242802,I696044,I696038);
and I_14123 (I242819,I242802,I696050);
DFFARX1 I_14124 (I242819,I2683,I242768,I242845,);
nor I_14125 (I242736,I242845,I242794);
not I_14126 (I242867,I242845);
DFFARX1 I_14127 (I696053,I2683,I242768,I242893,);
nand I_14128 (I242901,I242893,I696044);
not I_14129 (I242918,I242901);
DFFARX1 I_14130 (I242918,I2683,I242768,I242944,);
not I_14131 (I242760,I242944);
nor I_14132 (I242966,I242794,I242901);
nor I_14133 (I242742,I242845,I242966);
DFFARX1 I_14134 (I696056,I2683,I242768,I243006,);
DFFARX1 I_14135 (I243006,I2683,I242768,I243023,);
not I_14136 (I243031,I243023);
not I_14137 (I243048,I243006);
nand I_14138 (I242745,I243048,I242867);
nand I_14139 (I243079,I696038,I696047);
and I_14140 (I243096,I243079,I696041);
DFFARX1 I_14141 (I243096,I2683,I242768,I243122,);
nor I_14142 (I243130,I243122,I242794);
DFFARX1 I_14143 (I243130,I2683,I242768,I242733,);
DFFARX1 I_14144 (I243122,I2683,I242768,I242751,);
nor I_14145 (I243175,I696059,I696047);
not I_14146 (I243192,I243175);
nor I_14147 (I242754,I243031,I243192);
nand I_14148 (I242739,I243048,I243192);
nor I_14149 (I242748,I242794,I243175);
DFFARX1 I_14150 (I243175,I2683,I242768,I242757,);
not I_14151 (I243295,I2690);
DFFARX1 I_14152 (I75915,I2683,I243295,I243321,);
nand I_14153 (I243329,I75927,I75936);
and I_14154 (I243346,I243329,I75915);
DFFARX1 I_14155 (I243346,I2683,I243295,I243372,);
nor I_14156 (I243263,I243372,I243321);
not I_14157 (I243394,I243372);
DFFARX1 I_14158 (I75930,I2683,I243295,I243420,);
nand I_14159 (I243428,I243420,I75918);
not I_14160 (I243445,I243428);
DFFARX1 I_14161 (I243445,I2683,I243295,I243471,);
not I_14162 (I243287,I243471);
nor I_14163 (I243493,I243321,I243428);
nor I_14164 (I243269,I243372,I243493);
DFFARX1 I_14165 (I75921,I2683,I243295,I243533,);
DFFARX1 I_14166 (I243533,I2683,I243295,I243550,);
not I_14167 (I243558,I243550);
not I_14168 (I243575,I243533);
nand I_14169 (I243272,I243575,I243394);
nand I_14170 (I243606,I75912,I75912);
and I_14171 (I243623,I243606,I75924);
DFFARX1 I_14172 (I243623,I2683,I243295,I243649,);
nor I_14173 (I243657,I243649,I243321);
DFFARX1 I_14174 (I243657,I2683,I243295,I243260,);
DFFARX1 I_14175 (I243649,I2683,I243295,I243278,);
nor I_14176 (I243702,I75933,I75912);
not I_14177 (I243719,I243702);
nor I_14178 (I243281,I243558,I243719);
nand I_14179 (I243266,I243575,I243719);
nor I_14180 (I243275,I243321,I243702);
DFFARX1 I_14181 (I243702,I2683,I243295,I243284,);
not I_14182 (I243822,I2690);
DFFARX1 I_14183 (I537610,I2683,I243822,I243848,);
nand I_14184 (I243856,I537601,I537616);
and I_14185 (I243873,I243856,I537622);
DFFARX1 I_14186 (I243873,I2683,I243822,I243899,);
nor I_14187 (I243790,I243899,I243848);
not I_14188 (I243921,I243899);
DFFARX1 I_14189 (I537607,I2683,I243822,I243947,);
nand I_14190 (I243955,I243947,I537601);
not I_14191 (I243972,I243955);
DFFARX1 I_14192 (I243972,I2683,I243822,I243998,);
not I_14193 (I243814,I243998);
nor I_14194 (I244020,I243848,I243955);
nor I_14195 (I243796,I243899,I244020);
DFFARX1 I_14196 (I537604,I2683,I243822,I244060,);
DFFARX1 I_14197 (I244060,I2683,I243822,I244077,);
not I_14198 (I244085,I244077);
not I_14199 (I244102,I244060);
nand I_14200 (I243799,I244102,I243921);
nand I_14201 (I244133,I537598,I537613);
and I_14202 (I244150,I244133,I537598);
DFFARX1 I_14203 (I244150,I2683,I243822,I244176,);
nor I_14204 (I244184,I244176,I243848);
DFFARX1 I_14205 (I244184,I2683,I243822,I243787,);
DFFARX1 I_14206 (I244176,I2683,I243822,I243805,);
nor I_14207 (I244229,I537619,I537613);
not I_14208 (I244246,I244229);
nor I_14209 (I243808,I244085,I244246);
nand I_14210 (I243793,I244102,I244246);
nor I_14211 (I243802,I243848,I244229);
DFFARX1 I_14212 (I244229,I2683,I243822,I243811,);
not I_14213 (I244349,I2690);
DFFARX1 I_14214 (I162850,I2683,I244349,I244375,);
nand I_14215 (I244383,I162850,I162856);
and I_14216 (I244400,I244383,I162874);
DFFARX1 I_14217 (I244400,I2683,I244349,I244426,);
nor I_14218 (I244317,I244426,I244375);
not I_14219 (I244448,I244426);
DFFARX1 I_14220 (I162862,I2683,I244349,I244474,);
nand I_14221 (I244482,I244474,I162859);
not I_14222 (I244499,I244482);
DFFARX1 I_14223 (I244499,I2683,I244349,I244525,);
not I_14224 (I244341,I244525);
nor I_14225 (I244547,I244375,I244482);
nor I_14226 (I244323,I244426,I244547);
DFFARX1 I_14227 (I162868,I2683,I244349,I244587,);
DFFARX1 I_14228 (I244587,I2683,I244349,I244604,);
not I_14229 (I244612,I244604);
not I_14230 (I244629,I244587);
nand I_14231 (I244326,I244629,I244448);
nand I_14232 (I244660,I162853,I162853);
and I_14233 (I244677,I244660,I162865);
DFFARX1 I_14234 (I244677,I2683,I244349,I244703,);
nor I_14235 (I244711,I244703,I244375);
DFFARX1 I_14236 (I244711,I2683,I244349,I244314,);
DFFARX1 I_14237 (I244703,I2683,I244349,I244332,);
nor I_14238 (I244756,I162871,I162853);
not I_14239 (I244773,I244756);
nor I_14240 (I244335,I244612,I244773);
nand I_14241 (I244320,I244629,I244773);
nor I_14242 (I244329,I244375,I244756);
DFFARX1 I_14243 (I244756,I2683,I244349,I244338,);
not I_14244 (I244876,I2690);
DFFARX1 I_14245 (I564198,I2683,I244876,I244902,);
nand I_14246 (I244910,I564189,I564204);
and I_14247 (I244927,I244910,I564210);
DFFARX1 I_14248 (I244927,I2683,I244876,I244953,);
nor I_14249 (I244844,I244953,I244902);
not I_14250 (I244975,I244953);
DFFARX1 I_14251 (I564195,I2683,I244876,I245001,);
nand I_14252 (I245009,I245001,I564189);
not I_14253 (I245026,I245009);
DFFARX1 I_14254 (I245026,I2683,I244876,I245052,);
not I_14255 (I244868,I245052);
nor I_14256 (I245074,I244902,I245009);
nor I_14257 (I244850,I244953,I245074);
DFFARX1 I_14258 (I564192,I2683,I244876,I245114,);
DFFARX1 I_14259 (I245114,I2683,I244876,I245131,);
not I_14260 (I245139,I245131);
not I_14261 (I245156,I245114);
nand I_14262 (I244853,I245156,I244975);
nand I_14263 (I245187,I564186,I564201);
and I_14264 (I245204,I245187,I564186);
DFFARX1 I_14265 (I245204,I2683,I244876,I245230,);
nor I_14266 (I245238,I245230,I244902);
DFFARX1 I_14267 (I245238,I2683,I244876,I244841,);
DFFARX1 I_14268 (I245230,I2683,I244876,I244859,);
nor I_14269 (I245283,I564207,I564201);
not I_14270 (I245300,I245283);
nor I_14271 (I244862,I245139,I245300);
nand I_14272 (I244847,I245156,I245300);
nor I_14273 (I244856,I244902,I245283);
DFFARX1 I_14274 (I245283,I2683,I244876,I244865,);
not I_14275 (I245403,I2690);
DFFARX1 I_14276 (I85401,I2683,I245403,I245429,);
nand I_14277 (I245437,I85413,I85422);
and I_14278 (I245454,I245437,I85401);
DFFARX1 I_14279 (I245454,I2683,I245403,I245480,);
nor I_14280 (I245371,I245480,I245429);
not I_14281 (I245502,I245480);
DFFARX1 I_14282 (I85416,I2683,I245403,I245528,);
nand I_14283 (I245536,I245528,I85404);
not I_14284 (I245553,I245536);
DFFARX1 I_14285 (I245553,I2683,I245403,I245579,);
not I_14286 (I245395,I245579);
nor I_14287 (I245601,I245429,I245536);
nor I_14288 (I245377,I245480,I245601);
DFFARX1 I_14289 (I85407,I2683,I245403,I245641,);
DFFARX1 I_14290 (I245641,I2683,I245403,I245658,);
not I_14291 (I245666,I245658);
not I_14292 (I245683,I245641);
nand I_14293 (I245380,I245683,I245502);
nand I_14294 (I245714,I85398,I85398);
and I_14295 (I245731,I245714,I85410);
DFFARX1 I_14296 (I245731,I2683,I245403,I245757,);
nor I_14297 (I245765,I245757,I245429);
DFFARX1 I_14298 (I245765,I2683,I245403,I245368,);
DFFARX1 I_14299 (I245757,I2683,I245403,I245386,);
nor I_14300 (I245810,I85419,I85398);
not I_14301 (I245827,I245810);
nor I_14302 (I245389,I245666,I245827);
nand I_14303 (I245374,I245683,I245827);
nor I_14304 (I245383,I245429,I245810);
DFFARX1 I_14305 (I245810,I2683,I245403,I245392,);
not I_14306 (I245930,I2690);
DFFARX1 I_14307 (I78550,I2683,I245930,I245956,);
nand I_14308 (I245964,I78562,I78571);
and I_14309 (I245981,I245964,I78550);
DFFARX1 I_14310 (I245981,I2683,I245930,I246007,);
nor I_14311 (I245898,I246007,I245956);
not I_14312 (I246029,I246007);
DFFARX1 I_14313 (I78565,I2683,I245930,I246055,);
nand I_14314 (I246063,I246055,I78553);
not I_14315 (I246080,I246063);
DFFARX1 I_14316 (I246080,I2683,I245930,I246106,);
not I_14317 (I245922,I246106);
nor I_14318 (I246128,I245956,I246063);
nor I_14319 (I245904,I246007,I246128);
DFFARX1 I_14320 (I78556,I2683,I245930,I246168,);
DFFARX1 I_14321 (I246168,I2683,I245930,I246185,);
not I_14322 (I246193,I246185);
not I_14323 (I246210,I246168);
nand I_14324 (I245907,I246210,I246029);
nand I_14325 (I246241,I78547,I78547);
and I_14326 (I246258,I246241,I78559);
DFFARX1 I_14327 (I246258,I2683,I245930,I246284,);
nor I_14328 (I246292,I246284,I245956);
DFFARX1 I_14329 (I246292,I2683,I245930,I245895,);
DFFARX1 I_14330 (I246284,I2683,I245930,I245913,);
nor I_14331 (I246337,I78568,I78547);
not I_14332 (I246354,I246337);
nor I_14333 (I245916,I246193,I246354);
nand I_14334 (I245901,I246210,I246354);
nor I_14335 (I245910,I245956,I246337);
DFFARX1 I_14336 (I246337,I2683,I245930,I245919,);
not I_14337 (I246457,I2690);
DFFARX1 I_14338 (I951888,I2683,I246457,I246483,);
nand I_14339 (I246491,I951903,I951888);
and I_14340 (I246508,I246491,I951906);
DFFARX1 I_14341 (I246508,I2683,I246457,I246534,);
nor I_14342 (I246425,I246534,I246483);
not I_14343 (I246556,I246534);
DFFARX1 I_14344 (I951912,I2683,I246457,I246582,);
nand I_14345 (I246590,I246582,I951894);
not I_14346 (I246607,I246590);
DFFARX1 I_14347 (I246607,I2683,I246457,I246633,);
not I_14348 (I246449,I246633);
nor I_14349 (I246655,I246483,I246590);
nor I_14350 (I246431,I246534,I246655);
DFFARX1 I_14351 (I951891,I2683,I246457,I246695,);
DFFARX1 I_14352 (I246695,I2683,I246457,I246712,);
not I_14353 (I246720,I246712);
not I_14354 (I246737,I246695);
nand I_14355 (I246434,I246737,I246556);
nand I_14356 (I246768,I951891,I951897);
and I_14357 (I246785,I246768,I951909);
DFFARX1 I_14358 (I246785,I2683,I246457,I246811,);
nor I_14359 (I246819,I246811,I246483);
DFFARX1 I_14360 (I246819,I2683,I246457,I246422,);
DFFARX1 I_14361 (I246811,I2683,I246457,I246440,);
nor I_14362 (I246864,I951900,I951897);
not I_14363 (I246881,I246864);
nor I_14364 (I246443,I246720,I246881);
nand I_14365 (I246428,I246737,I246881);
nor I_14366 (I246437,I246483,I246864);
DFFARX1 I_14367 (I246864,I2683,I246457,I246446,);
not I_14368 (I246984,I2690);
DFFARX1 I_14369 (I1101305,I2683,I246984,I247010,);
nand I_14370 (I247018,I1101284,I1101284);
and I_14371 (I247035,I247018,I1101311);
DFFARX1 I_14372 (I247035,I2683,I246984,I247061,);
nor I_14373 (I246952,I247061,I247010);
not I_14374 (I247083,I247061);
DFFARX1 I_14375 (I1101299,I2683,I246984,I247109,);
nand I_14376 (I247117,I247109,I1101302);
not I_14377 (I247134,I247117);
DFFARX1 I_14378 (I247134,I2683,I246984,I247160,);
not I_14379 (I246976,I247160);
nor I_14380 (I247182,I247010,I247117);
nor I_14381 (I246958,I247061,I247182);
DFFARX1 I_14382 (I1101293,I2683,I246984,I247222,);
DFFARX1 I_14383 (I247222,I2683,I246984,I247239,);
not I_14384 (I247247,I247239);
not I_14385 (I247264,I247222);
nand I_14386 (I246961,I247264,I247083);
nand I_14387 (I247295,I1101290,I1101287);
and I_14388 (I247312,I247295,I1101308);
DFFARX1 I_14389 (I247312,I2683,I246984,I247338,);
nor I_14390 (I247346,I247338,I247010);
DFFARX1 I_14391 (I247346,I2683,I246984,I246949,);
DFFARX1 I_14392 (I247338,I2683,I246984,I246967,);
nor I_14393 (I247391,I1101296,I1101287);
not I_14394 (I247408,I247391);
nor I_14395 (I246970,I247247,I247408);
nand I_14396 (I246955,I247264,I247408);
nor I_14397 (I246964,I247010,I247391);
DFFARX1 I_14398 (I247391,I2683,I246984,I246973,);
not I_14399 (I247511,I2690);
DFFARX1 I_14400 (I419315,I2683,I247511,I247537,);
nand I_14401 (I247545,I419315,I419327);
and I_14402 (I247562,I247545,I419312);
DFFARX1 I_14403 (I247562,I2683,I247511,I247588,);
nor I_14404 (I247479,I247588,I247537);
not I_14405 (I247610,I247588);
DFFARX1 I_14406 (I419336,I2683,I247511,I247636,);
nand I_14407 (I247644,I247636,I419333);
not I_14408 (I247661,I247644);
DFFARX1 I_14409 (I247661,I2683,I247511,I247687,);
not I_14410 (I247503,I247687);
nor I_14411 (I247709,I247537,I247644);
nor I_14412 (I247485,I247588,I247709);
DFFARX1 I_14413 (I419324,I2683,I247511,I247749,);
DFFARX1 I_14414 (I247749,I2683,I247511,I247766,);
not I_14415 (I247774,I247766);
not I_14416 (I247791,I247749);
nand I_14417 (I247488,I247791,I247610);
nand I_14418 (I247822,I419312,I419321);
and I_14419 (I247839,I247822,I419330);
DFFARX1 I_14420 (I247839,I2683,I247511,I247865,);
nor I_14421 (I247873,I247865,I247537);
DFFARX1 I_14422 (I247873,I2683,I247511,I247476,);
DFFARX1 I_14423 (I247865,I2683,I247511,I247494,);
nor I_14424 (I247918,I419318,I419321);
not I_14425 (I247935,I247918);
nor I_14426 (I247497,I247774,I247935);
nand I_14427 (I247482,I247791,I247935);
nor I_14428 (I247491,I247537,I247918);
DFFARX1 I_14429 (I247918,I2683,I247511,I247500,);
not I_14430 (I248038,I2690);
DFFARX1 I_14431 (I876748,I2683,I248038,I248064,);
nand I_14432 (I248072,I876763,I876748);
and I_14433 (I248089,I248072,I876766);
DFFARX1 I_14434 (I248089,I2683,I248038,I248115,);
nor I_14435 (I248006,I248115,I248064);
not I_14436 (I248137,I248115);
DFFARX1 I_14437 (I876772,I2683,I248038,I248163,);
nand I_14438 (I248171,I248163,I876754);
not I_14439 (I248188,I248171);
DFFARX1 I_14440 (I248188,I2683,I248038,I248214,);
not I_14441 (I248030,I248214);
nor I_14442 (I248236,I248064,I248171);
nor I_14443 (I248012,I248115,I248236);
DFFARX1 I_14444 (I876751,I2683,I248038,I248276,);
DFFARX1 I_14445 (I248276,I2683,I248038,I248293,);
not I_14446 (I248301,I248293);
not I_14447 (I248318,I248276);
nand I_14448 (I248015,I248318,I248137);
nand I_14449 (I248349,I876751,I876757);
and I_14450 (I248366,I248349,I876769);
DFFARX1 I_14451 (I248366,I2683,I248038,I248392,);
nor I_14452 (I248400,I248392,I248064);
DFFARX1 I_14453 (I248400,I2683,I248038,I248003,);
DFFARX1 I_14454 (I248392,I2683,I248038,I248021,);
nor I_14455 (I248445,I876760,I876757);
not I_14456 (I248462,I248445);
nor I_14457 (I248024,I248301,I248462);
nand I_14458 (I248009,I248318,I248462);
nor I_14459 (I248018,I248064,I248445);
DFFARX1 I_14460 (I248445,I2683,I248038,I248027,);
not I_14461 (I248565,I2690);
DFFARX1 I_14462 (I949576,I2683,I248565,I248591,);
nand I_14463 (I248599,I949591,I949576);
and I_14464 (I248616,I248599,I949594);
DFFARX1 I_14465 (I248616,I2683,I248565,I248642,);
nor I_14466 (I248533,I248642,I248591);
not I_14467 (I248664,I248642);
DFFARX1 I_14468 (I949600,I2683,I248565,I248690,);
nand I_14469 (I248698,I248690,I949582);
not I_14470 (I248715,I248698);
DFFARX1 I_14471 (I248715,I2683,I248565,I248741,);
not I_14472 (I248557,I248741);
nor I_14473 (I248763,I248591,I248698);
nor I_14474 (I248539,I248642,I248763);
DFFARX1 I_14475 (I949579,I2683,I248565,I248803,);
DFFARX1 I_14476 (I248803,I2683,I248565,I248820,);
not I_14477 (I248828,I248820);
not I_14478 (I248845,I248803);
nand I_14479 (I248542,I248845,I248664);
nand I_14480 (I248876,I949579,I949585);
and I_14481 (I248893,I248876,I949597);
DFFARX1 I_14482 (I248893,I2683,I248565,I248919,);
nor I_14483 (I248927,I248919,I248591);
DFFARX1 I_14484 (I248927,I2683,I248565,I248530,);
DFFARX1 I_14485 (I248919,I2683,I248565,I248548,);
nor I_14486 (I248972,I949588,I949585);
not I_14487 (I248989,I248972);
nor I_14488 (I248551,I248828,I248989);
nand I_14489 (I248536,I248845,I248989);
nor I_14490 (I248545,I248591,I248972);
DFFARX1 I_14491 (I248972,I2683,I248565,I248554,);
not I_14492 (I249092,I2690);
DFFARX1 I_14493 (I605814,I2683,I249092,I249118,);
nand I_14494 (I249126,I605805,I605820);
and I_14495 (I249143,I249126,I605826);
DFFARX1 I_14496 (I249143,I2683,I249092,I249169,);
nor I_14497 (I249060,I249169,I249118);
not I_14498 (I249191,I249169);
DFFARX1 I_14499 (I605811,I2683,I249092,I249217,);
nand I_14500 (I249225,I249217,I605805);
not I_14501 (I249242,I249225);
DFFARX1 I_14502 (I249242,I2683,I249092,I249268,);
not I_14503 (I249084,I249268);
nor I_14504 (I249290,I249118,I249225);
nor I_14505 (I249066,I249169,I249290);
DFFARX1 I_14506 (I605808,I2683,I249092,I249330,);
DFFARX1 I_14507 (I249330,I2683,I249092,I249347,);
not I_14508 (I249355,I249347);
not I_14509 (I249372,I249330);
nand I_14510 (I249069,I249372,I249191);
nand I_14511 (I249403,I605802,I605817);
and I_14512 (I249420,I249403,I605802);
DFFARX1 I_14513 (I249420,I2683,I249092,I249446,);
nor I_14514 (I249454,I249446,I249118);
DFFARX1 I_14515 (I249454,I2683,I249092,I249057,);
DFFARX1 I_14516 (I249446,I2683,I249092,I249075,);
nor I_14517 (I249499,I605823,I605817);
not I_14518 (I249516,I249499);
nor I_14519 (I249078,I249355,I249516);
nand I_14520 (I249063,I249372,I249516);
nor I_14521 (I249072,I249118,I249499);
DFFARX1 I_14522 (I249499,I2683,I249092,I249081,);
not I_14523 (I249619,I2690);
DFFARX1 I_14524 (I722578,I2683,I249619,I249645,);
nand I_14525 (I249653,I722575,I722593);
and I_14526 (I249670,I249653,I722584);
DFFARX1 I_14527 (I249670,I2683,I249619,I249696,);
nor I_14528 (I249587,I249696,I249645);
not I_14529 (I249718,I249696);
DFFARX1 I_14530 (I722599,I2683,I249619,I249744,);
nand I_14531 (I249752,I249744,I722581);
not I_14532 (I249769,I249752);
DFFARX1 I_14533 (I249769,I2683,I249619,I249795,);
not I_14534 (I249611,I249795);
nor I_14535 (I249817,I249645,I249752);
nor I_14536 (I249593,I249696,I249817);
DFFARX1 I_14537 (I722587,I2683,I249619,I249857,);
DFFARX1 I_14538 (I249857,I2683,I249619,I249874,);
not I_14539 (I249882,I249874);
not I_14540 (I249899,I249857);
nand I_14541 (I249596,I249899,I249718);
nand I_14542 (I249930,I722575,I722602);
and I_14543 (I249947,I249930,I722590);
DFFARX1 I_14544 (I249947,I2683,I249619,I249973,);
nor I_14545 (I249981,I249973,I249645);
DFFARX1 I_14546 (I249981,I2683,I249619,I249584,);
DFFARX1 I_14547 (I249973,I2683,I249619,I249602,);
nor I_14548 (I250026,I722596,I722602);
not I_14549 (I250043,I250026);
nor I_14550 (I249605,I249882,I250043);
nand I_14551 (I249590,I249899,I250043);
nor I_14552 (I249599,I249645,I250026);
DFFARX1 I_14553 (I250026,I2683,I249619,I249608,);
not I_14554 (I250146,I2690);
DFFARX1 I_14555 (I924722,I2683,I250146,I250172,);
nand I_14556 (I250180,I924737,I924722);
and I_14557 (I250197,I250180,I924740);
DFFARX1 I_14558 (I250197,I2683,I250146,I250223,);
nor I_14559 (I250114,I250223,I250172);
not I_14560 (I250245,I250223);
DFFARX1 I_14561 (I924746,I2683,I250146,I250271,);
nand I_14562 (I250279,I250271,I924728);
not I_14563 (I250296,I250279);
DFFARX1 I_14564 (I250296,I2683,I250146,I250322,);
not I_14565 (I250138,I250322);
nor I_14566 (I250344,I250172,I250279);
nor I_14567 (I250120,I250223,I250344);
DFFARX1 I_14568 (I924725,I2683,I250146,I250384,);
DFFARX1 I_14569 (I250384,I2683,I250146,I250401,);
not I_14570 (I250409,I250401);
not I_14571 (I250426,I250384);
nand I_14572 (I250123,I250426,I250245);
nand I_14573 (I250457,I924725,I924731);
and I_14574 (I250474,I250457,I924743);
DFFARX1 I_14575 (I250474,I2683,I250146,I250500,);
nor I_14576 (I250508,I250500,I250172);
DFFARX1 I_14577 (I250508,I2683,I250146,I250111,);
DFFARX1 I_14578 (I250500,I2683,I250146,I250129,);
nor I_14579 (I250553,I924734,I924731);
not I_14580 (I250570,I250553);
nor I_14581 (I250132,I250409,I250570);
nand I_14582 (I250117,I250426,I250570);
nor I_14583 (I250126,I250172,I250553);
DFFARX1 I_14584 (I250553,I2683,I250146,I250135,);
not I_14585 (I250673,I2690);
DFFARX1 I_14586 (I792346,I2683,I250673,I250699,);
nand I_14587 (I250707,I792343,I792361);
and I_14588 (I250724,I250707,I792352);
DFFARX1 I_14589 (I250724,I2683,I250673,I250750,);
nor I_14590 (I250641,I250750,I250699);
not I_14591 (I250772,I250750);
DFFARX1 I_14592 (I792367,I2683,I250673,I250798,);
nand I_14593 (I250806,I250798,I792349);
not I_14594 (I250823,I250806);
DFFARX1 I_14595 (I250823,I2683,I250673,I250849,);
not I_14596 (I250665,I250849);
nor I_14597 (I250871,I250699,I250806);
nor I_14598 (I250647,I250750,I250871);
DFFARX1 I_14599 (I792355,I2683,I250673,I250911,);
DFFARX1 I_14600 (I250911,I2683,I250673,I250928,);
not I_14601 (I250936,I250928);
not I_14602 (I250953,I250911);
nand I_14603 (I250650,I250953,I250772);
nand I_14604 (I250984,I792343,I792370);
and I_14605 (I251001,I250984,I792358);
DFFARX1 I_14606 (I251001,I2683,I250673,I251027,);
nor I_14607 (I251035,I251027,I250699);
DFFARX1 I_14608 (I251035,I2683,I250673,I250638,);
DFFARX1 I_14609 (I251027,I2683,I250673,I250656,);
nor I_14610 (I251080,I792364,I792370);
not I_14611 (I251097,I251080);
nor I_14612 (I250659,I250936,I251097);
nand I_14613 (I250644,I250953,I251097);
nor I_14614 (I250653,I250699,I251080);
DFFARX1 I_14615 (I251080,I2683,I250673,I250662,);
not I_14616 (I251200,I2690);
DFFARX1 I_14617 (I610438,I2683,I251200,I251226,);
nand I_14618 (I251234,I610429,I610444);
and I_14619 (I251251,I251234,I610450);
DFFARX1 I_14620 (I251251,I2683,I251200,I251277,);
nor I_14621 (I251168,I251277,I251226);
not I_14622 (I251299,I251277);
DFFARX1 I_14623 (I610435,I2683,I251200,I251325,);
nand I_14624 (I251333,I251325,I610429);
not I_14625 (I251350,I251333);
DFFARX1 I_14626 (I251350,I2683,I251200,I251376,);
not I_14627 (I251192,I251376);
nor I_14628 (I251398,I251226,I251333);
nor I_14629 (I251174,I251277,I251398);
DFFARX1 I_14630 (I610432,I2683,I251200,I251438,);
DFFARX1 I_14631 (I251438,I2683,I251200,I251455,);
not I_14632 (I251463,I251455);
not I_14633 (I251480,I251438);
nand I_14634 (I251177,I251480,I251299);
nand I_14635 (I251511,I610426,I610441);
and I_14636 (I251528,I251511,I610426);
DFFARX1 I_14637 (I251528,I2683,I251200,I251554,);
nor I_14638 (I251562,I251554,I251226);
DFFARX1 I_14639 (I251562,I2683,I251200,I251165,);
DFFARX1 I_14640 (I251554,I2683,I251200,I251183,);
nor I_14641 (I251607,I610447,I610441);
not I_14642 (I251624,I251607);
nor I_14643 (I251186,I251463,I251624);
nand I_14644 (I251171,I251480,I251624);
nor I_14645 (I251180,I251226,I251607);
DFFARX1 I_14646 (I251607,I2683,I251200,I251189,);
not I_14647 (I251727,I2690);
DFFARX1 I_14648 (I68537,I2683,I251727,I251753,);
nand I_14649 (I251761,I68549,I68558);
and I_14650 (I251778,I251761,I68537);
DFFARX1 I_14651 (I251778,I2683,I251727,I251804,);
nor I_14652 (I251695,I251804,I251753);
not I_14653 (I251826,I251804);
DFFARX1 I_14654 (I68552,I2683,I251727,I251852,);
nand I_14655 (I251860,I251852,I68540);
not I_14656 (I251877,I251860);
DFFARX1 I_14657 (I251877,I2683,I251727,I251903,);
not I_14658 (I251719,I251903);
nor I_14659 (I251925,I251753,I251860);
nor I_14660 (I251701,I251804,I251925);
DFFARX1 I_14661 (I68543,I2683,I251727,I251965,);
DFFARX1 I_14662 (I251965,I2683,I251727,I251982,);
not I_14663 (I251990,I251982);
not I_14664 (I252007,I251965);
nand I_14665 (I251704,I252007,I251826);
nand I_14666 (I252038,I68534,I68534);
and I_14667 (I252055,I252038,I68546);
DFFARX1 I_14668 (I252055,I2683,I251727,I252081,);
nor I_14669 (I252089,I252081,I251753);
DFFARX1 I_14670 (I252089,I2683,I251727,I251692,);
DFFARX1 I_14671 (I252081,I2683,I251727,I251710,);
nor I_14672 (I252134,I68555,I68534);
not I_14673 (I252151,I252134);
nor I_14674 (I251713,I251990,I252151);
nand I_14675 (I251698,I252007,I252151);
nor I_14676 (I251707,I251753,I252134);
DFFARX1 I_14677 (I252134,I2683,I251727,I251716,);
not I_14678 (I252254,I2690);
DFFARX1 I_14679 (I568244,I2683,I252254,I252280,);
nand I_14680 (I252288,I568235,I568250);
and I_14681 (I252305,I252288,I568256);
DFFARX1 I_14682 (I252305,I2683,I252254,I252331,);
nor I_14683 (I252222,I252331,I252280);
not I_14684 (I252353,I252331);
DFFARX1 I_14685 (I568241,I2683,I252254,I252379,);
nand I_14686 (I252387,I252379,I568235);
not I_14687 (I252404,I252387);
DFFARX1 I_14688 (I252404,I2683,I252254,I252430,);
not I_14689 (I252246,I252430);
nor I_14690 (I252452,I252280,I252387);
nor I_14691 (I252228,I252331,I252452);
DFFARX1 I_14692 (I568238,I2683,I252254,I252492,);
DFFARX1 I_14693 (I252492,I2683,I252254,I252509,);
not I_14694 (I252517,I252509);
not I_14695 (I252534,I252492);
nand I_14696 (I252231,I252534,I252353);
nand I_14697 (I252565,I568232,I568247);
and I_14698 (I252582,I252565,I568232);
DFFARX1 I_14699 (I252582,I2683,I252254,I252608,);
nor I_14700 (I252616,I252608,I252280);
DFFARX1 I_14701 (I252616,I2683,I252254,I252219,);
DFFARX1 I_14702 (I252608,I2683,I252254,I252237,);
nor I_14703 (I252661,I568253,I568247);
not I_14704 (I252678,I252661);
nor I_14705 (I252240,I252517,I252678);
nand I_14706 (I252225,I252534,I252678);
nor I_14707 (I252234,I252280,I252661);
DFFARX1 I_14708 (I252661,I2683,I252254,I252243,);
not I_14709 (I252781,I2690);
DFFARX1 I_14710 (I487905,I2683,I252781,I252807,);
nand I_14711 (I252815,I487890,I487893);
and I_14712 (I252832,I252815,I487908);
DFFARX1 I_14713 (I252832,I2683,I252781,I252858,);
nor I_14714 (I252749,I252858,I252807);
not I_14715 (I252880,I252858);
DFFARX1 I_14716 (I487902,I2683,I252781,I252906,);
nand I_14717 (I252914,I252906,I487893);
not I_14718 (I252931,I252914);
DFFARX1 I_14719 (I252931,I2683,I252781,I252957,);
not I_14720 (I252773,I252957);
nor I_14721 (I252979,I252807,I252914);
nor I_14722 (I252755,I252858,I252979);
DFFARX1 I_14723 (I487899,I2683,I252781,I253019,);
DFFARX1 I_14724 (I253019,I2683,I252781,I253036,);
not I_14725 (I253044,I253036);
not I_14726 (I253061,I253019);
nand I_14727 (I252758,I253061,I252880);
nand I_14728 (I253092,I487914,I487890);
and I_14729 (I253109,I253092,I487911);
DFFARX1 I_14730 (I253109,I2683,I252781,I253135,);
nor I_14731 (I253143,I253135,I252807);
DFFARX1 I_14732 (I253143,I2683,I252781,I252746,);
DFFARX1 I_14733 (I253135,I2683,I252781,I252764,);
nor I_14734 (I253188,I487896,I487890);
not I_14735 (I253205,I253188);
nor I_14736 (I252767,I253044,I253205);
nand I_14737 (I252752,I253061,I253205);
nor I_14738 (I252761,I252807,I253188);
DFFARX1 I_14739 (I253188,I2683,I252781,I252770,);
not I_14740 (I253308,I2690);
DFFARX1 I_14741 (I507554,I2683,I253308,I253334,);
nand I_14742 (I253342,I507545,I507560);
and I_14743 (I253359,I253342,I507566);
DFFARX1 I_14744 (I253359,I2683,I253308,I253385,);
nor I_14745 (I253276,I253385,I253334);
not I_14746 (I253407,I253385);
DFFARX1 I_14747 (I507551,I2683,I253308,I253433,);
nand I_14748 (I253441,I253433,I507545);
not I_14749 (I253458,I253441);
DFFARX1 I_14750 (I253458,I2683,I253308,I253484,);
not I_14751 (I253300,I253484);
nor I_14752 (I253506,I253334,I253441);
nor I_14753 (I253282,I253385,I253506);
DFFARX1 I_14754 (I507548,I2683,I253308,I253546,);
DFFARX1 I_14755 (I253546,I2683,I253308,I253563,);
not I_14756 (I253571,I253563);
not I_14757 (I253588,I253546);
nand I_14758 (I253285,I253588,I253407);
nand I_14759 (I253619,I507542,I507557);
and I_14760 (I253636,I253619,I507542);
DFFARX1 I_14761 (I253636,I2683,I253308,I253662,);
nor I_14762 (I253670,I253662,I253334);
DFFARX1 I_14763 (I253670,I2683,I253308,I253273,);
DFFARX1 I_14764 (I253662,I2683,I253308,I253291,);
nor I_14765 (I253715,I507563,I507557);
not I_14766 (I253732,I253715);
nor I_14767 (I253294,I253571,I253732);
nand I_14768 (I253279,I253588,I253732);
nor I_14769 (I253288,I253334,I253715);
DFFARX1 I_14770 (I253715,I2683,I253308,I253297,);
not I_14771 (I253835,I2690);
DFFARX1 I_14772 (I721286,I2683,I253835,I253861,);
nand I_14773 (I253869,I721283,I721301);
and I_14774 (I253886,I253869,I721292);
DFFARX1 I_14775 (I253886,I2683,I253835,I253912,);
nor I_14776 (I253803,I253912,I253861);
not I_14777 (I253934,I253912);
DFFARX1 I_14778 (I721307,I2683,I253835,I253960,);
nand I_14779 (I253968,I253960,I721289);
not I_14780 (I253985,I253968);
DFFARX1 I_14781 (I253985,I2683,I253835,I254011,);
not I_14782 (I253827,I254011);
nor I_14783 (I254033,I253861,I253968);
nor I_14784 (I253809,I253912,I254033);
DFFARX1 I_14785 (I721295,I2683,I253835,I254073,);
DFFARX1 I_14786 (I254073,I2683,I253835,I254090,);
not I_14787 (I254098,I254090);
not I_14788 (I254115,I254073);
nand I_14789 (I253812,I254115,I253934);
nand I_14790 (I254146,I721283,I721310);
and I_14791 (I254163,I254146,I721298);
DFFARX1 I_14792 (I254163,I2683,I253835,I254189,);
nor I_14793 (I254197,I254189,I253861);
DFFARX1 I_14794 (I254197,I2683,I253835,I253800,);
DFFARX1 I_14795 (I254189,I2683,I253835,I253818,);
nor I_14796 (I254242,I721304,I721310);
not I_14797 (I254259,I254242);
nor I_14798 (I253821,I254098,I254259);
nand I_14799 (I253806,I254115,I254259);
nor I_14800 (I253815,I253861,I254242);
DFFARX1 I_14801 (I254242,I2683,I253835,I253824,);
not I_14802 (I254362,I2690);
DFFARX1 I_14803 (I658624,I2683,I254362,I254388,);
nand I_14804 (I254396,I658627,I658621);
and I_14805 (I254413,I254396,I658633);
DFFARX1 I_14806 (I254413,I2683,I254362,I254439,);
nor I_14807 (I254330,I254439,I254388);
not I_14808 (I254461,I254439);
DFFARX1 I_14809 (I658636,I2683,I254362,I254487,);
nand I_14810 (I254495,I254487,I658627);
not I_14811 (I254512,I254495);
DFFARX1 I_14812 (I254512,I2683,I254362,I254538,);
not I_14813 (I254354,I254538);
nor I_14814 (I254560,I254388,I254495);
nor I_14815 (I254336,I254439,I254560);
DFFARX1 I_14816 (I658639,I2683,I254362,I254600,);
DFFARX1 I_14817 (I254600,I2683,I254362,I254617,);
not I_14818 (I254625,I254617);
not I_14819 (I254642,I254600);
nand I_14820 (I254339,I254642,I254461);
nand I_14821 (I254673,I658621,I658630);
and I_14822 (I254690,I254673,I658624);
DFFARX1 I_14823 (I254690,I2683,I254362,I254716,);
nor I_14824 (I254724,I254716,I254388);
DFFARX1 I_14825 (I254724,I2683,I254362,I254327,);
DFFARX1 I_14826 (I254716,I2683,I254362,I254345,);
nor I_14827 (I254769,I658642,I658630);
not I_14828 (I254786,I254769);
nor I_14829 (I254348,I254625,I254786);
nand I_14830 (I254333,I254642,I254786);
nor I_14831 (I254342,I254388,I254769);
DFFARX1 I_14832 (I254769,I2683,I254362,I254351,);
not I_14833 (I254889,I2690);
DFFARX1 I_14834 (I531252,I2683,I254889,I254915,);
nand I_14835 (I254923,I531243,I531258);
and I_14836 (I254940,I254923,I531264);
DFFARX1 I_14837 (I254940,I2683,I254889,I254966,);
nor I_14838 (I254857,I254966,I254915);
not I_14839 (I254988,I254966);
DFFARX1 I_14840 (I531249,I2683,I254889,I255014,);
nand I_14841 (I255022,I255014,I531243);
not I_14842 (I255039,I255022);
DFFARX1 I_14843 (I255039,I2683,I254889,I255065,);
not I_14844 (I254881,I255065);
nor I_14845 (I255087,I254915,I255022);
nor I_14846 (I254863,I254966,I255087);
DFFARX1 I_14847 (I531246,I2683,I254889,I255127,);
DFFARX1 I_14848 (I255127,I2683,I254889,I255144,);
not I_14849 (I255152,I255144);
not I_14850 (I255169,I255127);
nand I_14851 (I254866,I255169,I254988);
nand I_14852 (I255200,I531240,I531255);
and I_14853 (I255217,I255200,I531240);
DFFARX1 I_14854 (I255217,I2683,I254889,I255243,);
nor I_14855 (I255251,I255243,I254915);
DFFARX1 I_14856 (I255251,I2683,I254889,I254854,);
DFFARX1 I_14857 (I255243,I2683,I254889,I254872,);
nor I_14858 (I255296,I531261,I531255);
not I_14859 (I255313,I255296);
nor I_14860 (I254875,I255152,I255313);
nand I_14861 (I254860,I255169,I255313);
nor I_14862 (I254869,I254915,I255296);
DFFARX1 I_14863 (I255296,I2683,I254889,I254878,);
not I_14864 (I255416,I2690);
DFFARX1 I_14865 (I971728,I2683,I255416,I255442,);
nand I_14866 (I255450,I971710,I971734);
and I_14867 (I255467,I255450,I971725);
DFFARX1 I_14868 (I255467,I2683,I255416,I255493,);
nor I_14869 (I255384,I255493,I255442);
not I_14870 (I255515,I255493);
DFFARX1 I_14871 (I971731,I2683,I255416,I255541,);
nand I_14872 (I255549,I255541,I971719);
not I_14873 (I255566,I255549);
DFFARX1 I_14874 (I255566,I2683,I255416,I255592,);
not I_14875 (I255408,I255592);
nor I_14876 (I255614,I255442,I255549);
nor I_14877 (I255390,I255493,I255614);
DFFARX1 I_14878 (I971710,I2683,I255416,I255654,);
DFFARX1 I_14879 (I255654,I2683,I255416,I255671,);
not I_14880 (I255679,I255671);
not I_14881 (I255696,I255654);
nand I_14882 (I255393,I255696,I255515);
nand I_14883 (I255727,I971716,I971713);
and I_14884 (I255744,I255727,I971722);
DFFARX1 I_14885 (I255744,I2683,I255416,I255770,);
nor I_14886 (I255778,I255770,I255442);
DFFARX1 I_14887 (I255778,I2683,I255416,I255381,);
DFFARX1 I_14888 (I255770,I2683,I255416,I255399,);
nor I_14889 (I255823,I971713,I971713);
not I_14890 (I255840,I255823);
nor I_14891 (I255402,I255679,I255840);
nand I_14892 (I255387,I255696,I255840);
nor I_14893 (I255396,I255442,I255823);
DFFARX1 I_14894 (I255823,I2683,I255416,I255405,);
not I_14895 (I255943,I2690);
DFFARX1 I_14896 (I641760,I2683,I255943,I255969,);
nand I_14897 (I255977,I641763,I641757);
and I_14898 (I255994,I255977,I641769);
DFFARX1 I_14899 (I255994,I2683,I255943,I256020,);
nor I_14900 (I255911,I256020,I255969);
not I_14901 (I256042,I256020);
DFFARX1 I_14902 (I641772,I2683,I255943,I256068,);
nand I_14903 (I256076,I256068,I641763);
not I_14904 (I256093,I256076);
DFFARX1 I_14905 (I256093,I2683,I255943,I256119,);
not I_14906 (I255935,I256119);
nor I_14907 (I256141,I255969,I256076);
nor I_14908 (I255917,I256020,I256141);
DFFARX1 I_14909 (I641775,I2683,I255943,I256181,);
DFFARX1 I_14910 (I256181,I2683,I255943,I256198,);
not I_14911 (I256206,I256198);
not I_14912 (I256223,I256181);
nand I_14913 (I255920,I256223,I256042);
nand I_14914 (I256254,I641757,I641766);
and I_14915 (I256271,I256254,I641760);
DFFARX1 I_14916 (I256271,I2683,I255943,I256297,);
nor I_14917 (I256305,I256297,I255969);
DFFARX1 I_14918 (I256305,I2683,I255943,I255908,);
DFFARX1 I_14919 (I256297,I2683,I255943,I255926,);
nor I_14920 (I256350,I641778,I641766);
not I_14921 (I256367,I256350);
nor I_14922 (I255929,I256206,I256367);
nand I_14923 (I255914,I256223,I256367);
nor I_14924 (I255923,I255969,I256350);
DFFARX1 I_14925 (I256350,I2683,I255943,I255932,);
not I_14926 (I256470,I2690);
DFFARX1 I_14927 (I579226,I2683,I256470,I256496,);
nand I_14928 (I256504,I579217,I579232);
and I_14929 (I256521,I256504,I579238);
DFFARX1 I_14930 (I256521,I2683,I256470,I256547,);
nor I_14931 (I256438,I256547,I256496);
not I_14932 (I256569,I256547);
DFFARX1 I_14933 (I579223,I2683,I256470,I256595,);
nand I_14934 (I256603,I256595,I579217);
not I_14935 (I256620,I256603);
DFFARX1 I_14936 (I256620,I2683,I256470,I256646,);
not I_14937 (I256462,I256646);
nor I_14938 (I256668,I256496,I256603);
nor I_14939 (I256444,I256547,I256668);
DFFARX1 I_14940 (I579220,I2683,I256470,I256708,);
DFFARX1 I_14941 (I256708,I2683,I256470,I256725,);
not I_14942 (I256733,I256725);
not I_14943 (I256750,I256708);
nand I_14944 (I256447,I256750,I256569);
nand I_14945 (I256781,I579214,I579229);
and I_14946 (I256798,I256781,I579214);
DFFARX1 I_14947 (I256798,I2683,I256470,I256824,);
nor I_14948 (I256832,I256824,I256496);
DFFARX1 I_14949 (I256832,I2683,I256470,I256435,);
DFFARX1 I_14950 (I256824,I2683,I256470,I256453,);
nor I_14951 (I256877,I579235,I579229);
not I_14952 (I256894,I256877);
nor I_14953 (I256456,I256733,I256894);
nand I_14954 (I256441,I256750,I256894);
nor I_14955 (I256450,I256496,I256877);
DFFARX1 I_14956 (I256877,I2683,I256470,I256459,);
not I_14957 (I256997,I2690);
DFFARX1 I_14958 (I155710,I2683,I256997,I257023,);
nand I_14959 (I257031,I155710,I155716);
and I_14960 (I257048,I257031,I155734);
DFFARX1 I_14961 (I257048,I2683,I256997,I257074,);
nor I_14962 (I256965,I257074,I257023);
not I_14963 (I257096,I257074);
DFFARX1 I_14964 (I155722,I2683,I256997,I257122,);
nand I_14965 (I257130,I257122,I155719);
not I_14966 (I257147,I257130);
DFFARX1 I_14967 (I257147,I2683,I256997,I257173,);
not I_14968 (I256989,I257173);
nor I_14969 (I257195,I257023,I257130);
nor I_14970 (I256971,I257074,I257195);
DFFARX1 I_14971 (I155728,I2683,I256997,I257235,);
DFFARX1 I_14972 (I257235,I2683,I256997,I257252,);
not I_14973 (I257260,I257252);
not I_14974 (I257277,I257235);
nand I_14975 (I256974,I257277,I257096);
nand I_14976 (I257308,I155713,I155713);
and I_14977 (I257325,I257308,I155725);
DFFARX1 I_14978 (I257325,I2683,I256997,I257351,);
nor I_14979 (I257359,I257351,I257023);
DFFARX1 I_14980 (I257359,I2683,I256997,I256962,);
DFFARX1 I_14981 (I257351,I2683,I256997,I256980,);
nor I_14982 (I257404,I155731,I155713);
not I_14983 (I257421,I257404);
nor I_14984 (I256983,I257260,I257421);
nand I_14985 (I256968,I257277,I257421);
nor I_14986 (I256977,I257023,I257404);
DFFARX1 I_14987 (I257404,I2683,I256997,I256986,);
not I_14988 (I257524,I2690);
DFFARX1 I_14989 (I882528,I2683,I257524,I257550,);
nand I_14990 (I257558,I882543,I882528);
and I_14991 (I257575,I257558,I882546);
DFFARX1 I_14992 (I257575,I2683,I257524,I257601,);
nor I_14993 (I257492,I257601,I257550);
not I_14994 (I257623,I257601);
DFFARX1 I_14995 (I882552,I2683,I257524,I257649,);
nand I_14996 (I257657,I257649,I882534);
not I_14997 (I257674,I257657);
DFFARX1 I_14998 (I257674,I2683,I257524,I257700,);
not I_14999 (I257516,I257700);
nor I_15000 (I257722,I257550,I257657);
nor I_15001 (I257498,I257601,I257722);
DFFARX1 I_15002 (I882531,I2683,I257524,I257762,);
DFFARX1 I_15003 (I257762,I2683,I257524,I257779,);
not I_15004 (I257787,I257779);
not I_15005 (I257804,I257762);
nand I_15006 (I257501,I257804,I257623);
nand I_15007 (I257835,I882531,I882537);
and I_15008 (I257852,I257835,I882549);
DFFARX1 I_15009 (I257852,I2683,I257524,I257878,);
nor I_15010 (I257886,I257878,I257550);
DFFARX1 I_15011 (I257886,I2683,I257524,I257489,);
DFFARX1 I_15012 (I257878,I2683,I257524,I257507,);
nor I_15013 (I257931,I882540,I882537);
not I_15014 (I257948,I257931);
nor I_15015 (I257510,I257787,I257948);
nand I_15016 (I257495,I257804,I257948);
nor I_15017 (I257504,I257550,I257931);
DFFARX1 I_15018 (I257931,I2683,I257524,I257513,);
not I_15019 (I258051,I2690);
DFFARX1 I_15020 (I571712,I2683,I258051,I258077,);
nand I_15021 (I258085,I571703,I571718);
and I_15022 (I258102,I258085,I571724);
DFFARX1 I_15023 (I258102,I2683,I258051,I258128,);
nor I_15024 (I258019,I258128,I258077);
not I_15025 (I258150,I258128);
DFFARX1 I_15026 (I571709,I2683,I258051,I258176,);
nand I_15027 (I258184,I258176,I571703);
not I_15028 (I258201,I258184);
DFFARX1 I_15029 (I258201,I2683,I258051,I258227,);
not I_15030 (I258043,I258227);
nor I_15031 (I258249,I258077,I258184);
nor I_15032 (I258025,I258128,I258249);
DFFARX1 I_15033 (I571706,I2683,I258051,I258289,);
DFFARX1 I_15034 (I258289,I2683,I258051,I258306,);
not I_15035 (I258314,I258306);
not I_15036 (I258331,I258289);
nand I_15037 (I258028,I258331,I258150);
nand I_15038 (I258362,I571700,I571715);
and I_15039 (I258379,I258362,I571700);
DFFARX1 I_15040 (I258379,I2683,I258051,I258405,);
nor I_15041 (I258413,I258405,I258077);
DFFARX1 I_15042 (I258413,I2683,I258051,I258016,);
DFFARX1 I_15043 (I258405,I2683,I258051,I258034,);
nor I_15044 (I258458,I571721,I571715);
not I_15045 (I258475,I258458);
nor I_15046 (I258037,I258314,I258475);
nand I_15047 (I258022,I258331,I258475);
nor I_15048 (I258031,I258077,I258458);
DFFARX1 I_15049 (I258458,I2683,I258051,I258040,);
not I_15050 (I258578,I2690);
DFFARX1 I_15051 (I603502,I2683,I258578,I258604,);
nand I_15052 (I258612,I603493,I603508);
and I_15053 (I258629,I258612,I603514);
DFFARX1 I_15054 (I258629,I2683,I258578,I258655,);
nor I_15055 (I258546,I258655,I258604);
not I_15056 (I258677,I258655);
DFFARX1 I_15057 (I603499,I2683,I258578,I258703,);
nand I_15058 (I258711,I258703,I603493);
not I_15059 (I258728,I258711);
DFFARX1 I_15060 (I258728,I2683,I258578,I258754,);
not I_15061 (I258570,I258754);
nor I_15062 (I258776,I258604,I258711);
nor I_15063 (I258552,I258655,I258776);
DFFARX1 I_15064 (I603496,I2683,I258578,I258816,);
DFFARX1 I_15065 (I258816,I2683,I258578,I258833,);
not I_15066 (I258841,I258833);
not I_15067 (I258858,I258816);
nand I_15068 (I258555,I258858,I258677);
nand I_15069 (I258889,I603490,I603505);
and I_15070 (I258906,I258889,I603490);
DFFARX1 I_15071 (I258906,I2683,I258578,I258932,);
nor I_15072 (I258940,I258932,I258604);
DFFARX1 I_15073 (I258940,I2683,I258578,I258543,);
DFFARX1 I_15074 (I258932,I2683,I258578,I258561,);
nor I_15075 (I258985,I603511,I603505);
not I_15076 (I259002,I258985);
nor I_15077 (I258564,I258841,I259002);
nand I_15078 (I258549,I258858,I259002);
nor I_15079 (I258558,I258604,I258985);
DFFARX1 I_15080 (I258985,I2683,I258578,I258567,);
not I_15081 (I259105,I2690);
DFFARX1 I_15082 (I818662,I2683,I259105,I259131,);
nand I_15083 (I259139,I818659,I818662);
and I_15084 (I259156,I259139,I818671);
DFFARX1 I_15085 (I259156,I2683,I259105,I259182,);
nor I_15086 (I259073,I259182,I259131);
not I_15087 (I259204,I259182);
DFFARX1 I_15088 (I818659,I2683,I259105,I259230,);
nand I_15089 (I259238,I259230,I818677);
not I_15090 (I259255,I259238);
DFFARX1 I_15091 (I259255,I2683,I259105,I259281,);
not I_15092 (I259097,I259281);
nor I_15093 (I259303,I259131,I259238);
nor I_15094 (I259079,I259182,I259303);
DFFARX1 I_15095 (I818665,I2683,I259105,I259343,);
DFFARX1 I_15096 (I259343,I2683,I259105,I259360,);
not I_15097 (I259368,I259360);
not I_15098 (I259385,I259343);
nand I_15099 (I259082,I259385,I259204);
nand I_15100 (I259416,I818674,I818680);
and I_15101 (I259433,I259416,I818665);
DFFARX1 I_15102 (I259433,I2683,I259105,I259459,);
nor I_15103 (I259467,I259459,I259131);
DFFARX1 I_15104 (I259467,I2683,I259105,I259070,);
DFFARX1 I_15105 (I259459,I2683,I259105,I259088,);
nor I_15106 (I259512,I818668,I818680);
not I_15107 (I259529,I259512);
nor I_15108 (I259091,I259368,I259529);
nand I_15109 (I259076,I259385,I259529);
nor I_15110 (I259085,I259131,I259512);
DFFARX1 I_15111 (I259512,I2683,I259105,I259094,);
not I_15112 (I259632,I2690);
DFFARX1 I_15113 (I392158,I2683,I259632,I259658,);
nand I_15114 (I259666,I392170,I392149);
and I_15115 (I259683,I259666,I392173);
DFFARX1 I_15116 (I259683,I2683,I259632,I259709,);
nor I_15117 (I259600,I259709,I259658);
not I_15118 (I259731,I259709);
DFFARX1 I_15119 (I392164,I2683,I259632,I259757,);
nand I_15120 (I259765,I259757,I392146);
not I_15121 (I259782,I259765);
DFFARX1 I_15122 (I259782,I2683,I259632,I259808,);
not I_15123 (I259624,I259808);
nor I_15124 (I259830,I259658,I259765);
nor I_15125 (I259606,I259709,I259830);
DFFARX1 I_15126 (I392161,I2683,I259632,I259870,);
DFFARX1 I_15127 (I259870,I2683,I259632,I259887,);
not I_15128 (I259895,I259887);
not I_15129 (I259912,I259870);
nand I_15130 (I259609,I259912,I259731);
nand I_15131 (I259943,I392146,I392152);
and I_15132 (I259960,I259943,I392155);
DFFARX1 I_15133 (I259960,I2683,I259632,I259986,);
nor I_15134 (I259994,I259986,I259658);
DFFARX1 I_15135 (I259994,I2683,I259632,I259597,);
DFFARX1 I_15136 (I259986,I2683,I259632,I259615,);
nor I_15137 (I260039,I392167,I392152);
not I_15138 (I260056,I260039);
nor I_15139 (I259618,I259895,I260056);
nand I_15140 (I259603,I259912,I260056);
nor I_15141 (I259612,I259658,I260039);
DFFARX1 I_15142 (I260039,I2683,I259632,I259621,);
not I_15143 (I260159,I2690);
DFFARX1 I_15144 (I1057275,I2683,I260159,I260185,);
nand I_15145 (I260193,I1057254,I1057254);
and I_15146 (I260210,I260193,I1057281);
DFFARX1 I_15147 (I260210,I2683,I260159,I260236,);
nor I_15148 (I260127,I260236,I260185);
not I_15149 (I260258,I260236);
DFFARX1 I_15150 (I1057269,I2683,I260159,I260284,);
nand I_15151 (I260292,I260284,I1057272);
not I_15152 (I260309,I260292);
DFFARX1 I_15153 (I260309,I2683,I260159,I260335,);
not I_15154 (I260151,I260335);
nor I_15155 (I260357,I260185,I260292);
nor I_15156 (I260133,I260236,I260357);
DFFARX1 I_15157 (I1057263,I2683,I260159,I260397,);
DFFARX1 I_15158 (I260397,I2683,I260159,I260414,);
not I_15159 (I260422,I260414);
not I_15160 (I260439,I260397);
nand I_15161 (I260136,I260439,I260258);
nand I_15162 (I260470,I1057260,I1057257);
and I_15163 (I260487,I260470,I1057278);
DFFARX1 I_15164 (I260487,I2683,I260159,I260513,);
nor I_15165 (I260521,I260513,I260185);
DFFARX1 I_15166 (I260521,I2683,I260159,I260124,);
DFFARX1 I_15167 (I260513,I2683,I260159,I260142,);
nor I_15168 (I260566,I1057266,I1057257);
not I_15169 (I260583,I260566);
nor I_15170 (I260145,I260422,I260583);
nand I_15171 (I260130,I260439,I260583);
nor I_15172 (I260139,I260185,I260566);
DFFARX1 I_15173 (I260566,I2683,I260159,I260148,);
not I_15174 (I260686,I2690);
DFFARX1 I_15175 (I802954,I2683,I260686,I260712,);
nand I_15176 (I260720,I802951,I802954);
and I_15177 (I260737,I260720,I802963);
DFFARX1 I_15178 (I260737,I2683,I260686,I260763,);
nor I_15179 (I260654,I260763,I260712);
not I_15180 (I260785,I260763);
DFFARX1 I_15181 (I802951,I2683,I260686,I260811,);
nand I_15182 (I260819,I260811,I802969);
not I_15183 (I260836,I260819);
DFFARX1 I_15184 (I260836,I2683,I260686,I260862,);
not I_15185 (I260678,I260862);
nor I_15186 (I260884,I260712,I260819);
nor I_15187 (I260660,I260763,I260884);
DFFARX1 I_15188 (I802957,I2683,I260686,I260924,);
DFFARX1 I_15189 (I260924,I2683,I260686,I260941,);
not I_15190 (I260949,I260941);
not I_15191 (I260966,I260924);
nand I_15192 (I260663,I260966,I260785);
nand I_15193 (I260997,I802966,I802972);
and I_15194 (I261014,I260997,I802957);
DFFARX1 I_15195 (I261014,I2683,I260686,I261040,);
nor I_15196 (I261048,I261040,I260712);
DFFARX1 I_15197 (I261048,I2683,I260686,I260651,);
DFFARX1 I_15198 (I261040,I2683,I260686,I260669,);
nor I_15199 (I261093,I802960,I802972);
not I_15200 (I261110,I261093);
nor I_15201 (I260672,I260949,I261110);
nand I_15202 (I260657,I260966,I261110);
nor I_15203 (I260666,I260712,I261093);
DFFARX1 I_15204 (I261093,I2683,I260686,I260675,);
not I_15205 (I261213,I2690);
DFFARX1 I_15206 (I100684,I2683,I261213,I261239,);
nand I_15207 (I261247,I100696,I100705);
and I_15208 (I261264,I261247,I100684);
DFFARX1 I_15209 (I261264,I2683,I261213,I261290,);
nor I_15210 (I261181,I261290,I261239);
not I_15211 (I261312,I261290);
DFFARX1 I_15212 (I100699,I2683,I261213,I261338,);
nand I_15213 (I261346,I261338,I100687);
not I_15214 (I261363,I261346);
DFFARX1 I_15215 (I261363,I2683,I261213,I261389,);
not I_15216 (I261205,I261389);
nor I_15217 (I261411,I261239,I261346);
nor I_15218 (I261187,I261290,I261411);
DFFARX1 I_15219 (I100690,I2683,I261213,I261451,);
DFFARX1 I_15220 (I261451,I2683,I261213,I261468,);
not I_15221 (I261476,I261468);
not I_15222 (I261493,I261451);
nand I_15223 (I261190,I261493,I261312);
nand I_15224 (I261524,I100681,I100681);
and I_15225 (I261541,I261524,I100693);
DFFARX1 I_15226 (I261541,I2683,I261213,I261567,);
nor I_15227 (I261575,I261567,I261239);
DFFARX1 I_15228 (I261575,I2683,I261213,I261178,);
DFFARX1 I_15229 (I261567,I2683,I261213,I261196,);
nor I_15230 (I261620,I100702,I100681);
not I_15231 (I261637,I261620);
nor I_15232 (I261199,I261476,I261637);
nand I_15233 (I261184,I261493,I261637);
nor I_15234 (I261193,I261239,I261620);
DFFARX1 I_15235 (I261620,I2683,I261213,I261202,);
not I_15236 (I261740,I2690);
DFFARX1 I_15237 (I458427,I2683,I261740,I261766,);
nand I_15238 (I261774,I458412,I458415);
and I_15239 (I261791,I261774,I458430);
DFFARX1 I_15240 (I261791,I2683,I261740,I261817,);
nor I_15241 (I261708,I261817,I261766);
not I_15242 (I261839,I261817);
DFFARX1 I_15243 (I458424,I2683,I261740,I261865,);
nand I_15244 (I261873,I261865,I458415);
not I_15245 (I261890,I261873);
DFFARX1 I_15246 (I261890,I2683,I261740,I261916,);
not I_15247 (I261732,I261916);
nor I_15248 (I261938,I261766,I261873);
nor I_15249 (I261714,I261817,I261938);
DFFARX1 I_15250 (I458421,I2683,I261740,I261978,);
DFFARX1 I_15251 (I261978,I2683,I261740,I261995,);
not I_15252 (I262003,I261995);
not I_15253 (I262020,I261978);
nand I_15254 (I261717,I262020,I261839);
nand I_15255 (I262051,I458436,I458412);
and I_15256 (I262068,I262051,I458433);
DFFARX1 I_15257 (I262068,I2683,I261740,I262094,);
nor I_15258 (I262102,I262094,I261766);
DFFARX1 I_15259 (I262102,I2683,I261740,I261705,);
DFFARX1 I_15260 (I262094,I2683,I261740,I261723,);
nor I_15261 (I262147,I458418,I458412);
not I_15262 (I262164,I262147);
nor I_15263 (I261726,I262003,I262164);
nand I_15264 (I261711,I262020,I262164);
nor I_15265 (I261720,I261766,I262147);
DFFARX1 I_15266 (I262147,I2683,I261740,I261729,);
not I_15267 (I262267,I2690);
DFFARX1 I_15268 (I387262,I2683,I262267,I262293,);
nand I_15269 (I262301,I387274,I387253);
and I_15270 (I262318,I262301,I387277);
DFFARX1 I_15271 (I262318,I2683,I262267,I262344,);
nor I_15272 (I262235,I262344,I262293);
not I_15273 (I262366,I262344);
DFFARX1 I_15274 (I387268,I2683,I262267,I262392,);
nand I_15275 (I262400,I262392,I387250);
not I_15276 (I262417,I262400);
DFFARX1 I_15277 (I262417,I2683,I262267,I262443,);
not I_15278 (I262259,I262443);
nor I_15279 (I262465,I262293,I262400);
nor I_15280 (I262241,I262344,I262465);
DFFARX1 I_15281 (I387265,I2683,I262267,I262505,);
DFFARX1 I_15282 (I262505,I2683,I262267,I262522,);
not I_15283 (I262530,I262522);
not I_15284 (I262547,I262505);
nand I_15285 (I262244,I262547,I262366);
nand I_15286 (I262578,I387250,I387256);
and I_15287 (I262595,I262578,I387259);
DFFARX1 I_15288 (I262595,I2683,I262267,I262621,);
nor I_15289 (I262629,I262621,I262293);
DFFARX1 I_15290 (I262629,I2683,I262267,I262232,);
DFFARX1 I_15291 (I262621,I2683,I262267,I262250,);
nor I_15292 (I262674,I387271,I387256);
not I_15293 (I262691,I262674);
nor I_15294 (I262253,I262530,I262691);
nand I_15295 (I262238,I262547,I262691);
nor I_15296 (I262247,I262293,I262674);
DFFARX1 I_15297 (I262674,I2683,I262267,I262256,);
not I_15298 (I262794,I2690);
DFFARX1 I_15299 (I171180,I2683,I262794,I262820,);
nand I_15300 (I262828,I171180,I171186);
and I_15301 (I262845,I262828,I171204);
DFFARX1 I_15302 (I262845,I2683,I262794,I262871,);
nor I_15303 (I262762,I262871,I262820);
not I_15304 (I262893,I262871);
DFFARX1 I_15305 (I171192,I2683,I262794,I262919,);
nand I_15306 (I262927,I262919,I171189);
not I_15307 (I262944,I262927);
DFFARX1 I_15308 (I262944,I2683,I262794,I262970,);
not I_15309 (I262786,I262970);
nor I_15310 (I262992,I262820,I262927);
nor I_15311 (I262768,I262871,I262992);
DFFARX1 I_15312 (I171198,I2683,I262794,I263032,);
DFFARX1 I_15313 (I263032,I2683,I262794,I263049,);
not I_15314 (I263057,I263049);
not I_15315 (I263074,I263032);
nand I_15316 (I262771,I263074,I262893);
nand I_15317 (I263105,I171183,I171183);
and I_15318 (I263122,I263105,I171195);
DFFARX1 I_15319 (I263122,I2683,I262794,I263148,);
nor I_15320 (I263156,I263148,I262820);
DFFARX1 I_15321 (I263156,I2683,I262794,I262759,);
DFFARX1 I_15322 (I263148,I2683,I262794,I262777,);
nor I_15323 (I263201,I171201,I171183);
not I_15324 (I263218,I263201);
nor I_15325 (I262780,I263057,I263218);
nand I_15326 (I262765,I263074,I263218);
nor I_15327 (I262774,I262820,I263201);
DFFARX1 I_15328 (I263201,I2683,I262794,I262783,);
not I_15329 (I263321,I2690);
DFFARX1 I_15330 (I734206,I2683,I263321,I263347,);
nand I_15331 (I263355,I734203,I734221);
and I_15332 (I263372,I263355,I734212);
DFFARX1 I_15333 (I263372,I2683,I263321,I263398,);
nor I_15334 (I263289,I263398,I263347);
not I_15335 (I263420,I263398);
DFFARX1 I_15336 (I734227,I2683,I263321,I263446,);
nand I_15337 (I263454,I263446,I734209);
not I_15338 (I263471,I263454);
DFFARX1 I_15339 (I263471,I2683,I263321,I263497,);
not I_15340 (I263313,I263497);
nor I_15341 (I263519,I263347,I263454);
nor I_15342 (I263295,I263398,I263519);
DFFARX1 I_15343 (I734215,I2683,I263321,I263559,);
DFFARX1 I_15344 (I263559,I2683,I263321,I263576,);
not I_15345 (I263584,I263576);
not I_15346 (I263601,I263559);
nand I_15347 (I263298,I263601,I263420);
nand I_15348 (I263632,I734203,I734230);
and I_15349 (I263649,I263632,I734218);
DFFARX1 I_15350 (I263649,I2683,I263321,I263675,);
nor I_15351 (I263683,I263675,I263347);
DFFARX1 I_15352 (I263683,I2683,I263321,I263286,);
DFFARX1 I_15353 (I263675,I2683,I263321,I263304,);
nor I_15354 (I263728,I734224,I734230);
not I_15355 (I263745,I263728);
nor I_15356 (I263307,I263584,I263745);
nand I_15357 (I263292,I263601,I263745);
nor I_15358 (I263301,I263347,I263728);
DFFARX1 I_15359 (I263728,I2683,I263321,I263310,);
not I_15360 (I263848,I2690);
DFFARX1 I_15361 (I741312,I2683,I263848,I263874,);
nand I_15362 (I263882,I741309,I741327);
and I_15363 (I263899,I263882,I741318);
DFFARX1 I_15364 (I263899,I2683,I263848,I263925,);
nor I_15365 (I263816,I263925,I263874);
not I_15366 (I263947,I263925);
DFFARX1 I_15367 (I741333,I2683,I263848,I263973,);
nand I_15368 (I263981,I263973,I741315);
not I_15369 (I263998,I263981);
DFFARX1 I_15370 (I263998,I2683,I263848,I264024,);
not I_15371 (I263840,I264024);
nor I_15372 (I264046,I263874,I263981);
nor I_15373 (I263822,I263925,I264046);
DFFARX1 I_15374 (I741321,I2683,I263848,I264086,);
DFFARX1 I_15375 (I264086,I2683,I263848,I264103,);
not I_15376 (I264111,I264103);
not I_15377 (I264128,I264086);
nand I_15378 (I263825,I264128,I263947);
nand I_15379 (I264159,I741309,I741336);
and I_15380 (I264176,I264159,I741324);
DFFARX1 I_15381 (I264176,I2683,I263848,I264202,);
nor I_15382 (I264210,I264202,I263874);
DFFARX1 I_15383 (I264210,I2683,I263848,I263813,);
DFFARX1 I_15384 (I264202,I2683,I263848,I263831,);
nor I_15385 (I264255,I741330,I741336);
not I_15386 (I264272,I264255);
nor I_15387 (I263834,I264111,I264272);
nand I_15388 (I263819,I264128,I264272);
nor I_15389 (I263828,I263874,I264255);
DFFARX1 I_15390 (I264255,I2683,I263848,I263837,);
not I_15391 (I264375,I2690);
DFFARX1 I_15392 (I501196,I2683,I264375,I264401,);
nand I_15393 (I264409,I501187,I501202);
and I_15394 (I264426,I264409,I501208);
DFFARX1 I_15395 (I264426,I2683,I264375,I264452,);
nor I_15396 (I264343,I264452,I264401);
not I_15397 (I264474,I264452);
DFFARX1 I_15398 (I501193,I2683,I264375,I264500,);
nand I_15399 (I264508,I264500,I501187);
not I_15400 (I264525,I264508);
DFFARX1 I_15401 (I264525,I2683,I264375,I264551,);
not I_15402 (I264367,I264551);
nor I_15403 (I264573,I264401,I264508);
nor I_15404 (I264349,I264452,I264573);
DFFARX1 I_15405 (I501190,I2683,I264375,I264613,);
DFFARX1 I_15406 (I264613,I2683,I264375,I264630,);
not I_15407 (I264638,I264630);
not I_15408 (I264655,I264613);
nand I_15409 (I264352,I264655,I264474);
nand I_15410 (I264686,I501184,I501199);
and I_15411 (I264703,I264686,I501184);
DFFARX1 I_15412 (I264703,I2683,I264375,I264729,);
nor I_15413 (I264737,I264729,I264401);
DFFARX1 I_15414 (I264737,I2683,I264375,I264340,);
DFFARX1 I_15415 (I264729,I2683,I264375,I264358,);
nor I_15416 (I264782,I501205,I501199);
not I_15417 (I264799,I264782);
nor I_15418 (I264361,I264638,I264799);
nand I_15419 (I264346,I264655,I264799);
nor I_15420 (I264355,I264401,I264782);
DFFARX1 I_15421 (I264782,I2683,I264375,I264364,);
not I_15422 (I264902,I2690);
DFFARX1 I_15423 (I188435,I2683,I264902,I264928,);
nand I_15424 (I264936,I188435,I188441);
and I_15425 (I264953,I264936,I188459);
DFFARX1 I_15426 (I264953,I2683,I264902,I264979,);
nor I_15427 (I264870,I264979,I264928);
not I_15428 (I265001,I264979);
DFFARX1 I_15429 (I188447,I2683,I264902,I265027,);
nand I_15430 (I265035,I265027,I188444);
not I_15431 (I265052,I265035);
DFFARX1 I_15432 (I265052,I2683,I264902,I265078,);
not I_15433 (I264894,I265078);
nor I_15434 (I265100,I264928,I265035);
nor I_15435 (I264876,I264979,I265100);
DFFARX1 I_15436 (I188453,I2683,I264902,I265140,);
DFFARX1 I_15437 (I265140,I2683,I264902,I265157,);
not I_15438 (I265165,I265157);
not I_15439 (I265182,I265140);
nand I_15440 (I264879,I265182,I265001);
nand I_15441 (I265213,I188438,I188438);
and I_15442 (I265230,I265213,I188450);
DFFARX1 I_15443 (I265230,I2683,I264902,I265256,);
nor I_15444 (I265264,I265256,I264928);
DFFARX1 I_15445 (I265264,I2683,I264902,I264867,);
DFFARX1 I_15446 (I265256,I2683,I264902,I264885,);
nor I_15447 (I265309,I188456,I188438);
not I_15448 (I265326,I265309);
nor I_15449 (I264888,I265165,I265326);
nand I_15450 (I264873,I265182,I265326);
nor I_15451 (I264882,I264928,I265309);
DFFARX1 I_15452 (I265309,I2683,I264902,I264891,);
not I_15453 (I265429,I2690);
DFFARX1 I_15454 (I137265,I2683,I265429,I265455,);
nand I_15455 (I265463,I137265,I137271);
and I_15456 (I265480,I265463,I137289);
DFFARX1 I_15457 (I265480,I2683,I265429,I265506,);
nor I_15458 (I265397,I265506,I265455);
not I_15459 (I265528,I265506);
DFFARX1 I_15460 (I137277,I2683,I265429,I265554,);
nand I_15461 (I265562,I265554,I137274);
not I_15462 (I265579,I265562);
DFFARX1 I_15463 (I265579,I2683,I265429,I265605,);
not I_15464 (I265421,I265605);
nor I_15465 (I265627,I265455,I265562);
nor I_15466 (I265403,I265506,I265627);
DFFARX1 I_15467 (I137283,I2683,I265429,I265667,);
DFFARX1 I_15468 (I265667,I2683,I265429,I265684,);
not I_15469 (I265692,I265684);
not I_15470 (I265709,I265667);
nand I_15471 (I265406,I265709,I265528);
nand I_15472 (I265740,I137268,I137268);
and I_15473 (I265757,I265740,I137280);
DFFARX1 I_15474 (I265757,I2683,I265429,I265783,);
nor I_15475 (I265791,I265783,I265455);
DFFARX1 I_15476 (I265791,I2683,I265429,I265394,);
DFFARX1 I_15477 (I265783,I2683,I265429,I265412,);
nor I_15478 (I265836,I137286,I137268);
not I_15479 (I265853,I265836);
nor I_15480 (I265415,I265692,I265853);
nand I_15481 (I265400,I265709,I265853);
nor I_15482 (I265409,I265455,I265836);
DFFARX1 I_15483 (I265836,I2683,I265429,I265418,);
not I_15484 (I265956,I2690);
DFFARX1 I_15485 (I807442,I2683,I265956,I265982,);
nand I_15486 (I265990,I807439,I807442);
and I_15487 (I266007,I265990,I807451);
DFFARX1 I_15488 (I266007,I2683,I265956,I266033,);
nor I_15489 (I265924,I266033,I265982);
not I_15490 (I266055,I266033);
DFFARX1 I_15491 (I807439,I2683,I265956,I266081,);
nand I_15492 (I266089,I266081,I807457);
not I_15493 (I266106,I266089);
DFFARX1 I_15494 (I266106,I2683,I265956,I266132,);
not I_15495 (I265948,I266132);
nor I_15496 (I266154,I265982,I266089);
nor I_15497 (I265930,I266033,I266154);
DFFARX1 I_15498 (I807445,I2683,I265956,I266194,);
DFFARX1 I_15499 (I266194,I2683,I265956,I266211,);
not I_15500 (I266219,I266211);
not I_15501 (I266236,I266194);
nand I_15502 (I265933,I266236,I266055);
nand I_15503 (I266267,I807454,I807460);
and I_15504 (I266284,I266267,I807445);
DFFARX1 I_15505 (I266284,I2683,I265956,I266310,);
nor I_15506 (I266318,I266310,I265982);
DFFARX1 I_15507 (I266318,I2683,I265956,I265921,);
DFFARX1 I_15508 (I266310,I2683,I265956,I265939,);
nor I_15509 (I266363,I807448,I807460);
not I_15510 (I266380,I266363);
nor I_15511 (I265942,I266219,I266380);
nand I_15512 (I265927,I266236,I266380);
nor I_15513 (I265936,I265982,I266363);
DFFARX1 I_15514 (I266363,I2683,I265956,I265945,);
not I_15515 (I266483,I2690);
DFFARX1 I_15516 (I778134,I2683,I266483,I266509,);
nand I_15517 (I266517,I778131,I778149);
and I_15518 (I266534,I266517,I778140);
DFFARX1 I_15519 (I266534,I2683,I266483,I266560,);
nor I_15520 (I266451,I266560,I266509);
not I_15521 (I266582,I266560);
DFFARX1 I_15522 (I778155,I2683,I266483,I266608,);
nand I_15523 (I266616,I266608,I778137);
not I_15524 (I266633,I266616);
DFFARX1 I_15525 (I266633,I2683,I266483,I266659,);
not I_15526 (I266475,I266659);
nor I_15527 (I266681,I266509,I266616);
nor I_15528 (I266457,I266560,I266681);
DFFARX1 I_15529 (I778143,I2683,I266483,I266721,);
DFFARX1 I_15530 (I266721,I2683,I266483,I266738,);
not I_15531 (I266746,I266738);
not I_15532 (I266763,I266721);
nand I_15533 (I266460,I266763,I266582);
nand I_15534 (I266794,I778131,I778158);
and I_15535 (I266811,I266794,I778146);
DFFARX1 I_15536 (I266811,I2683,I266483,I266837,);
nor I_15537 (I266845,I266837,I266509);
DFFARX1 I_15538 (I266845,I2683,I266483,I266448,);
DFFARX1 I_15539 (I266837,I2683,I266483,I266466,);
nor I_15540 (I266890,I778152,I778158);
not I_15541 (I266907,I266890);
nor I_15542 (I266469,I266746,I266907);
nand I_15543 (I266454,I266763,I266907);
nor I_15544 (I266463,I266509,I266890);
DFFARX1 I_15545 (I266890,I2683,I266483,I266472,);
not I_15546 (I267010,I2690);
DFFARX1 I_15547 (I567666,I2683,I267010,I267036,);
nand I_15548 (I267044,I567657,I567672);
and I_15549 (I267061,I267044,I567678);
DFFARX1 I_15550 (I267061,I2683,I267010,I267087,);
nor I_15551 (I266978,I267087,I267036);
not I_15552 (I267109,I267087);
DFFARX1 I_15553 (I567663,I2683,I267010,I267135,);
nand I_15554 (I267143,I267135,I567657);
not I_15555 (I267160,I267143);
DFFARX1 I_15556 (I267160,I2683,I267010,I267186,);
not I_15557 (I267002,I267186);
nor I_15558 (I267208,I267036,I267143);
nor I_15559 (I266984,I267087,I267208);
DFFARX1 I_15560 (I567660,I2683,I267010,I267248,);
DFFARX1 I_15561 (I267248,I2683,I267010,I267265,);
not I_15562 (I267273,I267265);
not I_15563 (I267290,I267248);
nand I_15564 (I266987,I267290,I267109);
nand I_15565 (I267321,I567654,I567669);
and I_15566 (I267338,I267321,I567654);
DFFARX1 I_15567 (I267338,I2683,I267010,I267364,);
nor I_15568 (I267372,I267364,I267036);
DFFARX1 I_15569 (I267372,I2683,I267010,I266975,);
DFFARX1 I_15570 (I267364,I2683,I267010,I266993,);
nor I_15571 (I267417,I567675,I567669);
not I_15572 (I267434,I267417);
nor I_15573 (I266996,I267273,I267434);
nand I_15574 (I266981,I267290,I267434);
nor I_15575 (I266990,I267036,I267417);
DFFARX1 I_15576 (I267417,I2683,I267010,I266999,);
not I_15577 (I267537,I2690);
DFFARX1 I_15578 (I791054,I2683,I267537,I267563,);
nand I_15579 (I267571,I791051,I791069);
and I_15580 (I267588,I267571,I791060);
DFFARX1 I_15581 (I267588,I2683,I267537,I267614,);
nor I_15582 (I267505,I267614,I267563);
not I_15583 (I267636,I267614);
DFFARX1 I_15584 (I791075,I2683,I267537,I267662,);
nand I_15585 (I267670,I267662,I791057);
not I_15586 (I267687,I267670);
DFFARX1 I_15587 (I267687,I2683,I267537,I267713,);
not I_15588 (I267529,I267713);
nor I_15589 (I267735,I267563,I267670);
nor I_15590 (I267511,I267614,I267735);
DFFARX1 I_15591 (I791063,I2683,I267537,I267775,);
DFFARX1 I_15592 (I267775,I2683,I267537,I267792,);
not I_15593 (I267800,I267792);
not I_15594 (I267817,I267775);
nand I_15595 (I267514,I267817,I267636);
nand I_15596 (I267848,I791051,I791078);
and I_15597 (I267865,I267848,I791066);
DFFARX1 I_15598 (I267865,I2683,I267537,I267891,);
nor I_15599 (I267899,I267891,I267563);
DFFARX1 I_15600 (I267899,I2683,I267537,I267502,);
DFFARX1 I_15601 (I267891,I2683,I267537,I267520,);
nor I_15602 (I267944,I791072,I791078);
not I_15603 (I267961,I267944);
nor I_15604 (I267523,I267800,I267961);
nand I_15605 (I267508,I267817,I267961);
nor I_15606 (I267517,I267563,I267944);
DFFARX1 I_15607 (I267944,I2683,I267537,I267526,);
not I_15608 (I268064,I2690);
DFFARX1 I_15609 (I1084645,I2683,I268064,I268090,);
nand I_15610 (I268098,I1084624,I1084624);
and I_15611 (I268115,I268098,I1084651);
DFFARX1 I_15612 (I268115,I2683,I268064,I268141,);
nor I_15613 (I268032,I268141,I268090);
not I_15614 (I268163,I268141);
DFFARX1 I_15615 (I1084639,I2683,I268064,I268189,);
nand I_15616 (I268197,I268189,I1084642);
not I_15617 (I268214,I268197);
DFFARX1 I_15618 (I268214,I2683,I268064,I268240,);
not I_15619 (I268056,I268240);
nor I_15620 (I268262,I268090,I268197);
nor I_15621 (I268038,I268141,I268262);
DFFARX1 I_15622 (I1084633,I2683,I268064,I268302,);
DFFARX1 I_15623 (I268302,I2683,I268064,I268319,);
not I_15624 (I268327,I268319);
not I_15625 (I268344,I268302);
nand I_15626 (I268041,I268344,I268163);
nand I_15627 (I268375,I1084630,I1084627);
and I_15628 (I268392,I268375,I1084648);
DFFARX1 I_15629 (I268392,I2683,I268064,I268418,);
nor I_15630 (I268426,I268418,I268090);
DFFARX1 I_15631 (I268426,I2683,I268064,I268029,);
DFFARX1 I_15632 (I268418,I2683,I268064,I268047,);
nor I_15633 (I268471,I1084636,I1084627);
not I_15634 (I268488,I268471);
nor I_15635 (I268050,I268327,I268488);
nand I_15636 (I268035,I268344,I268488);
nor I_15637 (I268044,I268090,I268471);
DFFARX1 I_15638 (I268471,I2683,I268064,I268053,);
not I_15639 (I268591,I2690);
DFFARX1 I_15640 (I1037640,I2683,I268591,I268617,);
nand I_15641 (I268625,I1037619,I1037619);
and I_15642 (I268642,I268625,I1037646);
DFFARX1 I_15643 (I268642,I2683,I268591,I268668,);
nor I_15644 (I268559,I268668,I268617);
not I_15645 (I268690,I268668);
DFFARX1 I_15646 (I1037634,I2683,I268591,I268716,);
nand I_15647 (I268724,I268716,I1037637);
not I_15648 (I268741,I268724);
DFFARX1 I_15649 (I268741,I2683,I268591,I268767,);
not I_15650 (I268583,I268767);
nor I_15651 (I268789,I268617,I268724);
nor I_15652 (I268565,I268668,I268789);
DFFARX1 I_15653 (I1037628,I2683,I268591,I268829,);
DFFARX1 I_15654 (I268829,I2683,I268591,I268846,);
not I_15655 (I268854,I268846);
not I_15656 (I268871,I268829);
nand I_15657 (I268568,I268871,I268690);
nand I_15658 (I268902,I1037625,I1037622);
and I_15659 (I268919,I268902,I1037643);
DFFARX1 I_15660 (I268919,I2683,I268591,I268945,);
nor I_15661 (I268953,I268945,I268617);
DFFARX1 I_15662 (I268953,I2683,I268591,I268556,);
DFFARX1 I_15663 (I268945,I2683,I268591,I268574,);
nor I_15664 (I268998,I1037631,I1037622);
not I_15665 (I269015,I268998);
nor I_15666 (I268577,I268854,I269015);
nand I_15667 (I268562,I268871,I269015);
nor I_15668 (I268571,I268617,I268998);
DFFARX1 I_15669 (I268998,I2683,I268591,I268580,);
not I_15670 (I269118,I2690);
DFFARX1 I_15671 (I972272,I2683,I269118,I269144,);
nand I_15672 (I269152,I972254,I972278);
and I_15673 (I269169,I269152,I972269);
DFFARX1 I_15674 (I269169,I2683,I269118,I269195,);
nor I_15675 (I269086,I269195,I269144);
not I_15676 (I269217,I269195);
DFFARX1 I_15677 (I972275,I2683,I269118,I269243,);
nand I_15678 (I269251,I269243,I972263);
not I_15679 (I269268,I269251);
DFFARX1 I_15680 (I269268,I2683,I269118,I269294,);
not I_15681 (I269110,I269294);
nor I_15682 (I269316,I269144,I269251);
nor I_15683 (I269092,I269195,I269316);
DFFARX1 I_15684 (I972254,I2683,I269118,I269356,);
DFFARX1 I_15685 (I269356,I2683,I269118,I269373,);
not I_15686 (I269381,I269373);
not I_15687 (I269398,I269356);
nand I_15688 (I269095,I269398,I269217);
nand I_15689 (I269429,I972260,I972257);
and I_15690 (I269446,I269429,I972266);
DFFARX1 I_15691 (I269446,I2683,I269118,I269472,);
nor I_15692 (I269480,I269472,I269144);
DFFARX1 I_15693 (I269480,I2683,I269118,I269083,);
DFFARX1 I_15694 (I269472,I2683,I269118,I269101,);
nor I_15695 (I269525,I972257,I972257);
not I_15696 (I269542,I269525);
nor I_15697 (I269104,I269381,I269542);
nand I_15698 (I269089,I269398,I269542);
nor I_15699 (I269098,I269144,I269525);
DFFARX1 I_15700 (I269525,I2683,I269118,I269107,);
not I_15701 (I269645,I2690);
DFFARX1 I_15702 (I634909,I2683,I269645,I269671,);
nand I_15703 (I269679,I634912,I634906);
and I_15704 (I269696,I269679,I634918);
DFFARX1 I_15705 (I269696,I2683,I269645,I269722,);
nor I_15706 (I269613,I269722,I269671);
not I_15707 (I269744,I269722);
DFFARX1 I_15708 (I634921,I2683,I269645,I269770,);
nand I_15709 (I269778,I269770,I634912);
not I_15710 (I269795,I269778);
DFFARX1 I_15711 (I269795,I2683,I269645,I269821,);
not I_15712 (I269637,I269821);
nor I_15713 (I269843,I269671,I269778);
nor I_15714 (I269619,I269722,I269843);
DFFARX1 I_15715 (I634924,I2683,I269645,I269883,);
DFFARX1 I_15716 (I269883,I2683,I269645,I269900,);
not I_15717 (I269908,I269900);
not I_15718 (I269925,I269883);
nand I_15719 (I269622,I269925,I269744);
nand I_15720 (I269956,I634906,I634915);
and I_15721 (I269973,I269956,I634909);
DFFARX1 I_15722 (I269973,I2683,I269645,I269999,);
nor I_15723 (I270007,I269999,I269671);
DFFARX1 I_15724 (I270007,I2683,I269645,I269610,);
DFFARX1 I_15725 (I269999,I2683,I269645,I269628,);
nor I_15726 (I270052,I634927,I634915);
not I_15727 (I270069,I270052);
nor I_15728 (I269631,I269908,I270069);
nand I_15729 (I269616,I269925,I270069);
nor I_15730 (I269625,I269671,I270052);
DFFARX1 I_15731 (I270052,I2683,I269645,I269634,);
not I_15732 (I270172,I2690);
DFFARX1 I_15733 (I339390,I2683,I270172,I270198,);
nand I_15734 (I270206,I339402,I339381);
and I_15735 (I270223,I270206,I339405);
DFFARX1 I_15736 (I270223,I2683,I270172,I270249,);
nor I_15737 (I270140,I270249,I270198);
not I_15738 (I270271,I270249);
DFFARX1 I_15739 (I339396,I2683,I270172,I270297,);
nand I_15740 (I270305,I270297,I339378);
not I_15741 (I270322,I270305);
DFFARX1 I_15742 (I270322,I2683,I270172,I270348,);
not I_15743 (I270164,I270348);
nor I_15744 (I270370,I270198,I270305);
nor I_15745 (I270146,I270249,I270370);
DFFARX1 I_15746 (I339393,I2683,I270172,I270410,);
DFFARX1 I_15747 (I270410,I2683,I270172,I270427,);
not I_15748 (I270435,I270427);
not I_15749 (I270452,I270410);
nand I_15750 (I270149,I270452,I270271);
nand I_15751 (I270483,I339378,I339384);
and I_15752 (I270500,I270483,I339387);
DFFARX1 I_15753 (I270500,I2683,I270172,I270526,);
nor I_15754 (I270534,I270526,I270198);
DFFARX1 I_15755 (I270534,I2683,I270172,I270137,);
DFFARX1 I_15756 (I270526,I2683,I270172,I270155,);
nor I_15757 (I270579,I339399,I339384);
not I_15758 (I270596,I270579);
nor I_15759 (I270158,I270435,I270596);
nand I_15760 (I270143,I270452,I270596);
nor I_15761 (I270152,I270198,I270579);
DFFARX1 I_15762 (I270579,I2683,I270172,I270161,);
not I_15763 (I270699,I2690);
DFFARX1 I_15764 (I479235,I2683,I270699,I270725,);
nand I_15765 (I270733,I479220,I479223);
and I_15766 (I270750,I270733,I479238);
DFFARX1 I_15767 (I270750,I2683,I270699,I270776,);
nor I_15768 (I270667,I270776,I270725);
not I_15769 (I270798,I270776);
DFFARX1 I_15770 (I479232,I2683,I270699,I270824,);
nand I_15771 (I270832,I270824,I479223);
not I_15772 (I270849,I270832);
DFFARX1 I_15773 (I270849,I2683,I270699,I270875,);
not I_15774 (I270691,I270875);
nor I_15775 (I270897,I270725,I270832);
nor I_15776 (I270673,I270776,I270897);
DFFARX1 I_15777 (I479229,I2683,I270699,I270937,);
DFFARX1 I_15778 (I270937,I2683,I270699,I270954,);
not I_15779 (I270962,I270954);
not I_15780 (I270979,I270937);
nand I_15781 (I270676,I270979,I270798);
nand I_15782 (I271010,I479244,I479220);
and I_15783 (I271027,I271010,I479241);
DFFARX1 I_15784 (I271027,I2683,I270699,I271053,);
nor I_15785 (I271061,I271053,I270725);
DFFARX1 I_15786 (I271061,I2683,I270699,I270664,);
DFFARX1 I_15787 (I271053,I2683,I270699,I270682,);
nor I_15788 (I271106,I479226,I479220);
not I_15789 (I271123,I271106);
nor I_15790 (I270685,I270962,I271123);
nand I_15791 (I270670,I270979,I271123);
nor I_15792 (I270679,I270725,I271106);
DFFARX1 I_15793 (I271106,I2683,I270699,I270688,);
not I_15794 (I271226,I2690);
DFFARX1 I_15795 (I440509,I2683,I271226,I271252,);
nand I_15796 (I271260,I440494,I440497);
and I_15797 (I271277,I271260,I440512);
DFFARX1 I_15798 (I271277,I2683,I271226,I271303,);
nor I_15799 (I271194,I271303,I271252);
not I_15800 (I271325,I271303);
DFFARX1 I_15801 (I440506,I2683,I271226,I271351,);
nand I_15802 (I271359,I271351,I440497);
not I_15803 (I271376,I271359);
DFFARX1 I_15804 (I271376,I2683,I271226,I271402,);
not I_15805 (I271218,I271402);
nor I_15806 (I271424,I271252,I271359);
nor I_15807 (I271200,I271303,I271424);
DFFARX1 I_15808 (I440503,I2683,I271226,I271464,);
DFFARX1 I_15809 (I271464,I2683,I271226,I271481,);
not I_15810 (I271489,I271481);
not I_15811 (I271506,I271464);
nand I_15812 (I271203,I271506,I271325);
nand I_15813 (I271537,I440518,I440494);
and I_15814 (I271554,I271537,I440515);
DFFARX1 I_15815 (I271554,I2683,I271226,I271580,);
nor I_15816 (I271588,I271580,I271252);
DFFARX1 I_15817 (I271588,I2683,I271226,I271191,);
DFFARX1 I_15818 (I271580,I2683,I271226,I271209,);
nor I_15819 (I271633,I440500,I440494);
not I_15820 (I271650,I271633);
nor I_15821 (I271212,I271489,I271650);
nand I_15822 (I271197,I271506,I271650);
nor I_15823 (I271206,I271252,I271633);
DFFARX1 I_15824 (I271633,I2683,I271226,I271215,);
not I_15825 (I271753,I2690);
DFFARX1 I_15826 (I690244,I2683,I271753,I271779,);
nand I_15827 (I271787,I690247,I690241);
and I_15828 (I271804,I271787,I690253);
DFFARX1 I_15829 (I271804,I2683,I271753,I271830,);
nor I_15830 (I271721,I271830,I271779);
not I_15831 (I271852,I271830);
DFFARX1 I_15832 (I690256,I2683,I271753,I271878,);
nand I_15833 (I271886,I271878,I690247);
not I_15834 (I271903,I271886);
DFFARX1 I_15835 (I271903,I2683,I271753,I271929,);
not I_15836 (I271745,I271929);
nor I_15837 (I271951,I271779,I271886);
nor I_15838 (I271727,I271830,I271951);
DFFARX1 I_15839 (I690259,I2683,I271753,I271991,);
DFFARX1 I_15840 (I271991,I2683,I271753,I272008,);
not I_15841 (I272016,I272008);
not I_15842 (I272033,I271991);
nand I_15843 (I271730,I272033,I271852);
nand I_15844 (I272064,I690241,I690250);
and I_15845 (I272081,I272064,I690244);
DFFARX1 I_15846 (I272081,I2683,I271753,I272107,);
nor I_15847 (I272115,I272107,I271779);
DFFARX1 I_15848 (I272115,I2683,I271753,I271718,);
DFFARX1 I_15849 (I272107,I2683,I271753,I271736,);
nor I_15850 (I272160,I690262,I690250);
not I_15851 (I272177,I272160);
nor I_15852 (I271739,I272016,I272177);
nand I_15853 (I271724,I272033,I272177);
nor I_15854 (I271733,I271779,I272160);
DFFARX1 I_15855 (I272160,I2683,I271753,I271742,);
not I_15856 (I272280,I2690);
DFFARX1 I_15857 (I76442,I2683,I272280,I272306,);
nand I_15858 (I272314,I76454,I76463);
and I_15859 (I272331,I272314,I76442);
DFFARX1 I_15860 (I272331,I2683,I272280,I272357,);
nor I_15861 (I272248,I272357,I272306);
not I_15862 (I272379,I272357);
DFFARX1 I_15863 (I76457,I2683,I272280,I272405,);
nand I_15864 (I272413,I272405,I76445);
not I_15865 (I272430,I272413);
DFFARX1 I_15866 (I272430,I2683,I272280,I272456,);
not I_15867 (I272272,I272456);
nor I_15868 (I272478,I272306,I272413);
nor I_15869 (I272254,I272357,I272478);
DFFARX1 I_15870 (I76448,I2683,I272280,I272518,);
DFFARX1 I_15871 (I272518,I2683,I272280,I272535,);
not I_15872 (I272543,I272535);
not I_15873 (I272560,I272518);
nand I_15874 (I272257,I272560,I272379);
nand I_15875 (I272591,I76439,I76439);
and I_15876 (I272608,I272591,I76451);
DFFARX1 I_15877 (I272608,I2683,I272280,I272634,);
nor I_15878 (I272642,I272634,I272306);
DFFARX1 I_15879 (I272642,I2683,I272280,I272245,);
DFFARX1 I_15880 (I272634,I2683,I272280,I272263,);
nor I_15881 (I272687,I76460,I76439);
not I_15882 (I272704,I272687);
nor I_15883 (I272266,I272543,I272704);
nand I_15884 (I272251,I272560,I272704);
nor I_15885 (I272260,I272306,I272687);
DFFARX1 I_15886 (I272687,I2683,I272280,I272269,);
not I_15887 (I272807,I2690);
DFFARX1 I_15888 (I741958,I2683,I272807,I272833,);
nand I_15889 (I272841,I741955,I741973);
and I_15890 (I272858,I272841,I741964);
DFFARX1 I_15891 (I272858,I2683,I272807,I272884,);
nor I_15892 (I272775,I272884,I272833);
not I_15893 (I272906,I272884);
DFFARX1 I_15894 (I741979,I2683,I272807,I272932,);
nand I_15895 (I272940,I272932,I741961);
not I_15896 (I272957,I272940);
DFFARX1 I_15897 (I272957,I2683,I272807,I272983,);
not I_15898 (I272799,I272983);
nor I_15899 (I273005,I272833,I272940);
nor I_15900 (I272781,I272884,I273005);
DFFARX1 I_15901 (I741967,I2683,I272807,I273045,);
DFFARX1 I_15902 (I273045,I2683,I272807,I273062,);
not I_15903 (I273070,I273062);
not I_15904 (I273087,I273045);
nand I_15905 (I272784,I273087,I272906);
nand I_15906 (I273118,I741955,I741982);
and I_15907 (I273135,I273118,I741970);
DFFARX1 I_15908 (I273135,I2683,I272807,I273161,);
nor I_15909 (I273169,I273161,I272833);
DFFARX1 I_15910 (I273169,I2683,I272807,I272772,);
DFFARX1 I_15911 (I273161,I2683,I272807,I272790,);
nor I_15912 (I273214,I741976,I741982);
not I_15913 (I273231,I273214);
nor I_15914 (I272793,I273070,I273231);
nand I_15915 (I272778,I273087,I273231);
nor I_15916 (I272787,I272833,I273214);
DFFARX1 I_15917 (I273214,I2683,I272807,I272796,);
not I_15918 (I273334,I2690);
DFFARX1 I_15919 (I370942,I2683,I273334,I273360,);
nand I_15920 (I273368,I370954,I370933);
and I_15921 (I273385,I273368,I370957);
DFFARX1 I_15922 (I273385,I2683,I273334,I273411,);
nor I_15923 (I273302,I273411,I273360);
not I_15924 (I273433,I273411);
DFFARX1 I_15925 (I370948,I2683,I273334,I273459,);
nand I_15926 (I273467,I273459,I370930);
not I_15927 (I273484,I273467);
DFFARX1 I_15928 (I273484,I2683,I273334,I273510,);
not I_15929 (I273326,I273510);
nor I_15930 (I273532,I273360,I273467);
nor I_15931 (I273308,I273411,I273532);
DFFARX1 I_15932 (I370945,I2683,I273334,I273572,);
DFFARX1 I_15933 (I273572,I2683,I273334,I273589,);
not I_15934 (I273597,I273589);
not I_15935 (I273614,I273572);
nand I_15936 (I273311,I273614,I273433);
nand I_15937 (I273645,I370930,I370936);
and I_15938 (I273662,I273645,I370939);
DFFARX1 I_15939 (I273662,I2683,I273334,I273688,);
nor I_15940 (I273696,I273688,I273360);
DFFARX1 I_15941 (I273696,I2683,I273334,I273299,);
DFFARX1 I_15942 (I273688,I2683,I273334,I273317,);
nor I_15943 (I273741,I370951,I370936);
not I_15944 (I273758,I273741);
nor I_15945 (I273320,I273597,I273758);
nand I_15946 (I273305,I273614,I273758);
nor I_15947 (I273314,I273360,I273741);
DFFARX1 I_15948 (I273741,I2683,I273334,I273323,);
not I_15949 (I273861,I2690);
DFFARX1 I_15950 (I983152,I2683,I273861,I273887,);
nand I_15951 (I273895,I983134,I983158);
and I_15952 (I273912,I273895,I983149);
DFFARX1 I_15953 (I273912,I2683,I273861,I273938,);
nor I_15954 (I273829,I273938,I273887);
not I_15955 (I273960,I273938);
DFFARX1 I_15956 (I983155,I2683,I273861,I273986,);
nand I_15957 (I273994,I273986,I983143);
not I_15958 (I274011,I273994);
DFFARX1 I_15959 (I274011,I2683,I273861,I274037,);
not I_15960 (I273853,I274037);
nor I_15961 (I274059,I273887,I273994);
nor I_15962 (I273835,I273938,I274059);
DFFARX1 I_15963 (I983134,I2683,I273861,I274099,);
DFFARX1 I_15964 (I274099,I2683,I273861,I274116,);
not I_15965 (I274124,I274116);
not I_15966 (I274141,I274099);
nand I_15967 (I273838,I274141,I273960);
nand I_15968 (I274172,I983140,I983137);
and I_15969 (I274189,I274172,I983146);
DFFARX1 I_15970 (I274189,I2683,I273861,I274215,);
nor I_15971 (I274223,I274215,I273887);
DFFARX1 I_15972 (I274223,I2683,I273861,I273826,);
DFFARX1 I_15973 (I274215,I2683,I273861,I273844,);
nor I_15974 (I274268,I983137,I983137);
not I_15975 (I274285,I274268);
nor I_15976 (I273847,I274124,I274285);
nand I_15977 (I273832,I274141,I274285);
nor I_15978 (I273841,I273887,I274268);
DFFARX1 I_15979 (I274268,I2683,I273861,I273850,);
not I_15980 (I274388,I2690);
DFFARX1 I_15981 (I743896,I2683,I274388,I274414,);
nand I_15982 (I274422,I743893,I743911);
and I_15983 (I274439,I274422,I743902);
DFFARX1 I_15984 (I274439,I2683,I274388,I274465,);
nor I_15985 (I274356,I274465,I274414);
not I_15986 (I274487,I274465);
DFFARX1 I_15987 (I743917,I2683,I274388,I274513,);
nand I_15988 (I274521,I274513,I743899);
not I_15989 (I274538,I274521);
DFFARX1 I_15990 (I274538,I2683,I274388,I274564,);
not I_15991 (I274380,I274564);
nor I_15992 (I274586,I274414,I274521);
nor I_15993 (I274362,I274465,I274586);
DFFARX1 I_15994 (I743905,I2683,I274388,I274626,);
DFFARX1 I_15995 (I274626,I2683,I274388,I274643,);
not I_15996 (I274651,I274643);
not I_15997 (I274668,I274626);
nand I_15998 (I274365,I274668,I274487);
nand I_15999 (I274699,I743893,I743920);
and I_16000 (I274716,I274699,I743908);
DFFARX1 I_16001 (I274716,I2683,I274388,I274742,);
nor I_16002 (I274750,I274742,I274414);
DFFARX1 I_16003 (I274750,I2683,I274388,I274353,);
DFFARX1 I_16004 (I274742,I2683,I274388,I274371,);
nor I_16005 (I274795,I743914,I743920);
not I_16006 (I274812,I274795);
nor I_16007 (I274374,I274651,I274812);
nand I_16008 (I274359,I274668,I274812);
nor I_16009 (I274368,I274414,I274795);
DFFARX1 I_16010 (I274795,I2683,I274388,I274377,);
not I_16011 (I274915,I2690);
DFFARX1 I_16012 (I874436,I2683,I274915,I274941,);
nand I_16013 (I274949,I874451,I874436);
and I_16014 (I274966,I274949,I874454);
DFFARX1 I_16015 (I274966,I2683,I274915,I274992,);
nor I_16016 (I274883,I274992,I274941);
not I_16017 (I275014,I274992);
DFFARX1 I_16018 (I874460,I2683,I274915,I275040,);
nand I_16019 (I275048,I275040,I874442);
not I_16020 (I275065,I275048);
DFFARX1 I_16021 (I275065,I2683,I274915,I275091,);
not I_16022 (I274907,I275091);
nor I_16023 (I275113,I274941,I275048);
nor I_16024 (I274889,I274992,I275113);
DFFARX1 I_16025 (I874439,I2683,I274915,I275153,);
DFFARX1 I_16026 (I275153,I2683,I274915,I275170,);
not I_16027 (I275178,I275170);
not I_16028 (I275195,I275153);
nand I_16029 (I274892,I275195,I275014);
nand I_16030 (I275226,I874439,I874445);
and I_16031 (I275243,I275226,I874457);
DFFARX1 I_16032 (I275243,I2683,I274915,I275269,);
nor I_16033 (I275277,I275269,I274941);
DFFARX1 I_16034 (I275277,I2683,I274915,I274880,);
DFFARX1 I_16035 (I275269,I2683,I274915,I274898,);
nor I_16036 (I275322,I874448,I874445);
not I_16037 (I275339,I275322);
nor I_16038 (I274901,I275178,I275339);
nand I_16039 (I274886,I275195,I275339);
nor I_16040 (I274895,I274941,I275322);
DFFARX1 I_16041 (I275322,I2683,I274915,I274904,);
not I_16042 (I275442,I2690);
DFFARX1 I_16043 (I543390,I2683,I275442,I275468,);
nand I_16044 (I275476,I543381,I543396);
and I_16045 (I275493,I275476,I543402);
DFFARX1 I_16046 (I275493,I2683,I275442,I275519,);
nor I_16047 (I275410,I275519,I275468);
not I_16048 (I275541,I275519);
DFFARX1 I_16049 (I543387,I2683,I275442,I275567,);
nand I_16050 (I275575,I275567,I543381);
not I_16051 (I275592,I275575);
DFFARX1 I_16052 (I275592,I2683,I275442,I275618,);
not I_16053 (I275434,I275618);
nor I_16054 (I275640,I275468,I275575);
nor I_16055 (I275416,I275519,I275640);
DFFARX1 I_16056 (I543384,I2683,I275442,I275680,);
DFFARX1 I_16057 (I275680,I2683,I275442,I275697,);
not I_16058 (I275705,I275697);
not I_16059 (I275722,I275680);
nand I_16060 (I275419,I275722,I275541);
nand I_16061 (I275753,I543378,I543393);
and I_16062 (I275770,I275753,I543378);
DFFARX1 I_16063 (I275770,I2683,I275442,I275796,);
nor I_16064 (I275804,I275796,I275468);
DFFARX1 I_16065 (I275804,I2683,I275442,I275407,);
DFFARX1 I_16066 (I275796,I2683,I275442,I275425,);
nor I_16067 (I275849,I543399,I543393);
not I_16068 (I275866,I275849);
nor I_16069 (I275428,I275705,I275866);
nand I_16070 (I275413,I275722,I275866);
nor I_16071 (I275422,I275468,I275849);
DFFARX1 I_16072 (I275849,I2683,I275442,I275431,);
not I_16073 (I275969,I2690);
DFFARX1 I_16074 (I622788,I2683,I275969,I275995,);
nand I_16075 (I276003,I622791,I622785);
and I_16076 (I276020,I276003,I622797);
DFFARX1 I_16077 (I276020,I2683,I275969,I276046,);
nor I_16078 (I275937,I276046,I275995);
not I_16079 (I276068,I276046);
DFFARX1 I_16080 (I622800,I2683,I275969,I276094,);
nand I_16081 (I276102,I276094,I622791);
not I_16082 (I276119,I276102);
DFFARX1 I_16083 (I276119,I2683,I275969,I276145,);
not I_16084 (I275961,I276145);
nor I_16085 (I276167,I275995,I276102);
nor I_16086 (I275943,I276046,I276167);
DFFARX1 I_16087 (I622803,I2683,I275969,I276207,);
DFFARX1 I_16088 (I276207,I2683,I275969,I276224,);
not I_16089 (I276232,I276224);
not I_16090 (I276249,I276207);
nand I_16091 (I275946,I276249,I276068);
nand I_16092 (I276280,I622785,I622794);
and I_16093 (I276297,I276280,I622788);
DFFARX1 I_16094 (I276297,I2683,I275969,I276323,);
nor I_16095 (I276331,I276323,I275995);
DFFARX1 I_16096 (I276331,I2683,I275969,I275934,);
DFFARX1 I_16097 (I276323,I2683,I275969,I275952,);
nor I_16098 (I276376,I622806,I622794);
not I_16099 (I276393,I276376);
nor I_16100 (I275955,I276232,I276393);
nand I_16101 (I275940,I276249,I276393);
nor I_16102 (I275949,I275995,I276376);
DFFARX1 I_16103 (I276376,I2683,I275969,I275958,);
not I_16104 (I276496,I2690);
DFFARX1 I_16105 (I877904,I2683,I276496,I276522,);
nand I_16106 (I276530,I877919,I877904);
and I_16107 (I276547,I276530,I877922);
DFFARX1 I_16108 (I276547,I2683,I276496,I276573,);
nor I_16109 (I276464,I276573,I276522);
not I_16110 (I276595,I276573);
DFFARX1 I_16111 (I877928,I2683,I276496,I276621,);
nand I_16112 (I276629,I276621,I877910);
not I_16113 (I276646,I276629);
DFFARX1 I_16114 (I276646,I2683,I276496,I276672,);
not I_16115 (I276488,I276672);
nor I_16116 (I276694,I276522,I276629);
nor I_16117 (I276470,I276573,I276694);
DFFARX1 I_16118 (I877907,I2683,I276496,I276734,);
DFFARX1 I_16119 (I276734,I2683,I276496,I276751,);
not I_16120 (I276759,I276751);
not I_16121 (I276776,I276734);
nand I_16122 (I276473,I276776,I276595);
nand I_16123 (I276807,I877907,I877913);
and I_16124 (I276824,I276807,I877925);
DFFARX1 I_16125 (I276824,I2683,I276496,I276850,);
nor I_16126 (I276858,I276850,I276522);
DFFARX1 I_16127 (I276858,I2683,I276496,I276461,);
DFFARX1 I_16128 (I276850,I2683,I276496,I276479,);
nor I_16129 (I276903,I877916,I877913);
not I_16130 (I276920,I276903);
nor I_16131 (I276482,I276759,I276920);
nand I_16132 (I276467,I276776,I276920);
nor I_16133 (I276476,I276522,I276903);
DFFARX1 I_16134 (I276903,I2683,I276496,I276485,);
not I_16135 (I277023,I2690);
DFFARX1 I_16136 (I403845,I2683,I277023,I277049,);
nand I_16137 (I277057,I403845,I403857);
and I_16138 (I277074,I277057,I403842);
DFFARX1 I_16139 (I277074,I2683,I277023,I277100,);
nor I_16140 (I276991,I277100,I277049);
not I_16141 (I277122,I277100);
DFFARX1 I_16142 (I403866,I2683,I277023,I277148,);
nand I_16143 (I277156,I277148,I403863);
not I_16144 (I277173,I277156);
DFFARX1 I_16145 (I277173,I2683,I277023,I277199,);
not I_16146 (I277015,I277199);
nor I_16147 (I277221,I277049,I277156);
nor I_16148 (I276997,I277100,I277221);
DFFARX1 I_16149 (I403854,I2683,I277023,I277261,);
DFFARX1 I_16150 (I277261,I2683,I277023,I277278,);
not I_16151 (I277286,I277278);
not I_16152 (I277303,I277261);
nand I_16153 (I277000,I277303,I277122);
nand I_16154 (I277334,I403842,I403851);
and I_16155 (I277351,I277334,I403860);
DFFARX1 I_16156 (I277351,I2683,I277023,I277377,);
nor I_16157 (I277385,I277377,I277049);
DFFARX1 I_16158 (I277385,I2683,I277023,I276988,);
DFFARX1 I_16159 (I277377,I2683,I277023,I277006,);
nor I_16160 (I277430,I403848,I403851);
not I_16161 (I277447,I277430);
nor I_16162 (I277009,I277286,I277447);
nand I_16163 (I276994,I277303,I277447);
nor I_16164 (I277003,I277049,I277430);
DFFARX1 I_16165 (I277430,I2683,I277023,I277012,);
not I_16166 (I277550,I2690);
DFFARX1 I_16167 (I680231,I2683,I277550,I277576,);
nand I_16168 (I277584,I680234,I680228);
and I_16169 (I277601,I277584,I680240);
DFFARX1 I_16170 (I277601,I2683,I277550,I277627,);
nor I_16171 (I277518,I277627,I277576);
not I_16172 (I277649,I277627);
DFFARX1 I_16173 (I680243,I2683,I277550,I277675,);
nand I_16174 (I277683,I277675,I680234);
not I_16175 (I277700,I277683);
DFFARX1 I_16176 (I277700,I2683,I277550,I277726,);
not I_16177 (I277542,I277726);
nor I_16178 (I277748,I277576,I277683);
nor I_16179 (I277524,I277627,I277748);
DFFARX1 I_16180 (I680246,I2683,I277550,I277788,);
DFFARX1 I_16181 (I277788,I2683,I277550,I277805,);
not I_16182 (I277813,I277805);
not I_16183 (I277830,I277788);
nand I_16184 (I277527,I277830,I277649);
nand I_16185 (I277861,I680228,I680237);
and I_16186 (I277878,I277861,I680231);
DFFARX1 I_16187 (I277878,I2683,I277550,I277904,);
nor I_16188 (I277912,I277904,I277576);
DFFARX1 I_16189 (I277912,I2683,I277550,I277515,);
DFFARX1 I_16190 (I277904,I2683,I277550,I277533,);
nor I_16191 (I277957,I680249,I680237);
not I_16192 (I277974,I277957);
nor I_16193 (I277536,I277813,I277974);
nand I_16194 (I277521,I277830,I277974);
nor I_16195 (I277530,I277576,I277957);
DFFARX1 I_16196 (I277957,I2683,I277550,I277539,);
not I_16197 (I278077,I2690);
DFFARX1 I_16198 (I352990,I2683,I278077,I278103,);
nand I_16199 (I278111,I353002,I352981);
and I_16200 (I278128,I278111,I353005);
DFFARX1 I_16201 (I278128,I2683,I278077,I278154,);
nor I_16202 (I278045,I278154,I278103);
not I_16203 (I278176,I278154);
DFFARX1 I_16204 (I352996,I2683,I278077,I278202,);
nand I_16205 (I278210,I278202,I352978);
not I_16206 (I278227,I278210);
DFFARX1 I_16207 (I278227,I2683,I278077,I278253,);
not I_16208 (I278069,I278253);
nor I_16209 (I278275,I278103,I278210);
nor I_16210 (I278051,I278154,I278275);
DFFARX1 I_16211 (I352993,I2683,I278077,I278315,);
DFFARX1 I_16212 (I278315,I2683,I278077,I278332,);
not I_16213 (I278340,I278332);
not I_16214 (I278357,I278315);
nand I_16215 (I278054,I278357,I278176);
nand I_16216 (I278388,I352978,I352984);
and I_16217 (I278405,I278388,I352987);
DFFARX1 I_16218 (I278405,I2683,I278077,I278431,);
nor I_16219 (I278439,I278431,I278103);
DFFARX1 I_16220 (I278439,I2683,I278077,I278042,);
DFFARX1 I_16221 (I278431,I2683,I278077,I278060,);
nor I_16222 (I278484,I352999,I352984);
not I_16223 (I278501,I278484);
nor I_16224 (I278063,I278340,I278501);
nand I_16225 (I278048,I278357,I278501);
nor I_16226 (I278057,I278103,I278484);
DFFARX1 I_16227 (I278484,I2683,I278077,I278066,);
not I_16228 (I278604,I2690);
DFFARX1 I_16229 (I958128,I2683,I278604,I278630,);
nand I_16230 (I278638,I958110,I958134);
and I_16231 (I278655,I278638,I958125);
DFFARX1 I_16232 (I278655,I2683,I278604,I278681,);
nor I_16233 (I278572,I278681,I278630);
not I_16234 (I278703,I278681);
DFFARX1 I_16235 (I958131,I2683,I278604,I278729,);
nand I_16236 (I278737,I278729,I958119);
not I_16237 (I278754,I278737);
DFFARX1 I_16238 (I278754,I2683,I278604,I278780,);
not I_16239 (I278596,I278780);
nor I_16240 (I278802,I278630,I278737);
nor I_16241 (I278578,I278681,I278802);
DFFARX1 I_16242 (I958110,I2683,I278604,I278842,);
DFFARX1 I_16243 (I278842,I2683,I278604,I278859,);
not I_16244 (I278867,I278859);
not I_16245 (I278884,I278842);
nand I_16246 (I278581,I278884,I278703);
nand I_16247 (I278915,I958116,I958113);
and I_16248 (I278932,I278915,I958122);
DFFARX1 I_16249 (I278932,I2683,I278604,I278958,);
nor I_16250 (I278966,I278958,I278630);
DFFARX1 I_16251 (I278966,I2683,I278604,I278569,);
DFFARX1 I_16252 (I278958,I2683,I278604,I278587,);
nor I_16253 (I279011,I958113,I958113);
not I_16254 (I279028,I279011);
nor I_16255 (I278590,I278867,I279028);
nand I_16256 (I278575,I278884,I279028);
nor I_16257 (I278584,I278630,I279011);
DFFARX1 I_16258 (I279011,I2683,I278604,I278593,);
not I_16259 (I279131,I2690);
DFFARX1 I_16260 (I161065,I2683,I279131,I279157,);
nand I_16261 (I279165,I161065,I161071);
and I_16262 (I279182,I279165,I161089);
DFFARX1 I_16263 (I279182,I2683,I279131,I279208,);
nor I_16264 (I279099,I279208,I279157);
not I_16265 (I279230,I279208);
DFFARX1 I_16266 (I161077,I2683,I279131,I279256,);
nand I_16267 (I279264,I279256,I161074);
not I_16268 (I279281,I279264);
DFFARX1 I_16269 (I279281,I2683,I279131,I279307,);
not I_16270 (I279123,I279307);
nor I_16271 (I279329,I279157,I279264);
nor I_16272 (I279105,I279208,I279329);
DFFARX1 I_16273 (I161083,I2683,I279131,I279369,);
DFFARX1 I_16274 (I279369,I2683,I279131,I279386,);
not I_16275 (I279394,I279386);
not I_16276 (I279411,I279369);
nand I_16277 (I279108,I279411,I279230);
nand I_16278 (I279442,I161068,I161068);
and I_16279 (I279459,I279442,I161080);
DFFARX1 I_16280 (I279459,I2683,I279131,I279485,);
nor I_16281 (I279493,I279485,I279157);
DFFARX1 I_16282 (I279493,I2683,I279131,I279096,);
DFFARX1 I_16283 (I279485,I2683,I279131,I279114,);
nor I_16284 (I279538,I161086,I161068);
not I_16285 (I279555,I279538);
nor I_16286 (I279117,I279394,I279555);
nand I_16287 (I279102,I279411,I279555);
nor I_16288 (I279111,I279157,I279538);
DFFARX1 I_16289 (I279538,I2683,I279131,I279120,);
not I_16290 (I279658,I2690);
DFFARX1 I_16291 (I61159,I2683,I279658,I279684,);
nand I_16292 (I279692,I61171,I61180);
and I_16293 (I279709,I279692,I61159);
DFFARX1 I_16294 (I279709,I2683,I279658,I279735,);
nor I_16295 (I279626,I279735,I279684);
not I_16296 (I279757,I279735);
DFFARX1 I_16297 (I61174,I2683,I279658,I279783,);
nand I_16298 (I279791,I279783,I61162);
not I_16299 (I279808,I279791);
DFFARX1 I_16300 (I279808,I2683,I279658,I279834,);
not I_16301 (I279650,I279834);
nor I_16302 (I279856,I279684,I279791);
nor I_16303 (I279632,I279735,I279856);
DFFARX1 I_16304 (I61165,I2683,I279658,I279896,);
DFFARX1 I_16305 (I279896,I2683,I279658,I279913,);
not I_16306 (I279921,I279913);
not I_16307 (I279938,I279896);
nand I_16308 (I279635,I279938,I279757);
nand I_16309 (I279969,I61156,I61156);
and I_16310 (I279986,I279969,I61168);
DFFARX1 I_16311 (I279986,I2683,I279658,I280012,);
nor I_16312 (I280020,I280012,I279684);
DFFARX1 I_16313 (I280020,I2683,I279658,I279623,);
DFFARX1 I_16314 (I280012,I2683,I279658,I279641,);
nor I_16315 (I280065,I61177,I61156);
not I_16316 (I280082,I280065);
nor I_16317 (I279644,I279921,I280082);
nand I_16318 (I279629,I279938,I280082);
nor I_16319 (I279638,I279684,I280065);
DFFARX1 I_16320 (I280065,I2683,I279658,I279647,);
not I_16321 (I280185,I2690);
DFFARX1 I_16322 (I89090,I2683,I280185,I280211,);
nand I_16323 (I280219,I89102,I89111);
and I_16324 (I280236,I280219,I89090);
DFFARX1 I_16325 (I280236,I2683,I280185,I280262,);
nor I_16326 (I280153,I280262,I280211);
not I_16327 (I280284,I280262);
DFFARX1 I_16328 (I89105,I2683,I280185,I280310,);
nand I_16329 (I280318,I280310,I89093);
not I_16330 (I280335,I280318);
DFFARX1 I_16331 (I280335,I2683,I280185,I280361,);
not I_16332 (I280177,I280361);
nor I_16333 (I280383,I280211,I280318);
nor I_16334 (I280159,I280262,I280383);
DFFARX1 I_16335 (I89096,I2683,I280185,I280423,);
DFFARX1 I_16336 (I280423,I2683,I280185,I280440,);
not I_16337 (I280448,I280440);
not I_16338 (I280465,I280423);
nand I_16339 (I280162,I280465,I280284);
nand I_16340 (I280496,I89087,I89087);
and I_16341 (I280513,I280496,I89099);
DFFARX1 I_16342 (I280513,I2683,I280185,I280539,);
nor I_16343 (I280547,I280539,I280211);
DFFARX1 I_16344 (I280547,I2683,I280185,I280150,);
DFFARX1 I_16345 (I280539,I2683,I280185,I280168,);
nor I_16346 (I280592,I89108,I89087);
not I_16347 (I280609,I280592);
nor I_16348 (I280171,I280448,I280609);
nand I_16349 (I280156,I280465,I280609);
nor I_16350 (I280165,I280211,I280592);
DFFARX1 I_16351 (I280592,I2683,I280185,I280174,);
not I_16352 (I280712,I2690);
DFFARX1 I_16353 (I668637,I2683,I280712,I280738,);
nand I_16354 (I280746,I668640,I668634);
and I_16355 (I280763,I280746,I668646);
DFFARX1 I_16356 (I280763,I2683,I280712,I280789,);
nor I_16357 (I280680,I280789,I280738);
not I_16358 (I280811,I280789);
DFFARX1 I_16359 (I668649,I2683,I280712,I280837,);
nand I_16360 (I280845,I280837,I668640);
not I_16361 (I280862,I280845);
DFFARX1 I_16362 (I280862,I2683,I280712,I280888,);
not I_16363 (I280704,I280888);
nor I_16364 (I280910,I280738,I280845);
nor I_16365 (I280686,I280789,I280910);
DFFARX1 I_16366 (I668652,I2683,I280712,I280950,);
DFFARX1 I_16367 (I280950,I2683,I280712,I280967,);
not I_16368 (I280975,I280967);
not I_16369 (I280992,I280950);
nand I_16370 (I280689,I280992,I280811);
nand I_16371 (I281023,I668634,I668643);
and I_16372 (I281040,I281023,I668637);
DFFARX1 I_16373 (I281040,I2683,I280712,I281066,);
nor I_16374 (I281074,I281066,I280738);
DFFARX1 I_16375 (I281074,I2683,I280712,I280677,);
DFFARX1 I_16376 (I281066,I2683,I280712,I280695,);
nor I_16377 (I281119,I668655,I668643);
not I_16378 (I281136,I281119);
nor I_16379 (I280698,I280975,I281136);
nand I_16380 (I280683,I280992,I281136);
nor I_16381 (I280692,I280738,I281119);
DFFARX1 I_16382 (I281119,I2683,I280712,I280701,);
not I_16383 (I281239,I2690);
DFFARX1 I_16384 (I823150,I2683,I281239,I281265,);
nand I_16385 (I281273,I823147,I823150);
and I_16386 (I281290,I281273,I823159);
DFFARX1 I_16387 (I281290,I2683,I281239,I281316,);
nor I_16388 (I281207,I281316,I281265);
not I_16389 (I281338,I281316);
DFFARX1 I_16390 (I823147,I2683,I281239,I281364,);
nand I_16391 (I281372,I281364,I823165);
not I_16392 (I281389,I281372);
DFFARX1 I_16393 (I281389,I2683,I281239,I281415,);
not I_16394 (I281231,I281415);
nor I_16395 (I281437,I281265,I281372);
nor I_16396 (I281213,I281316,I281437);
DFFARX1 I_16397 (I823153,I2683,I281239,I281477,);
DFFARX1 I_16398 (I281477,I2683,I281239,I281494,);
not I_16399 (I281502,I281494);
not I_16400 (I281519,I281477);
nand I_16401 (I281216,I281519,I281338);
nand I_16402 (I281550,I823162,I823168);
and I_16403 (I281567,I281550,I823153);
DFFARX1 I_16404 (I281567,I2683,I281239,I281593,);
nor I_16405 (I281601,I281593,I281265);
DFFARX1 I_16406 (I281601,I2683,I281239,I281204,);
DFFARX1 I_16407 (I281593,I2683,I281239,I281222,);
nor I_16408 (I281646,I823156,I823168);
not I_16409 (I281663,I281646);
nor I_16410 (I281225,I281502,I281663);
nand I_16411 (I281210,I281519,I281663);
nor I_16412 (I281219,I281265,I281646);
DFFARX1 I_16413 (I281646,I2683,I281239,I281228,);
not I_16414 (I281766,I2690);
DFFARX1 I_16415 (I961936,I2683,I281766,I281792,);
nand I_16416 (I281800,I961918,I961942);
and I_16417 (I281817,I281800,I961933);
DFFARX1 I_16418 (I281817,I2683,I281766,I281843,);
nor I_16419 (I281734,I281843,I281792);
not I_16420 (I281865,I281843);
DFFARX1 I_16421 (I961939,I2683,I281766,I281891,);
nand I_16422 (I281899,I281891,I961927);
not I_16423 (I281916,I281899);
DFFARX1 I_16424 (I281916,I2683,I281766,I281942,);
not I_16425 (I281758,I281942);
nor I_16426 (I281964,I281792,I281899);
nor I_16427 (I281740,I281843,I281964);
DFFARX1 I_16428 (I961918,I2683,I281766,I282004,);
DFFARX1 I_16429 (I282004,I2683,I281766,I282021,);
not I_16430 (I282029,I282021);
not I_16431 (I282046,I282004);
nand I_16432 (I281743,I282046,I281865);
nand I_16433 (I282077,I961924,I961921);
and I_16434 (I282094,I282077,I961930);
DFFARX1 I_16435 (I282094,I2683,I281766,I282120,);
nor I_16436 (I282128,I282120,I281792);
DFFARX1 I_16437 (I282128,I2683,I281766,I281731,);
DFFARX1 I_16438 (I282120,I2683,I281766,I281749,);
nor I_16439 (I282173,I961921,I961921);
not I_16440 (I282190,I282173);
nor I_16441 (I281752,I282029,I282190);
nand I_16442 (I281737,I282046,I282190);
nor I_16443 (I281746,I281792,I282173);
DFFARX1 I_16444 (I282173,I2683,I281766,I281755,);
not I_16445 (I282293,I2690);
DFFARX1 I_16446 (I127150,I2683,I282293,I282319,);
nand I_16447 (I282327,I127150,I127156);
and I_16448 (I282344,I282327,I127174);
DFFARX1 I_16449 (I282344,I2683,I282293,I282370,);
nor I_16450 (I282261,I282370,I282319);
not I_16451 (I282392,I282370);
DFFARX1 I_16452 (I127162,I2683,I282293,I282418,);
nand I_16453 (I282426,I282418,I127159);
not I_16454 (I282443,I282426);
DFFARX1 I_16455 (I282443,I2683,I282293,I282469,);
not I_16456 (I282285,I282469);
nor I_16457 (I282491,I282319,I282426);
nor I_16458 (I282267,I282370,I282491);
DFFARX1 I_16459 (I127168,I2683,I282293,I282531,);
DFFARX1 I_16460 (I282531,I2683,I282293,I282548,);
not I_16461 (I282556,I282548);
not I_16462 (I282573,I282531);
nand I_16463 (I282270,I282573,I282392);
nand I_16464 (I282604,I127153,I127153);
and I_16465 (I282621,I282604,I127165);
DFFARX1 I_16466 (I282621,I2683,I282293,I282647,);
nor I_16467 (I282655,I282647,I282319);
DFFARX1 I_16468 (I282655,I2683,I282293,I282258,);
DFFARX1 I_16469 (I282647,I2683,I282293,I282276,);
nor I_16470 (I282700,I127171,I127153);
not I_16471 (I282717,I282700);
nor I_16472 (I282279,I282556,I282717);
nand I_16473 (I282264,I282573,I282717);
nor I_16474 (I282273,I282319,I282700);
DFFARX1 I_16475 (I282700,I2683,I282293,I282282,);
not I_16476 (I282820,I2690);
DFFARX1 I_16477 (I753586,I2683,I282820,I282846,);
nand I_16478 (I282854,I753583,I753601);
and I_16479 (I282871,I282854,I753592);
DFFARX1 I_16480 (I282871,I2683,I282820,I282897,);
nor I_16481 (I282788,I282897,I282846);
not I_16482 (I282919,I282897);
DFFARX1 I_16483 (I753607,I2683,I282820,I282945,);
nand I_16484 (I282953,I282945,I753589);
not I_16485 (I282970,I282953);
DFFARX1 I_16486 (I282970,I2683,I282820,I282996,);
not I_16487 (I282812,I282996);
nor I_16488 (I283018,I282846,I282953);
nor I_16489 (I282794,I282897,I283018);
DFFARX1 I_16490 (I753595,I2683,I282820,I283058,);
DFFARX1 I_16491 (I283058,I2683,I282820,I283075,);
not I_16492 (I283083,I283075);
not I_16493 (I283100,I283058);
nand I_16494 (I282797,I283100,I282919);
nand I_16495 (I283131,I753583,I753610);
and I_16496 (I283148,I283131,I753598);
DFFARX1 I_16497 (I283148,I2683,I282820,I283174,);
nor I_16498 (I283182,I283174,I282846);
DFFARX1 I_16499 (I283182,I2683,I282820,I282785,);
DFFARX1 I_16500 (I283174,I2683,I282820,I282803,);
nor I_16501 (I283227,I753604,I753610);
not I_16502 (I283244,I283227);
nor I_16503 (I282806,I283083,I283244);
nand I_16504 (I282791,I283100,I283244);
nor I_16505 (I282800,I282846,I283227);
DFFARX1 I_16506 (I283227,I2683,I282820,I282809,);
not I_16507 (I283347,I2690);
DFFARX1 I_16508 (I824272,I2683,I283347,I283373,);
nand I_16509 (I283381,I824269,I824272);
and I_16510 (I283398,I283381,I824281);
DFFARX1 I_16511 (I283398,I2683,I283347,I283424,);
nor I_16512 (I283315,I283424,I283373);
not I_16513 (I283446,I283424);
DFFARX1 I_16514 (I824269,I2683,I283347,I283472,);
nand I_16515 (I283480,I283472,I824287);
not I_16516 (I283497,I283480);
DFFARX1 I_16517 (I283497,I2683,I283347,I283523,);
not I_16518 (I283339,I283523);
nor I_16519 (I283545,I283373,I283480);
nor I_16520 (I283321,I283424,I283545);
DFFARX1 I_16521 (I824275,I2683,I283347,I283585,);
DFFARX1 I_16522 (I283585,I2683,I283347,I283602,);
not I_16523 (I283610,I283602);
not I_16524 (I283627,I283585);
nand I_16525 (I283324,I283627,I283446);
nand I_16526 (I283658,I824284,I824290);
and I_16527 (I283675,I283658,I824275);
DFFARX1 I_16528 (I283675,I2683,I283347,I283701,);
nor I_16529 (I283709,I283701,I283373);
DFFARX1 I_16530 (I283709,I2683,I283347,I283312,);
DFFARX1 I_16531 (I283701,I2683,I283347,I283330,);
nor I_16532 (I283754,I824278,I824290);
not I_16533 (I283771,I283754);
nor I_16534 (I283333,I283610,I283771);
nand I_16535 (I283318,I283627,I283771);
nor I_16536 (I283327,I283373,I283754);
DFFARX1 I_16537 (I283754,I2683,I283347,I283336,);
not I_16538 (I283874,I2690);
DFFARX1 I_16539 (I1013443,I2683,I283874,I283900,);
nand I_16540 (I283908,I1013440,I1013431);
and I_16541 (I283925,I283908,I1013428);
DFFARX1 I_16542 (I283925,I2683,I283874,I283951,);
nor I_16543 (I283842,I283951,I283900);
not I_16544 (I283973,I283951);
DFFARX1 I_16545 (I1013437,I2683,I283874,I283999,);
nand I_16546 (I284007,I283999,I1013446);
not I_16547 (I284024,I284007);
DFFARX1 I_16548 (I284024,I2683,I283874,I284050,);
not I_16549 (I283866,I284050);
nor I_16550 (I284072,I283900,I284007);
nor I_16551 (I283848,I283951,I284072);
DFFARX1 I_16552 (I1013449,I2683,I283874,I284112,);
DFFARX1 I_16553 (I284112,I2683,I283874,I284129,);
not I_16554 (I284137,I284129);
not I_16555 (I284154,I284112);
nand I_16556 (I283851,I284154,I283973);
nand I_16557 (I284185,I1013428,I1013434);
and I_16558 (I284202,I284185,I1013452);
DFFARX1 I_16559 (I284202,I2683,I283874,I284228,);
nor I_16560 (I284236,I284228,I283900);
DFFARX1 I_16561 (I284236,I2683,I283874,I283839,);
DFFARX1 I_16562 (I284228,I2683,I283874,I283857,);
nor I_16563 (I284281,I1013431,I1013434);
not I_16564 (I284298,I284281);
nor I_16565 (I283860,I284137,I284298);
nand I_16566 (I283845,I284154,I284298);
nor I_16567 (I283854,I283900,I284281);
DFFARX1 I_16568 (I284281,I2683,I283874,I283863,);
not I_16569 (I284401,I2690);
DFFARX1 I_16570 (I575180,I2683,I284401,I284427,);
nand I_16571 (I284435,I575171,I575186);
and I_16572 (I284452,I284435,I575192);
DFFARX1 I_16573 (I284452,I2683,I284401,I284478,);
nor I_16574 (I284369,I284478,I284427);
not I_16575 (I284500,I284478);
DFFARX1 I_16576 (I575177,I2683,I284401,I284526,);
nand I_16577 (I284534,I284526,I575171);
not I_16578 (I284551,I284534);
DFFARX1 I_16579 (I284551,I2683,I284401,I284577,);
not I_16580 (I284393,I284577);
nor I_16581 (I284599,I284427,I284534);
nor I_16582 (I284375,I284478,I284599);
DFFARX1 I_16583 (I575174,I2683,I284401,I284639,);
DFFARX1 I_16584 (I284639,I2683,I284401,I284656,);
not I_16585 (I284664,I284656);
not I_16586 (I284681,I284639);
nand I_16587 (I284378,I284681,I284500);
nand I_16588 (I284712,I575168,I575183);
and I_16589 (I284729,I284712,I575168);
DFFARX1 I_16590 (I284729,I2683,I284401,I284755,);
nor I_16591 (I284763,I284755,I284427);
DFFARX1 I_16592 (I284763,I2683,I284401,I284366,);
DFFARX1 I_16593 (I284755,I2683,I284401,I284384,);
nor I_16594 (I284808,I575189,I575183);
not I_16595 (I284825,I284808);
nor I_16596 (I284387,I284664,I284825);
nand I_16597 (I284372,I284681,I284825);
nor I_16598 (I284381,I284427,I284808);
DFFARX1 I_16599 (I284808,I2683,I284401,I284390,);
not I_16600 (I284928,I2690);
DFFARX1 I_16601 (I167610,I2683,I284928,I284954,);
nand I_16602 (I284962,I167610,I167616);
and I_16603 (I284979,I284962,I167634);
DFFARX1 I_16604 (I284979,I2683,I284928,I285005,);
nor I_16605 (I284896,I285005,I284954);
not I_16606 (I285027,I285005);
DFFARX1 I_16607 (I167622,I2683,I284928,I285053,);
nand I_16608 (I285061,I285053,I167619);
not I_16609 (I285078,I285061);
DFFARX1 I_16610 (I285078,I2683,I284928,I285104,);
not I_16611 (I284920,I285104);
nor I_16612 (I285126,I284954,I285061);
nor I_16613 (I284902,I285005,I285126);
DFFARX1 I_16614 (I167628,I2683,I284928,I285166,);
DFFARX1 I_16615 (I285166,I2683,I284928,I285183,);
not I_16616 (I285191,I285183);
not I_16617 (I285208,I285166);
nand I_16618 (I284905,I285208,I285027);
nand I_16619 (I285239,I167613,I167613);
and I_16620 (I285256,I285239,I167625);
DFFARX1 I_16621 (I285256,I2683,I284928,I285282,);
nor I_16622 (I285290,I285282,I284954);
DFFARX1 I_16623 (I285290,I2683,I284928,I284893,);
DFFARX1 I_16624 (I285282,I2683,I284928,I284911,);
nor I_16625 (I285335,I167631,I167613);
not I_16626 (I285352,I285335);
nor I_16627 (I284914,I285191,I285352);
nand I_16628 (I284899,I285208,I285352);
nor I_16629 (I284908,I284954,I285335);
DFFARX1 I_16630 (I285335,I2683,I284928,I284917,);
not I_16631 (I285455,I2690);
DFFARX1 I_16632 (I831086,I2683,I285455,I285481,);
nand I_16633 (I285489,I831101,I831086);
and I_16634 (I285506,I285489,I831104);
DFFARX1 I_16635 (I285506,I2683,I285455,I285532,);
nor I_16636 (I285423,I285532,I285481);
not I_16637 (I285554,I285532);
DFFARX1 I_16638 (I831110,I2683,I285455,I285580,);
nand I_16639 (I285588,I285580,I831092);
not I_16640 (I285605,I285588);
DFFARX1 I_16641 (I285605,I2683,I285455,I285631,);
not I_16642 (I285447,I285631);
nor I_16643 (I285653,I285481,I285588);
nor I_16644 (I285429,I285532,I285653);
DFFARX1 I_16645 (I831089,I2683,I285455,I285693,);
DFFARX1 I_16646 (I285693,I2683,I285455,I285710,);
not I_16647 (I285718,I285710);
not I_16648 (I285735,I285693);
nand I_16649 (I285432,I285735,I285554);
nand I_16650 (I285766,I831089,I831095);
and I_16651 (I285783,I285766,I831107);
DFFARX1 I_16652 (I285783,I2683,I285455,I285809,);
nor I_16653 (I285817,I285809,I285481);
DFFARX1 I_16654 (I285817,I2683,I285455,I285420,);
DFFARX1 I_16655 (I285809,I2683,I285455,I285438,);
nor I_16656 (I285862,I831098,I831095);
not I_16657 (I285879,I285862);
nor I_16658 (I285441,I285718,I285879);
nand I_16659 (I285426,I285735,I285879);
nor I_16660 (I285435,I285481,I285862);
DFFARX1 I_16661 (I285862,I2683,I285455,I285444,);
not I_16662 (I285982,I2690);
DFFARX1 I_16663 (I56416,I2683,I285982,I286008,);
nand I_16664 (I286016,I56428,I56437);
and I_16665 (I286033,I286016,I56416);
DFFARX1 I_16666 (I286033,I2683,I285982,I286059,);
nor I_16667 (I285950,I286059,I286008);
not I_16668 (I286081,I286059);
DFFARX1 I_16669 (I56431,I2683,I285982,I286107,);
nand I_16670 (I286115,I286107,I56419);
not I_16671 (I286132,I286115);
DFFARX1 I_16672 (I286132,I2683,I285982,I286158,);
not I_16673 (I285974,I286158);
nor I_16674 (I286180,I286008,I286115);
nor I_16675 (I285956,I286059,I286180);
DFFARX1 I_16676 (I56422,I2683,I285982,I286220,);
DFFARX1 I_16677 (I286220,I2683,I285982,I286237,);
not I_16678 (I286245,I286237);
not I_16679 (I286262,I286220);
nand I_16680 (I285959,I286262,I286081);
nand I_16681 (I286293,I56413,I56413);
and I_16682 (I286310,I286293,I56425);
DFFARX1 I_16683 (I286310,I2683,I285982,I286336,);
nor I_16684 (I286344,I286336,I286008);
DFFARX1 I_16685 (I286344,I2683,I285982,I285947,);
DFFARX1 I_16686 (I286336,I2683,I285982,I285965,);
nor I_16687 (I286389,I56434,I56413);
not I_16688 (I286406,I286389);
nor I_16689 (I285968,I286245,I286406);
nand I_16690 (I285953,I286262,I286406);
nor I_16691 (I285962,I286008,I286389);
DFFARX1 I_16692 (I286389,I2683,I285982,I285971,);
not I_16693 (I286509,I2690);
DFFARX1 I_16694 (I713534,I2683,I286509,I286535,);
nand I_16695 (I286543,I713531,I713549);
and I_16696 (I286560,I286543,I713540);
DFFARX1 I_16697 (I286560,I2683,I286509,I286586,);
nor I_16698 (I286477,I286586,I286535);
not I_16699 (I286608,I286586);
DFFARX1 I_16700 (I713555,I2683,I286509,I286634,);
nand I_16701 (I286642,I286634,I713537);
not I_16702 (I286659,I286642);
DFFARX1 I_16703 (I286659,I2683,I286509,I286685,);
not I_16704 (I286501,I286685);
nor I_16705 (I286707,I286535,I286642);
nor I_16706 (I286483,I286586,I286707);
DFFARX1 I_16707 (I713543,I2683,I286509,I286747,);
DFFARX1 I_16708 (I286747,I2683,I286509,I286764,);
not I_16709 (I286772,I286764);
not I_16710 (I286789,I286747);
nand I_16711 (I286486,I286789,I286608);
nand I_16712 (I286820,I713531,I713558);
and I_16713 (I286837,I286820,I713546);
DFFARX1 I_16714 (I286837,I2683,I286509,I286863,);
nor I_16715 (I286871,I286863,I286535);
DFFARX1 I_16716 (I286871,I2683,I286509,I286474,);
DFFARX1 I_16717 (I286863,I2683,I286509,I286492,);
nor I_16718 (I286916,I713552,I713558);
not I_16719 (I286933,I286916);
nor I_16720 (I286495,I286772,I286933);
nand I_16721 (I286480,I286789,I286933);
nor I_16722 (I286489,I286535,I286916);
DFFARX1 I_16723 (I286916,I2683,I286509,I286498,);
not I_16724 (I287036,I2690);
DFFARX1 I_16725 (I679177,I2683,I287036,I287062,);
nand I_16726 (I287070,I679180,I679174);
and I_16727 (I287087,I287070,I679186);
DFFARX1 I_16728 (I287087,I2683,I287036,I287113,);
nor I_16729 (I287004,I287113,I287062);
not I_16730 (I287135,I287113);
DFFARX1 I_16731 (I679189,I2683,I287036,I287161,);
nand I_16732 (I287169,I287161,I679180);
not I_16733 (I287186,I287169);
DFFARX1 I_16734 (I287186,I2683,I287036,I287212,);
not I_16735 (I287028,I287212);
nor I_16736 (I287234,I287062,I287169);
nor I_16737 (I287010,I287113,I287234);
DFFARX1 I_16738 (I679192,I2683,I287036,I287274,);
DFFARX1 I_16739 (I287274,I2683,I287036,I287291,);
not I_16740 (I287299,I287291);
not I_16741 (I287316,I287274);
nand I_16742 (I287013,I287316,I287135);
nand I_16743 (I287347,I679174,I679183);
and I_16744 (I287364,I287347,I679177);
DFFARX1 I_16745 (I287364,I2683,I287036,I287390,);
nor I_16746 (I287398,I287390,I287062);
DFFARX1 I_16747 (I287398,I2683,I287036,I287001,);
DFFARX1 I_16748 (I287390,I2683,I287036,I287019,);
nor I_16749 (I287443,I679195,I679183);
not I_16750 (I287460,I287443);
nor I_16751 (I287022,I287299,I287460);
nand I_16752 (I287007,I287316,I287460);
nor I_16753 (I287016,I287062,I287443);
DFFARX1 I_16754 (I287443,I2683,I287036,I287025,);
not I_16755 (I287563,I2690);
DFFARX1 I_16756 (I110170,I2683,I287563,I287589,);
nand I_16757 (I287597,I110182,I110191);
and I_16758 (I287614,I287597,I110170);
DFFARX1 I_16759 (I287614,I2683,I287563,I287640,);
nor I_16760 (I287531,I287640,I287589);
not I_16761 (I287662,I287640);
DFFARX1 I_16762 (I110185,I2683,I287563,I287688,);
nand I_16763 (I287696,I287688,I110173);
not I_16764 (I287713,I287696);
DFFARX1 I_16765 (I287713,I2683,I287563,I287739,);
not I_16766 (I287555,I287739);
nor I_16767 (I287761,I287589,I287696);
nor I_16768 (I287537,I287640,I287761);
DFFARX1 I_16769 (I110176,I2683,I287563,I287801,);
DFFARX1 I_16770 (I287801,I2683,I287563,I287818,);
not I_16771 (I287826,I287818);
not I_16772 (I287843,I287801);
nand I_16773 (I287540,I287843,I287662);
nand I_16774 (I287874,I110167,I110167);
and I_16775 (I287891,I287874,I110179);
DFFARX1 I_16776 (I287891,I2683,I287563,I287917,);
nor I_16777 (I287925,I287917,I287589);
DFFARX1 I_16778 (I287925,I2683,I287563,I287528,);
DFFARX1 I_16779 (I287917,I2683,I287563,I287546,);
nor I_16780 (I287970,I110188,I110167);
not I_16781 (I287987,I287970);
nor I_16782 (I287549,I287826,I287987);
nand I_16783 (I287534,I287843,I287987);
nor I_16784 (I287543,I287589,I287970);
DFFARX1 I_16785 (I287970,I2683,I287563,I287552,);
not I_16786 (I288090,I2690);
DFFARX1 I_16787 (I861720,I2683,I288090,I288116,);
nand I_16788 (I288124,I861735,I861720);
and I_16789 (I288141,I288124,I861738);
DFFARX1 I_16790 (I288141,I2683,I288090,I288167,);
nor I_16791 (I288058,I288167,I288116);
not I_16792 (I288189,I288167);
DFFARX1 I_16793 (I861744,I2683,I288090,I288215,);
nand I_16794 (I288223,I288215,I861726);
not I_16795 (I288240,I288223);
DFFARX1 I_16796 (I288240,I2683,I288090,I288266,);
not I_16797 (I288082,I288266);
nor I_16798 (I288288,I288116,I288223);
nor I_16799 (I288064,I288167,I288288);
DFFARX1 I_16800 (I861723,I2683,I288090,I288328,);
DFFARX1 I_16801 (I288328,I2683,I288090,I288345,);
not I_16802 (I288353,I288345);
not I_16803 (I288370,I288328);
nand I_16804 (I288067,I288370,I288189);
nand I_16805 (I288401,I861723,I861729);
and I_16806 (I288418,I288401,I861741);
DFFARX1 I_16807 (I288418,I2683,I288090,I288444,);
nor I_16808 (I288452,I288444,I288116);
DFFARX1 I_16809 (I288452,I2683,I288090,I288055,);
DFFARX1 I_16810 (I288444,I2683,I288090,I288073,);
nor I_16811 (I288497,I861732,I861729);
not I_16812 (I288514,I288497);
nor I_16813 (I288076,I288353,I288514);
nand I_16814 (I288061,I288370,I288514);
nor I_16815 (I288070,I288116,I288497);
DFFARX1 I_16816 (I288497,I2683,I288090,I288079,);
not I_16817 (I288617,I2690);
DFFARX1 I_16818 (I899868,I2683,I288617,I288643,);
nand I_16819 (I288651,I899883,I899868);
and I_16820 (I288668,I288651,I899886);
DFFARX1 I_16821 (I288668,I2683,I288617,I288694,);
nor I_16822 (I288585,I288694,I288643);
not I_16823 (I288716,I288694);
DFFARX1 I_16824 (I899892,I2683,I288617,I288742,);
nand I_16825 (I288750,I288742,I899874);
not I_16826 (I288767,I288750);
DFFARX1 I_16827 (I288767,I2683,I288617,I288793,);
not I_16828 (I288609,I288793);
nor I_16829 (I288815,I288643,I288750);
nor I_16830 (I288591,I288694,I288815);
DFFARX1 I_16831 (I899871,I2683,I288617,I288855,);
DFFARX1 I_16832 (I288855,I2683,I288617,I288872,);
not I_16833 (I288880,I288872);
not I_16834 (I288897,I288855);
nand I_16835 (I288594,I288897,I288716);
nand I_16836 (I288928,I899871,I899877);
and I_16837 (I288945,I288928,I899889);
DFFARX1 I_16838 (I288945,I2683,I288617,I288971,);
nor I_16839 (I288979,I288971,I288643);
DFFARX1 I_16840 (I288979,I2683,I288617,I288582,);
DFFARX1 I_16841 (I288971,I2683,I288617,I288600,);
nor I_16842 (I289024,I899880,I899877);
not I_16843 (I289041,I289024);
nor I_16844 (I288603,I288880,I289041);
nand I_16845 (I288588,I288897,I289041);
nor I_16846 (I288597,I288643,I289024);
DFFARX1 I_16847 (I289024,I2683,I288617,I288606,);
not I_16848 (I289144,I2690);
DFFARX1 I_16849 (I851894,I2683,I289144,I289170,);
nand I_16850 (I289178,I851909,I851894);
and I_16851 (I289195,I289178,I851912);
DFFARX1 I_16852 (I289195,I2683,I289144,I289221,);
nor I_16853 (I289112,I289221,I289170);
not I_16854 (I289243,I289221);
DFFARX1 I_16855 (I851918,I2683,I289144,I289269,);
nand I_16856 (I289277,I289269,I851900);
not I_16857 (I289294,I289277);
DFFARX1 I_16858 (I289294,I2683,I289144,I289320,);
not I_16859 (I289136,I289320);
nor I_16860 (I289342,I289170,I289277);
nor I_16861 (I289118,I289221,I289342);
DFFARX1 I_16862 (I851897,I2683,I289144,I289382,);
DFFARX1 I_16863 (I289382,I2683,I289144,I289399,);
not I_16864 (I289407,I289399);
not I_16865 (I289424,I289382);
nand I_16866 (I289121,I289424,I289243);
nand I_16867 (I289455,I851897,I851903);
and I_16868 (I289472,I289455,I851915);
DFFARX1 I_16869 (I289472,I2683,I289144,I289498,);
nor I_16870 (I289506,I289498,I289170);
DFFARX1 I_16871 (I289506,I2683,I289144,I289109,);
DFFARX1 I_16872 (I289498,I2683,I289144,I289127,);
nor I_16873 (I289551,I851906,I851903);
not I_16874 (I289568,I289551);
nor I_16875 (I289130,I289407,I289568);
nand I_16876 (I289115,I289424,I289568);
nor I_16877 (I289124,I289170,I289551);
DFFARX1 I_16878 (I289551,I2683,I289144,I289133,);
not I_16879 (I289671,I2690);
DFFARX1 I_16880 (I955356,I2683,I289671,I289697,);
nand I_16881 (I289705,I955371,I955356);
and I_16882 (I289722,I289705,I955374);
DFFARX1 I_16883 (I289722,I2683,I289671,I289748,);
nor I_16884 (I289639,I289748,I289697);
not I_16885 (I289770,I289748);
DFFARX1 I_16886 (I955380,I2683,I289671,I289796,);
nand I_16887 (I289804,I289796,I955362);
not I_16888 (I289821,I289804);
DFFARX1 I_16889 (I289821,I2683,I289671,I289847,);
not I_16890 (I289663,I289847);
nor I_16891 (I289869,I289697,I289804);
nor I_16892 (I289645,I289748,I289869);
DFFARX1 I_16893 (I955359,I2683,I289671,I289909,);
DFFARX1 I_16894 (I289909,I2683,I289671,I289926,);
not I_16895 (I289934,I289926);
not I_16896 (I289951,I289909);
nand I_16897 (I289648,I289951,I289770);
nand I_16898 (I289982,I955359,I955365);
and I_16899 (I289999,I289982,I955377);
DFFARX1 I_16900 (I289999,I2683,I289671,I290025,);
nor I_16901 (I290033,I290025,I289697);
DFFARX1 I_16902 (I290033,I2683,I289671,I289636,);
DFFARX1 I_16903 (I290025,I2683,I289671,I289654,);
nor I_16904 (I290078,I955368,I955365);
not I_16905 (I290095,I290078);
nor I_16906 (I289657,I289934,I290095);
nand I_16907 (I289642,I289951,I290095);
nor I_16908 (I289651,I289697,I290078);
DFFARX1 I_16909 (I290078,I2683,I289671,I289660,);
not I_16910 (I290198,I2690);
DFFARX1 I_16911 (I456693,I2683,I290198,I290224,);
nand I_16912 (I290232,I456678,I456681);
and I_16913 (I290249,I290232,I456696);
DFFARX1 I_16914 (I290249,I2683,I290198,I290275,);
nor I_16915 (I290166,I290275,I290224);
not I_16916 (I290297,I290275);
DFFARX1 I_16917 (I456690,I2683,I290198,I290323,);
nand I_16918 (I290331,I290323,I456681);
not I_16919 (I290348,I290331);
DFFARX1 I_16920 (I290348,I2683,I290198,I290374,);
not I_16921 (I290190,I290374);
nor I_16922 (I290396,I290224,I290331);
nor I_16923 (I290172,I290275,I290396);
DFFARX1 I_16924 (I456687,I2683,I290198,I290436,);
DFFARX1 I_16925 (I290436,I2683,I290198,I290453,);
not I_16926 (I290461,I290453);
not I_16927 (I290478,I290436);
nand I_16928 (I290175,I290478,I290297);
nand I_16929 (I290509,I456702,I456678);
and I_16930 (I290526,I290509,I456699);
DFFARX1 I_16931 (I290526,I2683,I290198,I290552,);
nor I_16932 (I290560,I290552,I290224);
DFFARX1 I_16933 (I290560,I2683,I290198,I290163,);
DFFARX1 I_16934 (I290552,I2683,I290198,I290181,);
nor I_16935 (I290605,I456684,I456678);
not I_16936 (I290622,I290605);
nor I_16937 (I290184,I290461,I290622);
nand I_16938 (I290169,I290478,I290622);
nor I_16939 (I290178,I290224,I290605);
DFFARX1 I_16940 (I290605,I2683,I290198,I290187,);
not I_16941 (I290725,I2690);
DFFARX1 I_16942 (I137860,I2683,I290725,I290751,);
nand I_16943 (I290759,I137860,I137866);
and I_16944 (I290776,I290759,I137884);
DFFARX1 I_16945 (I290776,I2683,I290725,I290802,);
nor I_16946 (I290693,I290802,I290751);
not I_16947 (I290824,I290802);
DFFARX1 I_16948 (I137872,I2683,I290725,I290850,);
nand I_16949 (I290858,I290850,I137869);
not I_16950 (I290875,I290858);
DFFARX1 I_16951 (I290875,I2683,I290725,I290901,);
not I_16952 (I290717,I290901);
nor I_16953 (I290923,I290751,I290858);
nor I_16954 (I290699,I290802,I290923);
DFFARX1 I_16955 (I137878,I2683,I290725,I290963,);
DFFARX1 I_16956 (I290963,I2683,I290725,I290980,);
not I_16957 (I290988,I290980);
not I_16958 (I291005,I290963);
nand I_16959 (I290702,I291005,I290824);
nand I_16960 (I291036,I137863,I137863);
and I_16961 (I291053,I291036,I137875);
DFFARX1 I_16962 (I291053,I2683,I290725,I291079,);
nor I_16963 (I291087,I291079,I290751);
DFFARX1 I_16964 (I291087,I2683,I290725,I290690,);
DFFARX1 I_16965 (I291079,I2683,I290725,I290708,);
nor I_16966 (I291132,I137881,I137863);
not I_16967 (I291149,I291132);
nor I_16968 (I290711,I290988,I291149);
nand I_16969 (I290696,I291005,I291149);
nor I_16970 (I290705,I290751,I291132);
DFFARX1 I_16971 (I291132,I2683,I290725,I290714,);
not I_16972 (I291252,I2690);
DFFARX1 I_16973 (I205690,I2683,I291252,I291278,);
nand I_16974 (I291286,I205690,I205696);
and I_16975 (I291303,I291286,I205714);
DFFARX1 I_16976 (I291303,I2683,I291252,I291329,);
nor I_16977 (I291220,I291329,I291278);
not I_16978 (I291351,I291329);
DFFARX1 I_16979 (I205702,I2683,I291252,I291377,);
nand I_16980 (I291385,I291377,I205699);
not I_16981 (I291402,I291385);
DFFARX1 I_16982 (I291402,I2683,I291252,I291428,);
not I_16983 (I291244,I291428);
nor I_16984 (I291450,I291278,I291385);
nor I_16985 (I291226,I291329,I291450);
DFFARX1 I_16986 (I205708,I2683,I291252,I291490,);
DFFARX1 I_16987 (I291490,I2683,I291252,I291507,);
not I_16988 (I291515,I291507);
not I_16989 (I291532,I291490);
nand I_16990 (I291229,I291532,I291351);
nand I_16991 (I291563,I205693,I205693);
and I_16992 (I291580,I291563,I205705);
DFFARX1 I_16993 (I291580,I2683,I291252,I291606,);
nor I_16994 (I291614,I291606,I291278);
DFFARX1 I_16995 (I291614,I2683,I291252,I291217,);
DFFARX1 I_16996 (I291606,I2683,I291252,I291235,);
nor I_16997 (I291659,I205711,I205693);
not I_16998 (I291676,I291659);
nor I_16999 (I291238,I291515,I291676);
nand I_17000 (I291223,I291532,I291676);
nor I_17001 (I291232,I291278,I291659);
DFFARX1 I_17002 (I291659,I2683,I291252,I291241,);
not I_17003 (I291779,I2690);
DFFARX1 I_17004 (I914896,I2683,I291779,I291805,);
nand I_17005 (I291813,I914911,I914896);
and I_17006 (I291830,I291813,I914914);
DFFARX1 I_17007 (I291830,I2683,I291779,I291856,);
nor I_17008 (I291747,I291856,I291805);
not I_17009 (I291878,I291856);
DFFARX1 I_17010 (I914920,I2683,I291779,I291904,);
nand I_17011 (I291912,I291904,I914902);
not I_17012 (I291929,I291912);
DFFARX1 I_17013 (I291929,I2683,I291779,I291955,);
not I_17014 (I291771,I291955);
nor I_17015 (I291977,I291805,I291912);
nor I_17016 (I291753,I291856,I291977);
DFFARX1 I_17017 (I914899,I2683,I291779,I292017,);
DFFARX1 I_17018 (I292017,I2683,I291779,I292034,);
not I_17019 (I292042,I292034);
not I_17020 (I292059,I292017);
nand I_17021 (I291756,I292059,I291878);
nand I_17022 (I292090,I914899,I914905);
and I_17023 (I292107,I292090,I914917);
DFFARX1 I_17024 (I292107,I2683,I291779,I292133,);
nor I_17025 (I292141,I292133,I291805);
DFFARX1 I_17026 (I292141,I2683,I291779,I291744,);
DFFARX1 I_17027 (I292133,I2683,I291779,I291762,);
nor I_17028 (I292186,I914908,I914905);
not I_17029 (I292203,I292186);
nor I_17030 (I291765,I292042,I292203);
nand I_17031 (I291750,I292059,I292203);
nor I_17032 (I291759,I291805,I292186);
DFFARX1 I_17033 (I292186,I2683,I291779,I291768,);
not I_17034 (I292306,I2690);
DFFARX1 I_17035 (I410985,I2683,I292306,I292332,);
nand I_17036 (I292340,I410985,I410997);
and I_17037 (I292357,I292340,I410982);
DFFARX1 I_17038 (I292357,I2683,I292306,I292383,);
nor I_17039 (I292274,I292383,I292332);
not I_17040 (I292405,I292383);
DFFARX1 I_17041 (I411006,I2683,I292306,I292431,);
nand I_17042 (I292439,I292431,I411003);
not I_17043 (I292456,I292439);
DFFARX1 I_17044 (I292456,I2683,I292306,I292482,);
not I_17045 (I292298,I292482);
nor I_17046 (I292504,I292332,I292439);
nor I_17047 (I292280,I292383,I292504);
DFFARX1 I_17048 (I410994,I2683,I292306,I292544,);
DFFARX1 I_17049 (I292544,I2683,I292306,I292561,);
not I_17050 (I292569,I292561);
not I_17051 (I292586,I292544);
nand I_17052 (I292283,I292586,I292405);
nand I_17053 (I292617,I410982,I410991);
and I_17054 (I292634,I292617,I411000);
DFFARX1 I_17055 (I292634,I2683,I292306,I292660,);
nor I_17056 (I292668,I292660,I292332);
DFFARX1 I_17057 (I292668,I2683,I292306,I292271,);
DFFARX1 I_17058 (I292660,I2683,I292306,I292289,);
nor I_17059 (I292713,I410988,I410991);
not I_17060 (I292730,I292713);
nor I_17061 (I292292,I292569,I292730);
nand I_17062 (I292277,I292586,I292730);
nor I_17063 (I292286,I292332,I292713);
DFFARX1 I_17064 (I292713,I2683,I292306,I292295,);
not I_17065 (I292833,I2690);
DFFARX1 I_17066 (I88036,I2683,I292833,I292859,);
nand I_17067 (I292867,I88048,I88057);
and I_17068 (I292884,I292867,I88036);
DFFARX1 I_17069 (I292884,I2683,I292833,I292910,);
nor I_17070 (I292801,I292910,I292859);
not I_17071 (I292932,I292910);
DFFARX1 I_17072 (I88051,I2683,I292833,I292958,);
nand I_17073 (I292966,I292958,I88039);
not I_17074 (I292983,I292966);
DFFARX1 I_17075 (I292983,I2683,I292833,I293009,);
not I_17076 (I292825,I293009);
nor I_17077 (I293031,I292859,I292966);
nor I_17078 (I292807,I292910,I293031);
DFFARX1 I_17079 (I88042,I2683,I292833,I293071,);
DFFARX1 I_17080 (I293071,I2683,I292833,I293088,);
not I_17081 (I293096,I293088);
not I_17082 (I293113,I293071);
nand I_17083 (I292810,I293113,I292932);
nand I_17084 (I293144,I88033,I88033);
and I_17085 (I293161,I293144,I88045);
DFFARX1 I_17086 (I293161,I2683,I292833,I293187,);
nor I_17087 (I293195,I293187,I292859);
DFFARX1 I_17088 (I293195,I2683,I292833,I292798,);
DFFARX1 I_17089 (I293187,I2683,I292833,I292816,);
nor I_17090 (I293240,I88054,I88033);
not I_17091 (I293257,I293240);
nor I_17092 (I292819,I293096,I293257);
nand I_17093 (I292804,I293113,I293257);
nor I_17094 (I292813,I292859,I293240);
DFFARX1 I_17095 (I293240,I2683,I292833,I292822,);
not I_17096 (I293360,I2690);
DFFARX1 I_17097 (I986416,I2683,I293360,I293386,);
nand I_17098 (I293394,I986398,I986422);
and I_17099 (I293411,I293394,I986413);
DFFARX1 I_17100 (I293411,I2683,I293360,I293437,);
nor I_17101 (I293328,I293437,I293386);
not I_17102 (I293459,I293437);
DFFARX1 I_17103 (I986419,I2683,I293360,I293485,);
nand I_17104 (I293493,I293485,I986407);
not I_17105 (I293510,I293493);
DFFARX1 I_17106 (I293510,I2683,I293360,I293536,);
not I_17107 (I293352,I293536);
nor I_17108 (I293558,I293386,I293493);
nor I_17109 (I293334,I293437,I293558);
DFFARX1 I_17110 (I986398,I2683,I293360,I293598,);
DFFARX1 I_17111 (I293598,I2683,I293360,I293615,);
not I_17112 (I293623,I293615);
not I_17113 (I293640,I293598);
nand I_17114 (I293337,I293640,I293459);
nand I_17115 (I293671,I986404,I986401);
and I_17116 (I293688,I293671,I986410);
DFFARX1 I_17117 (I293688,I2683,I293360,I293714,);
nor I_17118 (I293722,I293714,I293386);
DFFARX1 I_17119 (I293722,I2683,I293360,I293325,);
DFFARX1 I_17120 (I293714,I2683,I293360,I293343,);
nor I_17121 (I293767,I986401,I986401);
not I_17122 (I293784,I293767);
nor I_17123 (I293346,I293623,I293784);
nand I_17124 (I293331,I293640,I293784);
nor I_17125 (I293340,I293386,I293767);
DFFARX1 I_17126 (I293767,I2683,I293360,I293349,);
not I_17127 (I293887,I2690);
DFFARX1 I_17128 (I701260,I2683,I293887,I293913,);
nand I_17129 (I293921,I701257,I701275);
and I_17130 (I293938,I293921,I701266);
DFFARX1 I_17131 (I293938,I2683,I293887,I293964,);
nor I_17132 (I293855,I293964,I293913);
not I_17133 (I293986,I293964);
DFFARX1 I_17134 (I701281,I2683,I293887,I294012,);
nand I_17135 (I294020,I294012,I701263);
not I_17136 (I294037,I294020);
DFFARX1 I_17137 (I294037,I2683,I293887,I294063,);
not I_17138 (I293879,I294063);
nor I_17139 (I294085,I293913,I294020);
nor I_17140 (I293861,I293964,I294085);
DFFARX1 I_17141 (I701269,I2683,I293887,I294125,);
DFFARX1 I_17142 (I294125,I2683,I293887,I294142,);
not I_17143 (I294150,I294142);
not I_17144 (I294167,I294125);
nand I_17145 (I293864,I294167,I293986);
nand I_17146 (I294198,I701257,I701284);
and I_17147 (I294215,I294198,I701272);
DFFARX1 I_17148 (I294215,I2683,I293887,I294241,);
nor I_17149 (I294249,I294241,I293913);
DFFARX1 I_17150 (I294249,I2683,I293887,I293852,);
DFFARX1 I_17151 (I294241,I2683,I293887,I293870,);
nor I_17152 (I294294,I701278,I701284);
not I_17153 (I294311,I294294);
nor I_17154 (I293873,I294150,I294311);
nand I_17155 (I293858,I294167,I294311);
nor I_17156 (I293867,I293913,I294294);
DFFARX1 I_17157 (I294294,I2683,I293887,I293876,);
not I_17158 (I294414,I2690);
DFFARX1 I_17159 (I872124,I2683,I294414,I294440,);
nand I_17160 (I294448,I872139,I872124);
and I_17161 (I294465,I294448,I872142);
DFFARX1 I_17162 (I294465,I2683,I294414,I294491,);
nor I_17163 (I294382,I294491,I294440);
not I_17164 (I294513,I294491);
DFFARX1 I_17165 (I872148,I2683,I294414,I294539,);
nand I_17166 (I294547,I294539,I872130);
not I_17167 (I294564,I294547);
DFFARX1 I_17168 (I294564,I2683,I294414,I294590,);
not I_17169 (I294406,I294590);
nor I_17170 (I294612,I294440,I294547);
nor I_17171 (I294388,I294491,I294612);
DFFARX1 I_17172 (I872127,I2683,I294414,I294652,);
DFFARX1 I_17173 (I294652,I2683,I294414,I294669,);
not I_17174 (I294677,I294669);
not I_17175 (I294694,I294652);
nand I_17176 (I294391,I294694,I294513);
nand I_17177 (I294725,I872127,I872133);
and I_17178 (I294742,I294725,I872145);
DFFARX1 I_17179 (I294742,I2683,I294414,I294768,);
nor I_17180 (I294776,I294768,I294440);
DFFARX1 I_17181 (I294776,I2683,I294414,I294379,);
DFFARX1 I_17182 (I294768,I2683,I294414,I294397,);
nor I_17183 (I294821,I872136,I872133);
not I_17184 (I294838,I294821);
nor I_17185 (I294400,I294677,I294838);
nand I_17186 (I294385,I294694,I294838);
nor I_17187 (I294394,I294440,I294821);
DFFARX1 I_17188 (I294821,I2683,I294414,I294403,);
not I_17189 (I294941,I2690);
DFFARX1 I_17190 (I554950,I2683,I294941,I294967,);
nand I_17191 (I294975,I554941,I554956);
and I_17192 (I294992,I294975,I554962);
DFFARX1 I_17193 (I294992,I2683,I294941,I295018,);
nor I_17194 (I294909,I295018,I294967);
not I_17195 (I295040,I295018);
DFFARX1 I_17196 (I554947,I2683,I294941,I295066,);
nand I_17197 (I295074,I295066,I554941);
not I_17198 (I295091,I295074);
DFFARX1 I_17199 (I295091,I2683,I294941,I295117,);
not I_17200 (I294933,I295117);
nor I_17201 (I295139,I294967,I295074);
nor I_17202 (I294915,I295018,I295139);
DFFARX1 I_17203 (I554944,I2683,I294941,I295179,);
DFFARX1 I_17204 (I295179,I2683,I294941,I295196,);
not I_17205 (I295204,I295196);
not I_17206 (I295221,I295179);
nand I_17207 (I294918,I295221,I295040);
nand I_17208 (I295252,I554938,I554953);
and I_17209 (I295269,I295252,I554938);
DFFARX1 I_17210 (I295269,I2683,I294941,I295295,);
nor I_17211 (I295303,I295295,I294967);
DFFARX1 I_17212 (I295303,I2683,I294941,I294906,);
DFFARX1 I_17213 (I295295,I2683,I294941,I294924,);
nor I_17214 (I295348,I554959,I554953);
not I_17215 (I295365,I295348);
nor I_17216 (I294927,I295204,I295365);
nand I_17217 (I294912,I295221,I295365);
nor I_17218 (I294921,I294967,I295348);
DFFARX1 I_17219 (I295348,I2683,I294941,I294930,);
not I_17220 (I295468,I2690);
DFFARX1 I_17221 (I594254,I2683,I295468,I295494,);
nand I_17222 (I295502,I594245,I594260);
and I_17223 (I295519,I295502,I594266);
DFFARX1 I_17224 (I295519,I2683,I295468,I295545,);
nor I_17225 (I295436,I295545,I295494);
not I_17226 (I295567,I295545);
DFFARX1 I_17227 (I594251,I2683,I295468,I295593,);
nand I_17228 (I295601,I295593,I594245);
not I_17229 (I295618,I295601);
DFFARX1 I_17230 (I295618,I2683,I295468,I295644,);
not I_17231 (I295460,I295644);
nor I_17232 (I295666,I295494,I295601);
nor I_17233 (I295442,I295545,I295666);
DFFARX1 I_17234 (I594248,I2683,I295468,I295706,);
DFFARX1 I_17235 (I295706,I2683,I295468,I295723,);
not I_17236 (I295731,I295723);
not I_17237 (I295748,I295706);
nand I_17238 (I295445,I295748,I295567);
nand I_17239 (I295779,I594242,I594257);
and I_17240 (I295796,I295779,I594242);
DFFARX1 I_17241 (I295796,I2683,I295468,I295822,);
nor I_17242 (I295830,I295822,I295494);
DFFARX1 I_17243 (I295830,I2683,I295468,I295433,);
DFFARX1 I_17244 (I295822,I2683,I295468,I295451,);
nor I_17245 (I295875,I594263,I594257);
not I_17246 (I295892,I295875);
nor I_17247 (I295454,I295731,I295892);
nand I_17248 (I295439,I295748,I295892);
nor I_17249 (I295448,I295494,I295875);
DFFARX1 I_17250 (I295875,I2683,I295468,I295457,);
not I_17251 (I295995,I2690);
DFFARX1 I_17252 (I752940,I2683,I295995,I296021,);
nand I_17253 (I296029,I752937,I752955);
and I_17254 (I296046,I296029,I752946);
DFFARX1 I_17255 (I296046,I2683,I295995,I296072,);
nor I_17256 (I295963,I296072,I296021);
not I_17257 (I296094,I296072);
DFFARX1 I_17258 (I752961,I2683,I295995,I296120,);
nand I_17259 (I296128,I296120,I752943);
not I_17260 (I296145,I296128);
DFFARX1 I_17261 (I296145,I2683,I295995,I296171,);
not I_17262 (I295987,I296171);
nor I_17263 (I296193,I296021,I296128);
nor I_17264 (I295969,I296072,I296193);
DFFARX1 I_17265 (I752949,I2683,I295995,I296233,);
DFFARX1 I_17266 (I296233,I2683,I295995,I296250,);
not I_17267 (I296258,I296250);
not I_17268 (I296275,I296233);
nand I_17269 (I295972,I296275,I296094);
nand I_17270 (I296306,I752937,I752964);
and I_17271 (I296323,I296306,I752952);
DFFARX1 I_17272 (I296323,I2683,I295995,I296349,);
nor I_17273 (I296357,I296349,I296021);
DFFARX1 I_17274 (I296357,I2683,I295995,I295960,);
DFFARX1 I_17275 (I296349,I2683,I295995,I295978,);
nor I_17276 (I296402,I752958,I752964);
not I_17277 (I296419,I296402);
nor I_17278 (I295981,I296258,I296419);
nand I_17279 (I295966,I296275,I296419);
nor I_17280 (I295975,I296021,I296402);
DFFARX1 I_17281 (I296402,I2683,I295995,I295984,);
not I_17282 (I296522,I2690);
DFFARX1 I_17283 (I408605,I2683,I296522,I296548,);
nand I_17284 (I296556,I408605,I408617);
and I_17285 (I296573,I296556,I408602);
DFFARX1 I_17286 (I296573,I2683,I296522,I296599,);
nor I_17287 (I296490,I296599,I296548);
not I_17288 (I296621,I296599);
DFFARX1 I_17289 (I408626,I2683,I296522,I296647,);
nand I_17290 (I296655,I296647,I408623);
not I_17291 (I296672,I296655);
DFFARX1 I_17292 (I296672,I2683,I296522,I296698,);
not I_17293 (I296514,I296698);
nor I_17294 (I296720,I296548,I296655);
nor I_17295 (I296496,I296599,I296720);
DFFARX1 I_17296 (I408614,I2683,I296522,I296760,);
DFFARX1 I_17297 (I296760,I2683,I296522,I296777,);
not I_17298 (I296785,I296777);
not I_17299 (I296802,I296760);
nand I_17300 (I296499,I296802,I296621);
nand I_17301 (I296833,I408602,I408611);
and I_17302 (I296850,I296833,I408620);
DFFARX1 I_17303 (I296850,I2683,I296522,I296876,);
nor I_17304 (I296884,I296876,I296548);
DFFARX1 I_17305 (I296884,I2683,I296522,I296487,);
DFFARX1 I_17306 (I296876,I2683,I296522,I296505,);
nor I_17307 (I296929,I408608,I408611);
not I_17308 (I296946,I296929);
nor I_17309 (I296508,I296785,I296946);
nand I_17310 (I296493,I296802,I296946);
nor I_17311 (I296502,I296548,I296929);
DFFARX1 I_17312 (I296929,I2683,I296522,I296511,);
not I_17313 (I297049,I2690);
DFFARX1 I_17314 (I905648,I2683,I297049,I297075,);
nand I_17315 (I297083,I905663,I905648);
and I_17316 (I297100,I297083,I905666);
DFFARX1 I_17317 (I297100,I2683,I297049,I297126,);
nor I_17318 (I297017,I297126,I297075);
not I_17319 (I297148,I297126);
DFFARX1 I_17320 (I905672,I2683,I297049,I297174,);
nand I_17321 (I297182,I297174,I905654);
not I_17322 (I297199,I297182);
DFFARX1 I_17323 (I297199,I2683,I297049,I297225,);
not I_17324 (I297041,I297225);
nor I_17325 (I297247,I297075,I297182);
nor I_17326 (I297023,I297126,I297247);
DFFARX1 I_17327 (I905651,I2683,I297049,I297287,);
DFFARX1 I_17328 (I297287,I2683,I297049,I297304,);
not I_17329 (I297312,I297304);
not I_17330 (I297329,I297287);
nand I_17331 (I297026,I297329,I297148);
nand I_17332 (I297360,I905651,I905657);
and I_17333 (I297377,I297360,I905669);
DFFARX1 I_17334 (I297377,I2683,I297049,I297403,);
nor I_17335 (I297411,I297403,I297075);
DFFARX1 I_17336 (I297411,I2683,I297049,I297014,);
DFFARX1 I_17337 (I297403,I2683,I297049,I297032,);
nor I_17338 (I297456,I905660,I905657);
not I_17339 (I297473,I297456);
nor I_17340 (I297035,I297312,I297473);
nand I_17341 (I297020,I297329,I297473);
nor I_17342 (I297029,I297075,I297456);
DFFARX1 I_17343 (I297456,I2683,I297049,I297038,);
not I_17344 (I297576,I2690);
DFFARX1 I_17345 (I711596,I2683,I297576,I297602,);
nand I_17346 (I297610,I711593,I711611);
and I_17347 (I297627,I297610,I711602);
DFFARX1 I_17348 (I297627,I2683,I297576,I297653,);
nor I_17349 (I297544,I297653,I297602);
not I_17350 (I297675,I297653);
DFFARX1 I_17351 (I711617,I2683,I297576,I297701,);
nand I_17352 (I297709,I297701,I711599);
not I_17353 (I297726,I297709);
DFFARX1 I_17354 (I297726,I2683,I297576,I297752,);
not I_17355 (I297568,I297752);
nor I_17356 (I297774,I297602,I297709);
nor I_17357 (I297550,I297653,I297774);
DFFARX1 I_17358 (I711605,I2683,I297576,I297814,);
DFFARX1 I_17359 (I297814,I2683,I297576,I297831,);
not I_17360 (I297839,I297831);
not I_17361 (I297856,I297814);
nand I_17362 (I297553,I297856,I297675);
nand I_17363 (I297887,I711593,I711620);
and I_17364 (I297904,I297887,I711608);
DFFARX1 I_17365 (I297904,I2683,I297576,I297930,);
nor I_17366 (I297938,I297930,I297602);
DFFARX1 I_17367 (I297938,I2683,I297576,I297541,);
DFFARX1 I_17368 (I297930,I2683,I297576,I297559,);
nor I_17369 (I297983,I711614,I711620);
not I_17370 (I298000,I297983);
nor I_17371 (I297562,I297839,I298000);
nand I_17372 (I297547,I297856,I298000);
nor I_17373 (I297556,I297602,I297983);
DFFARX1 I_17374 (I297983,I2683,I297576,I297565,);
not I_17375 (I298103,I2690);
DFFARX1 I_17376 (I991479,I2683,I298103,I298129,);
nand I_17377 (I298137,I991476,I991467);
and I_17378 (I298154,I298137,I991464);
DFFARX1 I_17379 (I298154,I2683,I298103,I298180,);
nor I_17380 (I298071,I298180,I298129);
not I_17381 (I298202,I298180);
DFFARX1 I_17382 (I991473,I2683,I298103,I298228,);
nand I_17383 (I298236,I298228,I991482);
not I_17384 (I298253,I298236);
DFFARX1 I_17385 (I298253,I2683,I298103,I298279,);
not I_17386 (I298095,I298279);
nor I_17387 (I298301,I298129,I298236);
nor I_17388 (I298077,I298180,I298301);
DFFARX1 I_17389 (I991485,I2683,I298103,I298341,);
DFFARX1 I_17390 (I298341,I2683,I298103,I298358,);
not I_17391 (I298366,I298358);
not I_17392 (I298383,I298341);
nand I_17393 (I298080,I298383,I298202);
nand I_17394 (I298414,I991464,I991470);
and I_17395 (I298431,I298414,I991488);
DFFARX1 I_17396 (I298431,I2683,I298103,I298457,);
nor I_17397 (I298465,I298457,I298129);
DFFARX1 I_17398 (I298465,I2683,I298103,I298068,);
DFFARX1 I_17399 (I298457,I2683,I298103,I298086,);
nor I_17400 (I298510,I991467,I991470);
not I_17401 (I298527,I298510);
nor I_17402 (I298089,I298366,I298527);
nand I_17403 (I298074,I298383,I298527);
nor I_17404 (I298083,I298129,I298510);
DFFARX1 I_17405 (I298510,I2683,I298103,I298092,);
not I_17406 (I298630,I2690);
DFFARX1 I_17407 (I840334,I2683,I298630,I298656,);
nand I_17408 (I298664,I840349,I840334);
and I_17409 (I298681,I298664,I840352);
DFFARX1 I_17410 (I298681,I2683,I298630,I298707,);
nor I_17411 (I298598,I298707,I298656);
not I_17412 (I298729,I298707);
DFFARX1 I_17413 (I840358,I2683,I298630,I298755,);
nand I_17414 (I298763,I298755,I840340);
not I_17415 (I298780,I298763);
DFFARX1 I_17416 (I298780,I2683,I298630,I298806,);
not I_17417 (I298622,I298806);
nor I_17418 (I298828,I298656,I298763);
nor I_17419 (I298604,I298707,I298828);
DFFARX1 I_17420 (I840337,I2683,I298630,I298868,);
DFFARX1 I_17421 (I298868,I2683,I298630,I298885,);
not I_17422 (I298893,I298885);
not I_17423 (I298910,I298868);
nand I_17424 (I298607,I298910,I298729);
nand I_17425 (I298941,I840337,I840343);
and I_17426 (I298958,I298941,I840355);
DFFARX1 I_17427 (I298958,I2683,I298630,I298984,);
nor I_17428 (I298992,I298984,I298656);
DFFARX1 I_17429 (I298992,I2683,I298630,I298595,);
DFFARX1 I_17430 (I298984,I2683,I298630,I298613,);
nor I_17431 (I299037,I840346,I840343);
not I_17432 (I299054,I299037);
nor I_17433 (I298616,I298893,I299054);
nand I_17434 (I298601,I298910,I299054);
nor I_17435 (I298610,I298656,I299037);
DFFARX1 I_17436 (I299037,I2683,I298630,I298619,);
not I_17437 (I299157,I2690);
DFFARX1 I_17438 (I118249,I2683,I299157,I299183,);
nand I_17439 (I299191,I118234,I118225);
and I_17440 (I299208,I299191,I118240);
DFFARX1 I_17441 (I299208,I2683,I299157,I299234,);
nor I_17442 (I299125,I299234,I299183);
not I_17443 (I299256,I299234);
DFFARX1 I_17444 (I118252,I2683,I299157,I299282,);
nand I_17445 (I299290,I299282,I118243);
not I_17446 (I299307,I299290);
DFFARX1 I_17447 (I299307,I2683,I299157,I299333,);
not I_17448 (I299149,I299333);
nor I_17449 (I299355,I299183,I299290);
nor I_17450 (I299131,I299234,I299355);
DFFARX1 I_17451 (I118231,I2683,I299157,I299395,);
DFFARX1 I_17452 (I299395,I2683,I299157,I299412,);
not I_17453 (I299420,I299412);
not I_17454 (I299437,I299395);
nand I_17455 (I299134,I299437,I299256);
nand I_17456 (I299468,I118237,I118228);
and I_17457 (I299485,I299468,I118225);
DFFARX1 I_17458 (I299485,I2683,I299157,I299511,);
nor I_17459 (I299519,I299511,I299183);
DFFARX1 I_17460 (I299519,I2683,I299157,I299122,);
DFFARX1 I_17461 (I299511,I2683,I299157,I299140,);
nor I_17462 (I299564,I118246,I118228);
not I_17463 (I299581,I299564);
nor I_17464 (I299143,I299420,I299581);
nand I_17465 (I299128,I299437,I299581);
nor I_17466 (I299137,I299183,I299564);
DFFARX1 I_17467 (I299564,I2683,I299157,I299146,);
not I_17468 (I299684,I2690);
DFFARX1 I_17469 (I959760,I2683,I299684,I299710,);
nand I_17470 (I299718,I959742,I959766);
and I_17471 (I299735,I299718,I959757);
DFFARX1 I_17472 (I299735,I2683,I299684,I299761,);
nor I_17473 (I299652,I299761,I299710);
not I_17474 (I299783,I299761);
DFFARX1 I_17475 (I959763,I2683,I299684,I299809,);
nand I_17476 (I299817,I299809,I959751);
not I_17477 (I299834,I299817);
DFFARX1 I_17478 (I299834,I2683,I299684,I299860,);
not I_17479 (I299676,I299860);
nor I_17480 (I299882,I299710,I299817);
nor I_17481 (I299658,I299761,I299882);
DFFARX1 I_17482 (I959742,I2683,I299684,I299922,);
DFFARX1 I_17483 (I299922,I2683,I299684,I299939,);
not I_17484 (I299947,I299939);
not I_17485 (I299964,I299922);
nand I_17486 (I299661,I299964,I299783);
nand I_17487 (I299995,I959748,I959745);
and I_17488 (I300012,I299995,I959754);
DFFARX1 I_17489 (I300012,I2683,I299684,I300038,);
nor I_17490 (I300046,I300038,I299710);
DFFARX1 I_17491 (I300046,I2683,I299684,I299649,);
DFFARX1 I_17492 (I300038,I2683,I299684,I299667,);
nor I_17493 (I300091,I959745,I959745);
not I_17494 (I300108,I300091);
nor I_17495 (I299670,I299947,I300108);
nand I_17496 (I299655,I299964,I300108);
nor I_17497 (I299664,I299710,I300091);
DFFARX1 I_17498 (I300091,I2683,I299684,I299673,);
not I_17499 (I300211,I2690);
DFFARX1 I_17500 (I152140,I2683,I300211,I300237,);
nand I_17501 (I300245,I152140,I152146);
and I_17502 (I300262,I300245,I152164);
DFFARX1 I_17503 (I300262,I2683,I300211,I300288,);
nor I_17504 (I300179,I300288,I300237);
not I_17505 (I300310,I300288);
DFFARX1 I_17506 (I152152,I2683,I300211,I300336,);
nand I_17507 (I300344,I300336,I152149);
not I_17508 (I300361,I300344);
DFFARX1 I_17509 (I300361,I2683,I300211,I300387,);
not I_17510 (I300203,I300387);
nor I_17511 (I300409,I300237,I300344);
nor I_17512 (I300185,I300288,I300409);
DFFARX1 I_17513 (I152158,I2683,I300211,I300449,);
DFFARX1 I_17514 (I300449,I2683,I300211,I300466,);
not I_17515 (I300474,I300466);
not I_17516 (I300491,I300449);
nand I_17517 (I300188,I300491,I300310);
nand I_17518 (I300522,I152143,I152143);
and I_17519 (I300539,I300522,I152155);
DFFARX1 I_17520 (I300539,I2683,I300211,I300565,);
nor I_17521 (I300573,I300565,I300237);
DFFARX1 I_17522 (I300573,I2683,I300211,I300176,);
DFFARX1 I_17523 (I300565,I2683,I300211,I300194,);
nor I_17524 (I300618,I152161,I152143);
not I_17525 (I300635,I300618);
nor I_17526 (I300197,I300474,I300635);
nand I_17527 (I300182,I300491,I300635);
nor I_17528 (I300191,I300237,I300618);
DFFARX1 I_17529 (I300618,I2683,I300211,I300200,);
not I_17530 (I300738,I2690);
DFFARX1 I_17531 (I113489,I2683,I300738,I300764,);
nand I_17532 (I300772,I113474,I113465);
and I_17533 (I300789,I300772,I113480);
DFFARX1 I_17534 (I300789,I2683,I300738,I300815,);
nor I_17535 (I300706,I300815,I300764);
not I_17536 (I300837,I300815);
DFFARX1 I_17537 (I113492,I2683,I300738,I300863,);
nand I_17538 (I300871,I300863,I113483);
not I_17539 (I300888,I300871);
DFFARX1 I_17540 (I300888,I2683,I300738,I300914,);
not I_17541 (I300730,I300914);
nor I_17542 (I300936,I300764,I300871);
nor I_17543 (I300712,I300815,I300936);
DFFARX1 I_17544 (I113471,I2683,I300738,I300976,);
DFFARX1 I_17545 (I300976,I2683,I300738,I300993,);
not I_17546 (I301001,I300993);
not I_17547 (I301018,I300976);
nand I_17548 (I300715,I301018,I300837);
nand I_17549 (I301049,I113477,I113468);
and I_17550 (I301066,I301049,I113465);
DFFARX1 I_17551 (I301066,I2683,I300738,I301092,);
nor I_17552 (I301100,I301092,I300764);
DFFARX1 I_17553 (I301100,I2683,I300738,I300703,);
DFFARX1 I_17554 (I301092,I2683,I300738,I300721,);
nor I_17555 (I301145,I113486,I113468);
not I_17556 (I301162,I301145);
nor I_17557 (I300724,I301001,I301162);
nand I_17558 (I300709,I301018,I301162);
nor I_17559 (I300718,I300764,I301145);
DFFARX1 I_17560 (I301145,I2683,I300738,I300727,);
not I_17561 (I301265,I2690);
DFFARX1 I_17562 (I693933,I2683,I301265,I301291,);
nand I_17563 (I301299,I693936,I693930);
and I_17564 (I301316,I301299,I693942);
DFFARX1 I_17565 (I301316,I2683,I301265,I301342,);
nor I_17566 (I301233,I301342,I301291);
not I_17567 (I301364,I301342);
DFFARX1 I_17568 (I693945,I2683,I301265,I301390,);
nand I_17569 (I301398,I301390,I693936);
not I_17570 (I301415,I301398);
DFFARX1 I_17571 (I301415,I2683,I301265,I301441,);
not I_17572 (I301257,I301441);
nor I_17573 (I301463,I301291,I301398);
nor I_17574 (I301239,I301342,I301463);
DFFARX1 I_17575 (I693948,I2683,I301265,I301503,);
DFFARX1 I_17576 (I301503,I2683,I301265,I301520,);
not I_17577 (I301528,I301520);
not I_17578 (I301545,I301503);
nand I_17579 (I301242,I301545,I301364);
nand I_17580 (I301576,I693930,I693939);
and I_17581 (I301593,I301576,I693933);
DFFARX1 I_17582 (I301593,I2683,I301265,I301619,);
nor I_17583 (I301627,I301619,I301291);
DFFARX1 I_17584 (I301627,I2683,I301265,I301230,);
DFFARX1 I_17585 (I301619,I2683,I301265,I301248,);
nor I_17586 (I301672,I693951,I693939);
not I_17587 (I301689,I301672);
nor I_17588 (I301251,I301528,I301689);
nand I_17589 (I301236,I301545,I301689);
nor I_17590 (I301245,I301291,I301672);
DFFARX1 I_17591 (I301672,I2683,I301265,I301254,);
not I_17592 (I301792,I2690);
DFFARX1 I_17593 (I1095950,I2683,I301792,I301818,);
nand I_17594 (I301826,I1095929,I1095929);
and I_17595 (I301843,I301826,I1095956);
DFFARX1 I_17596 (I301843,I2683,I301792,I301869,);
nor I_17597 (I301760,I301869,I301818);
not I_17598 (I301891,I301869);
DFFARX1 I_17599 (I1095944,I2683,I301792,I301917,);
nand I_17600 (I301925,I301917,I1095947);
not I_17601 (I301942,I301925);
DFFARX1 I_17602 (I301942,I2683,I301792,I301968,);
not I_17603 (I301784,I301968);
nor I_17604 (I301990,I301818,I301925);
nor I_17605 (I301766,I301869,I301990);
DFFARX1 I_17606 (I1095938,I2683,I301792,I302030,);
DFFARX1 I_17607 (I302030,I2683,I301792,I302047,);
not I_17608 (I302055,I302047);
not I_17609 (I302072,I302030);
nand I_17610 (I301769,I302072,I301891);
nand I_17611 (I302103,I1095935,I1095932);
and I_17612 (I302120,I302103,I1095953);
DFFARX1 I_17613 (I302120,I2683,I301792,I302146,);
nor I_17614 (I302154,I302146,I301818);
DFFARX1 I_17615 (I302154,I2683,I301792,I301757,);
DFFARX1 I_17616 (I302146,I2683,I301792,I301775,);
nor I_17617 (I302199,I1095941,I1095932);
not I_17618 (I302216,I302199);
nor I_17619 (I301778,I302055,I302216);
nand I_17620 (I301763,I302072,I302216);
nor I_17621 (I301772,I301818,I302199);
DFFARX1 I_17622 (I302199,I2683,I301792,I301781,);
not I_17623 (I302319,I2690);
DFFARX1 I_17624 (I811930,I2683,I302319,I302345,);
nand I_17625 (I302353,I811927,I811930);
and I_17626 (I302370,I302353,I811939);
DFFARX1 I_17627 (I302370,I2683,I302319,I302396,);
nor I_17628 (I302287,I302396,I302345);
not I_17629 (I302418,I302396);
DFFARX1 I_17630 (I811927,I2683,I302319,I302444,);
nand I_17631 (I302452,I302444,I811945);
not I_17632 (I302469,I302452);
DFFARX1 I_17633 (I302469,I2683,I302319,I302495,);
not I_17634 (I302311,I302495);
nor I_17635 (I302517,I302345,I302452);
nor I_17636 (I302293,I302396,I302517);
DFFARX1 I_17637 (I811933,I2683,I302319,I302557,);
DFFARX1 I_17638 (I302557,I2683,I302319,I302574,);
not I_17639 (I302582,I302574);
not I_17640 (I302599,I302557);
nand I_17641 (I302296,I302599,I302418);
nand I_17642 (I302630,I811942,I811948);
and I_17643 (I302647,I302630,I811933);
DFFARX1 I_17644 (I302647,I2683,I302319,I302673,);
nor I_17645 (I302681,I302673,I302345);
DFFARX1 I_17646 (I302681,I2683,I302319,I302284,);
DFFARX1 I_17647 (I302673,I2683,I302319,I302302,);
nor I_17648 (I302726,I811936,I811948);
not I_17649 (I302743,I302726);
nor I_17650 (I302305,I302582,I302743);
nand I_17651 (I302290,I302599,I302743);
nor I_17652 (I302299,I302345,I302726);
DFFARX1 I_17653 (I302726,I2683,I302319,I302308,);
not I_17654 (I302846,I2690);
DFFARX1 I_17655 (I448023,I2683,I302846,I302872,);
nand I_17656 (I302880,I448008,I448011);
and I_17657 (I302897,I302880,I448026);
DFFARX1 I_17658 (I302897,I2683,I302846,I302923,);
nor I_17659 (I302814,I302923,I302872);
not I_17660 (I302945,I302923);
DFFARX1 I_17661 (I448020,I2683,I302846,I302971,);
nand I_17662 (I302979,I302971,I448011);
not I_17663 (I302996,I302979);
DFFARX1 I_17664 (I302996,I2683,I302846,I303022,);
not I_17665 (I302838,I303022);
nor I_17666 (I303044,I302872,I302979);
nor I_17667 (I302820,I302923,I303044);
DFFARX1 I_17668 (I448017,I2683,I302846,I303084,);
DFFARX1 I_17669 (I303084,I2683,I302846,I303101,);
not I_17670 (I303109,I303101);
not I_17671 (I303126,I303084);
nand I_17672 (I302823,I303126,I302945);
nand I_17673 (I303157,I448032,I448008);
and I_17674 (I303174,I303157,I448029);
DFFARX1 I_17675 (I303174,I2683,I302846,I303200,);
nor I_17676 (I303208,I303200,I302872);
DFFARX1 I_17677 (I303208,I2683,I302846,I302811,);
DFFARX1 I_17678 (I303200,I2683,I302846,I302829,);
nor I_17679 (I303253,I448014,I448008);
not I_17680 (I303270,I303253);
nor I_17681 (I302832,I303109,I303270);
nand I_17682 (I302817,I303126,I303270);
nor I_17683 (I302826,I302872,I303253);
DFFARX1 I_17684 (I303253,I2683,I302846,I302835,);
not I_17685 (I303373,I2690);
DFFARX1 I_17686 (I492529,I2683,I303373,I303399,);
nand I_17687 (I303407,I492514,I492517);
and I_17688 (I303424,I303407,I492532);
DFFARX1 I_17689 (I303424,I2683,I303373,I303450,);
nor I_17690 (I303341,I303450,I303399);
not I_17691 (I303472,I303450);
DFFARX1 I_17692 (I492526,I2683,I303373,I303498,);
nand I_17693 (I303506,I303498,I492517);
not I_17694 (I303523,I303506);
DFFARX1 I_17695 (I303523,I2683,I303373,I303549,);
not I_17696 (I303365,I303549);
nor I_17697 (I303571,I303399,I303506);
nor I_17698 (I303347,I303450,I303571);
DFFARX1 I_17699 (I492523,I2683,I303373,I303611,);
DFFARX1 I_17700 (I303611,I2683,I303373,I303628,);
not I_17701 (I303636,I303628);
not I_17702 (I303653,I303611);
nand I_17703 (I303350,I303653,I303472);
nand I_17704 (I303684,I492538,I492514);
and I_17705 (I303701,I303684,I492535);
DFFARX1 I_17706 (I303701,I2683,I303373,I303727,);
nor I_17707 (I303735,I303727,I303399);
DFFARX1 I_17708 (I303735,I2683,I303373,I303338,);
DFFARX1 I_17709 (I303727,I2683,I303373,I303356,);
nor I_17710 (I303780,I492520,I492514);
not I_17711 (I303797,I303780);
nor I_17712 (I303359,I303636,I303797);
nand I_17713 (I303344,I303653,I303797);
nor I_17714 (I303353,I303399,I303780);
DFFARX1 I_17715 (I303780,I2683,I303373,I303362,);
not I_17716 (I303900,I2690);
DFFARX1 I_17717 (I825394,I2683,I303900,I303926,);
nand I_17718 (I303934,I825391,I825394);
and I_17719 (I303951,I303934,I825403);
DFFARX1 I_17720 (I303951,I2683,I303900,I303977,);
nor I_17721 (I303868,I303977,I303926);
not I_17722 (I303999,I303977);
DFFARX1 I_17723 (I825391,I2683,I303900,I304025,);
nand I_17724 (I304033,I304025,I825409);
not I_17725 (I304050,I304033);
DFFARX1 I_17726 (I304050,I2683,I303900,I304076,);
not I_17727 (I303892,I304076);
nor I_17728 (I304098,I303926,I304033);
nor I_17729 (I303874,I303977,I304098);
DFFARX1 I_17730 (I825397,I2683,I303900,I304138,);
DFFARX1 I_17731 (I304138,I2683,I303900,I304155,);
not I_17732 (I304163,I304155);
not I_17733 (I304180,I304138);
nand I_17734 (I303877,I304180,I303999);
nand I_17735 (I304211,I825406,I825412);
and I_17736 (I304228,I304211,I825397);
DFFARX1 I_17737 (I304228,I2683,I303900,I304254,);
nor I_17738 (I304262,I304254,I303926);
DFFARX1 I_17739 (I304262,I2683,I303900,I303865,);
DFFARX1 I_17740 (I304254,I2683,I303900,I303883,);
nor I_17741 (I304307,I825400,I825412);
not I_17742 (I304324,I304307);
nor I_17743 (I303886,I304163,I304324);
nand I_17744 (I303871,I304180,I304324);
nor I_17745 (I303880,I303926,I304307);
DFFARX1 I_17746 (I304307,I2683,I303900,I303889,);
not I_17747 (I304427,I2690);
DFFARX1 I_17748 (I813613,I2683,I304427,I304453,);
nand I_17749 (I304461,I813610,I813613);
and I_17750 (I304478,I304461,I813622);
DFFARX1 I_17751 (I304478,I2683,I304427,I304504,);
nor I_17752 (I304395,I304504,I304453);
not I_17753 (I304526,I304504);
DFFARX1 I_17754 (I813610,I2683,I304427,I304552,);
nand I_17755 (I304560,I304552,I813628);
not I_17756 (I304577,I304560);
DFFARX1 I_17757 (I304577,I2683,I304427,I304603,);
not I_17758 (I304419,I304603);
nor I_17759 (I304625,I304453,I304560);
nor I_17760 (I304401,I304504,I304625);
DFFARX1 I_17761 (I813616,I2683,I304427,I304665,);
DFFARX1 I_17762 (I304665,I2683,I304427,I304682,);
not I_17763 (I304690,I304682);
not I_17764 (I304707,I304665);
nand I_17765 (I304404,I304707,I304526);
nand I_17766 (I304738,I813625,I813631);
and I_17767 (I304755,I304738,I813616);
DFFARX1 I_17768 (I304755,I2683,I304427,I304781,);
nor I_17769 (I304789,I304781,I304453);
DFFARX1 I_17770 (I304789,I2683,I304427,I304392,);
DFFARX1 I_17771 (I304781,I2683,I304427,I304410,);
nor I_17772 (I304834,I813619,I813631);
not I_17773 (I304851,I304834);
nor I_17774 (I304413,I304690,I304851);
nand I_17775 (I304398,I304707,I304851);
nor I_17776 (I304407,I304453,I304834);
DFFARX1 I_17777 (I304834,I2683,I304427,I304416,);
not I_17778 (I304954,I2690);
DFFARX1 I_17779 (I1030500,I2683,I304954,I304980,);
nand I_17780 (I304988,I1030479,I1030479);
and I_17781 (I305005,I304988,I1030506);
DFFARX1 I_17782 (I305005,I2683,I304954,I305031,);
nor I_17783 (I304922,I305031,I304980);
not I_17784 (I305053,I305031);
DFFARX1 I_17785 (I1030494,I2683,I304954,I305079,);
nand I_17786 (I305087,I305079,I1030497);
not I_17787 (I305104,I305087);
DFFARX1 I_17788 (I305104,I2683,I304954,I305130,);
not I_17789 (I304946,I305130);
nor I_17790 (I305152,I304980,I305087);
nor I_17791 (I304928,I305031,I305152);
DFFARX1 I_17792 (I1030488,I2683,I304954,I305192,);
DFFARX1 I_17793 (I305192,I2683,I304954,I305209,);
not I_17794 (I305217,I305209);
not I_17795 (I305234,I305192);
nand I_17796 (I304931,I305234,I305053);
nand I_17797 (I305265,I1030485,I1030482);
and I_17798 (I305282,I305265,I1030503);
DFFARX1 I_17799 (I305282,I2683,I304954,I305308,);
nor I_17800 (I305316,I305308,I304980);
DFFARX1 I_17801 (I305316,I2683,I304954,I304919,);
DFFARX1 I_17802 (I305308,I2683,I304954,I304937,);
nor I_17803 (I305361,I1030491,I1030482);
not I_17804 (I305378,I305361);
nor I_17805 (I304940,I305217,I305378);
nand I_17806 (I304925,I305234,I305378);
nor I_17807 (I304934,I304980,I305361);
DFFARX1 I_17808 (I305361,I2683,I304954,I304943,);
not I_17809 (I305481,I2690);
DFFARX1 I_17810 (I14253,I2683,I305481,I305507,);
nand I_17811 (I305515,I14277,I14256);
and I_17812 (I305532,I305515,I14253);
DFFARX1 I_17813 (I305532,I2683,I305481,I305558,);
nor I_17814 (I305449,I305558,I305507);
not I_17815 (I305580,I305558);
DFFARX1 I_17816 (I14259,I2683,I305481,I305606,);
nand I_17817 (I305614,I305606,I14268);
not I_17818 (I305631,I305614);
DFFARX1 I_17819 (I305631,I2683,I305481,I305657,);
not I_17820 (I305473,I305657);
nor I_17821 (I305679,I305507,I305614);
nor I_17822 (I305455,I305558,I305679);
DFFARX1 I_17823 (I14262,I2683,I305481,I305719,);
DFFARX1 I_17824 (I305719,I2683,I305481,I305736,);
not I_17825 (I305744,I305736);
not I_17826 (I305761,I305719);
nand I_17827 (I305458,I305761,I305580);
nand I_17828 (I305792,I14274,I14256);
and I_17829 (I305809,I305792,I14265);
DFFARX1 I_17830 (I305809,I2683,I305481,I305835,);
nor I_17831 (I305843,I305835,I305507);
DFFARX1 I_17832 (I305843,I2683,I305481,I305446,);
DFFARX1 I_17833 (I305835,I2683,I305481,I305464,);
nor I_17834 (I305888,I14271,I14256);
not I_17835 (I305905,I305888);
nor I_17836 (I305467,I305744,I305905);
nand I_17837 (I305452,I305761,I305905);
nor I_17838 (I305461,I305507,I305888);
DFFARX1 I_17839 (I305888,I2683,I305481,I305470,);
not I_17840 (I306008,I2690);
DFFARX1 I_17841 (I650719,I2683,I306008,I306034,);
nand I_17842 (I306042,I650722,I650716);
and I_17843 (I306059,I306042,I650728);
DFFARX1 I_17844 (I306059,I2683,I306008,I306085,);
nor I_17845 (I305976,I306085,I306034);
not I_17846 (I306107,I306085);
DFFARX1 I_17847 (I650731,I2683,I306008,I306133,);
nand I_17848 (I306141,I306133,I650722);
not I_17849 (I306158,I306141);
DFFARX1 I_17850 (I306158,I2683,I306008,I306184,);
not I_17851 (I306000,I306184);
nor I_17852 (I306206,I306034,I306141);
nor I_17853 (I305982,I306085,I306206);
DFFARX1 I_17854 (I650734,I2683,I306008,I306246,);
DFFARX1 I_17855 (I306246,I2683,I306008,I306263,);
not I_17856 (I306271,I306263);
not I_17857 (I306288,I306246);
nand I_17858 (I305985,I306288,I306107);
nand I_17859 (I306319,I650716,I650725);
and I_17860 (I306336,I306319,I650719);
DFFARX1 I_17861 (I306336,I2683,I306008,I306362,);
nor I_17862 (I306370,I306362,I306034);
DFFARX1 I_17863 (I306370,I2683,I306008,I305973,);
DFFARX1 I_17864 (I306362,I2683,I306008,I305991,);
nor I_17865 (I306415,I650737,I650725);
not I_17866 (I306432,I306415);
nor I_17867 (I305994,I306271,I306432);
nand I_17868 (I305979,I306288,I306432);
nor I_17869 (I305988,I306034,I306415);
DFFARX1 I_17870 (I306415,I2683,I306008,I305997,);
not I_17871 (I306535,I2690);
DFFARX1 I_17872 (I1029918,I2683,I306535,I306561,);
nand I_17873 (I306569,I1029945,I1029921);
and I_17874 (I306586,I306569,I1029930);
DFFARX1 I_17875 (I306586,I2683,I306535,I306612,);
nor I_17876 (I306503,I306612,I306561);
not I_17877 (I306634,I306612);
DFFARX1 I_17878 (I1029918,I2683,I306535,I306660,);
nand I_17879 (I306668,I306660,I1029942);
not I_17880 (I306685,I306668);
DFFARX1 I_17881 (I306685,I2683,I306535,I306711,);
not I_17882 (I306527,I306711);
nor I_17883 (I306733,I306561,I306668);
nor I_17884 (I306509,I306612,I306733);
DFFARX1 I_17885 (I1029924,I2683,I306535,I306773,);
DFFARX1 I_17886 (I306773,I2683,I306535,I306790,);
not I_17887 (I306798,I306790);
not I_17888 (I306815,I306773);
nand I_17889 (I306512,I306815,I306634);
nand I_17890 (I306846,I1029939,I1029927);
and I_17891 (I306863,I306846,I1029933);
DFFARX1 I_17892 (I306863,I2683,I306535,I306889,);
nor I_17893 (I306897,I306889,I306561);
DFFARX1 I_17894 (I306897,I2683,I306535,I306500,);
DFFARX1 I_17895 (I306889,I2683,I306535,I306518,);
nor I_17896 (I306942,I1029936,I1029927);
not I_17897 (I306959,I306942);
nor I_17898 (I306521,I306798,I306959);
nand I_17899 (I306506,I306815,I306959);
nor I_17900 (I306515,I306561,I306942);
DFFARX1 I_17901 (I306942,I2683,I306535,I306524,);
not I_17902 (I307062,I2690);
DFFARX1 I_17903 (I661786,I2683,I307062,I307088,);
nand I_17904 (I307096,I661789,I661783);
and I_17905 (I307113,I307096,I661795);
DFFARX1 I_17906 (I307113,I2683,I307062,I307139,);
nor I_17907 (I307030,I307139,I307088);
not I_17908 (I307161,I307139);
DFFARX1 I_17909 (I661798,I2683,I307062,I307187,);
nand I_17910 (I307195,I307187,I661789);
not I_17911 (I307212,I307195);
DFFARX1 I_17912 (I307212,I2683,I307062,I307238,);
not I_17913 (I307054,I307238);
nor I_17914 (I307260,I307088,I307195);
nor I_17915 (I307036,I307139,I307260);
DFFARX1 I_17916 (I661801,I2683,I307062,I307300,);
DFFARX1 I_17917 (I307300,I2683,I307062,I307317,);
not I_17918 (I307325,I307317);
not I_17919 (I307342,I307300);
nand I_17920 (I307039,I307342,I307161);
nand I_17921 (I307373,I661783,I661792);
and I_17922 (I307390,I307373,I661786);
DFFARX1 I_17923 (I307390,I2683,I307062,I307416,);
nor I_17924 (I307424,I307416,I307088);
DFFARX1 I_17925 (I307424,I2683,I307062,I307027,);
DFFARX1 I_17926 (I307416,I2683,I307062,I307045,);
nor I_17927 (I307469,I661804,I661792);
not I_17928 (I307486,I307469);
nor I_17929 (I307048,I307325,I307486);
nand I_17930 (I307033,I307342,I307486);
nor I_17931 (I307042,I307088,I307469);
DFFARX1 I_17932 (I307469,I2683,I307062,I307051,);
not I_17933 (I307589,I2690);
DFFARX1 I_17934 (I33752,I2683,I307589,I307615,);
nand I_17935 (I307623,I33776,I33755);
and I_17936 (I307640,I307623,I33752);
DFFARX1 I_17937 (I307640,I2683,I307589,I307666,);
nor I_17938 (I307557,I307666,I307615);
not I_17939 (I307688,I307666);
DFFARX1 I_17940 (I33758,I2683,I307589,I307714,);
nand I_17941 (I307722,I307714,I33767);
not I_17942 (I307739,I307722);
DFFARX1 I_17943 (I307739,I2683,I307589,I307765,);
not I_17944 (I307581,I307765);
nor I_17945 (I307787,I307615,I307722);
nor I_17946 (I307563,I307666,I307787);
DFFARX1 I_17947 (I33761,I2683,I307589,I307827,);
DFFARX1 I_17948 (I307827,I2683,I307589,I307844,);
not I_17949 (I307852,I307844);
not I_17950 (I307869,I307827);
nand I_17951 (I307566,I307869,I307688);
nand I_17952 (I307900,I33773,I33755);
and I_17953 (I307917,I307900,I33764);
DFFARX1 I_17954 (I307917,I2683,I307589,I307943,);
nor I_17955 (I307951,I307943,I307615);
DFFARX1 I_17956 (I307951,I2683,I307589,I307554,);
DFFARX1 I_17957 (I307943,I2683,I307589,I307572,);
nor I_17958 (I307996,I33770,I33755);
not I_17959 (I308013,I307996);
nor I_17960 (I307575,I307852,I308013);
nand I_17961 (I307560,I307869,I308013);
nor I_17962 (I307569,I307615,I307996);
DFFARX1 I_17963 (I307996,I2683,I307589,I307578,);
not I_17964 (I308116,I2690);
DFFARX1 I_17965 (I723224,I2683,I308116,I308142,);
nand I_17966 (I308150,I723221,I723239);
and I_17967 (I308167,I308150,I723230);
DFFARX1 I_17968 (I308167,I2683,I308116,I308193,);
nor I_17969 (I308084,I308193,I308142);
not I_17970 (I308215,I308193);
DFFARX1 I_17971 (I723245,I2683,I308116,I308241,);
nand I_17972 (I308249,I308241,I723227);
not I_17973 (I308266,I308249);
DFFARX1 I_17974 (I308266,I2683,I308116,I308292,);
not I_17975 (I308108,I308292);
nor I_17976 (I308314,I308142,I308249);
nor I_17977 (I308090,I308193,I308314);
DFFARX1 I_17978 (I723233,I2683,I308116,I308354,);
DFFARX1 I_17979 (I308354,I2683,I308116,I308371,);
not I_17980 (I308379,I308371);
not I_17981 (I308396,I308354);
nand I_17982 (I308093,I308396,I308215);
nand I_17983 (I308427,I723221,I723248);
and I_17984 (I308444,I308427,I723236);
DFFARX1 I_17985 (I308444,I2683,I308116,I308470,);
nor I_17986 (I308478,I308470,I308142);
DFFARX1 I_17987 (I308478,I2683,I308116,I308081,);
DFFARX1 I_17988 (I308470,I2683,I308116,I308099,);
nor I_17989 (I308523,I723242,I723248);
not I_17990 (I308540,I308523);
nor I_17991 (I308102,I308379,I308540);
nand I_17992 (I308087,I308396,I308540);
nor I_17993 (I308096,I308142,I308523);
DFFARX1 I_17994 (I308523,I2683,I308116,I308105,);
not I_17995 (I308643,I2690);
DFFARX1 I_17996 (I329054,I2683,I308643,I308669,);
nand I_17997 (I308677,I329066,I329045);
and I_17998 (I308694,I308677,I329069);
DFFARX1 I_17999 (I308694,I2683,I308643,I308720,);
nor I_18000 (I308611,I308720,I308669);
not I_18001 (I308742,I308720);
DFFARX1 I_18002 (I329060,I2683,I308643,I308768,);
nand I_18003 (I308776,I308768,I329042);
not I_18004 (I308793,I308776);
DFFARX1 I_18005 (I308793,I2683,I308643,I308819,);
not I_18006 (I308635,I308819);
nor I_18007 (I308841,I308669,I308776);
nor I_18008 (I308617,I308720,I308841);
DFFARX1 I_18009 (I329057,I2683,I308643,I308881,);
DFFARX1 I_18010 (I308881,I2683,I308643,I308898,);
not I_18011 (I308906,I308898);
not I_18012 (I308923,I308881);
nand I_18013 (I308620,I308923,I308742);
nand I_18014 (I308954,I329042,I329048);
and I_18015 (I308971,I308954,I329051);
DFFARX1 I_18016 (I308971,I2683,I308643,I308997,);
nor I_18017 (I309005,I308997,I308669);
DFFARX1 I_18018 (I309005,I2683,I308643,I308608,);
DFFARX1 I_18019 (I308997,I2683,I308643,I308626,);
nor I_18020 (I309050,I329063,I329048);
not I_18021 (I309067,I309050);
nor I_18022 (I308629,I308906,I309067);
nand I_18023 (I308614,I308923,I309067);
nor I_18024 (I308623,I308669,I309050);
DFFARX1 I_18025 (I309050,I2683,I308643,I308632,);
not I_18026 (I309170,I2690);
DFFARX1 I_18027 (I135480,I2683,I309170,I309196,);
nand I_18028 (I309204,I135480,I135486);
and I_18029 (I309221,I309204,I135504);
DFFARX1 I_18030 (I309221,I2683,I309170,I309247,);
nor I_18031 (I309138,I309247,I309196);
not I_18032 (I309269,I309247);
DFFARX1 I_18033 (I135492,I2683,I309170,I309295,);
nand I_18034 (I309303,I309295,I135489);
not I_18035 (I309320,I309303);
DFFARX1 I_18036 (I309320,I2683,I309170,I309346,);
not I_18037 (I309162,I309346);
nor I_18038 (I309368,I309196,I309303);
nor I_18039 (I309144,I309247,I309368);
DFFARX1 I_18040 (I135498,I2683,I309170,I309408,);
DFFARX1 I_18041 (I309408,I2683,I309170,I309425,);
not I_18042 (I309433,I309425);
not I_18043 (I309450,I309408);
nand I_18044 (I309147,I309450,I309269);
nand I_18045 (I309481,I135483,I135483);
and I_18046 (I309498,I309481,I135495);
DFFARX1 I_18047 (I309498,I2683,I309170,I309524,);
nor I_18048 (I309532,I309524,I309196);
DFFARX1 I_18049 (I309532,I2683,I309170,I309135,);
DFFARX1 I_18050 (I309524,I2683,I309170,I309153,);
nor I_18051 (I309577,I135501,I135483);
not I_18052 (I309594,I309577);
nor I_18053 (I309156,I309433,I309594);
nand I_18054 (I309141,I309450,I309594);
nor I_18055 (I309150,I309196,I309577);
DFFARX1 I_18056 (I309577,I2683,I309170,I309159,);
not I_18057 (I309697,I2690);
DFFARX1 I_18058 (I14780,I2683,I309697,I309723,);
nand I_18059 (I309731,I14804,I14783);
and I_18060 (I309748,I309731,I14780);
DFFARX1 I_18061 (I309748,I2683,I309697,I309774,);
nor I_18062 (I309665,I309774,I309723);
not I_18063 (I309796,I309774);
DFFARX1 I_18064 (I14786,I2683,I309697,I309822,);
nand I_18065 (I309830,I309822,I14795);
not I_18066 (I309847,I309830);
DFFARX1 I_18067 (I309847,I2683,I309697,I309873,);
not I_18068 (I309689,I309873);
nor I_18069 (I309895,I309723,I309830);
nor I_18070 (I309671,I309774,I309895);
DFFARX1 I_18071 (I14789,I2683,I309697,I309935,);
DFFARX1 I_18072 (I309935,I2683,I309697,I309952,);
not I_18073 (I309960,I309952);
not I_18074 (I309977,I309935);
nand I_18075 (I309674,I309977,I309796);
nand I_18076 (I310008,I14801,I14783);
and I_18077 (I310025,I310008,I14792);
DFFARX1 I_18078 (I310025,I2683,I309697,I310051,);
nor I_18079 (I310059,I310051,I309723);
DFFARX1 I_18080 (I310059,I2683,I309697,I309662,);
DFFARX1 I_18081 (I310051,I2683,I309697,I309680,);
nor I_18082 (I310104,I14798,I14783);
not I_18083 (I310121,I310104);
nor I_18084 (I309683,I309960,I310121);
nand I_18085 (I309668,I309977,I310121);
nor I_18086 (I309677,I309723,I310104);
DFFARX1 I_18087 (I310104,I2683,I309697,I309686,);
not I_18088 (I310224,I2690);
DFFARX1 I_18089 (I489639,I2683,I310224,I310250,);
nand I_18090 (I310258,I489624,I489627);
and I_18091 (I310275,I310258,I489642);
DFFARX1 I_18092 (I310275,I2683,I310224,I310301,);
nor I_18093 (I310192,I310301,I310250);
not I_18094 (I310323,I310301);
DFFARX1 I_18095 (I489636,I2683,I310224,I310349,);
nand I_18096 (I310357,I310349,I489627);
not I_18097 (I310374,I310357);
DFFARX1 I_18098 (I310374,I2683,I310224,I310400,);
not I_18099 (I310216,I310400);
nor I_18100 (I310422,I310250,I310357);
nor I_18101 (I310198,I310301,I310422);
DFFARX1 I_18102 (I489633,I2683,I310224,I310462,);
DFFARX1 I_18103 (I310462,I2683,I310224,I310479,);
not I_18104 (I310487,I310479);
not I_18105 (I310504,I310462);
nand I_18106 (I310201,I310504,I310323);
nand I_18107 (I310535,I489648,I489624);
and I_18108 (I310552,I310535,I489645);
DFFARX1 I_18109 (I310552,I2683,I310224,I310578,);
nor I_18110 (I310586,I310578,I310250);
DFFARX1 I_18111 (I310586,I2683,I310224,I310189,);
DFFARX1 I_18112 (I310578,I2683,I310224,I310207,);
nor I_18113 (I310631,I489630,I489624);
not I_18114 (I310648,I310631);
nor I_18115 (I310210,I310487,I310648);
nand I_18116 (I310195,I310504,I310648);
nor I_18117 (I310204,I310250,I310631);
DFFARX1 I_18118 (I310631,I2683,I310224,I310213,);
not I_18119 (I310751,I2690);
DFFARX1 I_18120 (I965744,I2683,I310751,I310777,);
nand I_18121 (I310785,I965726,I965750);
and I_18122 (I310802,I310785,I965741);
DFFARX1 I_18123 (I310802,I2683,I310751,I310828,);
nor I_18124 (I310719,I310828,I310777);
not I_18125 (I310850,I310828);
DFFARX1 I_18126 (I965747,I2683,I310751,I310876,);
nand I_18127 (I310884,I310876,I965735);
not I_18128 (I310901,I310884);
DFFARX1 I_18129 (I310901,I2683,I310751,I310927,);
not I_18130 (I310743,I310927);
nor I_18131 (I310949,I310777,I310884);
nor I_18132 (I310725,I310828,I310949);
DFFARX1 I_18133 (I965726,I2683,I310751,I310989,);
DFFARX1 I_18134 (I310989,I2683,I310751,I311006,);
not I_18135 (I311014,I311006);
not I_18136 (I311031,I310989);
nand I_18137 (I310728,I311031,I310850);
nand I_18138 (I311062,I965732,I965729);
and I_18139 (I311079,I311062,I965738);
DFFARX1 I_18140 (I311079,I2683,I310751,I311105,);
nor I_18141 (I311113,I311105,I310777);
DFFARX1 I_18142 (I311113,I2683,I310751,I310716,);
DFFARX1 I_18143 (I311105,I2683,I310751,I310734,);
nor I_18144 (I311158,I965729,I965729);
not I_18145 (I311175,I311158);
nor I_18146 (I310737,I311014,I311175);
nand I_18147 (I310722,I311031,I311175);
nor I_18148 (I310731,I310777,I311158);
DFFARX1 I_18149 (I311158,I2683,I310751,I310740,);
not I_18150 (I311278,I2690);
DFFARX1 I_18151 (I988589,I2683,I311278,I311304,);
nand I_18152 (I311312,I988586,I988577);
and I_18153 (I311329,I311312,I988574);
DFFARX1 I_18154 (I311329,I2683,I311278,I311355,);
nor I_18155 (I311246,I311355,I311304);
not I_18156 (I311377,I311355);
DFFARX1 I_18157 (I988583,I2683,I311278,I311403,);
nand I_18158 (I311411,I311403,I988592);
not I_18159 (I311428,I311411);
DFFARX1 I_18160 (I311428,I2683,I311278,I311454,);
not I_18161 (I311270,I311454);
nor I_18162 (I311476,I311304,I311411);
nor I_18163 (I311252,I311355,I311476);
DFFARX1 I_18164 (I988595,I2683,I311278,I311516,);
DFFARX1 I_18165 (I311516,I2683,I311278,I311533,);
not I_18166 (I311541,I311533);
not I_18167 (I311558,I311516);
nand I_18168 (I311255,I311558,I311377);
nand I_18169 (I311589,I988574,I988580);
and I_18170 (I311606,I311589,I988598);
DFFARX1 I_18171 (I311606,I2683,I311278,I311632,);
nor I_18172 (I311640,I311632,I311304);
DFFARX1 I_18173 (I311640,I2683,I311278,I311243,);
DFFARX1 I_18174 (I311632,I2683,I311278,I311261,);
nor I_18175 (I311685,I988577,I988580);
not I_18176 (I311702,I311685);
nor I_18177 (I311264,I311541,I311702);
nand I_18178 (I311249,I311558,I311702);
nor I_18179 (I311258,I311304,I311685);
DFFARX1 I_18180 (I311685,I2683,I311278,I311267,);
not I_18181 (I311805,I2690);
DFFARX1 I_18182 (I637544,I2683,I311805,I311831,);
nand I_18183 (I311839,I637547,I637541);
and I_18184 (I311856,I311839,I637553);
DFFARX1 I_18185 (I311856,I2683,I311805,I311882,);
nor I_18186 (I311773,I311882,I311831);
not I_18187 (I311904,I311882);
DFFARX1 I_18188 (I637556,I2683,I311805,I311930,);
nand I_18189 (I311938,I311930,I637547);
not I_18190 (I311955,I311938);
DFFARX1 I_18191 (I311955,I2683,I311805,I311981,);
not I_18192 (I311797,I311981);
nor I_18193 (I312003,I311831,I311938);
nor I_18194 (I311779,I311882,I312003);
DFFARX1 I_18195 (I637559,I2683,I311805,I312043,);
DFFARX1 I_18196 (I312043,I2683,I311805,I312060,);
not I_18197 (I312068,I312060);
not I_18198 (I312085,I312043);
nand I_18199 (I311782,I312085,I311904);
nand I_18200 (I312116,I637541,I637550);
and I_18201 (I312133,I312116,I637544);
DFFARX1 I_18202 (I312133,I2683,I311805,I312159,);
nor I_18203 (I312167,I312159,I311831);
DFFARX1 I_18204 (I312167,I2683,I311805,I311770,);
DFFARX1 I_18205 (I312159,I2683,I311805,I311788,);
nor I_18206 (I312212,I637562,I637550);
not I_18207 (I312229,I312212);
nor I_18208 (I311791,I312068,I312229);
nand I_18209 (I311776,I312085,I312229);
nor I_18210 (I311785,I311831,I312212);
DFFARX1 I_18211 (I312212,I2683,I311805,I311794,);
not I_18212 (I312332,I2690);
DFFARX1 I_18213 (I1096545,I2683,I312332,I312358,);
nand I_18214 (I312366,I1096524,I1096524);
and I_18215 (I312383,I312366,I1096551);
DFFARX1 I_18216 (I312383,I2683,I312332,I312409,);
nor I_18217 (I312300,I312409,I312358);
not I_18218 (I312431,I312409);
DFFARX1 I_18219 (I1096539,I2683,I312332,I312457,);
nand I_18220 (I312465,I312457,I1096542);
not I_18221 (I312482,I312465);
DFFARX1 I_18222 (I312482,I2683,I312332,I312508,);
not I_18223 (I312324,I312508);
nor I_18224 (I312530,I312358,I312465);
nor I_18225 (I312306,I312409,I312530);
DFFARX1 I_18226 (I1096533,I2683,I312332,I312570,);
DFFARX1 I_18227 (I312570,I2683,I312332,I312587,);
not I_18228 (I312595,I312587);
not I_18229 (I312612,I312570);
nand I_18230 (I312309,I312612,I312431);
nand I_18231 (I312643,I1096530,I1096527);
and I_18232 (I312660,I312643,I1096548);
DFFARX1 I_18233 (I312660,I2683,I312332,I312686,);
nor I_18234 (I312694,I312686,I312358);
DFFARX1 I_18235 (I312694,I2683,I312332,I312297,);
DFFARX1 I_18236 (I312686,I2683,I312332,I312315,);
nor I_18237 (I312739,I1096536,I1096527);
not I_18238 (I312756,I312739);
nor I_18239 (I312318,I312595,I312756);
nand I_18240 (I312303,I312612,I312756);
nor I_18241 (I312312,I312358,I312739);
DFFARX1 I_18242 (I312739,I2683,I312332,I312321,);
not I_18243 (I312859,I2690);
DFFARX1 I_18244 (I446867,I2683,I312859,I312885,);
nand I_18245 (I312893,I446852,I446855);
and I_18246 (I312910,I312893,I446870);
DFFARX1 I_18247 (I312910,I2683,I312859,I312936,);
nor I_18248 (I312827,I312936,I312885);
not I_18249 (I312958,I312936);
DFFARX1 I_18250 (I446864,I2683,I312859,I312984,);
nand I_18251 (I312992,I312984,I446855);
not I_18252 (I313009,I312992);
DFFARX1 I_18253 (I313009,I2683,I312859,I313035,);
not I_18254 (I312851,I313035);
nor I_18255 (I313057,I312885,I312992);
nor I_18256 (I312833,I312936,I313057);
DFFARX1 I_18257 (I446861,I2683,I312859,I313097,);
DFFARX1 I_18258 (I313097,I2683,I312859,I313114,);
not I_18259 (I313122,I313114);
not I_18260 (I313139,I313097);
nand I_18261 (I312836,I313139,I312958);
nand I_18262 (I313170,I446876,I446852);
and I_18263 (I313187,I313170,I446873);
DFFARX1 I_18264 (I313187,I2683,I312859,I313213,);
nor I_18265 (I313221,I313213,I312885);
DFFARX1 I_18266 (I313221,I2683,I312859,I312824,);
DFFARX1 I_18267 (I313213,I2683,I312859,I312842,);
nor I_18268 (I313266,I446858,I446852);
not I_18269 (I313283,I313266);
nor I_18270 (I312845,I313122,I313283);
nand I_18271 (I312830,I313139,I313283);
nor I_18272 (I312839,I312885,I313266);
DFFARX1 I_18273 (I313266,I2683,I312859,I312848,);
not I_18274 (I313386,I2690);
DFFARX1 I_18275 (I32698,I2683,I313386,I313412,);
nand I_18276 (I313420,I32722,I32701);
and I_18277 (I313437,I313420,I32698);
DFFARX1 I_18278 (I313437,I2683,I313386,I313463,);
nor I_18279 (I313354,I313463,I313412);
not I_18280 (I313485,I313463);
DFFARX1 I_18281 (I32704,I2683,I313386,I313511,);
nand I_18282 (I313519,I313511,I32713);
not I_18283 (I313536,I313519);
DFFARX1 I_18284 (I313536,I2683,I313386,I313562,);
not I_18285 (I313378,I313562);
nor I_18286 (I313584,I313412,I313519);
nor I_18287 (I313360,I313463,I313584);
DFFARX1 I_18288 (I32707,I2683,I313386,I313624,);
DFFARX1 I_18289 (I313624,I2683,I313386,I313641,);
not I_18290 (I313649,I313641);
not I_18291 (I313666,I313624);
nand I_18292 (I313363,I313666,I313485);
nand I_18293 (I313697,I32719,I32701);
and I_18294 (I313714,I313697,I32710);
DFFARX1 I_18295 (I313714,I2683,I313386,I313740,);
nor I_18296 (I313748,I313740,I313412);
DFFARX1 I_18297 (I313748,I2683,I313386,I313351,);
DFFARX1 I_18298 (I313740,I2683,I313386,I313369,);
nor I_18299 (I313793,I32716,I32701);
not I_18300 (I313810,I313793);
nor I_18301 (I313372,I313649,I313810);
nand I_18302 (I313357,I313666,I313810);
nor I_18303 (I313366,I313412,I313793);
DFFARX1 I_18304 (I313793,I2683,I313386,I313375,);
not I_18305 (I313913,I2690);
DFFARX1 I_18306 (I1066795,I2683,I313913,I313939,);
nand I_18307 (I313947,I1066774,I1066774);
and I_18308 (I313964,I313947,I1066801);
DFFARX1 I_18309 (I313964,I2683,I313913,I313990,);
nor I_18310 (I313881,I313990,I313939);
not I_18311 (I314012,I313990);
DFFARX1 I_18312 (I1066789,I2683,I313913,I314038,);
nand I_18313 (I314046,I314038,I1066792);
not I_18314 (I314063,I314046);
DFFARX1 I_18315 (I314063,I2683,I313913,I314089,);
not I_18316 (I313905,I314089);
nor I_18317 (I314111,I313939,I314046);
nor I_18318 (I313887,I313990,I314111);
DFFARX1 I_18319 (I1066783,I2683,I313913,I314151,);
DFFARX1 I_18320 (I314151,I2683,I313913,I314168,);
not I_18321 (I314176,I314168);
not I_18322 (I314193,I314151);
nand I_18323 (I313890,I314193,I314012);
nand I_18324 (I314224,I1066780,I1066777);
and I_18325 (I314241,I314224,I1066798);
DFFARX1 I_18326 (I314241,I2683,I313913,I314267,);
nor I_18327 (I314275,I314267,I313939);
DFFARX1 I_18328 (I314275,I2683,I313913,I313878,);
DFFARX1 I_18329 (I314267,I2683,I313913,I313896,);
nor I_18330 (I314320,I1066786,I1066777);
not I_18331 (I314337,I314320);
nor I_18332 (I313899,I314176,I314337);
nand I_18333 (I313884,I314193,I314337);
nor I_18334 (I313893,I313939,I314320);
DFFARX1 I_18335 (I314320,I2683,I313913,I313902,);
not I_18336 (I314440,I2690);
DFFARX1 I_18337 (I473455,I2683,I314440,I314466,);
nand I_18338 (I314474,I473440,I473443);
and I_18339 (I314491,I314474,I473458);
DFFARX1 I_18340 (I314491,I2683,I314440,I314517,);
nor I_18341 (I314408,I314517,I314466);
not I_18342 (I314539,I314517);
DFFARX1 I_18343 (I473452,I2683,I314440,I314565,);
nand I_18344 (I314573,I314565,I473443);
not I_18345 (I314590,I314573);
DFFARX1 I_18346 (I314590,I2683,I314440,I314616,);
not I_18347 (I314432,I314616);
nor I_18348 (I314638,I314466,I314573);
nor I_18349 (I314414,I314517,I314638);
DFFARX1 I_18350 (I473449,I2683,I314440,I314678,);
DFFARX1 I_18351 (I314678,I2683,I314440,I314695,);
not I_18352 (I314703,I314695);
not I_18353 (I314720,I314678);
nand I_18354 (I314417,I314720,I314539);
nand I_18355 (I314751,I473464,I473440);
and I_18356 (I314768,I314751,I473461);
DFFARX1 I_18357 (I314768,I2683,I314440,I314794,);
nor I_18358 (I314802,I314794,I314466);
DFFARX1 I_18359 (I314802,I2683,I314440,I314405,);
DFFARX1 I_18360 (I314794,I2683,I314440,I314423,);
nor I_18361 (I314847,I473446,I473440);
not I_18362 (I314864,I314847);
nor I_18363 (I314426,I314703,I314864);
nand I_18364 (I314411,I314720,I314864);
nor I_18365 (I314420,I314466,I314847);
DFFARX1 I_18366 (I314847,I2683,I314440,I314429,);
not I_18367 (I314967,I2690);
DFFARX1 I_18368 (I17415,I2683,I314967,I314993,);
nand I_18369 (I315001,I17439,I17418);
and I_18370 (I315018,I315001,I17415);
DFFARX1 I_18371 (I315018,I2683,I314967,I315044,);
nor I_18372 (I314935,I315044,I314993);
not I_18373 (I315066,I315044);
DFFARX1 I_18374 (I17421,I2683,I314967,I315092,);
nand I_18375 (I315100,I315092,I17430);
not I_18376 (I315117,I315100);
DFFARX1 I_18377 (I315117,I2683,I314967,I315143,);
not I_18378 (I314959,I315143);
nor I_18379 (I315165,I314993,I315100);
nor I_18380 (I314941,I315044,I315165);
DFFARX1 I_18381 (I17424,I2683,I314967,I315205,);
DFFARX1 I_18382 (I315205,I2683,I314967,I315222,);
not I_18383 (I315230,I315222);
not I_18384 (I315247,I315205);
nand I_18385 (I314944,I315247,I315066);
nand I_18386 (I315278,I17436,I17418);
and I_18387 (I315295,I315278,I17427);
DFFARX1 I_18388 (I315295,I2683,I314967,I315321,);
nor I_18389 (I315329,I315321,I314993);
DFFARX1 I_18390 (I315329,I2683,I314967,I314932,);
DFFARX1 I_18391 (I315321,I2683,I314967,I314950,);
nor I_18392 (I315374,I17433,I17418);
not I_18393 (I315391,I315374);
nor I_18394 (I314953,I315230,I315391);
nand I_18395 (I314938,I315247,I315391);
nor I_18396 (I314947,I314993,I315374);
DFFARX1 I_18397 (I315374,I2683,I314967,I314956,);
not I_18398 (I315494,I2690);
DFFARX1 I_18399 (I123580,I2683,I315494,I315520,);
nand I_18400 (I315528,I123580,I123586);
and I_18401 (I315545,I315528,I123604);
DFFARX1 I_18402 (I315545,I2683,I315494,I315571,);
nor I_18403 (I315462,I315571,I315520);
not I_18404 (I315593,I315571);
DFFARX1 I_18405 (I123592,I2683,I315494,I315619,);
nand I_18406 (I315627,I315619,I123589);
not I_18407 (I315644,I315627);
DFFARX1 I_18408 (I315644,I2683,I315494,I315670,);
not I_18409 (I315486,I315670);
nor I_18410 (I315692,I315520,I315627);
nor I_18411 (I315468,I315571,I315692);
DFFARX1 I_18412 (I123598,I2683,I315494,I315732,);
DFFARX1 I_18413 (I315732,I2683,I315494,I315749,);
not I_18414 (I315757,I315749);
not I_18415 (I315774,I315732);
nand I_18416 (I315471,I315774,I315593);
nand I_18417 (I315805,I123583,I123583);
and I_18418 (I315822,I315805,I123595);
DFFARX1 I_18419 (I315822,I2683,I315494,I315848,);
nor I_18420 (I315856,I315848,I315520);
DFFARX1 I_18421 (I315856,I2683,I315494,I315459,);
DFFARX1 I_18422 (I315848,I2683,I315494,I315477,);
nor I_18423 (I315901,I123601,I123583);
not I_18424 (I315918,I315901);
nor I_18425 (I315480,I315757,I315918);
nand I_18426 (I315465,I315774,I315918);
nor I_18427 (I315474,I315520,I315901);
DFFARX1 I_18428 (I315901,I2683,I315494,I315483,);
not I_18429 (I316021,I2690);
DFFARX1 I_18430 (I395515,I2683,I316021,I316047,);
DFFARX1 I_18431 (I316047,I2683,I316021,I316064,);
not I_18432 (I316013,I316064);
not I_18433 (I316086,I316047);
nand I_18434 (I316103,I395518,I395536);
and I_18435 (I316120,I316103,I395524);
DFFARX1 I_18436 (I316120,I2683,I316021,I316146,);
not I_18437 (I316154,I316146);
DFFARX1 I_18438 (I395515,I2683,I316021,I316180,);
and I_18439 (I316188,I316180,I395533);
nand I_18440 (I316205,I316180,I395533);
nand I_18441 (I315992,I316154,I316205);
DFFARX1 I_18442 (I395527,I2683,I316021,I316245,);
nor I_18443 (I316253,I316245,I316188);
DFFARX1 I_18444 (I316253,I2683,I316021,I315986,);
nor I_18445 (I316001,I316245,I316146);
nand I_18446 (I316298,I395530,I395512);
and I_18447 (I316315,I316298,I395521);
DFFARX1 I_18448 (I316315,I2683,I316021,I316341,);
nor I_18449 (I315989,I316341,I316245);
not I_18450 (I316363,I316341);
nor I_18451 (I316380,I316363,I316154);
nor I_18452 (I316397,I316086,I316380);
DFFARX1 I_18453 (I316397,I2683,I316021,I316004,);
nor I_18454 (I316428,I316363,I316245);
nor I_18455 (I316445,I395512,I395512);
nor I_18456 (I315995,I316445,I316428);
not I_18457 (I316476,I316445);
nand I_18458 (I315998,I316205,I316476);
DFFARX1 I_18459 (I316445,I2683,I316021,I316010,);
DFFARX1 I_18460 (I316445,I2683,I316021,I316007,);
not I_18461 (I316565,I2690);
DFFARX1 I_18462 (I673916,I2683,I316565,I316591,);
DFFARX1 I_18463 (I316591,I2683,I316565,I316608,);
not I_18464 (I316557,I316608);
not I_18465 (I316630,I316591);
nand I_18466 (I316647,I673910,I673907);
and I_18467 (I316664,I316647,I673922);
DFFARX1 I_18468 (I316664,I2683,I316565,I316690,);
not I_18469 (I316698,I316690);
DFFARX1 I_18470 (I673910,I2683,I316565,I316724,);
and I_18471 (I316732,I316724,I673904);
nand I_18472 (I316749,I316724,I673904);
nand I_18473 (I316536,I316698,I316749);
DFFARX1 I_18474 (I673904,I2683,I316565,I316789,);
nor I_18475 (I316797,I316789,I316732);
DFFARX1 I_18476 (I316797,I2683,I316565,I316530,);
nor I_18477 (I316545,I316789,I316690);
nand I_18478 (I316842,I673919,I673913);
and I_18479 (I316859,I316842,I673907);
DFFARX1 I_18480 (I316859,I2683,I316565,I316885,);
nor I_18481 (I316533,I316885,I316789);
not I_18482 (I316907,I316885);
nor I_18483 (I316924,I316907,I316698);
nor I_18484 (I316941,I316630,I316924);
DFFARX1 I_18485 (I316941,I2683,I316565,I316548,);
nor I_18486 (I316972,I316907,I316789);
nor I_18487 (I316989,I673925,I673913);
nor I_18488 (I316539,I316989,I316972);
not I_18489 (I317020,I316989);
nand I_18490 (I316542,I316749,I317020);
DFFARX1 I_18491 (I316989,I2683,I316565,I316554,);
DFFARX1 I_18492 (I316989,I2683,I316565,I316551,);
not I_18493 (I317109,I2690);
DFFARX1 I_18494 (I432983,I2683,I317109,I317135,);
DFFARX1 I_18495 (I317135,I2683,I317109,I317152,);
not I_18496 (I317101,I317152);
not I_18497 (I317174,I317135);
nand I_18498 (I317191,I432980,I433001);
and I_18499 (I317208,I317191,I433004);
DFFARX1 I_18500 (I317208,I2683,I317109,I317234,);
not I_18501 (I317242,I317234);
DFFARX1 I_18502 (I432989,I2683,I317109,I317268,);
and I_18503 (I317276,I317268,I432992);
nand I_18504 (I317293,I317268,I432992);
nand I_18505 (I317080,I317242,I317293);
DFFARX1 I_18506 (I432995,I2683,I317109,I317333,);
nor I_18507 (I317341,I317333,I317276);
DFFARX1 I_18508 (I317341,I2683,I317109,I317074,);
nor I_18509 (I317089,I317333,I317234);
nand I_18510 (I317386,I432980,I432986);
and I_18511 (I317403,I317386,I432998);
DFFARX1 I_18512 (I317403,I2683,I317109,I317429,);
nor I_18513 (I317077,I317429,I317333);
not I_18514 (I317451,I317429);
nor I_18515 (I317468,I317451,I317242);
nor I_18516 (I317485,I317174,I317468);
DFFARX1 I_18517 (I317485,I2683,I317109,I317092,);
nor I_18518 (I317516,I317451,I317333);
nor I_18519 (I317533,I432983,I432986);
nor I_18520 (I317083,I317533,I317516);
not I_18521 (I317564,I317533);
nand I_18522 (I317086,I317293,I317564);
DFFARX1 I_18523 (I317533,I2683,I317109,I317098,);
DFFARX1 I_18524 (I317533,I2683,I317109,I317095,);
not I_18525 (I317653,I2690);
DFFARX1 I_18526 (I981505,I2683,I317653,I317679,);
DFFARX1 I_18527 (I317679,I2683,I317653,I317696,);
not I_18528 (I317645,I317696);
not I_18529 (I317718,I317679);
nand I_18530 (I317735,I981517,I981520);
and I_18531 (I317752,I317735,I981523);
DFFARX1 I_18532 (I317752,I2683,I317653,I317778,);
not I_18533 (I317786,I317778);
DFFARX1 I_18534 (I981508,I2683,I317653,I317812,);
and I_18535 (I317820,I317812,I981514);
nand I_18536 (I317837,I317812,I981514);
nand I_18537 (I317624,I317786,I317837);
DFFARX1 I_18538 (I981502,I2683,I317653,I317877,);
nor I_18539 (I317885,I317877,I317820);
DFFARX1 I_18540 (I317885,I2683,I317653,I317618,);
nor I_18541 (I317633,I317877,I317778);
nand I_18542 (I317930,I981505,I981526);
and I_18543 (I317947,I317930,I981511);
DFFARX1 I_18544 (I317947,I2683,I317653,I317973,);
nor I_18545 (I317621,I317973,I317877);
not I_18546 (I317995,I317973);
nor I_18547 (I318012,I317995,I317786);
nor I_18548 (I318029,I317718,I318012);
DFFARX1 I_18549 (I318029,I2683,I317653,I317636,);
nor I_18550 (I318060,I317995,I317877);
nor I_18551 (I318077,I981502,I981526);
nor I_18552 (I317627,I318077,I318060);
not I_18553 (I318108,I318077);
nand I_18554 (I317630,I317837,I318108);
DFFARX1 I_18555 (I318077,I2683,I317653,I317642,);
DFFARX1 I_18556 (I318077,I2683,I317653,I317639,);
not I_18557 (I318197,I2690);
DFFARX1 I_18558 (I998418,I2683,I318197,I318223,);
DFFARX1 I_18559 (I318223,I2683,I318197,I318240,);
not I_18560 (I318189,I318240);
not I_18561 (I318262,I318223);
nand I_18562 (I318279,I998415,I998412);
and I_18563 (I318296,I318279,I998400);
DFFARX1 I_18564 (I318296,I2683,I318197,I318322,);
not I_18565 (I318330,I318322);
DFFARX1 I_18566 (I998424,I2683,I318197,I318356,);
and I_18567 (I318364,I318356,I998409);
nand I_18568 (I318381,I318356,I998409);
nand I_18569 (I318168,I318330,I318381);
DFFARX1 I_18570 (I998403,I2683,I318197,I318421,);
nor I_18571 (I318429,I318421,I318364);
DFFARX1 I_18572 (I318429,I2683,I318197,I318162,);
nor I_18573 (I318177,I318421,I318322);
nand I_18574 (I318474,I998400,I998406);
and I_18575 (I318491,I318474,I998421);
DFFARX1 I_18576 (I318491,I2683,I318197,I318517,);
nor I_18577 (I318165,I318517,I318421);
not I_18578 (I318539,I318517);
nor I_18579 (I318556,I318539,I318330);
nor I_18580 (I318573,I318262,I318556);
DFFARX1 I_18581 (I318573,I2683,I318197,I318180,);
nor I_18582 (I318604,I318539,I318421);
nor I_18583 (I318621,I998403,I998406);
nor I_18584 (I318171,I318621,I318604);
not I_18585 (I318652,I318621);
nand I_18586 (I318174,I318381,I318652);
DFFARX1 I_18587 (I318621,I2683,I318197,I318186,);
DFFARX1 I_18588 (I318621,I2683,I318197,I318183,);
not I_18589 (I318741,I2690);
DFFARX1 I_18590 (I207484,I2683,I318741,I318767,);
DFFARX1 I_18591 (I318767,I2683,I318741,I318784,);
not I_18592 (I318733,I318784);
not I_18593 (I318806,I318767);
nand I_18594 (I318823,I207496,I207475);
and I_18595 (I318840,I318823,I207478);
DFFARX1 I_18596 (I318840,I2683,I318741,I318866,);
not I_18597 (I318874,I318866);
DFFARX1 I_18598 (I207487,I2683,I318741,I318900,);
and I_18599 (I318908,I318900,I207499);
nand I_18600 (I318925,I318900,I207499);
nand I_18601 (I318712,I318874,I318925);
DFFARX1 I_18602 (I207493,I2683,I318741,I318965,);
nor I_18603 (I318973,I318965,I318908);
DFFARX1 I_18604 (I318973,I2683,I318741,I318706,);
nor I_18605 (I318721,I318965,I318866);
nand I_18606 (I319018,I207481,I207478);
and I_18607 (I319035,I319018,I207490);
DFFARX1 I_18608 (I319035,I2683,I318741,I319061,);
nor I_18609 (I318709,I319061,I318965);
not I_18610 (I319083,I319061);
nor I_18611 (I319100,I319083,I318874);
nor I_18612 (I319117,I318806,I319100);
DFFARX1 I_18613 (I319117,I2683,I318741,I318724,);
nor I_18614 (I319148,I319083,I318965);
nor I_18615 (I319165,I207475,I207478);
nor I_18616 (I318715,I319165,I319148);
not I_18617 (I319196,I319165);
nand I_18618 (I318718,I318925,I319196);
DFFARX1 I_18619 (I319165,I2683,I318741,I318730,);
DFFARX1 I_18620 (I319165,I2683,I318741,I318727,);
not I_18621 (I319285,I2690);
DFFARX1 I_18622 (I709661,I2683,I319285,I319311,);
DFFARX1 I_18623 (I319311,I2683,I319285,I319328,);
not I_18624 (I319277,I319328);
not I_18625 (I319350,I319311);
nand I_18626 (I319367,I709676,I709664);
and I_18627 (I319384,I319367,I709655);
DFFARX1 I_18628 (I319384,I2683,I319285,I319410,);
not I_18629 (I319418,I319410);
DFFARX1 I_18630 (I709667,I2683,I319285,I319444,);
and I_18631 (I319452,I319444,I709658);
nand I_18632 (I319469,I319444,I709658);
nand I_18633 (I319256,I319418,I319469);
DFFARX1 I_18634 (I709673,I2683,I319285,I319509,);
nor I_18635 (I319517,I319509,I319452);
DFFARX1 I_18636 (I319517,I2683,I319285,I319250,);
nor I_18637 (I319265,I319509,I319410);
nand I_18638 (I319562,I709682,I709670);
and I_18639 (I319579,I319562,I709679);
DFFARX1 I_18640 (I319579,I2683,I319285,I319605,);
nor I_18641 (I319253,I319605,I319509);
not I_18642 (I319627,I319605);
nor I_18643 (I319644,I319627,I319418);
nor I_18644 (I319661,I319350,I319644);
DFFARX1 I_18645 (I319661,I2683,I319285,I319268,);
nor I_18646 (I319692,I319627,I319509);
nor I_18647 (I319709,I709655,I709670);
nor I_18648 (I319259,I319709,I319692);
not I_18649 (I319740,I319709);
nand I_18650 (I319262,I319469,I319740);
DFFARX1 I_18651 (I319709,I2683,I319285,I319274,);
DFFARX1 I_18652 (I319709,I2683,I319285,I319271,);
not I_18653 (I319829,I2690);
DFFARX1 I_18654 (I394325,I2683,I319829,I319855,);
DFFARX1 I_18655 (I319855,I2683,I319829,I319872,);
not I_18656 (I319821,I319872);
not I_18657 (I319894,I319855);
nand I_18658 (I319911,I394328,I394346);
and I_18659 (I319928,I319911,I394334);
DFFARX1 I_18660 (I319928,I2683,I319829,I319954,);
not I_18661 (I319962,I319954);
DFFARX1 I_18662 (I394325,I2683,I319829,I319988,);
and I_18663 (I319996,I319988,I394343);
nand I_18664 (I320013,I319988,I394343);
nand I_18665 (I319800,I319962,I320013);
DFFARX1 I_18666 (I394337,I2683,I319829,I320053,);
nor I_18667 (I320061,I320053,I319996);
DFFARX1 I_18668 (I320061,I2683,I319829,I319794,);
nor I_18669 (I319809,I320053,I319954);
nand I_18670 (I320106,I394340,I394322);
and I_18671 (I320123,I320106,I394331);
DFFARX1 I_18672 (I320123,I2683,I319829,I320149,);
nor I_18673 (I319797,I320149,I320053);
not I_18674 (I320171,I320149);
nor I_18675 (I320188,I320171,I319962);
nor I_18676 (I320205,I319894,I320188);
DFFARX1 I_18677 (I320205,I2683,I319829,I319812,);
nor I_18678 (I320236,I320171,I320053);
nor I_18679 (I320253,I394322,I394322);
nor I_18680 (I319803,I320253,I320236);
not I_18681 (I320284,I320253);
nand I_18682 (I319806,I320013,I320284);
DFFARX1 I_18683 (I320253,I2683,I319829,I319818,);
DFFARX1 I_18684 (I320253,I2683,I319829,I319815,);
not I_18685 (I320373,I2690);
DFFARX1 I_18686 (I150959,I2683,I320373,I320399,);
DFFARX1 I_18687 (I320399,I2683,I320373,I320416,);
not I_18688 (I320365,I320416);
not I_18689 (I320438,I320399);
nand I_18690 (I320455,I150971,I150950);
and I_18691 (I320472,I320455,I150953);
DFFARX1 I_18692 (I320472,I2683,I320373,I320498,);
not I_18693 (I320506,I320498);
DFFARX1 I_18694 (I150962,I2683,I320373,I320532,);
and I_18695 (I320540,I320532,I150974);
nand I_18696 (I320557,I320532,I150974);
nand I_18697 (I320344,I320506,I320557);
DFFARX1 I_18698 (I150968,I2683,I320373,I320597,);
nor I_18699 (I320605,I320597,I320540);
DFFARX1 I_18700 (I320605,I2683,I320373,I320338,);
nor I_18701 (I320353,I320597,I320498);
nand I_18702 (I320650,I150956,I150953);
and I_18703 (I320667,I320650,I150965);
DFFARX1 I_18704 (I320667,I2683,I320373,I320693,);
nor I_18705 (I320341,I320693,I320597);
not I_18706 (I320715,I320693);
nor I_18707 (I320732,I320715,I320506);
nor I_18708 (I320749,I320438,I320732);
DFFARX1 I_18709 (I320749,I2683,I320373,I320356,);
nor I_18710 (I320780,I320715,I320597);
nor I_18711 (I320797,I150950,I150953);
nor I_18712 (I320347,I320797,I320780);
not I_18713 (I320828,I320797);
nand I_18714 (I320350,I320557,I320828);
DFFARX1 I_18715 (I320797,I2683,I320373,I320362,);
DFFARX1 I_18716 (I320797,I2683,I320373,I320359,);
not I_18717 (I320917,I2690);
DFFARX1 I_18718 (I724519,I2683,I320917,I320943,);
DFFARX1 I_18719 (I320943,I2683,I320917,I320960,);
not I_18720 (I320909,I320960);
not I_18721 (I320982,I320943);
nand I_18722 (I320999,I724534,I724522);
and I_18723 (I321016,I320999,I724513);
DFFARX1 I_18724 (I321016,I2683,I320917,I321042,);
not I_18725 (I321050,I321042);
DFFARX1 I_18726 (I724525,I2683,I320917,I321076,);
and I_18727 (I321084,I321076,I724516);
nand I_18728 (I321101,I321076,I724516);
nand I_18729 (I320888,I321050,I321101);
DFFARX1 I_18730 (I724531,I2683,I320917,I321141,);
nor I_18731 (I321149,I321141,I321084);
DFFARX1 I_18732 (I321149,I2683,I320917,I320882,);
nor I_18733 (I320897,I321141,I321042);
nand I_18734 (I321194,I724540,I724528);
and I_18735 (I321211,I321194,I724537);
DFFARX1 I_18736 (I321211,I2683,I320917,I321237,);
nor I_18737 (I320885,I321237,I321141);
not I_18738 (I321259,I321237);
nor I_18739 (I321276,I321259,I321050);
nor I_18740 (I321293,I320982,I321276);
DFFARX1 I_18741 (I321293,I2683,I320917,I320900,);
nor I_18742 (I321324,I321259,I321141);
nor I_18743 (I321341,I724513,I724528);
nor I_18744 (I320891,I321341,I321324);
not I_18745 (I321372,I321341);
nand I_18746 (I320894,I321101,I321372);
DFFARX1 I_18747 (I321341,I2683,I320917,I320906,);
DFFARX1 I_18748 (I321341,I2683,I320917,I320903,);
not I_18749 (I321461,I2690);
DFFARX1 I_18750 (I843227,I2683,I321461,I321487,);
DFFARX1 I_18751 (I321487,I2683,I321461,I321504,);
not I_18752 (I321453,I321504);
not I_18753 (I321526,I321487);
nand I_18754 (I321543,I843239,I843227);
and I_18755 (I321560,I321543,I843230);
DFFARX1 I_18756 (I321560,I2683,I321461,I321586,);
not I_18757 (I321594,I321586);
DFFARX1 I_18758 (I843248,I2683,I321461,I321620,);
and I_18759 (I321628,I321620,I843224);
nand I_18760 (I321645,I321620,I843224);
nand I_18761 (I321432,I321594,I321645);
DFFARX1 I_18762 (I843242,I2683,I321461,I321685,);
nor I_18763 (I321693,I321685,I321628);
DFFARX1 I_18764 (I321693,I2683,I321461,I321426,);
nor I_18765 (I321441,I321685,I321586);
nand I_18766 (I321738,I843236,I843233);
and I_18767 (I321755,I321738,I843245);
DFFARX1 I_18768 (I321755,I2683,I321461,I321781,);
nor I_18769 (I321429,I321781,I321685);
not I_18770 (I321803,I321781);
nor I_18771 (I321820,I321803,I321594);
nor I_18772 (I321837,I321526,I321820);
DFFARX1 I_18773 (I321837,I2683,I321461,I321444,);
nor I_18774 (I321868,I321803,I321685);
nor I_18775 (I321885,I843224,I843233);
nor I_18776 (I321435,I321885,I321868);
not I_18777 (I321916,I321885);
nand I_18778 (I321438,I321645,I321916);
DFFARX1 I_18779 (I321885,I2683,I321461,I321450,);
DFFARX1 I_18780 (I321885,I2683,I321461,I321447,);
not I_18781 (I322005,I2690);
DFFARX1 I_18782 (I28494,I2683,I322005,I322031,);
DFFARX1 I_18783 (I322031,I2683,I322005,I322048,);
not I_18784 (I321997,I322048);
not I_18785 (I322070,I322031);
nand I_18786 (I322087,I28482,I28497);
and I_18787 (I322104,I322087,I28485);
DFFARX1 I_18788 (I322104,I2683,I322005,I322130,);
not I_18789 (I322138,I322130);
DFFARX1 I_18790 (I28506,I2683,I322005,I322164,);
and I_18791 (I322172,I322164,I28500);
nand I_18792 (I322189,I322164,I28500);
nand I_18793 (I321976,I322138,I322189);
DFFARX1 I_18794 (I28503,I2683,I322005,I322229,);
nor I_18795 (I322237,I322229,I322172);
DFFARX1 I_18796 (I322237,I2683,I322005,I321970,);
nor I_18797 (I321985,I322229,I322130);
nand I_18798 (I322282,I28482,I28485);
and I_18799 (I322299,I322282,I28488);
DFFARX1 I_18800 (I322299,I2683,I322005,I322325,);
nor I_18801 (I321973,I322325,I322229);
not I_18802 (I322347,I322325);
nor I_18803 (I322364,I322347,I322138);
nor I_18804 (I322381,I322070,I322364);
DFFARX1 I_18805 (I322381,I2683,I322005,I321988,);
nor I_18806 (I322412,I322347,I322229);
nor I_18807 (I322429,I28491,I28485);
nor I_18808 (I321979,I322429,I322412);
not I_18809 (I322460,I322429);
nand I_18810 (I321982,I322189,I322460);
DFFARX1 I_18811 (I322429,I2683,I322005,I321994,);
DFFARX1 I_18812 (I322429,I2683,I322005,I321991,);
not I_18813 (I322549,I2690);
DFFARX1 I_18814 (I892935,I2683,I322549,I322575,);
DFFARX1 I_18815 (I322575,I2683,I322549,I322592,);
not I_18816 (I322541,I322592);
not I_18817 (I322614,I322575);
nand I_18818 (I322631,I892947,I892935);
and I_18819 (I322648,I322631,I892938);
DFFARX1 I_18820 (I322648,I2683,I322549,I322674,);
not I_18821 (I322682,I322674);
DFFARX1 I_18822 (I892956,I2683,I322549,I322708,);
and I_18823 (I322716,I322708,I892932);
nand I_18824 (I322733,I322708,I892932);
nand I_18825 (I322520,I322682,I322733);
DFFARX1 I_18826 (I892950,I2683,I322549,I322773,);
nor I_18827 (I322781,I322773,I322716);
DFFARX1 I_18828 (I322781,I2683,I322549,I322514,);
nor I_18829 (I322529,I322773,I322674);
nand I_18830 (I322826,I892944,I892941);
and I_18831 (I322843,I322826,I892953);
DFFARX1 I_18832 (I322843,I2683,I322549,I322869,);
nor I_18833 (I322517,I322869,I322773);
not I_18834 (I322891,I322869);
nor I_18835 (I322908,I322891,I322682);
nor I_18836 (I322925,I322614,I322908);
DFFARX1 I_18837 (I322925,I2683,I322549,I322532,);
nor I_18838 (I322956,I322891,I322773);
nor I_18839 (I322973,I892932,I892941);
nor I_18840 (I322523,I322973,I322956);
not I_18841 (I323004,I322973);
nand I_18842 (I322526,I322733,I323004);
DFFARX1 I_18843 (I322973,I2683,I322549,I322538,);
DFFARX1 I_18844 (I322973,I2683,I322549,I322535,);
not I_18845 (I323093,I2690);
DFFARX1 I_18846 (I714829,I2683,I323093,I323119,);
DFFARX1 I_18847 (I323119,I2683,I323093,I323136,);
not I_18848 (I323085,I323136);
not I_18849 (I323158,I323119);
nand I_18850 (I323175,I714844,I714832);
and I_18851 (I323192,I323175,I714823);
DFFARX1 I_18852 (I323192,I2683,I323093,I323218,);
not I_18853 (I323226,I323218);
DFFARX1 I_18854 (I714835,I2683,I323093,I323252,);
and I_18855 (I323260,I323252,I714826);
nand I_18856 (I323277,I323252,I714826);
nand I_18857 (I323064,I323226,I323277);
DFFARX1 I_18858 (I714841,I2683,I323093,I323317,);
nor I_18859 (I323325,I323317,I323260);
DFFARX1 I_18860 (I323325,I2683,I323093,I323058,);
nor I_18861 (I323073,I323317,I323218);
nand I_18862 (I323370,I714850,I714838);
and I_18863 (I323387,I323370,I714847);
DFFARX1 I_18864 (I323387,I2683,I323093,I323413,);
nor I_18865 (I323061,I323413,I323317);
not I_18866 (I323435,I323413);
nor I_18867 (I323452,I323435,I323226);
nor I_18868 (I323469,I323158,I323452);
DFFARX1 I_18869 (I323469,I2683,I323093,I323076,);
nor I_18870 (I323500,I323435,I323317);
nor I_18871 (I323517,I714823,I714838);
nor I_18872 (I323067,I323517,I323500);
not I_18873 (I323548,I323517);
nand I_18874 (I323070,I323277,I323548);
DFFARX1 I_18875 (I323517,I2683,I323093,I323082,);
DFFARX1 I_18876 (I323517,I2683,I323093,I323079,);
not I_18877 (I323637,I2690);
DFFARX1 I_18878 (I964641,I2683,I323637,I323663,);
DFFARX1 I_18879 (I323663,I2683,I323637,I323680,);
not I_18880 (I323629,I323680);
not I_18881 (I323702,I323663);
nand I_18882 (I323719,I964653,I964656);
and I_18883 (I323736,I323719,I964659);
DFFARX1 I_18884 (I323736,I2683,I323637,I323762,);
not I_18885 (I323770,I323762);
DFFARX1 I_18886 (I964644,I2683,I323637,I323796,);
and I_18887 (I323804,I323796,I964650);
nand I_18888 (I323821,I323796,I964650);
nand I_18889 (I323608,I323770,I323821);
DFFARX1 I_18890 (I964638,I2683,I323637,I323861,);
nor I_18891 (I323869,I323861,I323804);
DFFARX1 I_18892 (I323869,I2683,I323637,I323602,);
nor I_18893 (I323617,I323861,I323762);
nand I_18894 (I323914,I964641,I964662);
and I_18895 (I323931,I323914,I964647);
DFFARX1 I_18896 (I323931,I2683,I323637,I323957,);
nor I_18897 (I323605,I323957,I323861);
not I_18898 (I323979,I323957);
nor I_18899 (I323996,I323979,I323770);
nor I_18900 (I324013,I323702,I323996);
DFFARX1 I_18901 (I324013,I2683,I323637,I323620,);
nor I_18902 (I324044,I323979,I323861);
nor I_18903 (I324061,I964638,I964662);
nor I_18904 (I323611,I324061,I324044);
not I_18905 (I324092,I324061);
nand I_18906 (I323614,I323821,I324092);
DFFARX1 I_18907 (I324061,I2683,I323637,I323626,);
DFFARX1 I_18908 (I324061,I2683,I323637,I323623,);
not I_18909 (I324181,I2690);
DFFARX1 I_18910 (I1003042,I2683,I324181,I324207,);
DFFARX1 I_18911 (I324207,I2683,I324181,I324224,);
not I_18912 (I324173,I324224);
not I_18913 (I324246,I324207);
nand I_18914 (I324263,I1003039,I1003036);
and I_18915 (I324280,I324263,I1003024);
DFFARX1 I_18916 (I324280,I2683,I324181,I324306,);
not I_18917 (I324314,I324306);
DFFARX1 I_18918 (I1003048,I2683,I324181,I324340,);
and I_18919 (I324348,I324340,I1003033);
nand I_18920 (I324365,I324340,I1003033);
nand I_18921 (I324152,I324314,I324365);
DFFARX1 I_18922 (I1003027,I2683,I324181,I324405,);
nor I_18923 (I324413,I324405,I324348);
DFFARX1 I_18924 (I324413,I2683,I324181,I324146,);
nor I_18925 (I324161,I324405,I324306);
nand I_18926 (I324458,I1003024,I1003030);
and I_18927 (I324475,I324458,I1003045);
DFFARX1 I_18928 (I324475,I2683,I324181,I324501,);
nor I_18929 (I324149,I324501,I324405);
not I_18930 (I324523,I324501);
nor I_18931 (I324540,I324523,I324314);
nor I_18932 (I324557,I324246,I324540);
DFFARX1 I_18933 (I324557,I2683,I324181,I324164,);
nor I_18934 (I324588,I324523,I324405);
nor I_18935 (I324605,I1003027,I1003030);
nor I_18936 (I324155,I324605,I324588);
not I_18937 (I324636,I324605);
nand I_18938 (I324158,I324365,I324636);
DFFARX1 I_18939 (I324605,I2683,I324181,I324170,);
DFFARX1 I_18940 (I324605,I2683,I324181,I324167,);
not I_18941 (I324725,I2690);
DFFARX1 I_18942 (I221674,I2683,I324725,I324751,);
DFFARX1 I_18943 (I324751,I2683,I324725,I324768,);
not I_18944 (I324717,I324768);
not I_18945 (I324790,I324751);
nand I_18946 (I324807,I221653,I221677);
and I_18947 (I324824,I324807,I221680);
DFFARX1 I_18948 (I324824,I2683,I324725,I324850,);
not I_18949 (I324858,I324850);
DFFARX1 I_18950 (I221662,I2683,I324725,I324884,);
and I_18951 (I324892,I324884,I221668);
nand I_18952 (I324909,I324884,I221668);
nand I_18953 (I324696,I324858,I324909);
DFFARX1 I_18954 (I221656,I2683,I324725,I324949,);
nor I_18955 (I324957,I324949,I324892);
DFFARX1 I_18956 (I324957,I2683,I324725,I324690,);
nor I_18957 (I324705,I324949,I324850);
nand I_18958 (I325002,I221665,I221653);
and I_18959 (I325019,I325002,I221659);
DFFARX1 I_18960 (I325019,I2683,I324725,I325045,);
nor I_18961 (I324693,I325045,I324949);
not I_18962 (I325067,I325045);
nor I_18963 (I325084,I325067,I324858);
nor I_18964 (I325101,I324790,I325084);
DFFARX1 I_18965 (I325101,I2683,I324725,I324708,);
nor I_18966 (I325132,I325067,I324949);
nor I_18967 (I325149,I221671,I221653);
nor I_18968 (I324699,I325149,I325132);
not I_18969 (I325180,I325149);
nand I_18970 (I324702,I324909,I325180);
DFFARX1 I_18971 (I325149,I2683,I324725,I324714,);
DFFARX1 I_18972 (I325149,I2683,I324725,I324711,);
not I_18973 (I325269,I2690);
DFFARX1 I_18974 (I739377,I2683,I325269,I325295,);
DFFARX1 I_18975 (I325295,I2683,I325269,I325312,);
not I_18976 (I325261,I325312);
not I_18977 (I325334,I325295);
nand I_18978 (I325351,I739392,I739380);
and I_18979 (I325368,I325351,I739371);
DFFARX1 I_18980 (I325368,I2683,I325269,I325394,);
not I_18981 (I325402,I325394);
DFFARX1 I_18982 (I739383,I2683,I325269,I325428,);
and I_18983 (I325436,I325428,I739374);
nand I_18984 (I325453,I325428,I739374);
nand I_18985 (I325240,I325402,I325453);
DFFARX1 I_18986 (I739389,I2683,I325269,I325493,);
nor I_18987 (I325501,I325493,I325436);
DFFARX1 I_18988 (I325501,I2683,I325269,I325234,);
nor I_18989 (I325249,I325493,I325394);
nand I_18990 (I325546,I739398,I739386);
and I_18991 (I325563,I325546,I739395);
DFFARX1 I_18992 (I325563,I2683,I325269,I325589,);
nor I_18993 (I325237,I325589,I325493);
not I_18994 (I325611,I325589);
nor I_18995 (I325628,I325611,I325402);
nor I_18996 (I325645,I325334,I325628);
DFFARX1 I_18997 (I325645,I2683,I325269,I325252,);
nor I_18998 (I325676,I325611,I325493);
nor I_18999 (I325693,I739371,I739386);
nor I_19000 (I325243,I325693,I325676);
not I_19001 (I325724,I325693);
nand I_19002 (I325246,I325453,I325724);
DFFARX1 I_19003 (I325693,I2683,I325269,I325258,);
DFFARX1 I_19004 (I325693,I2683,I325269,I325255,);
not I_19005 (I325813,I2690);
DFFARX1 I_19006 (I718705,I2683,I325813,I325839,);
DFFARX1 I_19007 (I325839,I2683,I325813,I325856,);
not I_19008 (I325805,I325856);
not I_19009 (I325878,I325839);
nand I_19010 (I325895,I718720,I718708);
and I_19011 (I325912,I325895,I718699);
DFFARX1 I_19012 (I325912,I2683,I325813,I325938,);
not I_19013 (I325946,I325938);
DFFARX1 I_19014 (I718711,I2683,I325813,I325972,);
and I_19015 (I325980,I325972,I718702);
nand I_19016 (I325997,I325972,I718702);
nand I_19017 (I325784,I325946,I325997);
DFFARX1 I_19018 (I718717,I2683,I325813,I326037,);
nor I_19019 (I326045,I326037,I325980);
DFFARX1 I_19020 (I326045,I2683,I325813,I325778,);
nor I_19021 (I325793,I326037,I325938);
nand I_19022 (I326090,I718726,I718714);
and I_19023 (I326107,I326090,I718723);
DFFARX1 I_19024 (I326107,I2683,I325813,I326133,);
nor I_19025 (I325781,I326133,I326037);
not I_19026 (I326155,I326133);
nor I_19027 (I326172,I326155,I325946);
nor I_19028 (I326189,I325878,I326172);
DFFARX1 I_19029 (I326189,I2683,I325813,I325796,);
nor I_19030 (I326220,I326155,I326037);
nor I_19031 (I326237,I718699,I718714);
nor I_19032 (I325787,I326237,I326220);
not I_19033 (I326268,I326237);
nand I_19034 (I325790,I325997,I326268);
DFFARX1 I_19035 (I326237,I2683,I325813,I325802,);
DFFARX1 I_19036 (I326237,I2683,I325813,I325799,);
not I_19037 (I326357,I2690);
DFFARX1 I_19038 (I1057876,I2683,I326357,I326383,);
DFFARX1 I_19039 (I326383,I2683,I326357,I326400,);
not I_19040 (I326349,I326400);
not I_19041 (I326422,I326383);
nand I_19042 (I326439,I1057852,I1057873);
and I_19043 (I326456,I326439,I1057870);
DFFARX1 I_19044 (I326456,I2683,I326357,I326482,);
not I_19045 (I326490,I326482);
DFFARX1 I_19046 (I1057849,I2683,I326357,I326516,);
and I_19047 (I326524,I326516,I1057861);
nand I_19048 (I326541,I326516,I1057861);
nand I_19049 (I326328,I326490,I326541);
DFFARX1 I_19050 (I1057864,I2683,I326357,I326581,);
nor I_19051 (I326589,I326581,I326524);
DFFARX1 I_19052 (I326589,I2683,I326357,I326322,);
nor I_19053 (I326337,I326581,I326482);
nand I_19054 (I326634,I1057867,I1057855);
and I_19055 (I326651,I326634,I1057858);
DFFARX1 I_19056 (I326651,I2683,I326357,I326677,);
nor I_19057 (I326325,I326677,I326581);
not I_19058 (I326699,I326677);
nor I_19059 (I326716,I326699,I326490);
nor I_19060 (I326733,I326422,I326716);
DFFARX1 I_19061 (I326733,I2683,I326357,I326340,);
nor I_19062 (I326764,I326699,I326581);
nor I_19063 (I326781,I1057849,I1057855);
nor I_19064 (I326331,I326781,I326764);
not I_19065 (I326812,I326781);
nand I_19066 (I326334,I326541,I326812);
DFFARX1 I_19067 (I326781,I2683,I326357,I326346,);
DFFARX1 I_19068 (I326781,I2683,I326357,I326343,);
not I_19069 (I326901,I2690);
DFFARX1 I_19070 (I772969,I2683,I326901,I326927,);
DFFARX1 I_19071 (I326927,I2683,I326901,I326944,);
not I_19072 (I326893,I326944);
not I_19073 (I326966,I326927);
nand I_19074 (I326983,I772984,I772972);
and I_19075 (I327000,I326983,I772963);
DFFARX1 I_19076 (I327000,I2683,I326901,I327026,);
not I_19077 (I327034,I327026);
DFFARX1 I_19078 (I772975,I2683,I326901,I327060,);
and I_19079 (I327068,I327060,I772966);
nand I_19080 (I327085,I327060,I772966);
nand I_19081 (I326872,I327034,I327085);
DFFARX1 I_19082 (I772981,I2683,I326901,I327125,);
nor I_19083 (I327133,I327125,I327068);
DFFARX1 I_19084 (I327133,I2683,I326901,I326866,);
nor I_19085 (I326881,I327125,I327026);
nand I_19086 (I327178,I772990,I772978);
and I_19087 (I327195,I327178,I772987);
DFFARX1 I_19088 (I327195,I2683,I326901,I327221,);
nor I_19089 (I326869,I327221,I327125);
not I_19090 (I327243,I327221);
nor I_19091 (I327260,I327243,I327034);
nor I_19092 (I327277,I326966,I327260);
DFFARX1 I_19093 (I327277,I2683,I326901,I326884,);
nor I_19094 (I327308,I327243,I327125);
nor I_19095 (I327325,I772963,I772978);
nor I_19096 (I326875,I327325,I327308);
not I_19097 (I327356,I327325);
nand I_19098 (I326878,I327085,I327356);
DFFARX1 I_19099 (I327325,I2683,I326901,I326890,);
DFFARX1 I_19100 (I327325,I2683,I326901,I326887,);
not I_19101 (I327445,I2690);
DFFARX1 I_19102 (I435873,I2683,I327445,I327471,);
DFFARX1 I_19103 (I327471,I2683,I327445,I327488,);
not I_19104 (I327437,I327488);
not I_19105 (I327510,I327471);
nand I_19106 (I327527,I435870,I435891);
and I_19107 (I327544,I327527,I435894);
DFFARX1 I_19108 (I327544,I2683,I327445,I327570,);
not I_19109 (I327578,I327570);
DFFARX1 I_19110 (I435879,I2683,I327445,I327604,);
and I_19111 (I327612,I327604,I435882);
nand I_19112 (I327629,I327604,I435882);
nand I_19113 (I327416,I327578,I327629);
DFFARX1 I_19114 (I435885,I2683,I327445,I327669,);
nor I_19115 (I327677,I327669,I327612);
DFFARX1 I_19116 (I327677,I2683,I327445,I327410,);
nor I_19117 (I327425,I327669,I327570);
nand I_19118 (I327722,I435870,I435876);
and I_19119 (I327739,I327722,I435888);
DFFARX1 I_19120 (I327739,I2683,I327445,I327765,);
nor I_19121 (I327413,I327765,I327669);
not I_19122 (I327787,I327765);
nor I_19123 (I327804,I327787,I327578);
nor I_19124 (I327821,I327510,I327804);
DFFARX1 I_19125 (I327821,I2683,I327445,I327428,);
nor I_19126 (I327852,I327787,I327669);
nor I_19127 (I327869,I435873,I435876);
nor I_19128 (I327419,I327869,I327852);
not I_19129 (I327900,I327869);
nand I_19130 (I327422,I327629,I327900);
DFFARX1 I_19131 (I327869,I2683,I327445,I327434,);
DFFARX1 I_19132 (I327869,I2683,I327445,I327431,);
not I_19133 (I327989,I2690);
DFFARX1 I_19134 (I1033481,I2683,I327989,I328015,);
DFFARX1 I_19135 (I328015,I2683,I327989,I328032,);
not I_19136 (I327981,I328032);
not I_19137 (I328054,I328015);
nand I_19138 (I328071,I1033457,I1033478);
and I_19139 (I328088,I328071,I1033475);
DFFARX1 I_19140 (I328088,I2683,I327989,I328114,);
not I_19141 (I328122,I328114);
DFFARX1 I_19142 (I1033454,I2683,I327989,I328148,);
and I_19143 (I328156,I328148,I1033466);
nand I_19144 (I328173,I328148,I1033466);
nand I_19145 (I327960,I328122,I328173);
DFFARX1 I_19146 (I1033469,I2683,I327989,I328213,);
nor I_19147 (I328221,I328213,I328156);
DFFARX1 I_19148 (I328221,I2683,I327989,I327954,);
nor I_19149 (I327969,I328213,I328114);
nand I_19150 (I328266,I1033472,I1033460);
and I_19151 (I328283,I328266,I1033463);
DFFARX1 I_19152 (I328283,I2683,I327989,I328309,);
nor I_19153 (I327957,I328309,I328213);
not I_19154 (I328331,I328309);
nor I_19155 (I328348,I328331,I328122);
nor I_19156 (I328365,I328054,I328348);
DFFARX1 I_19157 (I328365,I2683,I327989,I327972,);
nor I_19158 (I328396,I328331,I328213);
nor I_19159 (I328413,I1033454,I1033460);
nor I_19160 (I327963,I328413,I328396);
not I_19161 (I328444,I328413);
nand I_19162 (I327966,I328173,I328444);
DFFARX1 I_19163 (I328413,I2683,I327989,I327978,);
DFFARX1 I_19164 (I328413,I2683,I327989,I327975,);
not I_19165 (I328533,I2690);
DFFARX1 I_19166 (I121804,I2683,I328533,I328559,);
DFFARX1 I_19167 (I328559,I2683,I328533,I328576,);
not I_19168 (I328525,I328576);
not I_19169 (I328598,I328559);
nand I_19170 (I328615,I121816,I121795);
and I_19171 (I328632,I328615,I121798);
DFFARX1 I_19172 (I328632,I2683,I328533,I328658,);
not I_19173 (I328666,I328658);
DFFARX1 I_19174 (I121807,I2683,I328533,I328692,);
and I_19175 (I328700,I328692,I121819);
nand I_19176 (I328717,I328692,I121819);
nand I_19177 (I328504,I328666,I328717);
DFFARX1 I_19178 (I121813,I2683,I328533,I328757,);
nor I_19179 (I328765,I328757,I328700);
DFFARX1 I_19180 (I328765,I2683,I328533,I328498,);
nor I_19181 (I328513,I328757,I328658);
nand I_19182 (I328810,I121801,I121798);
and I_19183 (I328827,I328810,I121810);
DFFARX1 I_19184 (I328827,I2683,I328533,I328853,);
nor I_19185 (I328501,I328853,I328757);
not I_19186 (I328875,I328853);
nor I_19187 (I328892,I328875,I328666);
nor I_19188 (I328909,I328598,I328892);
DFFARX1 I_19189 (I328909,I2683,I328533,I328516,);
nor I_19190 (I328940,I328875,I328757);
nor I_19191 (I328957,I121795,I121798);
nor I_19192 (I328507,I328957,I328940);
not I_19193 (I328988,I328957);
nand I_19194 (I328510,I328717,I328988);
DFFARX1 I_19195 (I328957,I2683,I328533,I328522,);
DFFARX1 I_19196 (I328957,I2683,I328533,I328519,);
not I_19197 (I329077,I2690);
DFFARX1 I_19198 (I1098931,I2683,I329077,I329103,);
DFFARX1 I_19199 (I329103,I2683,I329077,I329120,);
not I_19200 (I329069,I329120);
not I_19201 (I329142,I329103);
nand I_19202 (I329159,I1098907,I1098928);
and I_19203 (I329176,I329159,I1098925);
DFFARX1 I_19204 (I329176,I2683,I329077,I329202,);
not I_19205 (I329210,I329202);
DFFARX1 I_19206 (I1098904,I2683,I329077,I329236,);
and I_19207 (I329244,I329236,I1098916);
nand I_19208 (I329261,I329236,I1098916);
nand I_19209 (I329048,I329210,I329261);
DFFARX1 I_19210 (I1098919,I2683,I329077,I329301,);
nor I_19211 (I329309,I329301,I329244);
DFFARX1 I_19212 (I329309,I2683,I329077,I329042,);
nor I_19213 (I329057,I329301,I329202);
nand I_19214 (I329354,I1098922,I1098910);
and I_19215 (I329371,I329354,I1098913);
DFFARX1 I_19216 (I329371,I2683,I329077,I329397,);
nor I_19217 (I329045,I329397,I329301);
not I_19218 (I329419,I329397);
nor I_19219 (I329436,I329419,I329210);
nor I_19220 (I329453,I329142,I329436);
DFFARX1 I_19221 (I329453,I2683,I329077,I329060,);
nor I_19222 (I329484,I329419,I329301);
nor I_19223 (I329501,I1098904,I1098910);
nor I_19224 (I329051,I329501,I329484);
not I_19225 (I329532,I329501);
nand I_19226 (I329054,I329261,I329532);
DFFARX1 I_19227 (I329501,I2683,I329077,I329066,);
DFFARX1 I_19228 (I329501,I2683,I329077,I329063,);
not I_19229 (I329621,I2690);
DFFARX1 I_19230 (I669700,I2683,I329621,I329647,);
DFFARX1 I_19231 (I329647,I2683,I329621,I329664,);
not I_19232 (I329613,I329664);
not I_19233 (I329686,I329647);
nand I_19234 (I329703,I669694,I669691);
and I_19235 (I329720,I329703,I669706);
DFFARX1 I_19236 (I329720,I2683,I329621,I329746,);
not I_19237 (I329754,I329746);
DFFARX1 I_19238 (I669694,I2683,I329621,I329780,);
and I_19239 (I329788,I329780,I669688);
nand I_19240 (I329805,I329780,I669688);
nand I_19241 (I329592,I329754,I329805);
DFFARX1 I_19242 (I669688,I2683,I329621,I329845,);
nor I_19243 (I329853,I329845,I329788);
DFFARX1 I_19244 (I329853,I2683,I329621,I329586,);
nor I_19245 (I329601,I329845,I329746);
nand I_19246 (I329898,I669703,I669697);
and I_19247 (I329915,I329898,I669691);
DFFARX1 I_19248 (I329915,I2683,I329621,I329941,);
nor I_19249 (I329589,I329941,I329845);
not I_19250 (I329963,I329941);
nor I_19251 (I329980,I329963,I329754);
nor I_19252 (I329997,I329686,I329980);
DFFARX1 I_19253 (I329997,I2683,I329621,I329604,);
nor I_19254 (I330028,I329963,I329845);
nor I_19255 (I330045,I669709,I669697);
nor I_19256 (I329595,I330045,I330028);
not I_19257 (I330076,I330045);
nand I_19258 (I329598,I329805,I330076);
DFFARX1 I_19259 (I330045,I2683,I329621,I329610,);
DFFARX1 I_19260 (I330045,I2683,I329621,I329607,);
not I_19261 (I330165,I2690);
DFFARX1 I_19262 (I876173,I2683,I330165,I330191,);
DFFARX1 I_19263 (I330191,I2683,I330165,I330208,);
not I_19264 (I330157,I330208);
not I_19265 (I330230,I330191);
nand I_19266 (I330247,I876185,I876173);
and I_19267 (I330264,I330247,I876176);
DFFARX1 I_19268 (I330264,I2683,I330165,I330290,);
not I_19269 (I330298,I330290);
DFFARX1 I_19270 (I876194,I2683,I330165,I330324,);
and I_19271 (I330332,I330324,I876170);
nand I_19272 (I330349,I330324,I876170);
nand I_19273 (I330136,I330298,I330349);
DFFARX1 I_19274 (I876188,I2683,I330165,I330389,);
nor I_19275 (I330397,I330389,I330332);
DFFARX1 I_19276 (I330397,I2683,I330165,I330130,);
nor I_19277 (I330145,I330389,I330290);
nand I_19278 (I330442,I876182,I876179);
and I_19279 (I330459,I330442,I876191);
DFFARX1 I_19280 (I330459,I2683,I330165,I330485,);
nor I_19281 (I330133,I330485,I330389);
not I_19282 (I330507,I330485);
nor I_19283 (I330524,I330507,I330298);
nor I_19284 (I330541,I330230,I330524);
DFFARX1 I_19285 (I330541,I2683,I330165,I330148,);
nor I_19286 (I330572,I330507,I330389);
nor I_19287 (I330589,I876170,I876179);
nor I_19288 (I330139,I330589,I330572);
not I_19289 (I330620,I330589);
nand I_19290 (I330142,I330349,I330620);
DFFARX1 I_19291 (I330589,I2683,I330165,I330154,);
DFFARX1 I_19292 (I330589,I2683,I330165,I330151,);
not I_19293 (I330709,I2690);
DFFARX1 I_19294 (I90674,I2683,I330709,I330735,);
DFFARX1 I_19295 (I330735,I2683,I330709,I330752,);
not I_19296 (I330701,I330752);
not I_19297 (I330774,I330735);
nand I_19298 (I330791,I90689,I90668);
and I_19299 (I330808,I330791,I90671);
DFFARX1 I_19300 (I330808,I2683,I330709,I330834,);
not I_19301 (I330842,I330834);
DFFARX1 I_19302 (I90677,I2683,I330709,I330868,);
and I_19303 (I330876,I330868,I90671);
nand I_19304 (I330893,I330868,I90671);
nand I_19305 (I330680,I330842,I330893);
DFFARX1 I_19306 (I90686,I2683,I330709,I330933,);
nor I_19307 (I330941,I330933,I330876);
DFFARX1 I_19308 (I330941,I2683,I330709,I330674,);
nor I_19309 (I330689,I330933,I330834);
nand I_19310 (I330986,I90668,I90683);
and I_19311 (I331003,I330986,I90680);
DFFARX1 I_19312 (I331003,I2683,I330709,I331029,);
nor I_19313 (I330677,I331029,I330933);
not I_19314 (I331051,I331029);
nor I_19315 (I331068,I331051,I330842);
nor I_19316 (I331085,I330774,I331068);
DFFARX1 I_19317 (I331085,I2683,I330709,I330692,);
nor I_19318 (I331116,I331051,I330933);
nor I_19319 (I331133,I90692,I90683);
nor I_19320 (I330683,I331133,I331116);
not I_19321 (I331164,I331133);
nand I_19322 (I330686,I330893,I331164);
DFFARX1 I_19323 (I331133,I2683,I330709,I330698,);
DFFARX1 I_19324 (I331133,I2683,I330709,I330695,);
not I_19325 (I331253,I2690);
DFFARX1 I_19326 (I825952,I2683,I331253,I331279,);
DFFARX1 I_19327 (I331279,I2683,I331253,I331296,);
not I_19328 (I331245,I331296);
not I_19329 (I331318,I331279);
nand I_19330 (I331335,I825952,I825970);
and I_19331 (I331352,I331335,I825964);
DFFARX1 I_19332 (I331352,I2683,I331253,I331378,);
not I_19333 (I331386,I331378);
DFFARX1 I_19334 (I825958,I2683,I331253,I331412,);
and I_19335 (I331420,I331412,I825967);
nand I_19336 (I331437,I331412,I825967);
nand I_19337 (I331224,I331386,I331437);
DFFARX1 I_19338 (I825955,I2683,I331253,I331477,);
nor I_19339 (I331485,I331477,I331420);
DFFARX1 I_19340 (I331485,I2683,I331253,I331218,);
nor I_19341 (I331233,I331477,I331378);
nand I_19342 (I331530,I825955,I825973);
and I_19343 (I331547,I331530,I825958);
DFFARX1 I_19344 (I331547,I2683,I331253,I331573,);
nor I_19345 (I331221,I331573,I331477);
not I_19346 (I331595,I331573);
nor I_19347 (I331612,I331595,I331386);
nor I_19348 (I331629,I331318,I331612);
DFFARX1 I_19349 (I331629,I2683,I331253,I331236,);
nor I_19350 (I331660,I331595,I331477);
nor I_19351 (I331677,I825961,I825973);
nor I_19352 (I331227,I331677,I331660);
not I_19353 (I331708,I331677);
nand I_19354 (I331230,I331437,I331708);
DFFARX1 I_19355 (I331677,I2683,I331253,I331242,);
DFFARX1 I_19356 (I331677,I2683,I331253,I331239,);
not I_19357 (I331797,I2690);
DFFARX1 I_19358 (I59054,I2683,I331797,I331823,);
DFFARX1 I_19359 (I331823,I2683,I331797,I331840,);
not I_19360 (I331789,I331840);
not I_19361 (I331862,I331823);
nand I_19362 (I331879,I59069,I59048);
and I_19363 (I331896,I331879,I59051);
DFFARX1 I_19364 (I331896,I2683,I331797,I331922,);
not I_19365 (I331930,I331922);
DFFARX1 I_19366 (I59057,I2683,I331797,I331956,);
and I_19367 (I331964,I331956,I59051);
nand I_19368 (I331981,I331956,I59051);
nand I_19369 (I331768,I331930,I331981);
DFFARX1 I_19370 (I59066,I2683,I331797,I332021,);
nor I_19371 (I332029,I332021,I331964);
DFFARX1 I_19372 (I332029,I2683,I331797,I331762,);
nor I_19373 (I331777,I332021,I331922);
nand I_19374 (I332074,I59048,I59063);
and I_19375 (I332091,I332074,I59060);
DFFARX1 I_19376 (I332091,I2683,I331797,I332117,);
nor I_19377 (I331765,I332117,I332021);
not I_19378 (I332139,I332117);
nor I_19379 (I332156,I332139,I331930);
nor I_19380 (I332173,I331862,I332156);
DFFARX1 I_19381 (I332173,I2683,I331797,I331780,);
nor I_19382 (I332204,I332139,I332021);
nor I_19383 (I332221,I59072,I59063);
nor I_19384 (I331771,I332221,I332204);
not I_19385 (I332252,I332221);
nand I_19386 (I331774,I331981,I332252);
DFFARX1 I_19387 (I332221,I2683,I331797,I331786,);
DFFARX1 I_19388 (I332221,I2683,I331797,I331783,);
not I_19389 (I332341,I2690);
DFFARX1 I_19390 (I174759,I2683,I332341,I332367,);
DFFARX1 I_19391 (I332367,I2683,I332341,I332384,);
not I_19392 (I332333,I332384);
not I_19393 (I332406,I332367);
nand I_19394 (I332423,I174771,I174750);
and I_19395 (I332440,I332423,I174753);
DFFARX1 I_19396 (I332440,I2683,I332341,I332466,);
not I_19397 (I332474,I332466);
DFFARX1 I_19398 (I174762,I2683,I332341,I332500,);
and I_19399 (I332508,I332500,I174774);
nand I_19400 (I332525,I332500,I174774);
nand I_19401 (I332312,I332474,I332525);
DFFARX1 I_19402 (I174768,I2683,I332341,I332565,);
nor I_19403 (I332573,I332565,I332508);
DFFARX1 I_19404 (I332573,I2683,I332341,I332306,);
nor I_19405 (I332321,I332565,I332466);
nand I_19406 (I332618,I174756,I174753);
and I_19407 (I332635,I332618,I174765);
DFFARX1 I_19408 (I332635,I2683,I332341,I332661,);
nor I_19409 (I332309,I332661,I332565);
not I_19410 (I332683,I332661);
nor I_19411 (I332700,I332683,I332474);
nor I_19412 (I332717,I332406,I332700);
DFFARX1 I_19413 (I332717,I2683,I332341,I332324,);
nor I_19414 (I332748,I332683,I332565);
nor I_19415 (I332765,I174750,I174753);
nor I_19416 (I332315,I332765,I332748);
not I_19417 (I332796,I332765);
nand I_19418 (I332318,I332525,I332796);
DFFARX1 I_19419 (I332765,I2683,I332341,I332330,);
DFFARX1 I_19420 (I332765,I2683,I332341,I332327,);
not I_19421 (I332885,I2690);
DFFARX1 I_19422 (I35872,I2683,I332885,I332911,);
DFFARX1 I_19423 (I332911,I2683,I332885,I332928,);
not I_19424 (I332877,I332928);
not I_19425 (I332950,I332911);
nand I_19426 (I332967,I35860,I35875);
and I_19427 (I332984,I332967,I35863);
DFFARX1 I_19428 (I332984,I2683,I332885,I333010,);
not I_19429 (I333018,I333010);
DFFARX1 I_19430 (I35884,I2683,I332885,I333044,);
and I_19431 (I333052,I333044,I35878);
nand I_19432 (I333069,I333044,I35878);
nand I_19433 (I332856,I333018,I333069);
DFFARX1 I_19434 (I35881,I2683,I332885,I333109,);
nor I_19435 (I333117,I333109,I333052);
DFFARX1 I_19436 (I333117,I2683,I332885,I332850,);
nor I_19437 (I332865,I333109,I333010);
nand I_19438 (I333162,I35860,I35863);
and I_19439 (I333179,I333162,I35866);
DFFARX1 I_19440 (I333179,I2683,I332885,I333205,);
nor I_19441 (I332853,I333205,I333109);
not I_19442 (I333227,I333205);
nor I_19443 (I333244,I333227,I333018);
nor I_19444 (I333261,I332950,I333244);
DFFARX1 I_19445 (I333261,I2683,I332885,I332868,);
nor I_19446 (I333292,I333227,I333109);
nor I_19447 (I333309,I35869,I35863);
nor I_19448 (I332859,I333309,I333292);
not I_19449 (I333340,I333309);
nand I_19450 (I332862,I333069,I333340);
DFFARX1 I_19451 (I333309,I2683,I332885,I332874,);
DFFARX1 I_19452 (I333309,I2683,I332885,I332871,);
not I_19453 (I333429,I2690);
DFFARX1 I_19454 (I727103,I2683,I333429,I333455,);
DFFARX1 I_19455 (I333455,I2683,I333429,I333472,);
not I_19456 (I333421,I333472);
not I_19457 (I333494,I333455);
nand I_19458 (I333511,I727118,I727106);
and I_19459 (I333528,I333511,I727097);
DFFARX1 I_19460 (I333528,I2683,I333429,I333554,);
not I_19461 (I333562,I333554);
DFFARX1 I_19462 (I727109,I2683,I333429,I333588,);
and I_19463 (I333596,I333588,I727100);
nand I_19464 (I333613,I333588,I727100);
nand I_19465 (I333400,I333562,I333613);
DFFARX1 I_19466 (I727115,I2683,I333429,I333653,);
nor I_19467 (I333661,I333653,I333596);
DFFARX1 I_19468 (I333661,I2683,I333429,I333394,);
nor I_19469 (I333409,I333653,I333554);
nand I_19470 (I333706,I727124,I727112);
and I_19471 (I333723,I333706,I727121);
DFFARX1 I_19472 (I333723,I2683,I333429,I333749,);
nor I_19473 (I333397,I333749,I333653);
not I_19474 (I333771,I333749);
nor I_19475 (I333788,I333771,I333562);
nor I_19476 (I333805,I333494,I333788);
DFFARX1 I_19477 (I333805,I2683,I333429,I333412,);
nor I_19478 (I333836,I333771,I333653);
nor I_19479 (I333853,I727097,I727112);
nor I_19480 (I333403,I333853,I333836);
not I_19481 (I333884,I333853);
nand I_19482 (I333406,I333613,I333884);
DFFARX1 I_19483 (I333853,I2683,I333429,I333418,);
DFFARX1 I_19484 (I333853,I2683,I333429,I333415,);
not I_19485 (I333973,I2690);
DFFARX1 I_19486 (I894091,I2683,I333973,I333999,);
DFFARX1 I_19487 (I333999,I2683,I333973,I334016,);
not I_19488 (I333965,I334016);
not I_19489 (I334038,I333999);
nand I_19490 (I334055,I894103,I894091);
and I_19491 (I334072,I334055,I894094);
DFFARX1 I_19492 (I334072,I2683,I333973,I334098,);
not I_19493 (I334106,I334098);
DFFARX1 I_19494 (I894112,I2683,I333973,I334132,);
and I_19495 (I334140,I334132,I894088);
nand I_19496 (I334157,I334132,I894088);
nand I_19497 (I333944,I334106,I334157);
DFFARX1 I_19498 (I894106,I2683,I333973,I334197,);
nor I_19499 (I334205,I334197,I334140);
DFFARX1 I_19500 (I334205,I2683,I333973,I333938,);
nor I_19501 (I333953,I334197,I334098);
nand I_19502 (I334250,I894100,I894097);
and I_19503 (I334267,I334250,I894109);
DFFARX1 I_19504 (I334267,I2683,I333973,I334293,);
nor I_19505 (I333941,I334293,I334197);
not I_19506 (I334315,I334293);
nor I_19507 (I334332,I334315,I334106);
nor I_19508 (I334349,I334038,I334332);
DFFARX1 I_19509 (I334349,I2683,I333973,I333956,);
nor I_19510 (I334380,I334315,I334197);
nor I_19511 (I334397,I894088,I894097);
nor I_19512 (I333947,I334397,I334380);
not I_19513 (I334428,I334397);
nand I_19514 (I333950,I334157,I334428);
DFFARX1 I_19515 (I334397,I2683,I333973,I333962,);
DFFARX1 I_19516 (I334397,I2683,I333973,I333959,);
not I_19517 (I334517,I2690);
DFFARX1 I_19518 (I1097146,I2683,I334517,I334543,);
DFFARX1 I_19519 (I334543,I2683,I334517,I334560,);
not I_19520 (I334509,I334560);
not I_19521 (I334582,I334543);
nand I_19522 (I334599,I1097122,I1097143);
and I_19523 (I334616,I334599,I1097140);
DFFARX1 I_19524 (I334616,I2683,I334517,I334642,);
not I_19525 (I334650,I334642);
DFFARX1 I_19526 (I1097119,I2683,I334517,I334676,);
and I_19527 (I334684,I334676,I1097131);
nand I_19528 (I334701,I334676,I1097131);
nand I_19529 (I334488,I334650,I334701);
DFFARX1 I_19530 (I1097134,I2683,I334517,I334741,);
nor I_19531 (I334749,I334741,I334684);
DFFARX1 I_19532 (I334749,I2683,I334517,I334482,);
nor I_19533 (I334497,I334741,I334642);
nand I_19534 (I334794,I1097137,I1097125);
and I_19535 (I334811,I334794,I1097128);
DFFARX1 I_19536 (I334811,I2683,I334517,I334837,);
nor I_19537 (I334485,I334837,I334741);
not I_19538 (I334859,I334837);
nor I_19539 (I334876,I334859,I334650);
nor I_19540 (I334893,I334582,I334876);
DFFARX1 I_19541 (I334893,I2683,I334517,I334500,);
nor I_19542 (I334924,I334859,I334741);
nor I_19543 (I334941,I1097119,I1097125);
nor I_19544 (I334491,I334941,I334924);
not I_19545 (I334972,I334941);
nand I_19546 (I334494,I334701,I334972);
DFFARX1 I_19547 (I334941,I2683,I334517,I334506,);
DFFARX1 I_19548 (I334941,I2683,I334517,I334503,);
not I_19549 (I335061,I2690);
DFFARX1 I_19550 (I281752,I2683,I335061,I335087,);
DFFARX1 I_19551 (I335087,I2683,I335061,I335104,);
not I_19552 (I335053,I335104);
not I_19553 (I335126,I335087);
nand I_19554 (I335143,I281731,I281755);
and I_19555 (I335160,I335143,I281758);
DFFARX1 I_19556 (I335160,I2683,I335061,I335186,);
not I_19557 (I335194,I335186);
DFFARX1 I_19558 (I281740,I2683,I335061,I335220,);
and I_19559 (I335228,I335220,I281746);
nand I_19560 (I335245,I335220,I281746);
nand I_19561 (I335032,I335194,I335245);
DFFARX1 I_19562 (I281734,I2683,I335061,I335285,);
nor I_19563 (I335293,I335285,I335228);
DFFARX1 I_19564 (I335293,I2683,I335061,I335026,);
nor I_19565 (I335041,I335285,I335186);
nand I_19566 (I335338,I281743,I281731);
and I_19567 (I335355,I335338,I281737);
DFFARX1 I_19568 (I335355,I2683,I335061,I335381,);
nor I_19569 (I335029,I335381,I335285);
not I_19570 (I335403,I335381);
nor I_19571 (I335420,I335403,I335194);
nor I_19572 (I335437,I335126,I335420);
DFFARX1 I_19573 (I335437,I2683,I335061,I335044,);
nor I_19574 (I335468,I335403,I335285);
nor I_19575 (I335485,I281749,I281731);
nor I_19576 (I335035,I335485,I335468);
not I_19577 (I335516,I335485);
nand I_19578 (I335038,I335245,I335516);
DFFARX1 I_19579 (I335485,I2683,I335061,I335050,);
DFFARX1 I_19580 (I335485,I2683,I335061,I335047,);
not I_19581 (I335605,I2690);
DFFARX1 I_19582 (I579795,I2683,I335605,I335631,);
DFFARX1 I_19583 (I335631,I2683,I335605,I335648,);
not I_19584 (I335597,I335648);
not I_19585 (I335670,I335631);
nand I_19586 (I335687,I579816,I579807);
and I_19587 (I335704,I335687,I579795);
DFFARX1 I_19588 (I335704,I2683,I335605,I335730,);
not I_19589 (I335738,I335730);
DFFARX1 I_19590 (I579801,I2683,I335605,I335764,);
and I_19591 (I335772,I335764,I579798);
nand I_19592 (I335789,I335764,I579798);
nand I_19593 (I335576,I335738,I335789);
DFFARX1 I_19594 (I579792,I2683,I335605,I335829,);
nor I_19595 (I335837,I335829,I335772);
DFFARX1 I_19596 (I335837,I2683,I335605,I335570,);
nor I_19597 (I335585,I335829,I335730);
nand I_19598 (I335882,I579792,I579804);
and I_19599 (I335899,I335882,I579813);
DFFARX1 I_19600 (I335899,I2683,I335605,I335925,);
nor I_19601 (I335573,I335925,I335829);
not I_19602 (I335947,I335925);
nor I_19603 (I335964,I335947,I335738);
nor I_19604 (I335981,I335670,I335964);
DFFARX1 I_19605 (I335981,I2683,I335605,I335588,);
nor I_19606 (I336012,I335947,I335829);
nor I_19607 (I336029,I579810,I579804);
nor I_19608 (I335579,I336029,I336012);
not I_19609 (I336060,I336029);
nand I_19610 (I335582,I335789,I336060);
DFFARX1 I_19611 (I336029,I2683,I335605,I335594,);
DFFARX1 I_19612 (I336029,I2683,I335605,I335591,);
not I_19613 (I336149,I2690);
DFFARX1 I_19614 (I205104,I2683,I336149,I336175,);
DFFARX1 I_19615 (I336175,I2683,I336149,I336192,);
not I_19616 (I336141,I336192);
not I_19617 (I336214,I336175);
nand I_19618 (I336231,I205116,I205095);
and I_19619 (I336248,I336231,I205098);
DFFARX1 I_19620 (I336248,I2683,I336149,I336274,);
not I_19621 (I336282,I336274);
DFFARX1 I_19622 (I205107,I2683,I336149,I336308,);
and I_19623 (I336316,I336308,I205119);
nand I_19624 (I336333,I336308,I205119);
nand I_19625 (I336120,I336282,I336333);
DFFARX1 I_19626 (I205113,I2683,I336149,I336373,);
nor I_19627 (I336381,I336373,I336316);
DFFARX1 I_19628 (I336381,I2683,I336149,I336114,);
nor I_19629 (I336129,I336373,I336274);
nand I_19630 (I336426,I205101,I205098);
and I_19631 (I336443,I336426,I205110);
DFFARX1 I_19632 (I336443,I2683,I336149,I336469,);
nor I_19633 (I336117,I336469,I336373);
not I_19634 (I336491,I336469);
nor I_19635 (I336508,I336491,I336282);
nor I_19636 (I336525,I336214,I336508);
DFFARX1 I_19637 (I336525,I2683,I336149,I336132,);
nor I_19638 (I336556,I336491,I336373);
nor I_19639 (I336573,I205095,I205098);
nor I_19640 (I336123,I336573,I336556);
not I_19641 (I336604,I336573);
nand I_19642 (I336126,I336333,I336604);
DFFARX1 I_19643 (I336573,I2683,I336149,I336138,);
DFFARX1 I_19644 (I336573,I2683,I336149,I336135,);
not I_19645 (I336693,I2690);
DFFARX1 I_19646 (I1032291,I2683,I336693,I336719,);
DFFARX1 I_19647 (I336719,I2683,I336693,I336736,);
not I_19648 (I336685,I336736);
not I_19649 (I336758,I336719);
nand I_19650 (I336775,I1032267,I1032288);
and I_19651 (I336792,I336775,I1032285);
DFFARX1 I_19652 (I336792,I2683,I336693,I336818,);
not I_19653 (I336826,I336818);
DFFARX1 I_19654 (I1032264,I2683,I336693,I336852,);
and I_19655 (I336860,I336852,I1032276);
nand I_19656 (I336877,I336852,I1032276);
nand I_19657 (I336664,I336826,I336877);
DFFARX1 I_19658 (I1032279,I2683,I336693,I336917,);
nor I_19659 (I336925,I336917,I336860);
DFFARX1 I_19660 (I336925,I2683,I336693,I336658,);
nor I_19661 (I336673,I336917,I336818);
nand I_19662 (I336970,I1032282,I1032270);
and I_19663 (I336987,I336970,I1032273);
DFFARX1 I_19664 (I336987,I2683,I336693,I337013,);
nor I_19665 (I336661,I337013,I336917);
not I_19666 (I337035,I337013);
nor I_19667 (I337052,I337035,I336826);
nor I_19668 (I337069,I336758,I337052);
DFFARX1 I_19669 (I337069,I2683,I336693,I336676,);
nor I_19670 (I337100,I337035,I336917);
nor I_19671 (I337117,I1032264,I1032270);
nor I_19672 (I336667,I337117,I337100);
not I_19673 (I337148,I337117);
nand I_19674 (I336670,I336877,I337148);
DFFARX1 I_19675 (I337117,I2683,I336693,I336682,);
DFFARX1 I_19676 (I337117,I2683,I336693,I336679,);
not I_19677 (I337237,I2690);
DFFARX1 I_19678 (I1060851,I2683,I337237,I337263,);
DFFARX1 I_19679 (I337263,I2683,I337237,I337280,);
not I_19680 (I337229,I337280);
not I_19681 (I337302,I337263);
nand I_19682 (I337319,I1060827,I1060848);
and I_19683 (I337336,I337319,I1060845);
DFFARX1 I_19684 (I337336,I2683,I337237,I337362,);
not I_19685 (I337370,I337362);
DFFARX1 I_19686 (I1060824,I2683,I337237,I337396,);
and I_19687 (I337404,I337396,I1060836);
nand I_19688 (I337421,I337396,I1060836);
nand I_19689 (I337208,I337370,I337421);
DFFARX1 I_19690 (I1060839,I2683,I337237,I337461,);
nor I_19691 (I337469,I337461,I337404);
DFFARX1 I_19692 (I337469,I2683,I337237,I337202,);
nor I_19693 (I337217,I337461,I337362);
nand I_19694 (I337514,I1060842,I1060830);
and I_19695 (I337531,I337514,I1060833);
DFFARX1 I_19696 (I337531,I2683,I337237,I337557,);
nor I_19697 (I337205,I337557,I337461);
not I_19698 (I337579,I337557);
nor I_19699 (I337596,I337579,I337370);
nor I_19700 (I337613,I337302,I337596);
DFFARX1 I_19701 (I337613,I2683,I337237,I337220,);
nor I_19702 (I337644,I337579,I337461);
nor I_19703 (I337661,I1060824,I1060830);
nor I_19704 (I337211,I337661,I337644);
not I_19705 (I337692,I337661);
nand I_19706 (I337214,I337421,I337692);
DFFARX1 I_19707 (I337661,I2683,I337237,I337226,);
DFFARX1 I_19708 (I337661,I2683,I337237,I337223,);
not I_19709 (I337781,I2690);
DFFARX1 I_19710 (I583841,I2683,I337781,I337807,);
DFFARX1 I_19711 (I337807,I2683,I337781,I337824,);
not I_19712 (I337773,I337824);
not I_19713 (I337846,I337807);
nand I_19714 (I337863,I583862,I583853);
and I_19715 (I337880,I337863,I583841);
DFFARX1 I_19716 (I337880,I2683,I337781,I337906,);
not I_19717 (I337914,I337906);
DFFARX1 I_19718 (I583847,I2683,I337781,I337940,);
and I_19719 (I337948,I337940,I583844);
nand I_19720 (I337965,I337940,I583844);
nand I_19721 (I337752,I337914,I337965);
DFFARX1 I_19722 (I583838,I2683,I337781,I338005,);
nor I_19723 (I338013,I338005,I337948);
DFFARX1 I_19724 (I338013,I2683,I337781,I337746,);
nor I_19725 (I337761,I338005,I337906);
nand I_19726 (I338058,I583838,I583850);
and I_19727 (I338075,I338058,I583859);
DFFARX1 I_19728 (I338075,I2683,I337781,I338101,);
nor I_19729 (I337749,I338101,I338005);
not I_19730 (I338123,I338101);
nor I_19731 (I338140,I338123,I337914);
nor I_19732 (I338157,I337846,I338140);
DFFARX1 I_19733 (I338157,I2683,I337781,I337764,);
nor I_19734 (I338188,I338123,I338005);
nor I_19735 (I338205,I583856,I583850);
nor I_19736 (I337755,I338205,I338188);
not I_19737 (I338236,I338205);
nand I_19738 (I337758,I337965,I338236);
DFFARX1 I_19739 (I338205,I2683,I337781,I337770,);
DFFARX1 I_19740 (I338205,I2683,I337781,I337767,);
not I_19741 (I338325,I2690);
DFFARX1 I_19742 (I1054306,I2683,I338325,I338351,);
DFFARX1 I_19743 (I338351,I2683,I338325,I338368,);
not I_19744 (I338317,I338368);
not I_19745 (I338390,I338351);
nand I_19746 (I338407,I1054282,I1054303);
and I_19747 (I338424,I338407,I1054300);
DFFARX1 I_19748 (I338424,I2683,I338325,I338450,);
not I_19749 (I338458,I338450);
DFFARX1 I_19750 (I1054279,I2683,I338325,I338484,);
and I_19751 (I338492,I338484,I1054291);
nand I_19752 (I338509,I338484,I1054291);
nand I_19753 (I338296,I338458,I338509);
DFFARX1 I_19754 (I1054294,I2683,I338325,I338549,);
nor I_19755 (I338557,I338549,I338492);
DFFARX1 I_19756 (I338557,I2683,I338325,I338290,);
nor I_19757 (I338305,I338549,I338450);
nand I_19758 (I338602,I1054297,I1054285);
and I_19759 (I338619,I338602,I1054288);
DFFARX1 I_19760 (I338619,I2683,I338325,I338645,);
nor I_19761 (I338293,I338645,I338549);
not I_19762 (I338667,I338645);
nor I_19763 (I338684,I338667,I338458);
nor I_19764 (I338701,I338390,I338684);
DFFARX1 I_19765 (I338701,I2683,I338325,I338308,);
nor I_19766 (I338732,I338667,I338549);
nor I_19767 (I338749,I1054279,I1054285);
nor I_19768 (I338299,I338749,I338732);
not I_19769 (I338780,I338749);
nand I_19770 (I338302,I338509,I338780);
DFFARX1 I_19771 (I338749,I2683,I338325,I338314,);
DFFARX1 I_19772 (I338749,I2683,I338325,I338311,);
not I_19773 (I338869,I2690);
DFFARX1 I_19774 (I241173,I2683,I338869,I338895,);
DFFARX1 I_19775 (I338895,I2683,I338869,I338912,);
not I_19776 (I338861,I338912);
not I_19777 (I338934,I338895);
nand I_19778 (I338951,I241152,I241176);
and I_19779 (I338968,I338951,I241179);
DFFARX1 I_19780 (I338968,I2683,I338869,I338994,);
not I_19781 (I339002,I338994);
DFFARX1 I_19782 (I241161,I2683,I338869,I339028,);
and I_19783 (I339036,I339028,I241167);
nand I_19784 (I339053,I339028,I241167);
nand I_19785 (I338840,I339002,I339053);
DFFARX1 I_19786 (I241155,I2683,I338869,I339093,);
nor I_19787 (I339101,I339093,I339036);
DFFARX1 I_19788 (I339101,I2683,I338869,I338834,);
nor I_19789 (I338849,I339093,I338994);
nand I_19790 (I339146,I241164,I241152);
and I_19791 (I339163,I339146,I241158);
DFFARX1 I_19792 (I339163,I2683,I338869,I339189,);
nor I_19793 (I338837,I339189,I339093);
not I_19794 (I339211,I339189);
nor I_19795 (I339228,I339211,I339002);
nor I_19796 (I339245,I338934,I339228);
DFFARX1 I_19797 (I339245,I2683,I338869,I338852,);
nor I_19798 (I339276,I339211,I339093);
nor I_19799 (I339293,I241170,I241152);
nor I_19800 (I338843,I339293,I339276);
not I_19801 (I339324,I339293);
nand I_19802 (I338846,I339053,I339324);
DFFARX1 I_19803 (I339293,I2683,I338869,I338858,);
DFFARX1 I_19804 (I339293,I2683,I338869,I338855,);
not I_19805 (I339413,I2690);
DFFARX1 I_19806 (I1009400,I2683,I339413,I339439,);
DFFARX1 I_19807 (I339439,I2683,I339413,I339456,);
not I_19808 (I339405,I339456);
not I_19809 (I339478,I339439);
nand I_19810 (I339495,I1009397,I1009394);
and I_19811 (I339512,I339495,I1009382);
DFFARX1 I_19812 (I339512,I2683,I339413,I339538,);
not I_19813 (I339546,I339538);
DFFARX1 I_19814 (I1009406,I2683,I339413,I339572,);
and I_19815 (I339580,I339572,I1009391);
nand I_19816 (I339597,I339572,I1009391);
nand I_19817 (I339384,I339546,I339597);
DFFARX1 I_19818 (I1009385,I2683,I339413,I339637,);
nor I_19819 (I339645,I339637,I339580);
DFFARX1 I_19820 (I339645,I2683,I339413,I339378,);
nor I_19821 (I339393,I339637,I339538);
nand I_19822 (I339690,I1009382,I1009388);
and I_19823 (I339707,I339690,I1009403);
DFFARX1 I_19824 (I339707,I2683,I339413,I339733,);
nor I_19825 (I339381,I339733,I339637);
not I_19826 (I339755,I339733);
nor I_19827 (I339772,I339755,I339546);
nor I_19828 (I339789,I339478,I339772);
DFFARX1 I_19829 (I339789,I2683,I339413,I339396,);
nor I_19830 (I339820,I339755,I339637);
nor I_19831 (I339837,I1009385,I1009388);
nor I_19832 (I339387,I339837,I339820);
not I_19833 (I339868,I339837);
nand I_19834 (I339390,I339597,I339868);
DFFARX1 I_19835 (I339837,I2683,I339413,I339402,);
DFFARX1 I_19836 (I339837,I2683,I339413,I339399,);
not I_19837 (I339957,I2690);
DFFARX1 I_19838 (I1081676,I2683,I339957,I339983,);
DFFARX1 I_19839 (I339983,I2683,I339957,I340000,);
not I_19840 (I339949,I340000);
not I_19841 (I340022,I339983);
nand I_19842 (I340039,I1081652,I1081673);
and I_19843 (I340056,I340039,I1081670);
DFFARX1 I_19844 (I340056,I2683,I339957,I340082,);
not I_19845 (I340090,I340082);
DFFARX1 I_19846 (I1081649,I2683,I339957,I340116,);
and I_19847 (I340124,I340116,I1081661);
nand I_19848 (I340141,I340116,I1081661);
nand I_19849 (I339928,I340090,I340141);
DFFARX1 I_19850 (I1081664,I2683,I339957,I340181,);
nor I_19851 (I340189,I340181,I340124);
DFFARX1 I_19852 (I340189,I2683,I339957,I339922,);
nor I_19853 (I339937,I340181,I340082);
nand I_19854 (I340234,I1081667,I1081655);
and I_19855 (I340251,I340234,I1081658);
DFFARX1 I_19856 (I340251,I2683,I339957,I340277,);
nor I_19857 (I339925,I340277,I340181);
not I_19858 (I340299,I340277);
nor I_19859 (I340316,I340299,I340090);
nor I_19860 (I340333,I340022,I340316);
DFFARX1 I_19861 (I340333,I2683,I339957,I339940,);
nor I_19862 (I340364,I340299,I340181);
nor I_19863 (I340381,I1081649,I1081655);
nor I_19864 (I339931,I340381,I340364);
not I_19865 (I340412,I340381);
nand I_19866 (I339934,I340141,I340412);
DFFARX1 I_19867 (I340381,I2683,I339957,I339946,);
DFFARX1 I_19868 (I340381,I2683,I339957,I339943,);
not I_19869 (I340501,I2690);
DFFARX1 I_19870 (I252240,I2683,I340501,I340527,);
DFFARX1 I_19871 (I340527,I2683,I340501,I340544,);
not I_19872 (I340493,I340544);
not I_19873 (I340566,I340527);
nand I_19874 (I340583,I252219,I252243);
and I_19875 (I340600,I340583,I252246);
DFFARX1 I_19876 (I340600,I2683,I340501,I340626,);
not I_19877 (I340634,I340626);
DFFARX1 I_19878 (I252228,I2683,I340501,I340660,);
and I_19879 (I340668,I340660,I252234);
nand I_19880 (I340685,I340660,I252234);
nand I_19881 (I340472,I340634,I340685);
DFFARX1 I_19882 (I252222,I2683,I340501,I340725,);
nor I_19883 (I340733,I340725,I340668);
DFFARX1 I_19884 (I340733,I2683,I340501,I340466,);
nor I_19885 (I340481,I340725,I340626);
nand I_19886 (I340778,I252231,I252219);
and I_19887 (I340795,I340778,I252225);
DFFARX1 I_19888 (I340795,I2683,I340501,I340821,);
nor I_19889 (I340469,I340821,I340725);
not I_19890 (I340843,I340821);
nor I_19891 (I340860,I340843,I340634);
nor I_19892 (I340877,I340566,I340860);
DFFARX1 I_19893 (I340877,I2683,I340501,I340484,);
nor I_19894 (I340908,I340843,I340725);
nor I_19895 (I340925,I252237,I252219);
nor I_19896 (I340475,I340925,I340908);
not I_19897 (I340956,I340925);
nand I_19898 (I340478,I340685,I340956);
DFFARX1 I_19899 (I340925,I2683,I340501,I340490,);
DFFARX1 I_19900 (I340925,I2683,I340501,I340487,);
not I_19901 (I341045,I2690);
DFFARX1 I_19902 (I669173,I2683,I341045,I341071,);
DFFARX1 I_19903 (I341071,I2683,I341045,I341088,);
not I_19904 (I341037,I341088);
not I_19905 (I341110,I341071);
nand I_19906 (I341127,I669167,I669164);
and I_19907 (I341144,I341127,I669179);
DFFARX1 I_19908 (I341144,I2683,I341045,I341170,);
not I_19909 (I341178,I341170);
DFFARX1 I_19910 (I669167,I2683,I341045,I341204,);
and I_19911 (I341212,I341204,I669161);
nand I_19912 (I341229,I341204,I669161);
nand I_19913 (I341016,I341178,I341229);
DFFARX1 I_19914 (I669161,I2683,I341045,I341269,);
nor I_19915 (I341277,I341269,I341212);
DFFARX1 I_19916 (I341277,I2683,I341045,I341010,);
nor I_19917 (I341025,I341269,I341170);
nand I_19918 (I341322,I669176,I669170);
and I_19919 (I341339,I341322,I669164);
DFFARX1 I_19920 (I341339,I2683,I341045,I341365,);
nor I_19921 (I341013,I341365,I341269);
not I_19922 (I341387,I341365);
nor I_19923 (I341404,I341387,I341178);
nor I_19924 (I341421,I341110,I341404);
DFFARX1 I_19925 (I341421,I2683,I341045,I341028,);
nor I_19926 (I341452,I341387,I341269);
nor I_19927 (I341469,I669182,I669170);
nor I_19928 (I341019,I341469,I341452);
not I_19929 (I341500,I341469);
nand I_19930 (I341022,I341229,I341500);
DFFARX1 I_19931 (I341469,I2683,I341045,I341034,);
DFFARX1 I_19932 (I341469,I2683,I341045,I341031,);
not I_19933 (I341589,I2690);
DFFARX1 I_19934 (I181899,I2683,I341589,I341615,);
DFFARX1 I_19935 (I341615,I2683,I341589,I341632,);
not I_19936 (I341581,I341632);
not I_19937 (I341654,I341615);
nand I_19938 (I341671,I181911,I181890);
and I_19939 (I341688,I341671,I181893);
DFFARX1 I_19940 (I341688,I2683,I341589,I341714,);
not I_19941 (I341722,I341714);
DFFARX1 I_19942 (I181902,I2683,I341589,I341748,);
and I_19943 (I341756,I341748,I181914);
nand I_19944 (I341773,I341748,I181914);
nand I_19945 (I341560,I341722,I341773);
DFFARX1 I_19946 (I181908,I2683,I341589,I341813,);
nor I_19947 (I341821,I341813,I341756);
DFFARX1 I_19948 (I341821,I2683,I341589,I341554,);
nor I_19949 (I341569,I341813,I341714);
nand I_19950 (I341866,I181896,I181893);
and I_19951 (I341883,I341866,I181905);
DFFARX1 I_19952 (I341883,I2683,I341589,I341909,);
nor I_19953 (I341557,I341909,I341813);
not I_19954 (I341931,I341909);
nor I_19955 (I341948,I341931,I341722);
nor I_19956 (I341965,I341654,I341948);
DFFARX1 I_19957 (I341965,I2683,I341589,I341572,);
nor I_19958 (I341996,I341931,I341813);
nor I_19959 (I342013,I181890,I181893);
nor I_19960 (I341563,I342013,I341996);
not I_19961 (I342044,I342013);
nand I_19962 (I341566,I341773,I342044);
DFFARX1 I_19963 (I342013,I2683,I341589,I341578,);
DFFARX1 I_19964 (I342013,I2683,I341589,I341575,);
not I_19965 (I342133,I2690);
DFFARX1 I_19966 (I283333,I2683,I342133,I342159,);
DFFARX1 I_19967 (I342159,I2683,I342133,I342176,);
not I_19968 (I342125,I342176);
not I_19969 (I342198,I342159);
nand I_19970 (I342215,I283312,I283336);
and I_19971 (I342232,I342215,I283339);
DFFARX1 I_19972 (I342232,I2683,I342133,I342258,);
not I_19973 (I342266,I342258);
DFFARX1 I_19974 (I283321,I2683,I342133,I342292,);
and I_19975 (I342300,I342292,I283327);
nand I_19976 (I342317,I342292,I283327);
nand I_19977 (I342104,I342266,I342317);
DFFARX1 I_19978 (I283315,I2683,I342133,I342357,);
nor I_19979 (I342365,I342357,I342300);
DFFARX1 I_19980 (I342365,I2683,I342133,I342098,);
nor I_19981 (I342113,I342357,I342258);
nand I_19982 (I342410,I283324,I283312);
and I_19983 (I342427,I342410,I283318);
DFFARX1 I_19984 (I342427,I2683,I342133,I342453,);
nor I_19985 (I342101,I342453,I342357);
not I_19986 (I342475,I342453);
nor I_19987 (I342492,I342475,I342266);
nor I_19988 (I342509,I342198,I342492);
DFFARX1 I_19989 (I342509,I2683,I342133,I342116,);
nor I_19990 (I342540,I342475,I342357);
nor I_19991 (I342557,I283330,I283312);
nor I_19992 (I342107,I342557,I342540);
not I_19993 (I342588,I342557);
nand I_19994 (I342110,I342317,I342588);
DFFARX1 I_19995 (I342557,I2683,I342133,I342122,);
DFFARX1 I_19996 (I342557,I2683,I342133,I342119,);
not I_19997 (I342677,I2690);
DFFARX1 I_19998 (I459571,I2683,I342677,I342703,);
DFFARX1 I_19999 (I342703,I2683,I342677,I342720,);
not I_20000 (I342669,I342720);
not I_20001 (I342742,I342703);
nand I_20002 (I342759,I459568,I459589);
and I_20003 (I342776,I342759,I459592);
DFFARX1 I_20004 (I342776,I2683,I342677,I342802,);
not I_20005 (I342810,I342802);
DFFARX1 I_20006 (I459577,I2683,I342677,I342836,);
and I_20007 (I342844,I342836,I459580);
nand I_20008 (I342861,I342836,I459580);
nand I_20009 (I342648,I342810,I342861);
DFFARX1 I_20010 (I459583,I2683,I342677,I342901,);
nor I_20011 (I342909,I342901,I342844);
DFFARX1 I_20012 (I342909,I2683,I342677,I342642,);
nor I_20013 (I342657,I342901,I342802);
nand I_20014 (I342954,I459568,I459574);
and I_20015 (I342971,I342954,I459586);
DFFARX1 I_20016 (I342971,I2683,I342677,I342997,);
nor I_20017 (I342645,I342997,I342901);
not I_20018 (I343019,I342997);
nor I_20019 (I343036,I343019,I342810);
nor I_20020 (I343053,I342742,I343036);
DFFARX1 I_20021 (I343053,I2683,I342677,I342660,);
nor I_20022 (I343084,I343019,I342901);
nor I_20023 (I343101,I459571,I459574);
nor I_20024 (I342651,I343101,I343084);
not I_20025 (I343132,I343101);
nand I_20026 (I342654,I342861,I343132);
DFFARX1 I_20027 (I343101,I2683,I342677,I342666,);
DFFARX1 I_20028 (I343101,I2683,I342677,I342663,);
not I_20029 (I343221,I2690);
DFFARX1 I_20030 (I164049,I2683,I343221,I343247,);
DFFARX1 I_20031 (I343247,I2683,I343221,I343264,);
not I_20032 (I343213,I343264);
not I_20033 (I343286,I343247);
nand I_20034 (I343303,I164061,I164040);
and I_20035 (I343320,I343303,I164043);
DFFARX1 I_20036 (I343320,I2683,I343221,I343346,);
not I_20037 (I343354,I343346);
DFFARX1 I_20038 (I164052,I2683,I343221,I343380,);
and I_20039 (I343388,I343380,I164064);
nand I_20040 (I343405,I343380,I164064);
nand I_20041 (I343192,I343354,I343405);
DFFARX1 I_20042 (I164058,I2683,I343221,I343445,);
nor I_20043 (I343453,I343445,I343388);
DFFARX1 I_20044 (I343453,I2683,I343221,I343186,);
nor I_20045 (I343201,I343445,I343346);
nand I_20046 (I343498,I164046,I164043);
and I_20047 (I343515,I343498,I164055);
DFFARX1 I_20048 (I343515,I2683,I343221,I343541,);
nor I_20049 (I343189,I343541,I343445);
not I_20050 (I343563,I343541);
nor I_20051 (I343580,I343563,I343354);
nor I_20052 (I343597,I343286,I343580);
DFFARX1 I_20053 (I343597,I2683,I343221,I343204,);
nor I_20054 (I343628,I343563,I343445);
nor I_20055 (I343645,I164040,I164043);
nor I_20056 (I343195,I343645,I343628);
not I_20057 (I343676,I343645);
nand I_20058 (I343198,I343405,I343676);
DFFARX1 I_20059 (I343645,I2683,I343221,I343210,);
DFFARX1 I_20060 (I343645,I2683,I343221,I343207,);
not I_20061 (I343765,I2690);
DFFARX1 I_20062 (I584997,I2683,I343765,I343791,);
DFFARX1 I_20063 (I343791,I2683,I343765,I343808,);
not I_20064 (I343757,I343808);
not I_20065 (I343830,I343791);
nand I_20066 (I343847,I585018,I585009);
and I_20067 (I343864,I343847,I584997);
DFFARX1 I_20068 (I343864,I2683,I343765,I343890,);
not I_20069 (I343898,I343890);
DFFARX1 I_20070 (I585003,I2683,I343765,I343924,);
and I_20071 (I343932,I343924,I585000);
nand I_20072 (I343949,I343924,I585000);
nand I_20073 (I343736,I343898,I343949);
DFFARX1 I_20074 (I584994,I2683,I343765,I343989,);
nor I_20075 (I343997,I343989,I343932);
DFFARX1 I_20076 (I343997,I2683,I343765,I343730,);
nor I_20077 (I343745,I343989,I343890);
nand I_20078 (I344042,I584994,I585006);
and I_20079 (I344059,I344042,I585015);
DFFARX1 I_20080 (I344059,I2683,I343765,I344085,);
nor I_20081 (I343733,I344085,I343989);
not I_20082 (I344107,I344085);
nor I_20083 (I344124,I344107,I343898);
nor I_20084 (I344141,I343830,I344124);
DFFARX1 I_20085 (I344141,I2683,I343765,I343748,);
nor I_20086 (I344172,I344107,I343989);
nor I_20087 (I344189,I585012,I585006);
nor I_20088 (I343739,I344189,I344172);
not I_20089 (I344220,I344189);
nand I_20090 (I343742,I343949,I344220);
DFFARX1 I_20091 (I344189,I2683,I343765,I343754,);
DFFARX1 I_20092 (I344189,I2683,I343765,I343751,);
not I_20093 (I344309,I2690);
DFFARX1 I_20094 (I906229,I2683,I344309,I344335,);
DFFARX1 I_20095 (I344335,I2683,I344309,I344352,);
not I_20096 (I344301,I344352);
not I_20097 (I344374,I344335);
nand I_20098 (I344391,I906241,I906229);
and I_20099 (I344408,I344391,I906232);
DFFARX1 I_20100 (I344408,I2683,I344309,I344434,);
not I_20101 (I344442,I344434);
DFFARX1 I_20102 (I906250,I2683,I344309,I344468,);
and I_20103 (I344476,I344468,I906226);
nand I_20104 (I344493,I344468,I906226);
nand I_20105 (I344280,I344442,I344493);
DFFARX1 I_20106 (I906244,I2683,I344309,I344533,);
nor I_20107 (I344541,I344533,I344476);
DFFARX1 I_20108 (I344541,I2683,I344309,I344274,);
nor I_20109 (I344289,I344533,I344434);
nand I_20110 (I344586,I906238,I906235);
and I_20111 (I344603,I344586,I906247);
DFFARX1 I_20112 (I344603,I2683,I344309,I344629,);
nor I_20113 (I344277,I344629,I344533);
not I_20114 (I344651,I344629);
nor I_20115 (I344668,I344651,I344442);
nor I_20116 (I344685,I344374,I344668);
DFFARX1 I_20117 (I344685,I2683,I344309,I344292,);
nor I_20118 (I344716,I344651,I344533);
nor I_20119 (I344733,I906226,I906235);
nor I_20120 (I344283,I344733,I344716);
not I_20121 (I344764,I344733);
nand I_20122 (I344286,I344493,I344764);
DFFARX1 I_20123 (I344733,I2683,I344309,I344298,);
DFFARX1 I_20124 (I344733,I2683,I344309,I344295,);
not I_20125 (I344853,I2690);
DFFARX1 I_20126 (I175354,I2683,I344853,I344879,);
DFFARX1 I_20127 (I344879,I2683,I344853,I344896,);
not I_20128 (I344845,I344896);
not I_20129 (I344918,I344879);
nand I_20130 (I344935,I175366,I175345);
and I_20131 (I344952,I344935,I175348);
DFFARX1 I_20132 (I344952,I2683,I344853,I344978,);
not I_20133 (I344986,I344978);
DFFARX1 I_20134 (I175357,I2683,I344853,I345012,);
and I_20135 (I345020,I345012,I175369);
nand I_20136 (I345037,I345012,I175369);
nand I_20137 (I344824,I344986,I345037);
DFFARX1 I_20138 (I175363,I2683,I344853,I345077,);
nor I_20139 (I345085,I345077,I345020);
DFFARX1 I_20140 (I345085,I2683,I344853,I344818,);
nor I_20141 (I344833,I345077,I344978);
nand I_20142 (I345130,I175351,I175348);
and I_20143 (I345147,I345130,I175360);
DFFARX1 I_20144 (I345147,I2683,I344853,I345173,);
nor I_20145 (I344821,I345173,I345077);
not I_20146 (I345195,I345173);
nor I_20147 (I345212,I345195,I344986);
nor I_20148 (I345229,I344918,I345212);
DFFARX1 I_20149 (I345229,I2683,I344853,I344836,);
nor I_20150 (I345260,I345195,I345077);
nor I_20151 (I345277,I175345,I175348);
nor I_20152 (I344827,I345277,I345260);
not I_20153 (I345308,I345277);
nand I_20154 (I344830,I345037,I345308);
DFFARX1 I_20155 (I345277,I2683,I344853,I344842,);
DFFARX1 I_20156 (I345277,I2683,I344853,I344839,);
not I_20157 (I345397,I2690);
DFFARX1 I_20158 (I195584,I2683,I345397,I345423,);
DFFARX1 I_20159 (I345423,I2683,I345397,I345440,);
not I_20160 (I345389,I345440);
not I_20161 (I345462,I345423);
nand I_20162 (I345479,I195596,I195575);
and I_20163 (I345496,I345479,I195578);
DFFARX1 I_20164 (I345496,I2683,I345397,I345522,);
not I_20165 (I345530,I345522);
DFFARX1 I_20166 (I195587,I2683,I345397,I345556,);
and I_20167 (I345564,I345556,I195599);
nand I_20168 (I345581,I345556,I195599);
nand I_20169 (I345368,I345530,I345581);
DFFARX1 I_20170 (I195593,I2683,I345397,I345621,);
nor I_20171 (I345629,I345621,I345564);
DFFARX1 I_20172 (I345629,I2683,I345397,I345362,);
nor I_20173 (I345377,I345621,I345522);
nand I_20174 (I345674,I195581,I195578);
and I_20175 (I345691,I345674,I195590);
DFFARX1 I_20176 (I345691,I2683,I345397,I345717,);
nor I_20177 (I345365,I345717,I345621);
not I_20178 (I345739,I345717);
nor I_20179 (I345756,I345739,I345530);
nor I_20180 (I345773,I345462,I345756);
DFFARX1 I_20181 (I345773,I2683,I345397,I345380,);
nor I_20182 (I345804,I345739,I345621);
nor I_20183 (I345821,I195575,I195578);
nor I_20184 (I345371,I345821,I345804);
not I_20185 (I345852,I345821);
nand I_20186 (I345374,I345581,I345852);
DFFARX1 I_20187 (I345821,I2683,I345397,I345386,);
DFFARX1 I_20188 (I345821,I2683,I345397,I345383,);
not I_20189 (I345941,I2690);
DFFARX1 I_20190 (I942643,I2683,I345941,I345967,);
DFFARX1 I_20191 (I345967,I2683,I345941,I345984,);
not I_20192 (I345933,I345984);
not I_20193 (I346006,I345967);
nand I_20194 (I346023,I942655,I942643);
and I_20195 (I346040,I346023,I942646);
DFFARX1 I_20196 (I346040,I2683,I345941,I346066,);
not I_20197 (I346074,I346066);
DFFARX1 I_20198 (I942664,I2683,I345941,I346100,);
and I_20199 (I346108,I346100,I942640);
nand I_20200 (I346125,I346100,I942640);
nand I_20201 (I345912,I346074,I346125);
DFFARX1 I_20202 (I942658,I2683,I345941,I346165,);
nor I_20203 (I346173,I346165,I346108);
DFFARX1 I_20204 (I346173,I2683,I345941,I345906,);
nor I_20205 (I345921,I346165,I346066);
nand I_20206 (I346218,I942652,I942649);
and I_20207 (I346235,I346218,I942661);
DFFARX1 I_20208 (I346235,I2683,I345941,I346261,);
nor I_20209 (I345909,I346261,I346165);
not I_20210 (I346283,I346261);
nor I_20211 (I346300,I346283,I346074);
nor I_20212 (I346317,I346006,I346300);
DFFARX1 I_20213 (I346317,I2683,I345941,I345924,);
nor I_20214 (I346348,I346283,I346165);
nor I_20215 (I346365,I942640,I942649);
nor I_20216 (I345915,I346365,I346348);
not I_20217 (I346396,I346365);
nand I_20218 (I345918,I346125,I346396);
DFFARX1 I_20219 (I346365,I2683,I345941,I345930,);
DFFARX1 I_20220 (I346365,I2683,I345941,I345927,);
not I_20221 (I346485,I2690);
DFFARX1 I_20222 (I2460,I2683,I346485,I346511,);
DFFARX1 I_20223 (I346511,I2683,I346485,I346528,);
not I_20224 (I346477,I346528);
not I_20225 (I346550,I346511);
nand I_20226 (I346567,I2540,I2268);
and I_20227 (I346584,I346567,I1732);
DFFARX1 I_20228 (I346584,I2683,I346485,I346610,);
not I_20229 (I346618,I346610);
DFFARX1 I_20230 (I1428,I2683,I346485,I346644,);
and I_20231 (I346652,I346644,I1364);
nand I_20232 (I346669,I346644,I1364);
nand I_20233 (I346456,I346618,I346669);
DFFARX1 I_20234 (I1612,I2683,I346485,I346709,);
nor I_20235 (I346717,I346709,I346652);
DFFARX1 I_20236 (I346717,I2683,I346485,I346450,);
nor I_20237 (I346465,I346709,I346610);
nand I_20238 (I346762,I1892,I2556);
and I_20239 (I346779,I346762,I2452);
DFFARX1 I_20240 (I346779,I2683,I346485,I346805,);
nor I_20241 (I346453,I346805,I346709);
not I_20242 (I346827,I346805);
nor I_20243 (I346844,I346827,I346618);
nor I_20244 (I346861,I346550,I346844);
DFFARX1 I_20245 (I346861,I2683,I346485,I346468,);
nor I_20246 (I346892,I346827,I346709);
nor I_20247 (I346909,I2420,I2556);
nor I_20248 (I346459,I346909,I346892);
not I_20249 (I346940,I346909);
nand I_20250 (I346462,I346669,I346940);
DFFARX1 I_20251 (I346909,I2683,I346485,I346474,);
DFFARX1 I_20252 (I346909,I2683,I346485,I346471,);
not I_20253 (I347029,I2690);
DFFARX1 I_20254 (I557831,I2683,I347029,I347055,);
DFFARX1 I_20255 (I347055,I2683,I347029,I347072,);
not I_20256 (I347021,I347072);
not I_20257 (I347094,I347055);
nand I_20258 (I347111,I557852,I557843);
and I_20259 (I347128,I347111,I557831);
DFFARX1 I_20260 (I347128,I2683,I347029,I347154,);
not I_20261 (I347162,I347154);
DFFARX1 I_20262 (I557837,I2683,I347029,I347188,);
and I_20263 (I347196,I347188,I557834);
nand I_20264 (I347213,I347188,I557834);
nand I_20265 (I347000,I347162,I347213);
DFFARX1 I_20266 (I557828,I2683,I347029,I347253,);
nor I_20267 (I347261,I347253,I347196);
DFFARX1 I_20268 (I347261,I2683,I347029,I346994,);
nor I_20269 (I347009,I347253,I347154);
nand I_20270 (I347306,I557828,I557840);
and I_20271 (I347323,I347306,I557849);
DFFARX1 I_20272 (I347323,I2683,I347029,I347349,);
nor I_20273 (I346997,I347349,I347253);
not I_20274 (I347371,I347349);
nor I_20275 (I347388,I347371,I347162);
nor I_20276 (I347405,I347094,I347388);
DFFARX1 I_20277 (I347405,I2683,I347029,I347012,);
nor I_20278 (I347436,I347371,I347253);
nor I_20279 (I347453,I557846,I557840);
nor I_20280 (I347003,I347453,I347436);
not I_20281 (I347484,I347453);
nand I_20282 (I347006,I347213,I347484);
DFFARX1 I_20283 (I347453,I2683,I347029,I347018,);
DFFARX1 I_20284 (I347453,I2683,I347029,I347015,);
not I_20285 (I347573,I2690);
DFFARX1 I_20286 (I538757,I2683,I347573,I347599,);
DFFARX1 I_20287 (I347599,I2683,I347573,I347616,);
not I_20288 (I347565,I347616);
not I_20289 (I347638,I347599);
nand I_20290 (I347655,I538778,I538769);
and I_20291 (I347672,I347655,I538757);
DFFARX1 I_20292 (I347672,I2683,I347573,I347698,);
not I_20293 (I347706,I347698);
DFFARX1 I_20294 (I538763,I2683,I347573,I347732,);
and I_20295 (I347740,I347732,I538760);
nand I_20296 (I347757,I347732,I538760);
nand I_20297 (I347544,I347706,I347757);
DFFARX1 I_20298 (I538754,I2683,I347573,I347797,);
nor I_20299 (I347805,I347797,I347740);
DFFARX1 I_20300 (I347805,I2683,I347573,I347538,);
nor I_20301 (I347553,I347797,I347698);
nand I_20302 (I347850,I538754,I538766);
and I_20303 (I347867,I347850,I538775);
DFFARX1 I_20304 (I347867,I2683,I347573,I347893,);
nor I_20305 (I347541,I347893,I347797);
not I_20306 (I347915,I347893);
nor I_20307 (I347932,I347915,I347706);
nor I_20308 (I347949,I347638,I347932);
DFFARX1 I_20309 (I347949,I2683,I347573,I347556,);
nor I_20310 (I347980,I347915,I347797);
nor I_20311 (I347997,I538772,I538766);
nor I_20312 (I347547,I347997,I347980);
not I_20313 (I348028,I347997);
nand I_20314 (I347550,I347757,I348028);
DFFARX1 I_20315 (I347997,I2683,I347573,I347562,);
DFFARX1 I_20316 (I347997,I2683,I347573,I347559,);
not I_20317 (I348117,I2690);
DFFARX1 I_20318 (I766509,I2683,I348117,I348143,);
DFFARX1 I_20319 (I348143,I2683,I348117,I348160,);
not I_20320 (I348109,I348160);
not I_20321 (I348182,I348143);
nand I_20322 (I348199,I766524,I766512);
and I_20323 (I348216,I348199,I766503);
DFFARX1 I_20324 (I348216,I2683,I348117,I348242,);
not I_20325 (I348250,I348242);
DFFARX1 I_20326 (I766515,I2683,I348117,I348276,);
and I_20327 (I348284,I348276,I766506);
nand I_20328 (I348301,I348276,I766506);
nand I_20329 (I348088,I348250,I348301);
DFFARX1 I_20330 (I766521,I2683,I348117,I348341,);
nor I_20331 (I348349,I348341,I348284);
DFFARX1 I_20332 (I348349,I2683,I348117,I348082,);
nor I_20333 (I348097,I348341,I348242);
nand I_20334 (I348394,I766530,I766518);
and I_20335 (I348411,I348394,I766527);
DFFARX1 I_20336 (I348411,I2683,I348117,I348437,);
nor I_20337 (I348085,I348437,I348341);
not I_20338 (I348459,I348437);
nor I_20339 (I348476,I348459,I348250);
nor I_20340 (I348493,I348182,I348476);
DFFARX1 I_20341 (I348493,I2683,I348117,I348100,);
nor I_20342 (I348524,I348459,I348341);
nor I_20343 (I348541,I766503,I766518);
nor I_20344 (I348091,I348541,I348524);
not I_20345 (I348572,I348541);
nand I_20346 (I348094,I348301,I348572);
DFFARX1 I_20347 (I348541,I2683,I348117,I348106,);
DFFARX1 I_20348 (I348541,I2683,I348117,I348103,);
not I_20349 (I348661,I2690);
DFFARX1 I_20350 (I655998,I2683,I348661,I348687,);
DFFARX1 I_20351 (I348687,I2683,I348661,I348704,);
not I_20352 (I348653,I348704);
not I_20353 (I348726,I348687);
nand I_20354 (I348743,I655992,I655989);
and I_20355 (I348760,I348743,I656004);
DFFARX1 I_20356 (I348760,I2683,I348661,I348786,);
not I_20357 (I348794,I348786);
DFFARX1 I_20358 (I655992,I2683,I348661,I348820,);
and I_20359 (I348828,I348820,I655986);
nand I_20360 (I348845,I348820,I655986);
nand I_20361 (I348632,I348794,I348845);
DFFARX1 I_20362 (I655986,I2683,I348661,I348885,);
nor I_20363 (I348893,I348885,I348828);
DFFARX1 I_20364 (I348893,I2683,I348661,I348626,);
nor I_20365 (I348641,I348885,I348786);
nand I_20366 (I348938,I656001,I655995);
and I_20367 (I348955,I348938,I655989);
DFFARX1 I_20368 (I348955,I2683,I348661,I348981,);
nor I_20369 (I348629,I348981,I348885);
not I_20370 (I349003,I348981);
nor I_20371 (I349020,I349003,I348794);
nor I_20372 (I349037,I348726,I349020);
DFFARX1 I_20373 (I349037,I2683,I348661,I348644,);
nor I_20374 (I349068,I349003,I348885);
nor I_20375 (I349085,I656007,I655995);
nor I_20376 (I348635,I349085,I349068);
not I_20377 (I349116,I349085);
nand I_20378 (I348638,I348845,I349116);
DFFARX1 I_20379 (I349085,I2683,I348661,I348650,);
DFFARX1 I_20380 (I349085,I2683,I348661,I348647,);
not I_20381 (I349205,I2690);
DFFARX1 I_20382 (I213242,I2683,I349205,I349231,);
DFFARX1 I_20383 (I349231,I2683,I349205,I349248,);
not I_20384 (I349197,I349248);
not I_20385 (I349270,I349231);
nand I_20386 (I349287,I213221,I213245);
and I_20387 (I349304,I349287,I213248);
DFFARX1 I_20388 (I349304,I2683,I349205,I349330,);
not I_20389 (I349338,I349330);
DFFARX1 I_20390 (I213230,I2683,I349205,I349364,);
and I_20391 (I349372,I349364,I213236);
nand I_20392 (I349389,I349364,I213236);
nand I_20393 (I349176,I349338,I349389);
DFFARX1 I_20394 (I213224,I2683,I349205,I349429,);
nor I_20395 (I349437,I349429,I349372);
DFFARX1 I_20396 (I349437,I2683,I349205,I349170,);
nor I_20397 (I349185,I349429,I349330);
nand I_20398 (I349482,I213233,I213221);
and I_20399 (I349499,I349482,I213227);
DFFARX1 I_20400 (I349499,I2683,I349205,I349525,);
nor I_20401 (I349173,I349525,I349429);
not I_20402 (I349547,I349525);
nor I_20403 (I349564,I349547,I349338);
nor I_20404 (I349581,I349270,I349564);
DFFARX1 I_20405 (I349581,I2683,I349205,I349188,);
nor I_20406 (I349612,I349547,I349429);
nor I_20407 (I349629,I213239,I213221);
nor I_20408 (I349179,I349629,I349612);
not I_20409 (I349660,I349629);
nand I_20410 (I349182,I349389,I349660);
DFFARX1 I_20411 (I349629,I2683,I349205,I349194,);
DFFARX1 I_20412 (I349629,I2683,I349205,I349191,);
not I_20413 (I349749,I2690);
DFFARX1 I_20414 (I779429,I2683,I349749,I349775,);
DFFARX1 I_20415 (I349775,I2683,I349749,I349792,);
not I_20416 (I349741,I349792);
not I_20417 (I349814,I349775);
nand I_20418 (I349831,I779444,I779432);
and I_20419 (I349848,I349831,I779423);
DFFARX1 I_20420 (I349848,I2683,I349749,I349874,);
not I_20421 (I349882,I349874);
DFFARX1 I_20422 (I779435,I2683,I349749,I349908,);
and I_20423 (I349916,I349908,I779426);
nand I_20424 (I349933,I349908,I779426);
nand I_20425 (I349720,I349882,I349933);
DFFARX1 I_20426 (I779441,I2683,I349749,I349973,);
nor I_20427 (I349981,I349973,I349916);
DFFARX1 I_20428 (I349981,I2683,I349749,I349714,);
nor I_20429 (I349729,I349973,I349874);
nand I_20430 (I350026,I779450,I779438);
and I_20431 (I350043,I350026,I779447);
DFFARX1 I_20432 (I350043,I2683,I349749,I350069,);
nor I_20433 (I349717,I350069,I349973);
not I_20434 (I350091,I350069);
nor I_20435 (I350108,I350091,I349882);
nor I_20436 (I350125,I349814,I350108);
DFFARX1 I_20437 (I350125,I2683,I349749,I349732,);
nor I_20438 (I350156,I350091,I349973);
nor I_20439 (I350173,I779423,I779438);
nor I_20440 (I349723,I350173,I350156);
not I_20441 (I350204,I350173);
nand I_20442 (I349726,I349933,I350204);
DFFARX1 I_20443 (I350173,I2683,I349749,I349738,);
DFFARX1 I_20444 (I350173,I2683,I349749,I349735,);
not I_20445 (I350293,I2690);
DFFARX1 I_20446 (I143819,I2683,I350293,I350319,);
DFFARX1 I_20447 (I350319,I2683,I350293,I350336,);
not I_20448 (I350285,I350336);
not I_20449 (I350358,I350319);
nand I_20450 (I350375,I143831,I143810);
and I_20451 (I350392,I350375,I143813);
DFFARX1 I_20452 (I350392,I2683,I350293,I350418,);
not I_20453 (I350426,I350418);
DFFARX1 I_20454 (I143822,I2683,I350293,I350452,);
and I_20455 (I350460,I350452,I143834);
nand I_20456 (I350477,I350452,I143834);
nand I_20457 (I350264,I350426,I350477);
DFFARX1 I_20458 (I143828,I2683,I350293,I350517,);
nor I_20459 (I350525,I350517,I350460);
DFFARX1 I_20460 (I350525,I2683,I350293,I350258,);
nor I_20461 (I350273,I350517,I350418);
nand I_20462 (I350570,I143816,I143813);
and I_20463 (I350587,I350570,I143825);
DFFARX1 I_20464 (I350587,I2683,I350293,I350613,);
nor I_20465 (I350261,I350613,I350517);
not I_20466 (I350635,I350613);
nor I_20467 (I350652,I350635,I350426);
nor I_20468 (I350669,I350358,I350652);
DFFARX1 I_20469 (I350669,I2683,I350293,I350276,);
nor I_20470 (I350700,I350635,I350517);
nor I_20471 (I350717,I143810,I143813);
nor I_20472 (I350267,I350717,I350700);
not I_20473 (I350748,I350717);
nand I_20474 (I350270,I350477,I350748);
DFFARX1 I_20475 (I350717,I2683,I350293,I350282,);
DFFARX1 I_20476 (I350717,I2683,I350293,I350279,);
not I_20477 (I350837,I2690);
DFFARX1 I_20478 (I315480,I2683,I350837,I350863,);
DFFARX1 I_20479 (I350863,I2683,I350837,I350880,);
not I_20480 (I350829,I350880);
not I_20481 (I350902,I350863);
nand I_20482 (I350919,I315459,I315483);
and I_20483 (I350936,I350919,I315486);
DFFARX1 I_20484 (I350936,I2683,I350837,I350962,);
not I_20485 (I350970,I350962);
DFFARX1 I_20486 (I315468,I2683,I350837,I350996,);
and I_20487 (I351004,I350996,I315474);
nand I_20488 (I351021,I350996,I315474);
nand I_20489 (I350808,I350970,I351021);
DFFARX1 I_20490 (I315462,I2683,I350837,I351061,);
nor I_20491 (I351069,I351061,I351004);
DFFARX1 I_20492 (I351069,I2683,I350837,I350802,);
nor I_20493 (I350817,I351061,I350962);
nand I_20494 (I351114,I315471,I315459);
and I_20495 (I351131,I351114,I315465);
DFFARX1 I_20496 (I351131,I2683,I350837,I351157,);
nor I_20497 (I350805,I351157,I351061);
not I_20498 (I351179,I351157);
nor I_20499 (I351196,I351179,I350970);
nor I_20500 (I351213,I350902,I351196);
DFFARX1 I_20501 (I351213,I2683,I350837,I350820,);
nor I_20502 (I351244,I351179,I351061);
nor I_20503 (I351261,I315477,I315459);
nor I_20504 (I350811,I351261,I351244);
not I_20505 (I351292,I351261);
nand I_20506 (I350814,I351021,I351292);
DFFARX1 I_20507 (I351261,I2683,I350837,I350826,);
DFFARX1 I_20508 (I351261,I2683,I350837,I350823,);
not I_20509 (I351381,I2690);
DFFARX1 I_20510 (I37980,I2683,I351381,I351407,);
DFFARX1 I_20511 (I351407,I2683,I351381,I351424,);
not I_20512 (I351373,I351424);
not I_20513 (I351446,I351407);
nand I_20514 (I351463,I37968,I37983);
and I_20515 (I351480,I351463,I37971);
DFFARX1 I_20516 (I351480,I2683,I351381,I351506,);
not I_20517 (I351514,I351506);
DFFARX1 I_20518 (I37992,I2683,I351381,I351540,);
and I_20519 (I351548,I351540,I37986);
nand I_20520 (I351565,I351540,I37986);
nand I_20521 (I351352,I351514,I351565);
DFFARX1 I_20522 (I37989,I2683,I351381,I351605,);
nor I_20523 (I351613,I351605,I351548);
DFFARX1 I_20524 (I351613,I2683,I351381,I351346,);
nor I_20525 (I351361,I351605,I351506);
nand I_20526 (I351658,I37968,I37971);
and I_20527 (I351675,I351658,I37974);
DFFARX1 I_20528 (I351675,I2683,I351381,I351701,);
nor I_20529 (I351349,I351701,I351605);
not I_20530 (I351723,I351701);
nor I_20531 (I351740,I351723,I351514);
nor I_20532 (I351757,I351446,I351740);
DFFARX1 I_20533 (I351757,I2683,I351381,I351364,);
nor I_20534 (I351788,I351723,I351605);
nor I_20535 (I351805,I37977,I37971);
nor I_20536 (I351355,I351805,I351788);
not I_20537 (I351836,I351805);
nand I_20538 (I351358,I351565,I351836);
DFFARX1 I_20539 (I351805,I2683,I351381,I351370,);
DFFARX1 I_20540 (I351805,I2683,I351381,I351367,);
not I_20541 (I351925,I2690);
DFFARX1 I_20542 (I836291,I2683,I351925,I351951,);
DFFARX1 I_20543 (I351951,I2683,I351925,I351968,);
not I_20544 (I351917,I351968);
not I_20545 (I351990,I351951);
nand I_20546 (I352007,I836303,I836291);
and I_20547 (I352024,I352007,I836294);
DFFARX1 I_20548 (I352024,I2683,I351925,I352050,);
not I_20549 (I352058,I352050);
DFFARX1 I_20550 (I836312,I2683,I351925,I352084,);
and I_20551 (I352092,I352084,I836288);
nand I_20552 (I352109,I352084,I836288);
nand I_20553 (I351896,I352058,I352109);
DFFARX1 I_20554 (I836306,I2683,I351925,I352149,);
nor I_20555 (I352157,I352149,I352092);
DFFARX1 I_20556 (I352157,I2683,I351925,I351890,);
nor I_20557 (I351905,I352149,I352050);
nand I_20558 (I352202,I836300,I836297);
and I_20559 (I352219,I352202,I836309);
DFFARX1 I_20560 (I352219,I2683,I351925,I352245,);
nor I_20561 (I351893,I352245,I352149);
not I_20562 (I352267,I352245);
nor I_20563 (I352284,I352267,I352058);
nor I_20564 (I352301,I351990,I352284);
DFFARX1 I_20565 (I352301,I2683,I351925,I351908,);
nor I_20566 (I352332,I352267,I352149);
nor I_20567 (I352349,I836288,I836297);
nor I_20568 (I351899,I352349,I352332);
not I_20569 (I352380,I352349);
nand I_20570 (I351902,I352109,I352380);
DFFARX1 I_20571 (I352349,I2683,I351925,I351914,);
DFFARX1 I_20572 (I352349,I2683,I351925,I351911,);
not I_20573 (I352469,I2690);
DFFARX1 I_20574 (I625432,I2683,I352469,I352495,);
DFFARX1 I_20575 (I352495,I2683,I352469,I352512,);
not I_20576 (I352461,I352512);
not I_20577 (I352534,I352495);
nand I_20578 (I352551,I625426,I625423);
and I_20579 (I352568,I352551,I625438);
DFFARX1 I_20580 (I352568,I2683,I352469,I352594,);
not I_20581 (I352602,I352594);
DFFARX1 I_20582 (I625426,I2683,I352469,I352628,);
and I_20583 (I352636,I352628,I625420);
nand I_20584 (I352653,I352628,I625420);
nand I_20585 (I352440,I352602,I352653);
DFFARX1 I_20586 (I625420,I2683,I352469,I352693,);
nor I_20587 (I352701,I352693,I352636);
DFFARX1 I_20588 (I352701,I2683,I352469,I352434,);
nor I_20589 (I352449,I352693,I352594);
nand I_20590 (I352746,I625435,I625429);
and I_20591 (I352763,I352746,I625423);
DFFARX1 I_20592 (I352763,I2683,I352469,I352789,);
nor I_20593 (I352437,I352789,I352693);
not I_20594 (I352811,I352789);
nor I_20595 (I352828,I352811,I352602);
nor I_20596 (I352845,I352534,I352828);
DFFARX1 I_20597 (I352845,I2683,I352469,I352452,);
nor I_20598 (I352876,I352811,I352693);
nor I_20599 (I352893,I625441,I625429);
nor I_20600 (I352443,I352893,I352876);
not I_20601 (I352924,I352893);
nand I_20602 (I352446,I352653,I352924);
DFFARX1 I_20603 (I352893,I2683,I352469,I352458,);
DFFARX1 I_20604 (I352893,I2683,I352469,I352455,);
not I_20605 (I353013,I2690);
DFFARX1 I_20606 (I55892,I2683,I353013,I353039,);
DFFARX1 I_20607 (I353039,I2683,I353013,I353056,);
not I_20608 (I353005,I353056);
not I_20609 (I353078,I353039);
nand I_20610 (I353095,I55907,I55886);
and I_20611 (I353112,I353095,I55889);
DFFARX1 I_20612 (I353112,I2683,I353013,I353138,);
not I_20613 (I353146,I353138);
DFFARX1 I_20614 (I55895,I2683,I353013,I353172,);
and I_20615 (I353180,I353172,I55889);
nand I_20616 (I353197,I353172,I55889);
nand I_20617 (I352984,I353146,I353197);
DFFARX1 I_20618 (I55904,I2683,I353013,I353237,);
nor I_20619 (I353245,I353237,I353180);
DFFARX1 I_20620 (I353245,I2683,I353013,I352978,);
nor I_20621 (I352993,I353237,I353138);
nand I_20622 (I353290,I55886,I55901);
and I_20623 (I353307,I353290,I55898);
DFFARX1 I_20624 (I353307,I2683,I353013,I353333,);
nor I_20625 (I352981,I353333,I353237);
not I_20626 (I353355,I353333);
nor I_20627 (I353372,I353355,I353146);
nor I_20628 (I353389,I353078,I353372);
DFFARX1 I_20629 (I353389,I2683,I353013,I352996,);
nor I_20630 (I353420,I353355,I353237);
nor I_20631 (I353437,I55910,I55901);
nor I_20632 (I352987,I353437,I353420);
not I_20633 (I353468,I353437);
nand I_20634 (I352990,I353197,I353468);
DFFARX1 I_20635 (I353437,I2683,I353013,I353002,);
DFFARX1 I_20636 (I353437,I2683,I353013,I352999,);
not I_20637 (I353557,I2690);
DFFARX1 I_20638 (I632810,I2683,I353557,I353583,);
DFFARX1 I_20639 (I353583,I2683,I353557,I353600,);
not I_20640 (I353549,I353600);
not I_20641 (I353622,I353583);
nand I_20642 (I353639,I632804,I632801);
and I_20643 (I353656,I353639,I632816);
DFFARX1 I_20644 (I353656,I2683,I353557,I353682,);
not I_20645 (I353690,I353682);
DFFARX1 I_20646 (I632804,I2683,I353557,I353716,);
and I_20647 (I353724,I353716,I632798);
nand I_20648 (I353741,I353716,I632798);
nand I_20649 (I353528,I353690,I353741);
DFFARX1 I_20650 (I632798,I2683,I353557,I353781,);
nor I_20651 (I353789,I353781,I353724);
DFFARX1 I_20652 (I353789,I2683,I353557,I353522,);
nor I_20653 (I353537,I353781,I353682);
nand I_20654 (I353834,I632813,I632807);
and I_20655 (I353851,I353834,I632801);
DFFARX1 I_20656 (I353851,I2683,I353557,I353877,);
nor I_20657 (I353525,I353877,I353781);
not I_20658 (I353899,I353877);
nor I_20659 (I353916,I353899,I353690);
nor I_20660 (I353933,I353622,I353916);
DFFARX1 I_20661 (I353933,I2683,I353557,I353540,);
nor I_20662 (I353964,I353899,I353781);
nor I_20663 (I353981,I632819,I632807);
nor I_20664 (I353531,I353981,I353964);
not I_20665 (I354012,I353981);
nand I_20666 (I353534,I353741,I354012);
DFFARX1 I_20667 (I353981,I2683,I353557,I353546,);
DFFARX1 I_20668 (I353981,I2683,I353557,I353543,);
not I_20669 (I354101,I2690);
DFFARX1 I_20670 (I710953,I2683,I354101,I354127,);
DFFARX1 I_20671 (I354127,I2683,I354101,I354144,);
not I_20672 (I354093,I354144);
not I_20673 (I354166,I354127);
nand I_20674 (I354183,I710968,I710956);
and I_20675 (I354200,I354183,I710947);
DFFARX1 I_20676 (I354200,I2683,I354101,I354226,);
not I_20677 (I354234,I354226);
DFFARX1 I_20678 (I710959,I2683,I354101,I354260,);
and I_20679 (I354268,I354260,I710950);
nand I_20680 (I354285,I354260,I710950);
nand I_20681 (I354072,I354234,I354285);
DFFARX1 I_20682 (I710965,I2683,I354101,I354325,);
nor I_20683 (I354333,I354325,I354268);
DFFARX1 I_20684 (I354333,I2683,I354101,I354066,);
nor I_20685 (I354081,I354325,I354226);
nand I_20686 (I354378,I710974,I710962);
and I_20687 (I354395,I354378,I710971);
DFFARX1 I_20688 (I354395,I2683,I354101,I354421,);
nor I_20689 (I354069,I354421,I354325);
not I_20690 (I354443,I354421);
nor I_20691 (I354460,I354443,I354234);
nor I_20692 (I354477,I354166,I354460);
DFFARX1 I_20693 (I354477,I2683,I354101,I354084,);
nor I_20694 (I354508,I354443,I354325);
nor I_20695 (I354525,I710947,I710962);
nor I_20696 (I354075,I354525,I354508);
not I_20697 (I354556,I354525);
nand I_20698 (I354078,I354285,I354556);
DFFARX1 I_20699 (I354525,I2683,I354101,I354090,);
DFFARX1 I_20700 (I354525,I2683,I354101,I354087,);
not I_20701 (I354645,I2690);
DFFARX1 I_20702 (I136679,I2683,I354645,I354671,);
DFFARX1 I_20703 (I354671,I2683,I354645,I354688,);
not I_20704 (I354637,I354688);
not I_20705 (I354710,I354671);
nand I_20706 (I354727,I136691,I136670);
and I_20707 (I354744,I354727,I136673);
DFFARX1 I_20708 (I354744,I2683,I354645,I354770,);
not I_20709 (I354778,I354770);
DFFARX1 I_20710 (I136682,I2683,I354645,I354804,);
and I_20711 (I354812,I354804,I136694);
nand I_20712 (I354829,I354804,I136694);
nand I_20713 (I354616,I354778,I354829);
DFFARX1 I_20714 (I136688,I2683,I354645,I354869,);
nor I_20715 (I354877,I354869,I354812);
DFFARX1 I_20716 (I354877,I2683,I354645,I354610,);
nor I_20717 (I354625,I354869,I354770);
nand I_20718 (I354922,I136676,I136673);
and I_20719 (I354939,I354922,I136685);
DFFARX1 I_20720 (I354939,I2683,I354645,I354965,);
nor I_20721 (I354613,I354965,I354869);
not I_20722 (I354987,I354965);
nor I_20723 (I355004,I354987,I354778);
nor I_20724 (I355021,I354710,I355004);
DFFARX1 I_20725 (I355021,I2683,I354645,I354628,);
nor I_20726 (I355052,I354987,I354869);
nor I_20727 (I355069,I136670,I136673);
nor I_20728 (I354619,I355069,I355052);
not I_20729 (I355100,I355069);
nand I_20730 (I354622,I354829,I355100);
DFFARX1 I_20731 (I355069,I2683,I354645,I354634,);
DFFARX1 I_20732 (I355069,I2683,I354645,I354631,);
not I_20733 (I355189,I2690);
DFFARX1 I_20734 (I907963,I2683,I355189,I355215,);
DFFARX1 I_20735 (I355215,I2683,I355189,I355232,);
not I_20736 (I355181,I355232);
not I_20737 (I355254,I355215);
nand I_20738 (I355271,I907975,I907963);
and I_20739 (I355288,I355271,I907966);
DFFARX1 I_20740 (I355288,I2683,I355189,I355314,);
not I_20741 (I355322,I355314);
DFFARX1 I_20742 (I907984,I2683,I355189,I355348,);
and I_20743 (I355356,I355348,I907960);
nand I_20744 (I355373,I355348,I907960);
nand I_20745 (I355160,I355322,I355373);
DFFARX1 I_20746 (I907978,I2683,I355189,I355413,);
nor I_20747 (I355421,I355413,I355356);
DFFARX1 I_20748 (I355421,I2683,I355189,I355154,);
nor I_20749 (I355169,I355413,I355314);
nand I_20750 (I355466,I907972,I907969);
and I_20751 (I355483,I355466,I907981);
DFFARX1 I_20752 (I355483,I2683,I355189,I355509,);
nor I_20753 (I355157,I355509,I355413);
not I_20754 (I355531,I355509);
nor I_20755 (I355548,I355531,I355322);
nor I_20756 (I355565,I355254,I355548);
DFFARX1 I_20757 (I355565,I2683,I355189,I355172,);
nor I_20758 (I355596,I355531,I355413);
nor I_20759 (I355613,I907960,I907969);
nor I_20760 (I355163,I355613,I355596);
not I_20761 (I355644,I355613);
nand I_20762 (I355166,I355373,I355644);
DFFARX1 I_20763 (I355613,I2683,I355189,I355178,);
DFFARX1 I_20764 (I355613,I2683,I355189,I355175,);
not I_20765 (I355733,I2690);
DFFARX1 I_20766 (I710307,I2683,I355733,I355759,);
DFFARX1 I_20767 (I355759,I2683,I355733,I355776,);
not I_20768 (I355725,I355776);
not I_20769 (I355798,I355759);
nand I_20770 (I355815,I710322,I710310);
and I_20771 (I355832,I355815,I710301);
DFFARX1 I_20772 (I355832,I2683,I355733,I355858,);
not I_20773 (I355866,I355858);
DFFARX1 I_20774 (I710313,I2683,I355733,I355892,);
and I_20775 (I355900,I355892,I710304);
nand I_20776 (I355917,I355892,I710304);
nand I_20777 (I355704,I355866,I355917);
DFFARX1 I_20778 (I710319,I2683,I355733,I355957,);
nor I_20779 (I355965,I355957,I355900);
DFFARX1 I_20780 (I355965,I2683,I355733,I355698,);
nor I_20781 (I355713,I355957,I355858);
nand I_20782 (I356010,I710328,I710316);
and I_20783 (I356027,I356010,I710325);
DFFARX1 I_20784 (I356027,I2683,I355733,I356053,);
nor I_20785 (I355701,I356053,I355957);
not I_20786 (I356075,I356053);
nor I_20787 (I356092,I356075,I355866);
nor I_20788 (I356109,I355798,I356092);
DFFARX1 I_20789 (I356109,I2683,I355733,I355716,);
nor I_20790 (I356140,I356075,I355957);
nor I_20791 (I356157,I710301,I710316);
nor I_20792 (I355707,I356157,I356140);
not I_20793 (I356188,I356157);
nand I_20794 (I355710,I355917,I356188);
DFFARX1 I_20795 (I356157,I2683,I355733,I355722,);
DFFARX1 I_20796 (I356157,I2683,I355733,I355719,);
not I_20797 (I356277,I2690);
DFFARX1 I_20798 (I220093,I2683,I356277,I356303,);
DFFARX1 I_20799 (I356303,I2683,I356277,I356320,);
not I_20800 (I356269,I356320);
not I_20801 (I356342,I356303);
nand I_20802 (I356359,I220072,I220096);
and I_20803 (I356376,I356359,I220099);
DFFARX1 I_20804 (I356376,I2683,I356277,I356402,);
not I_20805 (I356410,I356402);
DFFARX1 I_20806 (I220081,I2683,I356277,I356436,);
and I_20807 (I356444,I356436,I220087);
nand I_20808 (I356461,I356436,I220087);
nand I_20809 (I356248,I356410,I356461);
DFFARX1 I_20810 (I220075,I2683,I356277,I356501,);
nor I_20811 (I356509,I356501,I356444);
DFFARX1 I_20812 (I356509,I2683,I356277,I356242,);
nor I_20813 (I356257,I356501,I356402);
nand I_20814 (I356554,I220084,I220072);
and I_20815 (I356571,I356554,I220078);
DFFARX1 I_20816 (I356571,I2683,I356277,I356597,);
nor I_20817 (I356245,I356597,I356501);
not I_20818 (I356619,I356597);
nor I_20819 (I356636,I356619,I356410);
nor I_20820 (I356653,I356342,I356636);
DFFARX1 I_20821 (I356653,I2683,I356277,I356260,);
nor I_20822 (I356684,I356619,I356501);
nor I_20823 (I356701,I220090,I220072);
nor I_20824 (I356251,I356701,I356684);
not I_20825 (I356732,I356701);
nand I_20826 (I356254,I356461,I356732);
DFFARX1 I_20827 (I356701,I2683,I356277,I356266,);
DFFARX1 I_20828 (I356701,I2683,I356277,I356263,);
not I_20829 (I356821,I2690);
DFFARX1 I_20830 (I1093576,I2683,I356821,I356847,);
DFFARX1 I_20831 (I356847,I2683,I356821,I356864,);
not I_20832 (I356813,I356864);
not I_20833 (I356886,I356847);
nand I_20834 (I356903,I1093552,I1093573);
and I_20835 (I356920,I356903,I1093570);
DFFARX1 I_20836 (I356920,I2683,I356821,I356946,);
not I_20837 (I356954,I356946);
DFFARX1 I_20838 (I1093549,I2683,I356821,I356980,);
and I_20839 (I356988,I356980,I1093561);
nand I_20840 (I357005,I356980,I1093561);
nand I_20841 (I356792,I356954,I357005);
DFFARX1 I_20842 (I1093564,I2683,I356821,I357045,);
nor I_20843 (I357053,I357045,I356988);
DFFARX1 I_20844 (I357053,I2683,I356821,I356786,);
nor I_20845 (I356801,I357045,I356946);
nand I_20846 (I357098,I1093567,I1093555);
and I_20847 (I357115,I357098,I1093558);
DFFARX1 I_20848 (I357115,I2683,I356821,I357141,);
nor I_20849 (I356789,I357141,I357045);
not I_20850 (I357163,I357141);
nor I_20851 (I357180,I357163,I356954);
nor I_20852 (I357197,I356886,I357180);
DFFARX1 I_20853 (I357197,I2683,I356821,I356804,);
nor I_20854 (I357228,I357163,I357045);
nor I_20855 (I357245,I1093549,I1093555);
nor I_20856 (I356795,I357245,I357228);
not I_20857 (I357276,I357245);
nand I_20858 (I356798,I357005,I357276);
DFFARX1 I_20859 (I357245,I2683,I356821,I356810,);
DFFARX1 I_20860 (I357245,I2683,I356821,I356807,);
not I_20861 (I357365,I2690);
DFFARX1 I_20862 (I838603,I2683,I357365,I357391,);
DFFARX1 I_20863 (I357391,I2683,I357365,I357408,);
not I_20864 (I357357,I357408);
not I_20865 (I357430,I357391);
nand I_20866 (I357447,I838615,I838603);
and I_20867 (I357464,I357447,I838606);
DFFARX1 I_20868 (I357464,I2683,I357365,I357490,);
not I_20869 (I357498,I357490);
DFFARX1 I_20870 (I838624,I2683,I357365,I357524,);
and I_20871 (I357532,I357524,I838600);
nand I_20872 (I357549,I357524,I838600);
nand I_20873 (I357336,I357498,I357549);
DFFARX1 I_20874 (I838618,I2683,I357365,I357589,);
nor I_20875 (I357597,I357589,I357532);
DFFARX1 I_20876 (I357597,I2683,I357365,I357330,);
nor I_20877 (I357345,I357589,I357490);
nand I_20878 (I357642,I838612,I838609);
and I_20879 (I357659,I357642,I838621);
DFFARX1 I_20880 (I357659,I2683,I357365,I357685,);
nor I_20881 (I357333,I357685,I357589);
not I_20882 (I357707,I357685);
nor I_20883 (I357724,I357707,I357498);
nor I_20884 (I357741,I357430,I357724);
DFFARX1 I_20885 (I357741,I2683,I357365,I357348,);
nor I_20886 (I357772,I357707,I357589);
nor I_20887 (I357789,I838600,I838609);
nor I_20888 (I357339,I357789,I357772);
not I_20889 (I357820,I357789);
nand I_20890 (I357342,I357549,I357820);
DFFARX1 I_20891 (I357789,I2683,I357365,I357354,);
DFFARX1 I_20892 (I357789,I2683,I357365,I357351,);
not I_20893 (I357909,I2690);
DFFARX1 I_20894 (I301251,I2683,I357909,I357935,);
DFFARX1 I_20895 (I357935,I2683,I357909,I357952,);
not I_20896 (I357901,I357952);
not I_20897 (I357974,I357935);
nand I_20898 (I357991,I301230,I301254);
and I_20899 (I358008,I357991,I301257);
DFFARX1 I_20900 (I358008,I2683,I357909,I358034,);
not I_20901 (I358042,I358034);
DFFARX1 I_20902 (I301239,I2683,I357909,I358068,);
and I_20903 (I358076,I358068,I301245);
nand I_20904 (I358093,I358068,I301245);
nand I_20905 (I357880,I358042,I358093);
DFFARX1 I_20906 (I301233,I2683,I357909,I358133,);
nor I_20907 (I358141,I358133,I358076);
DFFARX1 I_20908 (I358141,I2683,I357909,I357874,);
nor I_20909 (I357889,I358133,I358034);
nand I_20910 (I358186,I301242,I301230);
and I_20911 (I358203,I358186,I301236);
DFFARX1 I_20912 (I358203,I2683,I357909,I358229,);
nor I_20913 (I357877,I358229,I358133);
not I_20914 (I358251,I358229);
nor I_20915 (I358268,I358251,I358042);
nor I_20916 (I358285,I357974,I358268);
DFFARX1 I_20917 (I358285,I2683,I357909,I357892,);
nor I_20918 (I358316,I358251,I358133);
nor I_20919 (I358333,I301248,I301230);
nor I_20920 (I357883,I358333,I358316);
not I_20921 (I358364,I358333);
nand I_20922 (I357886,I358093,I358364);
DFFARX1 I_20923 (I358333,I2683,I357909,I357898,);
DFFARX1 I_20924 (I358333,I2683,I357909,I357895,);
not I_20925 (I358453,I2690);
DFFARX1 I_20926 (I154529,I2683,I358453,I358479,);
DFFARX1 I_20927 (I358479,I2683,I358453,I358496,);
not I_20928 (I358445,I358496);
not I_20929 (I358518,I358479);
nand I_20930 (I358535,I154541,I154520);
and I_20931 (I358552,I358535,I154523);
DFFARX1 I_20932 (I358552,I2683,I358453,I358578,);
not I_20933 (I358586,I358578);
DFFARX1 I_20934 (I154532,I2683,I358453,I358612,);
and I_20935 (I358620,I358612,I154544);
nand I_20936 (I358637,I358612,I154544);
nand I_20937 (I358424,I358586,I358637);
DFFARX1 I_20938 (I154538,I2683,I358453,I358677,);
nor I_20939 (I358685,I358677,I358620);
DFFARX1 I_20940 (I358685,I2683,I358453,I358418,);
nor I_20941 (I358433,I358677,I358578);
nand I_20942 (I358730,I154526,I154523);
and I_20943 (I358747,I358730,I154535);
DFFARX1 I_20944 (I358747,I2683,I358453,I358773,);
nor I_20945 (I358421,I358773,I358677);
not I_20946 (I358795,I358773);
nor I_20947 (I358812,I358795,I358586);
nor I_20948 (I358829,I358518,I358812);
DFFARX1 I_20949 (I358829,I2683,I358453,I358436,);
nor I_20950 (I358860,I358795,I358677);
nor I_20951 (I358877,I154520,I154523);
nor I_20952 (I358427,I358877,I358860);
not I_20953 (I358908,I358877);
nand I_20954 (I358430,I358637,I358908);
DFFARX1 I_20955 (I358877,I2683,I358453,I358442,);
DFFARX1 I_20956 (I358877,I2683,I358453,I358439,);
not I_20957 (I358997,I2690);
DFFARX1 I_20958 (I754235,I2683,I358997,I359023,);
DFFARX1 I_20959 (I359023,I2683,I358997,I359040,);
not I_20960 (I358989,I359040);
not I_20961 (I359062,I359023);
nand I_20962 (I359079,I754250,I754238);
and I_20963 (I359096,I359079,I754229);
DFFARX1 I_20964 (I359096,I2683,I358997,I359122,);
not I_20965 (I359130,I359122);
DFFARX1 I_20966 (I754241,I2683,I358997,I359156,);
and I_20967 (I359164,I359156,I754232);
nand I_20968 (I359181,I359156,I754232);
nand I_20969 (I358968,I359130,I359181);
DFFARX1 I_20970 (I754247,I2683,I358997,I359221,);
nor I_20971 (I359229,I359221,I359164);
DFFARX1 I_20972 (I359229,I2683,I358997,I358962,);
nor I_20973 (I358977,I359221,I359122);
nand I_20974 (I359274,I754256,I754244);
and I_20975 (I359291,I359274,I754253);
DFFARX1 I_20976 (I359291,I2683,I358997,I359317,);
nor I_20977 (I358965,I359317,I359221);
not I_20978 (I359339,I359317);
nor I_20979 (I359356,I359339,I359130);
nor I_20980 (I359373,I359062,I359356);
DFFARX1 I_20981 (I359373,I2683,I358997,I358980,);
nor I_20982 (I359404,I359339,I359221);
nor I_20983 (I359421,I754229,I754244);
nor I_20984 (I358971,I359421,I359404);
not I_20985 (I359452,I359421);
nand I_20986 (I358974,I359181,I359452);
DFFARX1 I_20987 (I359421,I2683,I358997,I358986,);
DFFARX1 I_20988 (I359421,I2683,I358997,I358983,);
not I_20989 (I359541,I2690);
DFFARX1 I_20990 (I305994,I2683,I359541,I359567,);
DFFARX1 I_20991 (I359567,I2683,I359541,I359584,);
not I_20992 (I359533,I359584);
not I_20993 (I359606,I359567);
nand I_20994 (I359623,I305973,I305997);
and I_20995 (I359640,I359623,I306000);
DFFARX1 I_20996 (I359640,I2683,I359541,I359666,);
not I_20997 (I359674,I359666);
DFFARX1 I_20998 (I305982,I2683,I359541,I359700,);
and I_20999 (I359708,I359700,I305988);
nand I_21000 (I359725,I359700,I305988);
nand I_21001 (I359512,I359674,I359725);
DFFARX1 I_21002 (I305976,I2683,I359541,I359765,);
nor I_21003 (I359773,I359765,I359708);
DFFARX1 I_21004 (I359773,I2683,I359541,I359506,);
nor I_21005 (I359521,I359765,I359666);
nand I_21006 (I359818,I305985,I305973);
and I_21007 (I359835,I359818,I305979);
DFFARX1 I_21008 (I359835,I2683,I359541,I359861,);
nor I_21009 (I359509,I359861,I359765);
not I_21010 (I359883,I359861);
nor I_21011 (I359900,I359883,I359674);
nor I_21012 (I359917,I359606,I359900);
DFFARX1 I_21013 (I359917,I2683,I359541,I359524,);
nor I_21014 (I359948,I359883,I359765);
nor I_21015 (I359965,I305991,I305973);
nor I_21016 (I359515,I359965,I359948);
not I_21017 (I359996,I359965);
nand I_21018 (I359518,I359725,I359996);
DFFARX1 I_21019 (I359965,I2683,I359541,I359530,);
DFFARX1 I_21020 (I359965,I2683,I359541,I359527,);
not I_21021 (I360085,I2690);
DFFARX1 I_21022 (I971169,I2683,I360085,I360111,);
DFFARX1 I_21023 (I360111,I2683,I360085,I360128,);
not I_21024 (I360077,I360128);
not I_21025 (I360150,I360111);
nand I_21026 (I360167,I971181,I971184);
and I_21027 (I360184,I360167,I971187);
DFFARX1 I_21028 (I360184,I2683,I360085,I360210,);
not I_21029 (I360218,I360210);
DFFARX1 I_21030 (I971172,I2683,I360085,I360244,);
and I_21031 (I360252,I360244,I971178);
nand I_21032 (I360269,I360244,I971178);
nand I_21033 (I360056,I360218,I360269);
DFFARX1 I_21034 (I971166,I2683,I360085,I360309,);
nor I_21035 (I360317,I360309,I360252);
DFFARX1 I_21036 (I360317,I2683,I360085,I360050,);
nor I_21037 (I360065,I360309,I360210);
nand I_21038 (I360362,I971169,I971190);
and I_21039 (I360379,I360362,I971175);
DFFARX1 I_21040 (I360379,I2683,I360085,I360405,);
nor I_21041 (I360053,I360405,I360309);
not I_21042 (I360427,I360405);
nor I_21043 (I360444,I360427,I360218);
nor I_21044 (I360461,I360150,I360444);
DFFARX1 I_21045 (I360461,I2683,I360085,I360068,);
nor I_21046 (I360492,I360427,I360309);
nor I_21047 (I360509,I971166,I971190);
nor I_21048 (I360059,I360509,I360492);
not I_21049 (I360540,I360509);
nand I_21050 (I360062,I360269,I360540);
DFFARX1 I_21051 (I360509,I2683,I360085,I360074,);
DFFARX1 I_21052 (I360509,I2683,I360085,I360071,);
not I_21053 (I360629,I2690);
DFFARX1 I_21054 (I31656,I2683,I360629,I360655,);
DFFARX1 I_21055 (I360655,I2683,I360629,I360672,);
not I_21056 (I360621,I360672);
not I_21057 (I360694,I360655);
nand I_21058 (I360711,I31644,I31659);
and I_21059 (I360728,I360711,I31647);
DFFARX1 I_21060 (I360728,I2683,I360629,I360754,);
not I_21061 (I360762,I360754);
DFFARX1 I_21062 (I31668,I2683,I360629,I360788,);
and I_21063 (I360796,I360788,I31662);
nand I_21064 (I360813,I360788,I31662);
nand I_21065 (I360600,I360762,I360813);
DFFARX1 I_21066 (I31665,I2683,I360629,I360853,);
nor I_21067 (I360861,I360853,I360796);
DFFARX1 I_21068 (I360861,I2683,I360629,I360594,);
nor I_21069 (I360609,I360853,I360754);
nand I_21070 (I360906,I31644,I31647);
and I_21071 (I360923,I360906,I31650);
DFFARX1 I_21072 (I360923,I2683,I360629,I360949,);
nor I_21073 (I360597,I360949,I360853);
not I_21074 (I360971,I360949);
nor I_21075 (I360988,I360971,I360762);
nor I_21076 (I361005,I360694,I360988);
DFFARX1 I_21077 (I361005,I2683,I360629,I360612,);
nor I_21078 (I361036,I360971,I360853);
nor I_21079 (I361053,I31653,I31647);
nor I_21080 (I360603,I361053,I361036);
not I_21081 (I361084,I361053);
nand I_21082 (I360606,I360813,I361084);
DFFARX1 I_21083 (I361053,I2683,I360629,I360618,);
DFFARX1 I_21084 (I361053,I2683,I360629,I360615,);
not I_21085 (I361173,I2690);
DFFARX1 I_21086 (I936285,I2683,I361173,I361199,);
DFFARX1 I_21087 (I361199,I2683,I361173,I361216,);
not I_21088 (I361165,I361216);
not I_21089 (I361238,I361199);
nand I_21090 (I361255,I936297,I936285);
and I_21091 (I361272,I361255,I936288);
DFFARX1 I_21092 (I361272,I2683,I361173,I361298,);
not I_21093 (I361306,I361298);
DFFARX1 I_21094 (I936306,I2683,I361173,I361332,);
and I_21095 (I361340,I361332,I936282);
nand I_21096 (I361357,I361332,I936282);
nand I_21097 (I361144,I361306,I361357);
DFFARX1 I_21098 (I936300,I2683,I361173,I361397,);
nor I_21099 (I361405,I361397,I361340);
DFFARX1 I_21100 (I361405,I2683,I361173,I361138,);
nor I_21101 (I361153,I361397,I361298);
nand I_21102 (I361450,I936294,I936291);
and I_21103 (I361467,I361450,I936303);
DFFARX1 I_21104 (I361467,I2683,I361173,I361493,);
nor I_21105 (I361141,I361493,I361397);
not I_21106 (I361515,I361493);
nor I_21107 (I361532,I361515,I361306);
nor I_21108 (I361549,I361238,I361532);
DFFARX1 I_21109 (I361549,I2683,I361173,I361156,);
nor I_21110 (I361580,I361515,I361397);
nor I_21111 (I361597,I936282,I936291);
nor I_21112 (I361147,I361597,I361580);
not I_21113 (I361628,I361597);
nand I_21114 (I361150,I361357,I361628);
DFFARX1 I_21115 (I361597,I2683,I361173,I361162,);
DFFARX1 I_21116 (I361597,I2683,I361173,I361159,);
not I_21117 (I361717,I2690);
DFFARX1 I_21118 (I484425,I2683,I361717,I361743,);
DFFARX1 I_21119 (I361743,I2683,I361717,I361760,);
not I_21120 (I361709,I361760);
not I_21121 (I361782,I361743);
nand I_21122 (I361799,I484422,I484443);
and I_21123 (I361816,I361799,I484446);
DFFARX1 I_21124 (I361816,I2683,I361717,I361842,);
not I_21125 (I361850,I361842);
DFFARX1 I_21126 (I484431,I2683,I361717,I361876,);
and I_21127 (I361884,I361876,I484434);
nand I_21128 (I361901,I361876,I484434);
nand I_21129 (I361688,I361850,I361901);
DFFARX1 I_21130 (I484437,I2683,I361717,I361941,);
nor I_21131 (I361949,I361941,I361884);
DFFARX1 I_21132 (I361949,I2683,I361717,I361682,);
nor I_21133 (I361697,I361941,I361842);
nand I_21134 (I361994,I484422,I484428);
and I_21135 (I362011,I361994,I484440);
DFFARX1 I_21136 (I362011,I2683,I361717,I362037,);
nor I_21137 (I361685,I362037,I361941);
not I_21138 (I362059,I362037);
nor I_21139 (I362076,I362059,I361850);
nor I_21140 (I362093,I361782,I362076);
DFFARX1 I_21141 (I362093,I2683,I361717,I361700,);
nor I_21142 (I362124,I362059,I361941);
nor I_21143 (I362141,I484425,I484428);
nor I_21144 (I361691,I362141,I362124);
not I_21145 (I362172,I362141);
nand I_21146 (I361694,I361901,I362172);
DFFARX1 I_21147 (I362141,I2683,I361717,I361706,);
DFFARX1 I_21148 (I362141,I2683,I361717,I361703,);
not I_21149 (I362261,I2690);
DFFARX1 I_21150 (I838025,I2683,I362261,I362287,);
DFFARX1 I_21151 (I362287,I2683,I362261,I362304,);
not I_21152 (I362253,I362304);
not I_21153 (I362326,I362287);
nand I_21154 (I362343,I838037,I838025);
and I_21155 (I362360,I362343,I838028);
DFFARX1 I_21156 (I362360,I2683,I362261,I362386,);
not I_21157 (I362394,I362386);
DFFARX1 I_21158 (I838046,I2683,I362261,I362420,);
and I_21159 (I362428,I362420,I838022);
nand I_21160 (I362445,I362420,I838022);
nand I_21161 (I362232,I362394,I362445);
DFFARX1 I_21162 (I838040,I2683,I362261,I362485,);
nor I_21163 (I362493,I362485,I362428);
DFFARX1 I_21164 (I362493,I2683,I362261,I362226,);
nor I_21165 (I362241,I362485,I362386);
nand I_21166 (I362538,I838034,I838031);
and I_21167 (I362555,I362538,I838043);
DFFARX1 I_21168 (I362555,I2683,I362261,I362581,);
nor I_21169 (I362229,I362581,I362485);
not I_21170 (I362603,I362581);
nor I_21171 (I362620,I362603,I362394);
nor I_21172 (I362637,I362326,I362620);
DFFARX1 I_21173 (I362637,I2683,I362261,I362244,);
nor I_21174 (I362668,I362603,I362485);
nor I_21175 (I362685,I838022,I838031);
nor I_21176 (I362235,I362685,I362668);
not I_21177 (I362716,I362685);
nand I_21178 (I362238,I362445,I362716);
DFFARX1 I_21179 (I362685,I2683,I362261,I362250,);
DFFARX1 I_21180 (I362685,I2683,I362261,I362247,);
not I_21181 (I362805,I2690);
DFFARX1 I_21182 (I672335,I2683,I362805,I362831,);
DFFARX1 I_21183 (I362831,I2683,I362805,I362848,);
not I_21184 (I362797,I362848);
not I_21185 (I362870,I362831);
nand I_21186 (I362887,I672329,I672326);
and I_21187 (I362904,I362887,I672341);
DFFARX1 I_21188 (I362904,I2683,I362805,I362930,);
not I_21189 (I362938,I362930);
DFFARX1 I_21190 (I672329,I2683,I362805,I362964,);
and I_21191 (I362972,I362964,I672323);
nand I_21192 (I362989,I362964,I672323);
nand I_21193 (I362776,I362938,I362989);
DFFARX1 I_21194 (I672323,I2683,I362805,I363029,);
nor I_21195 (I363037,I363029,I362972);
DFFARX1 I_21196 (I363037,I2683,I362805,I362770,);
nor I_21197 (I362785,I363029,I362930);
nand I_21198 (I363082,I672338,I672332);
and I_21199 (I363099,I363082,I672326);
DFFARX1 I_21200 (I363099,I2683,I362805,I363125,);
nor I_21201 (I362773,I363125,I363029);
not I_21202 (I363147,I363125);
nor I_21203 (I363164,I363147,I362938);
nor I_21204 (I363181,I362870,I363164);
DFFARX1 I_21205 (I363181,I2683,I362805,I362788,);
nor I_21206 (I363212,I363147,I363029);
nor I_21207 (I363229,I672344,I672332);
nor I_21208 (I362779,I363229,I363212);
not I_21209 (I363260,I363229);
nand I_21210 (I362782,I362989,I363260);
DFFARX1 I_21211 (I363229,I2683,I362805,I362794,);
DFFARX1 I_21212 (I363229,I2683,I362805,I362791,);
not I_21213 (I363349,I2690);
DFFARX1 I_21214 (I642296,I2683,I363349,I363375,);
DFFARX1 I_21215 (I363375,I2683,I363349,I363392,);
not I_21216 (I363341,I363392);
not I_21217 (I363414,I363375);
nand I_21218 (I363431,I642290,I642287);
and I_21219 (I363448,I363431,I642302);
DFFARX1 I_21220 (I363448,I2683,I363349,I363474,);
not I_21221 (I363482,I363474);
DFFARX1 I_21222 (I642290,I2683,I363349,I363508,);
and I_21223 (I363516,I363508,I642284);
nand I_21224 (I363533,I363508,I642284);
nand I_21225 (I363320,I363482,I363533);
DFFARX1 I_21226 (I642284,I2683,I363349,I363573,);
nor I_21227 (I363581,I363573,I363516);
DFFARX1 I_21228 (I363581,I2683,I363349,I363314,);
nor I_21229 (I363329,I363573,I363474);
nand I_21230 (I363626,I642299,I642293);
and I_21231 (I363643,I363626,I642287);
DFFARX1 I_21232 (I363643,I2683,I363349,I363669,);
nor I_21233 (I363317,I363669,I363573);
not I_21234 (I363691,I363669);
nor I_21235 (I363708,I363691,I363482);
nor I_21236 (I363725,I363414,I363708);
DFFARX1 I_21237 (I363725,I2683,I363349,I363332,);
nor I_21238 (I363756,I363691,I363573);
nor I_21239 (I363773,I642305,I642293);
nor I_21240 (I363323,I363773,I363756);
not I_21241 (I363804,I363773);
nand I_21242 (I363326,I363533,I363804);
DFFARX1 I_21243 (I363773,I2683,I363349,I363338,);
DFFARX1 I_21244 (I363773,I2683,I363349,I363335,);
not I_21245 (I363893,I2690);
DFFARX1 I_21246 (I820342,I2683,I363893,I363919,);
DFFARX1 I_21247 (I363919,I2683,I363893,I363936,);
not I_21248 (I363885,I363936);
not I_21249 (I363958,I363919);
nand I_21250 (I363975,I820342,I820360);
and I_21251 (I363992,I363975,I820354);
DFFARX1 I_21252 (I363992,I2683,I363893,I364018,);
not I_21253 (I364026,I364018);
DFFARX1 I_21254 (I820348,I2683,I363893,I364052,);
and I_21255 (I364060,I364052,I820357);
nand I_21256 (I364077,I364052,I820357);
nand I_21257 (I363864,I364026,I364077);
DFFARX1 I_21258 (I820345,I2683,I363893,I364117,);
nor I_21259 (I364125,I364117,I364060);
DFFARX1 I_21260 (I364125,I2683,I363893,I363858,);
nor I_21261 (I363873,I364117,I364018);
nand I_21262 (I364170,I820345,I820363);
and I_21263 (I364187,I364170,I820348);
DFFARX1 I_21264 (I364187,I2683,I363893,I364213,);
nor I_21265 (I363861,I364213,I364117);
not I_21266 (I364235,I364213);
nor I_21267 (I364252,I364235,I364026);
nor I_21268 (I364269,I363958,I364252);
DFFARX1 I_21269 (I364269,I2683,I363893,I363876,);
nor I_21270 (I364300,I364235,I364117);
nor I_21271 (I364317,I820351,I820363);
nor I_21272 (I363867,I364317,I364300);
not I_21273 (I364348,I364317);
nand I_21274 (I363870,I364077,I364348);
DFFARX1 I_21275 (I364317,I2683,I363893,I363882,);
DFFARX1 I_21276 (I364317,I2683,I363893,I363879,);
not I_21277 (I364437,I2690);
DFFARX1 I_21278 (I719997,I2683,I364437,I364463,);
DFFARX1 I_21279 (I364463,I2683,I364437,I364480,);
not I_21280 (I364429,I364480);
not I_21281 (I364502,I364463);
nand I_21282 (I364519,I720012,I720000);
and I_21283 (I364536,I364519,I719991);
DFFARX1 I_21284 (I364536,I2683,I364437,I364562,);
not I_21285 (I364570,I364562);
DFFARX1 I_21286 (I720003,I2683,I364437,I364596,);
and I_21287 (I364604,I364596,I719994);
nand I_21288 (I364621,I364596,I719994);
nand I_21289 (I364408,I364570,I364621);
DFFARX1 I_21290 (I720009,I2683,I364437,I364661,);
nor I_21291 (I364669,I364661,I364604);
DFFARX1 I_21292 (I364669,I2683,I364437,I364402,);
nor I_21293 (I364417,I364661,I364562);
nand I_21294 (I364714,I720018,I720006);
and I_21295 (I364731,I364714,I720015);
DFFARX1 I_21296 (I364731,I2683,I364437,I364757,);
nor I_21297 (I364405,I364757,I364661);
not I_21298 (I364779,I364757);
nor I_21299 (I364796,I364779,I364570);
nor I_21300 (I364813,I364502,I364796);
DFFARX1 I_21301 (I364813,I2683,I364437,I364420,);
nor I_21302 (I364844,I364779,I364661);
nor I_21303 (I364861,I719991,I720006);
nor I_21304 (I364411,I364861,I364844);
not I_21305 (I364892,I364861);
nand I_21306 (I364414,I364621,I364892);
DFFARX1 I_21307 (I364861,I2683,I364437,I364426,);
DFFARX1 I_21308 (I364861,I2683,I364437,I364423,);
not I_21309 (I364981,I2690);
DFFARX1 I_21310 (I760695,I2683,I364981,I365007,);
DFFARX1 I_21311 (I365007,I2683,I364981,I365024,);
not I_21312 (I364973,I365024);
not I_21313 (I365046,I365007);
nand I_21314 (I365063,I760710,I760698);
and I_21315 (I365080,I365063,I760689);
DFFARX1 I_21316 (I365080,I2683,I364981,I365106,);
not I_21317 (I365114,I365106);
DFFARX1 I_21318 (I760701,I2683,I364981,I365140,);
and I_21319 (I365148,I365140,I760692);
nand I_21320 (I365165,I365140,I760692);
nand I_21321 (I364952,I365114,I365165);
DFFARX1 I_21322 (I760707,I2683,I364981,I365205,);
nor I_21323 (I365213,I365205,I365148);
DFFARX1 I_21324 (I365213,I2683,I364981,I364946,);
nor I_21325 (I364961,I365205,I365106);
nand I_21326 (I365258,I760716,I760704);
and I_21327 (I365275,I365258,I760713);
DFFARX1 I_21328 (I365275,I2683,I364981,I365301,);
nor I_21329 (I364949,I365301,I365205);
not I_21330 (I365323,I365301);
nor I_21331 (I365340,I365323,I365114);
nor I_21332 (I365357,I365046,I365340);
DFFARX1 I_21333 (I365357,I2683,I364981,I364964,);
nor I_21334 (I365388,I365323,I365205);
nor I_21335 (I365405,I760689,I760704);
nor I_21336 (I364955,I365405,I365388);
not I_21337 (I365436,I365405);
nand I_21338 (I364958,I365165,I365436);
DFFARX1 I_21339 (I365405,I2683,I364981,I364970,);
DFFARX1 I_21340 (I365405,I2683,I364981,I364967,);
not I_21341 (I365525,I2690);
DFFARX1 I_21342 (I607539,I2683,I365525,I365551,);
DFFARX1 I_21343 (I365551,I2683,I365525,I365568,);
not I_21344 (I365517,I365568);
not I_21345 (I365590,I365551);
nand I_21346 (I365607,I607560,I607551);
and I_21347 (I365624,I365607,I607539);
DFFARX1 I_21348 (I365624,I2683,I365525,I365650,);
not I_21349 (I365658,I365650);
DFFARX1 I_21350 (I607545,I2683,I365525,I365684,);
and I_21351 (I365692,I365684,I607542);
nand I_21352 (I365709,I365684,I607542);
nand I_21353 (I365496,I365658,I365709);
DFFARX1 I_21354 (I607536,I2683,I365525,I365749,);
nor I_21355 (I365757,I365749,I365692);
DFFARX1 I_21356 (I365757,I2683,I365525,I365490,);
nor I_21357 (I365505,I365749,I365650);
nand I_21358 (I365802,I607536,I607548);
and I_21359 (I365819,I365802,I607557);
DFFARX1 I_21360 (I365819,I2683,I365525,I365845,);
nor I_21361 (I365493,I365845,I365749);
not I_21362 (I365867,I365845);
nor I_21363 (I365884,I365867,I365658);
nor I_21364 (I365901,I365590,I365884);
DFFARX1 I_21365 (I365901,I2683,I365525,I365508,);
nor I_21366 (I365932,I365867,I365749);
nor I_21367 (I365949,I607554,I607548);
nor I_21368 (I365499,I365949,I365932);
not I_21369 (I365980,I365949);
nand I_21370 (I365502,I365709,I365980);
DFFARX1 I_21371 (I365949,I2683,I365525,I365514,);
DFFARX1 I_21372 (I365949,I2683,I365525,I365511,);
not I_21373 (I366069,I2690);
DFFARX1 I_21374 (I577483,I2683,I366069,I366095,);
DFFARX1 I_21375 (I366095,I2683,I366069,I366112,);
not I_21376 (I366061,I366112);
not I_21377 (I366134,I366095);
nand I_21378 (I366151,I577504,I577495);
and I_21379 (I366168,I366151,I577483);
DFFARX1 I_21380 (I366168,I2683,I366069,I366194,);
not I_21381 (I366202,I366194);
DFFARX1 I_21382 (I577489,I2683,I366069,I366228,);
and I_21383 (I366236,I366228,I577486);
nand I_21384 (I366253,I366228,I577486);
nand I_21385 (I366040,I366202,I366253);
DFFARX1 I_21386 (I577480,I2683,I366069,I366293,);
nor I_21387 (I366301,I366293,I366236);
DFFARX1 I_21388 (I366301,I2683,I366069,I366034,);
nor I_21389 (I366049,I366293,I366194);
nand I_21390 (I366346,I577480,I577492);
and I_21391 (I366363,I366346,I577501);
DFFARX1 I_21392 (I366363,I2683,I366069,I366389,);
nor I_21393 (I366037,I366389,I366293);
not I_21394 (I366411,I366389);
nor I_21395 (I366428,I366411,I366202);
nor I_21396 (I366445,I366134,I366428);
DFFARX1 I_21397 (I366445,I2683,I366069,I366052,);
nor I_21398 (I366476,I366411,I366293);
nor I_21399 (I366493,I577498,I577492);
nor I_21400 (I366043,I366493,I366476);
not I_21401 (I366524,I366493);
nand I_21402 (I366046,I366253,I366524);
DFFARX1 I_21403 (I366493,I2683,I366069,I366058,);
DFFARX1 I_21404 (I366493,I2683,I366069,I366055,);
not I_21405 (I366613,I2690);
DFFARX1 I_21406 (I841493,I2683,I366613,I366639,);
DFFARX1 I_21407 (I366639,I2683,I366613,I366656,);
not I_21408 (I366605,I366656);
not I_21409 (I366678,I366639);
nand I_21410 (I366695,I841505,I841493);
and I_21411 (I366712,I366695,I841496);
DFFARX1 I_21412 (I366712,I2683,I366613,I366738,);
not I_21413 (I366746,I366738);
DFFARX1 I_21414 (I841514,I2683,I366613,I366772,);
and I_21415 (I366780,I366772,I841490);
nand I_21416 (I366797,I366772,I841490);
nand I_21417 (I366584,I366746,I366797);
DFFARX1 I_21418 (I841508,I2683,I366613,I366837,);
nor I_21419 (I366845,I366837,I366780);
DFFARX1 I_21420 (I366845,I2683,I366613,I366578,);
nor I_21421 (I366593,I366837,I366738);
nand I_21422 (I366890,I841502,I841499);
and I_21423 (I366907,I366890,I841511);
DFFARX1 I_21424 (I366907,I2683,I366613,I366933,);
nor I_21425 (I366581,I366933,I366837);
not I_21426 (I366955,I366933);
nor I_21427 (I366972,I366955,I366746);
nor I_21428 (I366989,I366678,I366972);
DFFARX1 I_21429 (I366989,I2683,I366613,I366596,);
nor I_21430 (I367020,I366955,I366837);
nor I_21431 (I367037,I841490,I841499);
nor I_21432 (I366587,I367037,I367020);
not I_21433 (I367068,I367037);
nand I_21434 (I366590,I366797,I367068);
DFFARX1 I_21435 (I367037,I2683,I366613,I366602,);
DFFARX1 I_21436 (I367037,I2683,I366613,I366599,);
not I_21437 (I367157,I2690);
DFFARX1 I_21438 (I89620,I2683,I367157,I367183,);
DFFARX1 I_21439 (I367183,I2683,I367157,I367200,);
not I_21440 (I367149,I367200);
not I_21441 (I367222,I367183);
nand I_21442 (I367239,I89635,I89614);
and I_21443 (I367256,I367239,I89617);
DFFARX1 I_21444 (I367256,I2683,I367157,I367282,);
not I_21445 (I367290,I367282);
DFFARX1 I_21446 (I89623,I2683,I367157,I367316,);
and I_21447 (I367324,I367316,I89617);
nand I_21448 (I367341,I367316,I89617);
nand I_21449 (I367128,I367290,I367341);
DFFARX1 I_21450 (I89632,I2683,I367157,I367381,);
nor I_21451 (I367389,I367381,I367324);
DFFARX1 I_21452 (I367389,I2683,I367157,I367122,);
nor I_21453 (I367137,I367381,I367282);
nand I_21454 (I367434,I89614,I89629);
and I_21455 (I367451,I367434,I89626);
DFFARX1 I_21456 (I367451,I2683,I367157,I367477,);
nor I_21457 (I367125,I367477,I367381);
not I_21458 (I367499,I367477);
nor I_21459 (I367516,I367499,I367290);
nor I_21460 (I367533,I367222,I367516);
DFFARX1 I_21461 (I367533,I2683,I367157,I367140,);
nor I_21462 (I367564,I367499,I367381);
nor I_21463 (I367581,I89638,I89629);
nor I_21464 (I367131,I367581,I367564);
not I_21465 (I367612,I367581);
nand I_21466 (I367134,I367341,I367612);
DFFARX1 I_21467 (I367581,I2683,I367157,I367146,);
DFFARX1 I_21468 (I367581,I2683,I367157,I367143,);
not I_21469 (I367701,I2690);
DFFARX1 I_21470 (I749713,I2683,I367701,I367727,);
DFFARX1 I_21471 (I367727,I2683,I367701,I367744,);
not I_21472 (I367693,I367744);
not I_21473 (I367766,I367727);
nand I_21474 (I367783,I749728,I749716);
and I_21475 (I367800,I367783,I749707);
DFFARX1 I_21476 (I367800,I2683,I367701,I367826,);
not I_21477 (I367834,I367826);
DFFARX1 I_21478 (I749719,I2683,I367701,I367860,);
and I_21479 (I367868,I367860,I749710);
nand I_21480 (I367885,I367860,I749710);
nand I_21481 (I367672,I367834,I367885);
DFFARX1 I_21482 (I749725,I2683,I367701,I367925,);
nor I_21483 (I367933,I367925,I367868);
DFFARX1 I_21484 (I367933,I2683,I367701,I367666,);
nor I_21485 (I367681,I367925,I367826);
nand I_21486 (I367978,I749734,I749722);
and I_21487 (I367995,I367978,I749731);
DFFARX1 I_21488 (I367995,I2683,I367701,I368021,);
nor I_21489 (I367669,I368021,I367925);
not I_21490 (I368043,I368021);
nor I_21491 (I368060,I368043,I367834);
nor I_21492 (I368077,I367766,I368060);
DFFARX1 I_21493 (I368077,I2683,I367701,I367684,);
nor I_21494 (I368108,I368043,I367925);
nor I_21495 (I368125,I749707,I749722);
nor I_21496 (I367675,I368125,I368108);
not I_21497 (I368156,I368125);
nand I_21498 (I367678,I367885,I368156);
DFFARX1 I_21499 (I368125,I2683,I367701,I367690,);
DFFARX1 I_21500 (I368125,I2683,I367701,I367687,);
not I_21501 (I368245,I2690);
DFFARX1 I_21502 (I163454,I2683,I368245,I368271,);
DFFARX1 I_21503 (I368271,I2683,I368245,I368288,);
not I_21504 (I368237,I368288);
not I_21505 (I368310,I368271);
nand I_21506 (I368327,I163466,I163445);
and I_21507 (I368344,I368327,I163448);
DFFARX1 I_21508 (I368344,I2683,I368245,I368370,);
not I_21509 (I368378,I368370);
DFFARX1 I_21510 (I163457,I2683,I368245,I368404,);
and I_21511 (I368412,I368404,I163469);
nand I_21512 (I368429,I368404,I163469);
nand I_21513 (I368216,I368378,I368429);
DFFARX1 I_21514 (I163463,I2683,I368245,I368469,);
nor I_21515 (I368477,I368469,I368412);
DFFARX1 I_21516 (I368477,I2683,I368245,I368210,);
nor I_21517 (I368225,I368469,I368370);
nand I_21518 (I368522,I163451,I163448);
and I_21519 (I368539,I368522,I163460);
DFFARX1 I_21520 (I368539,I2683,I368245,I368565,);
nor I_21521 (I368213,I368565,I368469);
not I_21522 (I368587,I368565);
nor I_21523 (I368604,I368587,I368378);
nor I_21524 (I368621,I368310,I368604);
DFFARX1 I_21525 (I368621,I2683,I368245,I368228,);
nor I_21526 (I368652,I368587,I368469);
nor I_21527 (I368669,I163445,I163448);
nor I_21528 (I368219,I368669,I368652);
not I_21529 (I368700,I368669);
nand I_21530 (I368222,I368429,I368700);
DFFARX1 I_21531 (I368669,I2683,I368245,I368234,);
DFFARX1 I_21532 (I368669,I2683,I368245,I368231,);
not I_21533 (I368789,I2690);
DFFARX1 I_21534 (I49041,I2683,I368789,I368815,);
DFFARX1 I_21535 (I368815,I2683,I368789,I368832,);
not I_21536 (I368781,I368832);
not I_21537 (I368854,I368815);
nand I_21538 (I368871,I49056,I49035);
and I_21539 (I368888,I368871,I49038);
DFFARX1 I_21540 (I368888,I2683,I368789,I368914,);
not I_21541 (I368922,I368914);
DFFARX1 I_21542 (I49044,I2683,I368789,I368948,);
and I_21543 (I368956,I368948,I49038);
nand I_21544 (I368973,I368948,I49038);
nand I_21545 (I368760,I368922,I368973);
DFFARX1 I_21546 (I49053,I2683,I368789,I369013,);
nor I_21547 (I369021,I369013,I368956);
DFFARX1 I_21548 (I369021,I2683,I368789,I368754,);
nor I_21549 (I368769,I369013,I368914);
nand I_21550 (I369066,I49035,I49050);
and I_21551 (I369083,I369066,I49047);
DFFARX1 I_21552 (I369083,I2683,I368789,I369109,);
nor I_21553 (I368757,I369109,I369013);
not I_21554 (I369131,I369109);
nor I_21555 (I369148,I369131,I368922);
nor I_21556 (I369165,I368854,I369148);
DFFARX1 I_21557 (I369165,I2683,I368789,I368772,);
nor I_21558 (I369196,I369131,I369013);
nor I_21559 (I369213,I49059,I49050);
nor I_21560 (I368763,I369213,I369196);
not I_21561 (I369244,I369213);
nand I_21562 (I368766,I368973,I369244);
DFFARX1 I_21563 (I369213,I2683,I368789,I368778,);
DFFARX1 I_21564 (I369213,I2683,I368789,I368775,);
not I_21565 (I369333,I2690);
DFFARX1 I_21566 (I984769,I2683,I369333,I369359,);
DFFARX1 I_21567 (I369359,I2683,I369333,I369376,);
not I_21568 (I369325,I369376);
not I_21569 (I369398,I369359);
nand I_21570 (I369415,I984781,I984784);
and I_21571 (I369432,I369415,I984787);
DFFARX1 I_21572 (I369432,I2683,I369333,I369458,);
not I_21573 (I369466,I369458);
DFFARX1 I_21574 (I984772,I2683,I369333,I369492,);
and I_21575 (I369500,I369492,I984778);
nand I_21576 (I369517,I369492,I984778);
nand I_21577 (I369304,I369466,I369517);
DFFARX1 I_21578 (I984766,I2683,I369333,I369557,);
nor I_21579 (I369565,I369557,I369500);
DFFARX1 I_21580 (I369565,I2683,I369333,I369298,);
nor I_21581 (I369313,I369557,I369458);
nand I_21582 (I369610,I984769,I984790);
and I_21583 (I369627,I369610,I984775);
DFFARX1 I_21584 (I369627,I2683,I369333,I369653,);
nor I_21585 (I369301,I369653,I369557);
not I_21586 (I369675,I369653);
nor I_21587 (I369692,I369675,I369466);
nor I_21588 (I369709,I369398,I369692);
DFFARX1 I_21589 (I369709,I2683,I369333,I369316,);
nor I_21590 (I369740,I369675,I369557);
nor I_21591 (I369757,I984766,I984790);
nor I_21592 (I369307,I369757,I369740);
not I_21593 (I369788,I369757);
nand I_21594 (I369310,I369517,I369788);
DFFARX1 I_21595 (I369757,I2683,I369333,I369322,);
DFFARX1 I_21596 (I369757,I2683,I369333,I369319,);
not I_21597 (I369877,I2690);
DFFARX1 I_21598 (I620689,I2683,I369877,I369903,);
DFFARX1 I_21599 (I369903,I2683,I369877,I369920,);
not I_21600 (I369869,I369920);
not I_21601 (I369942,I369903);
nand I_21602 (I369959,I620683,I620680);
and I_21603 (I369976,I369959,I620695);
DFFARX1 I_21604 (I369976,I2683,I369877,I370002,);
not I_21605 (I370010,I370002);
DFFARX1 I_21606 (I620683,I2683,I369877,I370036,);
and I_21607 (I370044,I370036,I620677);
nand I_21608 (I370061,I370036,I620677);
nand I_21609 (I369848,I370010,I370061);
DFFARX1 I_21610 (I620677,I2683,I369877,I370101,);
nor I_21611 (I370109,I370101,I370044);
DFFARX1 I_21612 (I370109,I2683,I369877,I369842,);
nor I_21613 (I369857,I370101,I370002);
nand I_21614 (I370154,I620692,I620686);
and I_21615 (I370171,I370154,I620680);
DFFARX1 I_21616 (I370171,I2683,I369877,I370197,);
nor I_21617 (I369845,I370197,I370101);
not I_21618 (I370219,I370197);
nor I_21619 (I370236,I370219,I370010);
nor I_21620 (I370253,I369942,I370236);
DFFARX1 I_21621 (I370253,I2683,I369877,I369860,);
nor I_21622 (I370284,I370219,I370101);
nor I_21623 (I370301,I620698,I620686);
nor I_21624 (I369851,I370301,I370284);
not I_21625 (I370332,I370301);
nand I_21626 (I369854,I370061,I370332);
DFFARX1 I_21627 (I370301,I2683,I369877,I369866,);
DFFARX1 I_21628 (I370301,I2683,I369877,I369863,);
not I_21629 (I370421,I2690);
DFFARX1 I_21630 (I557253,I2683,I370421,I370447,);
DFFARX1 I_21631 (I370447,I2683,I370421,I370464,);
not I_21632 (I370413,I370464);
not I_21633 (I370486,I370447);
nand I_21634 (I370503,I557274,I557265);
and I_21635 (I370520,I370503,I557253);
DFFARX1 I_21636 (I370520,I2683,I370421,I370546,);
not I_21637 (I370554,I370546);
DFFARX1 I_21638 (I557259,I2683,I370421,I370580,);
and I_21639 (I370588,I370580,I557256);
nand I_21640 (I370605,I370580,I557256);
nand I_21641 (I370392,I370554,I370605);
DFFARX1 I_21642 (I557250,I2683,I370421,I370645,);
nor I_21643 (I370653,I370645,I370588);
DFFARX1 I_21644 (I370653,I2683,I370421,I370386,);
nor I_21645 (I370401,I370645,I370546);
nand I_21646 (I370698,I557250,I557262);
and I_21647 (I370715,I370698,I557271);
DFFARX1 I_21648 (I370715,I2683,I370421,I370741,);
nor I_21649 (I370389,I370741,I370645);
not I_21650 (I370763,I370741);
nor I_21651 (I370780,I370763,I370554);
nor I_21652 (I370797,I370486,I370780);
DFFARX1 I_21653 (I370797,I2683,I370421,I370404,);
nor I_21654 (I370828,I370763,I370645);
nor I_21655 (I370845,I557268,I557262);
nor I_21656 (I370395,I370845,I370828);
not I_21657 (I370876,I370845);
nand I_21658 (I370398,I370605,I370876);
DFFARX1 I_21659 (I370845,I2683,I370421,I370410,);
DFFARX1 I_21660 (I370845,I2683,I370421,I370407,);
not I_21661 (I370965,I2690);
DFFARX1 I_21662 (I504077,I2683,I370965,I370991,);
DFFARX1 I_21663 (I370991,I2683,I370965,I371008,);
not I_21664 (I370957,I371008);
not I_21665 (I371030,I370991);
nand I_21666 (I371047,I504098,I504089);
and I_21667 (I371064,I371047,I504077);
DFFARX1 I_21668 (I371064,I2683,I370965,I371090,);
not I_21669 (I371098,I371090);
DFFARX1 I_21670 (I504083,I2683,I370965,I371124,);
and I_21671 (I371132,I371124,I504080);
nand I_21672 (I371149,I371124,I504080);
nand I_21673 (I370936,I371098,I371149);
DFFARX1 I_21674 (I504074,I2683,I370965,I371189,);
nor I_21675 (I371197,I371189,I371132);
DFFARX1 I_21676 (I371197,I2683,I370965,I370930,);
nor I_21677 (I370945,I371189,I371090);
nand I_21678 (I371242,I504074,I504086);
and I_21679 (I371259,I371242,I504095);
DFFARX1 I_21680 (I371259,I2683,I370965,I371285,);
nor I_21681 (I370933,I371285,I371189);
not I_21682 (I371307,I371285);
nor I_21683 (I371324,I371307,I371098);
nor I_21684 (I371341,I371030,I371324);
DFFARX1 I_21685 (I371341,I2683,I370965,I370948,);
nor I_21686 (I371372,I371307,I371189);
nor I_21687 (I371389,I504092,I504086);
nor I_21688 (I370939,I371389,I371372);
not I_21689 (I371420,I371389);
nand I_21690 (I370942,I371149,I371420);
DFFARX1 I_21691 (I371389,I2683,I370965,I370954,);
DFFARX1 I_21692 (I371389,I2683,I370965,I370951,);
not I_21693 (I371509,I2690);
DFFARX1 I_21694 (I33237,I2683,I371509,I371535,);
DFFARX1 I_21695 (I371535,I2683,I371509,I371552,);
not I_21696 (I371501,I371552);
not I_21697 (I371574,I371535);
nand I_21698 (I371591,I33225,I33240);
and I_21699 (I371608,I371591,I33228);
DFFARX1 I_21700 (I371608,I2683,I371509,I371634,);
not I_21701 (I371642,I371634);
DFFARX1 I_21702 (I33249,I2683,I371509,I371668,);
and I_21703 (I371676,I371668,I33243);
nand I_21704 (I371693,I371668,I33243);
nand I_21705 (I371480,I371642,I371693);
DFFARX1 I_21706 (I33246,I2683,I371509,I371733,);
nor I_21707 (I371741,I371733,I371676);
DFFARX1 I_21708 (I371741,I2683,I371509,I371474,);
nor I_21709 (I371489,I371733,I371634);
nand I_21710 (I371786,I33225,I33228);
and I_21711 (I371803,I371786,I33231);
DFFARX1 I_21712 (I371803,I2683,I371509,I371829,);
nor I_21713 (I371477,I371829,I371733);
not I_21714 (I371851,I371829);
nor I_21715 (I371868,I371851,I371642);
nor I_21716 (I371885,I371574,I371868);
DFFARX1 I_21717 (I371885,I2683,I371509,I371492,);
nor I_21718 (I371916,I371851,I371733);
nor I_21719 (I371933,I33234,I33228);
nor I_21720 (I371483,I371933,I371916);
not I_21721 (I371964,I371933);
nand I_21722 (I371486,I371693,I371964);
DFFARX1 I_21723 (I371933,I2683,I371509,I371498,);
DFFARX1 I_21724 (I371933,I2683,I371509,I371495,);
not I_21725 (I372053,I2690);
DFFARX1 I_21726 (I1014024,I2683,I372053,I372079,);
DFFARX1 I_21727 (I372079,I2683,I372053,I372096,);
not I_21728 (I372045,I372096);
not I_21729 (I372118,I372079);
nand I_21730 (I372135,I1014021,I1014018);
and I_21731 (I372152,I372135,I1014006);
DFFARX1 I_21732 (I372152,I2683,I372053,I372178,);
not I_21733 (I372186,I372178);
DFFARX1 I_21734 (I1014030,I2683,I372053,I372212,);
and I_21735 (I372220,I372212,I1014015);
nand I_21736 (I372237,I372212,I1014015);
nand I_21737 (I372024,I372186,I372237);
DFFARX1 I_21738 (I1014009,I2683,I372053,I372277,);
nor I_21739 (I372285,I372277,I372220);
DFFARX1 I_21740 (I372285,I2683,I372053,I372018,);
nor I_21741 (I372033,I372277,I372178);
nand I_21742 (I372330,I1014006,I1014012);
and I_21743 (I372347,I372330,I1014027);
DFFARX1 I_21744 (I372347,I2683,I372053,I372373,);
nor I_21745 (I372021,I372373,I372277);
not I_21746 (I372395,I372373);
nor I_21747 (I372412,I372395,I372186);
nor I_21748 (I372429,I372118,I372412);
DFFARX1 I_21749 (I372429,I2683,I372053,I372036,);
nor I_21750 (I372460,I372395,I372277);
nor I_21751 (I372477,I1014009,I1014012);
nor I_21752 (I372027,I372477,I372460);
not I_21753 (I372508,I372477);
nand I_21754 (I372030,I372237,I372508);
DFFARX1 I_21755 (I372477,I2683,I372053,I372042,);
DFFARX1 I_21756 (I372477,I2683,I372053,I372039,);
not I_21757 (I372597,I2690);
DFFARX1 I_21758 (I1048356,I2683,I372597,I372623,);
DFFARX1 I_21759 (I372623,I2683,I372597,I372640,);
not I_21760 (I372589,I372640);
not I_21761 (I372662,I372623);
nand I_21762 (I372679,I1048332,I1048353);
and I_21763 (I372696,I372679,I1048350);
DFFARX1 I_21764 (I372696,I2683,I372597,I372722,);
not I_21765 (I372730,I372722);
DFFARX1 I_21766 (I1048329,I2683,I372597,I372756,);
and I_21767 (I372764,I372756,I1048341);
nand I_21768 (I372781,I372756,I1048341);
nand I_21769 (I372568,I372730,I372781);
DFFARX1 I_21770 (I1048344,I2683,I372597,I372821,);
nor I_21771 (I372829,I372821,I372764);
DFFARX1 I_21772 (I372829,I2683,I372597,I372562,);
nor I_21773 (I372577,I372821,I372722);
nand I_21774 (I372874,I1048347,I1048335);
and I_21775 (I372891,I372874,I1048338);
DFFARX1 I_21776 (I372891,I2683,I372597,I372917,);
nor I_21777 (I372565,I372917,I372821);
not I_21778 (I372939,I372917);
nor I_21779 (I372956,I372939,I372730);
nor I_21780 (I372973,I372662,I372956);
DFFARX1 I_21781 (I372973,I2683,I372597,I372580,);
nor I_21782 (I373004,I372939,I372821);
nor I_21783 (I373021,I1048329,I1048335);
nor I_21784 (I372571,I373021,I373004);
not I_21785 (I373052,I373021);
nand I_21786 (I372574,I372781,I373052);
DFFARX1 I_21787 (I373021,I2683,I372597,I372586,);
DFFARX1 I_21788 (I373021,I2683,I372597,I372583,);
not I_21789 (I373141,I2690);
DFFARX1 I_21790 (I1040026,I2683,I373141,I373167,);
DFFARX1 I_21791 (I373167,I2683,I373141,I373184,);
not I_21792 (I373133,I373184);
not I_21793 (I373206,I373167);
nand I_21794 (I373223,I1040002,I1040023);
and I_21795 (I373240,I373223,I1040020);
DFFARX1 I_21796 (I373240,I2683,I373141,I373266,);
not I_21797 (I373274,I373266);
DFFARX1 I_21798 (I1039999,I2683,I373141,I373300,);
and I_21799 (I373308,I373300,I1040011);
nand I_21800 (I373325,I373300,I1040011);
nand I_21801 (I373112,I373274,I373325);
DFFARX1 I_21802 (I1040014,I2683,I373141,I373365,);
nor I_21803 (I373373,I373365,I373308);
DFFARX1 I_21804 (I373373,I2683,I373141,I373106,);
nor I_21805 (I373121,I373365,I373266);
nand I_21806 (I373418,I1040017,I1040005);
and I_21807 (I373435,I373418,I1040008);
DFFARX1 I_21808 (I373435,I2683,I373141,I373461,);
nor I_21809 (I373109,I373461,I373365);
not I_21810 (I373483,I373461);
nor I_21811 (I373500,I373483,I373274);
nor I_21812 (I373517,I373206,I373500);
DFFARX1 I_21813 (I373517,I2683,I373141,I373124,);
nor I_21814 (I373548,I373483,I373365);
nor I_21815 (I373565,I1039999,I1040005);
nor I_21816 (I373115,I373565,I373548);
not I_21817 (I373596,I373565);
nand I_21818 (I373118,I373325,I373596);
DFFARX1 I_21819 (I373565,I2683,I373141,I373130,);
DFFARX1 I_21820 (I373565,I2683,I373141,I373127,);
not I_21821 (I373685,I2690);
DFFARX1 I_21822 (I687618,I2683,I373685,I373711,);
DFFARX1 I_21823 (I373711,I2683,I373685,I373728,);
not I_21824 (I373677,I373728);
not I_21825 (I373750,I373711);
nand I_21826 (I373767,I687612,I687609);
and I_21827 (I373784,I373767,I687624);
DFFARX1 I_21828 (I373784,I2683,I373685,I373810,);
not I_21829 (I373818,I373810);
DFFARX1 I_21830 (I687612,I2683,I373685,I373844,);
and I_21831 (I373852,I373844,I687606);
nand I_21832 (I373869,I373844,I687606);
nand I_21833 (I373656,I373818,I373869);
DFFARX1 I_21834 (I687606,I2683,I373685,I373909,);
nor I_21835 (I373917,I373909,I373852);
DFFARX1 I_21836 (I373917,I2683,I373685,I373650,);
nor I_21837 (I373665,I373909,I373810);
nand I_21838 (I373962,I687621,I687615);
and I_21839 (I373979,I373962,I687609);
DFFARX1 I_21840 (I373979,I2683,I373685,I374005,);
nor I_21841 (I373653,I374005,I373909);
not I_21842 (I374027,I374005);
nor I_21843 (I374044,I374027,I373818);
nor I_21844 (I374061,I373750,I374044);
DFFARX1 I_21845 (I374061,I2683,I373685,I373668,);
nor I_21846 (I374092,I374027,I373909);
nor I_21847 (I374109,I687627,I687615);
nor I_21848 (I373659,I374109,I374092);
not I_21849 (I374140,I374109);
nand I_21850 (I373662,I373869,I374140);
DFFARX1 I_21851 (I374109,I2683,I373685,I373674,);
DFFARX1 I_21852 (I374109,I2683,I373685,I373671,);
not I_21853 (I374229,I2690);
DFFARX1 I_21854 (I896403,I2683,I374229,I374255,);
DFFARX1 I_21855 (I374255,I2683,I374229,I374272,);
not I_21856 (I374221,I374272);
not I_21857 (I374294,I374255);
nand I_21858 (I374311,I896415,I896403);
and I_21859 (I374328,I374311,I896406);
DFFARX1 I_21860 (I374328,I2683,I374229,I374354,);
not I_21861 (I374362,I374354);
DFFARX1 I_21862 (I896424,I2683,I374229,I374388,);
and I_21863 (I374396,I374388,I896400);
nand I_21864 (I374413,I374388,I896400);
nand I_21865 (I374200,I374362,I374413);
DFFARX1 I_21866 (I896418,I2683,I374229,I374453,);
nor I_21867 (I374461,I374453,I374396);
DFFARX1 I_21868 (I374461,I2683,I374229,I374194,);
nor I_21869 (I374209,I374453,I374354);
nand I_21870 (I374506,I896412,I896409);
and I_21871 (I374523,I374506,I896421);
DFFARX1 I_21872 (I374523,I2683,I374229,I374549,);
nor I_21873 (I374197,I374549,I374453);
not I_21874 (I374571,I374549);
nor I_21875 (I374588,I374571,I374362);
nor I_21876 (I374605,I374294,I374588);
DFFARX1 I_21877 (I374605,I2683,I374229,I374212,);
nor I_21878 (I374636,I374571,I374453);
nor I_21879 (I374653,I896400,I896409);
nor I_21880 (I374203,I374653,I374636);
not I_21881 (I374684,I374653);
nand I_21882 (I374206,I374413,I374684);
DFFARX1 I_21883 (I374653,I2683,I374229,I374218,);
DFFARX1 I_21884 (I374653,I2683,I374229,I374215,);
not I_21885 (I374773,I2690);
DFFARX1 I_21886 (I615631,I2683,I374773,I374799,);
DFFARX1 I_21887 (I374799,I2683,I374773,I374816,);
not I_21888 (I374765,I374816);
not I_21889 (I374838,I374799);
nand I_21890 (I374855,I615652,I615643);
and I_21891 (I374872,I374855,I615631);
DFFARX1 I_21892 (I374872,I2683,I374773,I374898,);
not I_21893 (I374906,I374898);
DFFARX1 I_21894 (I615637,I2683,I374773,I374932,);
and I_21895 (I374940,I374932,I615634);
nand I_21896 (I374957,I374932,I615634);
nand I_21897 (I374744,I374906,I374957);
DFFARX1 I_21898 (I615628,I2683,I374773,I374997,);
nor I_21899 (I375005,I374997,I374940);
DFFARX1 I_21900 (I375005,I2683,I374773,I374738,);
nor I_21901 (I374753,I374997,I374898);
nand I_21902 (I375050,I615628,I615640);
and I_21903 (I375067,I375050,I615649);
DFFARX1 I_21904 (I375067,I2683,I374773,I375093,);
nor I_21905 (I374741,I375093,I374997);
not I_21906 (I375115,I375093);
nor I_21907 (I375132,I375115,I374906);
nor I_21908 (I375149,I374838,I375132);
DFFARX1 I_21909 (I375149,I2683,I374773,I374756,);
nor I_21910 (I375180,I375115,I374997);
nor I_21911 (I375197,I615646,I615640);
nor I_21912 (I374747,I375197,I375180);
not I_21913 (I375228,I375197);
nand I_21914 (I374750,I374957,I375228);
DFFARX1 I_21915 (I375197,I2683,I374773,I374762,);
DFFARX1 I_21916 (I375197,I2683,I374773,I374759,);
not I_21917 (I375317,I2690);
DFFARX1 I_21918 (I209864,I2683,I375317,I375343,);
DFFARX1 I_21919 (I375343,I2683,I375317,I375360,);
not I_21920 (I375309,I375360);
not I_21921 (I375382,I375343);
nand I_21922 (I375399,I209876,I209855);
and I_21923 (I375416,I375399,I209858);
DFFARX1 I_21924 (I375416,I2683,I375317,I375442,);
not I_21925 (I375450,I375442);
DFFARX1 I_21926 (I209867,I2683,I375317,I375476,);
and I_21927 (I375484,I375476,I209879);
nand I_21928 (I375501,I375476,I209879);
nand I_21929 (I375288,I375450,I375501);
DFFARX1 I_21930 (I209873,I2683,I375317,I375541,);
nor I_21931 (I375549,I375541,I375484);
DFFARX1 I_21932 (I375549,I2683,I375317,I375282,);
nor I_21933 (I375297,I375541,I375442);
nand I_21934 (I375594,I209861,I209858);
and I_21935 (I375611,I375594,I209870);
DFFARX1 I_21936 (I375611,I2683,I375317,I375637,);
nor I_21937 (I375285,I375637,I375541);
not I_21938 (I375659,I375637);
nor I_21939 (I375676,I375659,I375450);
nor I_21940 (I375693,I375382,I375676);
DFFARX1 I_21941 (I375693,I2683,I375317,I375300,);
nor I_21942 (I375724,I375659,I375541);
nor I_21943 (I375741,I209855,I209858);
nor I_21944 (I375291,I375741,I375724);
not I_21945 (I375772,I375741);
nand I_21946 (I375294,I375501,I375772);
DFFARX1 I_21947 (I375741,I2683,I375317,I375306,);
DFFARX1 I_21948 (I375741,I2683,I375317,I375303,);
not I_21949 (I375861,I2690);
DFFARX1 I_21950 (I941487,I2683,I375861,I375887,);
DFFARX1 I_21951 (I375887,I2683,I375861,I375904,);
not I_21952 (I375853,I375904);
not I_21953 (I375926,I375887);
nand I_21954 (I375943,I941499,I941487);
and I_21955 (I375960,I375943,I941490);
DFFARX1 I_21956 (I375960,I2683,I375861,I375986,);
not I_21957 (I375994,I375986);
DFFARX1 I_21958 (I941508,I2683,I375861,I376020,);
and I_21959 (I376028,I376020,I941484);
nand I_21960 (I376045,I376020,I941484);
nand I_21961 (I375832,I375994,I376045);
DFFARX1 I_21962 (I941502,I2683,I375861,I376085,);
nor I_21963 (I376093,I376085,I376028);
DFFARX1 I_21964 (I376093,I2683,I375861,I375826,);
nor I_21965 (I375841,I376085,I375986);
nand I_21966 (I376138,I941496,I941493);
and I_21967 (I376155,I376138,I941505);
DFFARX1 I_21968 (I376155,I2683,I375861,I376181,);
nor I_21969 (I375829,I376181,I376085);
not I_21970 (I376203,I376181);
nor I_21971 (I376220,I376203,I375994);
nor I_21972 (I376237,I375926,I376220);
DFFARX1 I_21973 (I376237,I2683,I375861,I375844,);
nor I_21974 (I376268,I376203,I376085);
nor I_21975 (I376285,I941484,I941493);
nor I_21976 (I375835,I376285,I376268);
not I_21977 (I376316,I376285);
nand I_21978 (I375838,I376045,I376316);
DFFARX1 I_21979 (I376285,I2683,I375861,I375850,);
DFFARX1 I_21980 (I376285,I2683,I375861,I375847,);
not I_21981 (I376405,I2690);
DFFARX1 I_21982 (I636499,I2683,I376405,I376431,);
DFFARX1 I_21983 (I376431,I2683,I376405,I376448,);
not I_21984 (I376397,I376448);
not I_21985 (I376470,I376431);
nand I_21986 (I376487,I636493,I636490);
and I_21987 (I376504,I376487,I636505);
DFFARX1 I_21988 (I376504,I2683,I376405,I376530,);
not I_21989 (I376538,I376530);
DFFARX1 I_21990 (I636493,I2683,I376405,I376564,);
and I_21991 (I376572,I376564,I636487);
nand I_21992 (I376589,I376564,I636487);
nand I_21993 (I376376,I376538,I376589);
DFFARX1 I_21994 (I636487,I2683,I376405,I376629,);
nor I_21995 (I376637,I376629,I376572);
DFFARX1 I_21996 (I376637,I2683,I376405,I376370,);
nor I_21997 (I376385,I376629,I376530);
nand I_21998 (I376682,I636502,I636496);
and I_21999 (I376699,I376682,I636490);
DFFARX1 I_22000 (I376699,I2683,I376405,I376725,);
nor I_22001 (I376373,I376725,I376629);
not I_22002 (I376747,I376725);
nor I_22003 (I376764,I376747,I376538);
nor I_22004 (I376781,I376470,I376764);
DFFARX1 I_22005 (I376781,I2683,I376405,I376388,);
nor I_22006 (I376812,I376747,I376629);
nor I_22007 (I376829,I636508,I636496);
nor I_22008 (I376379,I376829,I376812);
not I_22009 (I376860,I376829);
nand I_22010 (I376382,I376589,I376860);
DFFARX1 I_22011 (I376829,I2683,I376405,I376394,);
DFFARX1 I_22012 (I376829,I2683,I376405,I376391,);
not I_22013 (I376949,I2690);
DFFARX1 I_22014 (I110700,I2683,I376949,I376975,);
DFFARX1 I_22015 (I376975,I2683,I376949,I376992,);
not I_22016 (I376941,I376992);
not I_22017 (I377014,I376975);
nand I_22018 (I377031,I110715,I110694);
and I_22019 (I377048,I377031,I110697);
DFFARX1 I_22020 (I377048,I2683,I376949,I377074,);
not I_22021 (I377082,I377074);
DFFARX1 I_22022 (I110703,I2683,I376949,I377108,);
and I_22023 (I377116,I377108,I110697);
nand I_22024 (I377133,I377108,I110697);
nand I_22025 (I376920,I377082,I377133);
DFFARX1 I_22026 (I110712,I2683,I376949,I377173,);
nor I_22027 (I377181,I377173,I377116);
DFFARX1 I_22028 (I377181,I2683,I376949,I376914,);
nor I_22029 (I376929,I377173,I377074);
nand I_22030 (I377226,I110694,I110709);
and I_22031 (I377243,I377226,I110706);
DFFARX1 I_22032 (I377243,I2683,I376949,I377269,);
nor I_22033 (I376917,I377269,I377173);
not I_22034 (I377291,I377269);
nor I_22035 (I377308,I377291,I377082);
nor I_22036 (I377325,I377014,I377308);
DFFARX1 I_22037 (I377325,I2683,I376949,I376932,);
nor I_22038 (I377356,I377291,I377173);
nor I_22039 (I377373,I110718,I110709);
nor I_22040 (I376923,I377373,I377356);
not I_22041 (I377404,I377373);
nand I_22042 (I376926,I377133,I377404);
DFFARX1 I_22043 (I377373,I2683,I376949,I376938,);
DFFARX1 I_22044 (I377373,I2683,I376949,I376935,);
not I_22045 (I377493,I2690);
DFFARX1 I_22046 (I718059,I2683,I377493,I377519,);
DFFARX1 I_22047 (I377519,I2683,I377493,I377536,);
not I_22048 (I377485,I377536);
not I_22049 (I377558,I377519);
nand I_22050 (I377575,I718074,I718062);
and I_22051 (I377592,I377575,I718053);
DFFARX1 I_22052 (I377592,I2683,I377493,I377618,);
not I_22053 (I377626,I377618);
DFFARX1 I_22054 (I718065,I2683,I377493,I377652,);
and I_22055 (I377660,I377652,I718056);
nand I_22056 (I377677,I377652,I718056);
nand I_22057 (I377464,I377626,I377677);
DFFARX1 I_22058 (I718071,I2683,I377493,I377717,);
nor I_22059 (I377725,I377717,I377660);
DFFARX1 I_22060 (I377725,I2683,I377493,I377458,);
nor I_22061 (I377473,I377717,I377618);
nand I_22062 (I377770,I718080,I718068);
and I_22063 (I377787,I377770,I718077);
DFFARX1 I_22064 (I377787,I2683,I377493,I377813,);
nor I_22065 (I377461,I377813,I377717);
not I_22066 (I377835,I377813);
nor I_22067 (I377852,I377835,I377626);
nor I_22068 (I377869,I377558,I377852);
DFFARX1 I_22069 (I377869,I2683,I377493,I377476,);
nor I_22070 (I377900,I377835,I377717);
nor I_22071 (I377917,I718053,I718068);
nor I_22072 (I377467,I377917,I377900);
not I_22073 (I377948,I377917);
nand I_22074 (I377470,I377677,I377948);
DFFARX1 I_22075 (I377917,I2683,I377493,I377482,);
DFFARX1 I_22076 (I377917,I2683,I377493,I377479,);
not I_22077 (I378037,I2690);
DFFARX1 I_22078 (I1015180,I2683,I378037,I378063,);
DFFARX1 I_22079 (I378063,I2683,I378037,I378080,);
not I_22080 (I378029,I378080);
not I_22081 (I378102,I378063);
nand I_22082 (I378119,I1015177,I1015174);
and I_22083 (I378136,I378119,I1015162);
DFFARX1 I_22084 (I378136,I2683,I378037,I378162,);
not I_22085 (I378170,I378162);
DFFARX1 I_22086 (I1015186,I2683,I378037,I378196,);
and I_22087 (I378204,I378196,I1015171);
nand I_22088 (I378221,I378196,I1015171);
nand I_22089 (I378008,I378170,I378221);
DFFARX1 I_22090 (I1015165,I2683,I378037,I378261,);
nor I_22091 (I378269,I378261,I378204);
DFFARX1 I_22092 (I378269,I2683,I378037,I378002,);
nor I_22093 (I378017,I378261,I378162);
nand I_22094 (I378314,I1015162,I1015168);
and I_22095 (I378331,I378314,I1015183);
DFFARX1 I_22096 (I378331,I2683,I378037,I378357,);
nor I_22097 (I378005,I378357,I378261);
not I_22098 (I378379,I378357);
nor I_22099 (I378396,I378379,I378170);
nor I_22100 (I378413,I378102,I378396);
DFFARX1 I_22101 (I378413,I2683,I378037,I378020,);
nor I_22102 (I378444,I378379,I378261);
nor I_22103 (I378461,I1015165,I1015168);
nor I_22104 (I378011,I378461,I378444);
not I_22105 (I378492,I378461);
nand I_22106 (I378014,I378221,I378492);
DFFARX1 I_22107 (I378461,I2683,I378037,I378026,);
DFFARX1 I_22108 (I378461,I2683,I378037,I378023,);
not I_22109 (I378581,I2690);
DFFARX1 I_22110 (I832823,I2683,I378581,I378607,);
DFFARX1 I_22111 (I378607,I2683,I378581,I378624,);
not I_22112 (I378573,I378624);
not I_22113 (I378646,I378607);
nand I_22114 (I378663,I832835,I832823);
and I_22115 (I378680,I378663,I832826);
DFFARX1 I_22116 (I378680,I2683,I378581,I378706,);
not I_22117 (I378714,I378706);
DFFARX1 I_22118 (I832844,I2683,I378581,I378740,);
and I_22119 (I378748,I378740,I832820);
nand I_22120 (I378765,I378740,I832820);
nand I_22121 (I378552,I378714,I378765);
DFFARX1 I_22122 (I832838,I2683,I378581,I378805,);
nor I_22123 (I378813,I378805,I378748);
DFFARX1 I_22124 (I378813,I2683,I378581,I378546,);
nor I_22125 (I378561,I378805,I378706);
nand I_22126 (I378858,I832832,I832829);
and I_22127 (I378875,I378858,I832841);
DFFARX1 I_22128 (I378875,I2683,I378581,I378901,);
nor I_22129 (I378549,I378901,I378805);
not I_22130 (I378923,I378901);
nor I_22131 (I378940,I378923,I378714);
nor I_22132 (I378957,I378646,I378940);
DFFARX1 I_22133 (I378957,I2683,I378581,I378564,);
nor I_22134 (I378988,I378923,I378805);
nor I_22135 (I379005,I832820,I832829);
nor I_22136 (I378555,I379005,I378988);
not I_22137 (I379036,I379005);
nand I_22138 (I378558,I378765,I379036);
DFFARX1 I_22139 (I379005,I2683,I378581,I378570,);
DFFARX1 I_22140 (I379005,I2683,I378581,I378567,);
not I_22141 (I379125,I2690);
DFFARX1 I_22142 (I974977,I2683,I379125,I379151,);
DFFARX1 I_22143 (I379151,I2683,I379125,I379168,);
not I_22144 (I379117,I379168);
not I_22145 (I379190,I379151);
nand I_22146 (I379207,I974989,I974992);
and I_22147 (I379224,I379207,I974995);
DFFARX1 I_22148 (I379224,I2683,I379125,I379250,);
not I_22149 (I379258,I379250);
DFFARX1 I_22150 (I974980,I2683,I379125,I379284,);
and I_22151 (I379292,I379284,I974986);
nand I_22152 (I379309,I379284,I974986);
nand I_22153 (I379096,I379258,I379309);
DFFARX1 I_22154 (I974974,I2683,I379125,I379349,);
nor I_22155 (I379357,I379349,I379292);
DFFARX1 I_22156 (I379357,I2683,I379125,I379090,);
nor I_22157 (I379105,I379349,I379250);
nand I_22158 (I379402,I974977,I974998);
and I_22159 (I379419,I379402,I974983);
DFFARX1 I_22160 (I379419,I2683,I379125,I379445,);
nor I_22161 (I379093,I379445,I379349);
not I_22162 (I379467,I379445);
nor I_22163 (I379484,I379467,I379258);
nor I_22164 (I379501,I379190,I379484);
DFFARX1 I_22165 (I379501,I2683,I379125,I379108,);
nor I_22166 (I379532,I379467,I379349);
nor I_22167 (I379549,I974974,I974998);
nor I_22168 (I379099,I379549,I379532);
not I_22169 (I379580,I379549);
nand I_22170 (I379102,I379309,I379580);
DFFARX1 I_22171 (I379549,I2683,I379125,I379114,);
DFFARX1 I_22172 (I379549,I2683,I379125,I379111,);
not I_22173 (I379669,I2690);
DFFARX1 I_22174 (I245389,I2683,I379669,I379695,);
DFFARX1 I_22175 (I379695,I2683,I379669,I379712,);
not I_22176 (I379661,I379712);
not I_22177 (I379734,I379695);
nand I_22178 (I379751,I245368,I245392);
and I_22179 (I379768,I379751,I245395);
DFFARX1 I_22180 (I379768,I2683,I379669,I379794,);
not I_22181 (I379802,I379794);
DFFARX1 I_22182 (I245377,I2683,I379669,I379828,);
and I_22183 (I379836,I379828,I245383);
nand I_22184 (I379853,I379828,I245383);
nand I_22185 (I379640,I379802,I379853);
DFFARX1 I_22186 (I245371,I2683,I379669,I379893,);
nor I_22187 (I379901,I379893,I379836);
DFFARX1 I_22188 (I379901,I2683,I379669,I379634,);
nor I_22189 (I379649,I379893,I379794);
nand I_22190 (I379946,I245380,I245368);
and I_22191 (I379963,I379946,I245374);
DFFARX1 I_22192 (I379963,I2683,I379669,I379989,);
nor I_22193 (I379637,I379989,I379893);
not I_22194 (I380011,I379989);
nor I_22195 (I380028,I380011,I379802);
nor I_22196 (I380045,I379734,I380028);
DFFARX1 I_22197 (I380045,I2683,I379669,I379652,);
nor I_22198 (I380076,I380011,I379893);
nor I_22199 (I380093,I245386,I245368);
nor I_22200 (I379643,I380093,I380076);
not I_22201 (I380124,I380093);
nand I_22202 (I379646,I379853,I380124);
DFFARX1 I_22203 (I380093,I2683,I379669,I379658,);
DFFARX1 I_22204 (I380093,I2683,I379669,I379655,);
not I_22205 (I380213,I2690);
DFFARX1 I_22206 (I1014602,I2683,I380213,I380239,);
DFFARX1 I_22207 (I380239,I2683,I380213,I380256,);
not I_22208 (I380205,I380256);
not I_22209 (I380278,I380239);
nand I_22210 (I380295,I1014599,I1014596);
and I_22211 (I380312,I380295,I1014584);
DFFARX1 I_22212 (I380312,I2683,I380213,I380338,);
not I_22213 (I380346,I380338);
DFFARX1 I_22214 (I1014608,I2683,I380213,I380372,);
and I_22215 (I380380,I380372,I1014593);
nand I_22216 (I380397,I380372,I1014593);
nand I_22217 (I380184,I380346,I380397);
DFFARX1 I_22218 (I1014587,I2683,I380213,I380437,);
nor I_22219 (I380445,I380437,I380380);
DFFARX1 I_22220 (I380445,I2683,I380213,I380178,);
nor I_22221 (I380193,I380437,I380338);
nand I_22222 (I380490,I1014584,I1014590);
and I_22223 (I380507,I380490,I1014605);
DFFARX1 I_22224 (I380507,I2683,I380213,I380533,);
nor I_22225 (I380181,I380533,I380437);
not I_22226 (I380555,I380533);
nor I_22227 (I380572,I380555,I380346);
nor I_22228 (I380589,I380278,I380572);
DFFARX1 I_22229 (I380589,I2683,I380213,I380196,);
nor I_22230 (I380620,I380555,I380437);
nor I_22231 (I380637,I1014587,I1014590);
nor I_22232 (I380187,I380637,I380620);
not I_22233 (I380668,I380637);
nand I_22234 (I380190,I380397,I380668);
DFFARX1 I_22235 (I380637,I2683,I380213,I380202,);
DFFARX1 I_22236 (I380637,I2683,I380213,I380199,);
not I_22237 (I380757,I2690);
DFFARX1 I_22238 (I263834,I2683,I380757,I380783,);
DFFARX1 I_22239 (I380783,I2683,I380757,I380800,);
not I_22240 (I380749,I380800);
not I_22241 (I380822,I380783);
nand I_22242 (I380839,I263813,I263837);
and I_22243 (I380856,I380839,I263840);
DFFARX1 I_22244 (I380856,I2683,I380757,I380882,);
not I_22245 (I380890,I380882);
DFFARX1 I_22246 (I263822,I2683,I380757,I380916,);
and I_22247 (I380924,I380916,I263828);
nand I_22248 (I380941,I380916,I263828);
nand I_22249 (I380728,I380890,I380941);
DFFARX1 I_22250 (I263816,I2683,I380757,I380981,);
nor I_22251 (I380989,I380981,I380924);
DFFARX1 I_22252 (I380989,I2683,I380757,I380722,);
nor I_22253 (I380737,I380981,I380882);
nand I_22254 (I381034,I263825,I263813);
and I_22255 (I381051,I381034,I263819);
DFFARX1 I_22256 (I381051,I2683,I380757,I381077,);
nor I_22257 (I380725,I381077,I380981);
not I_22258 (I381099,I381077);
nor I_22259 (I381116,I381099,I380890);
nor I_22260 (I381133,I380822,I381116);
DFFARX1 I_22261 (I381133,I2683,I380757,I380740,);
nor I_22262 (I381164,I381099,I380981);
nor I_22263 (I381181,I263831,I263813);
nor I_22264 (I380731,I381181,I381164);
not I_22265 (I381212,I381181);
nand I_22266 (I380734,I380941,I381212);
DFFARX1 I_22267 (I381181,I2683,I380757,I380746,);
DFFARX1 I_22268 (I381181,I2683,I380757,I380743,);
not I_22269 (I381301,I2690);
DFFARX1 I_22270 (I475755,I2683,I381301,I381327,);
DFFARX1 I_22271 (I381327,I2683,I381301,I381344,);
not I_22272 (I381293,I381344);
not I_22273 (I381366,I381327);
nand I_22274 (I381383,I475752,I475773);
and I_22275 (I381400,I381383,I475776);
DFFARX1 I_22276 (I381400,I2683,I381301,I381426,);
not I_22277 (I381434,I381426);
DFFARX1 I_22278 (I475761,I2683,I381301,I381460,);
and I_22279 (I381468,I381460,I475764);
nand I_22280 (I381485,I381460,I475764);
nand I_22281 (I381272,I381434,I381485);
DFFARX1 I_22282 (I475767,I2683,I381301,I381525,);
nor I_22283 (I381533,I381525,I381468);
DFFARX1 I_22284 (I381533,I2683,I381301,I381266,);
nor I_22285 (I381281,I381525,I381426);
nand I_22286 (I381578,I475752,I475758);
and I_22287 (I381595,I381578,I475770);
DFFARX1 I_22288 (I381595,I2683,I381301,I381621,);
nor I_22289 (I381269,I381621,I381525);
not I_22290 (I381643,I381621);
nor I_22291 (I381660,I381643,I381434);
nor I_22292 (I381677,I381366,I381660);
DFFARX1 I_22293 (I381677,I2683,I381301,I381284,);
nor I_22294 (I381708,I381643,I381525);
nor I_22295 (I381725,I475755,I475758);
nor I_22296 (I381275,I381725,I381708);
not I_22297 (I381756,I381725);
nand I_22298 (I381278,I381485,I381756);
DFFARX1 I_22299 (I381725,I2683,I381301,I381290,);
DFFARX1 I_22300 (I381725,I2683,I381301,I381287,);
not I_22301 (I381845,I2690);
DFFARX1 I_22302 (I266996,I2683,I381845,I381871,);
DFFARX1 I_22303 (I381871,I2683,I381845,I381888,);
not I_22304 (I381837,I381888);
not I_22305 (I381910,I381871);
nand I_22306 (I381927,I266975,I266999);
and I_22307 (I381944,I381927,I267002);
DFFARX1 I_22308 (I381944,I2683,I381845,I381970,);
not I_22309 (I381978,I381970);
DFFARX1 I_22310 (I266984,I2683,I381845,I382004,);
and I_22311 (I382012,I382004,I266990);
nand I_22312 (I382029,I382004,I266990);
nand I_22313 (I381816,I381978,I382029);
DFFARX1 I_22314 (I266978,I2683,I381845,I382069,);
nor I_22315 (I382077,I382069,I382012);
DFFARX1 I_22316 (I382077,I2683,I381845,I381810,);
nor I_22317 (I381825,I382069,I381970);
nand I_22318 (I382122,I266987,I266975);
and I_22319 (I382139,I382122,I266981);
DFFARX1 I_22320 (I382139,I2683,I381845,I382165,);
nor I_22321 (I381813,I382165,I382069);
not I_22322 (I382187,I382165);
nor I_22323 (I382204,I382187,I381978);
nor I_22324 (I382221,I381910,I382204);
DFFARX1 I_22325 (I382221,I2683,I381845,I381828,);
nor I_22326 (I382252,I382187,I382069);
nor I_22327 (I382269,I266993,I266975);
nor I_22328 (I381819,I382269,I382252);
not I_22329 (I382300,I382269);
nand I_22330 (I381822,I382029,I382300);
DFFARX1 I_22331 (I382269,I2683,I381845,I381834,);
DFFARX1 I_22332 (I382269,I2683,I381845,I381831,);
not I_22333 (I382389,I2690);
DFFARX1 I_22334 (I291765,I2683,I382389,I382415,);
DFFARX1 I_22335 (I382415,I2683,I382389,I382432,);
not I_22336 (I382381,I382432);
not I_22337 (I382454,I382415);
nand I_22338 (I382471,I291744,I291768);
and I_22339 (I382488,I382471,I291771);
DFFARX1 I_22340 (I382488,I2683,I382389,I382514,);
not I_22341 (I382522,I382514);
DFFARX1 I_22342 (I291753,I2683,I382389,I382548,);
and I_22343 (I382556,I382548,I291759);
nand I_22344 (I382573,I382548,I291759);
nand I_22345 (I382360,I382522,I382573);
DFFARX1 I_22346 (I291747,I2683,I382389,I382613,);
nor I_22347 (I382621,I382613,I382556);
DFFARX1 I_22348 (I382621,I2683,I382389,I382354,);
nor I_22349 (I382369,I382613,I382514);
nand I_22350 (I382666,I291756,I291744);
and I_22351 (I382683,I382666,I291750);
DFFARX1 I_22352 (I382683,I2683,I382389,I382709,);
nor I_22353 (I382357,I382709,I382613);
not I_22354 (I382731,I382709);
nor I_22355 (I382748,I382731,I382522);
nor I_22356 (I382765,I382454,I382748);
DFFARX1 I_22357 (I382765,I2683,I382389,I382372,);
nor I_22358 (I382796,I382731,I382613);
nor I_22359 (I382813,I291762,I291744);
nor I_22360 (I382363,I382813,I382796);
not I_22361 (I382844,I382813);
nand I_22362 (I382366,I382573,I382844);
DFFARX1 I_22363 (I382813,I2683,I382389,I382378,);
DFFARX1 I_22364 (I382813,I2683,I382389,I382375,);
not I_22365 (I382933,I2690);
DFFARX1 I_22366 (I307048,I2683,I382933,I382959,);
DFFARX1 I_22367 (I382959,I2683,I382933,I382976,);
not I_22368 (I382925,I382976);
not I_22369 (I382998,I382959);
nand I_22370 (I383015,I307027,I307051);
and I_22371 (I383032,I383015,I307054);
DFFARX1 I_22372 (I383032,I2683,I382933,I383058,);
not I_22373 (I383066,I383058);
DFFARX1 I_22374 (I307036,I2683,I382933,I383092,);
and I_22375 (I383100,I383092,I307042);
nand I_22376 (I383117,I383092,I307042);
nand I_22377 (I382904,I383066,I383117);
DFFARX1 I_22378 (I307030,I2683,I382933,I383157,);
nor I_22379 (I383165,I383157,I383100);
DFFARX1 I_22380 (I383165,I2683,I382933,I382898,);
nor I_22381 (I382913,I383157,I383058);
nand I_22382 (I383210,I307039,I307027);
and I_22383 (I383227,I383210,I307033);
DFFARX1 I_22384 (I383227,I2683,I382933,I383253,);
nor I_22385 (I382901,I383253,I383157);
not I_22386 (I383275,I383253);
nor I_22387 (I383292,I383275,I383066);
nor I_22388 (I383309,I382998,I383292);
DFFARX1 I_22389 (I383309,I2683,I382933,I382916,);
nor I_22390 (I383340,I383275,I383157);
nor I_22391 (I383357,I307045,I307027);
nor I_22392 (I382907,I383357,I383340);
not I_22393 (I383388,I383357);
nand I_22394 (I382910,I383117,I383388);
DFFARX1 I_22395 (I383357,I2683,I382933,I382922,);
DFFARX1 I_22396 (I383357,I2683,I382933,I382919,);
not I_22397 (I383477,I2690);
DFFARX1 I_22398 (I480957,I2683,I383477,I383503,);
DFFARX1 I_22399 (I383503,I2683,I383477,I383520,);
not I_22400 (I383469,I383520);
not I_22401 (I383542,I383503);
nand I_22402 (I383559,I480954,I480975);
and I_22403 (I383576,I383559,I480978);
DFFARX1 I_22404 (I383576,I2683,I383477,I383602,);
not I_22405 (I383610,I383602);
DFFARX1 I_22406 (I480963,I2683,I383477,I383636,);
and I_22407 (I383644,I383636,I480966);
nand I_22408 (I383661,I383636,I480966);
nand I_22409 (I383448,I383610,I383661);
DFFARX1 I_22410 (I480969,I2683,I383477,I383701,);
nor I_22411 (I383709,I383701,I383644);
DFFARX1 I_22412 (I383709,I2683,I383477,I383442,);
nor I_22413 (I383457,I383701,I383602);
nand I_22414 (I383754,I480954,I480960);
and I_22415 (I383771,I383754,I480972);
DFFARX1 I_22416 (I383771,I2683,I383477,I383797,);
nor I_22417 (I383445,I383797,I383701);
not I_22418 (I383819,I383797);
nor I_22419 (I383836,I383819,I383610);
nor I_22420 (I383853,I383542,I383836);
DFFARX1 I_22421 (I383853,I2683,I383477,I383460,);
nor I_22422 (I383884,I383819,I383701);
nor I_22423 (I383901,I480957,I480960);
nor I_22424 (I383451,I383901,I383884);
not I_22425 (I383932,I383901);
nand I_22426 (I383454,I383661,I383932);
DFFARX1 I_22427 (I383901,I2683,I383477,I383466,);
DFFARX1 I_22428 (I383901,I2683,I383477,I383463,);
not I_22429 (I384021,I2690);
DFFARX1 I_22430 (I194989,I2683,I384021,I384047,);
DFFARX1 I_22431 (I384047,I2683,I384021,I384064,);
not I_22432 (I384013,I384064);
not I_22433 (I384086,I384047);
nand I_22434 (I384103,I195001,I194980);
and I_22435 (I384120,I384103,I194983);
DFFARX1 I_22436 (I384120,I2683,I384021,I384146,);
not I_22437 (I384154,I384146);
DFFARX1 I_22438 (I194992,I2683,I384021,I384180,);
and I_22439 (I384188,I384180,I195004);
nand I_22440 (I384205,I384180,I195004);
nand I_22441 (I383992,I384154,I384205);
DFFARX1 I_22442 (I194998,I2683,I384021,I384245,);
nor I_22443 (I384253,I384245,I384188);
DFFARX1 I_22444 (I384253,I2683,I384021,I383986,);
nor I_22445 (I384001,I384245,I384146);
nand I_22446 (I384298,I194986,I194983);
and I_22447 (I384315,I384298,I194995);
DFFARX1 I_22448 (I384315,I2683,I384021,I384341,);
nor I_22449 (I383989,I384341,I384245);
not I_22450 (I384363,I384341);
nor I_22451 (I384380,I384363,I384154);
nor I_22452 (I384397,I384086,I384380);
DFFARX1 I_22453 (I384397,I2683,I384021,I384004,);
nor I_22454 (I384428,I384363,I384245);
nor I_22455 (I384445,I194980,I194983);
nor I_22456 (I383995,I384445,I384428);
not I_22457 (I384476,I384445);
nand I_22458 (I383998,I384205,I384476);
DFFARX1 I_22459 (I384445,I2683,I384021,I384010,);
DFFARX1 I_22460 (I384445,I2683,I384021,I384007,);
not I_22461 (I384565,I2690);
DFFARX1 I_22462 (I9256,I2683,I384565,I384591,);
DFFARX1 I_22463 (I384591,I2683,I384565,I384608,);
not I_22464 (I384557,I384608);
not I_22465 (I384630,I384591);
nand I_22466 (I384647,I9259,I9247);
and I_22467 (I384664,I384647,I9253);
DFFARX1 I_22468 (I384664,I2683,I384565,I384690,);
not I_22469 (I384698,I384690);
DFFARX1 I_22470 (I9241,I2683,I384565,I384724,);
and I_22471 (I384732,I384724,I9238);
nand I_22472 (I384749,I384724,I9238);
nand I_22473 (I384536,I384698,I384749);
DFFARX1 I_22474 (I9244,I2683,I384565,I384789,);
nor I_22475 (I384797,I384789,I384732);
DFFARX1 I_22476 (I384797,I2683,I384565,I384530,);
nor I_22477 (I384545,I384789,I384690);
nand I_22478 (I384842,I9244,I9241);
and I_22479 (I384859,I384842,I9238);
DFFARX1 I_22480 (I384859,I2683,I384565,I384885,);
nor I_22481 (I384533,I384885,I384789);
not I_22482 (I384907,I384885);
nor I_22483 (I384924,I384907,I384698);
nor I_22484 (I384941,I384630,I384924);
DFFARX1 I_22485 (I384941,I2683,I384565,I384548,);
nor I_22486 (I384972,I384907,I384789);
nor I_22487 (I384989,I9250,I9241);
nor I_22488 (I384539,I384989,I384972);
not I_22489 (I385020,I384989);
nand I_22490 (I384542,I384749,I385020);
DFFARX1 I_22491 (I384989,I2683,I384565,I384554,);
DFFARX1 I_22492 (I384989,I2683,I384565,I384551,);
not I_22493 (I385109,I2690);
DFFARX1 I_22494 (I638607,I2683,I385109,I385135,);
DFFARX1 I_22495 (I385135,I2683,I385109,I385152,);
not I_22496 (I385101,I385152);
not I_22497 (I385174,I385135);
nand I_22498 (I385191,I638601,I638598);
and I_22499 (I385208,I385191,I638613);
DFFARX1 I_22500 (I385208,I2683,I385109,I385234,);
not I_22501 (I385242,I385234);
DFFARX1 I_22502 (I638601,I2683,I385109,I385268,);
and I_22503 (I385276,I385268,I638595);
nand I_22504 (I385293,I385268,I638595);
nand I_22505 (I385080,I385242,I385293);
DFFARX1 I_22506 (I638595,I2683,I385109,I385333,);
nor I_22507 (I385341,I385333,I385276);
DFFARX1 I_22508 (I385341,I2683,I385109,I385074,);
nor I_22509 (I385089,I385333,I385234);
nand I_22510 (I385386,I638610,I638604);
and I_22511 (I385403,I385386,I638598);
DFFARX1 I_22512 (I385403,I2683,I385109,I385429,);
nor I_22513 (I385077,I385429,I385333);
not I_22514 (I385451,I385429);
nor I_22515 (I385468,I385451,I385242);
nor I_22516 (I385485,I385174,I385468);
DFFARX1 I_22517 (I385485,I2683,I385109,I385092,);
nor I_22518 (I385516,I385451,I385333);
nor I_22519 (I385533,I638616,I638604);
nor I_22520 (I385083,I385533,I385516);
not I_22521 (I385564,I385533);
nand I_22522 (I385086,I385293,I385564);
DFFARX1 I_22523 (I385533,I2683,I385109,I385098,);
DFFARX1 I_22524 (I385533,I2683,I385109,I385095,);
not I_22525 (I385653,I2690);
DFFARX1 I_22526 (I676551,I2683,I385653,I385679,);
DFFARX1 I_22527 (I385679,I2683,I385653,I385696,);
not I_22528 (I385645,I385696);
not I_22529 (I385718,I385679);
nand I_22530 (I385735,I676545,I676542);
and I_22531 (I385752,I385735,I676557);
DFFARX1 I_22532 (I385752,I2683,I385653,I385778,);
not I_22533 (I385786,I385778);
DFFARX1 I_22534 (I676545,I2683,I385653,I385812,);
and I_22535 (I385820,I385812,I676539);
nand I_22536 (I385837,I385812,I676539);
nand I_22537 (I385624,I385786,I385837);
DFFARX1 I_22538 (I676539,I2683,I385653,I385877,);
nor I_22539 (I385885,I385877,I385820);
DFFARX1 I_22540 (I385885,I2683,I385653,I385618,);
nor I_22541 (I385633,I385877,I385778);
nand I_22542 (I385930,I676554,I676548);
and I_22543 (I385947,I385930,I676542);
DFFARX1 I_22544 (I385947,I2683,I385653,I385973,);
nor I_22545 (I385621,I385973,I385877);
not I_22546 (I385995,I385973);
nor I_22547 (I386012,I385995,I385786);
nor I_22548 (I386029,I385718,I386012);
DFFARX1 I_22549 (I386029,I2683,I385653,I385636,);
nor I_22550 (I386060,I385995,I385877);
nor I_22551 (I386077,I676560,I676548);
nor I_22552 (I385627,I386077,I386060);
not I_22553 (I386108,I386077);
nand I_22554 (I385630,I385837,I386108);
DFFARX1 I_22555 (I386077,I2683,I385653,I385642,);
DFFARX1 I_22556 (I386077,I2683,I385653,I385639,);
not I_22557 (I386197,I2690);
DFFARX1 I_22558 (I657579,I2683,I386197,I386223,);
DFFARX1 I_22559 (I386223,I2683,I386197,I386240,);
not I_22560 (I386189,I386240);
not I_22561 (I386262,I386223);
nand I_22562 (I386279,I657573,I657570);
and I_22563 (I386296,I386279,I657585);
DFFARX1 I_22564 (I386296,I2683,I386197,I386322,);
not I_22565 (I386330,I386322);
DFFARX1 I_22566 (I657573,I2683,I386197,I386356,);
and I_22567 (I386364,I386356,I657567);
nand I_22568 (I386381,I386356,I657567);
nand I_22569 (I386168,I386330,I386381);
DFFARX1 I_22570 (I657567,I2683,I386197,I386421,);
nor I_22571 (I386429,I386421,I386364);
DFFARX1 I_22572 (I386429,I2683,I386197,I386162,);
nor I_22573 (I386177,I386421,I386322);
nand I_22574 (I386474,I657582,I657576);
and I_22575 (I386491,I386474,I657570);
DFFARX1 I_22576 (I386491,I2683,I386197,I386517,);
nor I_22577 (I386165,I386517,I386421);
not I_22578 (I386539,I386517);
nor I_22579 (I386556,I386539,I386330);
nor I_22580 (I386573,I386262,I386556);
DFFARX1 I_22581 (I386573,I2683,I386197,I386180,);
nor I_22582 (I386604,I386539,I386421);
nor I_22583 (I386621,I657588,I657576);
nor I_22584 (I386171,I386621,I386604);
not I_22585 (I386652,I386621);
nand I_22586 (I386174,I386381,I386652);
DFFARX1 I_22587 (I386621,I2683,I386197,I386186,);
DFFARX1 I_22588 (I386621,I2683,I386197,I386183,);
not I_22589 (I386741,I2690);
DFFARX1 I_22590 (I558987,I2683,I386741,I386767,);
DFFARX1 I_22591 (I386767,I2683,I386741,I386784,);
not I_22592 (I386733,I386784);
not I_22593 (I386806,I386767);
nand I_22594 (I386823,I559008,I558999);
and I_22595 (I386840,I386823,I558987);
DFFARX1 I_22596 (I386840,I2683,I386741,I386866,);
not I_22597 (I386874,I386866);
DFFARX1 I_22598 (I558993,I2683,I386741,I386900,);
and I_22599 (I386908,I386900,I558990);
nand I_22600 (I386925,I386900,I558990);
nand I_22601 (I386712,I386874,I386925);
DFFARX1 I_22602 (I558984,I2683,I386741,I386965,);
nor I_22603 (I386973,I386965,I386908);
DFFARX1 I_22604 (I386973,I2683,I386741,I386706,);
nor I_22605 (I386721,I386965,I386866);
nand I_22606 (I387018,I558984,I558996);
and I_22607 (I387035,I387018,I559005);
DFFARX1 I_22608 (I387035,I2683,I386741,I387061,);
nor I_22609 (I386709,I387061,I386965);
not I_22610 (I387083,I387061);
nor I_22611 (I387100,I387083,I386874);
nor I_22612 (I387117,I386806,I387100);
DFFARX1 I_22613 (I387117,I2683,I386741,I386724,);
nor I_22614 (I387148,I387083,I386965);
nor I_22615 (I387165,I559002,I558996);
nor I_22616 (I386715,I387165,I387148);
not I_22617 (I387196,I387165);
nand I_22618 (I386718,I386925,I387196);
DFFARX1 I_22619 (I387165,I2683,I386741,I386730,);
DFFARX1 I_22620 (I387165,I2683,I386741,I386727,);
not I_22621 (I387285,I2690);
DFFARX1 I_22622 (I102795,I2683,I387285,I387311,);
DFFARX1 I_22623 (I387311,I2683,I387285,I387328,);
not I_22624 (I387277,I387328);
not I_22625 (I387350,I387311);
nand I_22626 (I387367,I102810,I102789);
and I_22627 (I387384,I387367,I102792);
DFFARX1 I_22628 (I387384,I2683,I387285,I387410,);
not I_22629 (I387418,I387410);
DFFARX1 I_22630 (I102798,I2683,I387285,I387444,);
and I_22631 (I387452,I387444,I102792);
nand I_22632 (I387469,I387444,I102792);
nand I_22633 (I387256,I387418,I387469);
DFFARX1 I_22634 (I102807,I2683,I387285,I387509,);
nor I_22635 (I387517,I387509,I387452);
DFFARX1 I_22636 (I387517,I2683,I387285,I387250,);
nor I_22637 (I387265,I387509,I387410);
nand I_22638 (I387562,I102789,I102804);
and I_22639 (I387579,I387562,I102801);
DFFARX1 I_22640 (I387579,I2683,I387285,I387605,);
nor I_22641 (I387253,I387605,I387509);
not I_22642 (I387627,I387605);
nor I_22643 (I387644,I387627,I387418);
nor I_22644 (I387661,I387350,I387644);
DFFARX1 I_22645 (I387661,I2683,I387285,I387268,);
nor I_22646 (I387692,I387627,I387509);
nor I_22647 (I387709,I102813,I102804);
nor I_22648 (I387259,I387709,I387692);
not I_22649 (I387740,I387709);
nand I_22650 (I387262,I387469,I387740);
DFFARX1 I_22651 (I387709,I2683,I387285,I387274,);
DFFARX1 I_22652 (I387709,I2683,I387285,I387271,);
not I_22653 (I387829,I2690);
DFFARX1 I_22654 (I260145,I2683,I387829,I387855,);
DFFARX1 I_22655 (I387855,I2683,I387829,I387872,);
not I_22656 (I387821,I387872);
not I_22657 (I387894,I387855);
nand I_22658 (I387911,I260124,I260148);
and I_22659 (I387928,I387911,I260151);
DFFARX1 I_22660 (I387928,I2683,I387829,I387954,);
not I_22661 (I387962,I387954);
DFFARX1 I_22662 (I260133,I2683,I387829,I387988,);
and I_22663 (I387996,I387988,I260139);
nand I_22664 (I388013,I387988,I260139);
nand I_22665 (I387800,I387962,I388013);
DFFARX1 I_22666 (I260127,I2683,I387829,I388053,);
nor I_22667 (I388061,I388053,I387996);
DFFARX1 I_22668 (I388061,I2683,I387829,I387794,);
nor I_22669 (I387809,I388053,I387954);
nand I_22670 (I388106,I260136,I260124);
and I_22671 (I388123,I388106,I260130);
DFFARX1 I_22672 (I388123,I2683,I387829,I388149,);
nor I_22673 (I387797,I388149,I388053);
not I_22674 (I388171,I388149);
nor I_22675 (I388188,I388171,I387962);
nor I_22676 (I388205,I387894,I388188);
DFFARX1 I_22677 (I388205,I2683,I387829,I387812,);
nor I_22678 (I388236,I388171,I388053);
nor I_22679 (I388253,I260142,I260124);
nor I_22680 (I387803,I388253,I388236);
not I_22681 (I388284,I388253);
nand I_22682 (I387806,I388013,I388284);
DFFARX1 I_22683 (I388253,I2683,I387829,I387818,);
DFFARX1 I_22684 (I388253,I2683,I387829,I387815,);
not I_22685 (I388373,I2690);
DFFARX1 I_22686 (I837447,I2683,I388373,I388399,);
DFFARX1 I_22687 (I388399,I2683,I388373,I388416,);
not I_22688 (I388365,I388416);
not I_22689 (I388438,I388399);
nand I_22690 (I388455,I837459,I837447);
and I_22691 (I388472,I388455,I837450);
DFFARX1 I_22692 (I388472,I2683,I388373,I388498,);
not I_22693 (I388506,I388498);
DFFARX1 I_22694 (I837468,I2683,I388373,I388532,);
and I_22695 (I388540,I388532,I837444);
nand I_22696 (I388557,I388532,I837444);
nand I_22697 (I388344,I388506,I388557);
DFFARX1 I_22698 (I837462,I2683,I388373,I388597,);
nor I_22699 (I388605,I388597,I388540);
DFFARX1 I_22700 (I388605,I2683,I388373,I388338,);
nor I_22701 (I388353,I388597,I388498);
nand I_22702 (I388650,I837456,I837453);
and I_22703 (I388667,I388650,I837465);
DFFARX1 I_22704 (I388667,I2683,I388373,I388693,);
nor I_22705 (I388341,I388693,I388597);
not I_22706 (I388715,I388693);
nor I_22707 (I388732,I388715,I388506);
nor I_22708 (I388749,I388438,I388732);
DFFARX1 I_22709 (I388749,I2683,I388373,I388356,);
nor I_22710 (I388780,I388715,I388597);
nor I_22711 (I388797,I837444,I837453);
nor I_22712 (I388347,I388797,I388780);
not I_22713 (I388828,I388797);
nand I_22714 (I388350,I388557,I388828);
DFFARX1 I_22715 (I388797,I2683,I388373,I388362,);
DFFARX1 I_22716 (I388797,I2683,I388373,I388359,);
not I_22717 (I388917,I2690);
DFFARX1 I_22718 (I870393,I2683,I388917,I388943,);
DFFARX1 I_22719 (I388943,I2683,I388917,I388960,);
not I_22720 (I388909,I388960);
not I_22721 (I388982,I388943);
nand I_22722 (I388999,I870405,I870393);
and I_22723 (I389016,I388999,I870396);
DFFARX1 I_22724 (I389016,I2683,I388917,I389042,);
not I_22725 (I389050,I389042);
DFFARX1 I_22726 (I870414,I2683,I388917,I389076,);
and I_22727 (I389084,I389076,I870390);
nand I_22728 (I389101,I389076,I870390);
nand I_22729 (I388888,I389050,I389101);
DFFARX1 I_22730 (I870408,I2683,I388917,I389141,);
nor I_22731 (I389149,I389141,I389084);
DFFARX1 I_22732 (I389149,I2683,I388917,I388882,);
nor I_22733 (I388897,I389141,I389042);
nand I_22734 (I389194,I870402,I870399);
and I_22735 (I389211,I389194,I870411);
DFFARX1 I_22736 (I389211,I2683,I388917,I389237,);
nor I_22737 (I388885,I389237,I389141);
not I_22738 (I389259,I389237);
nor I_22739 (I389276,I389259,I389050);
nor I_22740 (I389293,I388982,I389276);
DFFARX1 I_22741 (I389293,I2683,I388917,I388900,);
nor I_22742 (I389324,I389259,I389141);
nor I_22743 (I389341,I870390,I870399);
nor I_22744 (I388891,I389341,I389324);
not I_22745 (I389372,I389341);
nand I_22746 (I388894,I389101,I389372);
DFFARX1 I_22747 (I389341,I2683,I388917,I388906,);
DFFARX1 I_22748 (I389341,I2683,I388917,I388903,);
not I_22749 (I389461,I2690);
DFFARX1 I_22750 (I72756,I2683,I389461,I389487,);
DFFARX1 I_22751 (I389487,I2683,I389461,I389504,);
not I_22752 (I389453,I389504);
not I_22753 (I389526,I389487);
nand I_22754 (I389543,I72771,I72750);
and I_22755 (I389560,I389543,I72753);
DFFARX1 I_22756 (I389560,I2683,I389461,I389586,);
not I_22757 (I389594,I389586);
DFFARX1 I_22758 (I72759,I2683,I389461,I389620,);
and I_22759 (I389628,I389620,I72753);
nand I_22760 (I389645,I389620,I72753);
nand I_22761 (I389432,I389594,I389645);
DFFARX1 I_22762 (I72768,I2683,I389461,I389685,);
nor I_22763 (I389693,I389685,I389628);
DFFARX1 I_22764 (I389693,I2683,I389461,I389426,);
nor I_22765 (I389441,I389685,I389586);
nand I_22766 (I389738,I72750,I72765);
and I_22767 (I389755,I389738,I72762);
DFFARX1 I_22768 (I389755,I2683,I389461,I389781,);
nor I_22769 (I389429,I389781,I389685);
not I_22770 (I389803,I389781);
nor I_22771 (I389820,I389803,I389594);
nor I_22772 (I389837,I389526,I389820);
DFFARX1 I_22773 (I389837,I2683,I389461,I389444,);
nor I_22774 (I389868,I389803,I389685);
nor I_22775 (I389885,I72774,I72765);
nor I_22776 (I389435,I389885,I389868);
not I_22777 (I389916,I389885);
nand I_22778 (I389438,I389645,I389916);
DFFARX1 I_22779 (I389885,I2683,I389461,I389450,);
DFFARX1 I_22780 (I389885,I2683,I389461,I389447,);
not I_22781 (I390005,I2690);
DFFARX1 I_22782 (I692888,I2683,I390005,I390031,);
DFFARX1 I_22783 (I390031,I2683,I390005,I390048,);
not I_22784 (I389997,I390048);
not I_22785 (I390070,I390031);
nand I_22786 (I390087,I692882,I692879);
and I_22787 (I390104,I390087,I692894);
DFFARX1 I_22788 (I390104,I2683,I390005,I390130,);
not I_22789 (I390138,I390130);
DFFARX1 I_22790 (I692882,I2683,I390005,I390164,);
and I_22791 (I390172,I390164,I692876);
nand I_22792 (I390189,I390164,I692876);
nand I_22793 (I389976,I390138,I390189);
DFFARX1 I_22794 (I692876,I2683,I390005,I390229,);
nor I_22795 (I390237,I390229,I390172);
DFFARX1 I_22796 (I390237,I2683,I390005,I389970,);
nor I_22797 (I389985,I390229,I390130);
nand I_22798 (I390282,I692891,I692885);
and I_22799 (I390299,I390282,I692879);
DFFARX1 I_22800 (I390299,I2683,I390005,I390325,);
nor I_22801 (I389973,I390325,I390229);
not I_22802 (I390347,I390325);
nor I_22803 (I390364,I390347,I390138);
nor I_22804 (I390381,I390070,I390364);
DFFARX1 I_22805 (I390381,I2683,I390005,I389988,);
nor I_22806 (I390412,I390347,I390229);
nor I_22807 (I390429,I692897,I692885);
nor I_22808 (I389979,I390429,I390412);
not I_22809 (I390460,I390429);
nand I_22810 (I389982,I390189,I390460);
DFFARX1 I_22811 (I390429,I2683,I390005,I389994,);
DFFARX1 I_22812 (I390429,I2683,I390005,I389991,);
not I_22813 (I390549,I2690);
DFFARX1 I_22814 (I789765,I2683,I390549,I390575,);
DFFARX1 I_22815 (I390575,I2683,I390549,I390592,);
not I_22816 (I390541,I390592);
not I_22817 (I390614,I390575);
nand I_22818 (I390631,I789780,I789768);
and I_22819 (I390648,I390631,I789759);
DFFARX1 I_22820 (I390648,I2683,I390549,I390674,);
not I_22821 (I390682,I390674);
DFFARX1 I_22822 (I789771,I2683,I390549,I390708,);
and I_22823 (I390716,I390708,I789762);
nand I_22824 (I390733,I390708,I789762);
nand I_22825 (I390520,I390682,I390733);
DFFARX1 I_22826 (I789777,I2683,I390549,I390773,);
nor I_22827 (I390781,I390773,I390716);
DFFARX1 I_22828 (I390781,I2683,I390549,I390514,);
nor I_22829 (I390529,I390773,I390674);
nand I_22830 (I390826,I789786,I789774);
and I_22831 (I390843,I390826,I789783);
DFFARX1 I_22832 (I390843,I2683,I390549,I390869,);
nor I_22833 (I390517,I390869,I390773);
not I_22834 (I390891,I390869);
nor I_22835 (I390908,I390891,I390682);
nor I_22836 (I390925,I390614,I390908);
DFFARX1 I_22837 (I390925,I2683,I390549,I390532,);
nor I_22838 (I390956,I390891,I390773);
nor I_22839 (I390973,I789759,I789774);
nor I_22840 (I390523,I390973,I390956);
not I_22841 (I391004,I390973);
nand I_22842 (I390526,I390733,I391004);
DFFARX1 I_22843 (I390973,I2683,I390549,I390538,);
DFFARX1 I_22844 (I390973,I2683,I390549,I390535,);
not I_22845 (I391093,I2690);
DFFARX1 I_22846 (I747775,I2683,I391093,I391119,);
DFFARX1 I_22847 (I391119,I2683,I391093,I391136,);
not I_22848 (I391085,I391136);
not I_22849 (I391158,I391119);
nand I_22850 (I391175,I747790,I747778);
and I_22851 (I391192,I391175,I747769);
DFFARX1 I_22852 (I391192,I2683,I391093,I391218,);
not I_22853 (I391226,I391218);
DFFARX1 I_22854 (I747781,I2683,I391093,I391252,);
and I_22855 (I391260,I391252,I747772);
nand I_22856 (I391277,I391252,I747772);
nand I_22857 (I391064,I391226,I391277);
DFFARX1 I_22858 (I747787,I2683,I391093,I391317,);
nor I_22859 (I391325,I391317,I391260);
DFFARX1 I_22860 (I391325,I2683,I391093,I391058,);
nor I_22861 (I391073,I391317,I391218);
nand I_22862 (I391370,I747796,I747784);
and I_22863 (I391387,I391370,I747793);
DFFARX1 I_22864 (I391387,I2683,I391093,I391413,);
nor I_22865 (I391061,I391413,I391317);
not I_22866 (I391435,I391413);
nor I_22867 (I391452,I391435,I391226);
nor I_22868 (I391469,I391158,I391452);
DFFARX1 I_22869 (I391469,I2683,I391093,I391076,);
nor I_22870 (I391500,I391435,I391317);
nor I_22871 (I391517,I747769,I747784);
nor I_22872 (I391067,I391517,I391500);
not I_22873 (I391548,I391517);
nand I_22874 (I391070,I391277,I391548);
DFFARX1 I_22875 (I391517,I2683,I391093,I391082,);
DFFARX1 I_22876 (I391517,I2683,I391093,I391079,);
not I_22877 (I391637,I2690);
DFFARX1 I_22878 (I560721,I2683,I391637,I391663,);
DFFARX1 I_22879 (I391663,I2683,I391637,I391680,);
not I_22880 (I391629,I391680);
not I_22881 (I391702,I391663);
nand I_22882 (I391719,I560742,I560733);
and I_22883 (I391736,I391719,I560721);
DFFARX1 I_22884 (I391736,I2683,I391637,I391762,);
not I_22885 (I391770,I391762);
DFFARX1 I_22886 (I560727,I2683,I391637,I391796,);
and I_22887 (I391804,I391796,I560724);
nand I_22888 (I391821,I391796,I560724);
nand I_22889 (I391608,I391770,I391821);
DFFARX1 I_22890 (I560718,I2683,I391637,I391861,);
nor I_22891 (I391869,I391861,I391804);
DFFARX1 I_22892 (I391869,I2683,I391637,I391602,);
nor I_22893 (I391617,I391861,I391762);
nand I_22894 (I391914,I560718,I560730);
and I_22895 (I391931,I391914,I560739);
DFFARX1 I_22896 (I391931,I2683,I391637,I391957,);
nor I_22897 (I391605,I391957,I391861);
not I_22898 (I391979,I391957);
nor I_22899 (I391996,I391979,I391770);
nor I_22900 (I392013,I391702,I391996);
DFFARX1 I_22901 (I392013,I2683,I391637,I391620,);
nor I_22902 (I392044,I391979,I391861);
nor I_22903 (I392061,I560736,I560730);
nor I_22904 (I391611,I392061,I392044);
not I_22905 (I392092,I392061);
nand I_22906 (I391614,I391821,I392092);
DFFARX1 I_22907 (I392061,I2683,I391637,I391626,);
DFFARX1 I_22908 (I392061,I2683,I391637,I391623,);
not I_22909 (I392181,I2690);
DFFARX1 I_22910 (I425265,I2683,I392181,I392207,);
DFFARX1 I_22911 (I392207,I2683,I392181,I392224,);
not I_22912 (I392173,I392224);
not I_22913 (I392246,I392207);
nand I_22914 (I392263,I425268,I425286);
and I_22915 (I392280,I392263,I425274);
DFFARX1 I_22916 (I392280,I2683,I392181,I392306,);
not I_22917 (I392314,I392306);
DFFARX1 I_22918 (I425265,I2683,I392181,I392340,);
and I_22919 (I392348,I392340,I425283);
nand I_22920 (I392365,I392340,I425283);
nand I_22921 (I392152,I392314,I392365);
DFFARX1 I_22922 (I425277,I2683,I392181,I392405,);
nor I_22923 (I392413,I392405,I392348);
DFFARX1 I_22924 (I392413,I2683,I392181,I392146,);
nor I_22925 (I392161,I392405,I392306);
nand I_22926 (I392458,I425280,I425262);
and I_22927 (I392475,I392458,I425271);
DFFARX1 I_22928 (I392475,I2683,I392181,I392501,);
nor I_22929 (I392149,I392501,I392405);
not I_22930 (I392523,I392501);
nor I_22931 (I392540,I392523,I392314);
nor I_22932 (I392557,I392246,I392540);
DFFARX1 I_22933 (I392557,I2683,I392181,I392164,);
nor I_22934 (I392588,I392523,I392405);
nor I_22935 (I392605,I425262,I425262);
nor I_22936 (I392155,I392605,I392588);
not I_22937 (I392636,I392605);
nand I_22938 (I392158,I392365,I392636);
DFFARX1 I_22939 (I392605,I2683,I392181,I392170,);
DFFARX1 I_22940 (I392605,I2683,I392181,I392167,);
not I_22941 (I392725,I2690);
DFFARX1 I_22942 (I987489,I2683,I392725,I392751,);
DFFARX1 I_22943 (I392751,I2683,I392725,I392768,);
not I_22944 (I392717,I392768);
not I_22945 (I392790,I392751);
nand I_22946 (I392807,I987501,I987504);
and I_22947 (I392824,I392807,I987507);
DFFARX1 I_22948 (I392824,I2683,I392725,I392850,);
not I_22949 (I392858,I392850);
DFFARX1 I_22950 (I987492,I2683,I392725,I392884,);
and I_22951 (I392892,I392884,I987498);
nand I_22952 (I392909,I392884,I987498);
nand I_22953 (I392696,I392858,I392909);
DFFARX1 I_22954 (I987486,I2683,I392725,I392949,);
nor I_22955 (I392957,I392949,I392892);
DFFARX1 I_22956 (I392957,I2683,I392725,I392690,);
nor I_22957 (I392705,I392949,I392850);
nand I_22958 (I393002,I987489,I987510);
and I_22959 (I393019,I393002,I987495);
DFFARX1 I_22960 (I393019,I2683,I392725,I393045,);
nor I_22961 (I392693,I393045,I392949);
not I_22962 (I393067,I393045);
nor I_22963 (I393084,I393067,I392858);
nor I_22964 (I393101,I392790,I393084);
DFFARX1 I_22965 (I393101,I2683,I392725,I392708,);
nor I_22966 (I393132,I393067,I392949);
nor I_22967 (I393149,I987486,I987510);
nor I_22968 (I392699,I393149,I393132);
not I_22969 (I393180,I393149);
nand I_22970 (I392702,I392909,I393180);
DFFARX1 I_22971 (I393149,I2683,I392725,I392714,);
DFFARX1 I_22972 (I393149,I2683,I392725,I392711,);
not I_22973 (I393269,I2690);
DFFARX1 I_22974 (I235376,I2683,I393269,I393295,);
DFFARX1 I_22975 (I393295,I2683,I393269,I393312,);
not I_22976 (I393261,I393312);
not I_22977 (I393334,I393295);
nand I_22978 (I393351,I235355,I235379);
and I_22979 (I393368,I393351,I235382);
DFFARX1 I_22980 (I393368,I2683,I393269,I393394,);
not I_22981 (I393402,I393394);
DFFARX1 I_22982 (I235364,I2683,I393269,I393428,);
and I_22983 (I393436,I393428,I235370);
nand I_22984 (I393453,I393428,I235370);
nand I_22985 (I393240,I393402,I393453);
DFFARX1 I_22986 (I235358,I2683,I393269,I393493,);
nor I_22987 (I393501,I393493,I393436);
DFFARX1 I_22988 (I393501,I2683,I393269,I393234,);
nor I_22989 (I393249,I393493,I393394);
nand I_22990 (I393546,I235367,I235355);
and I_22991 (I393563,I393546,I235361);
DFFARX1 I_22992 (I393563,I2683,I393269,I393589,);
nor I_22993 (I393237,I393589,I393493);
not I_22994 (I393611,I393589);
nor I_22995 (I393628,I393611,I393402);
nor I_22996 (I393645,I393334,I393628);
DFFARX1 I_22997 (I393645,I2683,I393269,I393252,);
nor I_22998 (I393676,I393611,I393493);
nor I_22999 (I393693,I235373,I235355);
nor I_23000 (I393243,I393693,I393676);
not I_23001 (I393724,I393693);
nand I_23002 (I393246,I393453,I393724);
DFFARX1 I_23003 (I393693,I2683,I393269,I393258,);
DFFARX1 I_23004 (I393693,I2683,I393269,I393255,);
not I_23005 (I393813,I2690);
DFFARX1 I_23006 (I643877,I2683,I393813,I393839,);
DFFARX1 I_23007 (I393839,I2683,I393813,I393856,);
not I_23008 (I393805,I393856);
not I_23009 (I393878,I393839);
nand I_23010 (I393895,I643871,I643868);
and I_23011 (I393912,I393895,I643883);
DFFARX1 I_23012 (I393912,I2683,I393813,I393938,);
not I_23013 (I393946,I393938);
DFFARX1 I_23014 (I643871,I2683,I393813,I393972,);
and I_23015 (I393980,I393972,I643865);
nand I_23016 (I393997,I393972,I643865);
nand I_23017 (I393784,I393946,I393997);
DFFARX1 I_23018 (I643865,I2683,I393813,I394037,);
nor I_23019 (I394045,I394037,I393980);
DFFARX1 I_23020 (I394045,I2683,I393813,I393778,);
nor I_23021 (I393793,I394037,I393938);
nand I_23022 (I394090,I643880,I643874);
and I_23023 (I394107,I394090,I643868);
DFFARX1 I_23024 (I394107,I2683,I393813,I394133,);
nor I_23025 (I393781,I394133,I394037);
not I_23026 (I394155,I394133);
nor I_23027 (I394172,I394155,I393946);
nor I_23028 (I394189,I393878,I394172);
DFFARX1 I_23029 (I394189,I2683,I393813,I393796,);
nor I_23030 (I394220,I394155,I394037);
nor I_23031 (I394237,I643886,I643874);
nor I_23032 (I393787,I394237,I394220);
not I_23033 (I394268,I394237);
nand I_23034 (I393790,I393997,I394268);
DFFARX1 I_23035 (I394237,I2683,I393813,I393802,);
DFFARX1 I_23036 (I394237,I2683,I393813,I393799,);
not I_23037 (I394354,I2690);
DFFARX1 I_23038 (I256450,I2683,I394354,I394380,);
DFFARX1 I_23039 (I394380,I2683,I394354,I394397,);
not I_23040 (I394346,I394397);
DFFARX1 I_23041 (I256438,I2683,I394354,I394428,);
not I_23042 (I394436,I256441);
nor I_23043 (I394453,I394380,I394436);
not I_23044 (I394470,I256444);
not I_23045 (I394487,I256456);
nand I_23046 (I394504,I394487,I256444);
nor I_23047 (I394521,I394436,I394504);
nor I_23048 (I394538,I394428,I394521);
DFFARX1 I_23049 (I394487,I2683,I394354,I394343,);
nor I_23050 (I394569,I256456,I256447);
nand I_23051 (I394586,I394569,I256435);
nor I_23052 (I394603,I394586,I394470);
nand I_23053 (I394328,I394603,I256441);
DFFARX1 I_23054 (I394586,I2683,I394354,I394340,);
nand I_23055 (I394648,I394470,I256456);
nor I_23056 (I394665,I394470,I256456);
nand I_23057 (I394334,I394453,I394665);
not I_23058 (I394696,I256453);
nor I_23059 (I394713,I394696,I394648);
DFFARX1 I_23060 (I394713,I2683,I394354,I394322,);
nor I_23061 (I394744,I394696,I256459);
and I_23062 (I394761,I394744,I256462);
or I_23063 (I394778,I394761,I256435);
DFFARX1 I_23064 (I394778,I2683,I394354,I394804,);
nor I_23065 (I394812,I394804,I394428);
nor I_23066 (I394331,I394380,I394812);
not I_23067 (I394843,I394804);
nor I_23068 (I394860,I394843,I394538);
DFFARX1 I_23069 (I394860,I2683,I394354,I394337,);
nand I_23070 (I394891,I394843,I394470);
nor I_23071 (I394325,I394696,I394891);
not I_23072 (I394949,I2690);
DFFARX1 I_23073 (I127745,I2683,I394949,I394975,);
DFFARX1 I_23074 (I394975,I2683,I394949,I394992,);
not I_23075 (I394941,I394992);
DFFARX1 I_23076 (I127769,I2683,I394949,I395023,);
not I_23077 (I395031,I127763);
nor I_23078 (I395048,I394975,I395031);
not I_23079 (I395065,I127757);
not I_23080 (I395082,I127754);
nand I_23081 (I395099,I395082,I127757);
nor I_23082 (I395116,I395031,I395099);
nor I_23083 (I395133,I395023,I395116);
DFFARX1 I_23084 (I395082,I2683,I394949,I394938,);
nor I_23085 (I395164,I127754,I127748);
nand I_23086 (I395181,I395164,I127766);
nor I_23087 (I395198,I395181,I395065);
nand I_23088 (I394923,I395198,I127763);
DFFARX1 I_23089 (I395181,I2683,I394949,I394935,);
nand I_23090 (I395243,I395065,I127754);
nor I_23091 (I395260,I395065,I127754);
nand I_23092 (I394929,I395048,I395260);
not I_23093 (I395291,I127760);
nor I_23094 (I395308,I395291,I395243);
DFFARX1 I_23095 (I395308,I2683,I394949,I394917,);
nor I_23096 (I395339,I395291,I127745);
and I_23097 (I395356,I395339,I127751);
or I_23098 (I395373,I395356,I127748);
DFFARX1 I_23099 (I395373,I2683,I394949,I395399,);
nor I_23100 (I395407,I395399,I395023);
nor I_23101 (I394926,I394975,I395407);
not I_23102 (I395438,I395399);
nor I_23103 (I395455,I395438,I395133);
DFFARX1 I_23104 (I395455,I2683,I394949,I394932,);
nand I_23105 (I395486,I395438,I395065);
nor I_23106 (I394920,I395291,I395486);
not I_23107 (I395544,I2690);
DFFARX1 I_23108 (I319250,I2683,I395544,I395570,);
DFFARX1 I_23109 (I395570,I2683,I395544,I395587,);
not I_23110 (I395536,I395587);
DFFARX1 I_23111 (I319274,I2683,I395544,I395618,);
not I_23112 (I395626,I319253);
nor I_23113 (I395643,I395570,I395626);
not I_23114 (I395660,I319259);
not I_23115 (I395677,I319265);
nand I_23116 (I395694,I395677,I319259);
nor I_23117 (I395711,I395626,I395694);
nor I_23118 (I395728,I395618,I395711);
DFFARX1 I_23119 (I395677,I2683,I395544,I395533,);
nor I_23120 (I395759,I319265,I319277);
nand I_23121 (I395776,I395759,I319271);
nor I_23122 (I395793,I395776,I395660);
nand I_23123 (I395518,I395793,I319253);
DFFARX1 I_23124 (I395776,I2683,I395544,I395530,);
nand I_23125 (I395838,I395660,I319265);
nor I_23126 (I395855,I395660,I319265);
nand I_23127 (I395524,I395643,I395855);
not I_23128 (I395886,I319256);
nor I_23129 (I395903,I395886,I395838);
DFFARX1 I_23130 (I395903,I2683,I395544,I395512,);
nor I_23131 (I395934,I395886,I319250);
and I_23132 (I395951,I395934,I319268);
or I_23133 (I395968,I395951,I319262);
DFFARX1 I_23134 (I395968,I2683,I395544,I395994,);
nor I_23135 (I396002,I395994,I395618);
nor I_23136 (I395521,I395570,I396002);
not I_23137 (I396033,I395994);
nor I_23138 (I396050,I396033,I395728);
DFFARX1 I_23139 (I396050,I2683,I395544,I395527,);
nand I_23140 (I396081,I396033,I395660);
nor I_23141 (I395515,I395886,I396081);
not I_23142 (I396139,I2690);
DFFARX1 I_23143 (I573443,I2683,I396139,I396165,);
DFFARX1 I_23144 (I396165,I2683,I396139,I396182,);
not I_23145 (I396131,I396182);
DFFARX1 I_23146 (I573437,I2683,I396139,I396213,);
not I_23147 (I396221,I573434);
nor I_23148 (I396238,I396165,I396221);
not I_23149 (I396255,I573446);
not I_23150 (I396272,I573449);
nand I_23151 (I396289,I396272,I573446);
nor I_23152 (I396306,I396221,I396289);
nor I_23153 (I396323,I396213,I396306);
DFFARX1 I_23154 (I396272,I2683,I396139,I396128,);
nor I_23155 (I396354,I573449,I573458);
nand I_23156 (I396371,I396354,I573452);
nor I_23157 (I396388,I396371,I396255);
nand I_23158 (I396113,I396388,I573434);
DFFARX1 I_23159 (I396371,I2683,I396139,I396125,);
nand I_23160 (I396433,I396255,I573449);
nor I_23161 (I396450,I396255,I573449);
nand I_23162 (I396119,I396238,I396450);
not I_23163 (I396481,I573440);
nor I_23164 (I396498,I396481,I396433);
DFFARX1 I_23165 (I396498,I2683,I396139,I396107,);
nor I_23166 (I396529,I396481,I573455);
and I_23167 (I396546,I396529,I573434);
or I_23168 (I396563,I396546,I573437);
DFFARX1 I_23169 (I396563,I2683,I396139,I396589,);
nor I_23170 (I396597,I396589,I396213);
nor I_23171 (I396116,I396165,I396597);
not I_23172 (I396628,I396589);
nor I_23173 (I396645,I396628,I396323);
DFFARX1 I_23174 (I396645,I2683,I396139,I396122,);
nand I_23175 (I396676,I396628,I396255);
nor I_23176 (I396110,I396481,I396676);
not I_23177 (I396734,I2690);
DFFARX1 I_23178 (I692358,I2683,I396734,I396760,);
DFFARX1 I_23179 (I396760,I2683,I396734,I396777,);
not I_23180 (I396726,I396777);
DFFARX1 I_23181 (I692355,I2683,I396734,I396808,);
not I_23182 (I396816,I692355);
nor I_23183 (I396833,I396760,I396816);
not I_23184 (I396850,I692352);
not I_23185 (I396867,I692367);
nand I_23186 (I396884,I396867,I692352);
nor I_23187 (I396901,I396816,I396884);
nor I_23188 (I396918,I396808,I396901);
DFFARX1 I_23189 (I396867,I2683,I396734,I396723,);
nor I_23190 (I396949,I692367,I692361);
nand I_23191 (I396966,I396949,I692349);
nor I_23192 (I396983,I396966,I396850);
nand I_23193 (I396708,I396983,I692355);
DFFARX1 I_23194 (I396966,I2683,I396734,I396720,);
nand I_23195 (I397028,I396850,I692367);
nor I_23196 (I397045,I396850,I692367);
nand I_23197 (I396714,I396833,I397045);
not I_23198 (I397076,I692370);
nor I_23199 (I397093,I397076,I397028);
DFFARX1 I_23200 (I397093,I2683,I396734,I396702,);
nor I_23201 (I397124,I397076,I692349);
and I_23202 (I397141,I397124,I692364);
or I_23203 (I397158,I397141,I692352);
DFFARX1 I_23204 (I397158,I2683,I396734,I397184,);
nor I_23205 (I397192,I397184,I396808);
nor I_23206 (I396711,I396760,I397192);
not I_23207 (I397223,I397184);
nor I_23208 (I397240,I397223,I396918);
DFFARX1 I_23209 (I397240,I2683,I396734,I396717,);
nand I_23210 (I397271,I397223,I396850);
nor I_23211 (I396705,I397076,I397271);
not I_23212 (I397329,I2690);
DFFARX1 I_23213 (I102271,I2683,I397329,I397355,);
DFFARX1 I_23214 (I397355,I2683,I397329,I397372,);
not I_23215 (I397321,I397372);
DFFARX1 I_23216 (I102283,I2683,I397329,I397403,);
not I_23217 (I397411,I102274);
nor I_23218 (I397428,I397355,I397411);
not I_23219 (I397445,I102265);
not I_23220 (I397462,I102262);
nand I_23221 (I397479,I397462,I102265);
nor I_23222 (I397496,I397411,I397479);
nor I_23223 (I397513,I397403,I397496);
DFFARX1 I_23224 (I397462,I2683,I397329,I397318,);
nor I_23225 (I397544,I102262,I102262);
nand I_23226 (I397561,I397544,I102280);
nor I_23227 (I397578,I397561,I397445);
nand I_23228 (I397303,I397578,I102274);
DFFARX1 I_23229 (I397561,I2683,I397329,I397315,);
nand I_23230 (I397623,I397445,I102262);
nor I_23231 (I397640,I397445,I102262);
nand I_23232 (I397309,I397428,I397640);
not I_23233 (I397671,I102286);
nor I_23234 (I397688,I397671,I397623);
DFFARX1 I_23235 (I397688,I2683,I397329,I397297,);
nor I_23236 (I397719,I397671,I102265);
and I_23237 (I397736,I397719,I102268);
or I_23238 (I397753,I397736,I102277);
DFFARX1 I_23239 (I397753,I2683,I397329,I397779,);
nor I_23240 (I397787,I397779,I397403);
nor I_23241 (I397306,I397355,I397787);
not I_23242 (I397818,I397779);
nor I_23243 (I397835,I397818,I397513);
DFFARX1 I_23244 (I397835,I2683,I397329,I397312,);
nand I_23245 (I397866,I397818,I397445);
nor I_23246 (I397300,I397671,I397866);
not I_23247 (I397924,I2690);
DFFARX1 I_23248 (I908556,I2683,I397924,I397950,);
DFFARX1 I_23249 (I397950,I2683,I397924,I397967,);
not I_23250 (I397916,I397967);
DFFARX1 I_23251 (I908538,I2683,I397924,I397998,);
not I_23252 (I398006,I908544);
nor I_23253 (I398023,I397950,I398006);
not I_23254 (I398040,I908559);
not I_23255 (I398057,I908550);
nand I_23256 (I398074,I398057,I908559);
nor I_23257 (I398091,I398006,I398074);
nor I_23258 (I398108,I397998,I398091);
DFFARX1 I_23259 (I398057,I2683,I397924,I397913,);
nor I_23260 (I398139,I908550,I908562);
nand I_23261 (I398156,I398139,I908541);
nor I_23262 (I398173,I398156,I398040);
nand I_23263 (I397898,I398173,I908544);
DFFARX1 I_23264 (I398156,I2683,I397924,I397910,);
nand I_23265 (I398218,I398040,I908550);
nor I_23266 (I398235,I398040,I908550);
nand I_23267 (I397904,I398023,I398235);
not I_23268 (I398266,I908547);
nor I_23269 (I398283,I398266,I398218);
DFFARX1 I_23270 (I398283,I2683,I397924,I397892,);
nor I_23271 (I398314,I398266,I908553);
and I_23272 (I398331,I398314,I908538);
or I_23273 (I398348,I398331,I908541);
DFFARX1 I_23274 (I398348,I2683,I397924,I398374,);
nor I_23275 (I398382,I398374,I397998);
nor I_23276 (I397901,I397950,I398382);
not I_23277 (I398413,I398374);
nor I_23278 (I398430,I398413,I398108);
DFFARX1 I_23279 (I398430,I2683,I397924,I397907,);
nand I_23280 (I398461,I398413,I398040);
nor I_23281 (I397895,I398266,I398461);
not I_23282 (I398519,I2690);
DFFARX1 I_23283 (I928208,I2683,I398519,I398545,);
DFFARX1 I_23284 (I398545,I2683,I398519,I398562,);
not I_23285 (I398511,I398562);
DFFARX1 I_23286 (I928190,I2683,I398519,I398593,);
not I_23287 (I398601,I928196);
nor I_23288 (I398618,I398545,I398601);
not I_23289 (I398635,I928211);
not I_23290 (I398652,I928202);
nand I_23291 (I398669,I398652,I928211);
nor I_23292 (I398686,I398601,I398669);
nor I_23293 (I398703,I398593,I398686);
DFFARX1 I_23294 (I398652,I2683,I398519,I398508,);
nor I_23295 (I398734,I928202,I928214);
nand I_23296 (I398751,I398734,I928193);
nor I_23297 (I398768,I398751,I398635);
nand I_23298 (I398493,I398768,I928196);
DFFARX1 I_23299 (I398751,I2683,I398519,I398505,);
nand I_23300 (I398813,I398635,I928202);
nor I_23301 (I398830,I398635,I928202);
nand I_23302 (I398499,I398618,I398830);
not I_23303 (I398861,I928199);
nor I_23304 (I398878,I398861,I398813);
DFFARX1 I_23305 (I398878,I2683,I398519,I398487,);
nor I_23306 (I398909,I398861,I928205);
and I_23307 (I398926,I398909,I928190);
or I_23308 (I398943,I398926,I928193);
DFFARX1 I_23309 (I398943,I2683,I398519,I398969,);
nor I_23310 (I398977,I398969,I398593);
nor I_23311 (I398496,I398545,I398977);
not I_23312 (I399008,I398969);
nor I_23313 (I399025,I399008,I398703);
DFFARX1 I_23314 (I399025,I2683,I398519,I398502,);
nand I_23315 (I399056,I399008,I398635);
nor I_23316 (I398490,I398861,I399056);
not I_23317 (I399114,I2690);
DFFARX1 I_23318 (I954218,I2683,I399114,I399140,);
DFFARX1 I_23319 (I399140,I2683,I399114,I399157,);
not I_23320 (I399106,I399157);
DFFARX1 I_23321 (I954200,I2683,I399114,I399188,);
not I_23322 (I399196,I954206);
nor I_23323 (I399213,I399140,I399196);
not I_23324 (I399230,I954221);
not I_23325 (I399247,I954212);
nand I_23326 (I399264,I399247,I954221);
nor I_23327 (I399281,I399196,I399264);
nor I_23328 (I399298,I399188,I399281);
DFFARX1 I_23329 (I399247,I2683,I399114,I399103,);
nor I_23330 (I399329,I954212,I954224);
nand I_23331 (I399346,I399329,I954203);
nor I_23332 (I399363,I399346,I399230);
nand I_23333 (I399088,I399363,I954206);
DFFARX1 I_23334 (I399346,I2683,I399114,I399100,);
nand I_23335 (I399408,I399230,I954212);
nor I_23336 (I399425,I399230,I954212);
nand I_23337 (I399094,I399213,I399425);
not I_23338 (I399456,I954209);
nor I_23339 (I399473,I399456,I399408);
DFFARX1 I_23340 (I399473,I2683,I399114,I399082,);
nor I_23341 (I399504,I399456,I954215);
and I_23342 (I399521,I399504,I954200);
or I_23343 (I399538,I399521,I954203);
DFFARX1 I_23344 (I399538,I2683,I399114,I399564,);
nor I_23345 (I399572,I399564,I399188);
nor I_23346 (I399091,I399140,I399572);
not I_23347 (I399603,I399564);
nor I_23348 (I399620,I399603,I399298);
DFFARX1 I_23349 (I399620,I2683,I399114,I399097,);
nand I_23350 (I399651,I399603,I399230);
nor I_23351 (I399085,I399456,I399651);
not I_23352 (I399709,I2690);
DFFARX1 I_23353 (I1572,I2683,I399709,I399735,);
DFFARX1 I_23354 (I399735,I2683,I399709,I399752,);
not I_23355 (I399701,I399752);
DFFARX1 I_23356 (I1924,I2683,I399709,I399783,);
not I_23357 (I399791,I2068);
nor I_23358 (I399808,I399735,I399791);
not I_23359 (I399825,I2188);
not I_23360 (I399842,I2012);
nand I_23361 (I399859,I399842,I2188);
nor I_23362 (I399876,I399791,I399859);
nor I_23363 (I399893,I399783,I399876);
DFFARX1 I_23364 (I399842,I2683,I399709,I399698,);
nor I_23365 (I399924,I2012,I2060);
nand I_23366 (I399941,I399924,I1620);
nor I_23367 (I399958,I399941,I399825);
nand I_23368 (I399683,I399958,I2068);
DFFARX1 I_23369 (I399941,I2683,I399709,I399695,);
nand I_23370 (I400003,I399825,I2012);
nor I_23371 (I400020,I399825,I2012);
nand I_23372 (I399689,I399808,I400020);
not I_23373 (I400051,I1412);
nor I_23374 (I400068,I400051,I400003);
DFFARX1 I_23375 (I400068,I2683,I399709,I399677,);
nor I_23376 (I400099,I400051,I2332);
and I_23377 (I400116,I400099,I1916);
or I_23378 (I400133,I400116,I2676);
DFFARX1 I_23379 (I400133,I2683,I399709,I400159,);
nor I_23380 (I400167,I400159,I399783);
nor I_23381 (I399686,I399735,I400167);
not I_23382 (I400198,I400159);
nor I_23383 (I400215,I400198,I399893);
DFFARX1 I_23384 (I400215,I2683,I399709,I399692,);
nand I_23385 (I400246,I400198,I399825);
nor I_23386 (I399680,I400051,I400246);
not I_23387 (I400304,I2690);
DFFARX1 I_23388 (I73813,I2683,I400304,I400330,);
DFFARX1 I_23389 (I400330,I2683,I400304,I400347,);
not I_23390 (I400296,I400347);
DFFARX1 I_23391 (I73825,I2683,I400304,I400378,);
not I_23392 (I400386,I73816);
nor I_23393 (I400403,I400330,I400386);
not I_23394 (I400420,I73807);
not I_23395 (I400437,I73804);
nand I_23396 (I400454,I400437,I73807);
nor I_23397 (I400471,I400386,I400454);
nor I_23398 (I400488,I400378,I400471);
DFFARX1 I_23399 (I400437,I2683,I400304,I400293,);
nor I_23400 (I400519,I73804,I73804);
nand I_23401 (I400536,I400519,I73822);
nor I_23402 (I400553,I400536,I400420);
nand I_23403 (I400278,I400553,I73816);
DFFARX1 I_23404 (I400536,I2683,I400304,I400290,);
nand I_23405 (I400598,I400420,I73804);
nor I_23406 (I400615,I400420,I73804);
nand I_23407 (I400284,I400403,I400615);
not I_23408 (I400646,I73828);
nor I_23409 (I400663,I400646,I400598);
DFFARX1 I_23410 (I400663,I2683,I400304,I400272,);
nor I_23411 (I400694,I400646,I73807);
and I_23412 (I400711,I400694,I73810);
or I_23413 (I400728,I400711,I73819);
DFFARX1 I_23414 (I400728,I2683,I400304,I400754,);
nor I_23415 (I400762,I400754,I400378);
nor I_23416 (I400281,I400330,I400762);
not I_23417 (I400793,I400754);
nor I_23418 (I400810,I400793,I400488);
DFFARX1 I_23419 (I400810,I2683,I400304,I400287,);
nand I_23420 (I400841,I400793,I400420);
nor I_23421 (I400275,I400646,I400841);
not I_23422 (I400899,I2690);
DFFARX1 I_23423 (I560149,I2683,I400899,I400925,);
DFFARX1 I_23424 (I400925,I2683,I400899,I400942,);
not I_23425 (I400891,I400942);
DFFARX1 I_23426 (I560143,I2683,I400899,I400973,);
not I_23427 (I400981,I560140);
nor I_23428 (I400998,I400925,I400981);
not I_23429 (I401015,I560152);
not I_23430 (I401032,I560155);
nand I_23431 (I401049,I401032,I560152);
nor I_23432 (I401066,I400981,I401049);
nor I_23433 (I401083,I400973,I401066);
DFFARX1 I_23434 (I401032,I2683,I400899,I400888,);
nor I_23435 (I401114,I560155,I560164);
nand I_23436 (I401131,I401114,I560158);
nor I_23437 (I401148,I401131,I401015);
nand I_23438 (I400873,I401148,I560140);
DFFARX1 I_23439 (I401131,I2683,I400899,I400885,);
nand I_23440 (I401193,I401015,I560155);
nor I_23441 (I401210,I401015,I560155);
nand I_23442 (I400879,I400998,I401210);
not I_23443 (I401241,I560146);
nor I_23444 (I401258,I401241,I401193);
DFFARX1 I_23445 (I401258,I2683,I400899,I400867,);
nor I_23446 (I401289,I401241,I560161);
and I_23447 (I401306,I401289,I560140);
or I_23448 (I401323,I401306,I560143);
DFFARX1 I_23449 (I401323,I2683,I400899,I401349,);
nor I_23450 (I401357,I401349,I400973);
nor I_23451 (I400876,I400925,I401357);
not I_23452 (I401388,I401349);
nor I_23453 (I401405,I401388,I401083);
DFFARX1 I_23454 (I401405,I2683,I400899,I400882,);
nand I_23455 (I401436,I401388,I401015);
nor I_23456 (I400870,I401241,I401436);
not I_23457 (I401494,I2690);
DFFARX1 I_23458 (I256977,I2683,I401494,I401520,);
DFFARX1 I_23459 (I401520,I2683,I401494,I401537,);
not I_23460 (I401486,I401537);
DFFARX1 I_23461 (I256965,I2683,I401494,I401568,);
not I_23462 (I401576,I256968);
nor I_23463 (I401593,I401520,I401576);
not I_23464 (I401610,I256971);
not I_23465 (I401627,I256983);
nand I_23466 (I401644,I401627,I256971);
nor I_23467 (I401661,I401576,I401644);
nor I_23468 (I401678,I401568,I401661);
DFFARX1 I_23469 (I401627,I2683,I401494,I401483,);
nor I_23470 (I401709,I256983,I256974);
nand I_23471 (I401726,I401709,I256962);
nor I_23472 (I401743,I401726,I401610);
nand I_23473 (I401468,I401743,I256968);
DFFARX1 I_23474 (I401726,I2683,I401494,I401480,);
nand I_23475 (I401788,I401610,I256983);
nor I_23476 (I401805,I401610,I256983);
nand I_23477 (I401474,I401593,I401805);
not I_23478 (I401836,I256980);
nor I_23479 (I401853,I401836,I401788);
DFFARX1 I_23480 (I401853,I2683,I401494,I401462,);
nor I_23481 (I401884,I401836,I256986);
and I_23482 (I401901,I401884,I256989);
or I_23483 (I401918,I401901,I256962);
DFFARX1 I_23484 (I401918,I2683,I401494,I401944,);
nor I_23485 (I401952,I401944,I401568);
nor I_23486 (I401471,I401520,I401952);
not I_23487 (I401983,I401944);
nor I_23488 (I402000,I401983,I401678);
DFFARX1 I_23489 (I402000,I2683,I401494,I401477,);
nand I_23490 (I402031,I401983,I401610);
nor I_23491 (I401465,I401836,I402031);
not I_23492 (I402089,I2690);
DFFARX1 I_23493 (I889482,I2683,I402089,I402115,);
DFFARX1 I_23494 (I402115,I2683,I402089,I402132,);
not I_23495 (I402081,I402132);
DFFARX1 I_23496 (I889464,I2683,I402089,I402163,);
not I_23497 (I402171,I889470);
nor I_23498 (I402188,I402115,I402171);
not I_23499 (I402205,I889485);
not I_23500 (I402222,I889476);
nand I_23501 (I402239,I402222,I889485);
nor I_23502 (I402256,I402171,I402239);
nor I_23503 (I402273,I402163,I402256);
DFFARX1 I_23504 (I402222,I2683,I402089,I402078,);
nor I_23505 (I402304,I889476,I889488);
nand I_23506 (I402321,I402304,I889467);
nor I_23507 (I402338,I402321,I402205);
nand I_23508 (I402063,I402338,I889470);
DFFARX1 I_23509 (I402321,I2683,I402089,I402075,);
nand I_23510 (I402383,I402205,I889476);
nor I_23511 (I402400,I402205,I889476);
nand I_23512 (I402069,I402188,I402400);
not I_23513 (I402431,I889473);
nor I_23514 (I402448,I402431,I402383);
DFFARX1 I_23515 (I402448,I2683,I402089,I402057,);
nor I_23516 (I402479,I402431,I889479);
and I_23517 (I402496,I402479,I889464);
or I_23518 (I402513,I402496,I889467);
DFFARX1 I_23519 (I402513,I2683,I402089,I402539,);
nor I_23520 (I402547,I402539,I402163);
nor I_23521 (I402066,I402115,I402547);
not I_23522 (I402578,I402539);
nor I_23523 (I402595,I402578,I402273);
DFFARX1 I_23524 (I402595,I2683,I402089,I402072,);
nand I_23525 (I402626,I402578,I402205);
nor I_23526 (I402060,I402431,I402626);
not I_23527 (I402684,I2690);
DFFARX1 I_23528 (I297029,I2683,I402684,I402710,);
DFFARX1 I_23529 (I402710,I2683,I402684,I402727,);
not I_23530 (I402676,I402727);
DFFARX1 I_23531 (I297017,I2683,I402684,I402758,);
not I_23532 (I402766,I297020);
nor I_23533 (I402783,I402710,I402766);
not I_23534 (I402800,I297023);
not I_23535 (I402817,I297035);
nand I_23536 (I402834,I402817,I297023);
nor I_23537 (I402851,I402766,I402834);
nor I_23538 (I402868,I402758,I402851);
DFFARX1 I_23539 (I402817,I2683,I402684,I402673,);
nor I_23540 (I402899,I297035,I297026);
nand I_23541 (I402916,I402899,I297014);
nor I_23542 (I402933,I402916,I402800);
nand I_23543 (I402658,I402933,I297020);
DFFARX1 I_23544 (I402916,I2683,I402684,I402670,);
nand I_23545 (I402978,I402800,I297035);
nor I_23546 (I402995,I402800,I297035);
nand I_23547 (I402664,I402783,I402995);
not I_23548 (I403026,I297032);
nor I_23549 (I403043,I403026,I402978);
DFFARX1 I_23550 (I403043,I2683,I402684,I402652,);
nor I_23551 (I403074,I403026,I297038);
and I_23552 (I403091,I403074,I297041);
or I_23553 (I403108,I403091,I297014);
DFFARX1 I_23554 (I403108,I2683,I402684,I403134,);
nor I_23555 (I403142,I403134,I402758);
nor I_23556 (I402661,I402710,I403142);
not I_23557 (I403173,I403134);
nor I_23558 (I403190,I403173,I402868);
DFFARX1 I_23559 (I403190,I2683,I402684,I402667,);
nand I_23560 (I403221,I403173,I402800);
nor I_23561 (I402655,I403026,I403221);
not I_23562 (I403279,I2690);
DFFARX1 I_23563 (I933988,I2683,I403279,I403305,);
DFFARX1 I_23564 (I403305,I2683,I403279,I403322,);
not I_23565 (I403271,I403322);
DFFARX1 I_23566 (I933970,I2683,I403279,I403353,);
not I_23567 (I403361,I933976);
nor I_23568 (I403378,I403305,I403361);
not I_23569 (I403395,I933991);
not I_23570 (I403412,I933982);
nand I_23571 (I403429,I403412,I933991);
nor I_23572 (I403446,I403361,I403429);
nor I_23573 (I403463,I403353,I403446);
DFFARX1 I_23574 (I403412,I2683,I403279,I403268,);
nor I_23575 (I403494,I933982,I933994);
nand I_23576 (I403511,I403494,I933973);
nor I_23577 (I403528,I403511,I403395);
nand I_23578 (I403253,I403528,I933976);
DFFARX1 I_23579 (I403511,I2683,I403279,I403265,);
nand I_23580 (I403573,I403395,I933982);
nor I_23581 (I403590,I403395,I933982);
nand I_23582 (I403259,I403378,I403590);
not I_23583 (I403621,I933979);
nor I_23584 (I403638,I403621,I403573);
DFFARX1 I_23585 (I403638,I2683,I403279,I403247,);
nor I_23586 (I403669,I403621,I933985);
and I_23587 (I403686,I403669,I933970);
or I_23588 (I403703,I403686,I933973);
DFFARX1 I_23589 (I403703,I2683,I403279,I403729,);
nor I_23590 (I403737,I403729,I403353);
nor I_23591 (I403256,I403305,I403737);
not I_23592 (I403768,I403729);
nor I_23593 (I403785,I403768,I403463);
DFFARX1 I_23594 (I403785,I2683,I403279,I403262,);
nand I_23595 (I403816,I403768,I403395);
nor I_23596 (I403250,I403621,I403816);
not I_23597 (I403874,I2690);
DFFARX1 I_23598 (I775562,I2683,I403874,I403900,);
DFFARX1 I_23599 (I403900,I2683,I403874,I403917,);
not I_23600 (I403866,I403917);
DFFARX1 I_23601 (I775550,I2683,I403874,I403948,);
not I_23602 (I403956,I775547);
nor I_23603 (I403973,I403900,I403956);
not I_23604 (I403990,I775559);
not I_23605 (I404007,I775556);
nand I_23606 (I404024,I404007,I775559);
nor I_23607 (I404041,I403956,I404024);
nor I_23608 (I404058,I403948,I404041);
DFFARX1 I_23609 (I404007,I2683,I403874,I403863,);
nor I_23610 (I404089,I775556,I775565);
nand I_23611 (I404106,I404089,I775568);
nor I_23612 (I404123,I404106,I403990);
nand I_23613 (I403848,I404123,I775547);
DFFARX1 I_23614 (I404106,I2683,I403874,I403860,);
nand I_23615 (I404168,I403990,I775556);
nor I_23616 (I404185,I403990,I775556);
nand I_23617 (I403854,I403973,I404185);
not I_23618 (I404216,I775571);
nor I_23619 (I404233,I404216,I404168);
DFFARX1 I_23620 (I404233,I2683,I403874,I403842,);
nor I_23621 (I404264,I404216,I775574);
and I_23622 (I404281,I404264,I775553);
or I_23623 (I404298,I404281,I775547);
DFFARX1 I_23624 (I404298,I2683,I403874,I404324,);
nor I_23625 (I404332,I404324,I403948);
nor I_23626 (I403851,I403900,I404332);
not I_23627 (I404363,I404324);
nor I_23628 (I404380,I404363,I404058);
DFFARX1 I_23629 (I404380,I2683,I403874,I403857,);
nand I_23630 (I404411,I404363,I403990);
nor I_23631 (I403845,I404216,I404411);
not I_23632 (I404469,I2690);
DFFARX1 I_23633 (I1081054,I2683,I404469,I404495,);
DFFARX1 I_23634 (I404495,I2683,I404469,I404512,);
not I_23635 (I404461,I404512);
DFFARX1 I_23636 (I1081060,I2683,I404469,I404543,);
not I_23637 (I404551,I1081075);
nor I_23638 (I404568,I404495,I404551);
not I_23639 (I404585,I1081066);
not I_23640 (I404602,I1081063);
nand I_23641 (I404619,I404602,I1081066);
nor I_23642 (I404636,I404551,I404619);
nor I_23643 (I404653,I404543,I404636);
DFFARX1 I_23644 (I404602,I2683,I404469,I404458,);
nor I_23645 (I404684,I1081063,I1081054);
nand I_23646 (I404701,I404684,I1081078);
nor I_23647 (I404718,I404701,I404585);
nand I_23648 (I404443,I404718,I1081075);
DFFARX1 I_23649 (I404701,I2683,I404469,I404455,);
nand I_23650 (I404763,I404585,I1081063);
nor I_23651 (I404780,I404585,I1081063);
nand I_23652 (I404449,I404568,I404780);
not I_23653 (I404811,I1081072);
nor I_23654 (I404828,I404811,I404763);
DFFARX1 I_23655 (I404828,I2683,I404469,I404437,);
nor I_23656 (I404859,I404811,I1081057);
and I_23657 (I404876,I404859,I1081069);
or I_23658 (I404893,I404876,I1081081);
DFFARX1 I_23659 (I404893,I2683,I404469,I404919,);
nor I_23660 (I404927,I404919,I404543);
nor I_23661 (I404446,I404495,I404927);
not I_23662 (I404958,I404919);
nor I_23663 (I404975,I404958,I404653);
DFFARX1 I_23664 (I404975,I2683,I404469,I404452,);
nand I_23665 (I405006,I404958,I404585);
nor I_23666 (I404440,I404811,I405006);
not I_23667 (I405064,I2690);
DFFARX1 I_23668 (I1065584,I2683,I405064,I405090,);
DFFARX1 I_23669 (I405090,I2683,I405064,I405107,);
not I_23670 (I405056,I405107);
DFFARX1 I_23671 (I1065590,I2683,I405064,I405138,);
not I_23672 (I405146,I1065605);
nor I_23673 (I405163,I405090,I405146);
not I_23674 (I405180,I1065596);
not I_23675 (I405197,I1065593);
nand I_23676 (I405214,I405197,I1065596);
nor I_23677 (I405231,I405146,I405214);
nor I_23678 (I405248,I405138,I405231);
DFFARX1 I_23679 (I405197,I2683,I405064,I405053,);
nor I_23680 (I405279,I1065593,I1065584);
nand I_23681 (I405296,I405279,I1065608);
nor I_23682 (I405313,I405296,I405180);
nand I_23683 (I405038,I405313,I1065605);
DFFARX1 I_23684 (I405296,I2683,I405064,I405050,);
nand I_23685 (I405358,I405180,I1065593);
nor I_23686 (I405375,I405180,I1065593);
nand I_23687 (I405044,I405163,I405375);
not I_23688 (I405406,I1065602);
nor I_23689 (I405423,I405406,I405358);
DFFARX1 I_23690 (I405423,I2683,I405064,I405032,);
nor I_23691 (I405454,I405406,I1065587);
and I_23692 (I405471,I405454,I1065599);
or I_23693 (I405488,I405471,I1065611);
DFFARX1 I_23694 (I405488,I2683,I405064,I405514,);
nor I_23695 (I405522,I405514,I405138);
nor I_23696 (I405041,I405090,I405522);
not I_23697 (I405553,I405514);
nor I_23698 (I405570,I405553,I405248);
DFFARX1 I_23699 (I405570,I2683,I405064,I405047,);
nand I_23700 (I405601,I405553,I405180);
nor I_23701 (I405035,I405406,I405601);
not I_23702 (I405659,I2690);
DFFARX1 I_23703 (I582113,I2683,I405659,I405685,);
DFFARX1 I_23704 (I405685,I2683,I405659,I405702,);
not I_23705 (I405651,I405702);
DFFARX1 I_23706 (I582107,I2683,I405659,I405733,);
not I_23707 (I405741,I582104);
nor I_23708 (I405758,I405685,I405741);
not I_23709 (I405775,I582116);
not I_23710 (I405792,I582119);
nand I_23711 (I405809,I405792,I582116);
nor I_23712 (I405826,I405741,I405809);
nor I_23713 (I405843,I405733,I405826);
DFFARX1 I_23714 (I405792,I2683,I405659,I405648,);
nor I_23715 (I405874,I582119,I582128);
nand I_23716 (I405891,I405874,I582122);
nor I_23717 (I405908,I405891,I405775);
nand I_23718 (I405633,I405908,I582104);
DFFARX1 I_23719 (I405891,I2683,I405659,I405645,);
nand I_23720 (I405953,I405775,I582119);
nor I_23721 (I405970,I405775,I582119);
nand I_23722 (I405639,I405758,I405970);
not I_23723 (I406001,I582110);
nor I_23724 (I406018,I406001,I405953);
DFFARX1 I_23725 (I406018,I2683,I405659,I405627,);
nor I_23726 (I406049,I406001,I582125);
and I_23727 (I406066,I406049,I582104);
or I_23728 (I406083,I406066,I582107);
DFFARX1 I_23729 (I406083,I2683,I405659,I406109,);
nor I_23730 (I406117,I406109,I405733);
nor I_23731 (I405636,I405685,I406117);
not I_23732 (I406148,I406109);
nor I_23733 (I406165,I406148,I405843);
DFFARX1 I_23734 (I406165,I2683,I405659,I405642,);
nand I_23735 (I406196,I406148,I405775);
nor I_23736 (I405630,I406001,I406196);
not I_23737 (I406254,I2690);
DFFARX1 I_23738 (I565929,I2683,I406254,I406280,);
DFFARX1 I_23739 (I406280,I2683,I406254,I406297,);
not I_23740 (I406246,I406297);
DFFARX1 I_23741 (I565923,I2683,I406254,I406328,);
not I_23742 (I406336,I565920);
nor I_23743 (I406353,I406280,I406336);
not I_23744 (I406370,I565932);
not I_23745 (I406387,I565935);
nand I_23746 (I406404,I406387,I565932);
nor I_23747 (I406421,I406336,I406404);
nor I_23748 (I406438,I406328,I406421);
DFFARX1 I_23749 (I406387,I2683,I406254,I406243,);
nor I_23750 (I406469,I565935,I565944);
nand I_23751 (I406486,I406469,I565938);
nor I_23752 (I406503,I406486,I406370);
nand I_23753 (I406228,I406503,I565920);
DFFARX1 I_23754 (I406486,I2683,I406254,I406240,);
nand I_23755 (I406548,I406370,I565935);
nor I_23756 (I406565,I406370,I565935);
nand I_23757 (I406234,I406353,I406565);
not I_23758 (I406596,I565926);
nor I_23759 (I406613,I406596,I406548);
DFFARX1 I_23760 (I406613,I2683,I406254,I406222,);
nor I_23761 (I406644,I406596,I565941);
and I_23762 (I406661,I406644,I565920);
or I_23763 (I406678,I406661,I565923);
DFFARX1 I_23764 (I406678,I2683,I406254,I406704,);
nor I_23765 (I406712,I406704,I406328);
nor I_23766 (I406231,I406280,I406712);
not I_23767 (I406743,I406704);
nor I_23768 (I406760,I406743,I406438);
DFFARX1 I_23769 (I406760,I2683,I406254,I406237,);
nand I_23770 (I406791,I406743,I406370);
nor I_23771 (I406225,I406596,I406791);
not I_23772 (I406849,I2690);
DFFARX1 I_23773 (I36387,I2683,I406849,I406875,);
DFFARX1 I_23774 (I406875,I2683,I406849,I406892,);
not I_23775 (I406841,I406892);
DFFARX1 I_23776 (I36387,I2683,I406849,I406923,);
not I_23777 (I406931,I36402);
nor I_23778 (I406948,I406875,I406931);
not I_23779 (I406965,I36405);
not I_23780 (I406982,I36396);
nand I_23781 (I406999,I406982,I36405);
nor I_23782 (I407016,I406931,I406999);
nor I_23783 (I407033,I406923,I407016);
DFFARX1 I_23784 (I406982,I2683,I406849,I406838,);
nor I_23785 (I407064,I36396,I36408);
nand I_23786 (I407081,I407064,I36390);
nor I_23787 (I407098,I407081,I406965);
nand I_23788 (I406823,I407098,I36402);
DFFARX1 I_23789 (I407081,I2683,I406849,I406835,);
nand I_23790 (I407143,I406965,I36396);
nor I_23791 (I407160,I406965,I36396);
nand I_23792 (I406829,I406948,I407160);
not I_23793 (I407191,I36390);
nor I_23794 (I407208,I407191,I407143);
DFFARX1 I_23795 (I407208,I2683,I406849,I406817,);
nor I_23796 (I407239,I407191,I36399);
and I_23797 (I407256,I407239,I36393);
or I_23798 (I407273,I407256,I36411);
DFFARX1 I_23799 (I407273,I2683,I406849,I407299,);
nor I_23800 (I407307,I407299,I406923);
nor I_23801 (I406826,I406875,I407307);
not I_23802 (I407338,I407299);
nor I_23803 (I407355,I407338,I407033);
DFFARX1 I_23804 (I407355,I2683,I406849,I406832,);
nand I_23805 (I407386,I407338,I406965);
nor I_23806 (I406820,I407191,I407386);
not I_23807 (I407444,I2690);
DFFARX1 I_23808 (I147380,I2683,I407444,I407470,);
DFFARX1 I_23809 (I407470,I2683,I407444,I407487,);
not I_23810 (I407436,I407487);
DFFARX1 I_23811 (I147404,I2683,I407444,I407518,);
not I_23812 (I407526,I147398);
nor I_23813 (I407543,I407470,I407526);
not I_23814 (I407560,I147392);
not I_23815 (I407577,I147389);
nand I_23816 (I407594,I407577,I147392);
nor I_23817 (I407611,I407526,I407594);
nor I_23818 (I407628,I407518,I407611);
DFFARX1 I_23819 (I407577,I2683,I407444,I407433,);
nor I_23820 (I407659,I147389,I147383);
nand I_23821 (I407676,I407659,I147401);
nor I_23822 (I407693,I407676,I407560);
nand I_23823 (I407418,I407693,I147398);
DFFARX1 I_23824 (I407676,I2683,I407444,I407430,);
nand I_23825 (I407738,I407560,I147389);
nor I_23826 (I407755,I407560,I147389);
nand I_23827 (I407424,I407543,I407755);
not I_23828 (I407786,I147395);
nor I_23829 (I407803,I407786,I407738);
DFFARX1 I_23830 (I407803,I2683,I407444,I407412,);
nor I_23831 (I407834,I407786,I147380);
and I_23832 (I407851,I407834,I147386);
or I_23833 (I407868,I407851,I147383);
DFFARX1 I_23834 (I407868,I2683,I407444,I407894,);
nor I_23835 (I407902,I407894,I407518);
nor I_23836 (I407421,I407470,I407902);
not I_23837 (I407933,I407894);
nor I_23838 (I407950,I407933,I407628);
DFFARX1 I_23839 (I407950,I2683,I407444,I407427,);
nand I_23840 (I407981,I407933,I407560);
nor I_23841 (I407415,I407786,I407981);
not I_23842 (I408039,I2690);
DFFARX1 I_23843 (I556103,I2683,I408039,I408065,);
DFFARX1 I_23844 (I408065,I2683,I408039,I408082,);
not I_23845 (I408031,I408082);
DFFARX1 I_23846 (I556097,I2683,I408039,I408113,);
not I_23847 (I408121,I556094);
nor I_23848 (I408138,I408065,I408121);
not I_23849 (I408155,I556106);
not I_23850 (I408172,I556109);
nand I_23851 (I408189,I408172,I556106);
nor I_23852 (I408206,I408121,I408189);
nor I_23853 (I408223,I408113,I408206);
DFFARX1 I_23854 (I408172,I2683,I408039,I408028,);
nor I_23855 (I408254,I556109,I556118);
nand I_23856 (I408271,I408254,I556112);
nor I_23857 (I408288,I408271,I408155);
nand I_23858 (I408013,I408288,I556094);
DFFARX1 I_23859 (I408271,I2683,I408039,I408025,);
nand I_23860 (I408333,I408155,I556109);
nor I_23861 (I408350,I408155,I556109);
nand I_23862 (I408019,I408138,I408350);
not I_23863 (I408381,I556100);
nor I_23864 (I408398,I408381,I408333);
DFFARX1 I_23865 (I408398,I2683,I408039,I408007,);
nor I_23866 (I408429,I408381,I556115);
and I_23867 (I408446,I408429,I556094);
or I_23868 (I408463,I408446,I556097);
DFFARX1 I_23869 (I408463,I2683,I408039,I408489,);
nor I_23870 (I408497,I408489,I408113);
nor I_23871 (I408016,I408065,I408497);
not I_23872 (I408528,I408489);
nor I_23873 (I408545,I408528,I408223);
DFFARX1 I_23874 (I408545,I2683,I408039,I408022,);
nand I_23875 (I408576,I408528,I408155);
nor I_23876 (I408010,I408381,I408576);
not I_23877 (I408634,I2690);
DFFARX1 I_23878 (I784606,I2683,I408634,I408660,);
DFFARX1 I_23879 (I408660,I2683,I408634,I408677,);
not I_23880 (I408626,I408677);
DFFARX1 I_23881 (I784594,I2683,I408634,I408708,);
not I_23882 (I408716,I784591);
nor I_23883 (I408733,I408660,I408716);
not I_23884 (I408750,I784603);
not I_23885 (I408767,I784600);
nand I_23886 (I408784,I408767,I784603);
nor I_23887 (I408801,I408716,I408784);
nor I_23888 (I408818,I408708,I408801);
DFFARX1 I_23889 (I408767,I2683,I408634,I408623,);
nor I_23890 (I408849,I784600,I784609);
nand I_23891 (I408866,I408849,I784612);
nor I_23892 (I408883,I408866,I408750);
nand I_23893 (I408608,I408883,I784591);
DFFARX1 I_23894 (I408866,I2683,I408634,I408620,);
nand I_23895 (I408928,I408750,I784600);
nor I_23896 (I408945,I408750,I784600);
nand I_23897 (I408614,I408733,I408945);
not I_23898 (I408976,I784615);
nor I_23899 (I408993,I408976,I408928);
DFFARX1 I_23900 (I408993,I2683,I408634,I408602,);
nor I_23901 (I409024,I408976,I784618);
and I_23902 (I409041,I409024,I784597);
or I_23903 (I409058,I409041,I784591);
DFFARX1 I_23904 (I409058,I2683,I408634,I409084,);
nor I_23905 (I409092,I409084,I408708);
nor I_23906 (I408611,I408660,I409092);
not I_23907 (I409123,I409084);
nor I_23908 (I409140,I409123,I408818);
DFFARX1 I_23909 (I409140,I2683,I408634,I408617,);
nand I_23910 (I409171,I409123,I408750);
nor I_23911 (I408605,I408976,I409171);
not I_23912 (I409229,I2690);
DFFARX1 I_23913 (I460727,I2683,I409229,I409255,);
DFFARX1 I_23914 (I409255,I2683,I409229,I409272,);
not I_23915 (I409221,I409272);
DFFARX1 I_23916 (I460739,I2683,I409229,I409303,);
not I_23917 (I409311,I460724);
nor I_23918 (I409328,I409255,I409311);
not I_23919 (I409345,I460742);
not I_23920 (I409362,I460733);
nand I_23921 (I409379,I409362,I460742);
nor I_23922 (I409396,I409311,I409379);
nor I_23923 (I409413,I409303,I409396);
DFFARX1 I_23924 (I409362,I2683,I409229,I409218,);
nor I_23925 (I409444,I460733,I460745);
nand I_23926 (I409461,I409444,I460748);
nor I_23927 (I409478,I409461,I409345);
nand I_23928 (I409203,I409478,I460724);
DFFARX1 I_23929 (I409461,I2683,I409229,I409215,);
nand I_23930 (I409523,I409345,I460733);
nor I_23931 (I409540,I409345,I460733);
nand I_23932 (I409209,I409328,I409540);
not I_23933 (I409571,I460724);
nor I_23934 (I409588,I409571,I409523);
DFFARX1 I_23935 (I409588,I2683,I409229,I409197,);
nor I_23936 (I409619,I409571,I460736);
and I_23937 (I409636,I409619,I460730);
or I_23938 (I409653,I409636,I460727);
DFFARX1 I_23939 (I409653,I2683,I409229,I409679,);
nor I_23940 (I409687,I409679,I409303);
nor I_23941 (I409206,I409255,I409687);
not I_23942 (I409718,I409679);
nor I_23943 (I409735,I409718,I409413);
DFFARX1 I_23944 (I409735,I2683,I409229,I409212,);
nand I_23945 (I409766,I409718,I409345);
nor I_23946 (I409200,I409571,I409766);
not I_23947 (I409824,I2690);
DFFARX1 I_23948 (I675494,I2683,I409824,I409850,);
DFFARX1 I_23949 (I409850,I2683,I409824,I409867,);
not I_23950 (I409816,I409867);
DFFARX1 I_23951 (I675491,I2683,I409824,I409898,);
not I_23952 (I409906,I675491);
nor I_23953 (I409923,I409850,I409906);
not I_23954 (I409940,I675488);
not I_23955 (I409957,I675503);
nand I_23956 (I409974,I409957,I675488);
nor I_23957 (I409991,I409906,I409974);
nor I_23958 (I410008,I409898,I409991);
DFFARX1 I_23959 (I409957,I2683,I409824,I409813,);
nor I_23960 (I410039,I675503,I675497);
nand I_23961 (I410056,I410039,I675485);
nor I_23962 (I410073,I410056,I409940);
nand I_23963 (I409798,I410073,I675491);
DFFARX1 I_23964 (I410056,I2683,I409824,I409810,);
nand I_23965 (I410118,I409940,I675503);
nor I_23966 (I410135,I409940,I675503);
nand I_23967 (I409804,I409923,I410135);
not I_23968 (I410166,I675506);
nor I_23969 (I410183,I410166,I410118);
DFFARX1 I_23970 (I410183,I2683,I409824,I409792,);
nor I_23971 (I410214,I410166,I675485);
and I_23972 (I410231,I410214,I675500);
or I_23973 (I410248,I410231,I675488);
DFFARX1 I_23974 (I410248,I2683,I409824,I410274,);
nor I_23975 (I410282,I410274,I409898);
nor I_23976 (I409801,I409850,I410282);
not I_23977 (I410313,I410274);
nor I_23978 (I410330,I410313,I410008);
DFFARX1 I_23979 (I410330,I2683,I409824,I409807,);
nand I_23980 (I410361,I410313,I409940);
nor I_23981 (I409795,I410166,I410361);
not I_23982 (I410419,I2690);
DFFARX1 I_23983 (I261193,I2683,I410419,I410445,);
DFFARX1 I_23984 (I410445,I2683,I410419,I410462,);
not I_23985 (I410411,I410462);
DFFARX1 I_23986 (I261181,I2683,I410419,I410493,);
not I_23987 (I410501,I261184);
nor I_23988 (I410518,I410445,I410501);
not I_23989 (I410535,I261187);
not I_23990 (I410552,I261199);
nand I_23991 (I410569,I410552,I261187);
nor I_23992 (I410586,I410501,I410569);
nor I_23993 (I410603,I410493,I410586);
DFFARX1 I_23994 (I410552,I2683,I410419,I410408,);
nor I_23995 (I410634,I261199,I261190);
nand I_23996 (I410651,I410634,I261178);
nor I_23997 (I410668,I410651,I410535);
nand I_23998 (I410393,I410668,I261184);
DFFARX1 I_23999 (I410651,I2683,I410419,I410405,);
nand I_24000 (I410713,I410535,I261199);
nor I_24001 (I410730,I410535,I261199);
nand I_24002 (I410399,I410518,I410730);
not I_24003 (I410761,I261196);
nor I_24004 (I410778,I410761,I410713);
DFFARX1 I_24005 (I410778,I2683,I410419,I410387,);
nor I_24006 (I410809,I410761,I261202);
and I_24007 (I410826,I410809,I261205);
or I_24008 (I410843,I410826,I261178);
DFFARX1 I_24009 (I410843,I2683,I410419,I410869,);
nor I_24010 (I410877,I410869,I410493);
nor I_24011 (I410396,I410445,I410877);
not I_24012 (I410908,I410869);
nor I_24013 (I410925,I410908,I410603);
DFFARX1 I_24014 (I410925,I2683,I410419,I410402,);
nand I_24015 (I410956,I410908,I410535);
nor I_24016 (I410390,I410761,I410956);
not I_24017 (I411014,I2690);
DFFARX1 I_24018 (I463039,I2683,I411014,I411040,);
DFFARX1 I_24019 (I411040,I2683,I411014,I411057,);
not I_24020 (I411006,I411057);
DFFARX1 I_24021 (I463051,I2683,I411014,I411088,);
not I_24022 (I411096,I463036);
nor I_24023 (I411113,I411040,I411096);
not I_24024 (I411130,I463054);
not I_24025 (I411147,I463045);
nand I_24026 (I411164,I411147,I463054);
nor I_24027 (I411181,I411096,I411164);
nor I_24028 (I411198,I411088,I411181);
DFFARX1 I_24029 (I411147,I2683,I411014,I411003,);
nor I_24030 (I411229,I463045,I463057);
nand I_24031 (I411246,I411229,I463060);
nor I_24032 (I411263,I411246,I411130);
nand I_24033 (I410988,I411263,I463036);
DFFARX1 I_24034 (I411246,I2683,I411014,I411000,);
nand I_24035 (I411308,I411130,I463045);
nor I_24036 (I411325,I411130,I463045);
nand I_24037 (I410994,I411113,I411325);
not I_24038 (I411356,I463036);
nor I_24039 (I411373,I411356,I411308);
DFFARX1 I_24040 (I411373,I2683,I411014,I410982,);
nor I_24041 (I411404,I411356,I463048);
and I_24042 (I411421,I411404,I463042);
or I_24043 (I411438,I411421,I463039);
DFFARX1 I_24044 (I411438,I2683,I411014,I411464,);
nor I_24045 (I411472,I411464,I411088);
nor I_24046 (I410991,I411040,I411472);
not I_24047 (I411503,I411464);
nor I_24048 (I411520,I411503,I411198);
DFFARX1 I_24049 (I411520,I2683,I411014,I410997,);
nand I_24050 (I411551,I411503,I411130);
nor I_24051 (I410985,I411356,I411551);
not I_24052 (I411609,I2690);
DFFARX1 I_24053 (I910868,I2683,I411609,I411635,);
DFFARX1 I_24054 (I411635,I2683,I411609,I411652,);
not I_24055 (I411601,I411652);
DFFARX1 I_24056 (I910850,I2683,I411609,I411683,);
not I_24057 (I411691,I910856);
nor I_24058 (I411708,I411635,I411691);
not I_24059 (I411725,I910871);
not I_24060 (I411742,I910862);
nand I_24061 (I411759,I411742,I910871);
nor I_24062 (I411776,I411691,I411759);
nor I_24063 (I411793,I411683,I411776);
DFFARX1 I_24064 (I411742,I2683,I411609,I411598,);
nor I_24065 (I411824,I910862,I910874);
nand I_24066 (I411841,I411824,I910853);
nor I_24067 (I411858,I411841,I411725);
nand I_24068 (I411583,I411858,I910856);
DFFARX1 I_24069 (I411841,I2683,I411609,I411595,);
nand I_24070 (I411903,I411725,I910862);
nor I_24071 (I411920,I411725,I910862);
nand I_24072 (I411589,I411708,I411920);
not I_24073 (I411951,I910859);
nor I_24074 (I411968,I411951,I411903);
DFFARX1 I_24075 (I411968,I2683,I411609,I411577,);
nor I_24076 (I411999,I411951,I910865);
and I_24077 (I412016,I411999,I910850);
or I_24078 (I412033,I412016,I910853);
DFFARX1 I_24079 (I412033,I2683,I411609,I412059,);
nor I_24080 (I412067,I412059,I411683);
nor I_24081 (I411586,I411635,I412067);
not I_24082 (I412098,I412059);
nor I_24083 (I412115,I412098,I411793);
DFFARX1 I_24084 (I412115,I2683,I411609,I411592,);
nand I_24085 (I412146,I412098,I411725);
nor I_24086 (I411580,I411951,I412146);
not I_24087 (I412204,I2690);
DFFARX1 I_24088 (I239586,I2683,I412204,I412230,);
DFFARX1 I_24089 (I412230,I2683,I412204,I412247,);
not I_24090 (I412196,I412247);
DFFARX1 I_24091 (I239574,I2683,I412204,I412278,);
not I_24092 (I412286,I239577);
nor I_24093 (I412303,I412230,I412286);
not I_24094 (I412320,I239580);
not I_24095 (I412337,I239592);
nand I_24096 (I412354,I412337,I239580);
nor I_24097 (I412371,I412286,I412354);
nor I_24098 (I412388,I412278,I412371);
DFFARX1 I_24099 (I412337,I2683,I412204,I412193,);
nor I_24100 (I412419,I239592,I239583);
nand I_24101 (I412436,I412419,I239571);
nor I_24102 (I412453,I412436,I412320);
nand I_24103 (I412178,I412453,I239577);
DFFARX1 I_24104 (I412436,I2683,I412204,I412190,);
nand I_24105 (I412498,I412320,I239592);
nor I_24106 (I412515,I412320,I239592);
nand I_24107 (I412184,I412303,I412515);
not I_24108 (I412546,I239589);
nor I_24109 (I412563,I412546,I412498);
DFFARX1 I_24110 (I412563,I2683,I412204,I412172,);
nor I_24111 (I412594,I412546,I239595);
and I_24112 (I412611,I412594,I239598);
or I_24113 (I412628,I412611,I239571);
DFFARX1 I_24114 (I412628,I2683,I412204,I412654,);
nor I_24115 (I412662,I412654,I412278);
nor I_24116 (I412181,I412230,I412662);
not I_24117 (I412693,I412654);
nor I_24118 (I412710,I412693,I412388);
DFFARX1 I_24119 (I412710,I2683,I412204,I412187,);
nand I_24120 (I412741,I412693,I412320);
nor I_24121 (I412175,I412546,I412741);
not I_24122 (I412799,I2690);
DFFARX1 I_24123 (I224303,I2683,I412799,I412825,);
DFFARX1 I_24124 (I412825,I2683,I412799,I412842,);
not I_24125 (I412791,I412842);
DFFARX1 I_24126 (I224291,I2683,I412799,I412873,);
not I_24127 (I412881,I224294);
nor I_24128 (I412898,I412825,I412881);
not I_24129 (I412915,I224297);
not I_24130 (I412932,I224309);
nand I_24131 (I412949,I412932,I224297);
nor I_24132 (I412966,I412881,I412949);
nor I_24133 (I412983,I412873,I412966);
DFFARX1 I_24134 (I412932,I2683,I412799,I412788,);
nor I_24135 (I413014,I224309,I224300);
nand I_24136 (I413031,I413014,I224288);
nor I_24137 (I413048,I413031,I412915);
nand I_24138 (I412773,I413048,I224294);
DFFARX1 I_24139 (I413031,I2683,I412799,I412785,);
nand I_24140 (I413093,I412915,I224309);
nor I_24141 (I413110,I412915,I224309);
nand I_24142 (I412779,I412898,I413110);
not I_24143 (I413141,I224306);
nor I_24144 (I413158,I413141,I413093);
DFFARX1 I_24145 (I413158,I2683,I412799,I412767,);
nor I_24146 (I413189,I413141,I224312);
and I_24147 (I413206,I413189,I224315);
or I_24148 (I413223,I413206,I224288);
DFFARX1 I_24149 (I413223,I2683,I412799,I413249,);
nor I_24150 (I413257,I413249,I412873);
nor I_24151 (I412776,I412825,I413257);
not I_24152 (I413288,I413249);
nor I_24153 (I413305,I413288,I412983);
DFFARX1 I_24154 (I413305,I2683,I412799,I412782,);
nand I_24155 (I413336,I413288,I412915);
nor I_24156 (I412770,I413141,I413336);
not I_24157 (I413394,I2690);
DFFARX1 I_24158 (I827074,I2683,I413394,I413420,);
DFFARX1 I_24159 (I413420,I2683,I413394,I413437,);
not I_24160 (I413386,I413437);
DFFARX1 I_24161 (I827077,I2683,I413394,I413468,);
not I_24162 (I413476,I827080);
nor I_24163 (I413493,I413420,I413476);
not I_24164 (I413510,I827092);
not I_24165 (I413527,I827083);
nand I_24166 (I413544,I413527,I827092);
nor I_24167 (I413561,I413476,I413544);
nor I_24168 (I413578,I413468,I413561);
DFFARX1 I_24169 (I413527,I2683,I413394,I413383,);
nor I_24170 (I413609,I827083,I827089);
nand I_24171 (I413626,I413609,I827077);
nor I_24172 (I413643,I413626,I413510);
nand I_24173 (I413368,I413643,I827080);
DFFARX1 I_24174 (I413626,I2683,I413394,I413380,);
nand I_24175 (I413688,I413510,I827083);
nor I_24176 (I413705,I413510,I827083);
nand I_24177 (I413374,I413493,I413705);
not I_24178 (I413736,I827080);
nor I_24179 (I413753,I413736,I413688);
DFFARX1 I_24180 (I413753,I2683,I413394,I413362,);
nor I_24181 (I413784,I413736,I827086);
and I_24182 (I413801,I413784,I827074);
or I_24183 (I413818,I413801,I827095);
DFFARX1 I_24184 (I413818,I2683,I413394,I413844,);
nor I_24185 (I413852,I413844,I413468);
nor I_24186 (I413371,I413420,I413852);
not I_24187 (I413883,I413844);
nor I_24188 (I413900,I413883,I413578);
DFFARX1 I_24189 (I413900,I2683,I413394,I413377,);
nand I_24190 (I413931,I413883,I413510);
nor I_24191 (I413365,I413736,I413931);
not I_24192 (I413989,I2690);
DFFARX1 I_24193 (I816976,I2683,I413989,I414015,);
DFFARX1 I_24194 (I414015,I2683,I413989,I414032,);
not I_24195 (I413981,I414032);
DFFARX1 I_24196 (I816979,I2683,I413989,I414063,);
not I_24197 (I414071,I816982);
nor I_24198 (I414088,I414015,I414071);
not I_24199 (I414105,I816994);
not I_24200 (I414122,I816985);
nand I_24201 (I414139,I414122,I816994);
nor I_24202 (I414156,I414071,I414139);
nor I_24203 (I414173,I414063,I414156);
DFFARX1 I_24204 (I414122,I2683,I413989,I413978,);
nor I_24205 (I414204,I816985,I816991);
nand I_24206 (I414221,I414204,I816979);
nor I_24207 (I414238,I414221,I414105);
nand I_24208 (I413963,I414238,I816982);
DFFARX1 I_24209 (I414221,I2683,I413989,I413975,);
nand I_24210 (I414283,I414105,I816985);
nor I_24211 (I414300,I414105,I816985);
nand I_24212 (I413969,I414088,I414300);
not I_24213 (I414331,I816982);
nor I_24214 (I414348,I414331,I414283);
DFFARX1 I_24215 (I414348,I2683,I413989,I413957,);
nor I_24216 (I414379,I414331,I816988);
and I_24217 (I414396,I414379,I816976);
or I_24218 (I414413,I414396,I816997);
DFFARX1 I_24219 (I414413,I2683,I413989,I414439,);
nor I_24220 (I414447,I414439,I414063);
nor I_24221 (I413966,I414015,I414447);
not I_24222 (I414478,I414439);
nor I_24223 (I414495,I414478,I414173);
DFFARX1 I_24224 (I414495,I2683,I413989,I413972,);
nand I_24225 (I414526,I414478,I414105);
nor I_24226 (I413960,I414331,I414526);
not I_24227 (I414584,I2690);
DFFARX1 I_24228 (I932254,I2683,I414584,I414610,);
DFFARX1 I_24229 (I414610,I2683,I414584,I414627,);
not I_24230 (I414576,I414627);
DFFARX1 I_24231 (I932236,I2683,I414584,I414658,);
not I_24232 (I414666,I932242);
nor I_24233 (I414683,I414610,I414666);
not I_24234 (I414700,I932257);
not I_24235 (I414717,I932248);
nand I_24236 (I414734,I414717,I932257);
nor I_24237 (I414751,I414666,I414734);
nor I_24238 (I414768,I414658,I414751);
DFFARX1 I_24239 (I414717,I2683,I414584,I414573,);
nor I_24240 (I414799,I932248,I932260);
nand I_24241 (I414816,I414799,I932239);
nor I_24242 (I414833,I414816,I414700);
nand I_24243 (I414558,I414833,I932242);
DFFARX1 I_24244 (I414816,I2683,I414584,I414570,);
nand I_24245 (I414878,I414700,I932248);
nor I_24246 (I414895,I414700,I932248);
nand I_24247 (I414564,I414683,I414895);
not I_24248 (I414926,I932245);
nor I_24249 (I414943,I414926,I414878);
DFFARX1 I_24250 (I414943,I2683,I414584,I414552,);
nor I_24251 (I414974,I414926,I932251);
and I_24252 (I414991,I414974,I932236);
or I_24253 (I415008,I414991,I932239);
DFFARX1 I_24254 (I415008,I2683,I414584,I415034,);
nor I_24255 (I415042,I415034,I414658);
nor I_24256 (I414561,I414610,I415042);
not I_24257 (I415073,I415034);
nor I_24258 (I415090,I415073,I414768);
DFFARX1 I_24259 (I415090,I2683,I414584,I414567,);
nand I_24260 (I415121,I415073,I414700);
nor I_24261 (I414555,I414926,I415121);
not I_24262 (I415179,I2690);
DFFARX1 I_24263 (I659684,I2683,I415179,I415205,);
DFFARX1 I_24264 (I415205,I2683,I415179,I415222,);
not I_24265 (I415171,I415222);
DFFARX1 I_24266 (I659681,I2683,I415179,I415253,);
not I_24267 (I415261,I659681);
nor I_24268 (I415278,I415205,I415261);
not I_24269 (I415295,I659678);
not I_24270 (I415312,I659693);
nand I_24271 (I415329,I415312,I659678);
nor I_24272 (I415346,I415261,I415329);
nor I_24273 (I415363,I415253,I415346);
DFFARX1 I_24274 (I415312,I2683,I415179,I415168,);
nor I_24275 (I415394,I659693,I659687);
nand I_24276 (I415411,I415394,I659675);
nor I_24277 (I415428,I415411,I415295);
nand I_24278 (I415153,I415428,I659681);
DFFARX1 I_24279 (I415411,I2683,I415179,I415165,);
nand I_24280 (I415473,I415295,I659693);
nor I_24281 (I415490,I415295,I659693);
nand I_24282 (I415159,I415278,I415490);
not I_24283 (I415521,I659696);
nor I_24284 (I415538,I415521,I415473);
DFFARX1 I_24285 (I415538,I2683,I415179,I415147,);
nor I_24286 (I415569,I415521,I659675);
and I_24287 (I415586,I415569,I659690);
or I_24288 (I415603,I415586,I659678);
DFFARX1 I_24289 (I415603,I2683,I415179,I415629,);
nor I_24290 (I415637,I415629,I415253);
nor I_24291 (I415156,I415205,I415637);
not I_24292 (I415668,I415629);
nor I_24293 (I415685,I415668,I415363);
DFFARX1 I_24294 (I415685,I2683,I415179,I415162,);
nand I_24295 (I415716,I415668,I415295);
nor I_24296 (I415150,I415521,I415716);
not I_24297 (I415774,I2690);
DFFARX1 I_24298 (I297556,I2683,I415774,I415800,);
DFFARX1 I_24299 (I415800,I2683,I415774,I415817,);
not I_24300 (I415766,I415817);
DFFARX1 I_24301 (I297544,I2683,I415774,I415848,);
not I_24302 (I415856,I297547);
nor I_24303 (I415873,I415800,I415856);
not I_24304 (I415890,I297550);
not I_24305 (I415907,I297562);
nand I_24306 (I415924,I415907,I297550);
nor I_24307 (I415941,I415856,I415924);
nor I_24308 (I415958,I415848,I415941);
DFFARX1 I_24309 (I415907,I2683,I415774,I415763,);
nor I_24310 (I415989,I297562,I297553);
nand I_24311 (I416006,I415989,I297541);
nor I_24312 (I416023,I416006,I415890);
nand I_24313 (I415748,I416023,I297547);
DFFARX1 I_24314 (I416006,I2683,I415774,I415760,);
nand I_24315 (I416068,I415890,I297562);
nor I_24316 (I416085,I415890,I297562);
nand I_24317 (I415754,I415873,I416085);
not I_24318 (I416116,I297559);
nor I_24319 (I416133,I416116,I416068);
DFFARX1 I_24320 (I416133,I2683,I415774,I415742,);
nor I_24321 (I416164,I416116,I297565);
and I_24322 (I416181,I416164,I297568);
or I_24323 (I416198,I416181,I297541);
DFFARX1 I_24324 (I416198,I2683,I415774,I416224,);
nor I_24325 (I416232,I416224,I415848);
nor I_24326 (I415751,I415800,I416232);
not I_24327 (I416263,I416224);
nor I_24328 (I416280,I416263,I415958);
DFFARX1 I_24329 (I416280,I2683,I415774,I415757,);
nand I_24330 (I416311,I416263,I415890);
nor I_24331 (I415745,I416116,I416311);
not I_24332 (I416369,I2690);
DFFARX1 I_24333 (I556681,I2683,I416369,I416395,);
DFFARX1 I_24334 (I416395,I2683,I416369,I416412,);
not I_24335 (I416361,I416412);
DFFARX1 I_24336 (I556675,I2683,I416369,I416443,);
not I_24337 (I416451,I556672);
nor I_24338 (I416468,I416395,I416451);
not I_24339 (I416485,I556684);
not I_24340 (I416502,I556687);
nand I_24341 (I416519,I416502,I556684);
nor I_24342 (I416536,I416451,I416519);
nor I_24343 (I416553,I416443,I416536);
DFFARX1 I_24344 (I416502,I2683,I416369,I416358,);
nor I_24345 (I416584,I556687,I556696);
nand I_24346 (I416601,I416584,I556690);
nor I_24347 (I416618,I416601,I416485);
nand I_24348 (I416343,I416618,I556672);
DFFARX1 I_24349 (I416601,I2683,I416369,I416355,);
nand I_24350 (I416663,I416485,I556687);
nor I_24351 (I416680,I416485,I556687);
nand I_24352 (I416349,I416468,I416680);
not I_24353 (I416711,I556678);
nor I_24354 (I416728,I416711,I416663);
DFFARX1 I_24355 (I416728,I2683,I416369,I416337,);
nor I_24356 (I416759,I416711,I556693);
and I_24357 (I416776,I416759,I556672);
or I_24358 (I416793,I416776,I556675);
DFFARX1 I_24359 (I416793,I2683,I416369,I416819,);
nor I_24360 (I416827,I416819,I416443);
nor I_24361 (I416346,I416395,I416827);
not I_24362 (I416858,I416819);
nor I_24363 (I416875,I416858,I416553);
DFFARX1 I_24364 (I416875,I2683,I416369,I416352,);
nand I_24365 (I416906,I416858,I416485);
nor I_24366 (I416340,I416711,I416906);
not I_24367 (I416964,I2690);
DFFARX1 I_24368 (I376914,I2683,I416964,I416990,);
DFFARX1 I_24369 (I416990,I2683,I416964,I417007,);
not I_24370 (I416956,I417007);
DFFARX1 I_24371 (I376938,I2683,I416964,I417038,);
not I_24372 (I417046,I376917);
nor I_24373 (I417063,I416990,I417046);
not I_24374 (I417080,I376923);
not I_24375 (I417097,I376929);
nand I_24376 (I417114,I417097,I376923);
nor I_24377 (I417131,I417046,I417114);
nor I_24378 (I417148,I417038,I417131);
DFFARX1 I_24379 (I417097,I2683,I416964,I416953,);
nor I_24380 (I417179,I376929,I376941);
nand I_24381 (I417196,I417179,I376935);
nor I_24382 (I417213,I417196,I417080);
nand I_24383 (I416938,I417213,I376917);
DFFARX1 I_24384 (I417196,I2683,I416964,I416950,);
nand I_24385 (I417258,I417080,I376929);
nor I_24386 (I417275,I417080,I376929);
nand I_24387 (I416944,I417063,I417275);
not I_24388 (I417306,I376920);
nor I_24389 (I417323,I417306,I417258);
DFFARX1 I_24390 (I417323,I2683,I416964,I416932,);
nor I_24391 (I417354,I417306,I376914);
and I_24392 (I417371,I417354,I376932);
or I_24393 (I417388,I417371,I376926);
DFFARX1 I_24394 (I417388,I2683,I416964,I417414,);
nor I_24395 (I417422,I417414,I417038);
nor I_24396 (I416941,I416990,I417422);
not I_24397 (I417453,I417414);
nor I_24398 (I417470,I417453,I417148);
DFFARX1 I_24399 (I417470,I2683,I416964,I416947,);
nand I_24400 (I417501,I417453,I417080);
nor I_24401 (I416935,I417306,I417501);
not I_24402 (I417559,I2690);
DFFARX1 I_24403 (I828792,I2683,I417559,I417585,);
DFFARX1 I_24404 (I417585,I2683,I417559,I417602,);
not I_24405 (I417551,I417602);
DFFARX1 I_24406 (I828774,I2683,I417559,I417633,);
not I_24407 (I417641,I828780);
nor I_24408 (I417658,I417585,I417641);
not I_24409 (I417675,I828795);
not I_24410 (I417692,I828786);
nand I_24411 (I417709,I417692,I828795);
nor I_24412 (I417726,I417641,I417709);
nor I_24413 (I417743,I417633,I417726);
DFFARX1 I_24414 (I417692,I2683,I417559,I417548,);
nor I_24415 (I417774,I828786,I828798);
nand I_24416 (I417791,I417774,I828777);
nor I_24417 (I417808,I417791,I417675);
nand I_24418 (I417533,I417808,I828780);
DFFARX1 I_24419 (I417791,I2683,I417559,I417545,);
nand I_24420 (I417853,I417675,I828786);
nor I_24421 (I417870,I417675,I828786);
nand I_24422 (I417539,I417658,I417870);
not I_24423 (I417901,I828783);
nor I_24424 (I417918,I417901,I417853);
DFFARX1 I_24425 (I417918,I2683,I417559,I417527,);
nor I_24426 (I417949,I417901,I828789);
and I_24427 (I417966,I417949,I828774);
or I_24428 (I417983,I417966,I828777);
DFFARX1 I_24429 (I417983,I2683,I417559,I418009,);
nor I_24430 (I418017,I418009,I417633);
nor I_24431 (I417536,I417585,I418017);
not I_24432 (I418048,I418009);
nor I_24433 (I418065,I418048,I417743);
DFFARX1 I_24434 (I418065,I2683,I417559,I417542,);
nand I_24435 (I418096,I418048,I417675);
nor I_24436 (I417530,I417901,I418096);
not I_24437 (I418154,I2690);
DFFARX1 I_24438 (I125960,I2683,I418154,I418180,);
DFFARX1 I_24439 (I418180,I2683,I418154,I418197,);
not I_24440 (I418146,I418197);
DFFARX1 I_24441 (I125984,I2683,I418154,I418228,);
not I_24442 (I418236,I125978);
nor I_24443 (I418253,I418180,I418236);
not I_24444 (I418270,I125972);
not I_24445 (I418287,I125969);
nand I_24446 (I418304,I418287,I125972);
nor I_24447 (I418321,I418236,I418304);
nor I_24448 (I418338,I418228,I418321);
DFFARX1 I_24449 (I418287,I2683,I418154,I418143,);
nor I_24450 (I418369,I125969,I125963);
nand I_24451 (I418386,I418369,I125981);
nor I_24452 (I418403,I418386,I418270);
nand I_24453 (I418128,I418403,I125978);
DFFARX1 I_24454 (I418386,I2683,I418154,I418140,);
nand I_24455 (I418448,I418270,I125969);
nor I_24456 (I418465,I418270,I125969);
nand I_24457 (I418134,I418253,I418465);
not I_24458 (I418496,I125975);
nor I_24459 (I418513,I418496,I418448);
DFFARX1 I_24460 (I418513,I2683,I418154,I418122,);
nor I_24461 (I418544,I418496,I125960);
and I_24462 (I418561,I418544,I125966);
or I_24463 (I418578,I418561,I125963);
DFFARX1 I_24464 (I418578,I2683,I418154,I418604,);
nor I_24465 (I418612,I418604,I418228);
nor I_24466 (I418131,I418180,I418612);
not I_24467 (I418643,I418604);
nor I_24468 (I418660,I418643,I418338);
DFFARX1 I_24469 (I418660,I2683,I418154,I418137,);
nand I_24470 (I418691,I418643,I418270);
nor I_24471 (I418125,I418496,I418691);
not I_24472 (I418749,I2690);
DFFARX1 I_24473 (I748430,I2683,I418749,I418775,);
DFFARX1 I_24474 (I418775,I2683,I418749,I418792,);
not I_24475 (I418741,I418792);
DFFARX1 I_24476 (I748418,I2683,I418749,I418823,);
not I_24477 (I418831,I748415);
nor I_24478 (I418848,I418775,I418831);
not I_24479 (I418865,I748427);
not I_24480 (I418882,I748424);
nand I_24481 (I418899,I418882,I748427);
nor I_24482 (I418916,I418831,I418899);
nor I_24483 (I418933,I418823,I418916);
DFFARX1 I_24484 (I418882,I2683,I418749,I418738,);
nor I_24485 (I418964,I748424,I748433);
nand I_24486 (I418981,I418964,I748436);
nor I_24487 (I418998,I418981,I418865);
nand I_24488 (I418723,I418998,I748415);
DFFARX1 I_24489 (I418981,I2683,I418749,I418735,);
nand I_24490 (I419043,I418865,I748424);
nor I_24491 (I419060,I418865,I748424);
nand I_24492 (I418729,I418848,I419060);
not I_24493 (I419091,I748439);
nor I_24494 (I419108,I419091,I419043);
DFFARX1 I_24495 (I419108,I2683,I418749,I418717,);
nor I_24496 (I419139,I419091,I748442);
and I_24497 (I419156,I419139,I748421);
or I_24498 (I419173,I419156,I748415);
DFFARX1 I_24499 (I419173,I2683,I418749,I419199,);
nor I_24500 (I419207,I419199,I418823);
nor I_24501 (I418726,I418775,I419207);
not I_24502 (I419238,I419199);
nor I_24503 (I419255,I419238,I418933);
DFFARX1 I_24504 (I419255,I2683,I418749,I418732,);
nand I_24505 (I419286,I419238,I418865);
nor I_24506 (I418720,I419091,I419286);
not I_24507 (I419344,I2690);
DFFARX1 I_24508 (I939190,I2683,I419344,I419370,);
DFFARX1 I_24509 (I419370,I2683,I419344,I419387,);
not I_24510 (I419336,I419387);
DFFARX1 I_24511 (I939172,I2683,I419344,I419418,);
not I_24512 (I419426,I939178);
nor I_24513 (I419443,I419370,I419426);
not I_24514 (I419460,I939193);
not I_24515 (I419477,I939184);
nand I_24516 (I419494,I419477,I939193);
nor I_24517 (I419511,I419426,I419494);
nor I_24518 (I419528,I419418,I419511);
DFFARX1 I_24519 (I419477,I2683,I419344,I419333,);
nor I_24520 (I419559,I939184,I939196);
nand I_24521 (I419576,I419559,I939175);
nor I_24522 (I419593,I419576,I419460);
nand I_24523 (I419318,I419593,I939178);
DFFARX1 I_24524 (I419576,I2683,I419344,I419330,);
nand I_24525 (I419638,I419460,I939184);
nor I_24526 (I419655,I419460,I939184);
nand I_24527 (I419324,I419443,I419655);
not I_24528 (I419686,I939181);
nor I_24529 (I419703,I419686,I419638);
DFFARX1 I_24530 (I419703,I2683,I419344,I419312,);
nor I_24531 (I419734,I419686,I939187);
and I_24532 (I419751,I419734,I939172);
or I_24533 (I419768,I419751,I939175);
DFFARX1 I_24534 (I419768,I2683,I419344,I419794,);
nor I_24535 (I419802,I419794,I419418);
nor I_24536 (I419321,I419370,I419802);
not I_24537 (I419833,I419794);
nor I_24538 (I419850,I419833,I419528);
DFFARX1 I_24539 (I419850,I2683,I419344,I419327,);
nand I_24540 (I419881,I419833,I419460);
nor I_24541 (I419315,I419686,I419881);
not I_24542 (I419939,I2690);
DFFARX1 I_24543 (I866940,I2683,I419939,I419965,);
DFFARX1 I_24544 (I419965,I2683,I419939,I419982,);
not I_24545 (I419931,I419982);
DFFARX1 I_24546 (I866922,I2683,I419939,I420013,);
not I_24547 (I420021,I866928);
nor I_24548 (I420038,I419965,I420021);
not I_24549 (I420055,I866943);
not I_24550 (I420072,I866934);
nand I_24551 (I420089,I420072,I866943);
nor I_24552 (I420106,I420021,I420089);
nor I_24553 (I420123,I420013,I420106);
DFFARX1 I_24554 (I420072,I2683,I419939,I419928,);
nor I_24555 (I420154,I866934,I866946);
nand I_24556 (I420171,I420154,I866925);
nor I_24557 (I420188,I420171,I420055);
nand I_24558 (I419913,I420188,I866928);
DFFARX1 I_24559 (I420171,I2683,I419939,I419925,);
nand I_24560 (I420233,I420055,I866934);
nor I_24561 (I420250,I420055,I866934);
nand I_24562 (I419919,I420038,I420250);
not I_24563 (I420281,I866931);
nor I_24564 (I420298,I420281,I420233);
DFFARX1 I_24565 (I420298,I2683,I419939,I419907,);
nor I_24566 (I420329,I420281,I866937);
and I_24567 (I420346,I420329,I866922);
or I_24568 (I420363,I420346,I866925);
DFFARX1 I_24569 (I420363,I2683,I419939,I420389,);
nor I_24570 (I420397,I420389,I420013);
nor I_24571 (I419916,I419965,I420397);
not I_24572 (I420428,I420389);
nor I_24573 (I420445,I420428,I420123);
DFFARX1 I_24574 (I420445,I2683,I419939,I419922,);
nand I_24575 (I420476,I420428,I420055);
nor I_24576 (I419910,I420281,I420476);
not I_24577 (I420534,I2690);
DFFARX1 I_24578 (I174155,I2683,I420534,I420560,);
DFFARX1 I_24579 (I420560,I2683,I420534,I420577,);
not I_24580 (I420526,I420577);
DFFARX1 I_24581 (I174179,I2683,I420534,I420608,);
not I_24582 (I420616,I174173);
nor I_24583 (I420633,I420560,I420616);
not I_24584 (I420650,I174167);
not I_24585 (I420667,I174164);
nand I_24586 (I420684,I420667,I174167);
nor I_24587 (I420701,I420616,I420684);
nor I_24588 (I420718,I420608,I420701);
DFFARX1 I_24589 (I420667,I2683,I420534,I420523,);
nor I_24590 (I420749,I174164,I174158);
nand I_24591 (I420766,I420749,I174176);
nor I_24592 (I420783,I420766,I420650);
nand I_24593 (I420508,I420783,I174173);
DFFARX1 I_24594 (I420766,I2683,I420534,I420520,);
nand I_24595 (I420828,I420650,I174164);
nor I_24596 (I420845,I420650,I174164);
nand I_24597 (I420514,I420633,I420845);
not I_24598 (I420876,I174170);
nor I_24599 (I420893,I420876,I420828);
DFFARX1 I_24600 (I420893,I2683,I420534,I420502,);
nor I_24601 (I420924,I420876,I174155);
and I_24602 (I420941,I420924,I174161);
or I_24603 (I420958,I420941,I174158);
DFFARX1 I_24604 (I420958,I2683,I420534,I420984,);
nor I_24605 (I420992,I420984,I420608);
nor I_24606 (I420511,I420560,I420992);
not I_24607 (I421023,I420984);
nor I_24608 (I421040,I421023,I420718);
DFFARX1 I_24609 (I421040,I2683,I420534,I420517,);
nand I_24610 (I421071,I421023,I420650);
nor I_24611 (I420505,I420876,I421071);
not I_24612 (I421129,I2690);
DFFARX1 I_24613 (I1019795,I2683,I421129,I421155,);
DFFARX1 I_24614 (I421155,I2683,I421129,I421172,);
not I_24615 (I421121,I421172);
DFFARX1 I_24616 (I1019801,I2683,I421129,I421203,);
not I_24617 (I421211,I1019789);
nor I_24618 (I421228,I421155,I421211);
not I_24619 (I421245,I1019792);
not I_24620 (I421262,I1019798);
nand I_24621 (I421279,I421262,I1019792);
nor I_24622 (I421296,I421211,I421279);
nor I_24623 (I421313,I421203,I421296);
DFFARX1 I_24624 (I421262,I2683,I421129,I421118,);
nor I_24625 (I421344,I1019798,I1019789);
nand I_24626 (I421361,I421344,I1019807);
nor I_24627 (I421378,I421361,I421245);
nand I_24628 (I421103,I421378,I1019789);
DFFARX1 I_24629 (I421361,I2683,I421129,I421115,);
nand I_24630 (I421423,I421245,I1019798);
nor I_24631 (I421440,I421245,I1019798);
nand I_24632 (I421109,I421228,I421440);
not I_24633 (I421471,I1019786);
nor I_24634 (I421488,I421471,I421423);
DFFARX1 I_24635 (I421488,I2683,I421129,I421097,);
nor I_24636 (I421519,I421471,I1019810);
and I_24637 (I421536,I421519,I1019786);
or I_24638 (I421553,I421536,I1019804);
DFFARX1 I_24639 (I421553,I2683,I421129,I421579,);
nor I_24640 (I421587,I421579,I421203);
nor I_24641 (I421106,I421155,I421587);
not I_24642 (I421618,I421579);
nor I_24643 (I421635,I421618,I421313);
DFFARX1 I_24644 (I421635,I2683,I421129,I421112,);
nand I_24645 (I421666,I421618,I421245);
nor I_24646 (I421100,I421471,I421666);
not I_24647 (I421724,I2690);
DFFARX1 I_24648 (I996097,I2683,I421724,I421750,);
DFFARX1 I_24649 (I421750,I2683,I421724,I421767,);
not I_24650 (I421716,I421767);
DFFARX1 I_24651 (I996103,I2683,I421724,I421798,);
not I_24652 (I421806,I996091);
nor I_24653 (I421823,I421750,I421806);
not I_24654 (I421840,I996094);
not I_24655 (I421857,I996100);
nand I_24656 (I421874,I421857,I996094);
nor I_24657 (I421891,I421806,I421874);
nor I_24658 (I421908,I421798,I421891);
DFFARX1 I_24659 (I421857,I2683,I421724,I421713,);
nor I_24660 (I421939,I996100,I996091);
nand I_24661 (I421956,I421939,I996109);
nor I_24662 (I421973,I421956,I421840);
nand I_24663 (I421698,I421973,I996091);
DFFARX1 I_24664 (I421956,I2683,I421724,I421710,);
nand I_24665 (I422018,I421840,I996100);
nor I_24666 (I422035,I421840,I996100);
nand I_24667 (I421704,I421823,I422035);
not I_24668 (I422066,I996088);
nor I_24669 (I422083,I422066,I422018);
DFFARX1 I_24670 (I422083,I2683,I421724,I421692,);
nor I_24671 (I422114,I422066,I996112);
and I_24672 (I422131,I422114,I996088);
or I_24673 (I422148,I422131,I996106);
DFFARX1 I_24674 (I422148,I2683,I421724,I422174,);
nor I_24675 (I422182,I422174,I421798);
nor I_24676 (I421701,I421750,I422182);
not I_24677 (I422213,I422174);
nor I_24678 (I422230,I422213,I421908);
DFFARX1 I_24679 (I422230,I2683,I421724,I421707,);
nand I_24680 (I422261,I422213,I421840);
nor I_24681 (I421695,I422066,I422261);
not I_24682 (I422319,I2690);
DFFARX1 I_24683 (I442231,I2683,I422319,I422345,);
DFFARX1 I_24684 (I422345,I2683,I422319,I422362,);
not I_24685 (I422311,I422362);
DFFARX1 I_24686 (I442243,I2683,I422319,I422393,);
not I_24687 (I422401,I442228);
nor I_24688 (I422418,I422345,I422401);
not I_24689 (I422435,I442246);
not I_24690 (I422452,I442237);
nand I_24691 (I422469,I422452,I442246);
nor I_24692 (I422486,I422401,I422469);
nor I_24693 (I422503,I422393,I422486);
DFFARX1 I_24694 (I422452,I2683,I422319,I422308,);
nor I_24695 (I422534,I442237,I442249);
nand I_24696 (I422551,I422534,I442252);
nor I_24697 (I422568,I422551,I422435);
nand I_24698 (I422293,I422568,I442228);
DFFARX1 I_24699 (I422551,I2683,I422319,I422305,);
nand I_24700 (I422613,I422435,I442237);
nor I_24701 (I422630,I422435,I442237);
nand I_24702 (I422299,I422418,I422630);
not I_24703 (I422661,I442228);
nor I_24704 (I422678,I422661,I422613);
DFFARX1 I_24705 (I422678,I2683,I422319,I422287,);
nor I_24706 (I422709,I422661,I442240);
and I_24707 (I422726,I422709,I442234);
or I_24708 (I422743,I422726,I442231);
DFFARX1 I_24709 (I422743,I2683,I422319,I422769,);
nor I_24710 (I422777,I422769,I422393);
nor I_24711 (I422296,I422345,I422777);
not I_24712 (I422808,I422769);
nor I_24713 (I422825,I422808,I422503);
DFFARX1 I_24714 (I422825,I2683,I422319,I422302,);
nand I_24715 (I422856,I422808,I422435);
nor I_24716 (I422290,I422661,I422856);
not I_24717 (I422914,I2690);
DFFARX1 I_24718 (I122390,I2683,I422914,I422940,);
DFFARX1 I_24719 (I422940,I2683,I422914,I422957,);
not I_24720 (I422906,I422957);
DFFARX1 I_24721 (I122414,I2683,I422914,I422988,);
not I_24722 (I422996,I122408);
nor I_24723 (I423013,I422940,I422996);
not I_24724 (I423030,I122402);
not I_24725 (I423047,I122399);
nand I_24726 (I423064,I423047,I122402);
nor I_24727 (I423081,I422996,I423064);
nor I_24728 (I423098,I422988,I423081);
DFFARX1 I_24729 (I423047,I2683,I422914,I422903,);
nor I_24730 (I423129,I122399,I122393);
nand I_24731 (I423146,I423129,I122411);
nor I_24732 (I423163,I423146,I423030);
nand I_24733 (I422888,I423163,I122408);
DFFARX1 I_24734 (I423146,I2683,I422914,I422900,);
nand I_24735 (I423208,I423030,I122399);
nor I_24736 (I423225,I423030,I122399);
nand I_24737 (I422894,I423013,I423225);
not I_24738 (I423256,I122405);
nor I_24739 (I423273,I423256,I423208);
DFFARX1 I_24740 (I423273,I2683,I422914,I422882,);
nor I_24741 (I423304,I423256,I122390);
and I_24742 (I423321,I423304,I122396);
or I_24743 (I423338,I423321,I122393);
DFFARX1 I_24744 (I423338,I2683,I422914,I423364,);
nor I_24745 (I423372,I423364,I422988);
nor I_24746 (I422891,I422940,I423372);
not I_24747 (I423403,I423364);
nor I_24748 (I423420,I423403,I423098);
DFFARX1 I_24749 (I423420,I2683,I422914,I422897,);
nand I_24750 (I423451,I423403,I423030);
nor I_24751 (I422885,I423256,I423451);
not I_24752 (I423509,I2690);
DFFARX1 I_24753 (I13726,I2683,I423509,I423535,);
DFFARX1 I_24754 (I423535,I2683,I423509,I423552,);
not I_24755 (I423501,I423552);
DFFARX1 I_24756 (I13726,I2683,I423509,I423583,);
not I_24757 (I423591,I13741);
nor I_24758 (I423608,I423535,I423591);
not I_24759 (I423625,I13744);
not I_24760 (I423642,I13735);
nand I_24761 (I423659,I423642,I13744);
nor I_24762 (I423676,I423591,I423659);
nor I_24763 (I423693,I423583,I423676);
DFFARX1 I_24764 (I423642,I2683,I423509,I423498,);
nor I_24765 (I423724,I13735,I13747);
nand I_24766 (I423741,I423724,I13729);
nor I_24767 (I423758,I423741,I423625);
nand I_24768 (I423483,I423758,I13741);
DFFARX1 I_24769 (I423741,I2683,I423509,I423495,);
nand I_24770 (I423803,I423625,I13735);
nor I_24771 (I423820,I423625,I13735);
nand I_24772 (I423489,I423608,I423820);
not I_24773 (I423851,I13729);
nor I_24774 (I423868,I423851,I423803);
DFFARX1 I_24775 (I423868,I2683,I423509,I423477,);
nor I_24776 (I423899,I423851,I13738);
and I_24777 (I423916,I423899,I13732);
or I_24778 (I423933,I423916,I13750);
DFFARX1 I_24779 (I423933,I2683,I423509,I423959,);
nor I_24780 (I423967,I423959,I423583);
nor I_24781 (I423486,I423535,I423967);
not I_24782 (I423998,I423959);
nor I_24783 (I424015,I423998,I423693);
DFFARX1 I_24784 (I424015,I2683,I423509,I423492,);
nand I_24785 (I424046,I423998,I423625);
nor I_24786 (I423480,I423851,I424046);
not I_24787 (I424104,I2690);
DFFARX1 I_24788 (I534139,I2683,I424104,I424130,);
DFFARX1 I_24789 (I424130,I2683,I424104,I424147,);
not I_24790 (I424096,I424147);
DFFARX1 I_24791 (I534133,I2683,I424104,I424178,);
not I_24792 (I424186,I534130);
nor I_24793 (I424203,I424130,I424186);
not I_24794 (I424220,I534142);
not I_24795 (I424237,I534145);
nand I_24796 (I424254,I424237,I534142);
nor I_24797 (I424271,I424186,I424254);
nor I_24798 (I424288,I424178,I424271);
DFFARX1 I_24799 (I424237,I2683,I424104,I424093,);
nor I_24800 (I424319,I534145,I534154);
nand I_24801 (I424336,I424319,I534148);
nor I_24802 (I424353,I424336,I424220);
nand I_24803 (I424078,I424353,I534130);
DFFARX1 I_24804 (I424336,I2683,I424104,I424090,);
nand I_24805 (I424398,I424220,I534145);
nor I_24806 (I424415,I424220,I534145);
nand I_24807 (I424084,I424203,I424415);
not I_24808 (I424446,I534136);
nor I_24809 (I424463,I424446,I424398);
DFFARX1 I_24810 (I424463,I2683,I424104,I424072,);
nor I_24811 (I424494,I424446,I534151);
and I_24812 (I424511,I424494,I534130);
or I_24813 (I424528,I424511,I534133);
DFFARX1 I_24814 (I424528,I2683,I424104,I424554,);
nor I_24815 (I424562,I424554,I424178);
nor I_24816 (I424081,I424130,I424562);
not I_24817 (I424593,I424554);
nor I_24818 (I424610,I424593,I424288);
DFFARX1 I_24819 (I424610,I2683,I424104,I424087,);
nand I_24820 (I424641,I424593,I424220);
nor I_24821 (I424075,I424446,I424641);
not I_24822 (I424699,I2690);
DFFARX1 I_24823 (I42184,I2683,I424699,I424725,);
DFFARX1 I_24824 (I424725,I2683,I424699,I424742,);
not I_24825 (I424691,I424742);
DFFARX1 I_24826 (I42184,I2683,I424699,I424773,);
not I_24827 (I424781,I42199);
nor I_24828 (I424798,I424725,I424781);
not I_24829 (I424815,I42202);
not I_24830 (I424832,I42193);
nand I_24831 (I424849,I424832,I42202);
nor I_24832 (I424866,I424781,I424849);
nor I_24833 (I424883,I424773,I424866);
DFFARX1 I_24834 (I424832,I2683,I424699,I424688,);
nor I_24835 (I424914,I42193,I42205);
nand I_24836 (I424931,I424914,I42187);
nor I_24837 (I424948,I424931,I424815);
nand I_24838 (I424673,I424948,I42199);
DFFARX1 I_24839 (I424931,I2683,I424699,I424685,);
nand I_24840 (I424993,I424815,I42193);
nor I_24841 (I425010,I424815,I42193);
nand I_24842 (I424679,I424798,I425010);
not I_24843 (I425041,I42187);
nor I_24844 (I425058,I425041,I424993);
DFFARX1 I_24845 (I425058,I2683,I424699,I424667,);
nor I_24846 (I425089,I425041,I42196);
and I_24847 (I425106,I425089,I42190);
or I_24848 (I425123,I425106,I42208);
DFFARX1 I_24849 (I425123,I2683,I424699,I425149,);
nor I_24850 (I425157,I425149,I424773);
nor I_24851 (I424676,I424725,I425157);
not I_24852 (I425188,I425149);
nor I_24853 (I425205,I425188,I424883);
DFFARX1 I_24854 (I425205,I2683,I424699,I424682,);
nand I_24855 (I425236,I425188,I424815);
nor I_24856 (I424670,I425041,I425236);
not I_24857 (I425294,I2690);
DFFARX1 I_24858 (I250653,I2683,I425294,I425320,);
DFFARX1 I_24859 (I425320,I2683,I425294,I425337,);
not I_24860 (I425286,I425337);
DFFARX1 I_24861 (I250641,I2683,I425294,I425368,);
not I_24862 (I425376,I250644);
nor I_24863 (I425393,I425320,I425376);
not I_24864 (I425410,I250647);
not I_24865 (I425427,I250659);
nand I_24866 (I425444,I425427,I250647);
nor I_24867 (I425461,I425376,I425444);
nor I_24868 (I425478,I425368,I425461);
DFFARX1 I_24869 (I425427,I2683,I425294,I425283,);
nor I_24870 (I425509,I250659,I250650);
nand I_24871 (I425526,I425509,I250638);
nor I_24872 (I425543,I425526,I425410);
nand I_24873 (I425268,I425543,I250644);
DFFARX1 I_24874 (I425526,I2683,I425294,I425280,);
nand I_24875 (I425588,I425410,I250659);
nor I_24876 (I425605,I425410,I250659);
nand I_24877 (I425274,I425393,I425605);
not I_24878 (I425636,I250656);
nor I_24879 (I425653,I425636,I425588);
DFFARX1 I_24880 (I425653,I2683,I425294,I425262,);
nor I_24881 (I425684,I425636,I250662);
and I_24882 (I425701,I425684,I250665);
or I_24883 (I425718,I425701,I250638);
DFFARX1 I_24884 (I425718,I2683,I425294,I425744,);
nor I_24885 (I425752,I425744,I425368);
nor I_24886 (I425271,I425320,I425752);
not I_24887 (I425783,I425744);
nor I_24888 (I425800,I425783,I425478);
DFFARX1 I_24889 (I425800,I2683,I425294,I425277,);
nand I_24890 (I425831,I425783,I425410);
nor I_24891 (I425265,I425636,I425831);
not I_24892 (I425889,I2690);
DFFARX1 I_24893 (I762642,I2683,I425889,I425915,);
DFFARX1 I_24894 (I425915,I2683,I425889,I425932,);
not I_24895 (I425881,I425932);
DFFARX1 I_24896 (I762630,I2683,I425889,I425963,);
not I_24897 (I425971,I762627);
nor I_24898 (I425988,I425915,I425971);
not I_24899 (I426005,I762639);
not I_24900 (I426022,I762636);
nand I_24901 (I426039,I426022,I762639);
nor I_24902 (I426056,I425971,I426039);
nor I_24903 (I426073,I425963,I426056);
DFFARX1 I_24904 (I426022,I2683,I425889,I425878,);
nor I_24905 (I426104,I762636,I762645);
nand I_24906 (I426121,I426104,I762648);
nor I_24907 (I426138,I426121,I426005);
nand I_24908 (I425863,I426138,I762627);
DFFARX1 I_24909 (I426121,I2683,I425889,I425875,);
nand I_24910 (I426183,I426005,I762636);
nor I_24911 (I426200,I426005,I762636);
nand I_24912 (I425869,I425988,I426200);
not I_24913 (I426231,I762651);
nor I_24914 (I426248,I426231,I426183);
DFFARX1 I_24915 (I426248,I2683,I425889,I425857,);
nor I_24916 (I426279,I426231,I762654);
and I_24917 (I426296,I426279,I762633);
or I_24918 (I426313,I426296,I762627);
DFFARX1 I_24919 (I426313,I2683,I425889,I426339,);
nor I_24920 (I426347,I426339,I425963);
nor I_24921 (I425866,I425915,I426347);
not I_24922 (I426378,I426339);
nor I_24923 (I426395,I426378,I426073);
DFFARX1 I_24924 (I426395,I2683,I425889,I425872,);
nand I_24925 (I426426,I426378,I426005);
nor I_24926 (I425860,I426231,I426426);
not I_24927 (I426484,I2690);
DFFARX1 I_24928 (I53787,I2683,I426484,I426510,);
DFFARX1 I_24929 (I426510,I2683,I426484,I426527,);
not I_24930 (I426476,I426527);
DFFARX1 I_24931 (I53799,I2683,I426484,I426558,);
not I_24932 (I426566,I53790);
nor I_24933 (I426583,I426510,I426566);
not I_24934 (I426600,I53781);
not I_24935 (I426617,I53778);
nand I_24936 (I426634,I426617,I53781);
nor I_24937 (I426651,I426566,I426634);
nor I_24938 (I426668,I426558,I426651);
DFFARX1 I_24939 (I426617,I2683,I426484,I426473,);
nor I_24940 (I426699,I53778,I53778);
nand I_24941 (I426716,I426699,I53796);
nor I_24942 (I426733,I426716,I426600);
nand I_24943 (I426458,I426733,I53790);
DFFARX1 I_24944 (I426716,I2683,I426484,I426470,);
nand I_24945 (I426778,I426600,I53778);
nor I_24946 (I426795,I426600,I53778);
nand I_24947 (I426464,I426583,I426795);
not I_24948 (I426826,I53802);
nor I_24949 (I426843,I426826,I426778);
DFFARX1 I_24950 (I426843,I2683,I426484,I426452,);
nor I_24951 (I426874,I426826,I53781);
and I_24952 (I426891,I426874,I53784);
or I_24953 (I426908,I426891,I53793);
DFFARX1 I_24954 (I426908,I2683,I426484,I426934,);
nor I_24955 (I426942,I426934,I426558);
nor I_24956 (I426461,I426510,I426942);
not I_24957 (I426973,I426934);
nor I_24958 (I426990,I426973,I426668);
DFFARX1 I_24959 (I426990,I2683,I426484,I426467,);
nand I_24960 (I427021,I426973,I426600);
nor I_24961 (I426455,I426826,I427021);
not I_24962 (I427079,I2690);
DFFARX1 I_24963 (I707732,I2683,I427079,I427105,);
DFFARX1 I_24964 (I427105,I2683,I427079,I427122,);
not I_24965 (I427071,I427122);
DFFARX1 I_24966 (I707720,I2683,I427079,I427153,);
not I_24967 (I427161,I707717);
nor I_24968 (I427178,I427105,I427161);
not I_24969 (I427195,I707729);
not I_24970 (I427212,I707726);
nand I_24971 (I427229,I427212,I707729);
nor I_24972 (I427246,I427161,I427229);
nor I_24973 (I427263,I427153,I427246);
DFFARX1 I_24974 (I427212,I2683,I427079,I427068,);
nor I_24975 (I427294,I707726,I707735);
nand I_24976 (I427311,I427294,I707738);
nor I_24977 (I427328,I427311,I427195);
nand I_24978 (I427053,I427328,I707717);
DFFARX1 I_24979 (I427311,I2683,I427079,I427065,);
nand I_24980 (I427373,I427195,I707726);
nor I_24981 (I427390,I427195,I707726);
nand I_24982 (I427059,I427178,I427390);
not I_24983 (I427421,I707741);
nor I_24984 (I427438,I427421,I427373);
DFFARX1 I_24985 (I427438,I2683,I427079,I427047,);
nor I_24986 (I427469,I427421,I707744);
and I_24987 (I427486,I427469,I707723);
or I_24988 (I427503,I427486,I707717);
DFFARX1 I_24989 (I427503,I2683,I427079,I427529,);
nor I_24990 (I427537,I427529,I427153);
nor I_24991 (I427056,I427105,I427537);
not I_24992 (I427568,I427529);
nor I_24993 (I427585,I427568,I427263);
DFFARX1 I_24994 (I427585,I2683,I427079,I427062,);
nand I_24995 (I427616,I427568,I427195);
nor I_24996 (I427050,I427421,I427616);
not I_24997 (I427674,I2690);
DFFARX1 I_24998 (I6867,I2683,I427674,I427700,);
DFFARX1 I_24999 (I427700,I2683,I427674,I427717,);
not I_25000 (I427666,I427717);
DFFARX1 I_25001 (I6858,I2683,I427674,I427748,);
not I_25002 (I427756,I6861);
nor I_25003 (I427773,I427700,I427756);
not I_25004 (I427790,I6873);
not I_25005 (I427807,I6858);
nand I_25006 (I427824,I427807,I6873);
nor I_25007 (I427841,I427756,I427824);
nor I_25008 (I427858,I427748,I427841);
DFFARX1 I_25009 (I427807,I2683,I427674,I427663,);
nor I_25010 (I427889,I6858,I6864);
nand I_25011 (I427906,I427889,I6876);
nor I_25012 (I427923,I427906,I427790);
nand I_25013 (I427648,I427923,I6861);
DFFARX1 I_25014 (I427906,I2683,I427674,I427660,);
nand I_25015 (I427968,I427790,I6858);
nor I_25016 (I427985,I427790,I6858);
nand I_25017 (I427654,I427773,I427985);
not I_25018 (I428016,I6879);
nor I_25019 (I428033,I428016,I427968);
DFFARX1 I_25020 (I428033,I2683,I427674,I427642,);
nor I_25021 (I428064,I428016,I6861);
and I_25022 (I428081,I428064,I6870);
or I_25023 (I428098,I428081,I6864);
DFFARX1 I_25024 (I428098,I2683,I427674,I428124,);
nor I_25025 (I428132,I428124,I427748);
nor I_25026 (I427651,I427700,I428132);
not I_25027 (I428163,I428124);
nor I_25028 (I428180,I428163,I427858);
DFFARX1 I_25029 (I428180,I2683,I427674,I427657,);
nand I_25030 (I428211,I428163,I427790);
nor I_25031 (I427645,I428016,I428211);
not I_25032 (I428269,I2690);
DFFARX1 I_25033 (I667589,I2683,I428269,I428295,);
DFFARX1 I_25034 (I428295,I2683,I428269,I428312,);
not I_25035 (I428261,I428312);
DFFARX1 I_25036 (I667586,I2683,I428269,I428343,);
not I_25037 (I428351,I667586);
nor I_25038 (I428368,I428295,I428351);
not I_25039 (I428385,I667583);
not I_25040 (I428402,I667598);
nand I_25041 (I428419,I428402,I667583);
nor I_25042 (I428436,I428351,I428419);
nor I_25043 (I428453,I428343,I428436);
DFFARX1 I_25044 (I428402,I2683,I428269,I428258,);
nor I_25045 (I428484,I667598,I667592);
nand I_25046 (I428501,I428484,I667580);
nor I_25047 (I428518,I428501,I428385);
nand I_25048 (I428243,I428518,I667586);
DFFARX1 I_25049 (I428501,I2683,I428269,I428255,);
nand I_25050 (I428563,I428385,I667598);
nor I_25051 (I428580,I428385,I667598);
nand I_25052 (I428249,I428368,I428580);
not I_25053 (I428611,I667601);
nor I_25054 (I428628,I428611,I428563);
DFFARX1 I_25055 (I428628,I2683,I428269,I428237,);
nor I_25056 (I428659,I428611,I667580);
and I_25057 (I428676,I428659,I667595);
or I_25058 (I428693,I428676,I667583);
DFFARX1 I_25059 (I428693,I2683,I428269,I428719,);
nor I_25060 (I428727,I428719,I428343);
nor I_25061 (I428246,I428295,I428727);
not I_25062 (I428758,I428719);
nor I_25063 (I428775,I428758,I428453);
DFFARX1 I_25064 (I428775,I2683,I428269,I428252,);
nand I_25065 (I428806,I428758,I428385);
nor I_25066 (I428240,I428611,I428806);
not I_25067 (I428864,I2690);
DFFARX1 I_25068 (I528937,I2683,I428864,I428890,);
DFFARX1 I_25069 (I428890,I2683,I428864,I428907,);
not I_25070 (I428856,I428907);
DFFARX1 I_25071 (I528931,I2683,I428864,I428938,);
not I_25072 (I428946,I528928);
nor I_25073 (I428963,I428890,I428946);
not I_25074 (I428980,I528940);
not I_25075 (I428997,I528943);
nand I_25076 (I429014,I428997,I528940);
nor I_25077 (I429031,I428946,I429014);
nor I_25078 (I429048,I428938,I429031);
DFFARX1 I_25079 (I428997,I2683,I428864,I428853,);
nor I_25080 (I429079,I528943,I528952);
nand I_25081 (I429096,I429079,I528946);
nor I_25082 (I429113,I429096,I428980);
nand I_25083 (I428838,I429113,I528928);
DFFARX1 I_25084 (I429096,I2683,I428864,I428850,);
nand I_25085 (I429158,I428980,I528943);
nor I_25086 (I429175,I428980,I528943);
nand I_25087 (I428844,I428963,I429175);
not I_25088 (I429206,I528934);
nor I_25089 (I429223,I429206,I429158);
DFFARX1 I_25090 (I429223,I2683,I428864,I428832,);
nor I_25091 (I429254,I429206,I528949);
and I_25092 (I429271,I429254,I528928);
or I_25093 (I429288,I429271,I528931);
DFFARX1 I_25094 (I429288,I2683,I428864,I429314,);
nor I_25095 (I429322,I429314,I428938);
nor I_25096 (I428841,I428890,I429322);
not I_25097 (I429353,I429314);
nor I_25098 (I429370,I429353,I429048);
DFFARX1 I_25099 (I429370,I2683,I428864,I428847,);
nand I_25100 (I429401,I429353,I428980);
nor I_25101 (I428835,I429206,I429401);
not I_25102 (I429459,I2690);
DFFARX1 I_25103 (I687088,I2683,I429459,I429485,);
DFFARX1 I_25104 (I429485,I2683,I429459,I429502,);
not I_25105 (I429451,I429502);
DFFARX1 I_25106 (I687085,I2683,I429459,I429533,);
not I_25107 (I429541,I687085);
nor I_25108 (I429558,I429485,I429541);
not I_25109 (I429575,I687082);
not I_25110 (I429592,I687097);
nand I_25111 (I429609,I429592,I687082);
nor I_25112 (I429626,I429541,I429609);
nor I_25113 (I429643,I429533,I429626);
DFFARX1 I_25114 (I429592,I2683,I429459,I429448,);
nor I_25115 (I429674,I687097,I687091);
nand I_25116 (I429691,I429674,I687079);
nor I_25117 (I429708,I429691,I429575);
nand I_25118 (I429433,I429708,I687085);
DFFARX1 I_25119 (I429691,I2683,I429459,I429445,);
nand I_25120 (I429753,I429575,I687097);
nor I_25121 (I429770,I429575,I687097);
nand I_25122 (I429439,I429558,I429770);
not I_25123 (I429801,I687100);
nor I_25124 (I429818,I429801,I429753);
DFFARX1 I_25125 (I429818,I2683,I429459,I429427,);
nor I_25126 (I429849,I429801,I687079);
and I_25127 (I429866,I429849,I687094);
or I_25128 (I429883,I429866,I687082);
DFFARX1 I_25129 (I429883,I2683,I429459,I429909,);
nor I_25130 (I429917,I429909,I429533);
nor I_25131 (I429436,I429485,I429917);
not I_25132 (I429948,I429909);
nor I_25133 (I429965,I429948,I429643);
DFFARX1 I_25134 (I429965,I2683,I429459,I429442,);
nand I_25135 (I429996,I429948,I429575);
nor I_25136 (I429430,I429801,I429996);
not I_25137 (I430054,I2690);
DFFARX1 I_25138 (I363314,I2683,I430054,I430080,);
DFFARX1 I_25139 (I430080,I2683,I430054,I430097,);
not I_25140 (I430046,I430097);
DFFARX1 I_25141 (I363338,I2683,I430054,I430128,);
not I_25142 (I430136,I363317);
nor I_25143 (I430153,I430080,I430136);
not I_25144 (I430170,I363323);
not I_25145 (I430187,I363329);
nand I_25146 (I430204,I430187,I363323);
nor I_25147 (I430221,I430136,I430204);
nor I_25148 (I430238,I430128,I430221);
DFFARX1 I_25149 (I430187,I2683,I430054,I430043,);
nor I_25150 (I430269,I363329,I363341);
nand I_25151 (I430286,I430269,I363335);
nor I_25152 (I430303,I430286,I430170);
nand I_25153 (I430028,I430303,I363317);
DFFARX1 I_25154 (I430286,I2683,I430054,I430040,);
nand I_25155 (I430348,I430170,I363329);
nor I_25156 (I430365,I430170,I363329);
nand I_25157 (I430034,I430153,I430365);
not I_25158 (I430396,I363320);
nor I_25159 (I430413,I430396,I430348);
DFFARX1 I_25160 (I430413,I2683,I430054,I430022,);
nor I_25161 (I430444,I430396,I363314);
and I_25162 (I430461,I430444,I363332);
or I_25163 (I430478,I430461,I363326);
DFFARX1 I_25164 (I430478,I2683,I430054,I430504,);
nor I_25165 (I430512,I430504,I430128);
nor I_25166 (I430031,I430080,I430512);
not I_25167 (I430543,I430504);
nor I_25168 (I430560,I430543,I430238);
DFFARX1 I_25169 (I430560,I2683,I430054,I430037,);
nand I_25170 (I430591,I430543,I430170);
nor I_25171 (I430025,I430396,I430591);
not I_25172 (I430649,I2690);
DFFARX1 I_25173 (I887170,I2683,I430649,I430675,);
DFFARX1 I_25174 (I430675,I2683,I430649,I430692,);
not I_25175 (I430641,I430692);
DFFARX1 I_25176 (I887152,I2683,I430649,I430723,);
not I_25177 (I430731,I887158);
nor I_25178 (I430748,I430675,I430731);
not I_25179 (I430765,I887173);
not I_25180 (I430782,I887164);
nand I_25181 (I430799,I430782,I887173);
nor I_25182 (I430816,I430731,I430799);
nor I_25183 (I430833,I430723,I430816);
DFFARX1 I_25184 (I430782,I2683,I430649,I430638,);
nor I_25185 (I430864,I887164,I887176);
nand I_25186 (I430881,I430864,I887155);
nor I_25187 (I430898,I430881,I430765);
nand I_25188 (I430623,I430898,I887158);
DFFARX1 I_25189 (I430881,I2683,I430649,I430635,);
nand I_25190 (I430943,I430765,I887164);
nor I_25191 (I430960,I430765,I887164);
nand I_25192 (I430629,I430748,I430960);
not I_25193 (I430991,I887161);
nor I_25194 (I431008,I430991,I430943);
DFFARX1 I_25195 (I431008,I2683,I430649,I430617,);
nor I_25196 (I431039,I430991,I887167);
and I_25197 (I431056,I431039,I887152);
or I_25198 (I431073,I431056,I887155);
DFFARX1 I_25199 (I431073,I2683,I430649,I431099,);
nor I_25200 (I431107,I431099,I430723);
nor I_25201 (I430626,I430675,I431107);
not I_25202 (I431138,I431099);
nor I_25203 (I431155,I431138,I430833);
DFFARX1 I_25204 (I431155,I2683,I430649,I430632,);
nand I_25205 (I431186,I431138,I430765);
nor I_25206 (I430620,I430991,I431186);
not I_25207 (I431244,I2690);
DFFARX1 I_25208 (I60638,I2683,I431244,I431270,);
DFFARX1 I_25209 (I431270,I2683,I431244,I431287,);
not I_25210 (I431236,I431287);
DFFARX1 I_25211 (I60650,I2683,I431244,I431318,);
not I_25212 (I431326,I60641);
nor I_25213 (I431343,I431270,I431326);
not I_25214 (I431360,I60632);
not I_25215 (I431377,I60629);
nand I_25216 (I431394,I431377,I60632);
nor I_25217 (I431411,I431326,I431394);
nor I_25218 (I431428,I431318,I431411);
DFFARX1 I_25219 (I431377,I2683,I431244,I431233,);
nor I_25220 (I431459,I60629,I60629);
nand I_25221 (I431476,I431459,I60647);
nor I_25222 (I431493,I431476,I431360);
nand I_25223 (I431218,I431493,I60641);
DFFARX1 I_25224 (I431476,I2683,I431244,I431230,);
nand I_25225 (I431538,I431360,I60629);
nor I_25226 (I431555,I431360,I60629);
nand I_25227 (I431224,I431343,I431555);
not I_25228 (I431586,I60653);
nor I_25229 (I431603,I431586,I431538);
DFFARX1 I_25230 (I431603,I2683,I431244,I431212,);
nor I_25231 (I431634,I431586,I60632);
and I_25232 (I431651,I431634,I60635);
or I_25233 (I431668,I431651,I60644);
DFFARX1 I_25234 (I431668,I2683,I431244,I431694,);
nor I_25235 (I431702,I431694,I431318);
nor I_25236 (I431221,I431270,I431702);
not I_25237 (I431733,I431694);
nor I_25238 (I431750,I431733,I431428);
DFFARX1 I_25239 (I431750,I2683,I431244,I431227,);
nand I_25240 (I431781,I431733,I431360);
nor I_25241 (I431215,I431586,I431781);
not I_25242 (I431839,I2690);
DFFARX1 I_25243 (I103325,I2683,I431839,I431865,);
DFFARX1 I_25244 (I431865,I2683,I431839,I431882,);
not I_25245 (I431831,I431882);
DFFARX1 I_25246 (I103337,I2683,I431839,I431913,);
not I_25247 (I431921,I103328);
nor I_25248 (I431938,I431865,I431921);
not I_25249 (I431955,I103319);
not I_25250 (I431972,I103316);
nand I_25251 (I431989,I431972,I103319);
nor I_25252 (I432006,I431921,I431989);
nor I_25253 (I432023,I431913,I432006);
DFFARX1 I_25254 (I431972,I2683,I431839,I431828,);
nor I_25255 (I432054,I103316,I103316);
nand I_25256 (I432071,I432054,I103334);
nor I_25257 (I432088,I432071,I431955);
nand I_25258 (I431813,I432088,I103328);
DFFARX1 I_25259 (I432071,I2683,I431839,I431825,);
nand I_25260 (I432133,I431955,I103316);
nor I_25261 (I432150,I431955,I103316);
nand I_25262 (I431819,I431938,I432150);
not I_25263 (I432181,I103340);
nor I_25264 (I432198,I432181,I432133);
DFFARX1 I_25265 (I432198,I2683,I431839,I431807,);
nor I_25266 (I432229,I432181,I103319);
and I_25267 (I432246,I432229,I103322);
or I_25268 (I432263,I432246,I103331);
DFFARX1 I_25269 (I432263,I2683,I431839,I432289,);
nor I_25270 (I432297,I432289,I431913);
nor I_25271 (I431816,I431865,I432297);
not I_25272 (I432328,I432289);
nor I_25273 (I432345,I432328,I432023);
DFFARX1 I_25274 (I432345,I2683,I431839,I431822,);
nand I_25275 (I432376,I432328,I431955);
nor I_25276 (I431810,I432181,I432376);
not I_25277 (I432434,I2690);
DFFARX1 I_25278 (I968464,I2683,I432434,I432460,);
not I_25279 (I432468,I432460);
DFFARX1 I_25280 (I968458,I2683,I432434,I432494,);
not I_25281 (I432502,I968467);
nand I_25282 (I432519,I432502,I968446);
not I_25283 (I432536,I432519);
nor I_25284 (I432553,I432536,I968455);
nor I_25285 (I432570,I432468,I432553);
DFFARX1 I_25286 (I432570,I2683,I432434,I432420,);
not I_25287 (I432601,I968455);
nand I_25288 (I432618,I432601,I432536);
and I_25289 (I432635,I432601,I968470);
nand I_25290 (I432652,I432635,I968449);
nor I_25291 (I432417,I432652,I432601);
and I_25292 (I432408,I432494,I432652);
not I_25293 (I432697,I432652);
nand I_25294 (I432411,I432494,I432697);
nor I_25295 (I432405,I432460,I432652);
not I_25296 (I432742,I968452);
nor I_25297 (I432759,I432742,I968470);
nand I_25298 (I432776,I432759,I432601);
nor I_25299 (I432414,I432519,I432776);
nor I_25300 (I432807,I432742,I968461);
and I_25301 (I432824,I432807,I968449);
or I_25302 (I432841,I432824,I968446);
DFFARX1 I_25303 (I432841,I2683,I432434,I432867,);
nor I_25304 (I432875,I432867,I432618);
DFFARX1 I_25305 (I432875,I2683,I432434,I432402,);
DFFARX1 I_25306 (I432867,I2683,I432434,I432426,);
not I_25307 (I432920,I432867);
nor I_25308 (I432937,I432920,I432494);
nor I_25309 (I432954,I432759,I432937);
DFFARX1 I_25310 (I432954,I2683,I432434,I432423,);
not I_25311 (I433012,I2690);
DFFARX1 I_25312 (I200350,I2683,I433012,I433038,);
not I_25313 (I433046,I433038);
DFFARX1 I_25314 (I200335,I2683,I433012,I433072,);
not I_25315 (I433080,I200353);
nand I_25316 (I433097,I433080,I200338);
not I_25317 (I433114,I433097);
nor I_25318 (I433131,I433114,I200335);
nor I_25319 (I433148,I433046,I433131);
DFFARX1 I_25320 (I433148,I2683,I433012,I432998,);
not I_25321 (I433179,I200335);
nand I_25322 (I433196,I433179,I433114);
and I_25323 (I433213,I433179,I200338);
nand I_25324 (I433230,I433213,I200359);
nor I_25325 (I432995,I433230,I433179);
and I_25326 (I432986,I433072,I433230);
not I_25327 (I433275,I433230);
nand I_25328 (I432989,I433072,I433275);
nor I_25329 (I432983,I433038,I433230);
not I_25330 (I433320,I200347);
nor I_25331 (I433337,I433320,I200338);
nand I_25332 (I433354,I433337,I433179);
nor I_25333 (I432992,I433097,I433354);
nor I_25334 (I433385,I433320,I200341);
and I_25335 (I433402,I433385,I200356);
or I_25336 (I433419,I433402,I200344);
DFFARX1 I_25337 (I433419,I2683,I433012,I433445,);
nor I_25338 (I433453,I433445,I433196);
DFFARX1 I_25339 (I433453,I2683,I433012,I432980,);
DFFARX1 I_25340 (I433445,I2683,I433012,I433004,);
not I_25341 (I433498,I433445);
nor I_25342 (I433515,I433498,I433072);
nor I_25343 (I433532,I433337,I433515);
DFFARX1 I_25344 (I433532,I2683,I433012,I433001,);
not I_25345 (I433590,I2690);
DFFARX1 I_25346 (I817558,I2683,I433590,I433616,);
not I_25347 (I433624,I433616);
DFFARX1 I_25348 (I817549,I2683,I433590,I433650,);
not I_25349 (I433658,I817543);
nand I_25350 (I433675,I433658,I817555);
not I_25351 (I433692,I433675);
nor I_25352 (I433709,I433692,I817546);
nor I_25353 (I433726,I433624,I433709);
DFFARX1 I_25354 (I433726,I2683,I433590,I433576,);
not I_25355 (I433757,I817546);
nand I_25356 (I433774,I433757,I433692);
and I_25357 (I433791,I433757,I817552);
nand I_25358 (I433808,I433791,I817537);
nor I_25359 (I433573,I433808,I433757);
and I_25360 (I433564,I433650,I433808);
not I_25361 (I433853,I433808);
nand I_25362 (I433567,I433650,I433853);
nor I_25363 (I433561,I433616,I433808);
not I_25364 (I433898,I817537);
nor I_25365 (I433915,I433898,I817552);
nand I_25366 (I433932,I433915,I433757);
nor I_25367 (I433570,I433675,I433932);
nor I_25368 (I433963,I433898,I817540);
and I_25369 (I433980,I433963,I817543);
or I_25370 (I433997,I433980,I817540);
DFFARX1 I_25371 (I433997,I2683,I433590,I434023,);
nor I_25372 (I434031,I434023,I433774);
DFFARX1 I_25373 (I434031,I2683,I433590,I433558,);
DFFARX1 I_25374 (I434023,I2683,I433590,I433582,);
not I_25375 (I434076,I434023);
nor I_25376 (I434093,I434076,I433650);
nor I_25377 (I434110,I433915,I434093);
DFFARX1 I_25378 (I434110,I2683,I433590,I433579,);
not I_25379 (I434168,I2690);
DFFARX1 I_25380 (I664951,I2683,I434168,I434194,);
not I_25381 (I434202,I434194);
DFFARX1 I_25382 (I664951,I2683,I434168,I434228,);
not I_25383 (I434236,I664948);
nand I_25384 (I434253,I434236,I664963);
not I_25385 (I434270,I434253);
nor I_25386 (I434287,I434270,I664957);
nor I_25387 (I434304,I434202,I434287);
DFFARX1 I_25388 (I434304,I2683,I434168,I434154,);
not I_25389 (I434335,I664957);
nand I_25390 (I434352,I434335,I434270);
and I_25391 (I434369,I434335,I664954);
nand I_25392 (I434386,I434369,I664945);
nor I_25393 (I434151,I434386,I434335);
and I_25394 (I434142,I434228,I434386);
not I_25395 (I434431,I434386);
nand I_25396 (I434145,I434228,I434431);
nor I_25397 (I434139,I434194,I434386);
not I_25398 (I434476,I664966);
nor I_25399 (I434493,I434476,I664954);
nand I_25400 (I434510,I434493,I434335);
nor I_25401 (I434148,I434253,I434510);
nor I_25402 (I434541,I434476,I664945);
and I_25403 (I434558,I434541,I664948);
or I_25404 (I434575,I434558,I664960);
DFFARX1 I_25405 (I434575,I2683,I434168,I434601,);
nor I_25406 (I434609,I434601,I434352);
DFFARX1 I_25407 (I434609,I2683,I434168,I434136,);
DFFARX1 I_25408 (I434601,I2683,I434168,I434160,);
not I_25409 (I434654,I434601);
nor I_25410 (I434671,I434654,I434228);
nor I_25411 (I434688,I434493,I434671);
DFFARX1 I_25412 (I434688,I2683,I434168,I434157,);
not I_25413 (I434746,I2690);
DFFARX1 I_25414 (I121221,I2683,I434746,I434772,);
not I_25415 (I434780,I434772);
DFFARX1 I_25416 (I121200,I2683,I434746,I434806,);
not I_25417 (I434814,I121200);
nand I_25418 (I434831,I434814,I121227);
not I_25419 (I434848,I434831);
nor I_25420 (I434865,I434848,I121203);
nor I_25421 (I434882,I434780,I434865);
DFFARX1 I_25422 (I434882,I2683,I434746,I434732,);
not I_25423 (I434913,I121203);
nand I_25424 (I434930,I434913,I434848);
and I_25425 (I434947,I434913,I121224);
nand I_25426 (I434964,I434947,I121206);
nor I_25427 (I434729,I434964,I434913);
and I_25428 (I434720,I434806,I434964);
not I_25429 (I435009,I434964);
nand I_25430 (I434723,I434806,I435009);
nor I_25431 (I434717,I434772,I434964);
not I_25432 (I435054,I121209);
nor I_25433 (I435071,I435054,I121224);
nand I_25434 (I435088,I435071,I434913);
nor I_25435 (I434726,I434831,I435088);
nor I_25436 (I435119,I435054,I121215);
and I_25437 (I435136,I435119,I121212);
or I_25438 (I435153,I435136,I121218);
DFFARX1 I_25439 (I435153,I2683,I434746,I435179,);
nor I_25440 (I435187,I435179,I434930);
DFFARX1 I_25441 (I435187,I2683,I434746,I434714,);
DFFARX1 I_25442 (I435179,I2683,I434746,I434738,);
not I_25443 (I435232,I435179);
nor I_25444 (I435249,I435232,I434806);
nor I_25445 (I435266,I435071,I435249);
DFFARX1 I_25446 (I435266,I2683,I434746,I434735,);
not I_25447 (I435324,I2690);
DFFARX1 I_25448 (I431215,I2683,I435324,I435350,);
not I_25449 (I435358,I435350);
DFFARX1 I_25450 (I431227,I2683,I435324,I435384,);
not I_25451 (I435392,I431233);
nand I_25452 (I435409,I435392,I431224);
not I_25453 (I435426,I435409);
nor I_25454 (I435443,I435426,I431230);
nor I_25455 (I435460,I435358,I435443);
DFFARX1 I_25456 (I435460,I2683,I435324,I435310,);
not I_25457 (I435491,I431230);
nand I_25458 (I435508,I435491,I435426);
and I_25459 (I435525,I435491,I431221);
nand I_25460 (I435542,I435525,I431212);
nor I_25461 (I435307,I435542,I435491);
and I_25462 (I435298,I435384,I435542);
not I_25463 (I435587,I435542);
nand I_25464 (I435301,I435384,I435587);
nor I_25465 (I435295,I435350,I435542);
not I_25466 (I435632,I431218);
nor I_25467 (I435649,I435632,I431221);
nand I_25468 (I435666,I435649,I435491);
nor I_25469 (I435304,I435409,I435666);
nor I_25470 (I435697,I435632,I431215);
and I_25471 (I435714,I435697,I431212);
or I_25472 (I435731,I435714,I431236);
DFFARX1 I_25473 (I435731,I2683,I435324,I435757,);
nor I_25474 (I435765,I435757,I435508);
DFFARX1 I_25475 (I435765,I2683,I435324,I435292,);
DFFARX1 I_25476 (I435757,I2683,I435324,I435316,);
not I_25477 (I435810,I435757);
nor I_25478 (I435827,I435810,I435384);
nor I_25479 (I435844,I435649,I435827);
DFFARX1 I_25480 (I435844,I2683,I435324,I435313,);
not I_25481 (I435902,I2690);
DFFARX1 I_25482 (I246955,I2683,I435902,I435928,);
not I_25483 (I435936,I435928);
DFFARX1 I_25484 (I246970,I2683,I435902,I435962,);
not I_25485 (I435970,I246973);
nand I_25486 (I435987,I435970,I246952);
not I_25487 (I436004,I435987);
nor I_25488 (I436021,I436004,I246976);
nor I_25489 (I436038,I435936,I436021);
DFFARX1 I_25490 (I436038,I2683,I435902,I435888,);
not I_25491 (I436069,I246976);
nand I_25492 (I436086,I436069,I436004);
and I_25493 (I436103,I436069,I246958);
nand I_25494 (I436120,I436103,I246949);
nor I_25495 (I435885,I436120,I436069);
and I_25496 (I435876,I435962,I436120);
not I_25497 (I436165,I436120);
nand I_25498 (I435879,I435962,I436165);
nor I_25499 (I435873,I435928,I436120);
not I_25500 (I436210,I246949);
nor I_25501 (I436227,I436210,I246958);
nand I_25502 (I436244,I436227,I436069);
nor I_25503 (I435882,I435987,I436244);
nor I_25504 (I436275,I436210,I246964);
and I_25505 (I436292,I436275,I246967);
or I_25506 (I436309,I436292,I246961);
DFFARX1 I_25507 (I436309,I2683,I435902,I436335,);
nor I_25508 (I436343,I436335,I436086);
DFFARX1 I_25509 (I436343,I2683,I435902,I435870,);
DFFARX1 I_25510 (I436335,I2683,I435902,I435894,);
not I_25511 (I436388,I436335);
nor I_25512 (I436405,I436388,I435962);
nor I_25513 (I436422,I436227,I436405);
DFFARX1 I_25514 (I436422,I2683,I435902,I435891,);
not I_25515 (I436480,I2690);
DFFARX1 I_25516 (I219551,I2683,I436480,I436506,);
not I_25517 (I436514,I436506);
DFFARX1 I_25518 (I219566,I2683,I436480,I436540,);
not I_25519 (I436548,I219569);
nand I_25520 (I436565,I436548,I219548);
not I_25521 (I436582,I436565);
nor I_25522 (I436599,I436582,I219572);
nor I_25523 (I436616,I436514,I436599);
DFFARX1 I_25524 (I436616,I2683,I436480,I436466,);
not I_25525 (I436647,I219572);
nand I_25526 (I436664,I436647,I436582);
and I_25527 (I436681,I436647,I219554);
nand I_25528 (I436698,I436681,I219545);
nor I_25529 (I436463,I436698,I436647);
and I_25530 (I436454,I436540,I436698);
not I_25531 (I436743,I436698);
nand I_25532 (I436457,I436540,I436743);
nor I_25533 (I436451,I436506,I436698);
not I_25534 (I436788,I219545);
nor I_25535 (I436805,I436788,I219554);
nand I_25536 (I436822,I436805,I436647);
nor I_25537 (I436460,I436565,I436822);
nor I_25538 (I436853,I436788,I219560);
and I_25539 (I436870,I436853,I219563);
or I_25540 (I436887,I436870,I219557);
DFFARX1 I_25541 (I436887,I2683,I436480,I436913,);
nor I_25542 (I436921,I436913,I436664);
DFFARX1 I_25543 (I436921,I2683,I436480,I436448,);
DFFARX1 I_25544 (I436913,I2683,I436480,I436472,);
not I_25545 (I436966,I436913);
nor I_25546 (I436983,I436966,I436540);
nor I_25547 (I437000,I436805,I436983);
DFFARX1 I_25548 (I437000,I2683,I436480,I436469,);
not I_25549 (I437058,I2690);
DFFARX1 I_25550 (I1027113,I2683,I437058,I437084,);
not I_25551 (I437092,I437084);
DFFARX1 I_25552 (I1027131,I2683,I437058,I437118,);
not I_25553 (I437126,I1027128);
nand I_25554 (I437143,I437126,I1027119);
not I_25555 (I437160,I437143);
nor I_25556 (I437177,I437160,I1027116);
nor I_25557 (I437194,I437092,I437177);
DFFARX1 I_25558 (I437194,I2683,I437058,I437044,);
not I_25559 (I437225,I1027116);
nand I_25560 (I437242,I437225,I437160);
and I_25561 (I437259,I437225,I1027122);
nand I_25562 (I437276,I437259,I1027137);
nor I_25563 (I437041,I437276,I437225);
and I_25564 (I437032,I437118,I437276);
not I_25565 (I437321,I437276);
nand I_25566 (I437035,I437118,I437321);
nor I_25567 (I437029,I437084,I437276);
not I_25568 (I437366,I1027113);
nor I_25569 (I437383,I437366,I1027122);
nand I_25570 (I437400,I437383,I437225);
nor I_25571 (I437038,I437143,I437400);
nor I_25572 (I437431,I437366,I1027134);
and I_25573 (I437448,I437431,I1027125);
or I_25574 (I437465,I437448,I1027140);
DFFARX1 I_25575 (I437465,I2683,I437058,I437491,);
nor I_25576 (I437499,I437491,I437242);
DFFARX1 I_25577 (I437499,I2683,I437058,I437026,);
DFFARX1 I_25578 (I437491,I2683,I437058,I437050,);
not I_25579 (I437544,I437491);
nor I_25580 (I437561,I437544,I437118);
nor I_25581 (I437578,I437383,I437561);
DFFARX1 I_25582 (I437578,I2683,I437058,I437047,);
not I_25583 (I437636,I2690);
DFFARX1 I_25584 (I587306,I2683,I437636,I437662,);
not I_25585 (I437670,I437662);
DFFARX1 I_25586 (I587318,I2683,I437636,I437696,);
not I_25587 (I437704,I587309);
nand I_25588 (I437721,I437704,I587312);
not I_25589 (I437738,I437721);
nor I_25590 (I437755,I437738,I587315);
nor I_25591 (I437772,I437670,I437755);
DFFARX1 I_25592 (I437772,I2683,I437636,I437622,);
not I_25593 (I437803,I587315);
nand I_25594 (I437820,I437803,I437738);
and I_25595 (I437837,I437803,I587309);
nand I_25596 (I437854,I437837,I587321);
nor I_25597 (I437619,I437854,I437803);
and I_25598 (I437610,I437696,I437854);
not I_25599 (I437899,I437854);
nand I_25600 (I437613,I437696,I437899);
nor I_25601 (I437607,I437662,I437854);
not I_25602 (I437944,I587327);
nor I_25603 (I437961,I437944,I587309);
nand I_25604 (I437978,I437961,I437803);
nor I_25605 (I437616,I437721,I437978);
nor I_25606 (I438009,I437944,I587306);
and I_25607 (I438026,I438009,I587324);
or I_25608 (I438043,I438026,I587330);
DFFARX1 I_25609 (I438043,I2683,I437636,I438069,);
nor I_25610 (I438077,I438069,I437820);
DFFARX1 I_25611 (I438077,I2683,I437636,I437604,);
DFFARX1 I_25612 (I438069,I2683,I437636,I437628,);
not I_25613 (I438122,I438069);
nor I_25614 (I438139,I438122,I437696);
nor I_25615 (I438156,I437961,I438139);
DFFARX1 I_25616 (I438156,I2683,I437636,I437625,);
not I_25617 (I438214,I2690);
DFFARX1 I_25618 (I923566,I2683,I438214,I438240,);
not I_25619 (I438248,I438240);
DFFARX1 I_25620 (I923572,I2683,I438214,I438274,);
not I_25621 (I438282,I923566);
nand I_25622 (I438299,I438282,I923569);
not I_25623 (I438316,I438299);
nor I_25624 (I438333,I438316,I923587);
nor I_25625 (I438350,I438248,I438333);
DFFARX1 I_25626 (I438350,I2683,I438214,I438200,);
not I_25627 (I438381,I923587);
nand I_25628 (I438398,I438381,I438316);
and I_25629 (I438415,I438381,I923590);
nand I_25630 (I438432,I438415,I923569);
nor I_25631 (I438197,I438432,I438381);
and I_25632 (I438188,I438274,I438432);
not I_25633 (I438477,I438432);
nand I_25634 (I438191,I438274,I438477);
nor I_25635 (I438185,I438240,I438432);
not I_25636 (I438522,I923575);
nor I_25637 (I438539,I438522,I923590);
nand I_25638 (I438556,I438539,I438381);
nor I_25639 (I438194,I438299,I438556);
nor I_25640 (I438587,I438522,I923581);
and I_25641 (I438604,I438587,I923578);
or I_25642 (I438621,I438604,I923584);
DFFARX1 I_25643 (I438621,I2683,I438214,I438647,);
nor I_25644 (I438655,I438647,I438398);
DFFARX1 I_25645 (I438655,I2683,I438214,I438182,);
DFFARX1 I_25646 (I438647,I2683,I438214,I438206,);
not I_25647 (I438700,I438647);
nor I_25648 (I438717,I438700,I438274);
nor I_25649 (I438734,I438539,I438717);
DFFARX1 I_25650 (I438734,I2683,I438214,I438203,);
not I_25651 (I438792,I2690);
DFFARX1 I_25652 (I846114,I2683,I438792,I438818,);
not I_25653 (I438826,I438818);
DFFARX1 I_25654 (I846120,I2683,I438792,I438852,);
not I_25655 (I438860,I846114);
nand I_25656 (I438877,I438860,I846117);
not I_25657 (I438894,I438877);
nor I_25658 (I438911,I438894,I846135);
nor I_25659 (I438928,I438826,I438911);
DFFARX1 I_25660 (I438928,I2683,I438792,I438778,);
not I_25661 (I438959,I846135);
nand I_25662 (I438976,I438959,I438894);
and I_25663 (I438993,I438959,I846138);
nand I_25664 (I439010,I438993,I846117);
nor I_25665 (I438775,I439010,I438959);
and I_25666 (I438766,I438852,I439010);
not I_25667 (I439055,I439010);
nand I_25668 (I438769,I438852,I439055);
nor I_25669 (I438763,I438818,I439010);
not I_25670 (I439100,I846123);
nor I_25671 (I439117,I439100,I846138);
nand I_25672 (I439134,I439117,I438959);
nor I_25673 (I438772,I438877,I439134);
nor I_25674 (I439165,I439100,I846129);
and I_25675 (I439182,I439165,I846126);
or I_25676 (I439199,I439182,I846132);
DFFARX1 I_25677 (I439199,I2683,I438792,I439225,);
nor I_25678 (I439233,I439225,I438976);
DFFARX1 I_25679 (I439233,I2683,I438792,I438760,);
DFFARX1 I_25680 (I439225,I2683,I438792,I438784,);
not I_25681 (I439278,I439225);
nor I_25682 (I439295,I439278,I438852);
nor I_25683 (I439312,I439117,I439295);
DFFARX1 I_25684 (I439312,I2683,I438792,I438781,);
not I_25685 (I439370,I2690);
DFFARX1 I_25686 (I980432,I2683,I439370,I439396,);
not I_25687 (I439404,I439396);
DFFARX1 I_25688 (I980426,I2683,I439370,I439430,);
not I_25689 (I439438,I980435);
nand I_25690 (I439455,I439438,I980414);
not I_25691 (I439472,I439455);
nor I_25692 (I439489,I439472,I980423);
nor I_25693 (I439506,I439404,I439489);
DFFARX1 I_25694 (I439506,I2683,I439370,I439356,);
not I_25695 (I439537,I980423);
nand I_25696 (I439554,I439537,I439472);
and I_25697 (I439571,I439537,I980438);
nand I_25698 (I439588,I439571,I980417);
nor I_25699 (I439353,I439588,I439537);
and I_25700 (I439344,I439430,I439588);
not I_25701 (I439633,I439588);
nand I_25702 (I439347,I439430,I439633);
nor I_25703 (I439341,I439396,I439588);
not I_25704 (I439678,I980420);
nor I_25705 (I439695,I439678,I980438);
nand I_25706 (I439712,I439695,I439537);
nor I_25707 (I439350,I439455,I439712);
nor I_25708 (I439743,I439678,I980429);
and I_25709 (I439760,I439743,I980417);
or I_25710 (I439777,I439760,I980414);
DFFARX1 I_25711 (I439777,I2683,I439370,I439803,);
nor I_25712 (I439811,I439803,I439554);
DFFARX1 I_25713 (I439811,I2683,I439370,I439338,);
DFFARX1 I_25714 (I439803,I2683,I439370,I439362,);
not I_25715 (I439856,I439803);
nor I_25716 (I439873,I439856,I439430);
nor I_25717 (I439890,I439695,I439873);
DFFARX1 I_25718 (I439890,I2683,I439370,I439359,);
not I_25719 (I439948,I2690);
DFFARX1 I_25720 (I948420,I2683,I439948,I439974,);
not I_25721 (I439982,I439974);
DFFARX1 I_25722 (I948426,I2683,I439948,I440008,);
not I_25723 (I440016,I948420);
nand I_25724 (I440033,I440016,I948423);
not I_25725 (I440050,I440033);
nor I_25726 (I440067,I440050,I948441);
nor I_25727 (I440084,I439982,I440067);
DFFARX1 I_25728 (I440084,I2683,I439948,I439934,);
not I_25729 (I440115,I948441);
nand I_25730 (I440132,I440115,I440050);
and I_25731 (I440149,I440115,I948444);
nand I_25732 (I440166,I440149,I948423);
nor I_25733 (I439931,I440166,I440115);
and I_25734 (I439922,I440008,I440166);
not I_25735 (I440211,I440166);
nand I_25736 (I439925,I440008,I440211);
nor I_25737 (I439919,I439974,I440166);
not I_25738 (I440256,I948429);
nor I_25739 (I440273,I440256,I948444);
nand I_25740 (I440290,I440273,I440115);
nor I_25741 (I439928,I440033,I440290);
nor I_25742 (I440321,I440256,I948435);
and I_25743 (I440338,I440321,I948432);
or I_25744 (I440355,I440338,I948438);
DFFARX1 I_25745 (I440355,I2683,I439948,I440381,);
nor I_25746 (I440389,I440381,I440132);
DFFARX1 I_25747 (I440389,I2683,I439948,I439916,);
DFFARX1 I_25748 (I440381,I2683,I439948,I439940,);
not I_25749 (I440434,I440381);
nor I_25750 (I440451,I440434,I440008);
nor I_25751 (I440468,I440273,I440451);
DFFARX1 I_25752 (I440468,I2683,I439948,I439937,);
not I_25753 (I440526,I2690);
DFFARX1 I_25754 (I1021503,I2683,I440526,I440552,);
not I_25755 (I440560,I440552);
DFFARX1 I_25756 (I1021521,I2683,I440526,I440586,);
not I_25757 (I440594,I1021518);
nand I_25758 (I440611,I440594,I1021509);
not I_25759 (I440628,I440611);
nor I_25760 (I440645,I440628,I1021506);
nor I_25761 (I440662,I440560,I440645);
DFFARX1 I_25762 (I440662,I2683,I440526,I440512,);
not I_25763 (I440693,I1021506);
nand I_25764 (I440710,I440693,I440628);
and I_25765 (I440727,I440693,I1021512);
nand I_25766 (I440744,I440727,I1021527);
nor I_25767 (I440509,I440744,I440693);
and I_25768 (I440500,I440586,I440744);
not I_25769 (I440789,I440744);
nand I_25770 (I440503,I440586,I440789);
nor I_25771 (I440497,I440552,I440744);
not I_25772 (I440834,I1021503);
nor I_25773 (I440851,I440834,I1021512);
nand I_25774 (I440868,I440851,I440693);
nor I_25775 (I440506,I440611,I440868);
nor I_25776 (I440899,I440834,I1021524);
and I_25777 (I440916,I440899,I1021515);
or I_25778 (I440933,I440916,I1021530);
DFFARX1 I_25779 (I440933,I2683,I440526,I440959,);
nor I_25780 (I440967,I440959,I440710);
DFFARX1 I_25781 (I440967,I2683,I440526,I440494,);
DFFARX1 I_25782 (I440959,I2683,I440526,I440518,);
not I_25783 (I441012,I440959);
nor I_25784 (I441029,I441012,I440586);
nor I_25785 (I441046,I440851,I441029);
DFFARX1 I_25786 (I441046,I2683,I440526,I440515,);
not I_25787 (I441104,I2690);
DFFARX1 I_25788 (I312830,I2683,I441104,I441130,);
not I_25789 (I441138,I441130);
DFFARX1 I_25790 (I312845,I2683,I441104,I441164,);
not I_25791 (I441172,I312848);
nand I_25792 (I441189,I441172,I312827);
not I_25793 (I441206,I441189);
nor I_25794 (I441223,I441206,I312851);
nor I_25795 (I441240,I441138,I441223);
DFFARX1 I_25796 (I441240,I2683,I441104,I441090,);
not I_25797 (I441271,I312851);
nand I_25798 (I441288,I441271,I441206);
and I_25799 (I441305,I441271,I312833);
nand I_25800 (I441322,I441305,I312824);
nor I_25801 (I441087,I441322,I441271);
and I_25802 (I441078,I441164,I441322);
not I_25803 (I441367,I441322);
nand I_25804 (I441081,I441164,I441367);
nor I_25805 (I441075,I441130,I441322);
not I_25806 (I441412,I312824);
nor I_25807 (I441429,I441412,I312833);
nand I_25808 (I441446,I441429,I441271);
nor I_25809 (I441084,I441189,I441446);
nor I_25810 (I441477,I441412,I312839);
and I_25811 (I441494,I441477,I312842);
or I_25812 (I441511,I441494,I312836);
DFFARX1 I_25813 (I441511,I2683,I441104,I441537,);
nor I_25814 (I441545,I441537,I441288);
DFFARX1 I_25815 (I441545,I2683,I441104,I441072,);
DFFARX1 I_25816 (I441537,I2683,I441104,I441096,);
not I_25817 (I441590,I441537);
nor I_25818 (I441607,I441590,I441164);
nor I_25819 (I441624,I441429,I441607);
DFFARX1 I_25820 (I441624,I2683,I441104,I441093,);
not I_25821 (I441682,I2690);
DFFARX1 I_25822 (I523148,I2683,I441682,I441708,);
not I_25823 (I441716,I441708);
DFFARX1 I_25824 (I523160,I2683,I441682,I441742,);
not I_25825 (I441750,I523151);
nand I_25826 (I441767,I441750,I523154);
not I_25827 (I441784,I441767);
nor I_25828 (I441801,I441784,I523157);
nor I_25829 (I441818,I441716,I441801);
DFFARX1 I_25830 (I441818,I2683,I441682,I441668,);
not I_25831 (I441849,I523157);
nand I_25832 (I441866,I441849,I441784);
and I_25833 (I441883,I441849,I523151);
nand I_25834 (I441900,I441883,I523163);
nor I_25835 (I441665,I441900,I441849);
and I_25836 (I441656,I441742,I441900);
not I_25837 (I441945,I441900);
nand I_25838 (I441659,I441742,I441945);
nor I_25839 (I441653,I441708,I441900);
not I_25840 (I441990,I523169);
nor I_25841 (I442007,I441990,I523151);
nand I_25842 (I442024,I442007,I441849);
nor I_25843 (I441662,I441767,I442024);
nor I_25844 (I442055,I441990,I523148);
and I_25845 (I442072,I442055,I523166);
or I_25846 (I442089,I442072,I523172);
DFFARX1 I_25847 (I442089,I2683,I441682,I442115,);
nor I_25848 (I442123,I442115,I441866);
DFFARX1 I_25849 (I442123,I2683,I441682,I441650,);
DFFARX1 I_25850 (I442115,I2683,I441682,I441674,);
not I_25851 (I442168,I442115);
nor I_25852 (I442185,I442168,I441742);
nor I_25853 (I442202,I442007,I442185);
DFFARX1 I_25854 (I442202,I2683,I441682,I441671,);
not I_25855 (I442260,I2690);
DFFARX1 I_25856 (I415745,I2683,I442260,I442286,);
not I_25857 (I442294,I442286);
DFFARX1 I_25858 (I415757,I2683,I442260,I442320,);
not I_25859 (I442328,I415763);
nand I_25860 (I442345,I442328,I415754);
not I_25861 (I442362,I442345);
nor I_25862 (I442379,I442362,I415760);
nor I_25863 (I442396,I442294,I442379);
DFFARX1 I_25864 (I442396,I2683,I442260,I442246,);
not I_25865 (I442427,I415760);
nand I_25866 (I442444,I442427,I442362);
and I_25867 (I442461,I442427,I415751);
nand I_25868 (I442478,I442461,I415742);
nor I_25869 (I442243,I442478,I442427);
and I_25870 (I442234,I442320,I442478);
not I_25871 (I442523,I442478);
nand I_25872 (I442237,I442320,I442523);
nor I_25873 (I442231,I442286,I442478);
not I_25874 (I442568,I415748);
nor I_25875 (I442585,I442568,I415751);
nand I_25876 (I442602,I442585,I442427);
nor I_25877 (I442240,I442345,I442602);
nor I_25878 (I442633,I442568,I415745);
and I_25879 (I442650,I442633,I415742);
or I_25880 (I442667,I442650,I415766);
DFFARX1 I_25881 (I442667,I2683,I442260,I442693,);
nor I_25882 (I442701,I442693,I442444);
DFFARX1 I_25883 (I442701,I2683,I442260,I442228,);
DFFARX1 I_25884 (I442693,I2683,I442260,I442252,);
not I_25885 (I442746,I442693);
nor I_25886 (I442763,I442746,I442320);
nor I_25887 (I442780,I442585,I442763);
DFFARX1 I_25888 (I442780,I2683,I442260,I442249,);
not I_25889 (I442838,I2690);
DFFARX1 I_25890 (I953044,I2683,I442838,I442864,);
not I_25891 (I442872,I442864);
DFFARX1 I_25892 (I953050,I2683,I442838,I442898,);
not I_25893 (I442906,I953044);
nand I_25894 (I442923,I442906,I953047);
not I_25895 (I442940,I442923);
nor I_25896 (I442957,I442940,I953065);
nor I_25897 (I442974,I442872,I442957);
DFFARX1 I_25898 (I442974,I2683,I442838,I442824,);
not I_25899 (I443005,I953065);
nand I_25900 (I443022,I443005,I442940);
and I_25901 (I443039,I443005,I953068);
nand I_25902 (I443056,I443039,I953047);
nor I_25903 (I442821,I443056,I443005);
and I_25904 (I442812,I442898,I443056);
not I_25905 (I443101,I443056);
nand I_25906 (I442815,I442898,I443101);
nor I_25907 (I442809,I442864,I443056);
not I_25908 (I443146,I953053);
nor I_25909 (I443163,I443146,I953068);
nand I_25910 (I443180,I443163,I443005);
nor I_25911 (I442818,I442923,I443180);
nor I_25912 (I443211,I443146,I953059);
and I_25913 (I443228,I443211,I953056);
or I_25914 (I443245,I443228,I953062);
DFFARX1 I_25915 (I443245,I2683,I442838,I443271,);
nor I_25916 (I443279,I443271,I443022);
DFFARX1 I_25917 (I443279,I2683,I442838,I442806,);
DFFARX1 I_25918 (I443271,I2683,I442838,I442830,);
not I_25919 (I443324,I443271);
nor I_25920 (I443341,I443324,I442898);
nor I_25921 (I443358,I443163,I443341);
DFFARX1 I_25922 (I443358,I2683,I442838,I442827,);
not I_25923 (I443416,I2690);
DFFARX1 I_25924 (I913740,I2683,I443416,I443442,);
not I_25925 (I443450,I443442);
DFFARX1 I_25926 (I913746,I2683,I443416,I443476,);
not I_25927 (I443484,I913740);
nand I_25928 (I443501,I443484,I913743);
not I_25929 (I443518,I443501);
nor I_25930 (I443535,I443518,I913761);
nor I_25931 (I443552,I443450,I443535);
DFFARX1 I_25932 (I443552,I2683,I443416,I443402,);
not I_25933 (I443583,I913761);
nand I_25934 (I443600,I443583,I443518);
and I_25935 (I443617,I443583,I913764);
nand I_25936 (I443634,I443617,I913743);
nor I_25937 (I443399,I443634,I443583);
and I_25938 (I443390,I443476,I443634);
not I_25939 (I443679,I443634);
nand I_25940 (I443393,I443476,I443679);
nor I_25941 (I443387,I443442,I443634);
not I_25942 (I443724,I913749);
nor I_25943 (I443741,I443724,I913764);
nand I_25944 (I443758,I443741,I443583);
nor I_25945 (I443396,I443501,I443758);
nor I_25946 (I443789,I443724,I913755);
and I_25947 (I443806,I443789,I913752);
or I_25948 (I443823,I443806,I913758);
DFFARX1 I_25949 (I443823,I2683,I443416,I443849,);
nor I_25950 (I443857,I443849,I443600);
DFFARX1 I_25951 (I443857,I2683,I443416,I443384,);
DFFARX1 I_25952 (I443849,I2683,I443416,I443408,);
not I_25953 (I443902,I443849);
nor I_25954 (I443919,I443902,I443476);
nor I_25955 (I443936,I443741,I443919);
DFFARX1 I_25956 (I443936,I2683,I443416,I443405,);
not I_25957 (I443994,I2690);
DFFARX1 I_25958 (I854206,I2683,I443994,I444020,);
not I_25959 (I444028,I444020);
DFFARX1 I_25960 (I854212,I2683,I443994,I444054,);
not I_25961 (I444062,I854206);
nand I_25962 (I444079,I444062,I854209);
not I_25963 (I444096,I444079);
nor I_25964 (I444113,I444096,I854227);
nor I_25965 (I444130,I444028,I444113);
DFFARX1 I_25966 (I444130,I2683,I443994,I443980,);
not I_25967 (I444161,I854227);
nand I_25968 (I444178,I444161,I444096);
and I_25969 (I444195,I444161,I854230);
nand I_25970 (I444212,I444195,I854209);
nor I_25971 (I443977,I444212,I444161);
and I_25972 (I443968,I444054,I444212);
not I_25973 (I444257,I444212);
nand I_25974 (I443971,I444054,I444257);
nor I_25975 (I443965,I444020,I444212);
not I_25976 (I444302,I854215);
nor I_25977 (I444319,I444302,I854230);
nand I_25978 (I444336,I444319,I444161);
nor I_25979 (I443974,I444079,I444336);
nor I_25980 (I444367,I444302,I854221);
and I_25981 (I444384,I444367,I854218);
or I_25982 (I444401,I444384,I854224);
DFFARX1 I_25983 (I444401,I2683,I443994,I444427,);
nor I_25984 (I444435,I444427,I444178);
DFFARX1 I_25985 (I444435,I2683,I443994,I443962,);
DFFARX1 I_25986 (I444427,I2683,I443994,I443986,);
not I_25987 (I444480,I444427);
nor I_25988 (I444497,I444480,I444054);
nor I_25989 (I444514,I444319,I444497);
DFFARX1 I_25990 (I444514,I2683,I443994,I443983,);
not I_25991 (I444572,I2690);
DFFARX1 I_25992 (I979344,I2683,I444572,I444598,);
not I_25993 (I444606,I444598);
DFFARX1 I_25994 (I979338,I2683,I444572,I444632,);
not I_25995 (I444640,I979347);
nand I_25996 (I444657,I444640,I979326);
not I_25997 (I444674,I444657);
nor I_25998 (I444691,I444674,I979335);
nor I_25999 (I444708,I444606,I444691);
DFFARX1 I_26000 (I444708,I2683,I444572,I444558,);
not I_26001 (I444739,I979335);
nand I_26002 (I444756,I444739,I444674);
and I_26003 (I444773,I444739,I979350);
nand I_26004 (I444790,I444773,I979329);
nor I_26005 (I444555,I444790,I444739);
and I_26006 (I444546,I444632,I444790);
not I_26007 (I444835,I444790);
nand I_26008 (I444549,I444632,I444835);
nor I_26009 (I444543,I444598,I444790);
not I_26010 (I444880,I979332);
nor I_26011 (I444897,I444880,I979350);
nand I_26012 (I444914,I444897,I444739);
nor I_26013 (I444552,I444657,I444914);
nor I_26014 (I444945,I444880,I979341);
and I_26015 (I444962,I444945,I979329);
or I_26016 (I444979,I444962,I979326);
DFFARX1 I_26017 (I444979,I2683,I444572,I445005,);
nor I_26018 (I445013,I445005,I444756);
DFFARX1 I_26019 (I445013,I2683,I444572,I444540,);
DFFARX1 I_26020 (I445005,I2683,I444572,I444564,);
not I_26021 (I445058,I445005);
nor I_26022 (I445075,I445058,I444632);
nor I_26023 (I445092,I444897,I445075);
DFFARX1 I_26024 (I445092,I2683,I444572,I444561,);
not I_26025 (I445150,I2690);
DFFARX1 I_26026 (I1034644,I2683,I445150,I445176,);
not I_26027 (I445184,I445176);
DFFARX1 I_26028 (I1034644,I2683,I445150,I445210,);
not I_26029 (I445218,I1034668);
nand I_26030 (I445235,I445218,I1034650);
not I_26031 (I445252,I445235);
nor I_26032 (I445269,I445252,I1034665);
nor I_26033 (I445286,I445184,I445269);
DFFARX1 I_26034 (I445286,I2683,I445150,I445136,);
not I_26035 (I445317,I1034665);
nand I_26036 (I445334,I445317,I445252);
and I_26037 (I445351,I445317,I1034647);
nand I_26038 (I445368,I445351,I1034656);
nor I_26039 (I445133,I445368,I445317);
and I_26040 (I445124,I445210,I445368);
not I_26041 (I445413,I445368);
nand I_26042 (I445127,I445210,I445413);
nor I_26043 (I445121,I445176,I445368);
not I_26044 (I445458,I1034653);
nor I_26045 (I445475,I445458,I1034647);
nand I_26046 (I445492,I445475,I445317);
nor I_26047 (I445130,I445235,I445492);
nor I_26048 (I445523,I445458,I1034662);
and I_26049 (I445540,I445523,I1034671);
or I_26050 (I445557,I445540,I1034659);
DFFARX1 I_26051 (I445557,I2683,I445150,I445583,);
nor I_26052 (I445591,I445583,I445334);
DFFARX1 I_26053 (I445591,I2683,I445150,I445118,);
DFFARX1 I_26054 (I445583,I2683,I445150,I445142,);
not I_26055 (I445636,I445583);
nor I_26056 (I445653,I445636,I445210);
nor I_26057 (I445670,I445475,I445653);
DFFARX1 I_26058 (I445670,I2683,I445150,I445139,);
not I_26059 (I445728,I2690);
DFFARX1 I_26060 (I861142,I2683,I445728,I445754,);
not I_26061 (I445762,I445754);
DFFARX1 I_26062 (I861148,I2683,I445728,I445788,);
not I_26063 (I445796,I861142);
nand I_26064 (I445813,I445796,I861145);
not I_26065 (I445830,I445813);
nor I_26066 (I445847,I445830,I861163);
nor I_26067 (I445864,I445762,I445847);
DFFARX1 I_26068 (I445864,I2683,I445728,I445714,);
not I_26069 (I445895,I861163);
nand I_26070 (I445912,I445895,I445830);
and I_26071 (I445929,I445895,I861166);
nand I_26072 (I445946,I445929,I861145);
nor I_26073 (I445711,I445946,I445895);
and I_26074 (I445702,I445788,I445946);
not I_26075 (I445991,I445946);
nand I_26076 (I445705,I445788,I445991);
nor I_26077 (I445699,I445754,I445946);
not I_26078 (I446036,I861151);
nor I_26079 (I446053,I446036,I861166);
nand I_26080 (I446070,I446053,I445895);
nor I_26081 (I445708,I445813,I446070);
nor I_26082 (I446101,I446036,I861157);
and I_26083 (I446118,I446101,I861154);
or I_26084 (I446135,I446118,I861160);
DFFARX1 I_26085 (I446135,I2683,I445728,I446161,);
nor I_26086 (I446169,I446161,I445912);
DFFARX1 I_26087 (I446169,I2683,I445728,I445696,);
DFFARX1 I_26088 (I446161,I2683,I445728,I445720,);
not I_26089 (I446214,I446161);
nor I_26090 (I446231,I446214,I445788);
nor I_26091 (I446248,I446053,I446231);
DFFARX1 I_26092 (I446248,I2683,I445728,I445717,);
not I_26093 (I446306,I2690);
DFFARX1 I_26094 (I699971,I2683,I446306,I446332,);
not I_26095 (I446340,I446332);
DFFARX1 I_26096 (I699968,I2683,I446306,I446366,);
not I_26097 (I446374,I699965);
nand I_26098 (I446391,I446374,I699992);
not I_26099 (I446408,I446391);
nor I_26100 (I446425,I446408,I699980);
nor I_26101 (I446442,I446340,I446425);
DFFARX1 I_26102 (I446442,I2683,I446306,I446292,);
not I_26103 (I446473,I699980);
nand I_26104 (I446490,I446473,I446408);
and I_26105 (I446507,I446473,I699986);
nand I_26106 (I446524,I446507,I699977);
nor I_26107 (I446289,I446524,I446473);
and I_26108 (I446280,I446366,I446524);
not I_26109 (I446569,I446524);
nand I_26110 (I446283,I446366,I446569);
nor I_26111 (I446277,I446332,I446524);
not I_26112 (I446614,I699974);
nor I_26113 (I446631,I446614,I699986);
nand I_26114 (I446648,I446631,I446473);
nor I_26115 (I446286,I446391,I446648);
nor I_26116 (I446679,I446614,I699989);
and I_26117 (I446696,I446679,I699983);
or I_26118 (I446713,I446696,I699965);
DFFARX1 I_26119 (I446713,I2683,I446306,I446739,);
nor I_26120 (I446747,I446739,I446490);
DFFARX1 I_26121 (I446747,I2683,I446306,I446274,);
DFFARX1 I_26122 (I446739,I2683,I446306,I446298,);
not I_26123 (I446792,I446739);
nor I_26124 (I446809,I446792,I446366);
nor I_26125 (I446826,I446631,I446809);
DFFARX1 I_26126 (I446826,I2683,I446306,I446295,);
not I_26127 (I446884,I2690);
DFFARX1 I_26128 (I857096,I2683,I446884,I446910,);
not I_26129 (I446918,I446910);
DFFARX1 I_26130 (I857102,I2683,I446884,I446944,);
not I_26131 (I446952,I857096);
nand I_26132 (I446969,I446952,I857099);
not I_26133 (I446986,I446969);
nor I_26134 (I447003,I446986,I857117);
nor I_26135 (I447020,I446918,I447003);
DFFARX1 I_26136 (I447020,I2683,I446884,I446870,);
not I_26137 (I447051,I857117);
nand I_26138 (I447068,I447051,I446986);
and I_26139 (I447085,I447051,I857120);
nand I_26140 (I447102,I447085,I857099);
nor I_26141 (I446867,I447102,I447051);
and I_26142 (I446858,I446944,I447102);
not I_26143 (I447147,I447102);
nand I_26144 (I446861,I446944,I447147);
nor I_26145 (I446855,I446910,I447102);
not I_26146 (I447192,I857105);
nor I_26147 (I447209,I447192,I857120);
nand I_26148 (I447226,I447209,I447051);
nor I_26149 (I446864,I446969,I447226);
nor I_26150 (I447257,I447192,I857111);
and I_26151 (I447274,I447257,I857108);
or I_26152 (I447291,I447274,I857114);
DFFARX1 I_26153 (I447291,I2683,I446884,I447317,);
nor I_26154 (I447325,I447317,I447068);
DFFARX1 I_26155 (I447325,I2683,I446884,I446852,);
DFFARX1 I_26156 (I447317,I2683,I446884,I446876,);
not I_26157 (I447370,I447317);
nor I_26158 (I447387,I447370,I446944);
nor I_26159 (I447404,I447209,I447387);
DFFARX1 I_26160 (I447404,I2683,I446884,I446873,);
not I_26161 (I447462,I2690);
DFFARX1 I_26162 (I818119,I2683,I447462,I447488,);
not I_26163 (I447496,I447488);
DFFARX1 I_26164 (I818110,I2683,I447462,I447522,);
not I_26165 (I447530,I818104);
nand I_26166 (I447547,I447530,I818116);
not I_26167 (I447564,I447547);
nor I_26168 (I447581,I447564,I818107);
nor I_26169 (I447598,I447496,I447581);
DFFARX1 I_26170 (I447598,I2683,I447462,I447448,);
not I_26171 (I447629,I818107);
nand I_26172 (I447646,I447629,I447564);
and I_26173 (I447663,I447629,I818113);
nand I_26174 (I447680,I447663,I818098);
nor I_26175 (I447445,I447680,I447629);
and I_26176 (I447436,I447522,I447680);
not I_26177 (I447725,I447680);
nand I_26178 (I447439,I447522,I447725);
nor I_26179 (I447433,I447488,I447680);
not I_26180 (I447770,I818098);
nor I_26181 (I447787,I447770,I818113);
nand I_26182 (I447804,I447787,I447629);
nor I_26183 (I447442,I447547,I447804);
nor I_26184 (I447835,I447770,I818101);
and I_26185 (I447852,I447835,I818104);
or I_26186 (I447869,I447852,I818101);
DFFARX1 I_26187 (I447869,I2683,I447462,I447895,);
nor I_26188 (I447903,I447895,I447646);
DFFARX1 I_26189 (I447903,I2683,I447462,I447430,);
DFFARX1 I_26190 (I447895,I2683,I447462,I447454,);
not I_26191 (I447948,I447895);
nor I_26192 (I447965,I447948,I447522);
nor I_26193 (I447982,I447787,I447965);
DFFARX1 I_26194 (I447982,I2683,I447462,I447451,);
not I_26195 (I448040,I2690);
DFFARX1 I_26196 (I334494,I2683,I448040,I448066,);
not I_26197 (I448074,I448066);
DFFARX1 I_26198 (I334506,I2683,I448040,I448100,);
not I_26199 (I448108,I334482);
nand I_26200 (I448125,I448108,I334509);
not I_26201 (I448142,I448125);
nor I_26202 (I448159,I448142,I334497);
nor I_26203 (I448176,I448074,I448159);
DFFARX1 I_26204 (I448176,I2683,I448040,I448026,);
not I_26205 (I448207,I334497);
nand I_26206 (I448224,I448207,I448142);
and I_26207 (I448241,I448207,I334482);
nand I_26208 (I448258,I448241,I334485);
nor I_26209 (I448023,I448258,I448207);
and I_26210 (I448014,I448100,I448258);
not I_26211 (I448303,I448258);
nand I_26212 (I448017,I448100,I448303);
nor I_26213 (I448011,I448066,I448258);
not I_26214 (I448348,I334491);
nor I_26215 (I448365,I448348,I334482);
nand I_26216 (I448382,I448365,I448207);
nor I_26217 (I448020,I448125,I448382);
nor I_26218 (I448413,I448348,I334500);
and I_26219 (I448430,I448413,I334488);
or I_26220 (I448447,I448430,I334503);
DFFARX1 I_26221 (I448447,I2683,I448040,I448473,);
nor I_26222 (I448481,I448473,I448224);
DFFARX1 I_26223 (I448481,I2683,I448040,I448008,);
DFFARX1 I_26224 (I448473,I2683,I448040,I448032,);
not I_26225 (I448526,I448473);
nor I_26226 (I448543,I448526,I448100);
nor I_26227 (I448560,I448365,I448543);
DFFARX1 I_26228 (I448560,I2683,I448040,I448029,);
not I_26229 (I448618,I2690);
DFFARX1 I_26230 (I153345,I2683,I448618,I448644,);
not I_26231 (I448652,I448644);
DFFARX1 I_26232 (I153330,I2683,I448618,I448678,);
not I_26233 (I448686,I153348);
nand I_26234 (I448703,I448686,I153333);
not I_26235 (I448720,I448703);
nor I_26236 (I448737,I448720,I153330);
nor I_26237 (I448754,I448652,I448737);
DFFARX1 I_26238 (I448754,I2683,I448618,I448604,);
not I_26239 (I448785,I153330);
nand I_26240 (I448802,I448785,I448720);
and I_26241 (I448819,I448785,I153333);
nand I_26242 (I448836,I448819,I153354);
nor I_26243 (I448601,I448836,I448785);
and I_26244 (I448592,I448678,I448836);
not I_26245 (I448881,I448836);
nand I_26246 (I448595,I448678,I448881);
nor I_26247 (I448589,I448644,I448836);
not I_26248 (I448926,I153342);
nor I_26249 (I448943,I448926,I153333);
nand I_26250 (I448960,I448943,I448785);
nor I_26251 (I448598,I448703,I448960);
nor I_26252 (I448991,I448926,I153336);
and I_26253 (I449008,I448991,I153351);
or I_26254 (I449025,I449008,I153339);
DFFARX1 I_26255 (I449025,I2683,I448618,I449051,);
nor I_26256 (I449059,I449051,I448802);
DFFARX1 I_26257 (I449059,I2683,I448618,I448586,);
DFFARX1 I_26258 (I449051,I2683,I448618,I448610,);
not I_26259 (I449104,I449051);
nor I_26260 (I449121,I449104,I448678);
nor I_26261 (I449138,I448943,I449121);
DFFARX1 I_26262 (I449138,I2683,I448618,I448607,);
not I_26263 (I449196,I2690);
DFFARX1 I_26264 (I574012,I2683,I449196,I449222,);
not I_26265 (I449230,I449222);
DFFARX1 I_26266 (I574024,I2683,I449196,I449256,);
not I_26267 (I449264,I574015);
nand I_26268 (I449281,I449264,I574018);
not I_26269 (I449298,I449281);
nor I_26270 (I449315,I449298,I574021);
nor I_26271 (I449332,I449230,I449315);
DFFARX1 I_26272 (I449332,I2683,I449196,I449182,);
not I_26273 (I449363,I574021);
nand I_26274 (I449380,I449363,I449298);
and I_26275 (I449397,I449363,I574015);
nand I_26276 (I449414,I449397,I574027);
nor I_26277 (I449179,I449414,I449363);
and I_26278 (I449170,I449256,I449414);
not I_26279 (I449459,I449414);
nand I_26280 (I449173,I449256,I449459);
nor I_26281 (I449167,I449222,I449414);
not I_26282 (I449504,I574033);
nor I_26283 (I449521,I449504,I574015);
nand I_26284 (I449538,I449521,I449363);
nor I_26285 (I449176,I449281,I449538);
nor I_26286 (I449569,I449504,I574012);
and I_26287 (I449586,I449569,I574030);
or I_26288 (I449603,I449586,I574036);
DFFARX1 I_26289 (I449603,I2683,I449196,I449629,);
nor I_26290 (I449637,I449629,I449380);
DFFARX1 I_26291 (I449637,I2683,I449196,I449164,);
DFFARX1 I_26292 (I449629,I2683,I449196,I449188,);
not I_26293 (I449682,I449629);
nor I_26294 (I449699,I449682,I449256);
nor I_26295 (I449716,I449521,I449699);
DFFARX1 I_26296 (I449716,I2683,I449196,I449185,);
not I_26297 (I449774,I2690);
DFFARX1 I_26298 (I369310,I2683,I449774,I449800,);
not I_26299 (I449808,I449800);
DFFARX1 I_26300 (I369322,I2683,I449774,I449834,);
not I_26301 (I449842,I369298);
nand I_26302 (I449859,I449842,I369325);
not I_26303 (I449876,I449859);
nor I_26304 (I449893,I449876,I369313);
nor I_26305 (I449910,I449808,I449893);
DFFARX1 I_26306 (I449910,I2683,I449774,I449760,);
not I_26307 (I449941,I369313);
nand I_26308 (I449958,I449941,I449876);
and I_26309 (I449975,I449941,I369298);
nand I_26310 (I449992,I449975,I369301);
nor I_26311 (I449757,I449992,I449941);
and I_26312 (I449748,I449834,I449992);
not I_26313 (I450037,I449992);
nand I_26314 (I449751,I449834,I450037);
nor I_26315 (I449745,I449800,I449992);
not I_26316 (I450082,I369307);
nor I_26317 (I450099,I450082,I369298);
nand I_26318 (I450116,I450099,I449941);
nor I_26319 (I449754,I449859,I450116);
nor I_26320 (I450147,I450082,I369316);
and I_26321 (I450164,I450147,I369304);
or I_26322 (I450181,I450164,I369319);
DFFARX1 I_26323 (I450181,I2683,I449774,I450207,);
nor I_26324 (I450215,I450207,I449958);
DFFARX1 I_26325 (I450215,I2683,I449774,I449742,);
DFFARX1 I_26326 (I450207,I2683,I449774,I449766,);
not I_26327 (I450260,I450207);
nor I_26328 (I450277,I450260,I449834);
nor I_26329 (I450294,I450099,I450277);
DFFARX1 I_26330 (I450294,I2683,I449774,I449763,);
not I_26331 (I450352,I2690);
DFFARX1 I_26332 (I1036429,I2683,I450352,I450378,);
not I_26333 (I450386,I450378);
DFFARX1 I_26334 (I1036429,I2683,I450352,I450412,);
not I_26335 (I450420,I1036453);
nand I_26336 (I450437,I450420,I1036435);
not I_26337 (I450454,I450437);
nor I_26338 (I450471,I450454,I1036450);
nor I_26339 (I450488,I450386,I450471);
DFFARX1 I_26340 (I450488,I2683,I450352,I450338,);
not I_26341 (I450519,I1036450);
nand I_26342 (I450536,I450519,I450454);
and I_26343 (I450553,I450519,I1036432);
nand I_26344 (I450570,I450553,I1036441);
nor I_26345 (I450335,I450570,I450519);
and I_26346 (I450326,I450412,I450570);
not I_26347 (I450615,I450570);
nand I_26348 (I450329,I450412,I450615);
nor I_26349 (I450323,I450378,I450570);
not I_26350 (I450660,I1036438);
nor I_26351 (I450677,I450660,I1036432);
nand I_26352 (I450694,I450677,I450519);
nor I_26353 (I450332,I450437,I450694);
nor I_26354 (I450725,I450660,I1036447);
and I_26355 (I450742,I450725,I1036456);
or I_26356 (I450759,I450742,I1036444);
DFFARX1 I_26357 (I450759,I2683,I450352,I450785,);
nor I_26358 (I450793,I450785,I450536);
DFFARX1 I_26359 (I450793,I2683,I450352,I450320,);
DFFARX1 I_26360 (I450785,I2683,I450352,I450344,);
not I_26361 (I450838,I450785);
nor I_26362 (I450855,I450838,I450412);
nor I_26363 (I450872,I450677,I450855);
DFFARX1 I_26364 (I450872,I2683,I450352,I450341,);
not I_26365 (I450930,I2690);
DFFARX1 I_26366 (I511588,I2683,I450930,I450956,);
not I_26367 (I450964,I450956);
DFFARX1 I_26368 (I511600,I2683,I450930,I450990,);
not I_26369 (I450998,I511591);
nand I_26370 (I451015,I450998,I511594);
not I_26371 (I451032,I451015);
nor I_26372 (I451049,I451032,I511597);
nor I_26373 (I451066,I450964,I451049);
DFFARX1 I_26374 (I451066,I2683,I450930,I450916,);
not I_26375 (I451097,I511597);
nand I_26376 (I451114,I451097,I451032);
and I_26377 (I451131,I451097,I511591);
nand I_26378 (I451148,I451131,I511603);
nor I_26379 (I450913,I451148,I451097);
and I_26380 (I450904,I450990,I451148);
not I_26381 (I451193,I451148);
nand I_26382 (I450907,I450990,I451193);
nor I_26383 (I450901,I450956,I451148);
not I_26384 (I451238,I511609);
nor I_26385 (I451255,I451238,I511591);
nand I_26386 (I451272,I451255,I451097);
nor I_26387 (I450910,I451015,I451272);
nor I_26388 (I451303,I451238,I511588);
and I_26389 (I451320,I451303,I511606);
or I_26390 (I451337,I451320,I511612);
DFFARX1 I_26391 (I451337,I2683,I450930,I451363,);
nor I_26392 (I451371,I451363,I451114);
DFFARX1 I_26393 (I451371,I2683,I450930,I450898,);
DFFARX1 I_26394 (I451363,I2683,I450930,I450922,);
not I_26395 (I451416,I451363);
nor I_26396 (I451433,I451416,I450990);
nor I_26397 (I451450,I451255,I451433);
DFFARX1 I_26398 (I451450,I2683,I450930,I450919,);
not I_26399 (I451508,I2690);
DFFARX1 I_26400 (I659154,I2683,I451508,I451534,);
not I_26401 (I451542,I451534);
DFFARX1 I_26402 (I659154,I2683,I451508,I451568,);
not I_26403 (I451576,I659151);
nand I_26404 (I451593,I451576,I659166);
not I_26405 (I451610,I451593);
nor I_26406 (I451627,I451610,I659160);
nor I_26407 (I451644,I451542,I451627);
DFFARX1 I_26408 (I451644,I2683,I451508,I451494,);
not I_26409 (I451675,I659160);
nand I_26410 (I451692,I451675,I451610);
and I_26411 (I451709,I451675,I659157);
nand I_26412 (I451726,I451709,I659148);
nor I_26413 (I451491,I451726,I451675);
and I_26414 (I451482,I451568,I451726);
not I_26415 (I451771,I451726);
nand I_26416 (I451485,I451568,I451771);
nor I_26417 (I451479,I451534,I451726);
not I_26418 (I451816,I659169);
nor I_26419 (I451833,I451816,I659157);
nand I_26420 (I451850,I451833,I451675);
nor I_26421 (I451488,I451593,I451850);
nor I_26422 (I451881,I451816,I659148);
and I_26423 (I451898,I451881,I659151);
or I_26424 (I451915,I451898,I659163);
DFFARX1 I_26425 (I451915,I2683,I451508,I451941,);
nor I_26426 (I451949,I451941,I451692);
DFFARX1 I_26427 (I451949,I2683,I451508,I451476,);
DFFARX1 I_26428 (I451941,I2683,I451508,I451500,);
not I_26429 (I451994,I451941);
nor I_26430 (I452011,I451994,I451568);
nor I_26431 (I452028,I451833,I452011);
DFFARX1 I_26432 (I452028,I2683,I451508,I451497,);
not I_26433 (I452086,I2690);
DFFARX1 I_26434 (I707077,I2683,I452086,I452112,);
not I_26435 (I452120,I452112);
DFFARX1 I_26436 (I707074,I2683,I452086,I452146,);
not I_26437 (I452154,I707071);
nand I_26438 (I452171,I452154,I707098);
not I_26439 (I452188,I452171);
nor I_26440 (I452205,I452188,I707086);
nor I_26441 (I452222,I452120,I452205);
DFFARX1 I_26442 (I452222,I2683,I452086,I452072,);
not I_26443 (I452253,I707086);
nand I_26444 (I452270,I452253,I452188);
and I_26445 (I452287,I452253,I707092);
nand I_26446 (I452304,I452287,I707083);
nor I_26447 (I452069,I452304,I452253);
and I_26448 (I452060,I452146,I452304);
not I_26449 (I452349,I452304);
nand I_26450 (I452063,I452146,I452349);
nor I_26451 (I452057,I452112,I452304);
not I_26452 (I452394,I707080);
nor I_26453 (I452411,I452394,I707092);
nand I_26454 (I452428,I452411,I452253);
nor I_26455 (I452066,I452171,I452428);
nor I_26456 (I452459,I452394,I707095);
and I_26457 (I452476,I452459,I707089);
or I_26458 (I452493,I452476,I707071);
DFFARX1 I_26459 (I452493,I2683,I452086,I452519,);
nor I_26460 (I452527,I452519,I452270);
DFFARX1 I_26461 (I452527,I2683,I452086,I452054,);
DFFARX1 I_26462 (I452519,I2683,I452086,I452078,);
not I_26463 (I452572,I452519);
nor I_26464 (I452589,I452572,I452146);
nor I_26465 (I452606,I452411,I452589);
DFFARX1 I_26466 (I452606,I2683,I452086,I452075,);
not I_26467 (I452664,I2690);
DFFARX1 I_26468 (I635966,I2683,I452664,I452690,);
not I_26469 (I452698,I452690);
DFFARX1 I_26470 (I635966,I2683,I452664,I452724,);
not I_26471 (I452732,I635963);
nand I_26472 (I452749,I452732,I635978);
not I_26473 (I452766,I452749);
nor I_26474 (I452783,I452766,I635972);
nor I_26475 (I452800,I452698,I452783);
DFFARX1 I_26476 (I452800,I2683,I452664,I452650,);
not I_26477 (I452831,I635972);
nand I_26478 (I452848,I452831,I452766);
and I_26479 (I452865,I452831,I635969);
nand I_26480 (I452882,I452865,I635960);
nor I_26481 (I452647,I452882,I452831);
and I_26482 (I452638,I452724,I452882);
not I_26483 (I452927,I452882);
nand I_26484 (I452641,I452724,I452927);
nor I_26485 (I452635,I452690,I452882);
not I_26486 (I452972,I635981);
nor I_26487 (I452989,I452972,I635969);
nand I_26488 (I453006,I452989,I452831);
nor I_26489 (I452644,I452749,I453006);
nor I_26490 (I453037,I452972,I635960);
and I_26491 (I453054,I453037,I635963);
or I_26492 (I453071,I453054,I635975);
DFFARX1 I_26493 (I453071,I2683,I452664,I453097,);
nor I_26494 (I453105,I453097,I452848);
DFFARX1 I_26495 (I453105,I2683,I452664,I452632,);
DFFARX1 I_26496 (I453097,I2683,I452664,I452656,);
not I_26497 (I453150,I453097);
nor I_26498 (I453167,I453150,I452724);
nor I_26499 (I453184,I452989,I453167);
DFFARX1 I_26500 (I453184,I2683,I452664,I452653,);
not I_26501 (I453242,I2690);
DFFARX1 I_26502 (I978800,I2683,I453242,I453268,);
not I_26503 (I453276,I453268);
DFFARX1 I_26504 (I978794,I2683,I453242,I453302,);
not I_26505 (I453310,I978803);
nand I_26506 (I453327,I453310,I978782);
not I_26507 (I453344,I453327);
nor I_26508 (I453361,I453344,I978791);
nor I_26509 (I453378,I453276,I453361);
DFFARX1 I_26510 (I453378,I2683,I453242,I453228,);
not I_26511 (I453409,I978791);
nand I_26512 (I453426,I453409,I453344);
and I_26513 (I453443,I453409,I978806);
nand I_26514 (I453460,I453443,I978785);
nor I_26515 (I453225,I453460,I453409);
and I_26516 (I453216,I453302,I453460);
not I_26517 (I453505,I453460);
nand I_26518 (I453219,I453302,I453505);
nor I_26519 (I453213,I453268,I453460);
not I_26520 (I453550,I978788);
nor I_26521 (I453567,I453550,I978806);
nand I_26522 (I453584,I453567,I453409);
nor I_26523 (I453222,I453327,I453584);
nor I_26524 (I453615,I453550,I978797);
and I_26525 (I453632,I453615,I978785);
or I_26526 (I453649,I453632,I978782);
DFFARX1 I_26527 (I453649,I2683,I453242,I453675,);
nor I_26528 (I453683,I453675,I453426);
DFFARX1 I_26529 (I453683,I2683,I453242,I453210,);
DFFARX1 I_26530 (I453675,I2683,I453242,I453234,);
not I_26531 (I453728,I453675);
nor I_26532 (I453745,I453728,I453302);
nor I_26533 (I453762,I453567,I453745);
DFFARX1 I_26534 (I453762,I2683,I453242,I453231,);
not I_26535 (I453820,I2690);
DFFARX1 I_26536 (I218497,I2683,I453820,I453846,);
not I_26537 (I453854,I453846);
DFFARX1 I_26538 (I218512,I2683,I453820,I453880,);
not I_26539 (I453888,I218515);
nand I_26540 (I453905,I453888,I218494);
not I_26541 (I453922,I453905);
nor I_26542 (I453939,I453922,I218518);
nor I_26543 (I453956,I453854,I453939);
DFFARX1 I_26544 (I453956,I2683,I453820,I453806,);
not I_26545 (I453987,I218518);
nand I_26546 (I454004,I453987,I453922);
and I_26547 (I454021,I453987,I218500);
nand I_26548 (I454038,I454021,I218491);
nor I_26549 (I453803,I454038,I453987);
and I_26550 (I453794,I453880,I454038);
not I_26551 (I454083,I454038);
nand I_26552 (I453797,I453880,I454083);
nor I_26553 (I453791,I453846,I454038);
not I_26554 (I454128,I218491);
nor I_26555 (I454145,I454128,I218500);
nand I_26556 (I454162,I454145,I453987);
nor I_26557 (I453800,I453905,I454162);
nor I_26558 (I454193,I454128,I218506);
and I_26559 (I454210,I454193,I218509);
or I_26560 (I454227,I454210,I218503);
DFFARX1 I_26561 (I454227,I2683,I453820,I454253,);
nor I_26562 (I454261,I454253,I454004);
DFFARX1 I_26563 (I454261,I2683,I453820,I453788,);
DFFARX1 I_26564 (I454253,I2683,I453820,I453812,);
not I_26565 (I454306,I454253);
nor I_26566 (I454323,I454306,I453880);
nor I_26567 (I454340,I454145,I454323);
DFFARX1 I_26568 (I454340,I2683,I453820,I453809,);
not I_26569 (I454398,I2690);
DFFARX1 I_26570 (I963568,I2683,I454398,I454424,);
not I_26571 (I454432,I454424);
DFFARX1 I_26572 (I963562,I2683,I454398,I454458,);
not I_26573 (I454466,I963571);
nand I_26574 (I454483,I454466,I963550);
not I_26575 (I454500,I454483);
nor I_26576 (I454517,I454500,I963559);
nor I_26577 (I454534,I454432,I454517);
DFFARX1 I_26578 (I454534,I2683,I454398,I454384,);
not I_26579 (I454565,I963559);
nand I_26580 (I454582,I454565,I454500);
and I_26581 (I454599,I454565,I963574);
nand I_26582 (I454616,I454599,I963553);
nor I_26583 (I454381,I454616,I454565);
and I_26584 (I454372,I454458,I454616);
not I_26585 (I454661,I454616);
nand I_26586 (I454375,I454458,I454661);
nor I_26587 (I454369,I454424,I454616);
not I_26588 (I454706,I963556);
nor I_26589 (I454723,I454706,I963574);
nand I_26590 (I454740,I454723,I454565);
nor I_26591 (I454378,I454483,I454740);
nor I_26592 (I454771,I454706,I963565);
and I_26593 (I454788,I454771,I963553);
or I_26594 (I454805,I454788,I963550);
DFFARX1 I_26595 (I454805,I2683,I454398,I454831,);
nor I_26596 (I454839,I454831,I454582);
DFFARX1 I_26597 (I454839,I2683,I454398,I454366,);
DFFARX1 I_26598 (I454831,I2683,I454398,I454390,);
not I_26599 (I454884,I454831);
nor I_26600 (I454901,I454884,I454458);
nor I_26601 (I454918,I454723,I454901);
DFFARX1 I_26602 (I454918,I2683,I454398,I454387,);
not I_26603 (I454976,I2690);
DFFARX1 I_26604 (I735501,I2683,I454976,I455002,);
not I_26605 (I455010,I455002);
DFFARX1 I_26606 (I735498,I2683,I454976,I455036,);
not I_26607 (I455044,I735495);
nand I_26608 (I455061,I455044,I735522);
not I_26609 (I455078,I455061);
nor I_26610 (I455095,I455078,I735510);
nor I_26611 (I455112,I455010,I455095);
DFFARX1 I_26612 (I455112,I2683,I454976,I454962,);
not I_26613 (I455143,I735510);
nand I_26614 (I455160,I455143,I455078);
and I_26615 (I455177,I455143,I735516);
nand I_26616 (I455194,I455177,I735507);
nor I_26617 (I454959,I455194,I455143);
and I_26618 (I454950,I455036,I455194);
not I_26619 (I455239,I455194);
nand I_26620 (I454953,I455036,I455239);
nor I_26621 (I454947,I455002,I455194);
not I_26622 (I455284,I735504);
nor I_26623 (I455301,I455284,I735516);
nand I_26624 (I455318,I455301,I455143);
nor I_26625 (I454956,I455061,I455318);
nor I_26626 (I455349,I455284,I735519);
and I_26627 (I455366,I455349,I735513);
or I_26628 (I455383,I455366,I735495);
DFFARX1 I_26629 (I455383,I2683,I454976,I455409,);
nor I_26630 (I455417,I455409,I455160);
DFFARX1 I_26631 (I455417,I2683,I454976,I454944,);
DFFARX1 I_26632 (I455409,I2683,I454976,I454968,);
not I_26633 (I455462,I455409);
nor I_26634 (I455479,I455462,I455036);
nor I_26635 (I455496,I455301,I455479);
DFFARX1 I_26636 (I455496,I2683,I454976,I454965,);
not I_26637 (I455554,I2690);
DFFARX1 I_26638 (I524882,I2683,I455554,I455580,);
not I_26639 (I455588,I455580);
DFFARX1 I_26640 (I524894,I2683,I455554,I455614,);
not I_26641 (I455622,I524885);
nand I_26642 (I455639,I455622,I524888);
not I_26643 (I455656,I455639);
nor I_26644 (I455673,I455656,I524891);
nor I_26645 (I455690,I455588,I455673);
DFFARX1 I_26646 (I455690,I2683,I455554,I455540,);
not I_26647 (I455721,I524891);
nand I_26648 (I455738,I455721,I455656);
and I_26649 (I455755,I455721,I524885);
nand I_26650 (I455772,I455755,I524897);
nor I_26651 (I455537,I455772,I455721);
and I_26652 (I455528,I455614,I455772);
not I_26653 (I455817,I455772);
nand I_26654 (I455531,I455614,I455817);
nor I_26655 (I455525,I455580,I455772);
not I_26656 (I455862,I524903);
nor I_26657 (I455879,I455862,I524885);
nand I_26658 (I455896,I455879,I455721);
nor I_26659 (I455534,I455639,I455896);
nor I_26660 (I455927,I455862,I524882);
and I_26661 (I455944,I455927,I524900);
or I_26662 (I455961,I455944,I524906);
DFFARX1 I_26663 (I455961,I2683,I455554,I455987,);
nor I_26664 (I455995,I455987,I455738);
DFFARX1 I_26665 (I455995,I2683,I455554,I455522,);
DFFARX1 I_26666 (I455987,I2683,I455554,I455546,);
not I_26667 (I456040,I455987);
nor I_26668 (I456057,I456040,I455614);
nor I_26669 (I456074,I455879,I456057);
DFFARX1 I_26670 (I456074,I2683,I455554,I455543,);
not I_26671 (I456132,I2690);
DFFARX1 I_26672 (I1052494,I2683,I456132,I456158,);
not I_26673 (I456166,I456158);
DFFARX1 I_26674 (I1052494,I2683,I456132,I456192,);
not I_26675 (I456200,I1052518);
nand I_26676 (I456217,I456200,I1052500);
not I_26677 (I456234,I456217);
nor I_26678 (I456251,I456234,I1052515);
nor I_26679 (I456268,I456166,I456251);
DFFARX1 I_26680 (I456268,I2683,I456132,I456118,);
not I_26681 (I456299,I1052515);
nand I_26682 (I456316,I456299,I456234);
and I_26683 (I456333,I456299,I1052497);
nand I_26684 (I456350,I456333,I1052506);
nor I_26685 (I456115,I456350,I456299);
and I_26686 (I456106,I456192,I456350);
not I_26687 (I456395,I456350);
nand I_26688 (I456109,I456192,I456395);
nor I_26689 (I456103,I456158,I456350);
not I_26690 (I456440,I1052503);
nor I_26691 (I456457,I456440,I1052497);
nand I_26692 (I456474,I456457,I456299);
nor I_26693 (I456112,I456217,I456474);
nor I_26694 (I456505,I456440,I1052512);
and I_26695 (I456522,I456505,I1052521);
or I_26696 (I456539,I456522,I1052509);
DFFARX1 I_26697 (I456539,I2683,I456132,I456565,);
nor I_26698 (I456573,I456565,I456316);
DFFARX1 I_26699 (I456573,I2683,I456132,I456100,);
DFFARX1 I_26700 (I456565,I2683,I456132,I456124,);
not I_26701 (I456618,I456565);
nor I_26702 (I456635,I456618,I456192);
nor I_26703 (I456652,I456457,I456635);
DFFARX1 I_26704 (I456652,I2683,I456132,I456121,);
not I_26705 (I456710,I2690);
DFFARX1 I_26706 (I372030,I2683,I456710,I456736,);
not I_26707 (I456744,I456736);
DFFARX1 I_26708 (I372042,I2683,I456710,I456770,);
not I_26709 (I456778,I372018);
nand I_26710 (I456795,I456778,I372045);
not I_26711 (I456812,I456795);
nor I_26712 (I456829,I456812,I372033);
nor I_26713 (I456846,I456744,I456829);
DFFARX1 I_26714 (I456846,I2683,I456710,I456696,);
not I_26715 (I456877,I372033);
nand I_26716 (I456894,I456877,I456812);
and I_26717 (I456911,I456877,I372018);
nand I_26718 (I456928,I456911,I372021);
nor I_26719 (I456693,I456928,I456877);
and I_26720 (I456684,I456770,I456928);
not I_26721 (I456973,I456928);
nand I_26722 (I456687,I456770,I456973);
nor I_26723 (I456681,I456736,I456928);
not I_26724 (I457018,I372027);
nor I_26725 (I457035,I457018,I372018);
nand I_26726 (I457052,I457035,I456877);
nor I_26727 (I456690,I456795,I457052);
nor I_26728 (I457083,I457018,I372036);
and I_26729 (I457100,I457083,I372024);
or I_26730 (I457117,I457100,I372039);
DFFARX1 I_26731 (I457117,I2683,I456710,I457143,);
nor I_26732 (I457151,I457143,I456894);
DFFARX1 I_26733 (I457151,I2683,I456710,I456678,);
DFFARX1 I_26734 (I457143,I2683,I456710,I456702,);
not I_26735 (I457196,I457143);
nor I_26736 (I457213,I457196,I456770);
nor I_26737 (I457230,I457035,I457213);
DFFARX1 I_26738 (I457230,I2683,I456710,I456699,);
not I_26739 (I457288,I2690);
DFFARX1 I_26740 (I895244,I2683,I457288,I457314,);
not I_26741 (I457322,I457314);
DFFARX1 I_26742 (I895250,I2683,I457288,I457348,);
not I_26743 (I457356,I895244);
nand I_26744 (I457373,I457356,I895247);
not I_26745 (I457390,I457373);
nor I_26746 (I457407,I457390,I895265);
nor I_26747 (I457424,I457322,I457407);
DFFARX1 I_26748 (I457424,I2683,I457288,I457274,);
not I_26749 (I457455,I895265);
nand I_26750 (I457472,I457455,I457390);
and I_26751 (I457489,I457455,I895268);
nand I_26752 (I457506,I457489,I895247);
nor I_26753 (I457271,I457506,I457455);
and I_26754 (I457262,I457348,I457506);
not I_26755 (I457551,I457506);
nand I_26756 (I457265,I457348,I457551);
nor I_26757 (I457259,I457314,I457506);
not I_26758 (I457596,I895253);
nor I_26759 (I457613,I457596,I895268);
nand I_26760 (I457630,I457613,I457455);
nor I_26761 (I457268,I457373,I457630);
nor I_26762 (I457661,I457596,I895259);
and I_26763 (I457678,I457661,I895256);
or I_26764 (I457695,I457678,I895262);
DFFARX1 I_26765 (I457695,I2683,I457288,I457721,);
nor I_26766 (I457729,I457721,I457472);
DFFARX1 I_26767 (I457729,I2683,I457288,I457256,);
DFFARX1 I_26768 (I457721,I2683,I457288,I457280,);
not I_26769 (I457774,I457721);
nor I_26770 (I457791,I457774,I457348);
nor I_26771 (I457808,I457613,I457791);
DFFARX1 I_26772 (I457808,I2683,I457288,I457277,);
not I_26773 (I457866,I2690);
DFFARX1 I_26774 (I212700,I2683,I457866,I457892,);
not I_26775 (I457900,I457892);
DFFARX1 I_26776 (I212715,I2683,I457866,I457926,);
not I_26777 (I457934,I212718);
nand I_26778 (I457951,I457934,I212697);
not I_26779 (I457968,I457951);
nor I_26780 (I457985,I457968,I212721);
nor I_26781 (I458002,I457900,I457985);
DFFARX1 I_26782 (I458002,I2683,I457866,I457852,);
not I_26783 (I458033,I212721);
nand I_26784 (I458050,I458033,I457968);
and I_26785 (I458067,I458033,I212703);
nand I_26786 (I458084,I458067,I212694);
nor I_26787 (I457849,I458084,I458033);
and I_26788 (I457840,I457926,I458084);
not I_26789 (I458129,I458084);
nand I_26790 (I457843,I457926,I458129);
nor I_26791 (I457837,I457892,I458084);
not I_26792 (I458174,I212694);
nor I_26793 (I458191,I458174,I212703);
nand I_26794 (I458208,I458191,I458033);
nor I_26795 (I457846,I457951,I458208);
nor I_26796 (I458239,I458174,I212709);
and I_26797 (I458256,I458239,I212712);
or I_26798 (I458273,I458256,I212706);
DFFARX1 I_26799 (I458273,I2683,I457866,I458299,);
nor I_26800 (I458307,I458299,I458050);
DFFARX1 I_26801 (I458307,I2683,I457866,I457834,);
DFFARX1 I_26802 (I458299,I2683,I457866,I457858,);
not I_26803 (I458352,I458299);
nor I_26804 (I458369,I458352,I457926);
nor I_26805 (I458386,I458191,I458369);
DFFARX1 I_26806 (I458386,I2683,I457866,I457855,);
not I_26807 (I458444,I2690);
DFFARX1 I_26808 (I873280,I2683,I458444,I458470,);
not I_26809 (I458478,I458470);
DFFARX1 I_26810 (I873286,I2683,I458444,I458504,);
not I_26811 (I458512,I873280);
nand I_26812 (I458529,I458512,I873283);
not I_26813 (I458546,I458529);
nor I_26814 (I458563,I458546,I873301);
nor I_26815 (I458580,I458478,I458563);
DFFARX1 I_26816 (I458580,I2683,I458444,I458430,);
not I_26817 (I458611,I873301);
nand I_26818 (I458628,I458611,I458546);
and I_26819 (I458645,I458611,I873304);
nand I_26820 (I458662,I458645,I873283);
nor I_26821 (I458427,I458662,I458611);
and I_26822 (I458418,I458504,I458662);
not I_26823 (I458707,I458662);
nand I_26824 (I458421,I458504,I458707);
nor I_26825 (I458415,I458470,I458662);
not I_26826 (I458752,I873289);
nor I_26827 (I458769,I458752,I873304);
nand I_26828 (I458786,I458769,I458611);
nor I_26829 (I458424,I458529,I458786);
nor I_26830 (I458817,I458752,I873295);
and I_26831 (I458834,I458817,I873292);
or I_26832 (I458851,I458834,I873298);
DFFARX1 I_26833 (I458851,I2683,I458444,I458877,);
nor I_26834 (I458885,I458877,I458628);
DFFARX1 I_26835 (I458885,I2683,I458444,I458412,);
DFFARX1 I_26836 (I458877,I2683,I458444,I458436,);
not I_26837 (I458930,I458877);
nor I_26838 (I458947,I458930,I458504);
nor I_26839 (I458964,I458769,I458947);
DFFARX1 I_26840 (I458964,I2683,I458444,I458433,);
not I_26841 (I459022,I2690);
DFFARX1 I_26842 (I1010550,I2683,I459022,I459048,);
not I_26843 (I459056,I459048);
DFFARX1 I_26844 (I1010562,I2683,I459022,I459082,);
not I_26845 (I459090,I1010553);
nand I_26846 (I459107,I459090,I1010541);
not I_26847 (I459124,I459107);
nor I_26848 (I459141,I459124,I1010538);
nor I_26849 (I459158,I459056,I459141);
DFFARX1 I_26850 (I459158,I2683,I459022,I459008,);
not I_26851 (I459189,I1010538);
nand I_26852 (I459206,I459189,I459124);
and I_26853 (I459223,I459189,I1010544);
nand I_26854 (I459240,I459223,I1010541);
nor I_26855 (I459005,I459240,I459189);
and I_26856 (I458996,I459082,I459240);
not I_26857 (I459285,I459240);
nand I_26858 (I458999,I459082,I459285);
nor I_26859 (I458993,I459048,I459240);
not I_26860 (I459330,I1010559);
nor I_26861 (I459347,I459330,I1010544);
nand I_26862 (I459364,I459347,I459189);
nor I_26863 (I459002,I459107,I459364);
nor I_26864 (I459395,I459330,I1010547);
and I_26865 (I459412,I459395,I1010538);
or I_26866 (I459429,I459412,I1010556);
DFFARX1 I_26867 (I459429,I2683,I459022,I459455,);
nor I_26868 (I459463,I459455,I459206);
DFFARX1 I_26869 (I459463,I2683,I459022,I458990,);
DFFARX1 I_26870 (I459455,I2683,I459022,I459014,);
not I_26871 (I459508,I459455);
nor I_26872 (I459525,I459508,I459082);
nor I_26873 (I459542,I459347,I459525);
DFFARX1 I_26874 (I459542,I2683,I459022,I459011,);
not I_26875 (I459600,I2690);
DFFARX1 I_26876 (I156915,I2683,I459600,I459626,);
not I_26877 (I459634,I459626);
DFFARX1 I_26878 (I156900,I2683,I459600,I459660,);
not I_26879 (I459668,I156918);
nand I_26880 (I459685,I459668,I156903);
not I_26881 (I459702,I459685);
nor I_26882 (I459719,I459702,I156900);
nor I_26883 (I459736,I459634,I459719);
DFFARX1 I_26884 (I459736,I2683,I459600,I459586,);
not I_26885 (I459767,I156900);
nand I_26886 (I459784,I459767,I459702);
and I_26887 (I459801,I459767,I156903);
nand I_26888 (I459818,I459801,I156924);
nor I_26889 (I459583,I459818,I459767);
and I_26890 (I459574,I459660,I459818);
not I_26891 (I459863,I459818);
nand I_26892 (I459577,I459660,I459863);
nor I_26893 (I459571,I459626,I459818);
not I_26894 (I459908,I156912);
nor I_26895 (I459925,I459908,I156903);
nand I_26896 (I459942,I459925,I459767);
nor I_26897 (I459580,I459685,I459942);
nor I_26898 (I459973,I459908,I156906);
and I_26899 (I459990,I459973,I156921);
or I_26900 (I460007,I459990,I156909);
DFFARX1 I_26901 (I460007,I2683,I459600,I460033,);
nor I_26902 (I460041,I460033,I459784);
DFFARX1 I_26903 (I460041,I2683,I459600,I459568,);
DFFARX1 I_26904 (I460033,I2683,I459600,I459592,);
not I_26905 (I460086,I460033);
nor I_26906 (I460103,I460086,I459660);
nor I_26907 (I460120,I459925,I460103);
DFFARX1 I_26908 (I460120,I2683,I459600,I459589,);
not I_26909 (I460178,I2690);
DFFARX1 I_26910 (I425860,I2683,I460178,I460204,);
not I_26911 (I460212,I460204);
DFFARX1 I_26912 (I425872,I2683,I460178,I460238,);
not I_26913 (I460246,I425878);
nand I_26914 (I460263,I460246,I425869);
not I_26915 (I460280,I460263);
nor I_26916 (I460297,I460280,I425875);
nor I_26917 (I460314,I460212,I460297);
DFFARX1 I_26918 (I460314,I2683,I460178,I460164,);
not I_26919 (I460345,I425875);
nand I_26920 (I460362,I460345,I460280);
and I_26921 (I460379,I460345,I425866);
nand I_26922 (I460396,I460379,I425857);
nor I_26923 (I460161,I460396,I460345);
and I_26924 (I460152,I460238,I460396);
not I_26925 (I460441,I460396);
nand I_26926 (I460155,I460238,I460441);
nor I_26927 (I460149,I460204,I460396);
not I_26928 (I460486,I425863);
nor I_26929 (I460503,I460486,I425866);
nand I_26930 (I460520,I460503,I460345);
nor I_26931 (I460158,I460263,I460520);
nor I_26932 (I460551,I460486,I425860);
and I_26933 (I460568,I460551,I425857);
or I_26934 (I460585,I460568,I425881);
DFFARX1 I_26935 (I460585,I2683,I460178,I460611,);
nor I_26936 (I460619,I460611,I460362);
DFFARX1 I_26937 (I460619,I2683,I460178,I460146,);
DFFARX1 I_26938 (I460611,I2683,I460178,I460170,);
not I_26939 (I460664,I460611);
nor I_26940 (I460681,I460664,I460238);
nor I_26941 (I460698,I460503,I460681);
DFFARX1 I_26942 (I460698,I2683,I460178,I460167,);
not I_26943 (I460756,I2690);
DFFARX1 I_26944 (I884262,I2683,I460756,I460782,);
not I_26945 (I460790,I460782);
DFFARX1 I_26946 (I884268,I2683,I460756,I460816,);
not I_26947 (I460824,I884262);
nand I_26948 (I460841,I460824,I884265);
not I_26949 (I460858,I460841);
nor I_26950 (I460875,I460858,I884283);
nor I_26951 (I460892,I460790,I460875);
DFFARX1 I_26952 (I460892,I2683,I460756,I460742,);
not I_26953 (I460923,I884283);
nand I_26954 (I460940,I460923,I460858);
and I_26955 (I460957,I460923,I884286);
nand I_26956 (I460974,I460957,I884265);
nor I_26957 (I460739,I460974,I460923);
and I_26958 (I460730,I460816,I460974);
not I_26959 (I461019,I460974);
nand I_26960 (I460733,I460816,I461019);
nor I_26961 (I460727,I460782,I460974);
not I_26962 (I461064,I884271);
nor I_26963 (I461081,I461064,I884286);
nand I_26964 (I461098,I461081,I460923);
nor I_26965 (I460736,I460841,I461098);
nor I_26966 (I461129,I461064,I884277);
and I_26967 (I461146,I461129,I884274);
or I_26968 (I461163,I461146,I884280);
DFFARX1 I_26969 (I461163,I2683,I460756,I461189,);
nor I_26970 (I461197,I461189,I460940);
DFFARX1 I_26971 (I461197,I2683,I460756,I460724,);
DFFARX1 I_26972 (I461189,I2683,I460756,I460748,);
not I_26973 (I461242,I461189);
nor I_26974 (I461259,I461242,I460816);
nor I_26975 (I461276,I461081,I461259);
DFFARX1 I_26976 (I461276,I2683,I460756,I460745,);
not I_26977 (I461334,I2690);
DFFARX1 I_26978 (I712245,I2683,I461334,I461360,);
not I_26979 (I461368,I461360);
DFFARX1 I_26980 (I712242,I2683,I461334,I461394,);
not I_26981 (I461402,I712239);
nand I_26982 (I461419,I461402,I712266);
not I_26983 (I461436,I461419);
nor I_26984 (I461453,I461436,I712254);
nor I_26985 (I461470,I461368,I461453);
DFFARX1 I_26986 (I461470,I2683,I461334,I461320,);
not I_26987 (I461501,I712254);
nand I_26988 (I461518,I461501,I461436);
and I_26989 (I461535,I461501,I712260);
nand I_26990 (I461552,I461535,I712251);
nor I_26991 (I461317,I461552,I461501);
and I_26992 (I461308,I461394,I461552);
not I_26993 (I461597,I461552);
nand I_26994 (I461311,I461394,I461597);
nor I_26995 (I461305,I461360,I461552);
not I_26996 (I461642,I712248);
nor I_26997 (I461659,I461642,I712260);
nand I_26998 (I461676,I461659,I461501);
nor I_26999 (I461314,I461419,I461676);
nor I_27000 (I461707,I461642,I712263);
and I_27001 (I461724,I461707,I712257);
or I_27002 (I461741,I461724,I712239);
DFFARX1 I_27003 (I461741,I2683,I461334,I461767,);
nor I_27004 (I461775,I461767,I461518);
DFFARX1 I_27005 (I461775,I2683,I461334,I461302,);
DFFARX1 I_27006 (I461767,I2683,I461334,I461326,);
not I_27007 (I461820,I461767);
nor I_27008 (I461837,I461820,I461394);
nor I_27009 (I461854,I461659,I461837);
DFFARX1 I_27010 (I461854,I2683,I461334,I461323,);
not I_27011 (I461912,I2690);
DFFARX1 I_27012 (I428835,I2683,I461912,I461938,);
not I_27013 (I461946,I461938);
DFFARX1 I_27014 (I428847,I2683,I461912,I461972,);
not I_27015 (I461980,I428853);
nand I_27016 (I461997,I461980,I428844);
not I_27017 (I462014,I461997);
nor I_27018 (I462031,I462014,I428850);
nor I_27019 (I462048,I461946,I462031);
DFFARX1 I_27020 (I462048,I2683,I461912,I461898,);
not I_27021 (I462079,I428850);
nand I_27022 (I462096,I462079,I462014);
and I_27023 (I462113,I462079,I428841);
nand I_27024 (I462130,I462113,I428832);
nor I_27025 (I461895,I462130,I462079);
and I_27026 (I461886,I461972,I462130);
not I_27027 (I462175,I462130);
nand I_27028 (I461889,I461972,I462175);
nor I_27029 (I461883,I461938,I462130);
not I_27030 (I462220,I428838);
nor I_27031 (I462237,I462220,I428841);
nand I_27032 (I462254,I462237,I462079);
nor I_27033 (I461892,I461997,I462254);
nor I_27034 (I462285,I462220,I428835);
and I_27035 (I462302,I462285,I428832);
or I_27036 (I462319,I462302,I428856);
DFFARX1 I_27037 (I462319,I2683,I461912,I462345,);
nor I_27038 (I462353,I462345,I462096);
DFFARX1 I_27039 (I462353,I2683,I461912,I461880,);
DFFARX1 I_27040 (I462345,I2683,I461912,I461904,);
not I_27041 (I462398,I462345);
nor I_27042 (I462415,I462398,I461972);
nor I_27043 (I462432,I462237,I462415);
DFFARX1 I_27044 (I462432,I2683,I461912,I461901,);
not I_27045 (I462490,I2690);
DFFARX1 I_27046 (I1056659,I2683,I462490,I462516,);
not I_27047 (I462524,I462516);
DFFARX1 I_27048 (I1056659,I2683,I462490,I462550,);
not I_27049 (I462558,I1056683);
nand I_27050 (I462575,I462558,I1056665);
not I_27051 (I462592,I462575);
nor I_27052 (I462609,I462592,I1056680);
nor I_27053 (I462626,I462524,I462609);
DFFARX1 I_27054 (I462626,I2683,I462490,I462476,);
not I_27055 (I462657,I1056680);
nand I_27056 (I462674,I462657,I462592);
and I_27057 (I462691,I462657,I1056662);
nand I_27058 (I462708,I462691,I1056671);
nor I_27059 (I462473,I462708,I462657);
and I_27060 (I462464,I462550,I462708);
not I_27061 (I462753,I462708);
nand I_27062 (I462467,I462550,I462753);
nor I_27063 (I462461,I462516,I462708);
not I_27064 (I462798,I1056668);
nor I_27065 (I462815,I462798,I1056662);
nand I_27066 (I462832,I462815,I462657);
nor I_27067 (I462470,I462575,I462832);
nor I_27068 (I462863,I462798,I1056677);
and I_27069 (I462880,I462863,I1056686);
or I_27070 (I462897,I462880,I1056674);
DFFARX1 I_27071 (I462897,I2683,I462490,I462923,);
nor I_27072 (I462931,I462923,I462674);
DFFARX1 I_27073 (I462931,I2683,I462490,I462458,);
DFFARX1 I_27074 (I462923,I2683,I462490,I462482,);
not I_27075 (I462976,I462923);
nor I_27076 (I462993,I462976,I462550);
nor I_27077 (I463010,I462815,I462993);
DFFARX1 I_27078 (I463010,I2683,I462490,I462479,);
not I_27079 (I463068,I2690);
DFFARX1 I_27080 (I19526,I2683,I463068,I463094,);
not I_27081 (I463102,I463094);
DFFARX1 I_27082 (I19529,I2683,I463068,I463128,);
not I_27083 (I463136,I19523);
nand I_27084 (I463153,I463136,I19547);
not I_27085 (I463170,I463153);
nor I_27086 (I463187,I463170,I19526);
nor I_27087 (I463204,I463102,I463187);
DFFARX1 I_27088 (I463204,I2683,I463068,I463054,);
not I_27089 (I463235,I19526);
nand I_27090 (I463252,I463235,I463170);
and I_27091 (I463269,I463235,I19541);
nand I_27092 (I463286,I463269,I19535);
nor I_27093 (I463051,I463286,I463235);
and I_27094 (I463042,I463128,I463286);
not I_27095 (I463331,I463286);
nand I_27096 (I463045,I463128,I463331);
nor I_27097 (I463039,I463094,I463286);
not I_27098 (I463376,I19544);
nor I_27099 (I463393,I463376,I19541);
nand I_27100 (I463410,I463393,I463235);
nor I_27101 (I463048,I463153,I463410);
nor I_27102 (I463441,I463376,I19523);
and I_27103 (I463458,I463441,I19532);
or I_27104 (I463475,I463458,I19538);
DFFARX1 I_27105 (I463475,I2683,I463068,I463501,);
nor I_27106 (I463509,I463501,I463252);
DFFARX1 I_27107 (I463509,I2683,I463068,I463036,);
DFFARX1 I_27108 (I463501,I2683,I463068,I463060,);
not I_27109 (I463554,I463501);
nor I_27110 (I463571,I463554,I463128);
nor I_27111 (I463588,I463393,I463571);
DFFARX1 I_27112 (I463588,I2683,I463068,I463057,);
not I_27113 (I463646,I2690);
DFFARX1 I_27114 (I1047139,I2683,I463646,I463672,);
not I_27115 (I463680,I463672);
DFFARX1 I_27116 (I1047139,I2683,I463646,I463706,);
not I_27117 (I463714,I1047163);
nand I_27118 (I463731,I463714,I1047145);
not I_27119 (I463748,I463731);
nor I_27120 (I463765,I463748,I1047160);
nor I_27121 (I463782,I463680,I463765);
DFFARX1 I_27122 (I463782,I2683,I463646,I463632,);
not I_27123 (I463813,I1047160);
nand I_27124 (I463830,I463813,I463748);
and I_27125 (I463847,I463813,I1047142);
nand I_27126 (I463864,I463847,I1047151);
nor I_27127 (I463629,I463864,I463813);
and I_27128 (I463620,I463706,I463864);
not I_27129 (I463909,I463864);
nand I_27130 (I463623,I463706,I463909);
nor I_27131 (I463617,I463672,I463864);
not I_27132 (I463954,I1047148);
nor I_27133 (I463971,I463954,I1047142);
nand I_27134 (I463988,I463971,I463813);
nor I_27135 (I463626,I463731,I463988);
nor I_27136 (I464019,I463954,I1047157);
and I_27137 (I464036,I464019,I1047166);
or I_27138 (I464053,I464036,I1047154);
DFFARX1 I_27139 (I464053,I2683,I463646,I464079,);
nor I_27140 (I464087,I464079,I463830);
DFFARX1 I_27141 (I464087,I2683,I463646,I463614,);
DFFARX1 I_27142 (I464079,I2683,I463646,I463638,);
not I_27143 (I464132,I464079);
nor I_27144 (I464149,I464132,I463706);
nor I_27145 (I464166,I463971,I464149);
DFFARX1 I_27146 (I464166,I2683,I463646,I463635,);
not I_27147 (I464224,I2690);
DFFARX1 I_27148 (I554360,I2683,I464224,I464250,);
not I_27149 (I464258,I464250);
DFFARX1 I_27150 (I554372,I2683,I464224,I464284,);
not I_27151 (I464292,I554363);
nand I_27152 (I464309,I464292,I554366);
not I_27153 (I464326,I464309);
nor I_27154 (I464343,I464326,I554369);
nor I_27155 (I464360,I464258,I464343);
DFFARX1 I_27156 (I464360,I2683,I464224,I464210,);
not I_27157 (I464391,I554369);
nand I_27158 (I464408,I464391,I464326);
and I_27159 (I464425,I464391,I554363);
nand I_27160 (I464442,I464425,I554375);
nor I_27161 (I464207,I464442,I464391);
and I_27162 (I464198,I464284,I464442);
not I_27163 (I464487,I464442);
nand I_27164 (I464201,I464284,I464487);
nor I_27165 (I464195,I464250,I464442);
not I_27166 (I464532,I554381);
nor I_27167 (I464549,I464532,I554363);
nand I_27168 (I464566,I464549,I464391);
nor I_27169 (I464204,I464309,I464566);
nor I_27170 (I464597,I464532,I554360);
and I_27171 (I464614,I464597,I554378);
or I_27172 (I464631,I464614,I554384);
DFFARX1 I_27173 (I464631,I2683,I464224,I464657,);
nor I_27174 (I464665,I464657,I464408);
DFFARX1 I_27175 (I464665,I2683,I464224,I464192,);
DFFARX1 I_27176 (I464657,I2683,I464224,I464216,);
not I_27177 (I464710,I464657);
nor I_27178 (I464727,I464710,I464284);
nor I_27179 (I464744,I464549,I464727);
DFFARX1 I_27180 (I464744,I2683,I464224,I464213,);
not I_27181 (I464802,I2690);
DFFARX1 I_27182 (I189045,I2683,I464802,I464828,);
not I_27183 (I464836,I464828);
DFFARX1 I_27184 (I189030,I2683,I464802,I464862,);
not I_27185 (I464870,I189048);
nand I_27186 (I464887,I464870,I189033);
not I_27187 (I464904,I464887);
nor I_27188 (I464921,I464904,I189030);
nor I_27189 (I464938,I464836,I464921);
DFFARX1 I_27190 (I464938,I2683,I464802,I464788,);
not I_27191 (I464969,I189030);
nand I_27192 (I464986,I464969,I464904);
and I_27193 (I465003,I464969,I189033);
nand I_27194 (I465020,I465003,I189054);
nor I_27195 (I464785,I465020,I464969);
and I_27196 (I464776,I464862,I465020);
not I_27197 (I465065,I465020);
nand I_27198 (I464779,I464862,I465065);
nor I_27199 (I464773,I464828,I465020);
not I_27200 (I465110,I189042);
nor I_27201 (I465127,I465110,I189033);
nand I_27202 (I465144,I465127,I464969);
nor I_27203 (I464782,I464887,I465144);
nor I_27204 (I465175,I465110,I189036);
and I_27205 (I465192,I465175,I189051);
or I_27206 (I465209,I465192,I189039);
DFFARX1 I_27207 (I465209,I2683,I464802,I465235,);
nor I_27208 (I465243,I465235,I464986);
DFFARX1 I_27209 (I465243,I2683,I464802,I464770,);
DFFARX1 I_27210 (I465235,I2683,I464802,I464794,);
not I_27211 (I465288,I465235);
nor I_27212 (I465305,I465288,I464862);
nor I_27213 (I465322,I465127,I465305);
DFFARX1 I_27214 (I465322,I2683,I464802,I464791,);
not I_27215 (I465380,I2690);
DFFARX1 I_27216 (I1041784,I2683,I465380,I465406,);
not I_27217 (I465414,I465406);
DFFARX1 I_27218 (I1041784,I2683,I465380,I465440,);
not I_27219 (I465448,I1041808);
nand I_27220 (I465465,I465448,I1041790);
not I_27221 (I465482,I465465);
nor I_27222 (I465499,I465482,I1041805);
nor I_27223 (I465516,I465414,I465499);
DFFARX1 I_27224 (I465516,I2683,I465380,I465366,);
not I_27225 (I465547,I1041805);
nand I_27226 (I465564,I465547,I465482);
and I_27227 (I465581,I465547,I1041787);
nand I_27228 (I465598,I465581,I1041796);
nor I_27229 (I465363,I465598,I465547);
and I_27230 (I465354,I465440,I465598);
not I_27231 (I465643,I465598);
nand I_27232 (I465357,I465440,I465643);
nor I_27233 (I465351,I465406,I465598);
not I_27234 (I465688,I1041793);
nor I_27235 (I465705,I465688,I1041787);
nand I_27236 (I465722,I465705,I465547);
nor I_27237 (I465360,I465465,I465722);
nor I_27238 (I465753,I465688,I1041802);
and I_27239 (I465770,I465753,I1041811);
or I_27240 (I465787,I465770,I1041799);
DFFARX1 I_27241 (I465787,I2683,I465380,I465813,);
nor I_27242 (I465821,I465813,I465564);
DFFARX1 I_27243 (I465821,I2683,I465380,I465348,);
DFFARX1 I_27244 (I465813,I2683,I465380,I465372,);
not I_27245 (I465866,I465813);
nor I_27246 (I465883,I465866,I465440);
nor I_27247 (I465900,I465705,I465883);
DFFARX1 I_27248 (I465900,I2683,I465380,I465369,);
not I_27249 (I465958,I2690);
DFFARX1 I_27250 (I590196,I2683,I465958,I465984,);
not I_27251 (I465992,I465984);
DFFARX1 I_27252 (I590208,I2683,I465958,I466018,);
not I_27253 (I466026,I590199);
nand I_27254 (I466043,I466026,I590202);
not I_27255 (I466060,I466043);
nor I_27256 (I466077,I466060,I590205);
nor I_27257 (I466094,I465992,I466077);
DFFARX1 I_27258 (I466094,I2683,I465958,I465944,);
not I_27259 (I466125,I590205);
nand I_27260 (I466142,I466125,I466060);
and I_27261 (I466159,I466125,I590199);
nand I_27262 (I466176,I466159,I590211);
nor I_27263 (I465941,I466176,I466125);
and I_27264 (I465932,I466018,I466176);
not I_27265 (I466221,I466176);
nand I_27266 (I465935,I466018,I466221);
nor I_27267 (I465929,I465984,I466176);
not I_27268 (I466266,I590217);
nor I_27269 (I466283,I466266,I590199);
nand I_27270 (I466300,I466283,I466125);
nor I_27271 (I465938,I466043,I466300);
nor I_27272 (I466331,I466266,I590196);
and I_27273 (I466348,I466331,I590214);
or I_27274 (I466365,I466348,I590220);
DFFARX1 I_27275 (I466365,I2683,I465958,I466391,);
nor I_27276 (I466399,I466391,I466142);
DFFARX1 I_27277 (I466399,I2683,I465958,I465926,);
DFFARX1 I_27278 (I466391,I2683,I465958,I465950,);
not I_27279 (I466444,I466391);
nor I_27280 (I466461,I466444,I466018);
nor I_27281 (I466478,I466283,I466461);
DFFARX1 I_27282 (I466478,I2683,I465958,I465947,);
not I_27283 (I466536,I2690);
DFFARX1 I_27284 (I539332,I2683,I466536,I466562,);
not I_27285 (I466570,I466562);
DFFARX1 I_27286 (I539344,I2683,I466536,I466596,);
not I_27287 (I466604,I539335);
nand I_27288 (I466621,I466604,I539338);
not I_27289 (I466638,I466621);
nor I_27290 (I466655,I466638,I539341);
nor I_27291 (I466672,I466570,I466655);
DFFARX1 I_27292 (I466672,I2683,I466536,I466522,);
not I_27293 (I466703,I539341);
nand I_27294 (I466720,I466703,I466638);
and I_27295 (I466737,I466703,I539335);
nand I_27296 (I466754,I466737,I539347);
nor I_27297 (I466519,I466754,I466703);
and I_27298 (I466510,I466596,I466754);
not I_27299 (I466799,I466754);
nand I_27300 (I466513,I466596,I466799);
nor I_27301 (I466507,I466562,I466754);
not I_27302 (I466844,I539353);
nor I_27303 (I466861,I466844,I539335);
nand I_27304 (I466878,I466861,I466703);
nor I_27305 (I466516,I466621,I466878);
nor I_27306 (I466909,I466844,I539332);
and I_27307 (I466926,I466909,I539350);
or I_27308 (I466943,I466926,I539356);
DFFARX1 I_27309 (I466943,I2683,I466536,I466969,);
nor I_27310 (I466977,I466969,I466720);
DFFARX1 I_27311 (I466977,I2683,I466536,I466504,);
DFFARX1 I_27312 (I466969,I2683,I466536,I466528,);
not I_27313 (I467022,I466969);
nor I_27314 (I467039,I467022,I466596);
nor I_27315 (I467056,I466861,I467039);
DFFARX1 I_27316 (I467056,I2683,I466536,I466525,);
not I_27317 (I467114,I2690);
DFFARX1 I_27318 (I129545,I2683,I467114,I467140,);
not I_27319 (I467148,I467140);
DFFARX1 I_27320 (I129530,I2683,I467114,I467174,);
not I_27321 (I467182,I129548);
nand I_27322 (I467199,I467182,I129533);
not I_27323 (I467216,I467199);
nor I_27324 (I467233,I467216,I129530);
nor I_27325 (I467250,I467148,I467233);
DFFARX1 I_27326 (I467250,I2683,I467114,I467100,);
not I_27327 (I467281,I129530);
nand I_27328 (I467298,I467281,I467216);
and I_27329 (I467315,I467281,I129533);
nand I_27330 (I467332,I467315,I129554);
nor I_27331 (I467097,I467332,I467281);
and I_27332 (I467088,I467174,I467332);
not I_27333 (I467377,I467332);
nand I_27334 (I467091,I467174,I467377);
nor I_27335 (I467085,I467140,I467332);
not I_27336 (I467422,I129542);
nor I_27337 (I467439,I467422,I129533);
nand I_27338 (I467456,I467439,I467281);
nor I_27339 (I467094,I467199,I467456);
nor I_27340 (I467487,I467422,I129536);
and I_27341 (I467504,I467487,I129551);
or I_27342 (I467521,I467504,I129539);
DFFARX1 I_27343 (I467521,I2683,I467114,I467547,);
nor I_27344 (I467555,I467547,I467298);
DFFARX1 I_27345 (I467555,I2683,I467114,I467082,);
DFFARX1 I_27346 (I467547,I2683,I467114,I467106,);
not I_27347 (I467600,I467547);
nor I_27348 (I467617,I467600,I467174);
nor I_27349 (I467634,I467439,I467617);
DFFARX1 I_27350 (I467634,I2683,I467114,I467103,);
not I_27351 (I467692,I2690);
DFFARX1 I_27352 (I177145,I2683,I467692,I467718,);
not I_27353 (I467726,I467718);
DFFARX1 I_27354 (I177130,I2683,I467692,I467752,);
not I_27355 (I467760,I177148);
nand I_27356 (I467777,I467760,I177133);
not I_27357 (I467794,I467777);
nor I_27358 (I467811,I467794,I177130);
nor I_27359 (I467828,I467726,I467811);
DFFARX1 I_27360 (I467828,I2683,I467692,I467678,);
not I_27361 (I467859,I177130);
nand I_27362 (I467876,I467859,I467794);
and I_27363 (I467893,I467859,I177133);
nand I_27364 (I467910,I467893,I177154);
nor I_27365 (I467675,I467910,I467859);
and I_27366 (I467666,I467752,I467910);
not I_27367 (I467955,I467910);
nand I_27368 (I467669,I467752,I467955);
nor I_27369 (I467663,I467718,I467910);
not I_27370 (I468000,I177142);
nor I_27371 (I468017,I468000,I177133);
nand I_27372 (I468034,I468017,I467859);
nor I_27373 (I467672,I467777,I468034);
nor I_27374 (I468065,I468000,I177136);
and I_27375 (I468082,I468065,I177151);
or I_27376 (I468099,I468082,I177139);
DFFARX1 I_27377 (I468099,I2683,I467692,I468125,);
nor I_27378 (I468133,I468125,I467876);
DFFARX1 I_27379 (I468133,I2683,I467692,I467660,);
DFFARX1 I_27380 (I468125,I2683,I467692,I467684,);
not I_27381 (I468178,I468125);
nor I_27382 (I468195,I468178,I467752);
nor I_27383 (I468212,I468017,I468195);
DFFARX1 I_27384 (I468212,I2683,I467692,I467681,);
not I_27385 (I468270,I2690);
DFFARX1 I_27386 (I131925,I2683,I468270,I468296,);
not I_27387 (I468304,I468296);
DFFARX1 I_27388 (I131910,I2683,I468270,I468330,);
not I_27389 (I468338,I131928);
nand I_27390 (I468355,I468338,I131913);
not I_27391 (I468372,I468355);
nor I_27392 (I468389,I468372,I131910);
nor I_27393 (I468406,I468304,I468389);
DFFARX1 I_27394 (I468406,I2683,I468270,I468256,);
not I_27395 (I468437,I131910);
nand I_27396 (I468454,I468437,I468372);
and I_27397 (I468471,I468437,I131913);
nand I_27398 (I468488,I468471,I131934);
nor I_27399 (I468253,I468488,I468437);
and I_27400 (I468244,I468330,I468488);
not I_27401 (I468533,I468488);
nand I_27402 (I468247,I468330,I468533);
nor I_27403 (I468241,I468296,I468488);
not I_27404 (I468578,I131922);
nor I_27405 (I468595,I468578,I131913);
nand I_27406 (I468612,I468595,I468437);
nor I_27407 (I468250,I468355,I468612);
nor I_27408 (I468643,I468578,I131916);
and I_27409 (I468660,I468643,I131931);
or I_27410 (I468677,I468660,I131919);
DFFARX1 I_27411 (I468677,I2683,I468270,I468703,);
nor I_27412 (I468711,I468703,I468454);
DFFARX1 I_27413 (I468711,I2683,I468270,I468238,);
DFFARX1 I_27414 (I468703,I2683,I468270,I468262,);
not I_27415 (I468756,I468703);
nor I_27416 (I468773,I468756,I468330);
nor I_27417 (I468790,I468595,I468773);
DFFARX1 I_27418 (I468790,I2683,I468270,I468259,);
not I_27419 (I468848,I2690);
DFFARX1 I_27420 (I880794,I2683,I468848,I468874,);
not I_27421 (I468882,I468874);
DFFARX1 I_27422 (I880800,I2683,I468848,I468908,);
not I_27423 (I468916,I880794);
nand I_27424 (I468933,I468916,I880797);
not I_27425 (I468950,I468933);
nor I_27426 (I468967,I468950,I880815);
nor I_27427 (I468984,I468882,I468967);
DFFARX1 I_27428 (I468984,I2683,I468848,I468834,);
not I_27429 (I469015,I880815);
nand I_27430 (I469032,I469015,I468950);
and I_27431 (I469049,I469015,I880818);
nand I_27432 (I469066,I469049,I880797);
nor I_27433 (I468831,I469066,I469015);
and I_27434 (I468822,I468908,I469066);
not I_27435 (I469111,I469066);
nand I_27436 (I468825,I468908,I469111);
nor I_27437 (I468819,I468874,I469066);
not I_27438 (I469156,I880803);
nor I_27439 (I469173,I469156,I880818);
nand I_27440 (I469190,I469173,I469015);
nor I_27441 (I468828,I468933,I469190);
nor I_27442 (I469221,I469156,I880809);
and I_27443 (I469238,I469221,I880806);
or I_27444 (I469255,I469238,I880812);
DFFARX1 I_27445 (I469255,I2683,I468848,I469281,);
nor I_27446 (I469289,I469281,I469032);
DFFARX1 I_27447 (I469289,I2683,I468848,I468816,);
DFFARX1 I_27448 (I469281,I2683,I468848,I468840,);
not I_27449 (I469334,I469281);
nor I_27450 (I469351,I469334,I468908);
nor I_27451 (I469368,I469173,I469351);
DFFARX1 I_27452 (I469368,I2683,I468848,I468837,);
not I_27453 (I469426,I2690);
DFFARX1 I_27454 (I318718,I2683,I469426,I469452,);
not I_27455 (I469460,I469452);
DFFARX1 I_27456 (I318730,I2683,I469426,I469486,);
not I_27457 (I469494,I318706);
nand I_27458 (I469511,I469494,I318733);
not I_27459 (I469528,I469511);
nor I_27460 (I469545,I469528,I318721);
nor I_27461 (I469562,I469460,I469545);
DFFARX1 I_27462 (I469562,I2683,I469426,I469412,);
not I_27463 (I469593,I318721);
nand I_27464 (I469610,I469593,I469528);
and I_27465 (I469627,I469593,I318706);
nand I_27466 (I469644,I469627,I318709);
nor I_27467 (I469409,I469644,I469593);
and I_27468 (I469400,I469486,I469644);
not I_27469 (I469689,I469644);
nand I_27470 (I469403,I469486,I469689);
nor I_27471 (I469397,I469452,I469644);
not I_27472 (I469734,I318715);
nor I_27473 (I469751,I469734,I318706);
nand I_27474 (I469768,I469751,I469593);
nor I_27475 (I469406,I469511,I469768);
nor I_27476 (I469799,I469734,I318724);
and I_27477 (I469816,I469799,I318712);
or I_27478 (I469833,I469816,I318727);
DFFARX1 I_27479 (I469833,I2683,I469426,I469859,);
nor I_27480 (I469867,I469859,I469610);
DFFARX1 I_27481 (I469867,I2683,I469426,I469394,);
DFFARX1 I_27482 (I469859,I2683,I469426,I469418,);
not I_27483 (I469912,I469859);
nor I_27484 (I469929,I469912,I469486);
nor I_27485 (I469946,I469751,I469929);
DFFARX1 I_27486 (I469946,I2683,I469426,I469415,);
not I_27487 (I470004,I2690);
DFFARX1 I_27488 (I108610,I2683,I470004,I470030,);
not I_27489 (I470038,I470030);
DFFARX1 I_27490 (I108589,I2683,I470004,I470064,);
not I_27491 (I470072,I108586);
nand I_27492 (I470089,I470072,I108601);
not I_27493 (I470106,I470089);
nor I_27494 (I470123,I470106,I108589);
nor I_27495 (I470140,I470038,I470123);
DFFARX1 I_27496 (I470140,I2683,I470004,I469990,);
not I_27497 (I470171,I108589);
nand I_27498 (I470188,I470171,I470106);
and I_27499 (I470205,I470171,I108592);
nand I_27500 (I470222,I470205,I108607);
nor I_27501 (I469987,I470222,I470171);
and I_27502 (I469978,I470064,I470222);
not I_27503 (I470267,I470222);
nand I_27504 (I469981,I470064,I470267);
nor I_27505 (I469975,I470030,I470222);
not I_27506 (I470312,I108598);
nor I_27507 (I470329,I470312,I108592);
nand I_27508 (I470346,I470329,I470171);
nor I_27509 (I469984,I470089,I470346);
nor I_27510 (I470377,I470312,I108586);
and I_27511 (I470394,I470377,I108595);
or I_27512 (I470411,I470394,I108604);
DFFARX1 I_27513 (I470411,I2683,I470004,I470437,);
nor I_27514 (I470445,I470437,I470188);
DFFARX1 I_27515 (I470445,I2683,I470004,I469972,);
DFFARX1 I_27516 (I470437,I2683,I470004,I469996,);
not I_27517 (I470490,I470437);
nor I_27518 (I470507,I470490,I470064);
nor I_27519 (I470524,I470329,I470507);
DFFARX1 I_27520 (I470524,I2683,I470004,I469993,);
not I_27521 (I470582,I2690);
DFFARX1 I_27522 (I303344,I2683,I470582,I470608,);
not I_27523 (I470616,I470608);
DFFARX1 I_27524 (I303359,I2683,I470582,I470642,);
not I_27525 (I470650,I303362);
nand I_27526 (I470667,I470650,I303341);
not I_27527 (I470684,I470667);
nor I_27528 (I470701,I470684,I303365);
nor I_27529 (I470718,I470616,I470701);
DFFARX1 I_27530 (I470718,I2683,I470582,I470568,);
not I_27531 (I470749,I303365);
nand I_27532 (I470766,I470749,I470684);
and I_27533 (I470783,I470749,I303347);
nand I_27534 (I470800,I470783,I303338);
nor I_27535 (I470565,I470800,I470749);
and I_27536 (I470556,I470642,I470800);
not I_27537 (I470845,I470800);
nand I_27538 (I470559,I470642,I470845);
nor I_27539 (I470553,I470608,I470800);
not I_27540 (I470890,I303338);
nor I_27541 (I470907,I470890,I303347);
nand I_27542 (I470924,I470907,I470749);
nor I_27543 (I470562,I470667,I470924);
nor I_27544 (I470955,I470890,I303353);
and I_27545 (I470972,I470955,I303356);
or I_27546 (I470989,I470972,I303350);
DFFARX1 I_27547 (I470989,I2683,I470582,I471015,);
nor I_27548 (I471023,I471015,I470766);
DFFARX1 I_27549 (I471023,I2683,I470582,I470550,);
DFFARX1 I_27550 (I471015,I2683,I470582,I470574,);
not I_27551 (I471068,I471015);
nor I_27552 (I471085,I471068,I470642);
nor I_27553 (I471102,I470907,I471085);
DFFARX1 I_27554 (I471102,I2683,I470582,I470571,);
not I_27555 (I471160,I2690);
DFFARX1 I_27556 (I245901,I2683,I471160,I471186,);
not I_27557 (I471194,I471186);
DFFARX1 I_27558 (I245916,I2683,I471160,I471220,);
not I_27559 (I471228,I245919);
nand I_27560 (I471245,I471228,I245898);
not I_27561 (I471262,I471245);
nor I_27562 (I471279,I471262,I245922);
nor I_27563 (I471296,I471194,I471279);
DFFARX1 I_27564 (I471296,I2683,I471160,I471146,);
not I_27565 (I471327,I245922);
nand I_27566 (I471344,I471327,I471262);
and I_27567 (I471361,I471327,I245904);
nand I_27568 (I471378,I471361,I245895);
nor I_27569 (I471143,I471378,I471327);
and I_27570 (I471134,I471220,I471378);
not I_27571 (I471423,I471378);
nand I_27572 (I471137,I471220,I471423);
nor I_27573 (I471131,I471186,I471378);
not I_27574 (I471468,I245895);
nor I_27575 (I471485,I471468,I245904);
nand I_27576 (I471502,I471485,I471327);
nor I_27577 (I471140,I471245,I471502);
nor I_27578 (I471533,I471468,I245910);
and I_27579 (I471550,I471533,I245913);
or I_27580 (I471567,I471550,I245907);
DFFARX1 I_27581 (I471567,I2683,I471160,I471593,);
nor I_27582 (I471601,I471593,I471344);
DFFARX1 I_27583 (I471601,I2683,I471160,I471128,);
DFFARX1 I_27584 (I471593,I2683,I471160,I471152,);
not I_27585 (I471646,I471593);
nor I_27586 (I471663,I471646,I471220);
nor I_27587 (I471680,I471485,I471663);
DFFARX1 I_27588 (I471680,I2683,I471160,I471149,);
not I_27589 (I471738,I2690);
DFFARX1 I_27590 (I428240,I2683,I471738,I471764,);
not I_27591 (I471772,I471764);
DFFARX1 I_27592 (I428252,I2683,I471738,I471798,);
not I_27593 (I471806,I428258);
nand I_27594 (I471823,I471806,I428249);
not I_27595 (I471840,I471823);
nor I_27596 (I471857,I471840,I428255);
nor I_27597 (I471874,I471772,I471857);
DFFARX1 I_27598 (I471874,I2683,I471738,I471724,);
not I_27599 (I471905,I428255);
nand I_27600 (I471922,I471905,I471840);
and I_27601 (I471939,I471905,I428246);
nand I_27602 (I471956,I471939,I428237);
nor I_27603 (I471721,I471956,I471905);
and I_27604 (I471712,I471798,I471956);
not I_27605 (I472001,I471956);
nand I_27606 (I471715,I471798,I472001);
nor I_27607 (I471709,I471764,I471956);
not I_27608 (I472046,I428243);
nor I_27609 (I472063,I472046,I428246);
nand I_27610 (I472080,I472063,I471905);
nor I_27611 (I471718,I471823,I472080);
nor I_27612 (I472111,I472046,I428240);
and I_27613 (I472128,I472111,I428237);
or I_27614 (I472145,I472128,I428261);
DFFARX1 I_27615 (I472145,I2683,I471738,I472171,);
nor I_27616 (I472179,I472171,I471922);
DFFARX1 I_27617 (I472179,I2683,I471738,I471706,);
DFFARX1 I_27618 (I472171,I2683,I471738,I471730,);
not I_27619 (I472224,I472171);
nor I_27620 (I472241,I472224,I471798);
nor I_27621 (I472258,I472063,I472241);
DFFARX1 I_27622 (I472258,I2683,I471738,I471727,);
not I_27623 (I472316,I2690);
DFFARX1 I_27624 (I946686,I2683,I472316,I472342,);
not I_27625 (I472350,I472342);
DFFARX1 I_27626 (I946692,I2683,I472316,I472376,);
not I_27627 (I472384,I946686);
nand I_27628 (I472401,I472384,I946689);
not I_27629 (I472418,I472401);
nor I_27630 (I472435,I472418,I946707);
nor I_27631 (I472452,I472350,I472435);
DFFARX1 I_27632 (I472452,I2683,I472316,I472302,);
not I_27633 (I472483,I946707);
nand I_27634 (I472500,I472483,I472418);
and I_27635 (I472517,I472483,I946710);
nand I_27636 (I472534,I472517,I946689);
nor I_27637 (I472299,I472534,I472483);
and I_27638 (I472290,I472376,I472534);
not I_27639 (I472579,I472534);
nand I_27640 (I472293,I472376,I472579);
nor I_27641 (I472287,I472342,I472534);
not I_27642 (I472624,I946695);
nor I_27643 (I472641,I472624,I946710);
nand I_27644 (I472658,I472641,I472483);
nor I_27645 (I472296,I472401,I472658);
nor I_27646 (I472689,I472624,I946701);
and I_27647 (I472706,I472689,I946698);
or I_27648 (I472723,I472706,I946704);
DFFARX1 I_27649 (I472723,I2683,I472316,I472749,);
nor I_27650 (I472757,I472749,I472500);
DFFARX1 I_27651 (I472757,I2683,I472316,I472284,);
DFFARX1 I_27652 (I472749,I2683,I472316,I472308,);
not I_27653 (I472802,I472749);
nor I_27654 (I472819,I472802,I472376);
nor I_27655 (I472836,I472641,I472819);
DFFARX1 I_27656 (I472836,I2683,I472316,I472305,);
not I_27657 (I472894,I2690);
DFFARX1 I_27658 (I353534,I2683,I472894,I472920,);
not I_27659 (I472928,I472920);
DFFARX1 I_27660 (I353546,I2683,I472894,I472954,);
not I_27661 (I472962,I353522);
nand I_27662 (I472979,I472962,I353549);
not I_27663 (I472996,I472979);
nor I_27664 (I473013,I472996,I353537);
nor I_27665 (I473030,I472928,I473013);
DFFARX1 I_27666 (I473030,I2683,I472894,I472880,);
not I_27667 (I473061,I353537);
nand I_27668 (I473078,I473061,I472996);
and I_27669 (I473095,I473061,I353522);
nand I_27670 (I473112,I473095,I353525);
nor I_27671 (I472877,I473112,I473061);
and I_27672 (I472868,I472954,I473112);
not I_27673 (I473157,I473112);
nand I_27674 (I472871,I472954,I473157);
nor I_27675 (I472865,I472920,I473112);
not I_27676 (I473202,I353531);
nor I_27677 (I473219,I473202,I353522);
nand I_27678 (I473236,I473219,I473061);
nor I_27679 (I472874,I472979,I473236);
nor I_27680 (I473267,I473202,I353540);
and I_27681 (I473284,I473267,I353528);
or I_27682 (I473301,I473284,I353543);
DFFARX1 I_27683 (I473301,I2683,I472894,I473327,);
nor I_27684 (I473335,I473327,I473078);
DFFARX1 I_27685 (I473335,I2683,I472894,I472862,);
DFFARX1 I_27686 (I473327,I2683,I472894,I472886,);
not I_27687 (I473380,I473327);
nor I_27688 (I473397,I473380,I472954);
nor I_27689 (I473414,I473219,I473397);
DFFARX1 I_27690 (I473414,I2683,I472894,I472883,);
not I_27691 (I473472,I2690);
DFFARX1 I_27692 (I974448,I2683,I473472,I473498,);
not I_27693 (I473506,I473498);
DFFARX1 I_27694 (I974442,I2683,I473472,I473532,);
not I_27695 (I473540,I974451);
nand I_27696 (I473557,I473540,I974430);
not I_27697 (I473574,I473557);
nor I_27698 (I473591,I473574,I974439);
nor I_27699 (I473608,I473506,I473591);
DFFARX1 I_27700 (I473608,I2683,I473472,I473458,);
not I_27701 (I473639,I974439);
nand I_27702 (I473656,I473639,I473574);
and I_27703 (I473673,I473639,I974454);
nand I_27704 (I473690,I473673,I974433);
nor I_27705 (I473455,I473690,I473639);
and I_27706 (I473446,I473532,I473690);
not I_27707 (I473735,I473690);
nand I_27708 (I473449,I473532,I473735);
nor I_27709 (I473443,I473498,I473690);
not I_27710 (I473780,I974436);
nor I_27711 (I473797,I473780,I974454);
nand I_27712 (I473814,I473797,I473639);
nor I_27713 (I473452,I473557,I473814);
nor I_27714 (I473845,I473780,I974445);
and I_27715 (I473862,I473845,I974433);
or I_27716 (I473879,I473862,I974430);
DFFARX1 I_27717 (I473879,I2683,I473472,I473905,);
nor I_27718 (I473913,I473905,I473656);
DFFARX1 I_27719 (I473913,I2683,I473472,I473440,);
DFFARX1 I_27720 (I473905,I2683,I473472,I473464,);
not I_27721 (I473958,I473905);
nor I_27722 (I473975,I473958,I473532);
nor I_27723 (I473992,I473797,I473975);
DFFARX1 I_27724 (I473992,I2683,I473472,I473461,);
not I_27725 (I474050,I2690);
DFFARX1 I_27726 (I732917,I2683,I474050,I474076,);
not I_27727 (I474084,I474076);
DFFARX1 I_27728 (I732914,I2683,I474050,I474110,);
not I_27729 (I474118,I732911);
nand I_27730 (I474135,I474118,I732938);
not I_27731 (I474152,I474135);
nor I_27732 (I474169,I474152,I732926);
nor I_27733 (I474186,I474084,I474169);
DFFARX1 I_27734 (I474186,I2683,I474050,I474036,);
not I_27735 (I474217,I732926);
nand I_27736 (I474234,I474217,I474152);
and I_27737 (I474251,I474217,I732932);
nand I_27738 (I474268,I474251,I732923);
nor I_27739 (I474033,I474268,I474217);
and I_27740 (I474024,I474110,I474268);
not I_27741 (I474313,I474268);
nand I_27742 (I474027,I474110,I474313);
nor I_27743 (I474021,I474076,I474268);
not I_27744 (I474358,I732920);
nor I_27745 (I474375,I474358,I732932);
nand I_27746 (I474392,I474375,I474217);
nor I_27747 (I474030,I474135,I474392);
nor I_27748 (I474423,I474358,I732935);
and I_27749 (I474440,I474423,I732929);
or I_27750 (I474457,I474440,I732911);
DFFARX1 I_27751 (I474457,I2683,I474050,I474483,);
nor I_27752 (I474491,I474483,I474234);
DFFARX1 I_27753 (I474491,I2683,I474050,I474018,);
DFFARX1 I_27754 (I474483,I2683,I474050,I474042,);
not I_27755 (I474536,I474483);
nor I_27756 (I474553,I474536,I474110);
nor I_27757 (I474570,I474375,I474553);
DFFARX1 I_27758 (I474570,I2683,I474050,I474039,);
not I_27759 (I474628,I2690);
DFFARX1 I_27760 (I261711,I2683,I474628,I474654,);
not I_27761 (I474662,I474654);
DFFARX1 I_27762 (I261726,I2683,I474628,I474688,);
not I_27763 (I474696,I261729);
nand I_27764 (I474713,I474696,I261708);
not I_27765 (I474730,I474713);
nor I_27766 (I474747,I474730,I261732);
nor I_27767 (I474764,I474662,I474747);
DFFARX1 I_27768 (I474764,I2683,I474628,I474614,);
not I_27769 (I474795,I261732);
nand I_27770 (I474812,I474795,I474730);
and I_27771 (I474829,I474795,I261714);
nand I_27772 (I474846,I474829,I261705);
nor I_27773 (I474611,I474846,I474795);
and I_27774 (I474602,I474688,I474846);
not I_27775 (I474891,I474846);
nand I_27776 (I474605,I474688,I474891);
nor I_27777 (I474599,I474654,I474846);
not I_27778 (I474936,I261705);
nor I_27779 (I474953,I474936,I261714);
nand I_27780 (I474970,I474953,I474795);
nor I_27781 (I474608,I474713,I474970);
nor I_27782 (I475001,I474936,I261720);
and I_27783 (I475018,I475001,I261723);
or I_27784 (I475035,I475018,I261717);
DFFARX1 I_27785 (I475035,I2683,I474628,I475061,);
nor I_27786 (I475069,I475061,I474812);
DFFARX1 I_27787 (I475069,I2683,I474628,I474596,);
DFFARX1 I_27788 (I475061,I2683,I474628,I474620,);
not I_27789 (I475114,I475061);
nor I_27790 (I475131,I475114,I474688);
nor I_27791 (I475148,I474953,I475131);
DFFARX1 I_27792 (I475148,I2683,I474628,I474617,);
not I_27793 (I475206,I2690);
DFFARX1 I_27794 (I170005,I2683,I475206,I475232,);
not I_27795 (I475240,I475232);
DFFARX1 I_27796 (I169990,I2683,I475206,I475266,);
not I_27797 (I475274,I170008);
nand I_27798 (I475291,I475274,I169993);
not I_27799 (I475308,I475291);
nor I_27800 (I475325,I475308,I169990);
nor I_27801 (I475342,I475240,I475325);
DFFARX1 I_27802 (I475342,I2683,I475206,I475192,);
not I_27803 (I475373,I169990);
nand I_27804 (I475390,I475373,I475308);
and I_27805 (I475407,I475373,I169993);
nand I_27806 (I475424,I475407,I170014);
nor I_27807 (I475189,I475424,I475373);
and I_27808 (I475180,I475266,I475424);
not I_27809 (I475469,I475424);
nand I_27810 (I475183,I475266,I475469);
nor I_27811 (I475177,I475232,I475424);
not I_27812 (I475514,I170002);
nor I_27813 (I475531,I475514,I169993);
nand I_27814 (I475548,I475531,I475373);
nor I_27815 (I475186,I475291,I475548);
nor I_27816 (I475579,I475514,I169996);
and I_27817 (I475596,I475579,I170011);
or I_27818 (I475613,I475596,I169999);
DFFARX1 I_27819 (I475613,I2683,I475206,I475639,);
nor I_27820 (I475647,I475639,I475390);
DFFARX1 I_27821 (I475647,I2683,I475206,I475174,);
DFFARX1 I_27822 (I475639,I2683,I475206,I475198,);
not I_27823 (I475692,I475639);
nor I_27824 (I475709,I475692,I475266);
nor I_27825 (I475726,I475531,I475709);
DFFARX1 I_27826 (I475726,I2683,I475206,I475195,);
not I_27827 (I475784,I2690);
DFFARX1 I_27828 (I39025,I2683,I475784,I475810,);
not I_27829 (I475818,I475810);
DFFARX1 I_27830 (I39028,I2683,I475784,I475844,);
not I_27831 (I475852,I39022);
nand I_27832 (I475869,I475852,I39046);
not I_27833 (I475886,I475869);
nor I_27834 (I475903,I475886,I39025);
nor I_27835 (I475920,I475818,I475903);
DFFARX1 I_27836 (I475920,I2683,I475784,I475770,);
not I_27837 (I475951,I39025);
nand I_27838 (I475968,I475951,I475886);
and I_27839 (I475985,I475951,I39040);
nand I_27840 (I476002,I475985,I39034);
nor I_27841 (I475767,I476002,I475951);
and I_27842 (I475758,I475844,I476002);
not I_27843 (I476047,I476002);
nand I_27844 (I475761,I475844,I476047);
nor I_27845 (I475755,I475810,I476002);
not I_27846 (I476092,I39043);
nor I_27847 (I476109,I476092,I39040);
nand I_27848 (I476126,I476109,I475951);
nor I_27849 (I475764,I475869,I476126);
nor I_27850 (I476157,I476092,I39022);
and I_27851 (I476174,I476157,I39031);
or I_27852 (I476191,I476174,I39037);
DFFARX1 I_27853 (I476191,I2683,I475784,I476217,);
nor I_27854 (I476225,I476217,I475968);
DFFARX1 I_27855 (I476225,I2683,I475784,I475752,);
DFFARX1 I_27856 (I476217,I2683,I475784,I475776,);
not I_27857 (I476270,I476217);
nor I_27858 (I476287,I476270,I475844);
nor I_27859 (I476304,I476109,I476287);
DFFARX1 I_27860 (I476304,I2683,I475784,I475773,);
not I_27861 (I476362,I2690);
DFFARX1 I_27862 (I1023186,I2683,I476362,I476388,);
not I_27863 (I476396,I476388);
DFFARX1 I_27864 (I1023204,I2683,I476362,I476422,);
not I_27865 (I476430,I1023201);
nand I_27866 (I476447,I476430,I1023192);
not I_27867 (I476464,I476447);
nor I_27868 (I476481,I476464,I1023189);
nor I_27869 (I476498,I476396,I476481);
DFFARX1 I_27870 (I476498,I2683,I476362,I476348,);
not I_27871 (I476529,I1023189);
nand I_27872 (I476546,I476529,I476464);
and I_27873 (I476563,I476529,I1023195);
nand I_27874 (I476580,I476563,I1023210);
nor I_27875 (I476345,I476580,I476529);
and I_27876 (I476336,I476422,I476580);
not I_27877 (I476625,I476580);
nand I_27878 (I476339,I476422,I476625);
nor I_27879 (I476333,I476388,I476580);
not I_27880 (I476670,I1023186);
nor I_27881 (I476687,I476670,I1023195);
nand I_27882 (I476704,I476687,I476529);
nor I_27883 (I476342,I476447,I476704);
nor I_27884 (I476735,I476670,I1023207);
and I_27885 (I476752,I476735,I1023198);
or I_27886 (I476769,I476752,I1023213);
DFFARX1 I_27887 (I476769,I2683,I476362,I476795,);
nor I_27888 (I476803,I476795,I476546);
DFFARX1 I_27889 (I476803,I2683,I476362,I476330,);
DFFARX1 I_27890 (I476795,I2683,I476362,I476354,);
not I_27891 (I476848,I476795);
nor I_27892 (I476865,I476848,I476422);
nor I_27893 (I476882,I476687,I476865);
DFFARX1 I_27894 (I476882,I2683,I476362,I476351,);
not I_27895 (I476940,I2690);
DFFARX1 I_27896 (I138470,I2683,I476940,I476966,);
not I_27897 (I476974,I476966);
DFFARX1 I_27898 (I138455,I2683,I476940,I477000,);
not I_27899 (I477008,I138473);
nand I_27900 (I477025,I477008,I138458);
not I_27901 (I477042,I477025);
nor I_27902 (I477059,I477042,I138455);
nor I_27903 (I477076,I476974,I477059);
DFFARX1 I_27904 (I477076,I2683,I476940,I476926,);
not I_27905 (I477107,I138455);
nand I_27906 (I477124,I477107,I477042);
and I_27907 (I477141,I477107,I138458);
nand I_27908 (I477158,I477141,I138479);
nor I_27909 (I476923,I477158,I477107);
and I_27910 (I476914,I477000,I477158);
not I_27911 (I477203,I477158);
nand I_27912 (I476917,I477000,I477203);
nor I_27913 (I476911,I476966,I477158);
not I_27914 (I477248,I138467);
nor I_27915 (I477265,I477248,I138458);
nand I_27916 (I477282,I477265,I477107);
nor I_27917 (I476920,I477025,I477282);
nor I_27918 (I477313,I477248,I138461);
and I_27919 (I477330,I477313,I138476);
or I_27920 (I477347,I477330,I138464);
DFFARX1 I_27921 (I477347,I2683,I476940,I477373,);
nor I_27922 (I477381,I477373,I477124);
DFFARX1 I_27923 (I477381,I2683,I476940,I476908,);
DFFARX1 I_27924 (I477373,I2683,I476940,I476932,);
not I_27925 (I477426,I477373);
nor I_27926 (I477443,I477426,I477000);
nor I_27927 (I477460,I477265,I477443);
DFFARX1 I_27928 (I477460,I2683,I476940,I476929,);
not I_27929 (I477518,I2690);
DFFARX1 I_27930 (I714183,I2683,I477518,I477544,);
not I_27931 (I477552,I477544);
DFFARX1 I_27932 (I714180,I2683,I477518,I477578,);
not I_27933 (I477586,I714177);
nand I_27934 (I477603,I477586,I714204);
not I_27935 (I477620,I477603);
nor I_27936 (I477637,I477620,I714192);
nor I_27937 (I477654,I477552,I477637);
DFFARX1 I_27938 (I477654,I2683,I477518,I477504,);
not I_27939 (I477685,I714192);
nand I_27940 (I477702,I477685,I477620);
and I_27941 (I477719,I477685,I714198);
nand I_27942 (I477736,I477719,I714189);
nor I_27943 (I477501,I477736,I477685);
and I_27944 (I477492,I477578,I477736);
not I_27945 (I477781,I477736);
nand I_27946 (I477495,I477578,I477781);
nor I_27947 (I477489,I477544,I477736);
not I_27948 (I477826,I714186);
nor I_27949 (I477843,I477826,I714198);
nand I_27950 (I477860,I477843,I477685);
nor I_27951 (I477498,I477603,I477860);
nor I_27952 (I477891,I477826,I714201);
and I_27953 (I477908,I477891,I714195);
or I_27954 (I477925,I477908,I714177);
DFFARX1 I_27955 (I477925,I2683,I477518,I477951,);
nor I_27956 (I477959,I477951,I477702);
DFFARX1 I_27957 (I477959,I2683,I477518,I477486,);
DFFARX1 I_27958 (I477951,I2683,I477518,I477510,);
not I_27959 (I478004,I477951);
nor I_27960 (I478021,I478004,I477578);
nor I_27961 (I478038,I477843,I478021);
DFFARX1 I_27962 (I478038,I2683,I477518,I477507,);
not I_27963 (I478096,I2690);
DFFARX1 I_27964 (I85949,I2683,I478096,I478122,);
not I_27965 (I478130,I478122);
DFFARX1 I_27966 (I85928,I2683,I478096,I478156,);
not I_27967 (I478164,I85925);
nand I_27968 (I478181,I478164,I85940);
not I_27969 (I478198,I478181);
nor I_27970 (I478215,I478198,I85928);
nor I_27971 (I478232,I478130,I478215);
DFFARX1 I_27972 (I478232,I2683,I478096,I478082,);
not I_27973 (I478263,I85928);
nand I_27974 (I478280,I478263,I478198);
and I_27975 (I478297,I478263,I85931);
nand I_27976 (I478314,I478297,I85946);
nor I_27977 (I478079,I478314,I478263);
and I_27978 (I478070,I478156,I478314);
not I_27979 (I478359,I478314);
nand I_27980 (I478073,I478156,I478359);
nor I_27981 (I478067,I478122,I478314);
not I_27982 (I478404,I85937);
nor I_27983 (I478421,I478404,I85931);
nand I_27984 (I478438,I478421,I478263);
nor I_27985 (I478076,I478181,I478438);
nor I_27986 (I478469,I478404,I85925);
and I_27987 (I478486,I478469,I85934);
or I_27988 (I478503,I478486,I85943);
DFFARX1 I_27989 (I478503,I2683,I478096,I478529,);
nor I_27990 (I478537,I478529,I478280);
DFFARX1 I_27991 (I478537,I2683,I478096,I478064,);
DFFARX1 I_27992 (I478529,I2683,I478096,I478088,);
not I_27993 (I478582,I478529);
nor I_27994 (I478599,I478582,I478156);
nor I_27995 (I478616,I478421,I478599);
DFFARX1 I_27996 (I478616,I2683,I478096,I478085,);
not I_27997 (I478674,I2690);
DFFARX1 I_27998 (I602334,I2683,I478674,I478700,);
not I_27999 (I478708,I478700);
DFFARX1 I_28000 (I602346,I2683,I478674,I478734,);
not I_28001 (I478742,I602337);
nand I_28002 (I478759,I478742,I602340);
not I_28003 (I478776,I478759);
nor I_28004 (I478793,I478776,I602343);
nor I_28005 (I478810,I478708,I478793);
DFFARX1 I_28006 (I478810,I2683,I478674,I478660,);
not I_28007 (I478841,I602343);
nand I_28008 (I478858,I478841,I478776);
and I_28009 (I478875,I478841,I602337);
nand I_28010 (I478892,I478875,I602349);
nor I_28011 (I478657,I478892,I478841);
and I_28012 (I478648,I478734,I478892);
not I_28013 (I478937,I478892);
nand I_28014 (I478651,I478734,I478937);
nor I_28015 (I478645,I478700,I478892);
not I_28016 (I478982,I602355);
nor I_28017 (I478999,I478982,I602337);
nand I_28018 (I479016,I478999,I478841);
nor I_28019 (I478654,I478759,I479016);
nor I_28020 (I479047,I478982,I602334);
and I_28021 (I479064,I479047,I602352);
or I_28022 (I479081,I479064,I602358);
DFFARX1 I_28023 (I479081,I2683,I478674,I479107,);
nor I_28024 (I479115,I479107,I478858);
DFFARX1 I_28025 (I479115,I2683,I478674,I478642,);
DFFARX1 I_28026 (I479107,I2683,I478674,I478666,);
not I_28027 (I479160,I479107);
nor I_28028 (I479177,I479160,I478734);
nor I_28029 (I479194,I478999,I479177);
DFFARX1 I_28030 (I479194,I2683,I478674,I478663,);
not I_28031 (I479252,I2690);
DFFARX1 I_28032 (I705139,I2683,I479252,I479278,);
not I_28033 (I479286,I479278);
DFFARX1 I_28034 (I705136,I2683,I479252,I479312,);
not I_28035 (I479320,I705133);
nand I_28036 (I479337,I479320,I705160);
not I_28037 (I479354,I479337);
nor I_28038 (I479371,I479354,I705148);
nor I_28039 (I479388,I479286,I479371);
DFFARX1 I_28040 (I479388,I2683,I479252,I479238,);
not I_28041 (I479419,I705148);
nand I_28042 (I479436,I479419,I479354);
and I_28043 (I479453,I479419,I705154);
nand I_28044 (I479470,I479453,I705145);
nor I_28045 (I479235,I479470,I479419);
and I_28046 (I479226,I479312,I479470);
not I_28047 (I479515,I479470);
nand I_28048 (I479229,I479312,I479515);
nor I_28049 (I479223,I479278,I479470);
not I_28050 (I479560,I705142);
nor I_28051 (I479577,I479560,I705154);
nand I_28052 (I479594,I479577,I479419);
nor I_28053 (I479232,I479337,I479594);
nor I_28054 (I479625,I479560,I705157);
and I_28055 (I479642,I479625,I705151);
or I_28056 (I479659,I479642,I705133);
DFFARX1 I_28057 (I479659,I2683,I479252,I479685,);
nor I_28058 (I479693,I479685,I479436);
DFFARX1 I_28059 (I479693,I2683,I479252,I479220,);
DFFARX1 I_28060 (I479685,I2683,I479252,I479244,);
not I_28061 (I479738,I479685);
nor I_28062 (I479755,I479738,I479312);
nor I_28063 (I479772,I479577,I479755);
DFFARX1 I_28064 (I479772,I2683,I479252,I479241,);
not I_28065 (I479830,I2690);
DFFARX1 I_28066 (I285426,I2683,I479830,I479856,);
not I_28067 (I479864,I479856);
DFFARX1 I_28068 (I285441,I2683,I479830,I479890,);
not I_28069 (I479898,I285444);
nand I_28070 (I479915,I479898,I285423);
not I_28071 (I479932,I479915);
nor I_28072 (I479949,I479932,I285447);
nor I_28073 (I479966,I479864,I479949);
DFFARX1 I_28074 (I479966,I2683,I479830,I479816,);
not I_28075 (I479997,I285447);
nand I_28076 (I480014,I479997,I479932);
and I_28077 (I480031,I479997,I285429);
nand I_28078 (I480048,I480031,I285420);
nor I_28079 (I479813,I480048,I479997);
and I_28080 (I479804,I479890,I480048);
not I_28081 (I480093,I480048);
nand I_28082 (I479807,I479890,I480093);
nor I_28083 (I479801,I479856,I480048);
not I_28084 (I480138,I285420);
nor I_28085 (I480155,I480138,I285429);
nand I_28086 (I480172,I480155,I479997);
nor I_28087 (I479810,I479915,I480172);
nor I_28088 (I480203,I480138,I285435);
and I_28089 (I480220,I480203,I285438);
or I_28090 (I480237,I480220,I285432);
DFFARX1 I_28091 (I480237,I2683,I479830,I480263,);
nor I_28092 (I480271,I480263,I480014);
DFFARX1 I_28093 (I480271,I2683,I479830,I479798,);
DFFARX1 I_28094 (I480263,I2683,I479830,I479822,);
not I_28095 (I480316,I480263);
nor I_28096 (I480333,I480316,I479890);
nor I_28097 (I480350,I480155,I480333);
DFFARX1 I_28098 (I480350,I2683,I479830,I479819,);
not I_28099 (I480408,I2690);
DFFARX1 I_28100 (I1022625,I2683,I480408,I480434,);
not I_28101 (I480442,I480434);
DFFARX1 I_28102 (I1022643,I2683,I480408,I480468,);
not I_28103 (I480476,I1022640);
nand I_28104 (I480493,I480476,I1022631);
not I_28105 (I480510,I480493);
nor I_28106 (I480527,I480510,I1022628);
nor I_28107 (I480544,I480442,I480527);
DFFARX1 I_28108 (I480544,I2683,I480408,I480394,);
not I_28109 (I480575,I1022628);
nand I_28110 (I480592,I480575,I480510);
and I_28111 (I480609,I480575,I1022634);
nand I_28112 (I480626,I480609,I1022649);
nor I_28113 (I480391,I480626,I480575);
and I_28114 (I480382,I480468,I480626);
not I_28115 (I480671,I480626);
nand I_28116 (I480385,I480468,I480671);
nor I_28117 (I480379,I480434,I480626);
not I_28118 (I480716,I1022625);
nor I_28119 (I480733,I480716,I1022634);
nand I_28120 (I480750,I480733,I480575);
nor I_28121 (I480388,I480493,I480750);
nor I_28122 (I480781,I480716,I1022646);
and I_28123 (I480798,I480781,I1022637);
or I_28124 (I480815,I480798,I1022652);
DFFARX1 I_28125 (I480815,I2683,I480408,I480841,);
nor I_28126 (I480849,I480841,I480592);
DFFARX1 I_28127 (I480849,I2683,I480408,I480376,);
DFFARX1 I_28128 (I480841,I2683,I480408,I480400,);
not I_28129 (I480894,I480841);
nor I_28130 (I480911,I480894,I480468);
nor I_28131 (I480928,I480733,I480911);
DFFARX1 I_28132 (I480928,I2683,I480408,I480397,);
not I_28133 (I480986,I2690);
DFFARX1 I_28134 (I222713,I2683,I480986,I481012,);
not I_28135 (I481020,I481012);
DFFARX1 I_28136 (I222728,I2683,I480986,I481046,);
not I_28137 (I481054,I222731);
nand I_28138 (I481071,I481054,I222710);
not I_28139 (I481088,I481071);
nor I_28140 (I481105,I481088,I222734);
nor I_28141 (I481122,I481020,I481105);
DFFARX1 I_28142 (I481122,I2683,I480986,I480972,);
not I_28143 (I481153,I222734);
nand I_28144 (I481170,I481153,I481088);
and I_28145 (I481187,I481153,I222716);
nand I_28146 (I481204,I481187,I222707);
nor I_28147 (I480969,I481204,I481153);
and I_28148 (I480960,I481046,I481204);
not I_28149 (I481249,I481204);
nand I_28150 (I480963,I481046,I481249);
nor I_28151 (I480957,I481012,I481204);
not I_28152 (I481294,I222707);
nor I_28153 (I481311,I481294,I222716);
nand I_28154 (I481328,I481311,I481153);
nor I_28155 (I480966,I481071,I481328);
nor I_28156 (I481359,I481294,I222722);
and I_28157 (I481376,I481359,I222725);
or I_28158 (I481393,I481376,I222719);
DFFARX1 I_28159 (I481393,I2683,I480986,I481419,);
nor I_28160 (I481427,I481419,I481170);
DFFARX1 I_28161 (I481427,I2683,I480986,I480954,);
DFFARX1 I_28162 (I481419,I2683,I480986,I480978,);
not I_28163 (I481472,I481419);
nor I_28164 (I481489,I481472,I481046);
nor I_28165 (I481506,I481311,I481489);
DFFARX1 I_28166 (I481506,I2683,I480986,I480975,);
not I_28167 (I481564,I2690);
DFFARX1 I_28168 (I1073319,I2683,I481564,I481590,);
not I_28169 (I481598,I481590);
DFFARX1 I_28170 (I1073319,I2683,I481564,I481624,);
not I_28171 (I481632,I1073343);
nand I_28172 (I481649,I481632,I1073325);
not I_28173 (I481666,I481649);
nor I_28174 (I481683,I481666,I1073340);
nor I_28175 (I481700,I481598,I481683);
DFFARX1 I_28176 (I481700,I2683,I481564,I481550,);
not I_28177 (I481731,I1073340);
nand I_28178 (I481748,I481731,I481666);
and I_28179 (I481765,I481731,I1073322);
nand I_28180 (I481782,I481765,I1073331);
nor I_28181 (I481547,I481782,I481731);
and I_28182 (I481538,I481624,I481782);
not I_28183 (I481827,I481782);
nand I_28184 (I481541,I481624,I481827);
nor I_28185 (I481535,I481590,I481782);
not I_28186 (I481872,I1073328);
nor I_28187 (I481889,I481872,I1073322);
nand I_28188 (I481906,I481889,I481731);
nor I_28189 (I481544,I481649,I481906);
nor I_28190 (I481937,I481872,I1073337);
and I_28191 (I481954,I481937,I1073346);
or I_28192 (I481971,I481954,I1073334);
DFFARX1 I_28193 (I481971,I2683,I481564,I481997,);
nor I_28194 (I482005,I481997,I481748);
DFFARX1 I_28195 (I482005,I2683,I481564,I481532,);
DFFARX1 I_28196 (I481997,I2683,I481564,I481556,);
not I_28197 (I482050,I481997);
nor I_28198 (I482067,I482050,I481624);
nor I_28199 (I482084,I481889,I482067);
DFFARX1 I_28200 (I482084,I2683,I481564,I481553,);
not I_28201 (I482142,I2690);
DFFARX1 I_28202 (I268562,I2683,I482142,I482168,);
not I_28203 (I482176,I482168);
DFFARX1 I_28204 (I268577,I2683,I482142,I482202,);
not I_28205 (I482210,I268580);
nand I_28206 (I482227,I482210,I268559);
not I_28207 (I482244,I482227);
nor I_28208 (I482261,I482244,I268583);
nor I_28209 (I482278,I482176,I482261);
DFFARX1 I_28210 (I482278,I2683,I482142,I482128,);
not I_28211 (I482309,I268583);
nand I_28212 (I482326,I482309,I482244);
and I_28213 (I482343,I482309,I268565);
nand I_28214 (I482360,I482343,I268556);
nor I_28215 (I482125,I482360,I482309);
and I_28216 (I482116,I482202,I482360);
not I_28217 (I482405,I482360);
nand I_28218 (I482119,I482202,I482405);
nor I_28219 (I482113,I482168,I482360);
not I_28220 (I482450,I268556);
nor I_28221 (I482467,I482450,I268565);
nand I_28222 (I482484,I482467,I482309);
nor I_28223 (I482122,I482227,I482484);
nor I_28224 (I482515,I482450,I268571);
and I_28225 (I482532,I482515,I268574);
or I_28226 (I482549,I482532,I268568);
DFFARX1 I_28227 (I482549,I2683,I482142,I482575,);
nor I_28228 (I482583,I482575,I482326);
DFFARX1 I_28229 (I482583,I2683,I482142,I482110,);
DFFARX1 I_28230 (I482575,I2683,I482142,I482134,);
not I_28231 (I482628,I482575);
nor I_28232 (I482645,I482628,I482202);
nor I_28233 (I482662,I482467,I482645);
DFFARX1 I_28234 (I482662,I2683,I482142,I482131,);
not I_28235 (I482720,I2690);
DFFARX1 I_28236 (I130735,I2683,I482720,I482746,);
not I_28237 (I482754,I482746);
DFFARX1 I_28238 (I130720,I2683,I482720,I482780,);
not I_28239 (I482788,I130738);
nand I_28240 (I482805,I482788,I130723);
not I_28241 (I482822,I482805);
nor I_28242 (I482839,I482822,I130720);
nor I_28243 (I482856,I482754,I482839);
DFFARX1 I_28244 (I482856,I2683,I482720,I482706,);
not I_28245 (I482887,I130720);
nand I_28246 (I482904,I482887,I482822);
and I_28247 (I482921,I482887,I130723);
nand I_28248 (I482938,I482921,I130744);
nor I_28249 (I482703,I482938,I482887);
and I_28250 (I482694,I482780,I482938);
not I_28251 (I482983,I482938);
nand I_28252 (I482697,I482780,I482983);
nor I_28253 (I482691,I482746,I482938);
not I_28254 (I483028,I130732);
nor I_28255 (I483045,I483028,I130723);
nand I_28256 (I483062,I483045,I482887);
nor I_28257 (I482700,I482805,I483062);
nor I_28258 (I483093,I483028,I130726);
and I_28259 (I483110,I483093,I130741);
or I_28260 (I483127,I483110,I130729);
DFFARX1 I_28261 (I483127,I2683,I482720,I483153,);
nor I_28262 (I483161,I483153,I482904);
DFFARX1 I_28263 (I483161,I2683,I482720,I482688,);
DFFARX1 I_28264 (I483153,I2683,I482720,I482712,);
not I_28265 (I483206,I483153);
nor I_28266 (I483223,I483206,I482780);
nor I_28267 (I483240,I483045,I483223);
DFFARX1 I_28268 (I483240,I2683,I482720,I482709,);
not I_28269 (I483298,I2690);
DFFARX1 I_28270 (I516790,I2683,I483298,I483324,);
not I_28271 (I483332,I483324);
DFFARX1 I_28272 (I516802,I2683,I483298,I483358,);
not I_28273 (I483366,I516793);
nand I_28274 (I483383,I483366,I516796);
not I_28275 (I483400,I483383);
nor I_28276 (I483417,I483400,I516799);
nor I_28277 (I483434,I483332,I483417);
DFFARX1 I_28278 (I483434,I2683,I483298,I483284,);
not I_28279 (I483465,I516799);
nand I_28280 (I483482,I483465,I483400);
and I_28281 (I483499,I483465,I516793);
nand I_28282 (I483516,I483499,I516805);
nor I_28283 (I483281,I483516,I483465);
and I_28284 (I483272,I483358,I483516);
not I_28285 (I483561,I483516);
nand I_28286 (I483275,I483358,I483561);
nor I_28287 (I483269,I483324,I483516);
not I_28288 (I483606,I516811);
nor I_28289 (I483623,I483606,I516793);
nand I_28290 (I483640,I483623,I483465);
nor I_28291 (I483278,I483383,I483640);
nor I_28292 (I483671,I483606,I516790);
and I_28293 (I483688,I483671,I516808);
or I_28294 (I483705,I483688,I516814);
DFFARX1 I_28295 (I483705,I2683,I483298,I483731,);
nor I_28296 (I483739,I483731,I483482);
DFFARX1 I_28297 (I483739,I2683,I483298,I483266,);
DFFARX1 I_28298 (I483731,I2683,I483298,I483290,);
not I_28299 (I483784,I483731);
nor I_28300 (I483801,I483784,I483358);
nor I_28301 (I483818,I483623,I483801);
DFFARX1 I_28302 (I483818,I2683,I483298,I483287,);
not I_28303 (I483876,I2690);
DFFARX1 I_28304 (I633331,I2683,I483876,I483902,);
not I_28305 (I483910,I483902);
DFFARX1 I_28306 (I633331,I2683,I483876,I483936,);
not I_28307 (I483944,I633328);
nand I_28308 (I483961,I483944,I633343);
not I_28309 (I483978,I483961);
nor I_28310 (I483995,I483978,I633337);
nor I_28311 (I484012,I483910,I483995);
DFFARX1 I_28312 (I484012,I2683,I483876,I483862,);
not I_28313 (I484043,I633337);
nand I_28314 (I484060,I484043,I483978);
and I_28315 (I484077,I484043,I633334);
nand I_28316 (I484094,I484077,I633325);
nor I_28317 (I483859,I484094,I484043);
and I_28318 (I483850,I483936,I484094);
not I_28319 (I484139,I484094);
nand I_28320 (I483853,I483936,I484139);
nor I_28321 (I483847,I483902,I484094);
not I_28322 (I484184,I633346);
nor I_28323 (I484201,I484184,I633334);
nand I_28324 (I484218,I484201,I484043);
nor I_28325 (I483856,I483961,I484218);
nor I_28326 (I484249,I484184,I633325);
and I_28327 (I484266,I484249,I633328);
or I_28328 (I484283,I484266,I633340);
DFFARX1 I_28329 (I484283,I2683,I483876,I484309,);
nor I_28330 (I484317,I484309,I484060);
DFFARX1 I_28331 (I484317,I2683,I483876,I483844,);
DFFARX1 I_28332 (I484309,I2683,I483876,I483868,);
not I_28333 (I484362,I484309);
nor I_28334 (I484379,I484362,I483936);
nor I_28335 (I484396,I484201,I484379);
DFFARX1 I_28336 (I484396,I2683,I483876,I483865,);
not I_28337 (I484454,I2690);
DFFARX1 I_28338 (I24796,I2683,I484454,I484480,);
not I_28339 (I484488,I484480);
DFFARX1 I_28340 (I24799,I2683,I484454,I484514,);
not I_28341 (I484522,I24793);
nand I_28342 (I484539,I484522,I24817);
not I_28343 (I484556,I484539);
nor I_28344 (I484573,I484556,I24796);
nor I_28345 (I484590,I484488,I484573);
DFFARX1 I_28346 (I484590,I2683,I484454,I484440,);
not I_28347 (I484621,I24796);
nand I_28348 (I484638,I484621,I484556);
and I_28349 (I484655,I484621,I24811);
nand I_28350 (I484672,I484655,I24805);
nor I_28351 (I484437,I484672,I484621);
and I_28352 (I484428,I484514,I484672);
not I_28353 (I484717,I484672);
nand I_28354 (I484431,I484514,I484717);
nor I_28355 (I484425,I484480,I484672);
not I_28356 (I484762,I24814);
nor I_28357 (I484779,I484762,I24811);
nand I_28358 (I484796,I484779,I484621);
nor I_28359 (I484434,I484539,I484796);
nor I_28360 (I484827,I484762,I24793);
and I_28361 (I484844,I484827,I24802);
or I_28362 (I484861,I484844,I24808);
DFFARX1 I_28363 (I484861,I2683,I484454,I484887,);
nor I_28364 (I484895,I484887,I484638);
DFFARX1 I_28365 (I484895,I2683,I484454,I484422,);
DFFARX1 I_28366 (I484887,I2683,I484454,I484446,);
not I_28367 (I484940,I484887);
nor I_28368 (I484957,I484940,I484514);
nor I_28369 (I484974,I484779,I484957);
DFFARX1 I_28370 (I484974,I2683,I484454,I484443,);
not I_28371 (I485032,I2690);
DFFARX1 I_28372 (I989164,I2683,I485032,I485058,);
not I_28373 (I485066,I485058);
DFFARX1 I_28374 (I989176,I2683,I485032,I485092,);
not I_28375 (I485100,I989167);
nand I_28376 (I485117,I485100,I989155);
not I_28377 (I485134,I485117);
nor I_28378 (I485151,I485134,I989152);
nor I_28379 (I485168,I485066,I485151);
DFFARX1 I_28380 (I485168,I2683,I485032,I485018,);
not I_28381 (I485199,I989152);
nand I_28382 (I485216,I485199,I485134);
and I_28383 (I485233,I485199,I989158);
nand I_28384 (I485250,I485233,I989155);
nor I_28385 (I485015,I485250,I485199);
and I_28386 (I485006,I485092,I485250);
not I_28387 (I485295,I485250);
nand I_28388 (I485009,I485092,I485295);
nor I_28389 (I485003,I485058,I485250);
not I_28390 (I485340,I989173);
nor I_28391 (I485357,I485340,I989158);
nand I_28392 (I485374,I485357,I485199);
nor I_28393 (I485012,I485117,I485374);
nor I_28394 (I485405,I485340,I989161);
and I_28395 (I485422,I485405,I989152);
or I_28396 (I485439,I485422,I989170);
DFFARX1 I_28397 (I485439,I2683,I485032,I485465,);
nor I_28398 (I485473,I485465,I485216);
DFFARX1 I_28399 (I485473,I2683,I485032,I485000,);
DFFARX1 I_28400 (I485465,I2683,I485032,I485024,);
not I_28401 (I485518,I485465);
nor I_28402 (I485535,I485518,I485092);
nor I_28403 (I485552,I485357,I485535);
DFFARX1 I_28404 (I485552,I2683,I485032,I485021,);
not I_28405 (I485610,I2690);
DFFARX1 I_28406 (I409795,I2683,I485610,I485636,);
not I_28407 (I485644,I485636);
DFFARX1 I_28408 (I409807,I2683,I485610,I485670,);
not I_28409 (I485678,I409813);
nand I_28410 (I485695,I485678,I409804);
not I_28411 (I485712,I485695);
nor I_28412 (I485729,I485712,I409810);
nor I_28413 (I485746,I485644,I485729);
DFFARX1 I_28414 (I485746,I2683,I485610,I485596,);
not I_28415 (I485777,I409810);
nand I_28416 (I485794,I485777,I485712);
and I_28417 (I485811,I485777,I409801);
nand I_28418 (I485828,I485811,I409792);
nor I_28419 (I485593,I485828,I485777);
and I_28420 (I485584,I485670,I485828);
not I_28421 (I485873,I485828);
nand I_28422 (I485587,I485670,I485873);
nor I_28423 (I485581,I485636,I485828);
not I_28424 (I485918,I409798);
nor I_28425 (I485935,I485918,I409801);
nand I_28426 (I485952,I485935,I485777);
nor I_28427 (I485590,I485695,I485952);
nor I_28428 (I485983,I485918,I409795);
and I_28429 (I486000,I485983,I409792);
or I_28430 (I486017,I486000,I409816);
DFFARX1 I_28431 (I486017,I2683,I485610,I486043,);
nor I_28432 (I486051,I486043,I485794);
DFFARX1 I_28433 (I486051,I2683,I485610,I485578,);
DFFARX1 I_28434 (I486043,I2683,I485610,I485602,);
not I_28435 (I486096,I486043);
nor I_28436 (I486113,I486096,I485670);
nor I_28437 (I486130,I485935,I486113);
DFFARX1 I_28438 (I486130,I2683,I485610,I485599,);
not I_28439 (I486188,I2690);
DFFARX1 I_28440 (I247482,I2683,I486188,I486214,);
not I_28441 (I486222,I486214);
DFFARX1 I_28442 (I247497,I2683,I486188,I486248,);
not I_28443 (I486256,I247500);
nand I_28444 (I486273,I486256,I247479);
not I_28445 (I486290,I486273);
nor I_28446 (I486307,I486290,I247503);
nor I_28447 (I486324,I486222,I486307);
DFFARX1 I_28448 (I486324,I2683,I486188,I486174,);
not I_28449 (I486355,I247503);
nand I_28450 (I486372,I486355,I486290);
and I_28451 (I486389,I486355,I247485);
nand I_28452 (I486406,I486389,I247476);
nor I_28453 (I486171,I486406,I486355);
and I_28454 (I486162,I486248,I486406);
not I_28455 (I486451,I486406);
nand I_28456 (I486165,I486248,I486451);
nor I_28457 (I486159,I486214,I486406);
not I_28458 (I486496,I247476);
nor I_28459 (I486513,I486496,I247485);
nand I_28460 (I486530,I486513,I486355);
nor I_28461 (I486168,I486273,I486530);
nor I_28462 (I486561,I486496,I247491);
and I_28463 (I486578,I486561,I247494);
or I_28464 (I486595,I486578,I247488);
DFFARX1 I_28465 (I486595,I2683,I486188,I486621,);
nor I_28466 (I486629,I486621,I486372);
DFFARX1 I_28467 (I486629,I2683,I486188,I486156,);
DFFARX1 I_28468 (I486621,I2683,I486188,I486180,);
not I_28469 (I486674,I486621);
nor I_28470 (I486691,I486674,I486248);
nor I_28471 (I486708,I486513,I486691);
DFFARX1 I_28472 (I486708,I2683,I486188,I486177,);
not I_28473 (I486766,I2690);
DFFARX1 I_28474 (I156320,I2683,I486766,I486792,);
not I_28475 (I486800,I486792);
DFFARX1 I_28476 (I156305,I2683,I486766,I486826,);
not I_28477 (I486834,I156323);
nand I_28478 (I486851,I486834,I156308);
not I_28479 (I486868,I486851);
nor I_28480 (I486885,I486868,I156305);
nor I_28481 (I486902,I486800,I486885);
DFFARX1 I_28482 (I486902,I2683,I486766,I486752,);
not I_28483 (I486933,I156305);
nand I_28484 (I486950,I486933,I486868);
and I_28485 (I486967,I486933,I156308);
nand I_28486 (I486984,I486967,I156329);
nor I_28487 (I486749,I486984,I486933);
and I_28488 (I486740,I486826,I486984);
not I_28489 (I487029,I486984);
nand I_28490 (I486743,I486826,I487029);
nor I_28491 (I486737,I486792,I486984);
not I_28492 (I487074,I156317);
nor I_28493 (I487091,I487074,I156308);
nand I_28494 (I487108,I487091,I486933);
nor I_28495 (I486746,I486851,I487108);
nor I_28496 (I487139,I487074,I156311);
and I_28497 (I487156,I487139,I156326);
or I_28498 (I487173,I487156,I156314);
DFFARX1 I_28499 (I487173,I2683,I486766,I487199,);
nor I_28500 (I487207,I487199,I486950);
DFFARX1 I_28501 (I487207,I2683,I486766,I486734,);
DFFARX1 I_28502 (I487199,I2683,I486766,I486758,);
not I_28503 (I487252,I487199);
nor I_28504 (I487269,I487252,I486826);
nor I_28505 (I487286,I487091,I487269);
DFFARX1 I_28506 (I487286,I2683,I486766,I486755,);
not I_28507 (I487344,I2690);
DFFARX1 I_28508 (I677072,I2683,I487344,I487370,);
not I_28509 (I487378,I487370);
DFFARX1 I_28510 (I677072,I2683,I487344,I487404,);
not I_28511 (I487412,I677069);
nand I_28512 (I487429,I487412,I677084);
not I_28513 (I487446,I487429);
nor I_28514 (I487463,I487446,I677078);
nor I_28515 (I487480,I487378,I487463);
DFFARX1 I_28516 (I487480,I2683,I487344,I487330,);
not I_28517 (I487511,I677078);
nand I_28518 (I487528,I487511,I487446);
and I_28519 (I487545,I487511,I677075);
nand I_28520 (I487562,I487545,I677066);
nor I_28521 (I487327,I487562,I487511);
and I_28522 (I487318,I487404,I487562);
not I_28523 (I487607,I487562);
nand I_28524 (I487321,I487404,I487607);
nor I_28525 (I487315,I487370,I487562);
not I_28526 (I487652,I677087);
nor I_28527 (I487669,I487652,I677075);
nand I_28528 (I487686,I487669,I487511);
nor I_28529 (I487324,I487429,I487686);
nor I_28530 (I487717,I487652,I677066);
and I_28531 (I487734,I487717,I677069);
or I_28532 (I487751,I487734,I677081);
DFFARX1 I_28533 (I487751,I2683,I487344,I487777,);
nor I_28534 (I487785,I487777,I487528);
DFFARX1 I_28535 (I487785,I2683,I487344,I487312,);
DFFARX1 I_28536 (I487777,I2683,I487344,I487336,);
not I_28537 (I487830,I487777);
nor I_28538 (I487847,I487830,I487404);
nor I_28539 (I487864,I487669,I487847);
DFFARX1 I_28540 (I487864,I2683,I487344,I487333,);
not I_28541 (I487922,I2690);
DFFARX1 I_28542 (I146800,I2683,I487922,I487948,);
not I_28543 (I487956,I487948);
DFFARX1 I_28544 (I146785,I2683,I487922,I487982,);
not I_28545 (I487990,I146803);
nand I_28546 (I488007,I487990,I146788);
not I_28547 (I488024,I488007);
nor I_28548 (I488041,I488024,I146785);
nor I_28549 (I488058,I487956,I488041);
DFFARX1 I_28550 (I488058,I2683,I487922,I487908,);
not I_28551 (I488089,I146785);
nand I_28552 (I488106,I488089,I488024);
and I_28553 (I488123,I488089,I146788);
nand I_28554 (I488140,I488123,I146809);
nor I_28555 (I487905,I488140,I488089);
and I_28556 (I487896,I487982,I488140);
not I_28557 (I488185,I488140);
nand I_28558 (I487899,I487982,I488185);
nor I_28559 (I487893,I487948,I488140);
not I_28560 (I488230,I146797);
nor I_28561 (I488247,I488230,I146788);
nand I_28562 (I488264,I488247,I488089);
nor I_28563 (I487902,I488007,I488264);
nor I_28564 (I488295,I488230,I146791);
and I_28565 (I488312,I488295,I146806);
or I_28566 (I488329,I488312,I146794);
DFFARX1 I_28567 (I488329,I2683,I487922,I488355,);
nor I_28568 (I488363,I488355,I488106);
DFFARX1 I_28569 (I488363,I2683,I487922,I487890,);
DFFARX1 I_28570 (I488355,I2683,I487922,I487914,);
not I_28571 (I488408,I488355);
nor I_28572 (I488425,I488408,I487982);
nor I_28573 (I488442,I488247,I488425);
DFFARX1 I_28574 (I488442,I2683,I487922,I487911,);
not I_28575 (I488500,I2690);
DFFARX1 I_28576 (I57491,I2683,I488500,I488526,);
not I_28577 (I488534,I488526);
DFFARX1 I_28578 (I57470,I2683,I488500,I488560,);
not I_28579 (I488568,I57467);
nand I_28580 (I488585,I488568,I57482);
not I_28581 (I488602,I488585);
nor I_28582 (I488619,I488602,I57470);
nor I_28583 (I488636,I488534,I488619);
DFFARX1 I_28584 (I488636,I2683,I488500,I488486,);
not I_28585 (I488667,I57470);
nand I_28586 (I488684,I488667,I488602);
and I_28587 (I488701,I488667,I57473);
nand I_28588 (I488718,I488701,I57488);
nor I_28589 (I488483,I488718,I488667);
and I_28590 (I488474,I488560,I488718);
not I_28591 (I488763,I488718);
nand I_28592 (I488477,I488560,I488763);
nor I_28593 (I488471,I488526,I488718);
not I_28594 (I488808,I57479);
nor I_28595 (I488825,I488808,I57473);
nand I_28596 (I488842,I488825,I488667);
nor I_28597 (I488480,I488585,I488842);
nor I_28598 (I488873,I488808,I57467);
and I_28599 (I488890,I488873,I57476);
or I_28600 (I488907,I488890,I57485);
DFFARX1 I_28601 (I488907,I2683,I488500,I488933,);
nor I_28602 (I488941,I488933,I488684);
DFFARX1 I_28603 (I488941,I2683,I488500,I488468,);
DFFARX1 I_28604 (I488933,I2683,I488500,I488492,);
not I_28605 (I488986,I488933);
nor I_28606 (I489003,I488986,I488560);
nor I_28607 (I489020,I488825,I489003);
DFFARX1 I_28608 (I489020,I2683,I488500,I488489,);
not I_28609 (I489078,I2690);
DFFARX1 I_28610 (I393246,I2683,I489078,I489104,);
not I_28611 (I489112,I489104);
DFFARX1 I_28612 (I393258,I2683,I489078,I489138,);
not I_28613 (I489146,I393234);
nand I_28614 (I489163,I489146,I393261);
not I_28615 (I489180,I489163);
nor I_28616 (I489197,I489180,I393249);
nor I_28617 (I489214,I489112,I489197);
DFFARX1 I_28618 (I489214,I2683,I489078,I489064,);
not I_28619 (I489245,I393249);
nand I_28620 (I489262,I489245,I489180);
and I_28621 (I489279,I489245,I393234);
nand I_28622 (I489296,I489279,I393237);
nor I_28623 (I489061,I489296,I489245);
and I_28624 (I489052,I489138,I489296);
not I_28625 (I489341,I489296);
nand I_28626 (I489055,I489138,I489341);
nor I_28627 (I489049,I489104,I489296);
not I_28628 (I489386,I393243);
nor I_28629 (I489403,I489386,I393234);
nand I_28630 (I489420,I489403,I489245);
nor I_28631 (I489058,I489163,I489420);
nor I_28632 (I489451,I489386,I393252);
and I_28633 (I489468,I489451,I393240);
or I_28634 (I489485,I489468,I393255);
DFFARX1 I_28635 (I489485,I2683,I489078,I489511,);
nor I_28636 (I489519,I489511,I489262);
DFFARX1 I_28637 (I489519,I2683,I489078,I489046,);
DFFARX1 I_28638 (I489511,I2683,I489078,I489070,);
not I_28639 (I489564,I489511);
nor I_28640 (I489581,I489564,I489138);
nor I_28641 (I489598,I489403,I489581);
DFFARX1 I_28642 (I489598,I2683,I489078,I489067,);
not I_28643 (I489656,I2690);
DFFARX1 I_28644 (I1083434,I2683,I489656,I489682,);
not I_28645 (I489690,I489682);
DFFARX1 I_28646 (I1083434,I2683,I489656,I489716,);
not I_28647 (I489724,I1083458);
nand I_28648 (I489741,I489724,I1083440);
not I_28649 (I489758,I489741);
nor I_28650 (I489775,I489758,I1083455);
nor I_28651 (I489792,I489690,I489775);
DFFARX1 I_28652 (I489792,I2683,I489656,I489642,);
not I_28653 (I489823,I1083455);
nand I_28654 (I489840,I489823,I489758);
and I_28655 (I489857,I489823,I1083437);
nand I_28656 (I489874,I489857,I1083446);
nor I_28657 (I489639,I489874,I489823);
and I_28658 (I489630,I489716,I489874);
not I_28659 (I489919,I489874);
nand I_28660 (I489633,I489716,I489919);
nor I_28661 (I489627,I489682,I489874);
not I_28662 (I489964,I1083443);
nor I_28663 (I489981,I489964,I1083437);
nand I_28664 (I489998,I489981,I489823);
nor I_28665 (I489636,I489741,I489998);
nor I_28666 (I490029,I489964,I1083452);
and I_28667 (I490046,I490029,I1083461);
or I_28668 (I490063,I490046,I1083449);
DFFARX1 I_28669 (I490063,I2683,I489656,I490089,);
nor I_28670 (I490097,I490089,I489840);
DFFARX1 I_28671 (I490097,I2683,I489656,I489624,);
DFFARX1 I_28672 (I490089,I2683,I489656,I489648,);
not I_28673 (I490142,I490089);
nor I_28674 (I490159,I490142,I489716);
nor I_28675 (I490176,I489981,I490159);
DFFARX1 I_28676 (I490176,I2683,I489656,I489645,);
not I_28677 (I490234,I2690);
DFFARX1 I_28678 (I295966,I2683,I490234,I490260,);
not I_28679 (I490268,I490260);
DFFARX1 I_28680 (I295981,I2683,I490234,I490294,);
not I_28681 (I490302,I295984);
nand I_28682 (I490319,I490302,I295963);
not I_28683 (I490336,I490319);
nor I_28684 (I490353,I490336,I295987);
nor I_28685 (I490370,I490268,I490353);
DFFARX1 I_28686 (I490370,I2683,I490234,I490220,);
not I_28687 (I490401,I295987);
nand I_28688 (I490418,I490401,I490336);
and I_28689 (I490435,I490401,I295969);
nand I_28690 (I490452,I490435,I295960);
nor I_28691 (I490217,I490452,I490401);
and I_28692 (I490208,I490294,I490452);
not I_28693 (I490497,I490452);
nand I_28694 (I490211,I490294,I490497);
nor I_28695 (I490205,I490260,I490452);
not I_28696 (I490542,I295960);
nor I_28697 (I490559,I490542,I295969);
nand I_28698 (I490576,I490559,I490401);
nor I_28699 (I490214,I490319,I490576);
nor I_28700 (I490607,I490542,I295975);
and I_28701 (I490624,I490607,I295978);
or I_28702 (I490641,I490624,I295972);
DFFARX1 I_28703 (I490641,I2683,I490234,I490667,);
nor I_28704 (I490675,I490667,I490418);
DFFARX1 I_28705 (I490675,I2683,I490234,I490202,);
DFFARX1 I_28706 (I490667,I2683,I490234,I490226,);
not I_28707 (I490720,I490667);
nor I_28708 (I490737,I490720,I490294);
nor I_28709 (I490754,I490559,I490737);
DFFARX1 I_28710 (I490754,I2683,I490234,I490223,);
not I_28711 (I490812,I2690);
DFFARX1 I_28712 (I1007082,I2683,I490812,I490838,);
not I_28713 (I490846,I490838);
DFFARX1 I_28714 (I1007094,I2683,I490812,I490872,);
not I_28715 (I490880,I1007085);
nand I_28716 (I490897,I490880,I1007073);
not I_28717 (I490914,I490897);
nor I_28718 (I490931,I490914,I1007070);
nor I_28719 (I490948,I490846,I490931);
DFFARX1 I_28720 (I490948,I2683,I490812,I490798,);
not I_28721 (I490979,I1007070);
nand I_28722 (I490996,I490979,I490914);
and I_28723 (I491013,I490979,I1007076);
nand I_28724 (I491030,I491013,I1007073);
nor I_28725 (I490795,I491030,I490979);
and I_28726 (I490786,I490872,I491030);
not I_28727 (I491075,I491030);
nand I_28728 (I490789,I490872,I491075);
nor I_28729 (I490783,I490838,I491030);
not I_28730 (I491120,I1007091);
nor I_28731 (I491137,I491120,I1007076);
nand I_28732 (I491154,I491137,I490979);
nor I_28733 (I490792,I490897,I491154);
nor I_28734 (I491185,I491120,I1007079);
and I_28735 (I491202,I491185,I1007070);
or I_28736 (I491219,I491202,I1007088);
DFFARX1 I_28737 (I491219,I2683,I490812,I491245,);
nor I_28738 (I491253,I491245,I490996);
DFFARX1 I_28739 (I491253,I2683,I490812,I490780,);
DFFARX1 I_28740 (I491245,I2683,I490812,I490804,);
not I_28741 (I491298,I491245);
nor I_28742 (I491315,I491298,I490872);
nor I_28743 (I491332,I491137,I491315);
DFFARX1 I_28744 (I491332,I2683,I490812,I490801,);
not I_28745 (I491390,I2690);
DFFARX1 I_28746 (I548002,I2683,I491390,I491416,);
not I_28747 (I491424,I491416);
DFFARX1 I_28748 (I548014,I2683,I491390,I491450,);
not I_28749 (I491458,I548005);
nand I_28750 (I491475,I491458,I548008);
not I_28751 (I491492,I491475);
nor I_28752 (I491509,I491492,I548011);
nor I_28753 (I491526,I491424,I491509);
DFFARX1 I_28754 (I491526,I2683,I491390,I491376,);
not I_28755 (I491557,I548011);
nand I_28756 (I491574,I491557,I491492);
and I_28757 (I491591,I491557,I548005);
nand I_28758 (I491608,I491591,I548017);
nor I_28759 (I491373,I491608,I491557);
and I_28760 (I491364,I491450,I491608);
not I_28761 (I491653,I491608);
nand I_28762 (I491367,I491450,I491653);
nor I_28763 (I491361,I491416,I491608);
not I_28764 (I491698,I548023);
nor I_28765 (I491715,I491698,I548005);
nand I_28766 (I491732,I491715,I491557);
nor I_28767 (I491370,I491475,I491732);
nor I_28768 (I491763,I491698,I548002);
and I_28769 (I491780,I491763,I548020);
or I_28770 (I491797,I491780,I548026);
DFFARX1 I_28771 (I491797,I2683,I491390,I491823,);
nor I_28772 (I491831,I491823,I491574);
DFFARX1 I_28773 (I491831,I2683,I491390,I491358,);
DFFARX1 I_28774 (I491823,I2683,I491390,I491382,);
not I_28775 (I491876,I491823);
nor I_28776 (I491893,I491876,I491450);
nor I_28777 (I491910,I491715,I491893);
DFFARX1 I_28778 (I491910,I2683,I491390,I491379,);
not I_28779 (I491968,I2690);
DFFARX1 I_28780 (I146205,I2683,I491968,I491994,);
not I_28781 (I492002,I491994);
DFFARX1 I_28782 (I146190,I2683,I491968,I492028,);
not I_28783 (I492036,I146208);
nand I_28784 (I492053,I492036,I146193);
not I_28785 (I492070,I492053);
nor I_28786 (I492087,I492070,I146190);
nor I_28787 (I492104,I492002,I492087);
DFFARX1 I_28788 (I492104,I2683,I491968,I491954,);
not I_28789 (I492135,I146190);
nand I_28790 (I492152,I492135,I492070);
and I_28791 (I492169,I492135,I146193);
nand I_28792 (I492186,I492169,I146214);
nor I_28793 (I491951,I492186,I492135);
and I_28794 (I491942,I492028,I492186);
not I_28795 (I492231,I492186);
nand I_28796 (I491945,I492028,I492231);
nor I_28797 (I491939,I491994,I492186);
not I_28798 (I492276,I146202);
nor I_28799 (I492293,I492276,I146193);
nand I_28800 (I492310,I492293,I492135);
nor I_28801 (I491948,I492053,I492310);
nor I_28802 (I492341,I492276,I146196);
and I_28803 (I492358,I492341,I146211);
or I_28804 (I492375,I492358,I146199);
DFFARX1 I_28805 (I492375,I2683,I491968,I492401,);
nor I_28806 (I492409,I492401,I492152);
DFFARX1 I_28807 (I492409,I2683,I491968,I491936,);
DFFARX1 I_28808 (I492401,I2683,I491968,I491960,);
not I_28809 (I492454,I492401);
nor I_28810 (I492471,I492454,I492028);
nor I_28811 (I492488,I492293,I492471);
DFFARX1 I_28812 (I492488,I2683,I491968,I491957,);
not I_28813 (I492546,I2690);
DFFARX1 I_28814 (I613316,I2683,I492546,I492572,);
not I_28815 (I492580,I492572);
DFFARX1 I_28816 (I613328,I2683,I492546,I492606,);
not I_28817 (I492614,I613319);
nand I_28818 (I492631,I492614,I613322);
not I_28819 (I492648,I492631);
nor I_28820 (I492665,I492648,I613325);
nor I_28821 (I492682,I492580,I492665);
DFFARX1 I_28822 (I492682,I2683,I492546,I492532,);
not I_28823 (I492713,I613325);
nand I_28824 (I492730,I492713,I492648);
and I_28825 (I492747,I492713,I613319);
nand I_28826 (I492764,I492747,I613331);
nor I_28827 (I492529,I492764,I492713);
and I_28828 (I492520,I492606,I492764);
not I_28829 (I492809,I492764);
nand I_28830 (I492523,I492606,I492809);
nor I_28831 (I492517,I492572,I492764);
not I_28832 (I492854,I613337);
nor I_28833 (I492871,I492854,I613319);
nand I_28834 (I492888,I492871,I492713);
nor I_28835 (I492526,I492631,I492888);
nor I_28836 (I492919,I492854,I613316);
and I_28837 (I492936,I492919,I613334);
or I_28838 (I492953,I492936,I613340);
DFFARX1 I_28839 (I492953,I2683,I492546,I492979,);
nor I_28840 (I492987,I492979,I492730);
DFFARX1 I_28841 (I492987,I2683,I492546,I492514,);
DFFARX1 I_28842 (I492979,I2683,I492546,I492538,);
not I_28843 (I493032,I492979);
nor I_28844 (I493049,I493032,I492606);
nor I_28845 (I493066,I492871,I493049);
DFFARX1 I_28846 (I493066,I2683,I492546,I492535,);
not I_28847 (I493124,I2690);
DFFARX1 I_28848 (I117651,I2683,I493124,I493150,);
not I_28849 (I493158,I493150);
DFFARX1 I_28850 (I117630,I2683,I493124,I493184,);
not I_28851 (I493192,I117630);
nand I_28852 (I493209,I493192,I117657);
not I_28853 (I493226,I493209);
nor I_28854 (I493243,I493226,I117633);
nor I_28855 (I493260,I493158,I493243);
DFFARX1 I_28856 (I493260,I2683,I493124,I493110,);
not I_28857 (I493291,I117633);
nand I_28858 (I493308,I493291,I493226);
and I_28859 (I493325,I493291,I117654);
nand I_28860 (I493342,I493325,I117636);
nor I_28861 (I493107,I493342,I493291);
and I_28862 (I493098,I493184,I493342);
not I_28863 (I493387,I493342);
nand I_28864 (I493101,I493184,I493387);
nor I_28865 (I493095,I493150,I493342);
not I_28866 (I493432,I117639);
nor I_28867 (I493449,I493432,I117654);
nand I_28868 (I493466,I493449,I493291);
nor I_28869 (I493104,I493209,I493466);
nor I_28870 (I493497,I493432,I117645);
and I_28871 (I493514,I493497,I117642);
or I_28872 (I493531,I493514,I117648);
DFFARX1 I_28873 (I493531,I2683,I493124,I493557,);
nor I_28874 (I493565,I493557,I493308);
DFFARX1 I_28875 (I493565,I2683,I493124,I493092,);
DFFARX1 I_28876 (I493557,I2683,I493124,I493116,);
not I_28877 (I493610,I493557);
nor I_28878 (I493627,I493610,I493184);
nor I_28879 (I493644,I493449,I493627);
DFFARX1 I_28880 (I493644,I2683,I493124,I493113,);
not I_28881 (I493702,I2690);
DFFARX1 I_28882 (I587884,I2683,I493702,I493728,);
not I_28883 (I493736,I493728);
DFFARX1 I_28884 (I587896,I2683,I493702,I493762,);
not I_28885 (I493770,I587887);
nand I_28886 (I493787,I493770,I587890);
not I_28887 (I493804,I493787);
nor I_28888 (I493821,I493804,I587893);
nor I_28889 (I493838,I493736,I493821);
DFFARX1 I_28890 (I493838,I2683,I493702,I493688,);
not I_28891 (I493869,I587893);
nand I_28892 (I493886,I493869,I493804);
and I_28893 (I493903,I493869,I587887);
nand I_28894 (I493920,I493903,I587899);
nor I_28895 (I493685,I493920,I493869);
and I_28896 (I493676,I493762,I493920);
not I_28897 (I493965,I493920);
nand I_28898 (I493679,I493762,I493965);
nor I_28899 (I493673,I493728,I493920);
not I_28900 (I494010,I587905);
nor I_28901 (I494027,I494010,I587887);
nand I_28902 (I494044,I494027,I493869);
nor I_28903 (I493682,I493787,I494044);
nor I_28904 (I494075,I494010,I587884);
and I_28905 (I494092,I494075,I587902);
or I_28906 (I494109,I494092,I587908);
DFFARX1 I_28907 (I494109,I2683,I493702,I494135,);
nor I_28908 (I494143,I494135,I493886);
DFFARX1 I_28909 (I494143,I2683,I493702,I493670,);
DFFARX1 I_28910 (I494135,I2683,I493702,I493694,);
not I_28911 (I494188,I494135);
nor I_28912 (I494205,I494188,I493762);
nor I_28913 (I494222,I494027,I494205);
DFFARX1 I_28914 (I494222,I2683,I493702,I493691,);
not I_28915 (I494280,I2690);
DFFARX1 I_28916 (I869234,I2683,I494280,I494306,);
not I_28917 (I494314,I494306);
DFFARX1 I_28918 (I869240,I2683,I494280,I494340,);
not I_28919 (I494348,I869234);
nand I_28920 (I494365,I494348,I869237);
not I_28921 (I494382,I494365);
nor I_28922 (I494399,I494382,I869255);
nor I_28923 (I494416,I494314,I494399);
DFFARX1 I_28924 (I494416,I2683,I494280,I494266,);
not I_28925 (I494447,I869255);
nand I_28926 (I494464,I494447,I494382);
and I_28927 (I494481,I494447,I869258);
nand I_28928 (I494498,I494481,I869237);
nor I_28929 (I494263,I494498,I494447);
and I_28930 (I494254,I494340,I494498);
not I_28931 (I494543,I494498);
nand I_28932 (I494257,I494340,I494543);
nor I_28933 (I494251,I494306,I494498);
not I_28934 (I494588,I869243);
nor I_28935 (I494605,I494588,I869258);
nand I_28936 (I494622,I494605,I494447);
nor I_28937 (I494260,I494365,I494622);
nor I_28938 (I494653,I494588,I869249);
and I_28939 (I494670,I494653,I869246);
or I_28940 (I494687,I494670,I869252);
DFFARX1 I_28941 (I494687,I2683,I494280,I494713,);
nor I_28942 (I494721,I494713,I494464);
DFFARX1 I_28943 (I494721,I2683,I494280,I494248,);
DFFARX1 I_28944 (I494713,I2683,I494280,I494272,);
not I_28945 (I494766,I494713);
nor I_28946 (I494783,I494766,I494340);
nor I_28947 (I494800,I494605,I494783);
DFFARX1 I_28948 (I494800,I2683,I494280,I494269,);
not I_28949 (I494858,I2690);
DFFARX1 I_28950 (I799045,I2683,I494858,I494884,);
not I_28951 (I494892,I494884);
DFFARX1 I_28952 (I799036,I2683,I494858,I494918,);
not I_28953 (I494926,I799030);
nand I_28954 (I494943,I494926,I799042);
not I_28955 (I494960,I494943);
nor I_28956 (I494977,I494960,I799033);
nor I_28957 (I494994,I494892,I494977);
DFFARX1 I_28958 (I494994,I2683,I494858,I494844,);
not I_28959 (I495025,I799033);
nand I_28960 (I495042,I495025,I494960);
and I_28961 (I495059,I495025,I799039);
nand I_28962 (I495076,I495059,I799024);
nor I_28963 (I494841,I495076,I495025);
and I_28964 (I494832,I494918,I495076);
not I_28965 (I495121,I495076);
nand I_28966 (I494835,I494918,I495121);
nor I_28967 (I494829,I494884,I495076);
not I_28968 (I495166,I799024);
nor I_28969 (I495183,I495166,I799039);
nand I_28970 (I495200,I495183,I495025);
nor I_28971 (I494838,I494943,I495200);
nor I_28972 (I495231,I495166,I799027);
and I_28973 (I495248,I495231,I799030);
or I_28974 (I495265,I495248,I799027);
DFFARX1 I_28975 (I495265,I2683,I494858,I495291,);
nor I_28976 (I495299,I495291,I495042);
DFFARX1 I_28977 (I495299,I2683,I494858,I494826,);
DFFARX1 I_28978 (I495291,I2683,I494858,I494850,);
not I_28979 (I495344,I495291);
nor I_28980 (I495361,I495344,I494918);
nor I_28981 (I495378,I495183,I495361);
DFFARX1 I_28982 (I495378,I2683,I494858,I494847,);
not I_28983 (I495436,I2690);
DFFARX1 I_28984 (I367134,I2683,I495436,I495462,);
not I_28985 (I495470,I495462);
DFFARX1 I_28986 (I367146,I2683,I495436,I495496,);
not I_28987 (I495504,I367122);
nand I_28988 (I495521,I495504,I367149);
not I_28989 (I495538,I495521);
nor I_28990 (I495555,I495538,I367137);
nor I_28991 (I495572,I495470,I495555);
DFFARX1 I_28992 (I495572,I2683,I495436,I495422,);
not I_28993 (I495603,I367137);
nand I_28994 (I495620,I495603,I495538);
and I_28995 (I495637,I495603,I367122);
nand I_28996 (I495654,I495637,I367125);
nor I_28997 (I495419,I495654,I495603);
and I_28998 (I495410,I495496,I495654);
not I_28999 (I495699,I495654);
nand I_29000 (I495413,I495496,I495699);
nor I_29001 (I495407,I495462,I495654);
not I_29002 (I495744,I367131);
nor I_29003 (I495761,I495744,I367122);
nand I_29004 (I495778,I495761,I495603);
nor I_29005 (I495416,I495521,I495778);
nor I_29006 (I495809,I495744,I367140);
and I_29007 (I495826,I495809,I367128);
or I_29008 (I495843,I495826,I367143);
DFFARX1 I_29009 (I495843,I2683,I495436,I495869,);
nor I_29010 (I495877,I495869,I495620);
DFFARX1 I_29011 (I495877,I2683,I495436,I495404,);
DFFARX1 I_29012 (I495869,I2683,I495436,I495428,);
not I_29013 (I495922,I495869);
nor I_29014 (I495939,I495922,I495496);
nor I_29015 (I495956,I495761,I495939);
DFFARX1 I_29016 (I495956,I2683,I495436,I495425,);
not I_29017 (I496014,I2690);
DFFARX1 I_29018 (I200945,I2683,I496014,I496040,);
not I_29019 (I496048,I496040);
DFFARX1 I_29020 (I200930,I2683,I496014,I496074,);
not I_29021 (I496082,I200948);
nand I_29022 (I496099,I496082,I200933);
not I_29023 (I496116,I496099);
nor I_29024 (I496133,I496116,I200930);
nor I_29025 (I496150,I496048,I496133);
DFFARX1 I_29026 (I496150,I2683,I496014,I496000,);
not I_29027 (I496181,I200930);
nand I_29028 (I496198,I496181,I496116);
and I_29029 (I496215,I496181,I200933);
nand I_29030 (I496232,I496215,I200954);
nor I_29031 (I495997,I496232,I496181);
and I_29032 (I495988,I496074,I496232);
not I_29033 (I496277,I496232);
nand I_29034 (I495991,I496074,I496277);
nor I_29035 (I495985,I496040,I496232);
not I_29036 (I496322,I200942);
nor I_29037 (I496339,I496322,I200933);
nand I_29038 (I496356,I496339,I496181);
nor I_29039 (I495994,I496099,I496356);
nor I_29040 (I496387,I496322,I200936);
and I_29041 (I496404,I496387,I200951);
or I_29042 (I496421,I496404,I200939);
DFFARX1 I_29043 (I496421,I2683,I496014,I496447,);
nor I_29044 (I496455,I496447,I496198);
DFFARX1 I_29045 (I496455,I2683,I496014,I495982,);
DFFARX1 I_29046 (I496447,I2683,I496014,I496006,);
not I_29047 (I496500,I496447);
nor I_29048 (I496517,I496500,I496074);
nor I_29049 (I496534,I496339,I496517);
DFFARX1 I_29050 (I496534,I2683,I496014,I496003,);
not I_29051 (I496592,I2690);
DFFARX1 I_29052 (I892372,I2683,I496592,I496618,);
not I_29053 (I496626,I496618);
nand I_29054 (I496643,I892354,I892366);
and I_29055 (I496660,I496643,I892369);
DFFARX1 I_29056 (I496660,I2683,I496592,I496686,);
not I_29057 (I496694,I892363);
DFFARX1 I_29058 (I892360,I2683,I496592,I496720,);
not I_29059 (I496728,I496720);
nor I_29060 (I496745,I496728,I496626);
and I_29061 (I496762,I496745,I892363);
nor I_29062 (I496779,I496728,I496694);
nor I_29063 (I496575,I496686,I496779);
DFFARX1 I_29064 (I892378,I2683,I496592,I496819,);
nor I_29065 (I496827,I496819,I496686);
not I_29066 (I496844,I496827);
not I_29067 (I496861,I496819);
nor I_29068 (I496878,I496861,I496762);
DFFARX1 I_29069 (I496878,I2683,I496592,I496578,);
nand I_29070 (I496909,I892357,I892357);
and I_29071 (I496926,I496909,I892354);
DFFARX1 I_29072 (I496926,I2683,I496592,I496952,);
nor I_29073 (I496960,I496952,I496819);
DFFARX1 I_29074 (I496960,I2683,I496592,I496560,);
nand I_29075 (I496991,I496952,I496861);
nand I_29076 (I496569,I496844,I496991);
not I_29077 (I497022,I496952);
nor I_29078 (I497039,I497022,I496762);
DFFARX1 I_29079 (I497039,I2683,I496592,I496581,);
nor I_29080 (I497070,I892375,I892357);
or I_29081 (I496572,I496819,I497070);
nor I_29082 (I496563,I496952,I497070);
or I_29083 (I496566,I496686,I497070);
DFFARX1 I_29084 (I497070,I2683,I496592,I496584,);
not I_29085 (I497170,I2690);
DFFARX1 I_29086 (I331771,I2683,I497170,I497196,);
not I_29087 (I497204,I497196);
nand I_29088 (I497221,I331762,I331780);
and I_29089 (I497238,I497221,I331783);
DFFARX1 I_29090 (I497238,I2683,I497170,I497264,);
not I_29091 (I497272,I331777);
DFFARX1 I_29092 (I331765,I2683,I497170,I497298,);
not I_29093 (I497306,I497298);
nor I_29094 (I497323,I497306,I497204);
and I_29095 (I497340,I497323,I331777);
nor I_29096 (I497357,I497306,I497272);
nor I_29097 (I497153,I497264,I497357);
DFFARX1 I_29098 (I331774,I2683,I497170,I497397,);
nor I_29099 (I497405,I497397,I497264);
not I_29100 (I497422,I497405);
not I_29101 (I497439,I497397);
nor I_29102 (I497456,I497439,I497340);
DFFARX1 I_29103 (I497456,I2683,I497170,I497156,);
nand I_29104 (I497487,I331789,I331786);
and I_29105 (I497504,I497487,I331768);
DFFARX1 I_29106 (I497504,I2683,I497170,I497530,);
nor I_29107 (I497538,I497530,I497397);
DFFARX1 I_29108 (I497538,I2683,I497170,I497138,);
nand I_29109 (I497569,I497530,I497439);
nand I_29110 (I497147,I497422,I497569);
not I_29111 (I497600,I497530);
nor I_29112 (I497617,I497600,I497340);
DFFARX1 I_29113 (I497617,I2683,I497170,I497159,);
nor I_29114 (I497648,I331762,I331786);
or I_29115 (I497150,I497397,I497648);
nor I_29116 (I497141,I497530,I497648);
or I_29117 (I497144,I497264,I497648);
DFFARX1 I_29118 (I497648,I2683,I497170,I497162,);
not I_29119 (I497748,I2690);
DFFARX1 I_29120 (I351355,I2683,I497748,I497774,);
not I_29121 (I497782,I497774);
nand I_29122 (I497799,I351346,I351364);
and I_29123 (I497816,I497799,I351367);
DFFARX1 I_29124 (I497816,I2683,I497748,I497842,);
not I_29125 (I497850,I351361);
DFFARX1 I_29126 (I351349,I2683,I497748,I497876,);
not I_29127 (I497884,I497876);
nor I_29128 (I497901,I497884,I497782);
and I_29129 (I497918,I497901,I351361);
nor I_29130 (I497935,I497884,I497850);
nor I_29131 (I497731,I497842,I497935);
DFFARX1 I_29132 (I351358,I2683,I497748,I497975,);
nor I_29133 (I497983,I497975,I497842);
not I_29134 (I498000,I497983);
not I_29135 (I498017,I497975);
nor I_29136 (I498034,I498017,I497918);
DFFARX1 I_29137 (I498034,I2683,I497748,I497734,);
nand I_29138 (I498065,I351373,I351370);
and I_29139 (I498082,I498065,I351352);
DFFARX1 I_29140 (I498082,I2683,I497748,I498108,);
nor I_29141 (I498116,I498108,I497975);
DFFARX1 I_29142 (I498116,I2683,I497748,I497716,);
nand I_29143 (I498147,I498108,I498017);
nand I_29144 (I497725,I498000,I498147);
not I_29145 (I498178,I498108);
nor I_29146 (I498195,I498178,I497918);
DFFARX1 I_29147 (I498195,I2683,I497748,I497737,);
nor I_29148 (I498226,I351346,I351370);
or I_29149 (I497728,I497975,I498226);
nor I_29150 (I497719,I498108,I498226);
or I_29151 (I497722,I497842,I498226);
DFFARX1 I_29152 (I498226,I2683,I497748,I497740,);
not I_29153 (I498326,I2690);
DFFARX1 I_29154 (I1089411,I2683,I498326,I498352,);
not I_29155 (I498360,I498352);
nand I_29156 (I498377,I1089396,I1089384);
and I_29157 (I498394,I498377,I1089399);
DFFARX1 I_29158 (I498394,I2683,I498326,I498420,);
not I_29159 (I498428,I1089384);
DFFARX1 I_29160 (I1089402,I2683,I498326,I498454,);
not I_29161 (I498462,I498454);
nor I_29162 (I498479,I498462,I498360);
and I_29163 (I498496,I498479,I1089384);
nor I_29164 (I498513,I498462,I498428);
nor I_29165 (I498309,I498420,I498513);
DFFARX1 I_29166 (I1089390,I2683,I498326,I498553,);
nor I_29167 (I498561,I498553,I498420);
not I_29168 (I498578,I498561);
not I_29169 (I498595,I498553);
nor I_29170 (I498612,I498595,I498496);
DFFARX1 I_29171 (I498612,I2683,I498326,I498312,);
nand I_29172 (I498643,I1089387,I1089393);
and I_29173 (I498660,I498643,I1089408);
DFFARX1 I_29174 (I498660,I2683,I498326,I498686,);
nor I_29175 (I498694,I498686,I498553);
DFFARX1 I_29176 (I498694,I2683,I498326,I498294,);
nand I_29177 (I498725,I498686,I498595);
nand I_29178 (I498303,I498578,I498725);
not I_29179 (I498756,I498686);
nor I_29180 (I498773,I498756,I498496);
DFFARX1 I_29181 (I498773,I2683,I498326,I498315,);
nor I_29182 (I498804,I1089405,I1089393);
or I_29183 (I498306,I498553,I498804);
nor I_29184 (I498297,I498686,I498804);
or I_29185 (I498300,I498420,I498804);
DFFARX1 I_29186 (I498804,I2683,I498326,I498318,);
not I_29187 (I498904,I2690);
DFFARX1 I_29188 (I891794,I2683,I498904,I498930,);
not I_29189 (I498938,I498930);
nand I_29190 (I498955,I891776,I891788);
and I_29191 (I498972,I498955,I891791);
DFFARX1 I_29192 (I498972,I2683,I498904,I498998,);
not I_29193 (I499006,I891785);
DFFARX1 I_29194 (I891782,I2683,I498904,I499032,);
not I_29195 (I499040,I499032);
nor I_29196 (I499057,I499040,I498938);
and I_29197 (I499074,I499057,I891785);
nor I_29198 (I499091,I499040,I499006);
nor I_29199 (I498887,I498998,I499091);
DFFARX1 I_29200 (I891800,I2683,I498904,I499131,);
nor I_29201 (I499139,I499131,I498998);
not I_29202 (I499156,I499139);
not I_29203 (I499173,I499131);
nor I_29204 (I499190,I499173,I499074);
DFFARX1 I_29205 (I499190,I2683,I498904,I498890,);
nand I_29206 (I499221,I891779,I891779);
and I_29207 (I499238,I499221,I891776);
DFFARX1 I_29208 (I499238,I2683,I498904,I499264,);
nor I_29209 (I499272,I499264,I499131);
DFFARX1 I_29210 (I499272,I2683,I498904,I498872,);
nand I_29211 (I499303,I499264,I499173);
nand I_29212 (I498881,I499156,I499303);
not I_29213 (I499334,I499264);
nor I_29214 (I499351,I499334,I499074);
DFFARX1 I_29215 (I499351,I2683,I498904,I498893,);
nor I_29216 (I499382,I891797,I891779);
or I_29217 (I498884,I499131,I499382);
nor I_29218 (I498875,I499264,I499382);
or I_29219 (I498878,I498998,I499382);
DFFARX1 I_29220 (I499382,I2683,I498904,I498896,);
not I_29221 (I499482,I2690);
DFFARX1 I_29222 (I362235,I2683,I499482,I499508,);
not I_29223 (I499516,I499508);
nand I_29224 (I499533,I362226,I362244);
and I_29225 (I499550,I499533,I362247);
DFFARX1 I_29226 (I499550,I2683,I499482,I499576,);
not I_29227 (I499584,I362241);
DFFARX1 I_29228 (I362229,I2683,I499482,I499610,);
not I_29229 (I499618,I499610);
nor I_29230 (I499635,I499618,I499516);
and I_29231 (I499652,I499635,I362241);
nor I_29232 (I499669,I499618,I499584);
nor I_29233 (I499465,I499576,I499669);
DFFARX1 I_29234 (I362238,I2683,I499482,I499709,);
nor I_29235 (I499717,I499709,I499576);
not I_29236 (I499734,I499717);
not I_29237 (I499751,I499709);
nor I_29238 (I499768,I499751,I499652);
DFFARX1 I_29239 (I499768,I2683,I499482,I499468,);
nand I_29240 (I499799,I362253,I362250);
and I_29241 (I499816,I499799,I362232);
DFFARX1 I_29242 (I499816,I2683,I499482,I499842,);
nor I_29243 (I499850,I499842,I499709);
DFFARX1 I_29244 (I499850,I2683,I499482,I499450,);
nand I_29245 (I499881,I499842,I499751);
nand I_29246 (I499459,I499734,I499881);
not I_29247 (I499912,I499842);
nor I_29248 (I499929,I499912,I499652);
DFFARX1 I_29249 (I499929,I2683,I499482,I499471,);
nor I_29250 (I499960,I362226,I362250);
or I_29251 (I499462,I499709,I499960);
nor I_29252 (I499453,I499842,I499960);
or I_29253 (I499456,I499576,I499960);
DFFARX1 I_29254 (I499960,I2683,I499482,I499474,);
not I_29255 (I500060,I2690);
DFFARX1 I_29256 (I869830,I2683,I500060,I500086,);
not I_29257 (I500094,I500086);
nand I_29258 (I500111,I869812,I869824);
and I_29259 (I500128,I500111,I869827);
DFFARX1 I_29260 (I500128,I2683,I500060,I500154,);
not I_29261 (I500162,I869821);
DFFARX1 I_29262 (I869818,I2683,I500060,I500188,);
not I_29263 (I500196,I500188);
nor I_29264 (I500213,I500196,I500094);
and I_29265 (I500230,I500213,I869821);
nor I_29266 (I500247,I500196,I500162);
nor I_29267 (I500043,I500154,I500247);
DFFARX1 I_29268 (I869836,I2683,I500060,I500287,);
nor I_29269 (I500295,I500287,I500154);
not I_29270 (I500312,I500295);
not I_29271 (I500329,I500287);
nor I_29272 (I500346,I500329,I500230);
DFFARX1 I_29273 (I500346,I2683,I500060,I500046,);
nand I_29274 (I500377,I869815,I869815);
and I_29275 (I500394,I500377,I869812);
DFFARX1 I_29276 (I500394,I2683,I500060,I500420,);
nor I_29277 (I500428,I500420,I500287);
DFFARX1 I_29278 (I500428,I2683,I500060,I500028,);
nand I_29279 (I500459,I500420,I500329);
nand I_29280 (I500037,I500312,I500459);
not I_29281 (I500490,I500420);
nor I_29282 (I500507,I500490,I500230);
DFFARX1 I_29283 (I500507,I2683,I500060,I500049,);
nor I_29284 (I500538,I869833,I869815);
or I_29285 (I500040,I500287,I500538);
nor I_29286 (I500031,I500420,I500538);
or I_29287 (I500034,I500154,I500538);
DFFARX1 I_29288 (I500538,I2683,I500060,I500052,);
not I_29289 (I500638,I2690);
DFFARX1 I_29290 (I171775,I2683,I500638,I500664,);
not I_29291 (I500672,I500664);
nand I_29292 (I500689,I171778,I171799);
and I_29293 (I500706,I500689,I171787);
DFFARX1 I_29294 (I500706,I2683,I500638,I500732,);
not I_29295 (I500740,I171784);
DFFARX1 I_29296 (I171775,I2683,I500638,I500766,);
not I_29297 (I500774,I500766);
nor I_29298 (I500791,I500774,I500672);
and I_29299 (I500808,I500791,I171784);
nor I_29300 (I500825,I500774,I500740);
nor I_29301 (I500621,I500732,I500825);
DFFARX1 I_29302 (I171793,I2683,I500638,I500865,);
nor I_29303 (I500873,I500865,I500732);
not I_29304 (I500890,I500873);
not I_29305 (I500907,I500865);
nor I_29306 (I500924,I500907,I500808);
DFFARX1 I_29307 (I500924,I2683,I500638,I500624,);
nand I_29308 (I500955,I171778,I171781);
and I_29309 (I500972,I500955,I171790);
DFFARX1 I_29310 (I500972,I2683,I500638,I500998,);
nor I_29311 (I501006,I500998,I500865);
DFFARX1 I_29312 (I501006,I2683,I500638,I500606,);
nand I_29313 (I501037,I500998,I500907);
nand I_29314 (I500615,I500890,I501037);
not I_29315 (I501068,I500998);
nor I_29316 (I501085,I501068,I500808);
DFFARX1 I_29317 (I501085,I2683,I500638,I500627,);
nor I_29318 (I501116,I171796,I171781);
or I_29319 (I500618,I500865,I501116);
nor I_29320 (I500609,I500998,I501116);
or I_29321 (I500612,I500732,I501116);
DFFARX1 I_29322 (I501116,I2683,I500638,I500630,);
not I_29323 (I501216,I2690);
DFFARX1 I_29324 (I150355,I2683,I501216,I501242,);
not I_29325 (I501250,I501242);
nand I_29326 (I501267,I150358,I150379);
and I_29327 (I501284,I501267,I150367);
DFFARX1 I_29328 (I501284,I2683,I501216,I501310,);
not I_29329 (I501318,I150364);
DFFARX1 I_29330 (I150355,I2683,I501216,I501344,);
not I_29331 (I501352,I501344);
nor I_29332 (I501369,I501352,I501250);
and I_29333 (I501386,I501369,I150364);
nor I_29334 (I501403,I501352,I501318);
nor I_29335 (I501199,I501310,I501403);
DFFARX1 I_29336 (I150373,I2683,I501216,I501443,);
nor I_29337 (I501451,I501443,I501310);
not I_29338 (I501468,I501451);
not I_29339 (I501485,I501443);
nor I_29340 (I501502,I501485,I501386);
DFFARX1 I_29341 (I501502,I2683,I501216,I501202,);
nand I_29342 (I501533,I150358,I150361);
and I_29343 (I501550,I501533,I150370);
DFFARX1 I_29344 (I501550,I2683,I501216,I501576,);
nor I_29345 (I501584,I501576,I501443);
DFFARX1 I_29346 (I501584,I2683,I501216,I501184,);
nand I_29347 (I501615,I501576,I501485);
nand I_29348 (I501193,I501468,I501615);
not I_29349 (I501646,I501576);
nor I_29350 (I501663,I501646,I501386);
DFFARX1 I_29351 (I501663,I2683,I501216,I501205,);
nor I_29352 (I501694,I150376,I150361);
or I_29353 (I501196,I501443,I501694);
nor I_29354 (I501187,I501576,I501694);
or I_29355 (I501190,I501310,I501694);
DFFARX1 I_29356 (I501694,I2683,I501216,I501208,);
not I_29357 (I501794,I2690);
DFFARX1 I_29358 (I115262,I2683,I501794,I501820,);
not I_29359 (I501828,I501820);
nand I_29360 (I501845,I115277,I115250);
and I_29361 (I501862,I501845,I115265);
DFFARX1 I_29362 (I501862,I2683,I501794,I501888,);
not I_29363 (I501896,I115268);
DFFARX1 I_29364 (I115253,I2683,I501794,I501922,);
not I_29365 (I501930,I501922);
nor I_29366 (I501947,I501930,I501828);
and I_29367 (I501964,I501947,I115268);
nor I_29368 (I501981,I501930,I501896);
nor I_29369 (I501777,I501888,I501981);
DFFARX1 I_29370 (I115259,I2683,I501794,I502021,);
nor I_29371 (I502029,I502021,I501888);
not I_29372 (I502046,I502029);
not I_29373 (I502063,I502021);
nor I_29374 (I502080,I502063,I501964);
DFFARX1 I_29375 (I502080,I2683,I501794,I501780,);
nand I_29376 (I502111,I115274,I115256);
and I_29377 (I502128,I502111,I115271);
DFFARX1 I_29378 (I502128,I2683,I501794,I502154,);
nor I_29379 (I502162,I502154,I502021);
DFFARX1 I_29380 (I502162,I2683,I501794,I501762,);
nand I_29381 (I502193,I502154,I502063);
nand I_29382 (I501771,I502046,I502193);
not I_29383 (I502224,I502154);
nor I_29384 (I502241,I502224,I501964);
DFFARX1 I_29385 (I502241,I2683,I501794,I501783,);
nor I_29386 (I502272,I115250,I115256);
or I_29387 (I501774,I502021,I502272);
nor I_29388 (I501765,I502154,I502272);
or I_29389 (I501768,I501888,I502272);
DFFARX1 I_29390 (I502272,I2683,I501794,I501786,);
not I_29391 (I502372,I2690);
DFFARX1 I_29392 (I828214,I2683,I502372,I502398,);
not I_29393 (I502406,I502398);
nand I_29394 (I502423,I828196,I828208);
and I_29395 (I502440,I502423,I828211);
DFFARX1 I_29396 (I502440,I2683,I502372,I502466,);
not I_29397 (I502474,I828205);
DFFARX1 I_29398 (I828202,I2683,I502372,I502500,);
not I_29399 (I502508,I502500);
nor I_29400 (I502525,I502508,I502406);
and I_29401 (I502542,I502525,I828205);
nor I_29402 (I502559,I502508,I502474);
nor I_29403 (I502355,I502466,I502559);
DFFARX1 I_29404 (I828220,I2683,I502372,I502599,);
nor I_29405 (I502607,I502599,I502466);
not I_29406 (I502624,I502607);
not I_29407 (I502641,I502599);
nor I_29408 (I502658,I502641,I502542);
DFFARX1 I_29409 (I502658,I2683,I502372,I502358,);
nand I_29410 (I502689,I828199,I828199);
and I_29411 (I502706,I502689,I828196);
DFFARX1 I_29412 (I502706,I2683,I502372,I502732,);
nor I_29413 (I502740,I502732,I502599);
DFFARX1 I_29414 (I502740,I2683,I502372,I502340,);
nand I_29415 (I502771,I502732,I502641);
nand I_29416 (I502349,I502624,I502771);
not I_29417 (I502802,I502732);
nor I_29418 (I502819,I502802,I502542);
DFFARX1 I_29419 (I502819,I2683,I502372,I502361,);
nor I_29420 (I502850,I828217,I828199);
or I_29421 (I502352,I502599,I502850);
nor I_29422 (I502343,I502732,I502850);
or I_29423 (I502346,I502466,I502850);
DFFARX1 I_29424 (I502850,I2683,I502372,I502364,);
not I_29425 (I502950,I2690);
DFFARX1 I_29426 (I1076916,I2683,I502950,I502976,);
not I_29427 (I502984,I502976);
nand I_29428 (I503001,I1076901,I1076889);
and I_29429 (I503018,I503001,I1076904);
DFFARX1 I_29430 (I503018,I2683,I502950,I503044,);
not I_29431 (I503052,I1076889);
DFFARX1 I_29432 (I1076907,I2683,I502950,I503078,);
not I_29433 (I503086,I503078);
nor I_29434 (I503103,I503086,I502984);
and I_29435 (I503120,I503103,I1076889);
nor I_29436 (I503137,I503086,I503052);
nor I_29437 (I502933,I503044,I503137);
DFFARX1 I_29438 (I1076895,I2683,I502950,I503177,);
nor I_29439 (I503185,I503177,I503044);
not I_29440 (I503202,I503185);
not I_29441 (I503219,I503177);
nor I_29442 (I503236,I503219,I503120);
DFFARX1 I_29443 (I503236,I2683,I502950,I502936,);
nand I_29444 (I503267,I1076892,I1076898);
and I_29445 (I503284,I503267,I1076913);
DFFARX1 I_29446 (I503284,I2683,I502950,I503310,);
nor I_29447 (I503318,I503310,I503177);
DFFARX1 I_29448 (I503318,I2683,I502950,I502918,);
nand I_29449 (I503349,I503310,I503219);
nand I_29450 (I502927,I503202,I503349);
not I_29451 (I503380,I503310);
nor I_29452 (I503397,I503380,I503120);
DFFARX1 I_29453 (I503397,I2683,I502950,I502939,);
nor I_29454 (I503428,I1076910,I1076898);
or I_29455 (I502930,I503177,I503428);
nor I_29456 (I502921,I503310,I503428);
or I_29457 (I502924,I503044,I503428);
DFFARX1 I_29458 (I503428,I2683,I502950,I502942,);
not I_29459 (I503528,I2690);
DFFARX1 I_29460 (I382363,I2683,I503528,I503554,);
not I_29461 (I503562,I503554);
nand I_29462 (I503579,I382354,I382372);
and I_29463 (I503596,I503579,I382375);
DFFARX1 I_29464 (I503596,I2683,I503528,I503622,);
not I_29465 (I503630,I382369);
DFFARX1 I_29466 (I382357,I2683,I503528,I503656,);
not I_29467 (I503664,I503656);
nor I_29468 (I503681,I503664,I503562);
and I_29469 (I503698,I503681,I382369);
nor I_29470 (I503715,I503664,I503630);
nor I_29471 (I503511,I503622,I503715);
DFFARX1 I_29472 (I382366,I2683,I503528,I503755,);
nor I_29473 (I503763,I503755,I503622);
not I_29474 (I503780,I503763);
not I_29475 (I503797,I503755);
nor I_29476 (I503814,I503797,I503698);
DFFARX1 I_29477 (I503814,I2683,I503528,I503514,);
nand I_29478 (I503845,I382381,I382378);
and I_29479 (I503862,I503845,I382360);
DFFARX1 I_29480 (I503862,I2683,I503528,I503888,);
nor I_29481 (I503896,I503888,I503755);
DFFARX1 I_29482 (I503896,I2683,I503528,I503496,);
nand I_29483 (I503927,I503888,I503797);
nand I_29484 (I503505,I503780,I503927);
not I_29485 (I503958,I503888);
nor I_29486 (I503975,I503958,I503698);
DFFARX1 I_29487 (I503975,I2683,I503528,I503517,);
nor I_29488 (I504006,I382354,I382378);
or I_29489 (I503508,I503755,I504006);
nor I_29490 (I503499,I503888,I504006);
or I_29491 (I503502,I503622,I504006);
DFFARX1 I_29492 (I504006,I2683,I503528,I503520,);
not I_29493 (I504106,I2690);
DFFARX1 I_29494 (I232744,I2683,I504106,I504132,);
not I_29495 (I504140,I504132);
nand I_29496 (I504157,I232747,I232723);
and I_29497 (I504174,I504157,I232720);
DFFARX1 I_29498 (I504174,I2683,I504106,I504200,);
not I_29499 (I504208,I232726);
DFFARX1 I_29500 (I232720,I2683,I504106,I504234,);
not I_29501 (I504242,I504234);
nor I_29502 (I504259,I504242,I504140);
and I_29503 (I504276,I504259,I232726);
nor I_29504 (I504293,I504242,I504208);
nor I_29505 (I504089,I504200,I504293);
DFFARX1 I_29506 (I232729,I2683,I504106,I504333,);
nor I_29507 (I504341,I504333,I504200);
not I_29508 (I504358,I504341);
not I_29509 (I504375,I504333);
nor I_29510 (I504392,I504375,I504276);
DFFARX1 I_29511 (I504392,I2683,I504106,I504092,);
nand I_29512 (I504423,I232732,I232741);
and I_29513 (I504440,I504423,I232738);
DFFARX1 I_29514 (I504440,I2683,I504106,I504466,);
nor I_29515 (I504474,I504466,I504333);
DFFARX1 I_29516 (I504474,I2683,I504106,I504074,);
nand I_29517 (I504505,I504466,I504375);
nand I_29518 (I504083,I504358,I504505);
not I_29519 (I504536,I504466);
nor I_29520 (I504553,I504536,I504276);
DFFARX1 I_29521 (I504553,I2683,I504106,I504095,);
nor I_29522 (I504584,I232735,I232741);
or I_29523 (I504086,I504333,I504584);
nor I_29524 (I504077,I504466,I504584);
or I_29525 (I504080,I504200,I504584);
DFFARX1 I_29526 (I504584,I2683,I504106,I504098,);
not I_29527 (I504684,I2690);
DFFARX1 I_29528 (I145595,I2683,I504684,I504710,);
not I_29529 (I504718,I504710);
nand I_29530 (I504735,I145598,I145619);
and I_29531 (I504752,I504735,I145607);
DFFARX1 I_29532 (I504752,I2683,I504684,I504778,);
not I_29533 (I504786,I145604);
DFFARX1 I_29534 (I145595,I2683,I504684,I504812,);
not I_29535 (I504820,I504812);
nor I_29536 (I504837,I504820,I504718);
and I_29537 (I504854,I504837,I145604);
nor I_29538 (I504871,I504820,I504786);
nor I_29539 (I504667,I504778,I504871);
DFFARX1 I_29540 (I145613,I2683,I504684,I504911,);
nor I_29541 (I504919,I504911,I504778);
not I_29542 (I504936,I504919);
not I_29543 (I504953,I504911);
nor I_29544 (I504970,I504953,I504854);
DFFARX1 I_29545 (I504970,I2683,I504684,I504670,);
nand I_29546 (I505001,I145598,I145601);
and I_29547 (I505018,I505001,I145610);
DFFARX1 I_29548 (I505018,I2683,I504684,I505044,);
nor I_29549 (I505052,I505044,I504911);
DFFARX1 I_29550 (I505052,I2683,I504684,I504652,);
nand I_29551 (I505083,I505044,I504953);
nand I_29552 (I504661,I504936,I505083);
not I_29553 (I505114,I505044);
nor I_29554 (I505131,I505114,I504854);
DFFARX1 I_29555 (I505131,I2683,I504684,I504673,);
nor I_29556 (I505162,I145616,I145601);
or I_29557 (I504664,I504911,I505162);
nor I_29558 (I504655,I505044,I505162);
or I_29559 (I504658,I504778,I505162);
DFFARX1 I_29560 (I505162,I2683,I504684,I504676,);
not I_29561 (I505262,I2690);
DFFARX1 I_29562 (I34291,I2683,I505262,I505288,);
not I_29563 (I505296,I505288);
nand I_29564 (I505313,I34288,I34279);
and I_29565 (I505330,I505313,I34279);
DFFARX1 I_29566 (I505330,I2683,I505262,I505356,);
not I_29567 (I505364,I34282);
DFFARX1 I_29568 (I34297,I2683,I505262,I505390,);
not I_29569 (I505398,I505390);
nor I_29570 (I505415,I505398,I505296);
and I_29571 (I505432,I505415,I34282);
nor I_29572 (I505449,I505398,I505364);
nor I_29573 (I505245,I505356,I505449);
DFFARX1 I_29574 (I34282,I2683,I505262,I505489,);
nor I_29575 (I505497,I505489,I505356);
not I_29576 (I505514,I505497);
not I_29577 (I505531,I505489);
nor I_29578 (I505548,I505531,I505432);
DFFARX1 I_29579 (I505548,I2683,I505262,I505248,);
nand I_29580 (I505579,I34300,I34285);
and I_29581 (I505596,I505579,I34303);
DFFARX1 I_29582 (I505596,I2683,I505262,I505622,);
nor I_29583 (I505630,I505622,I505489);
DFFARX1 I_29584 (I505630,I2683,I505262,I505230,);
nand I_29585 (I505661,I505622,I505531);
nand I_29586 (I505239,I505514,I505661);
not I_29587 (I505692,I505622);
nor I_29588 (I505709,I505692,I505432);
DFFARX1 I_29589 (I505709,I2683,I505262,I505251,);
nor I_29590 (I505740,I34294,I34285);
or I_29591 (I505242,I505489,I505740);
nor I_29592 (I505233,I505622,I505740);
or I_29593 (I505236,I505356,I505740);
DFFARX1 I_29594 (I505740,I2683,I505262,I505254,);
not I_29595 (I505840,I2690);
DFFARX1 I_29596 (I143215,I2683,I505840,I505866,);
not I_29597 (I505874,I505866);
nand I_29598 (I505891,I143218,I143239);
and I_29599 (I505908,I505891,I143227);
DFFARX1 I_29600 (I505908,I2683,I505840,I505934,);
not I_29601 (I505942,I143224);
DFFARX1 I_29602 (I143215,I2683,I505840,I505968,);
not I_29603 (I505976,I505968);
nor I_29604 (I505993,I505976,I505874);
and I_29605 (I506010,I505993,I143224);
nor I_29606 (I506027,I505976,I505942);
nor I_29607 (I505823,I505934,I506027);
DFFARX1 I_29608 (I143233,I2683,I505840,I506067,);
nor I_29609 (I506075,I506067,I505934);
not I_29610 (I506092,I506075);
not I_29611 (I506109,I506067);
nor I_29612 (I506126,I506109,I506010);
DFFARX1 I_29613 (I506126,I2683,I505840,I505826,);
nand I_29614 (I506157,I143218,I143221);
and I_29615 (I506174,I506157,I143230);
DFFARX1 I_29616 (I506174,I2683,I505840,I506200,);
nor I_29617 (I506208,I506200,I506067);
DFFARX1 I_29618 (I506208,I2683,I505840,I505808,);
nand I_29619 (I506239,I506200,I506109);
nand I_29620 (I505817,I506092,I506239);
not I_29621 (I506270,I506200);
nor I_29622 (I506287,I506270,I506010);
DFFARX1 I_29623 (I506287,I2683,I505840,I505829,);
nor I_29624 (I506318,I143236,I143221);
or I_29625 (I505820,I506067,I506318);
nor I_29626 (I505811,I506200,I506318);
or I_29627 (I505814,I505934,I506318);
DFFARX1 I_29628 (I506318,I2683,I505840,I505832,);
not I_29629 (I506418,I2690);
DFFARX1 I_29630 (I213772,I2683,I506418,I506444,);
not I_29631 (I506452,I506444);
nand I_29632 (I506469,I213775,I213751);
and I_29633 (I506486,I506469,I213748);
DFFARX1 I_29634 (I506486,I2683,I506418,I506512,);
not I_29635 (I506520,I213754);
DFFARX1 I_29636 (I213748,I2683,I506418,I506546,);
not I_29637 (I506554,I506546);
nor I_29638 (I506571,I506554,I506452);
and I_29639 (I506588,I506571,I213754);
nor I_29640 (I506605,I506554,I506520);
nor I_29641 (I506401,I506512,I506605);
DFFARX1 I_29642 (I213757,I2683,I506418,I506645,);
nor I_29643 (I506653,I506645,I506512);
not I_29644 (I506670,I506653);
not I_29645 (I506687,I506645);
nor I_29646 (I506704,I506687,I506588);
DFFARX1 I_29647 (I506704,I2683,I506418,I506404,);
nand I_29648 (I506735,I213760,I213769);
and I_29649 (I506752,I506735,I213766);
DFFARX1 I_29650 (I506752,I2683,I506418,I506778,);
nor I_29651 (I506786,I506778,I506645);
DFFARX1 I_29652 (I506786,I2683,I506418,I506386,);
nand I_29653 (I506817,I506778,I506687);
nand I_29654 (I506395,I506670,I506817);
not I_29655 (I506848,I506778);
nor I_29656 (I506865,I506848,I506588);
DFFARX1 I_29657 (I506865,I2683,I506418,I506407,);
nor I_29658 (I506896,I213763,I213769);
or I_29659 (I506398,I506645,I506896);
nor I_29660 (I506389,I506778,I506896);
or I_29661 (I506392,I506512,I506896);
DFFARX1 I_29662 (I506896,I2683,I506418,I506410,);
not I_29663 (I506996,I2690);
DFFARX1 I_29664 (I801835,I2683,I506996,I507022,);
not I_29665 (I507030,I507022);
nand I_29666 (I507047,I801832,I801850);
and I_29667 (I507064,I507047,I801847);
DFFARX1 I_29668 (I507064,I2683,I506996,I507090,);
not I_29669 (I507098,I801829);
DFFARX1 I_29670 (I801832,I2683,I506996,I507124,);
not I_29671 (I507132,I507124);
nor I_29672 (I507149,I507132,I507030);
and I_29673 (I507166,I507149,I801829);
nor I_29674 (I507183,I507132,I507098);
nor I_29675 (I506979,I507090,I507183);
DFFARX1 I_29676 (I801841,I2683,I506996,I507223,);
nor I_29677 (I507231,I507223,I507090);
not I_29678 (I507248,I507231);
not I_29679 (I507265,I507223);
nor I_29680 (I507282,I507265,I507166);
DFFARX1 I_29681 (I507282,I2683,I506996,I506982,);
nand I_29682 (I507313,I801844,I801829);
and I_29683 (I507330,I507313,I801835);
DFFARX1 I_29684 (I507330,I2683,I506996,I507356,);
nor I_29685 (I507364,I507356,I507223);
DFFARX1 I_29686 (I507364,I2683,I506996,I506964,);
nand I_29687 (I507395,I507356,I507265);
nand I_29688 (I506973,I507248,I507395);
not I_29689 (I507426,I507356);
nor I_29690 (I507443,I507426,I507166);
DFFARX1 I_29691 (I507443,I2683,I506996,I506985,);
nor I_29692 (I507474,I801838,I801829);
or I_29693 (I506976,I507223,I507474);
nor I_29694 (I506967,I507356,I507474);
or I_29695 (I506970,I507090,I507474);
DFFARX1 I_29696 (I507474,I2683,I506996,I506988,);
not I_29697 (I507574,I2690);
DFFARX1 I_29698 (I833994,I2683,I507574,I507600,);
not I_29699 (I507608,I507600);
nand I_29700 (I507625,I833976,I833988);
and I_29701 (I507642,I507625,I833991);
DFFARX1 I_29702 (I507642,I2683,I507574,I507668,);
not I_29703 (I507676,I833985);
DFFARX1 I_29704 (I833982,I2683,I507574,I507702,);
not I_29705 (I507710,I507702);
nor I_29706 (I507727,I507710,I507608);
and I_29707 (I507744,I507727,I833985);
nor I_29708 (I507761,I507710,I507676);
nor I_29709 (I507557,I507668,I507761);
DFFARX1 I_29710 (I834000,I2683,I507574,I507801,);
nor I_29711 (I507809,I507801,I507668);
not I_29712 (I507826,I507809);
not I_29713 (I507843,I507801);
nor I_29714 (I507860,I507843,I507744);
DFFARX1 I_29715 (I507860,I2683,I507574,I507560,);
nand I_29716 (I507891,I833979,I833979);
and I_29717 (I507908,I507891,I833976);
DFFARX1 I_29718 (I507908,I2683,I507574,I507934,);
nor I_29719 (I507942,I507934,I507801);
DFFARX1 I_29720 (I507942,I2683,I507574,I507542,);
nand I_29721 (I507973,I507934,I507843);
nand I_29722 (I507551,I507826,I507973);
not I_29723 (I508004,I507934);
nor I_29724 (I508021,I508004,I507744);
DFFARX1 I_29725 (I508021,I2683,I507574,I507563,);
nor I_29726 (I508052,I833997,I833979);
or I_29727 (I507554,I507801,I508052);
nor I_29728 (I507545,I507934,I508052);
or I_29729 (I507548,I507668,I508052);
DFFARX1 I_29730 (I508052,I2683,I507574,I507566,);
not I_29731 (I508152,I2690);
DFFARX1 I_29732 (I493670,I2683,I508152,I508178,);
not I_29733 (I508186,I508178);
nand I_29734 (I508203,I493679,I493688);
and I_29735 (I508220,I508203,I493694);
DFFARX1 I_29736 (I508220,I2683,I508152,I508246,);
not I_29737 (I508254,I493691);
DFFARX1 I_29738 (I493676,I2683,I508152,I508280,);
not I_29739 (I508288,I508280);
nor I_29740 (I508305,I508288,I508186);
and I_29741 (I508322,I508305,I493691);
nor I_29742 (I508339,I508288,I508254);
nor I_29743 (I508135,I508246,I508339);
DFFARX1 I_29744 (I493685,I2683,I508152,I508379,);
nor I_29745 (I508387,I508379,I508246);
not I_29746 (I508404,I508387);
not I_29747 (I508421,I508379);
nor I_29748 (I508438,I508421,I508322);
DFFARX1 I_29749 (I508438,I2683,I508152,I508138,);
nand I_29750 (I508469,I493682,I493673);
and I_29751 (I508486,I508469,I493670);
DFFARX1 I_29752 (I508486,I2683,I508152,I508512,);
nor I_29753 (I508520,I508512,I508379);
DFFARX1 I_29754 (I508520,I2683,I508152,I508120,);
nand I_29755 (I508551,I508512,I508421);
nand I_29756 (I508129,I508404,I508551);
not I_29757 (I508582,I508512);
nor I_29758 (I508599,I508582,I508322);
DFFARX1 I_29759 (I508599,I2683,I508152,I508141,);
nor I_29760 (I508630,I493673,I493673);
or I_29761 (I508132,I508379,I508630);
nor I_29762 (I508123,I508512,I508630);
or I_29763 (I508126,I508246,I508630);
DFFARX1 I_29764 (I508630,I2683,I508152,I508144,);
not I_29765 (I508730,I2690);
DFFARX1 I_29766 (I95414,I2683,I508730,I508756,);
not I_29767 (I508764,I508756);
nand I_29768 (I508781,I95423,I95432);
and I_29769 (I508798,I508781,I95411);
DFFARX1 I_29770 (I508798,I2683,I508730,I508824,);
not I_29771 (I508832,I95414);
DFFARX1 I_29772 (I95429,I2683,I508730,I508858,);
not I_29773 (I508866,I508858);
nor I_29774 (I508883,I508866,I508764);
and I_29775 (I508900,I508883,I95414);
nor I_29776 (I508917,I508866,I508832);
nor I_29777 (I508713,I508824,I508917);
DFFARX1 I_29778 (I95420,I2683,I508730,I508957,);
nor I_29779 (I508965,I508957,I508824);
not I_29780 (I508982,I508965);
not I_29781 (I508999,I508957);
nor I_29782 (I509016,I508999,I508900);
DFFARX1 I_29783 (I509016,I2683,I508730,I508716,);
nand I_29784 (I509047,I95435,I95411);
and I_29785 (I509064,I509047,I95417);
DFFARX1 I_29786 (I509064,I2683,I508730,I509090,);
nor I_29787 (I509098,I509090,I508957);
DFFARX1 I_29788 (I509098,I2683,I508730,I508698,);
nand I_29789 (I509129,I509090,I508999);
nand I_29790 (I508707,I508982,I509129);
not I_29791 (I509160,I509090);
nor I_29792 (I509177,I509160,I508900);
DFFARX1 I_29793 (I509177,I2683,I508730,I508719,);
nor I_29794 (I509208,I95426,I95411);
or I_29795 (I508710,I508957,I509208);
nor I_29796 (I508701,I509090,I509208);
or I_29797 (I508704,I508824,I509208);
DFFARX1 I_29798 (I509208,I2683,I508730,I508722,);
not I_29799 (I509308,I2690);
DFFARX1 I_29800 (I312321,I2683,I509308,I509334,);
not I_29801 (I509342,I509334);
nand I_29802 (I509359,I312324,I312300);
and I_29803 (I509376,I509359,I312297);
DFFARX1 I_29804 (I509376,I2683,I509308,I509402,);
not I_29805 (I509410,I312303);
DFFARX1 I_29806 (I312297,I2683,I509308,I509436,);
not I_29807 (I509444,I509436);
nor I_29808 (I509461,I509444,I509342);
and I_29809 (I509478,I509461,I312303);
nor I_29810 (I509495,I509444,I509410);
nor I_29811 (I509291,I509402,I509495);
DFFARX1 I_29812 (I312306,I2683,I509308,I509535,);
nor I_29813 (I509543,I509535,I509402);
not I_29814 (I509560,I509543);
not I_29815 (I509577,I509535);
nor I_29816 (I509594,I509577,I509478);
DFFARX1 I_29817 (I509594,I2683,I509308,I509294,);
nand I_29818 (I509625,I312309,I312318);
and I_29819 (I509642,I509625,I312315);
DFFARX1 I_29820 (I509642,I2683,I509308,I509668,);
nor I_29821 (I509676,I509668,I509535);
DFFARX1 I_29822 (I509676,I2683,I509308,I509276,);
nand I_29823 (I509707,I509668,I509577);
nand I_29824 (I509285,I509560,I509707);
not I_29825 (I509738,I509668);
nor I_29826 (I509755,I509738,I509478);
DFFARX1 I_29827 (I509755,I2683,I509308,I509297,);
nor I_29828 (I509786,I312312,I312318);
or I_29829 (I509288,I509535,I509786);
nor I_29830 (I509279,I509668,I509786);
or I_29831 (I509282,I509402,I509786);
DFFARX1 I_29832 (I509786,I2683,I509308,I509300,);
not I_29833 (I509886,I2690);
DFFARX1 I_29834 (I918960,I2683,I509886,I509912,);
not I_29835 (I509920,I509912);
nand I_29836 (I509937,I918942,I918954);
and I_29837 (I509954,I509937,I918957);
DFFARX1 I_29838 (I509954,I2683,I509886,I509980,);
not I_29839 (I509988,I918951);
DFFARX1 I_29840 (I918948,I2683,I509886,I510014,);
not I_29841 (I510022,I510014);
nor I_29842 (I510039,I510022,I509920);
and I_29843 (I510056,I510039,I918951);
nor I_29844 (I510073,I510022,I509988);
nor I_29845 (I509869,I509980,I510073);
DFFARX1 I_29846 (I918966,I2683,I509886,I510113,);
nor I_29847 (I510121,I510113,I509980);
not I_29848 (I510138,I510121);
not I_29849 (I510155,I510113);
nor I_29850 (I510172,I510155,I510056);
DFFARX1 I_29851 (I510172,I2683,I509886,I509872,);
nand I_29852 (I510203,I918945,I918945);
and I_29853 (I510220,I510203,I918942);
DFFARX1 I_29854 (I510220,I2683,I509886,I510246,);
nor I_29855 (I510254,I510246,I510113);
DFFARX1 I_29856 (I510254,I2683,I509886,I509854,);
nand I_29857 (I510285,I510246,I510155);
nand I_29858 (I509863,I510138,I510285);
not I_29859 (I510316,I510246);
nor I_29860 (I510333,I510316,I510056);
DFFARX1 I_29861 (I510333,I2683,I509886,I509875,);
nor I_29862 (I510364,I918963,I918945);
or I_29863 (I509866,I510113,I510364);
nor I_29864 (I509857,I510246,I510364);
or I_29865 (I509860,I509980,I510364);
DFFARX1 I_29866 (I510364,I2683,I509886,I509878,);
not I_29867 (I510464,I2690);
DFFARX1 I_29868 (I956478,I2683,I510464,I510490,);
not I_29869 (I510498,I510490);
nand I_29870 (I510515,I956481,I956490);
and I_29871 (I510532,I510515,I956493);
DFFARX1 I_29872 (I510532,I2683,I510464,I510558,);
not I_29873 (I510566,I956502);
DFFARX1 I_29874 (I956484,I2683,I510464,I510592,);
not I_29875 (I510600,I510592);
nor I_29876 (I510617,I510600,I510498);
and I_29877 (I510634,I510617,I956502);
nor I_29878 (I510651,I510600,I510566);
nor I_29879 (I510447,I510558,I510651);
DFFARX1 I_29880 (I956481,I2683,I510464,I510691,);
nor I_29881 (I510699,I510691,I510558);
not I_29882 (I510716,I510699);
not I_29883 (I510733,I510691);
nor I_29884 (I510750,I510733,I510634);
DFFARX1 I_29885 (I510750,I2683,I510464,I510450,);
nand I_29886 (I510781,I956499,I956478);
and I_29887 (I510798,I510781,I956496);
DFFARX1 I_29888 (I510798,I2683,I510464,I510824,);
nor I_29889 (I510832,I510824,I510691);
DFFARX1 I_29890 (I510832,I2683,I510464,I510432,);
nand I_29891 (I510863,I510824,I510733);
nand I_29892 (I510441,I510716,I510863);
not I_29893 (I510894,I510824);
nor I_29894 (I510911,I510894,I510634);
DFFARX1 I_29895 (I510911,I2683,I510464,I510453,);
nor I_29896 (I510942,I956487,I956478);
or I_29897 (I510444,I510691,I510942);
nor I_29898 (I510435,I510824,I510942);
or I_29899 (I510438,I510558,I510942);
DFFARX1 I_29900 (I510942,I2683,I510464,I510456,);
not I_29901 (I511042,I2690);
DFFARX1 I_29902 (I472862,I2683,I511042,I511068,);
not I_29903 (I511076,I511068);
nand I_29904 (I511093,I472871,I472880);
and I_29905 (I511110,I511093,I472886);
DFFARX1 I_29906 (I511110,I2683,I511042,I511136,);
not I_29907 (I511144,I472883);
DFFARX1 I_29908 (I472868,I2683,I511042,I511170,);
not I_29909 (I511178,I511170);
nor I_29910 (I511195,I511178,I511076);
and I_29911 (I511212,I511195,I472883);
nor I_29912 (I511229,I511178,I511144);
nor I_29913 (I511025,I511136,I511229);
DFFARX1 I_29914 (I472877,I2683,I511042,I511269,);
nor I_29915 (I511277,I511269,I511136);
not I_29916 (I511294,I511277);
not I_29917 (I511311,I511269);
nor I_29918 (I511328,I511311,I511212);
DFFARX1 I_29919 (I511328,I2683,I511042,I511028,);
nand I_29920 (I511359,I472874,I472865);
and I_29921 (I511376,I511359,I472862);
DFFARX1 I_29922 (I511376,I2683,I511042,I511402,);
nor I_29923 (I511410,I511402,I511269);
DFFARX1 I_29924 (I511410,I2683,I511042,I511010,);
nand I_29925 (I511441,I511402,I511311);
nand I_29926 (I511019,I511294,I511441);
not I_29927 (I511472,I511402);
nor I_29928 (I511489,I511472,I511212);
DFFARX1 I_29929 (I511489,I2683,I511042,I511031,);
nor I_29930 (I511520,I472865,I472865);
or I_29931 (I511022,I511269,I511520);
nor I_29932 (I511013,I511402,I511520);
or I_29933 (I511016,I511136,I511520);
DFFARX1 I_29934 (I511520,I2683,I511042,I511034,);
not I_29935 (I511620,I2690);
DFFARX1 I_29936 (I104373,I2683,I511620,I511646,);
not I_29937 (I511654,I511646);
nand I_29938 (I511671,I104382,I104391);
and I_29939 (I511688,I511671,I104370);
DFFARX1 I_29940 (I511688,I2683,I511620,I511714,);
not I_29941 (I511722,I104373);
DFFARX1 I_29942 (I104388,I2683,I511620,I511748,);
not I_29943 (I511756,I511748);
nor I_29944 (I511773,I511756,I511654);
and I_29945 (I511790,I511773,I104373);
nor I_29946 (I511807,I511756,I511722);
nor I_29947 (I511603,I511714,I511807);
DFFARX1 I_29948 (I104379,I2683,I511620,I511847,);
nor I_29949 (I511855,I511847,I511714);
not I_29950 (I511872,I511855);
not I_29951 (I511889,I511847);
nor I_29952 (I511906,I511889,I511790);
DFFARX1 I_29953 (I511906,I2683,I511620,I511606,);
nand I_29954 (I511937,I104394,I104370);
and I_29955 (I511954,I511937,I104376);
DFFARX1 I_29956 (I511954,I2683,I511620,I511980,);
nor I_29957 (I511988,I511980,I511847);
DFFARX1 I_29958 (I511988,I2683,I511620,I511588,);
nand I_29959 (I512019,I511980,I511889);
nand I_29960 (I511597,I511872,I512019);
not I_29961 (I512050,I511980);
nor I_29962 (I512067,I512050,I511790);
DFFARX1 I_29963 (I512067,I2683,I511620,I511609,);
nor I_29964 (I512098,I104385,I104370);
or I_29965 (I511600,I511847,I512098);
nor I_29966 (I511591,I511980,I512098);
or I_29967 (I511594,I511714,I512098);
DFFARX1 I_29968 (I512098,I2683,I511620,I511612,);
not I_29969 (I512198,I2690);
DFFARX1 I_29970 (I279647,I2683,I512198,I512224,);
not I_29971 (I512232,I512224);
nand I_29972 (I512249,I279650,I279626);
and I_29973 (I512266,I512249,I279623);
DFFARX1 I_29974 (I512266,I2683,I512198,I512292,);
not I_29975 (I512300,I279629);
DFFARX1 I_29976 (I279623,I2683,I512198,I512326,);
not I_29977 (I512334,I512326);
nor I_29978 (I512351,I512334,I512232);
and I_29979 (I512368,I512351,I279629);
nor I_29980 (I512385,I512334,I512300);
nor I_29981 (I512181,I512292,I512385);
DFFARX1 I_29982 (I279632,I2683,I512198,I512425,);
nor I_29983 (I512433,I512425,I512292);
not I_29984 (I512450,I512433);
not I_29985 (I512467,I512425);
nor I_29986 (I512484,I512467,I512368);
DFFARX1 I_29987 (I512484,I2683,I512198,I512184,);
nand I_29988 (I512515,I279635,I279644);
and I_29989 (I512532,I512515,I279641);
DFFARX1 I_29990 (I512532,I2683,I512198,I512558,);
nor I_29991 (I512566,I512558,I512425);
DFFARX1 I_29992 (I512566,I2683,I512198,I512166,);
nand I_29993 (I512597,I512558,I512467);
nand I_29994 (I512175,I512450,I512597);
not I_29995 (I512628,I512558);
nor I_29996 (I512645,I512628,I512368);
DFFARX1 I_29997 (I512645,I2683,I512198,I512187,);
nor I_29998 (I512676,I279638,I279644);
or I_29999 (I512178,I512425,I512676);
nor I_30000 (I512169,I512558,I512676);
or I_30001 (I512172,I512292,I512676);
DFFARX1 I_30002 (I512676,I2683,I512198,I512190,);
not I_30003 (I512776,I2690);
DFFARX1 I_30004 (I52200,I2683,I512776,I512802,);
not I_30005 (I512810,I512802);
nand I_30006 (I512827,I52209,I52218);
and I_30007 (I512844,I512827,I52197);
DFFARX1 I_30008 (I512844,I2683,I512776,I512870,);
not I_30009 (I512878,I52200);
DFFARX1 I_30010 (I52215,I2683,I512776,I512904,);
not I_30011 (I512912,I512904);
nor I_30012 (I512929,I512912,I512810);
and I_30013 (I512946,I512929,I52200);
nor I_30014 (I512963,I512912,I512878);
nor I_30015 (I512759,I512870,I512963);
DFFARX1 I_30016 (I52206,I2683,I512776,I513003,);
nor I_30017 (I513011,I513003,I512870);
not I_30018 (I513028,I513011);
not I_30019 (I513045,I513003);
nor I_30020 (I513062,I513045,I512946);
DFFARX1 I_30021 (I513062,I2683,I512776,I512762,);
nand I_30022 (I513093,I52221,I52197);
and I_30023 (I513110,I513093,I52203);
DFFARX1 I_30024 (I513110,I2683,I512776,I513136,);
nor I_30025 (I513144,I513136,I513003);
DFFARX1 I_30026 (I513144,I2683,I512776,I512744,);
nand I_30027 (I513175,I513136,I513045);
nand I_30028 (I512753,I513028,I513175);
not I_30029 (I513206,I513136);
nor I_30030 (I513223,I513206,I512946);
DFFARX1 I_30031 (I513223,I2683,I512776,I512765,);
nor I_30032 (I513254,I52212,I52197);
or I_30033 (I512756,I513003,I513254);
nor I_30034 (I512747,I513136,I513254);
or I_30035 (I512750,I512870,I513254);
DFFARX1 I_30036 (I513254,I2683,I512776,I512768,);
not I_30037 (I513354,I2690);
DFFARX1 I_30038 (I235906,I2683,I513354,I513380,);
not I_30039 (I513388,I513380);
nand I_30040 (I513405,I235909,I235885);
and I_30041 (I513422,I513405,I235882);
DFFARX1 I_30042 (I513422,I2683,I513354,I513448,);
not I_30043 (I513456,I235888);
DFFARX1 I_30044 (I235882,I2683,I513354,I513482,);
not I_30045 (I513490,I513482);
nor I_30046 (I513507,I513490,I513388);
and I_30047 (I513524,I513507,I235888);
nor I_30048 (I513541,I513490,I513456);
nor I_30049 (I513337,I513448,I513541);
DFFARX1 I_30050 (I235891,I2683,I513354,I513581,);
nor I_30051 (I513589,I513581,I513448);
not I_30052 (I513606,I513589);
not I_30053 (I513623,I513581);
nor I_30054 (I513640,I513623,I513524);
DFFARX1 I_30055 (I513640,I2683,I513354,I513340,);
nand I_30056 (I513671,I235894,I235903);
and I_30057 (I513688,I513671,I235900);
DFFARX1 I_30058 (I513688,I2683,I513354,I513714,);
nor I_30059 (I513722,I513714,I513581);
DFFARX1 I_30060 (I513722,I2683,I513354,I513322,);
nand I_30061 (I513753,I513714,I513623);
nand I_30062 (I513331,I513606,I513753);
not I_30063 (I513784,I513714);
nor I_30064 (I513801,I513784,I513524);
DFFARX1 I_30065 (I513801,I2683,I513354,I513343,);
nor I_30066 (I513832,I235897,I235903);
or I_30067 (I513334,I513581,I513832);
nor I_30068 (I513325,I513714,I513832);
or I_30069 (I513328,I513448,I513832);
DFFARX1 I_30070 (I513832,I2683,I513354,I513346,);
not I_30071 (I513932,I2690);
DFFARX1 I_30072 (I80658,I2683,I513932,I513958,);
not I_30073 (I513966,I513958);
nand I_30074 (I513983,I80667,I80676);
and I_30075 (I514000,I513983,I80655);
DFFARX1 I_30076 (I514000,I2683,I513932,I514026,);
not I_30077 (I514034,I80658);
DFFARX1 I_30078 (I80673,I2683,I513932,I514060,);
not I_30079 (I514068,I514060);
nor I_30080 (I514085,I514068,I513966);
and I_30081 (I514102,I514085,I80658);
nor I_30082 (I514119,I514068,I514034);
nor I_30083 (I513915,I514026,I514119);
DFFARX1 I_30084 (I80664,I2683,I513932,I514159,);
nor I_30085 (I514167,I514159,I514026);
not I_30086 (I514184,I514167);
not I_30087 (I514201,I514159);
nor I_30088 (I514218,I514201,I514102);
DFFARX1 I_30089 (I514218,I2683,I513932,I513918,);
nand I_30090 (I514249,I80679,I80655);
and I_30091 (I514266,I514249,I80661);
DFFARX1 I_30092 (I514266,I2683,I513932,I514292,);
nor I_30093 (I514300,I514292,I514159);
DFFARX1 I_30094 (I514300,I2683,I513932,I513900,);
nand I_30095 (I514331,I514292,I514201);
nand I_30096 (I513909,I514184,I514331);
not I_30097 (I514362,I514292);
nor I_30098 (I514379,I514362,I514102);
DFFARX1 I_30099 (I514379,I2683,I513932,I513921,);
nor I_30100 (I514410,I80670,I80655);
or I_30101 (I513912,I514159,I514410);
nor I_30102 (I513903,I514292,I514410);
or I_30103 (I513906,I514026,I514410);
DFFARX1 I_30104 (I514410,I2683,I513932,I513924,);
not I_30105 (I514510,I2690);
DFFARX1 I_30106 (I378011,I2683,I514510,I514536,);
not I_30107 (I514544,I514536);
nand I_30108 (I514561,I378002,I378020);
and I_30109 (I514578,I514561,I378023);
DFFARX1 I_30110 (I514578,I2683,I514510,I514604,);
not I_30111 (I514612,I378017);
DFFARX1 I_30112 (I378005,I2683,I514510,I514638,);
not I_30113 (I514646,I514638);
nor I_30114 (I514663,I514646,I514544);
and I_30115 (I514680,I514663,I378017);
nor I_30116 (I514697,I514646,I514612);
nor I_30117 (I514493,I514604,I514697);
DFFARX1 I_30118 (I378014,I2683,I514510,I514737,);
nor I_30119 (I514745,I514737,I514604);
not I_30120 (I514762,I514745);
not I_30121 (I514779,I514737);
nor I_30122 (I514796,I514779,I514680);
DFFARX1 I_30123 (I514796,I2683,I514510,I514496,);
nand I_30124 (I514827,I378029,I378026);
and I_30125 (I514844,I514827,I378008);
DFFARX1 I_30126 (I514844,I2683,I514510,I514870,);
nor I_30127 (I514878,I514870,I514737);
DFFARX1 I_30128 (I514878,I2683,I514510,I514478,);
nand I_30129 (I514909,I514870,I514779);
nand I_30130 (I514487,I514762,I514909);
not I_30131 (I514940,I514870);
nor I_30132 (I514957,I514940,I514680);
DFFARX1 I_30133 (I514957,I2683,I514510,I514499,);
nor I_30134 (I514988,I378002,I378026);
or I_30135 (I514490,I514737,I514988);
nor I_30136 (I514481,I514870,I514988);
or I_30137 (I514484,I514604,I514988);
DFFARX1 I_30138 (I514988,I2683,I514510,I514502,);
not I_30139 (I515088,I2690);
DFFARX1 I_30140 (I830526,I2683,I515088,I515114,);
not I_30141 (I515122,I515114);
nand I_30142 (I515139,I830508,I830520);
and I_30143 (I515156,I515139,I830523);
DFFARX1 I_30144 (I515156,I2683,I515088,I515182,);
not I_30145 (I515190,I830517);
DFFARX1 I_30146 (I830514,I2683,I515088,I515216,);
not I_30147 (I515224,I515216);
nor I_30148 (I515241,I515224,I515122);
and I_30149 (I515258,I515241,I830517);
nor I_30150 (I515275,I515224,I515190);
nor I_30151 (I515071,I515182,I515275);
DFFARX1 I_30152 (I830532,I2683,I515088,I515315,);
nor I_30153 (I515323,I515315,I515182);
not I_30154 (I515340,I515323);
not I_30155 (I515357,I515315);
nor I_30156 (I515374,I515357,I515258);
DFFARX1 I_30157 (I515374,I2683,I515088,I515074,);
nand I_30158 (I515405,I830511,I830511);
and I_30159 (I515422,I515405,I830508);
DFFARX1 I_30160 (I515422,I2683,I515088,I515448,);
nor I_30161 (I515456,I515448,I515315);
DFFARX1 I_30162 (I515456,I2683,I515088,I515056,);
nand I_30163 (I515487,I515448,I515357);
nand I_30164 (I515065,I515340,I515487);
not I_30165 (I515518,I515448);
nor I_30166 (I515535,I515518,I515258);
DFFARX1 I_30167 (I515535,I2683,I515088,I515077,);
nor I_30168 (I515566,I830529,I830511);
or I_30169 (I515068,I515315,I515566);
nor I_30170 (I515059,I515448,I515566);
or I_30171 (I515062,I515182,I515566);
DFFARX1 I_30172 (I515566,I2683,I515088,I515080,);
not I_30173 (I515666,I2690);
DFFARX1 I_30174 (I1094171,I2683,I515666,I515692,);
not I_30175 (I515700,I515692);
nand I_30176 (I515717,I1094156,I1094144);
and I_30177 (I515734,I515717,I1094159);
DFFARX1 I_30178 (I515734,I2683,I515666,I515760,);
not I_30179 (I515768,I1094144);
DFFARX1 I_30180 (I1094162,I2683,I515666,I515794,);
not I_30181 (I515802,I515794);
nor I_30182 (I515819,I515802,I515700);
and I_30183 (I515836,I515819,I1094144);
nor I_30184 (I515853,I515802,I515768);
nor I_30185 (I515649,I515760,I515853);
DFFARX1 I_30186 (I1094150,I2683,I515666,I515893,);
nor I_30187 (I515901,I515893,I515760);
not I_30188 (I515918,I515901);
not I_30189 (I515935,I515893);
nor I_30190 (I515952,I515935,I515836);
DFFARX1 I_30191 (I515952,I2683,I515666,I515652,);
nand I_30192 (I515983,I1094147,I1094153);
and I_30193 (I516000,I515983,I1094168);
DFFARX1 I_30194 (I516000,I2683,I515666,I516026,);
nor I_30195 (I516034,I516026,I515893);
DFFARX1 I_30196 (I516034,I2683,I515666,I515634,);
nand I_30197 (I516065,I516026,I515935);
nand I_30198 (I515643,I515918,I516065);
not I_30199 (I516096,I516026);
nor I_30200 (I516113,I516096,I515836);
DFFARX1 I_30201 (I516113,I2683,I515666,I515655,);
nor I_30202 (I516144,I1094165,I1094153);
or I_30203 (I515646,I515893,I516144);
nor I_30204 (I515637,I516026,I516144);
or I_30205 (I515640,I515760,I516144);
DFFARX1 I_30206 (I516144,I2683,I515666,I515658,);
not I_30207 (I516244,I2690);
DFFARX1 I_30208 (I454366,I2683,I516244,I516270,);
not I_30209 (I516278,I516270);
nand I_30210 (I516295,I454375,I454384);
and I_30211 (I516312,I516295,I454390);
DFFARX1 I_30212 (I516312,I2683,I516244,I516338,);
not I_30213 (I516346,I454387);
DFFARX1 I_30214 (I454372,I2683,I516244,I516372,);
not I_30215 (I516380,I516372);
nor I_30216 (I516397,I516380,I516278);
and I_30217 (I516414,I516397,I454387);
nor I_30218 (I516431,I516380,I516346);
nor I_30219 (I516227,I516338,I516431);
DFFARX1 I_30220 (I454381,I2683,I516244,I516471,);
nor I_30221 (I516479,I516471,I516338);
not I_30222 (I516496,I516479);
not I_30223 (I516513,I516471);
nor I_30224 (I516530,I516513,I516414);
DFFARX1 I_30225 (I516530,I2683,I516244,I516230,);
nand I_30226 (I516561,I454378,I454369);
and I_30227 (I516578,I516561,I454366);
DFFARX1 I_30228 (I516578,I2683,I516244,I516604,);
nor I_30229 (I516612,I516604,I516471);
DFFARX1 I_30230 (I516612,I2683,I516244,I516212,);
nand I_30231 (I516643,I516604,I516513);
nand I_30232 (I516221,I516496,I516643);
not I_30233 (I516674,I516604);
nor I_30234 (I516691,I516674,I516414);
DFFARX1 I_30235 (I516691,I2683,I516244,I516233,);
nor I_30236 (I516722,I454369,I454369);
or I_30237 (I516224,I516471,I516722);
nor I_30238 (I516215,I516604,I516722);
or I_30239 (I516218,I516338,I516722);
DFFARX1 I_30240 (I516722,I2683,I516244,I516236,);
not I_30241 (I516822,I2690);
DFFARX1 I_30242 (I643353,I2683,I516822,I516848,);
not I_30243 (I516856,I516848);
nand I_30244 (I516873,I643341,I643359);
and I_30245 (I516890,I516873,I643356);
DFFARX1 I_30246 (I516890,I2683,I516822,I516916,);
not I_30247 (I516924,I643347);
DFFARX1 I_30248 (I643344,I2683,I516822,I516950,);
not I_30249 (I516958,I516950);
nor I_30250 (I516975,I516958,I516856);
and I_30251 (I516992,I516975,I643347);
nor I_30252 (I517009,I516958,I516924);
nor I_30253 (I516805,I516916,I517009);
DFFARX1 I_30254 (I643338,I2683,I516822,I517049,);
nor I_30255 (I517057,I517049,I516916);
not I_30256 (I517074,I517057);
not I_30257 (I517091,I517049);
nor I_30258 (I517108,I517091,I516992);
DFFARX1 I_30259 (I517108,I2683,I516822,I516808,);
nand I_30260 (I517139,I643338,I643341);
and I_30261 (I517156,I517139,I643344);
DFFARX1 I_30262 (I517156,I2683,I516822,I517182,);
nor I_30263 (I517190,I517182,I517049);
DFFARX1 I_30264 (I517190,I2683,I516822,I516790,);
nand I_30265 (I517221,I517182,I517091);
nand I_30266 (I516799,I517074,I517221);
not I_30267 (I517252,I517182);
nor I_30268 (I517269,I517252,I516992);
DFFARX1 I_30269 (I517269,I2683,I516822,I516811,);
nor I_30270 (I517300,I643350,I643341);
or I_30271 (I516802,I517049,I517300);
nor I_30272 (I516793,I517182,I517300);
or I_30273 (I516796,I516916,I517300);
DFFARX1 I_30274 (I517300,I2683,I516822,I516814,);
not I_30275 (I517400,I2690);
DFFARX1 I_30276 (I757483,I2683,I517400,I517426,);
not I_30277 (I517434,I517426);
nand I_30278 (I517451,I757459,I757474);
and I_30279 (I517468,I517451,I757486);
DFFARX1 I_30280 (I517468,I2683,I517400,I517494,);
not I_30281 (I517502,I757471);
DFFARX1 I_30282 (I757462,I2683,I517400,I517528,);
not I_30283 (I517536,I517528);
nor I_30284 (I517553,I517536,I517434);
and I_30285 (I517570,I517553,I757471);
nor I_30286 (I517587,I517536,I517502);
nor I_30287 (I517383,I517494,I517587);
DFFARX1 I_30288 (I757459,I2683,I517400,I517627,);
nor I_30289 (I517635,I517627,I517494);
not I_30290 (I517652,I517635);
not I_30291 (I517669,I517627);
nor I_30292 (I517686,I517669,I517570);
DFFARX1 I_30293 (I517686,I2683,I517400,I517386,);
nand I_30294 (I517717,I757477,I757468);
and I_30295 (I517734,I517717,I757480);
DFFARX1 I_30296 (I517734,I2683,I517400,I517760,);
nor I_30297 (I517768,I517760,I517627);
DFFARX1 I_30298 (I517768,I2683,I517400,I517368,);
nand I_30299 (I517799,I517760,I517669);
nand I_30300 (I517377,I517652,I517799);
not I_30301 (I517830,I517760);
nor I_30302 (I517847,I517830,I517570);
DFFARX1 I_30303 (I517847,I2683,I517400,I517389,);
nor I_30304 (I517878,I757465,I757468);
or I_30305 (I517380,I517627,I517878);
nor I_30306 (I517371,I517760,I517878);
or I_30307 (I517374,I517494,I517878);
DFFARX1 I_30308 (I517878,I2683,I517400,I517392,);
not I_30309 (I517978,I2690);
DFFARX1 I_30310 (I930520,I2683,I517978,I518004,);
not I_30311 (I518012,I518004);
nand I_30312 (I518029,I930502,I930514);
and I_30313 (I518046,I518029,I930517);
DFFARX1 I_30314 (I518046,I2683,I517978,I518072,);
not I_30315 (I518080,I930511);
DFFARX1 I_30316 (I930508,I2683,I517978,I518106,);
not I_30317 (I518114,I518106);
nor I_30318 (I518131,I518114,I518012);
and I_30319 (I518148,I518131,I930511);
nor I_30320 (I518165,I518114,I518080);
nor I_30321 (I517961,I518072,I518165);
DFFARX1 I_30322 (I930526,I2683,I517978,I518205,);
nor I_30323 (I518213,I518205,I518072);
not I_30324 (I518230,I518213);
not I_30325 (I518247,I518205);
nor I_30326 (I518264,I518247,I518148);
DFFARX1 I_30327 (I518264,I2683,I517978,I517964,);
nand I_30328 (I518295,I930505,I930505);
and I_30329 (I518312,I518295,I930502);
DFFARX1 I_30330 (I518312,I2683,I517978,I518338,);
nor I_30331 (I518346,I518338,I518205);
DFFARX1 I_30332 (I518346,I2683,I517978,I517946,);
nand I_30333 (I518377,I518338,I518247);
nand I_30334 (I517955,I518230,I518377);
not I_30335 (I518408,I518338);
nor I_30336 (I518425,I518408,I518148);
DFFARX1 I_30337 (I518425,I2683,I517978,I517967,);
nor I_30338 (I518456,I930523,I930505);
or I_30339 (I517958,I518205,I518456);
nor I_30340 (I517949,I518338,I518456);
or I_30341 (I517952,I518072,I518456);
DFFARX1 I_30342 (I518456,I2683,I517978,I517970,);
not I_30343 (I518556,I2690);
DFFARX1 I_30344 (I468238,I2683,I518556,I518582,);
not I_30345 (I518590,I518582);
nand I_30346 (I518607,I468247,I468256);
and I_30347 (I518624,I518607,I468262);
DFFARX1 I_30348 (I518624,I2683,I518556,I518650,);
not I_30349 (I518658,I468259);
DFFARX1 I_30350 (I468244,I2683,I518556,I518684,);
not I_30351 (I518692,I518684);
nor I_30352 (I518709,I518692,I518590);
and I_30353 (I518726,I518709,I468259);
nor I_30354 (I518743,I518692,I518658);
nor I_30355 (I518539,I518650,I518743);
DFFARX1 I_30356 (I468253,I2683,I518556,I518783,);
nor I_30357 (I518791,I518783,I518650);
not I_30358 (I518808,I518791);
not I_30359 (I518825,I518783);
nor I_30360 (I518842,I518825,I518726);
DFFARX1 I_30361 (I518842,I2683,I518556,I518542,);
nand I_30362 (I518873,I468250,I468241);
and I_30363 (I518890,I518873,I468238);
DFFARX1 I_30364 (I518890,I2683,I518556,I518916,);
nor I_30365 (I518924,I518916,I518783);
DFFARX1 I_30366 (I518924,I2683,I518556,I518524,);
nand I_30367 (I518955,I518916,I518825);
nand I_30368 (I518533,I518808,I518955);
not I_30369 (I518986,I518916);
nor I_30370 (I519003,I518986,I518726);
DFFARX1 I_30371 (I519003,I2683,I518556,I518545,);
nor I_30372 (I519034,I468241,I468241);
or I_30373 (I518536,I518783,I519034);
nor I_30374 (I518527,I518916,I519034);
or I_30375 (I518530,I518650,I519034);
DFFARX1 I_30376 (I519034,I2683,I518556,I518548,);
not I_30377 (I519134,I2690);
DFFARX1 I_30378 (I164635,I2683,I519134,I519160,);
not I_30379 (I519168,I519160);
nand I_30380 (I519185,I164638,I164659);
and I_30381 (I519202,I519185,I164647);
DFFARX1 I_30382 (I519202,I2683,I519134,I519228,);
not I_30383 (I519236,I164644);
DFFARX1 I_30384 (I164635,I2683,I519134,I519262,);
not I_30385 (I519270,I519262);
nor I_30386 (I519287,I519270,I519168);
and I_30387 (I519304,I519287,I164644);
nor I_30388 (I519321,I519270,I519236);
nor I_30389 (I519117,I519228,I519321);
DFFARX1 I_30390 (I164653,I2683,I519134,I519361,);
nor I_30391 (I519369,I519361,I519228);
not I_30392 (I519386,I519369);
not I_30393 (I519403,I519361);
nor I_30394 (I519420,I519403,I519304);
DFFARX1 I_30395 (I519420,I2683,I519134,I519120,);
nand I_30396 (I519451,I164638,I164641);
and I_30397 (I519468,I519451,I164650);
DFFARX1 I_30398 (I519468,I2683,I519134,I519494,);
nor I_30399 (I519502,I519494,I519361);
DFFARX1 I_30400 (I519502,I2683,I519134,I519102,);
nand I_30401 (I519533,I519494,I519403);
nand I_30402 (I519111,I519386,I519533);
not I_30403 (I519564,I519494);
nor I_30404 (I519581,I519564,I519304);
DFFARX1 I_30405 (I519581,I2683,I519134,I519123,);
nor I_30406 (I519612,I164656,I164641);
or I_30407 (I519114,I519361,I519612);
nor I_30408 (I519105,I519494,I519612);
or I_30409 (I519108,I519228,I519612);
DFFARX1 I_30410 (I519612,I2683,I519134,I519126,);
not I_30411 (I519712,I2690);
DFFARX1 I_30412 (I758775,I2683,I519712,I519738,);
not I_30413 (I519746,I519738);
nand I_30414 (I519763,I758751,I758766);
and I_30415 (I519780,I519763,I758778);
DFFARX1 I_30416 (I519780,I2683,I519712,I519806,);
not I_30417 (I519814,I758763);
DFFARX1 I_30418 (I758754,I2683,I519712,I519840,);
not I_30419 (I519848,I519840);
nor I_30420 (I519865,I519848,I519746);
and I_30421 (I519882,I519865,I758763);
nor I_30422 (I519899,I519848,I519814);
nor I_30423 (I519695,I519806,I519899);
DFFARX1 I_30424 (I758751,I2683,I519712,I519939,);
nor I_30425 (I519947,I519939,I519806);
not I_30426 (I519964,I519947);
not I_30427 (I519981,I519939);
nor I_30428 (I519998,I519981,I519882);
DFFARX1 I_30429 (I519998,I2683,I519712,I519698,);
nand I_30430 (I520029,I758769,I758760);
and I_30431 (I520046,I520029,I758772);
DFFARX1 I_30432 (I520046,I2683,I519712,I520072,);
nor I_30433 (I520080,I520072,I519939);
DFFARX1 I_30434 (I520080,I2683,I519712,I519680,);
nand I_30435 (I520111,I520072,I519981);
nand I_30436 (I519689,I519964,I520111);
not I_30437 (I520142,I520072);
nor I_30438 (I520159,I520142,I519882);
DFFARX1 I_30439 (I520159,I2683,I519712,I519701,);
nor I_30440 (I520190,I758757,I758760);
or I_30441 (I519692,I519939,I520190);
nor I_30442 (I519683,I520072,I520190);
or I_30443 (I519686,I519806,I520190);
DFFARX1 I_30444 (I520190,I2683,I519712,I519704,);
not I_30445 (I520290,I2690);
DFFARX1 I_30446 (I98049,I2683,I520290,I520316,);
not I_30447 (I520324,I520316);
nand I_30448 (I520341,I98058,I98067);
and I_30449 (I520358,I520341,I98046);
DFFARX1 I_30450 (I520358,I2683,I520290,I520384,);
not I_30451 (I520392,I98049);
DFFARX1 I_30452 (I98064,I2683,I520290,I520418,);
not I_30453 (I520426,I520418);
nor I_30454 (I520443,I520426,I520324);
and I_30455 (I520460,I520443,I98049);
nor I_30456 (I520477,I520426,I520392);
nor I_30457 (I520273,I520384,I520477);
DFFARX1 I_30458 (I98055,I2683,I520290,I520517,);
nor I_30459 (I520525,I520517,I520384);
not I_30460 (I520542,I520525);
not I_30461 (I520559,I520517);
nor I_30462 (I520576,I520559,I520460);
DFFARX1 I_30463 (I520576,I2683,I520290,I520276,);
nand I_30464 (I520607,I98070,I98046);
and I_30465 (I520624,I520607,I98052);
DFFARX1 I_30466 (I520624,I2683,I520290,I520650,);
nor I_30467 (I520658,I520650,I520517);
DFFARX1 I_30468 (I520658,I2683,I520290,I520258,);
nand I_30469 (I520689,I520650,I520559);
nand I_30470 (I520267,I520542,I520689);
not I_30471 (I520720,I520650);
nor I_30472 (I520737,I520720,I520460);
DFFARX1 I_30473 (I520737,I2683,I520290,I520279,);
nor I_30474 (I520768,I98061,I98046);
or I_30475 (I520270,I520517,I520768);
nor I_30476 (I520261,I520650,I520768);
or I_30477 (I520264,I520384,I520768);
DFFARX1 I_30478 (I520768,I2683,I520290,I520282,);
not I_30479 (I520868,I2690);
DFFARX1 I_30480 (I366043,I2683,I520868,I520894,);
not I_30481 (I520902,I520894);
nand I_30482 (I520919,I366034,I366052);
and I_30483 (I520936,I520919,I366055);
DFFARX1 I_30484 (I520936,I2683,I520868,I520962,);
not I_30485 (I520970,I366049);
DFFARX1 I_30486 (I366037,I2683,I520868,I520996,);
not I_30487 (I521004,I520996);
nor I_30488 (I521021,I521004,I520902);
and I_30489 (I521038,I521021,I366049);
nor I_30490 (I521055,I521004,I520970);
nor I_30491 (I520851,I520962,I521055);
DFFARX1 I_30492 (I366046,I2683,I520868,I521095,);
nor I_30493 (I521103,I521095,I520962);
not I_30494 (I521120,I521103);
not I_30495 (I521137,I521095);
nor I_30496 (I521154,I521137,I521038);
DFFARX1 I_30497 (I521154,I2683,I520868,I520854,);
nand I_30498 (I521185,I366061,I366058);
and I_30499 (I521202,I521185,I366040);
DFFARX1 I_30500 (I521202,I2683,I520868,I521228,);
nor I_30501 (I521236,I521228,I521095);
DFFARX1 I_30502 (I521236,I2683,I520868,I520836,);
nand I_30503 (I521267,I521228,I521137);
nand I_30504 (I520845,I521120,I521267);
not I_30505 (I521298,I521228);
nor I_30506 (I521315,I521298,I521038);
DFFARX1 I_30507 (I521315,I2683,I520868,I520857,);
nor I_30508 (I521346,I366034,I366058);
or I_30509 (I520848,I521095,I521346);
nor I_30510 (I520839,I521228,I521346);
or I_30511 (I520842,I520962,I521346);
DFFARX1 I_30512 (I521346,I2683,I520868,I520860,);
not I_30513 (I521446,I2690);
DFFARX1 I_30514 (I842086,I2683,I521446,I521472,);
not I_30515 (I521480,I521472);
nand I_30516 (I521497,I842068,I842080);
and I_30517 (I521514,I521497,I842083);
DFFARX1 I_30518 (I521514,I2683,I521446,I521540,);
not I_30519 (I521548,I842077);
DFFARX1 I_30520 (I842074,I2683,I521446,I521574,);
not I_30521 (I521582,I521574);
nor I_30522 (I521599,I521582,I521480);
and I_30523 (I521616,I521599,I842077);
nor I_30524 (I521633,I521582,I521548);
nor I_30525 (I521429,I521540,I521633);
DFFARX1 I_30526 (I842092,I2683,I521446,I521673,);
nor I_30527 (I521681,I521673,I521540);
not I_30528 (I521698,I521681);
not I_30529 (I521715,I521673);
nor I_30530 (I521732,I521715,I521616);
DFFARX1 I_30531 (I521732,I2683,I521446,I521432,);
nand I_30532 (I521763,I842071,I842071);
and I_30533 (I521780,I521763,I842068);
DFFARX1 I_30534 (I521780,I2683,I521446,I521806,);
nor I_30535 (I521814,I521806,I521673);
DFFARX1 I_30536 (I521814,I2683,I521446,I521414,);
nand I_30537 (I521845,I521806,I521715);
nand I_30538 (I521423,I521698,I521845);
not I_30539 (I521876,I521806);
nor I_30540 (I521893,I521876,I521616);
DFFARX1 I_30541 (I521893,I2683,I521446,I521435,);
nor I_30542 (I521924,I842089,I842071);
or I_30543 (I521426,I521673,I521924);
nor I_30544 (I521417,I521806,I521924);
or I_30545 (I521420,I521540,I521924);
DFFARX1 I_30546 (I521924,I2683,I521446,I521438,);
not I_30547 (I522024,I2690);
DFFARX1 I_30548 (I932832,I2683,I522024,I522050,);
not I_30549 (I522058,I522050);
nand I_30550 (I522075,I932814,I932826);
and I_30551 (I522092,I522075,I932829);
DFFARX1 I_30552 (I522092,I2683,I522024,I522118,);
not I_30553 (I522126,I932823);
DFFARX1 I_30554 (I932820,I2683,I522024,I522152,);
not I_30555 (I522160,I522152);
nor I_30556 (I522177,I522160,I522058);
and I_30557 (I522194,I522177,I932823);
nor I_30558 (I522211,I522160,I522126);
nor I_30559 (I522007,I522118,I522211);
DFFARX1 I_30560 (I932838,I2683,I522024,I522251,);
nor I_30561 (I522259,I522251,I522118);
not I_30562 (I522276,I522259);
not I_30563 (I522293,I522251);
nor I_30564 (I522310,I522293,I522194);
DFFARX1 I_30565 (I522310,I2683,I522024,I522010,);
nand I_30566 (I522341,I932817,I932817);
and I_30567 (I522358,I522341,I932814);
DFFARX1 I_30568 (I522358,I2683,I522024,I522384,);
nor I_30569 (I522392,I522384,I522251);
DFFARX1 I_30570 (I522392,I2683,I522024,I521992,);
nand I_30571 (I522423,I522384,I522293);
nand I_30572 (I522001,I522276,I522423);
not I_30573 (I522454,I522384);
nor I_30574 (I522471,I522454,I522194);
DFFARX1 I_30575 (I522471,I2683,I522024,I522013,);
nor I_30576 (I522502,I932835,I932817);
or I_30577 (I522004,I522251,I522502);
nor I_30578 (I521995,I522384,I522502);
or I_30579 (I521998,I522118,I522502);
DFFARX1 I_30580 (I522502,I2683,I522024,I522016,);
not I_30581 (I522602,I2690);
DFFARX1 I_30582 (I222204,I2683,I522602,I522628,);
not I_30583 (I522636,I522628);
nand I_30584 (I522653,I222207,I222183);
and I_30585 (I522670,I522653,I222180);
DFFARX1 I_30586 (I522670,I2683,I522602,I522696,);
not I_30587 (I522704,I222186);
DFFARX1 I_30588 (I222180,I2683,I522602,I522730,);
not I_30589 (I522738,I522730);
nor I_30590 (I522755,I522738,I522636);
and I_30591 (I522772,I522755,I222186);
nor I_30592 (I522789,I522738,I522704);
nor I_30593 (I522585,I522696,I522789);
DFFARX1 I_30594 (I222189,I2683,I522602,I522829,);
nor I_30595 (I522837,I522829,I522696);
not I_30596 (I522854,I522837);
not I_30597 (I522871,I522829);
nor I_30598 (I522888,I522871,I522772);
DFFARX1 I_30599 (I522888,I2683,I522602,I522588,);
nand I_30600 (I522919,I222192,I222201);
and I_30601 (I522936,I522919,I222198);
DFFARX1 I_30602 (I522936,I2683,I522602,I522962,);
nor I_30603 (I522970,I522962,I522829);
DFFARX1 I_30604 (I522970,I2683,I522602,I522570,);
nand I_30605 (I523001,I522962,I522871);
nand I_30606 (I522579,I522854,I523001);
not I_30607 (I523032,I522962);
nor I_30608 (I523049,I523032,I522772);
DFFARX1 I_30609 (I523049,I2683,I522602,I522591,);
nor I_30610 (I523080,I222195,I222201);
or I_30611 (I522582,I522829,I523080);
nor I_30612 (I522573,I522962,I523080);
or I_30613 (I522576,I522696,I523080);
DFFARX1 I_30614 (I523080,I2683,I522602,I522594,);
not I_30615 (I523180,I2690);
DFFARX1 I_30616 (I460146,I2683,I523180,I523206,);
not I_30617 (I523214,I523206);
nand I_30618 (I523231,I460155,I460164);
and I_30619 (I523248,I523231,I460170);
DFFARX1 I_30620 (I523248,I2683,I523180,I523274,);
not I_30621 (I523282,I460167);
DFFARX1 I_30622 (I460152,I2683,I523180,I523308,);
not I_30623 (I523316,I523308);
nor I_30624 (I523333,I523316,I523214);
and I_30625 (I523350,I523333,I460167);
nor I_30626 (I523367,I523316,I523282);
nor I_30627 (I523163,I523274,I523367);
DFFARX1 I_30628 (I460161,I2683,I523180,I523407,);
nor I_30629 (I523415,I523407,I523274);
not I_30630 (I523432,I523415);
not I_30631 (I523449,I523407);
nor I_30632 (I523466,I523449,I523350);
DFFARX1 I_30633 (I523466,I2683,I523180,I523166,);
nand I_30634 (I523497,I460158,I460149);
and I_30635 (I523514,I523497,I460146);
DFFARX1 I_30636 (I523514,I2683,I523180,I523540,);
nor I_30637 (I523548,I523540,I523407);
DFFARX1 I_30638 (I523548,I2683,I523180,I523148,);
nand I_30639 (I523579,I523540,I523449);
nand I_30640 (I523157,I523432,I523579);
not I_30641 (I523610,I523540);
nor I_30642 (I523627,I523610,I523350);
DFFARX1 I_30643 (I523627,I2683,I523180,I523169,);
nor I_30644 (I523658,I460149,I460149);
or I_30645 (I523160,I523407,I523658);
nor I_30646 (I523151,I523540,I523658);
or I_30647 (I523154,I523274,I523658);
DFFARX1 I_30648 (I523658,I2683,I523180,I523172,);
not I_30649 (I523758,I2690);
DFFARX1 I_30650 (I653893,I2683,I523758,I523784,);
not I_30651 (I523792,I523784);
nand I_30652 (I523809,I653881,I653899);
and I_30653 (I523826,I523809,I653896);
DFFARX1 I_30654 (I523826,I2683,I523758,I523852,);
not I_30655 (I523860,I653887);
DFFARX1 I_30656 (I653884,I2683,I523758,I523886,);
not I_30657 (I523894,I523886);
nor I_30658 (I523911,I523894,I523792);
and I_30659 (I523928,I523911,I653887);
nor I_30660 (I523945,I523894,I523860);
nor I_30661 (I523741,I523852,I523945);
DFFARX1 I_30662 (I653878,I2683,I523758,I523985,);
nor I_30663 (I523993,I523985,I523852);
not I_30664 (I524010,I523993);
not I_30665 (I524027,I523985);
nor I_30666 (I524044,I524027,I523928);
DFFARX1 I_30667 (I524044,I2683,I523758,I523744,);
nand I_30668 (I524075,I653878,I653881);
and I_30669 (I524092,I524075,I653884);
DFFARX1 I_30670 (I524092,I2683,I523758,I524118,);
nor I_30671 (I524126,I524118,I523985);
DFFARX1 I_30672 (I524126,I2683,I523758,I523726,);
nand I_30673 (I524157,I524118,I524027);
nand I_30674 (I523735,I524010,I524157);
not I_30675 (I524188,I524118);
nor I_30676 (I524205,I524188,I523928);
DFFARX1 I_30677 (I524205,I2683,I523758,I523747,);
nor I_30678 (I524236,I653890,I653881);
or I_30679 (I523738,I523985,I524236);
nor I_30680 (I523729,I524118,I524236);
or I_30681 (I523732,I523852,I524236);
DFFARX1 I_30682 (I524236,I2683,I523758,I523750,);
not I_30683 (I524336,I2690);
DFFARX1 I_30684 (I909134,I2683,I524336,I524362,);
not I_30685 (I524370,I524362);
nand I_30686 (I524387,I909116,I909128);
and I_30687 (I524404,I524387,I909131);
DFFARX1 I_30688 (I524404,I2683,I524336,I524430,);
not I_30689 (I524438,I909125);
DFFARX1 I_30690 (I909122,I2683,I524336,I524464,);
not I_30691 (I524472,I524464);
nor I_30692 (I524489,I524472,I524370);
and I_30693 (I524506,I524489,I909125);
nor I_30694 (I524523,I524472,I524438);
nor I_30695 (I524319,I524430,I524523);
DFFARX1 I_30696 (I909140,I2683,I524336,I524563,);
nor I_30697 (I524571,I524563,I524430);
not I_30698 (I524588,I524571);
not I_30699 (I524605,I524563);
nor I_30700 (I524622,I524605,I524506);
DFFARX1 I_30701 (I524622,I2683,I524336,I524322,);
nand I_30702 (I524653,I909119,I909119);
and I_30703 (I524670,I524653,I909116);
DFFARX1 I_30704 (I524670,I2683,I524336,I524696,);
nor I_30705 (I524704,I524696,I524563);
DFFARX1 I_30706 (I524704,I2683,I524336,I524304,);
nand I_30707 (I524735,I524696,I524605);
nand I_30708 (I524313,I524588,I524735);
not I_30709 (I524766,I524696);
nor I_30710 (I524783,I524766,I524506);
DFFARX1 I_30711 (I524783,I2683,I524336,I524325,);
nor I_30712 (I524814,I909137,I909119);
or I_30713 (I524316,I524563,I524814);
nor I_30714 (I524307,I524696,I524814);
or I_30715 (I524310,I524430,I524814);
DFFARX1 I_30716 (I524814,I2683,I524336,I524328,);
not I_30717 (I524914,I2690);
DFFARX1 I_30718 (I992620,I2683,I524914,I524940,);
not I_30719 (I524948,I524940);
nand I_30720 (I524965,I992644,I992626);
and I_30721 (I524982,I524965,I992632);
DFFARX1 I_30722 (I524982,I2683,I524914,I525008,);
not I_30723 (I525016,I992638);
DFFARX1 I_30724 (I992623,I2683,I524914,I525042,);
not I_30725 (I525050,I525042);
nor I_30726 (I525067,I525050,I524948);
and I_30727 (I525084,I525067,I992638);
nor I_30728 (I525101,I525050,I525016);
nor I_30729 (I524897,I525008,I525101);
DFFARX1 I_30730 (I992635,I2683,I524914,I525141,);
nor I_30731 (I525149,I525141,I525008);
not I_30732 (I525166,I525149);
not I_30733 (I525183,I525141);
nor I_30734 (I525200,I525183,I525084);
DFFARX1 I_30735 (I525200,I2683,I524914,I524900,);
nand I_30736 (I525231,I992641,I992629);
and I_30737 (I525248,I525231,I992623);
DFFARX1 I_30738 (I525248,I2683,I524914,I525274,);
nor I_30739 (I525282,I525274,I525141);
DFFARX1 I_30740 (I525282,I2683,I524914,I524882,);
nand I_30741 (I525313,I525274,I525183);
nand I_30742 (I524891,I525166,I525313);
not I_30743 (I525344,I525274);
nor I_30744 (I525361,I525344,I525084);
DFFARX1 I_30745 (I525361,I2683,I524914,I524903,);
nor I_30746 (I525392,I992620,I992629);
or I_30747 (I524894,I525141,I525392);
nor I_30748 (I524885,I525274,I525392);
or I_30749 (I524888,I525008,I525392);
DFFARX1 I_30750 (I525392,I2683,I524914,I524906,);
not I_30751 (I525492,I2690);
DFFARX1 I_30752 (I27967,I2683,I525492,I525518,);
not I_30753 (I525526,I525518);
nand I_30754 (I525543,I27964,I27955);
and I_30755 (I525560,I525543,I27955);
DFFARX1 I_30756 (I525560,I2683,I525492,I525586,);
not I_30757 (I525594,I27958);
DFFARX1 I_30758 (I27973,I2683,I525492,I525620,);
not I_30759 (I525628,I525620);
nor I_30760 (I525645,I525628,I525526);
and I_30761 (I525662,I525645,I27958);
nor I_30762 (I525679,I525628,I525594);
nor I_30763 (I525475,I525586,I525679);
DFFARX1 I_30764 (I27958,I2683,I525492,I525719,);
nor I_30765 (I525727,I525719,I525586);
not I_30766 (I525744,I525727);
not I_30767 (I525761,I525719);
nor I_30768 (I525778,I525761,I525662);
DFFARX1 I_30769 (I525778,I2683,I525492,I525478,);
nand I_30770 (I525809,I27976,I27961);
and I_30771 (I525826,I525809,I27979);
DFFARX1 I_30772 (I525826,I2683,I525492,I525852,);
nor I_30773 (I525860,I525852,I525719);
DFFARX1 I_30774 (I525860,I2683,I525492,I525460,);
nand I_30775 (I525891,I525852,I525761);
nand I_30776 (I525469,I525744,I525891);
not I_30777 (I525922,I525852);
nor I_30778 (I525939,I525922,I525662);
DFFARX1 I_30779 (I525939,I2683,I525492,I525481,);
nor I_30780 (I525970,I27970,I27961);
or I_30781 (I525472,I525719,I525970);
nor I_30782 (I525463,I525852,I525970);
or I_30783 (I525466,I525586,I525970);
DFFARX1 I_30784 (I525970,I2683,I525492,I525484,);
not I_30785 (I526070,I2690);
DFFARX1 I_30786 (I228001,I2683,I526070,I526096,);
not I_30787 (I526104,I526096);
nand I_30788 (I526121,I228004,I227980);
and I_30789 (I526138,I526121,I227977);
DFFARX1 I_30790 (I526138,I2683,I526070,I526164,);
not I_30791 (I526172,I227983);
DFFARX1 I_30792 (I227977,I2683,I526070,I526198,);
not I_30793 (I526206,I526198);
nor I_30794 (I526223,I526206,I526104);
and I_30795 (I526240,I526223,I227983);
nor I_30796 (I526257,I526206,I526172);
nor I_30797 (I526053,I526164,I526257);
DFFARX1 I_30798 (I227986,I2683,I526070,I526297,);
nor I_30799 (I526305,I526297,I526164);
not I_30800 (I526322,I526305);
not I_30801 (I526339,I526297);
nor I_30802 (I526356,I526339,I526240);
DFFARX1 I_30803 (I526356,I2683,I526070,I526056,);
nand I_30804 (I526387,I227989,I227998);
and I_30805 (I526404,I526387,I227995);
DFFARX1 I_30806 (I526404,I2683,I526070,I526430,);
nor I_30807 (I526438,I526430,I526297);
DFFARX1 I_30808 (I526438,I2683,I526070,I526038,);
nand I_30809 (I526469,I526430,I526339);
nand I_30810 (I526047,I526322,I526469);
not I_30811 (I526500,I526430);
nor I_30812 (I526517,I526500,I526240);
DFFARX1 I_30813 (I526517,I2683,I526070,I526059,);
nor I_30814 (I526548,I227992,I227998);
or I_30815 (I526050,I526297,I526548);
nor I_30816 (I526041,I526430,I526548);
or I_30817 (I526044,I526164,I526548);
DFFARX1 I_30818 (I526548,I2683,I526070,I526062,);
not I_30819 (I526648,I2690);
DFFARX1 I_30820 (I206880,I2683,I526648,I526674,);
not I_30821 (I526682,I526674);
nand I_30822 (I526699,I206883,I206904);
and I_30823 (I526716,I526699,I206892);
DFFARX1 I_30824 (I526716,I2683,I526648,I526742,);
not I_30825 (I526750,I206889);
DFFARX1 I_30826 (I206880,I2683,I526648,I526776,);
not I_30827 (I526784,I526776);
nor I_30828 (I526801,I526784,I526682);
and I_30829 (I526818,I526801,I206889);
nor I_30830 (I526835,I526784,I526750);
nor I_30831 (I526631,I526742,I526835);
DFFARX1 I_30832 (I206898,I2683,I526648,I526875,);
nor I_30833 (I526883,I526875,I526742);
not I_30834 (I526900,I526883);
not I_30835 (I526917,I526875);
nor I_30836 (I526934,I526917,I526818);
DFFARX1 I_30837 (I526934,I2683,I526648,I526634,);
nand I_30838 (I526965,I206883,I206886);
and I_30839 (I526982,I526965,I206895);
DFFARX1 I_30840 (I526982,I2683,I526648,I527008,);
nor I_30841 (I527016,I527008,I526875);
DFFARX1 I_30842 (I527016,I2683,I526648,I526616,);
nand I_30843 (I527047,I527008,I526917);
nand I_30844 (I526625,I526900,I527047);
not I_30845 (I527078,I527008);
nor I_30846 (I527095,I527078,I526818);
DFFARX1 I_30847 (I527095,I2683,I526648,I526637,);
nor I_30848 (I527126,I206901,I206886);
or I_30849 (I526628,I526875,I527126);
nor I_30850 (I526619,I527008,I527126);
or I_30851 (I526622,I526742,I527126);
DFFARX1 I_30852 (I527126,I2683,I526648,I526640,);
not I_30853 (I527226,I2690);
DFFARX1 I_30854 (I21643,I2683,I527226,I527252,);
not I_30855 (I527260,I527252);
nand I_30856 (I527277,I21640,I21631);
and I_30857 (I527294,I527277,I21631);
DFFARX1 I_30858 (I527294,I2683,I527226,I527320,);
not I_30859 (I527328,I21634);
DFFARX1 I_30860 (I21649,I2683,I527226,I527354,);
not I_30861 (I527362,I527354);
nor I_30862 (I527379,I527362,I527260);
and I_30863 (I527396,I527379,I21634);
nor I_30864 (I527413,I527362,I527328);
nor I_30865 (I527209,I527320,I527413);
DFFARX1 I_30866 (I21634,I2683,I527226,I527453,);
nor I_30867 (I527461,I527453,I527320);
not I_30868 (I527478,I527461);
not I_30869 (I527495,I527453);
nor I_30870 (I527512,I527495,I527396);
DFFARX1 I_30871 (I527512,I2683,I527226,I527212,);
nand I_30872 (I527543,I21652,I21637);
and I_30873 (I527560,I527543,I21655);
DFFARX1 I_30874 (I527560,I2683,I527226,I527586,);
nor I_30875 (I527594,I527586,I527453);
DFFARX1 I_30876 (I527594,I2683,I527226,I527194,);
nand I_30877 (I527625,I527586,I527495);
nand I_30878 (I527203,I527478,I527625);
not I_30879 (I527656,I527586);
nor I_30880 (I527673,I527656,I527396);
DFFARX1 I_30881 (I527673,I2683,I527226,I527215,);
nor I_30882 (I527704,I21646,I21637);
or I_30883 (I527206,I527453,I527704);
nor I_30884 (I527197,I527586,I527704);
or I_30885 (I527200,I527320,I527704);
DFFARX1 I_30886 (I527704,I2683,I527226,I527218,);
not I_30887 (I527804,I2690);
DFFARX1 I_30888 (I698697,I2683,I527804,I527830,);
not I_30889 (I527838,I527830);
nand I_30890 (I527855,I698673,I698688);
and I_30891 (I527872,I527855,I698700);
DFFARX1 I_30892 (I527872,I2683,I527804,I527898,);
not I_30893 (I527906,I698685);
DFFARX1 I_30894 (I698676,I2683,I527804,I527932,);
not I_30895 (I527940,I527932);
nor I_30896 (I527957,I527940,I527838);
and I_30897 (I527974,I527957,I698685);
nor I_30898 (I527991,I527940,I527906);
nor I_30899 (I527787,I527898,I527991);
DFFARX1 I_30900 (I698673,I2683,I527804,I528031,);
nor I_30901 (I528039,I528031,I527898);
not I_30902 (I528056,I528039);
not I_30903 (I528073,I528031);
nor I_30904 (I528090,I528073,I527974);
DFFARX1 I_30905 (I528090,I2683,I527804,I527790,);
nand I_30906 (I528121,I698691,I698682);
and I_30907 (I528138,I528121,I698694);
DFFARX1 I_30908 (I528138,I2683,I527804,I528164,);
nor I_30909 (I528172,I528164,I528031);
DFFARX1 I_30910 (I528172,I2683,I527804,I527772,);
nand I_30911 (I528203,I528164,I528073);
nand I_30912 (I527781,I528056,I528203);
not I_30913 (I528234,I528164);
nor I_30914 (I528251,I528234,I527974);
DFFARX1 I_30915 (I528251,I2683,I527804,I527793,);
nor I_30916 (I528282,I698679,I698682);
or I_30917 (I527784,I528031,I528282);
nor I_30918 (I527775,I528164,I528282);
or I_30919 (I527778,I527898,I528282);
DFFARX1 I_30920 (I528282,I2683,I527804,I527796,);
not I_30921 (I528382,I2690);
DFFARX1 I_30922 (I929942,I2683,I528382,I528408,);
not I_30923 (I528416,I528408);
nand I_30924 (I528433,I929924,I929936);
and I_30925 (I528450,I528433,I929939);
DFFARX1 I_30926 (I528450,I2683,I528382,I528476,);
not I_30927 (I528484,I929933);
DFFARX1 I_30928 (I929930,I2683,I528382,I528510,);
not I_30929 (I528518,I528510);
nor I_30930 (I528535,I528518,I528416);
and I_30931 (I528552,I528535,I929933);
nor I_30932 (I528569,I528518,I528484);
nor I_30933 (I528365,I528476,I528569);
DFFARX1 I_30934 (I929948,I2683,I528382,I528609,);
nor I_30935 (I528617,I528609,I528476);
not I_30936 (I528634,I528617);
not I_30937 (I528651,I528609);
nor I_30938 (I528668,I528651,I528552);
DFFARX1 I_30939 (I528668,I2683,I528382,I528368,);
nand I_30940 (I528699,I929927,I929927);
and I_30941 (I528716,I528699,I929924);
DFFARX1 I_30942 (I528716,I2683,I528382,I528742,);
nor I_30943 (I528750,I528742,I528609);
DFFARX1 I_30944 (I528750,I2683,I528382,I528350,);
nand I_30945 (I528781,I528742,I528651);
nand I_30946 (I528359,I528634,I528781);
not I_30947 (I528812,I528742);
nor I_30948 (I528829,I528812,I528552);
DFFARX1 I_30949 (I528829,I2683,I528382,I528371,);
nor I_30950 (I528860,I929945,I929927);
or I_30951 (I528362,I528609,I528860);
nor I_30952 (I528353,I528742,I528860);
or I_30953 (I528356,I528476,I528860);
DFFARX1 I_30954 (I528860,I2683,I528382,I528374,);
not I_30955 (I528960,I2690);
DFFARX1 I_30956 (I749085,I2683,I528960,I528986,);
not I_30957 (I528994,I528986);
nand I_30958 (I529011,I749061,I749076);
and I_30959 (I529028,I529011,I749088);
DFFARX1 I_30960 (I529028,I2683,I528960,I529054,);
not I_30961 (I529062,I749073);
DFFARX1 I_30962 (I749064,I2683,I528960,I529088,);
not I_30963 (I529096,I529088);
nor I_30964 (I529113,I529096,I528994);
and I_30965 (I529130,I529113,I749073);
nor I_30966 (I529147,I529096,I529062);
nor I_30967 (I528943,I529054,I529147);
DFFARX1 I_30968 (I749061,I2683,I528960,I529187,);
nor I_30969 (I529195,I529187,I529054);
not I_30970 (I529212,I529195);
not I_30971 (I529229,I529187);
nor I_30972 (I529246,I529229,I529130);
DFFARX1 I_30973 (I529246,I2683,I528960,I528946,);
nand I_30974 (I529277,I749079,I749070);
and I_30975 (I529294,I529277,I749082);
DFFARX1 I_30976 (I529294,I2683,I528960,I529320,);
nor I_30977 (I529328,I529320,I529187);
DFFARX1 I_30978 (I529328,I2683,I528960,I528928,);
nand I_30979 (I529359,I529320,I529229);
nand I_30980 (I528937,I529212,I529359);
not I_30981 (I529390,I529320);
nor I_30982 (I529407,I529390,I529130);
DFFARX1 I_30983 (I529407,I2683,I528960,I528949,);
nor I_30984 (I529438,I749067,I749070);
or I_30985 (I528940,I529187,I529438);
nor I_30986 (I528931,I529320,I529438);
or I_30987 (I528934,I529054,I529438);
DFFARX1 I_30988 (I529438,I2683,I528960,I528952,);
not I_30989 (I529538,I2690);
DFFARX1 I_30990 (I134290,I2683,I529538,I529564,);
not I_30991 (I529572,I529564);
nand I_30992 (I529589,I134293,I134314);
and I_30993 (I529606,I529589,I134302);
DFFARX1 I_30994 (I529606,I2683,I529538,I529632,);
not I_30995 (I529640,I134299);
DFFARX1 I_30996 (I134290,I2683,I529538,I529666,);
not I_30997 (I529674,I529666);
nor I_30998 (I529691,I529674,I529572);
and I_30999 (I529708,I529691,I134299);
nor I_31000 (I529725,I529674,I529640);
nor I_31001 (I529521,I529632,I529725);
DFFARX1 I_31002 (I134308,I2683,I529538,I529765,);
nor I_31003 (I529773,I529765,I529632);
not I_31004 (I529790,I529773);
not I_31005 (I529807,I529765);
nor I_31006 (I529824,I529807,I529708);
DFFARX1 I_31007 (I529824,I2683,I529538,I529524,);
nand I_31008 (I529855,I134293,I134296);
and I_31009 (I529872,I529855,I134305);
DFFARX1 I_31010 (I529872,I2683,I529538,I529898,);
nor I_31011 (I529906,I529898,I529765);
DFFARX1 I_31012 (I529906,I2683,I529538,I529506,);
nand I_31013 (I529937,I529898,I529807);
nand I_31014 (I529515,I529790,I529937);
not I_31015 (I529968,I529898);
nor I_31016 (I529985,I529968,I529708);
DFFARX1 I_31017 (I529985,I2683,I529538,I529527,);
nor I_31018 (I530016,I134311,I134296);
or I_31019 (I529518,I529765,I530016);
nor I_31020 (I529509,I529898,I530016);
or I_31021 (I529512,I529632,I530016);
DFFARX1 I_31022 (I530016,I2683,I529538,I529530,);
not I_31023 (I530116,I2690);
DFFARX1 I_31024 (I920116,I2683,I530116,I530142,);
not I_31025 (I530150,I530142);
nand I_31026 (I530167,I920098,I920110);
and I_31027 (I530184,I530167,I920113);
DFFARX1 I_31028 (I530184,I2683,I530116,I530210,);
not I_31029 (I530218,I920107);
DFFARX1 I_31030 (I920104,I2683,I530116,I530244,);
not I_31031 (I530252,I530244);
nor I_31032 (I530269,I530252,I530150);
and I_31033 (I530286,I530269,I920107);
nor I_31034 (I530303,I530252,I530218);
nor I_31035 (I530099,I530210,I530303);
DFFARX1 I_31036 (I920122,I2683,I530116,I530343,);
nor I_31037 (I530351,I530343,I530210);
not I_31038 (I530368,I530351);
not I_31039 (I530385,I530343);
nor I_31040 (I530402,I530385,I530286);
DFFARX1 I_31041 (I530402,I2683,I530116,I530102,);
nand I_31042 (I530433,I920101,I920101);
and I_31043 (I530450,I530433,I920098);
DFFARX1 I_31044 (I530450,I2683,I530116,I530476,);
nor I_31045 (I530484,I530476,I530343);
DFFARX1 I_31046 (I530484,I2683,I530116,I530084,);
nand I_31047 (I530515,I530476,I530385);
nand I_31048 (I530093,I530368,I530515);
not I_31049 (I530546,I530476);
nor I_31050 (I530563,I530546,I530286);
DFFARX1 I_31051 (I530563,I2683,I530116,I530105,);
nor I_31052 (I530594,I920119,I920101);
or I_31053 (I530096,I530343,I530594);
nor I_31054 (I530087,I530476,I530594);
or I_31055 (I530090,I530210,I530594);
DFFARX1 I_31056 (I530594,I2683,I530116,I530108,);
not I_31057 (I530694,I2690);
DFFARX1 I_31058 (I437604,I2683,I530694,I530720,);
not I_31059 (I530728,I530720);
nand I_31060 (I530745,I437613,I437622);
and I_31061 (I530762,I530745,I437628);
DFFARX1 I_31062 (I530762,I2683,I530694,I530788,);
not I_31063 (I530796,I437625);
DFFARX1 I_31064 (I437610,I2683,I530694,I530822,);
not I_31065 (I530830,I530822);
nor I_31066 (I530847,I530830,I530728);
and I_31067 (I530864,I530847,I437625);
nor I_31068 (I530881,I530830,I530796);
nor I_31069 (I530677,I530788,I530881);
DFFARX1 I_31070 (I437619,I2683,I530694,I530921,);
nor I_31071 (I530929,I530921,I530788);
not I_31072 (I530946,I530929);
not I_31073 (I530963,I530921);
nor I_31074 (I530980,I530963,I530864);
DFFARX1 I_31075 (I530980,I2683,I530694,I530680,);
nand I_31076 (I531011,I437616,I437607);
and I_31077 (I531028,I531011,I437604);
DFFARX1 I_31078 (I531028,I2683,I530694,I531054,);
nor I_31079 (I531062,I531054,I530921);
DFFARX1 I_31080 (I531062,I2683,I530694,I530662,);
nand I_31081 (I531093,I531054,I530963);
nand I_31082 (I530671,I530946,I531093);
not I_31083 (I531124,I531054);
nor I_31084 (I531141,I531124,I530864);
DFFARX1 I_31085 (I531141,I2683,I530694,I530683,);
nor I_31086 (I531172,I437607,I437607);
or I_31087 (I530674,I530921,I531172);
nor I_31088 (I530665,I531054,I531172);
or I_31089 (I530668,I530788,I531172);
DFFARX1 I_31090 (I531172,I2683,I530694,I530686,);
not I_31091 (I531272,I2690);
DFFARX1 I_31092 (I475174,I2683,I531272,I531298,);
not I_31093 (I531306,I531298);
nand I_31094 (I531323,I475183,I475192);
and I_31095 (I531340,I531323,I475198);
DFFARX1 I_31096 (I531340,I2683,I531272,I531366,);
not I_31097 (I531374,I475195);
DFFARX1 I_31098 (I475180,I2683,I531272,I531400,);
not I_31099 (I531408,I531400);
nor I_31100 (I531425,I531408,I531306);
and I_31101 (I531442,I531425,I475195);
nor I_31102 (I531459,I531408,I531374);
nor I_31103 (I531255,I531366,I531459);
DFFARX1 I_31104 (I475189,I2683,I531272,I531499,);
nor I_31105 (I531507,I531499,I531366);
not I_31106 (I531524,I531507);
not I_31107 (I531541,I531499);
nor I_31108 (I531558,I531541,I531442);
DFFARX1 I_31109 (I531558,I2683,I531272,I531258,);
nand I_31110 (I531589,I475186,I475177);
and I_31111 (I531606,I531589,I475174);
DFFARX1 I_31112 (I531606,I2683,I531272,I531632,);
nor I_31113 (I531640,I531632,I531499);
DFFARX1 I_31114 (I531640,I2683,I531272,I531240,);
nand I_31115 (I531671,I531632,I531541);
nand I_31116 (I531249,I531524,I531671);
not I_31117 (I531702,I531632);
nor I_31118 (I531719,I531702,I531442);
DFFARX1 I_31119 (I531719,I2683,I531272,I531261,);
nor I_31120 (I531750,I475177,I475177);
or I_31121 (I531252,I531499,I531750);
nor I_31122 (I531243,I531632,I531750);
or I_31123 (I531246,I531366,I531750);
DFFARX1 I_31124 (I531750,I2683,I531272,I531264,);
not I_31125 (I531850,I2690);
DFFARX1 I_31126 (I780739,I2683,I531850,I531876,);
not I_31127 (I531884,I531876);
nand I_31128 (I531901,I780715,I780730);
and I_31129 (I531918,I531901,I780742);
DFFARX1 I_31130 (I531918,I2683,I531850,I531944,);
not I_31131 (I531952,I780727);
DFFARX1 I_31132 (I780718,I2683,I531850,I531978,);
not I_31133 (I531986,I531978);
nor I_31134 (I532003,I531986,I531884);
and I_31135 (I532020,I532003,I780727);
nor I_31136 (I532037,I531986,I531952);
nor I_31137 (I531833,I531944,I532037);
DFFARX1 I_31138 (I780715,I2683,I531850,I532077,);
nor I_31139 (I532085,I532077,I531944);
not I_31140 (I532102,I532085);
not I_31141 (I532119,I532077);
nor I_31142 (I532136,I532119,I532020);
DFFARX1 I_31143 (I532136,I2683,I531850,I531836,);
nand I_31144 (I532167,I780733,I780724);
and I_31145 (I532184,I532167,I780736);
DFFARX1 I_31146 (I532184,I2683,I531850,I532210,);
nor I_31147 (I532218,I532210,I532077);
DFFARX1 I_31148 (I532218,I2683,I531850,I531818,);
nand I_31149 (I532249,I532210,I532119);
nand I_31150 (I531827,I532102,I532249);
not I_31151 (I532280,I532210);
nor I_31152 (I532297,I532280,I532020);
DFFARX1 I_31153 (I532297,I2683,I531850,I531839,);
nor I_31154 (I532328,I780721,I780724);
or I_31155 (I531830,I532077,I532328);
nor I_31156 (I531821,I532210,I532328);
or I_31157 (I531824,I531944,I532328);
DFFARX1 I_31158 (I532328,I2683,I531850,I531842,);
not I_31159 (I532428,I2690);
DFFARX1 I_31160 (I780093,I2683,I532428,I532454,);
not I_31161 (I532462,I532454);
nand I_31162 (I532479,I780069,I780084);
and I_31163 (I532496,I532479,I780096);
DFFARX1 I_31164 (I532496,I2683,I532428,I532522,);
not I_31165 (I532530,I780081);
DFFARX1 I_31166 (I780072,I2683,I532428,I532556,);
not I_31167 (I532564,I532556);
nor I_31168 (I532581,I532564,I532462);
and I_31169 (I532598,I532581,I780081);
nor I_31170 (I532615,I532564,I532530);
nor I_31171 (I532411,I532522,I532615);
DFFARX1 I_31172 (I780069,I2683,I532428,I532655,);
nor I_31173 (I532663,I532655,I532522);
not I_31174 (I532680,I532663);
not I_31175 (I532697,I532655);
nor I_31176 (I532714,I532697,I532598);
DFFARX1 I_31177 (I532714,I2683,I532428,I532414,);
nand I_31178 (I532745,I780087,I780078);
and I_31179 (I532762,I532745,I780090);
DFFARX1 I_31180 (I532762,I2683,I532428,I532788,);
nor I_31181 (I532796,I532788,I532655);
DFFARX1 I_31182 (I532796,I2683,I532428,I532396,);
nand I_31183 (I532827,I532788,I532697);
nand I_31184 (I532405,I532680,I532827);
not I_31185 (I532858,I532788);
nor I_31186 (I532875,I532858,I532598);
DFFARX1 I_31187 (I532875,I2683,I532428,I532417,);
nor I_31188 (I532906,I780075,I780078);
or I_31189 (I532408,I532655,I532906);
nor I_31190 (I532399,I532788,I532906);
or I_31191 (I532402,I532522,I532906);
DFFARX1 I_31192 (I532906,I2683,I532428,I532420,);
not I_31193 (I533006,I2690);
DFFARX1 I_31194 (I836884,I2683,I533006,I533032,);
not I_31195 (I533040,I533032);
nand I_31196 (I533057,I836866,I836878);
and I_31197 (I533074,I533057,I836881);
DFFARX1 I_31198 (I533074,I2683,I533006,I533100,);
not I_31199 (I533108,I836875);
DFFARX1 I_31200 (I836872,I2683,I533006,I533134,);
not I_31201 (I533142,I533134);
nor I_31202 (I533159,I533142,I533040);
and I_31203 (I533176,I533159,I836875);
nor I_31204 (I533193,I533142,I533108);
nor I_31205 (I532989,I533100,I533193);
DFFARX1 I_31206 (I836890,I2683,I533006,I533233,);
nor I_31207 (I533241,I533233,I533100);
not I_31208 (I533258,I533241);
not I_31209 (I533275,I533233);
nor I_31210 (I533292,I533275,I533176);
DFFARX1 I_31211 (I533292,I2683,I533006,I532992,);
nand I_31212 (I533323,I836869,I836869);
and I_31213 (I533340,I533323,I836866);
DFFARX1 I_31214 (I533340,I2683,I533006,I533366,);
nor I_31215 (I533374,I533366,I533233);
DFFARX1 I_31216 (I533374,I2683,I533006,I532974,);
nand I_31217 (I533405,I533366,I533275);
nand I_31218 (I532983,I533258,I533405);
not I_31219 (I533436,I533366);
nor I_31220 (I533453,I533436,I533176);
DFFARX1 I_31221 (I533453,I2683,I533006,I532995,);
nor I_31222 (I533484,I836887,I836869);
or I_31223 (I532986,I533233,I533484);
nor I_31224 (I532977,I533366,I533484);
or I_31225 (I532980,I533100,I533484);
DFFARX1 I_31226 (I533484,I2683,I533006,I532998,);
not I_31227 (I533584,I2690);
DFFARX1 I_31228 (I875032,I2683,I533584,I533610,);
not I_31229 (I533618,I533610);
nand I_31230 (I533635,I875014,I875026);
and I_31231 (I533652,I533635,I875029);
DFFARX1 I_31232 (I533652,I2683,I533584,I533678,);
not I_31233 (I533686,I875023);
DFFARX1 I_31234 (I875020,I2683,I533584,I533712,);
not I_31235 (I533720,I533712);
nor I_31236 (I533737,I533720,I533618);
and I_31237 (I533754,I533737,I875023);
nor I_31238 (I533771,I533720,I533686);
nor I_31239 (I533567,I533678,I533771);
DFFARX1 I_31240 (I875038,I2683,I533584,I533811,);
nor I_31241 (I533819,I533811,I533678);
not I_31242 (I533836,I533819);
not I_31243 (I533853,I533811);
nor I_31244 (I533870,I533853,I533754);
DFFARX1 I_31245 (I533870,I2683,I533584,I533570,);
nand I_31246 (I533901,I875017,I875017);
and I_31247 (I533918,I533901,I875014);
DFFARX1 I_31248 (I533918,I2683,I533584,I533944,);
nor I_31249 (I533952,I533944,I533811);
DFFARX1 I_31250 (I533952,I2683,I533584,I533552,);
nand I_31251 (I533983,I533944,I533853);
nand I_31252 (I533561,I533836,I533983);
not I_31253 (I534014,I533944);
nor I_31254 (I534031,I534014,I533754);
DFFARX1 I_31255 (I534031,I2683,I533584,I533573,);
nor I_31256 (I534062,I875035,I875017);
or I_31257 (I533564,I533811,I534062);
nor I_31258 (I533555,I533944,I534062);
or I_31259 (I533558,I533678,I534062);
DFFARX1 I_31260 (I534062,I2683,I533584,I533576,);
not I_31261 (I534162,I2690);
DFFARX1 I_31262 (I98576,I2683,I534162,I534188,);
not I_31263 (I534196,I534188);
nand I_31264 (I534213,I98585,I98594);
and I_31265 (I534230,I534213,I98573);
DFFARX1 I_31266 (I534230,I2683,I534162,I534256,);
not I_31267 (I534264,I98576);
DFFARX1 I_31268 (I98591,I2683,I534162,I534290,);
not I_31269 (I534298,I534290);
nor I_31270 (I534315,I534298,I534196);
and I_31271 (I534332,I534315,I98576);
nor I_31272 (I534349,I534298,I534264);
nor I_31273 (I534145,I534256,I534349);
DFFARX1 I_31274 (I98582,I2683,I534162,I534389,);
nor I_31275 (I534397,I534389,I534256);
not I_31276 (I534414,I534397);
not I_31277 (I534431,I534389);
nor I_31278 (I534448,I534431,I534332);
DFFARX1 I_31279 (I534448,I2683,I534162,I534148,);
nand I_31280 (I534479,I98597,I98573);
and I_31281 (I534496,I534479,I98579);
DFFARX1 I_31282 (I534496,I2683,I534162,I534522,);
nor I_31283 (I534530,I534522,I534389);
DFFARX1 I_31284 (I534530,I2683,I534162,I534130,);
nand I_31285 (I534561,I534522,I534431);
nand I_31286 (I534139,I534414,I534561);
not I_31287 (I534592,I534522);
nor I_31288 (I534609,I534592,I534332);
DFFARX1 I_31289 (I534609,I2683,I534162,I534151,);
nor I_31290 (I534640,I98588,I98573);
or I_31291 (I534142,I534389,I534640);
nor I_31292 (I534133,I534522,I534640);
or I_31293 (I534136,I534256,I534640);
DFFARX1 I_31294 (I534640,I2683,I534162,I534154,);
not I_31295 (I534740,I2690);
DFFARX1 I_31296 (I686567,I2683,I534740,I534766,);
not I_31297 (I534774,I534766);
nand I_31298 (I534791,I686555,I686573);
and I_31299 (I534808,I534791,I686570);
DFFARX1 I_31300 (I534808,I2683,I534740,I534834,);
not I_31301 (I534842,I686561);
DFFARX1 I_31302 (I686558,I2683,I534740,I534868,);
not I_31303 (I534876,I534868);
nor I_31304 (I534893,I534876,I534774);
and I_31305 (I534910,I534893,I686561);
nor I_31306 (I534927,I534876,I534842);
nor I_31307 (I534723,I534834,I534927);
DFFARX1 I_31308 (I686552,I2683,I534740,I534967,);
nor I_31309 (I534975,I534967,I534834);
not I_31310 (I534992,I534975);
not I_31311 (I535009,I534967);
nor I_31312 (I535026,I535009,I534910);
DFFARX1 I_31313 (I535026,I2683,I534740,I534726,);
nand I_31314 (I535057,I686552,I686555);
and I_31315 (I535074,I535057,I686558);
DFFARX1 I_31316 (I535074,I2683,I534740,I535100,);
nor I_31317 (I535108,I535100,I534967);
DFFARX1 I_31318 (I535108,I2683,I534740,I534708,);
nand I_31319 (I535139,I535100,I535009);
nand I_31320 (I534717,I534992,I535139);
not I_31321 (I535170,I535100);
nor I_31322 (I535187,I535170,I534910);
DFFARX1 I_31323 (I535187,I2683,I534740,I534729,);
nor I_31324 (I535218,I686564,I686555);
or I_31325 (I534720,I534967,I535218);
nor I_31326 (I534711,I535100,I535218);
or I_31327 (I534714,I534834,I535218);
DFFARX1 I_31328 (I535218,I2683,I534740,I534732,);
not I_31329 (I535318,I2690);
DFFARX1 I_31330 (I71172,I2683,I535318,I535344,);
not I_31331 (I535352,I535344);
nand I_31332 (I535369,I71181,I71190);
and I_31333 (I535386,I535369,I71169);
DFFARX1 I_31334 (I535386,I2683,I535318,I535412,);
not I_31335 (I535420,I71172);
DFFARX1 I_31336 (I71187,I2683,I535318,I535446,);
not I_31337 (I535454,I535446);
nor I_31338 (I535471,I535454,I535352);
and I_31339 (I535488,I535471,I71172);
nor I_31340 (I535505,I535454,I535420);
nor I_31341 (I535301,I535412,I535505);
DFFARX1 I_31342 (I71178,I2683,I535318,I535545,);
nor I_31343 (I535553,I535545,I535412);
not I_31344 (I535570,I535553);
not I_31345 (I535587,I535545);
nor I_31346 (I535604,I535587,I535488);
DFFARX1 I_31347 (I535604,I2683,I535318,I535304,);
nand I_31348 (I535635,I71193,I71169);
and I_31349 (I535652,I535635,I71175);
DFFARX1 I_31350 (I535652,I2683,I535318,I535678,);
nor I_31351 (I535686,I535678,I535545);
DFFARX1 I_31352 (I535686,I2683,I535318,I535286,);
nand I_31353 (I535717,I535678,I535587);
nand I_31354 (I535295,I535570,I535717);
not I_31355 (I535748,I535678);
nor I_31356 (I535765,I535748,I535488);
DFFARX1 I_31357 (I535765,I2683,I535318,I535307,);
nor I_31358 (I535796,I71184,I71169);
or I_31359 (I535298,I535545,I535796);
nor I_31360 (I535289,I535678,I535796);
or I_31361 (I535292,I535412,I535796);
DFFARX1 I_31362 (I535796,I2683,I535318,I535310,);
not I_31363 (I535896,I2690);
DFFARX1 I_31364 (I961374,I2683,I535896,I535922,);
not I_31365 (I535930,I535922);
nand I_31366 (I535947,I961377,I961386);
and I_31367 (I535964,I535947,I961389);
DFFARX1 I_31368 (I535964,I2683,I535896,I535990,);
not I_31369 (I535998,I961398);
DFFARX1 I_31370 (I961380,I2683,I535896,I536024,);
not I_31371 (I536032,I536024);
nor I_31372 (I536049,I536032,I535930);
and I_31373 (I536066,I536049,I961398);
nor I_31374 (I536083,I536032,I535998);
nor I_31375 (I535879,I535990,I536083);
DFFARX1 I_31376 (I961377,I2683,I535896,I536123,);
nor I_31377 (I536131,I536123,I535990);
not I_31378 (I536148,I536131);
not I_31379 (I536165,I536123);
nor I_31380 (I536182,I536165,I536066);
DFFARX1 I_31381 (I536182,I2683,I535896,I535882,);
nand I_31382 (I536213,I961395,I961374);
and I_31383 (I536230,I536213,I961392);
DFFARX1 I_31384 (I536230,I2683,I535896,I536256,);
nor I_31385 (I536264,I536256,I536123);
DFFARX1 I_31386 (I536264,I2683,I535896,I535864,);
nand I_31387 (I536295,I536256,I536165);
nand I_31388 (I535873,I536148,I536295);
not I_31389 (I536326,I536256);
nor I_31390 (I536343,I536326,I536066);
DFFARX1 I_31391 (I536343,I2683,I535896,I535885,);
nor I_31392 (I536374,I961383,I961374);
or I_31393 (I535876,I536123,I536374);
nor I_31394 (I535867,I536256,I536374);
or I_31395 (I535870,I535990,I536374);
DFFARX1 I_31396 (I536374,I2683,I535896,I535888,);
not I_31397 (I536474,I2690);
DFFARX1 I_31398 (I427642,I2683,I536474,I536500,);
not I_31399 (I536508,I536500);
nand I_31400 (I536525,I427657,I427642);
and I_31401 (I536542,I536525,I427645);
DFFARX1 I_31402 (I536542,I2683,I536474,I536568,);
not I_31403 (I536576,I427645);
DFFARX1 I_31404 (I427654,I2683,I536474,I536602,);
not I_31405 (I536610,I536602);
nor I_31406 (I536627,I536610,I536508);
and I_31407 (I536644,I536627,I427645);
nor I_31408 (I536661,I536610,I536576);
nor I_31409 (I536457,I536568,I536661);
DFFARX1 I_31410 (I427648,I2683,I536474,I536701,);
nor I_31411 (I536709,I536701,I536568);
not I_31412 (I536726,I536709);
not I_31413 (I536743,I536701);
nor I_31414 (I536760,I536743,I536644);
DFFARX1 I_31415 (I536760,I2683,I536474,I536460,);
nand I_31416 (I536791,I427651,I427660);
and I_31417 (I536808,I536791,I427666);
DFFARX1 I_31418 (I536808,I2683,I536474,I536834,);
nor I_31419 (I536842,I536834,I536701);
DFFARX1 I_31420 (I536842,I2683,I536474,I536442,);
nand I_31421 (I536873,I536834,I536743);
nand I_31422 (I536451,I536726,I536873);
not I_31423 (I536904,I536834);
nor I_31424 (I536921,I536904,I536644);
DFFARX1 I_31425 (I536921,I2683,I536474,I536463,);
nor I_31426 (I536952,I427663,I427660);
or I_31427 (I536454,I536701,I536952);
nor I_31428 (I536445,I536834,I536952);
or I_31429 (I536448,I536568,I536952);
DFFARX1 I_31430 (I536952,I2683,I536474,I536466,);
not I_31431 (I537052,I2690);
DFFARX1 I_31432 (I1035266,I2683,I537052,I537078,);
not I_31433 (I537086,I537078);
nand I_31434 (I537103,I1035251,I1035239);
and I_31435 (I537120,I537103,I1035254);
DFFARX1 I_31436 (I537120,I2683,I537052,I537146,);
not I_31437 (I537154,I1035239);
DFFARX1 I_31438 (I1035257,I2683,I537052,I537180,);
not I_31439 (I537188,I537180);
nor I_31440 (I537205,I537188,I537086);
and I_31441 (I537222,I537205,I1035239);
nor I_31442 (I537239,I537188,I537154);
nor I_31443 (I537035,I537146,I537239);
DFFARX1 I_31444 (I1035245,I2683,I537052,I537279,);
nor I_31445 (I537287,I537279,I537146);
not I_31446 (I537304,I537287);
not I_31447 (I537321,I537279);
nor I_31448 (I537338,I537321,I537222);
DFFARX1 I_31449 (I537338,I2683,I537052,I537038,);
nand I_31450 (I537369,I1035242,I1035248);
and I_31451 (I537386,I537369,I1035263);
DFFARX1 I_31452 (I537386,I2683,I537052,I537412,);
nor I_31453 (I537420,I537412,I537279);
DFFARX1 I_31454 (I537420,I2683,I537052,I537020,);
nand I_31455 (I537451,I537412,I537321);
nand I_31456 (I537029,I537304,I537451);
not I_31457 (I537482,I537412);
nor I_31458 (I537499,I537482,I537222);
DFFARX1 I_31459 (I537499,I2683,I537052,I537041,);
nor I_31460 (I537530,I1035260,I1035248);
or I_31461 (I537032,I537279,I537530);
nor I_31462 (I537023,I537412,I537530);
or I_31463 (I537026,I537146,I537530);
DFFARX1 I_31464 (I537530,I2683,I537052,I537044,);
not I_31465 (I537630,I2690);
DFFARX1 I_31466 (I183675,I2683,I537630,I537656,);
not I_31467 (I537664,I537656);
nand I_31468 (I537681,I183678,I183699);
and I_31469 (I537698,I537681,I183687);
DFFARX1 I_31470 (I537698,I2683,I537630,I537724,);
not I_31471 (I537732,I183684);
DFFARX1 I_31472 (I183675,I2683,I537630,I537758,);
not I_31473 (I537766,I537758);
nor I_31474 (I537783,I537766,I537664);
and I_31475 (I537800,I537783,I183684);
nor I_31476 (I537817,I537766,I537732);
nor I_31477 (I537613,I537724,I537817);
DFFARX1 I_31478 (I183693,I2683,I537630,I537857,);
nor I_31479 (I537865,I537857,I537724);
not I_31480 (I537882,I537865);
not I_31481 (I537899,I537857);
nor I_31482 (I537916,I537899,I537800);
DFFARX1 I_31483 (I537916,I2683,I537630,I537616,);
nand I_31484 (I537947,I183678,I183681);
and I_31485 (I537964,I537947,I183690);
DFFARX1 I_31486 (I537964,I2683,I537630,I537990,);
nor I_31487 (I537998,I537990,I537857);
DFFARX1 I_31488 (I537998,I2683,I537630,I537598,);
nand I_31489 (I538029,I537990,I537899);
nand I_31490 (I537607,I537882,I538029);
not I_31491 (I538060,I537990);
nor I_31492 (I538077,I538060,I537800);
DFFARX1 I_31493 (I538077,I2683,I537630,I537619,);
nor I_31494 (I538108,I183696,I183681);
or I_31495 (I537610,I537857,I538108);
nor I_31496 (I537601,I537990,I538108);
or I_31497 (I537604,I537724,I538108);
DFFARX1 I_31498 (I538108,I2683,I537630,I537622,);
not I_31499 (I538208,I2690);
DFFARX1 I_31500 (I238541,I2683,I538208,I538234,);
not I_31501 (I538242,I538234);
nand I_31502 (I538259,I238544,I238520);
and I_31503 (I538276,I538259,I238517);
DFFARX1 I_31504 (I538276,I2683,I538208,I538302,);
not I_31505 (I538310,I238523);
DFFARX1 I_31506 (I238517,I2683,I538208,I538336,);
not I_31507 (I538344,I538336);
nor I_31508 (I538361,I538344,I538242);
and I_31509 (I538378,I538361,I238523);
nor I_31510 (I538395,I538344,I538310);
nor I_31511 (I538191,I538302,I538395);
DFFARX1 I_31512 (I238526,I2683,I538208,I538435,);
nor I_31513 (I538443,I538435,I538302);
not I_31514 (I538460,I538443);
not I_31515 (I538477,I538435);
nor I_31516 (I538494,I538477,I538378);
DFFARX1 I_31517 (I538494,I2683,I538208,I538194,);
nand I_31518 (I538525,I238529,I238538);
and I_31519 (I538542,I538525,I238535);
DFFARX1 I_31520 (I538542,I2683,I538208,I538568,);
nor I_31521 (I538576,I538568,I538435);
DFFARX1 I_31522 (I538576,I2683,I538208,I538176,);
nand I_31523 (I538607,I538568,I538477);
nand I_31524 (I538185,I538460,I538607);
not I_31525 (I538638,I538568);
nor I_31526 (I538655,I538638,I538378);
DFFARX1 I_31527 (I538655,I2683,I538208,I538197,);
nor I_31528 (I538686,I238532,I238538);
or I_31529 (I538188,I538435,I538686);
nor I_31530 (I538179,I538568,I538686);
or I_31531 (I538182,I538302,I538686);
DFFARX1 I_31532 (I538686,I2683,I538208,I538200,);
not I_31533 (I538786,I2690);
DFFARX1 I_31534 (I226947,I2683,I538786,I538812,);
not I_31535 (I538820,I538812);
nand I_31536 (I538837,I226950,I226926);
and I_31537 (I538854,I538837,I226923);
DFFARX1 I_31538 (I538854,I2683,I538786,I538880,);
not I_31539 (I538888,I226929);
DFFARX1 I_31540 (I226923,I2683,I538786,I538914,);
not I_31541 (I538922,I538914);
nor I_31542 (I538939,I538922,I538820);
and I_31543 (I538956,I538939,I226929);
nor I_31544 (I538973,I538922,I538888);
nor I_31545 (I538769,I538880,I538973);
DFFARX1 I_31546 (I226932,I2683,I538786,I539013,);
nor I_31547 (I539021,I539013,I538880);
not I_31548 (I539038,I539021);
not I_31549 (I539055,I539013);
nor I_31550 (I539072,I539055,I538956);
DFFARX1 I_31551 (I539072,I2683,I538786,I538772,);
nand I_31552 (I539103,I226935,I226944);
and I_31553 (I539120,I539103,I226941);
DFFARX1 I_31554 (I539120,I2683,I538786,I539146,);
nor I_31555 (I539154,I539146,I539013);
DFFARX1 I_31556 (I539154,I2683,I538786,I538754,);
nand I_31557 (I539185,I539146,I539055);
nand I_31558 (I538763,I539038,I539185);
not I_31559 (I539216,I539146);
nor I_31560 (I539233,I539216,I538956);
DFFARX1 I_31561 (I539233,I2683,I538786,I538775,);
nor I_31562 (I539264,I226938,I226944);
or I_31563 (I538766,I539013,I539264);
nor I_31564 (I538757,I539146,I539264);
or I_31565 (I538760,I538880,I539264);
DFFARX1 I_31566 (I539264,I2683,I538786,I538778,);
not I_31567 (I539364,I2690);
DFFARX1 I_31568 (I273850,I2683,I539364,I539390,);
not I_31569 (I539398,I539390);
nand I_31570 (I539415,I273853,I273829);
and I_31571 (I539432,I539415,I273826);
DFFARX1 I_31572 (I539432,I2683,I539364,I539458,);
not I_31573 (I539466,I273832);
DFFARX1 I_31574 (I273826,I2683,I539364,I539492,);
not I_31575 (I539500,I539492);
nor I_31576 (I539517,I539500,I539398);
and I_31577 (I539534,I539517,I273832);
nor I_31578 (I539551,I539500,I539466);
nor I_31579 (I539347,I539458,I539551);
DFFARX1 I_31580 (I273835,I2683,I539364,I539591,);
nor I_31581 (I539599,I539591,I539458);
not I_31582 (I539616,I539599);
not I_31583 (I539633,I539591);
nor I_31584 (I539650,I539633,I539534);
DFFARX1 I_31585 (I539650,I2683,I539364,I539350,);
nand I_31586 (I539681,I273838,I273847);
and I_31587 (I539698,I539681,I273844);
DFFARX1 I_31588 (I539698,I2683,I539364,I539724,);
nor I_31589 (I539732,I539724,I539591);
DFFARX1 I_31590 (I539732,I2683,I539364,I539332,);
nand I_31591 (I539763,I539724,I539633);
nand I_31592 (I539341,I539616,I539763);
not I_31593 (I539794,I539724);
nor I_31594 (I539811,I539794,I539534);
DFFARX1 I_31595 (I539811,I2683,I539364,I539353,);
nor I_31596 (I539842,I273841,I273847);
or I_31597 (I539344,I539591,I539842);
nor I_31598 (I539335,I539724,I539842);
or I_31599 (I539338,I539458,I539842);
DFFARX1 I_31600 (I539842,I2683,I539364,I539356,);
not I_31601 (I539942,I2690);
DFFARX1 I_31602 (I282282,I2683,I539942,I539968,);
not I_31603 (I539976,I539968);
nand I_31604 (I539993,I282285,I282261);
and I_31605 (I540010,I539993,I282258);
DFFARX1 I_31606 (I540010,I2683,I539942,I540036,);
not I_31607 (I540044,I282264);
DFFARX1 I_31608 (I282258,I2683,I539942,I540070,);
not I_31609 (I540078,I540070);
nor I_31610 (I540095,I540078,I539976);
and I_31611 (I540112,I540095,I282264);
nor I_31612 (I540129,I540078,I540044);
nor I_31613 (I539925,I540036,I540129);
DFFARX1 I_31614 (I282267,I2683,I539942,I540169,);
nor I_31615 (I540177,I540169,I540036);
not I_31616 (I540194,I540177);
not I_31617 (I540211,I540169);
nor I_31618 (I540228,I540211,I540112);
DFFARX1 I_31619 (I540228,I2683,I539942,I539928,);
nand I_31620 (I540259,I282270,I282279);
and I_31621 (I540276,I540259,I282276);
DFFARX1 I_31622 (I540276,I2683,I539942,I540302,);
nor I_31623 (I540310,I540302,I540169);
DFFARX1 I_31624 (I540310,I2683,I539942,I539910,);
nand I_31625 (I540341,I540302,I540211);
nand I_31626 (I539919,I540194,I540341);
not I_31627 (I540372,I540302);
nor I_31628 (I540389,I540372,I540112);
DFFARX1 I_31629 (I540389,I2683,I539942,I539931,);
nor I_31630 (I540420,I282273,I282279);
or I_31631 (I539922,I540169,I540420);
nor I_31632 (I539913,I540302,I540420);
or I_31633 (I539916,I540036,I540420);
DFFARX1 I_31634 (I540420,I2683,I539942,I539934,);
not I_31635 (I540520,I2690);
DFFARX1 I_31636 (I668122,I2683,I540520,I540546,);
not I_31637 (I540554,I540546);
nand I_31638 (I540571,I668110,I668128);
and I_31639 (I540588,I540571,I668125);
DFFARX1 I_31640 (I540588,I2683,I540520,I540614,);
not I_31641 (I540622,I668116);
DFFARX1 I_31642 (I668113,I2683,I540520,I540648,);
not I_31643 (I540656,I540648);
nor I_31644 (I540673,I540656,I540554);
and I_31645 (I540690,I540673,I668116);
nor I_31646 (I540707,I540656,I540622);
nor I_31647 (I540503,I540614,I540707);
DFFARX1 I_31648 (I668107,I2683,I540520,I540747,);
nor I_31649 (I540755,I540747,I540614);
not I_31650 (I540772,I540755);
not I_31651 (I540789,I540747);
nor I_31652 (I540806,I540789,I540690);
DFFARX1 I_31653 (I540806,I2683,I540520,I540506,);
nand I_31654 (I540837,I668107,I668110);
and I_31655 (I540854,I540837,I668113);
DFFARX1 I_31656 (I540854,I2683,I540520,I540880,);
nor I_31657 (I540888,I540880,I540747);
DFFARX1 I_31658 (I540888,I2683,I540520,I540488,);
nand I_31659 (I540919,I540880,I540789);
nand I_31660 (I540497,I540772,I540919);
not I_31661 (I540950,I540880);
nor I_31662 (I540967,I540950,I540690);
DFFARX1 I_31663 (I540967,I2683,I540520,I540509,);
nor I_31664 (I540998,I668119,I668110);
or I_31665 (I540500,I540747,I540998);
nor I_31666 (I540491,I540880,I540998);
or I_31667 (I540494,I540614,I540998);
DFFARX1 I_31668 (I540998,I2683,I540520,I540512,);
not I_31669 (I541098,I2690);
DFFARX1 I_31670 (I344827,I2683,I541098,I541124,);
not I_31671 (I541132,I541124);
nand I_31672 (I541149,I344818,I344836);
and I_31673 (I541166,I541149,I344839);
DFFARX1 I_31674 (I541166,I2683,I541098,I541192,);
not I_31675 (I541200,I344833);
DFFARX1 I_31676 (I344821,I2683,I541098,I541226,);
not I_31677 (I541234,I541226);
nor I_31678 (I541251,I541234,I541132);
and I_31679 (I541268,I541251,I344833);
nor I_31680 (I541285,I541234,I541200);
nor I_31681 (I541081,I541192,I541285);
DFFARX1 I_31682 (I344830,I2683,I541098,I541325,);
nor I_31683 (I541333,I541325,I541192);
not I_31684 (I541350,I541333);
not I_31685 (I541367,I541325);
nor I_31686 (I541384,I541367,I541268);
DFFARX1 I_31687 (I541384,I2683,I541098,I541084,);
nand I_31688 (I541415,I344845,I344842);
and I_31689 (I541432,I541415,I344824);
DFFARX1 I_31690 (I541432,I2683,I541098,I541458,);
nor I_31691 (I541466,I541458,I541325);
DFFARX1 I_31692 (I541466,I2683,I541098,I541066,);
nand I_31693 (I541497,I541458,I541367);
nand I_31694 (I541075,I541350,I541497);
not I_31695 (I541528,I541458);
nor I_31696 (I541545,I541528,I541268);
DFFARX1 I_31697 (I541545,I2683,I541098,I541087,);
nor I_31698 (I541576,I344818,I344842);
or I_31699 (I541078,I541325,I541576);
nor I_31700 (I541069,I541458,I541576);
or I_31701 (I541072,I541192,I541576);
DFFARX1 I_31702 (I541576,I2683,I541098,I541090,);
not I_31703 (I541676,I2690);
DFFARX1 I_31704 (I672865,I2683,I541676,I541702,);
not I_31705 (I541710,I541702);
nand I_31706 (I541727,I672853,I672871);
and I_31707 (I541744,I541727,I672868);
DFFARX1 I_31708 (I541744,I2683,I541676,I541770,);
not I_31709 (I541778,I672859);
DFFARX1 I_31710 (I672856,I2683,I541676,I541804,);
not I_31711 (I541812,I541804);
nor I_31712 (I541829,I541812,I541710);
and I_31713 (I541846,I541829,I672859);
nor I_31714 (I541863,I541812,I541778);
nor I_31715 (I541659,I541770,I541863);
DFFARX1 I_31716 (I672850,I2683,I541676,I541903,);
nor I_31717 (I541911,I541903,I541770);
not I_31718 (I541928,I541911);
not I_31719 (I541945,I541903);
nor I_31720 (I541962,I541945,I541846);
DFFARX1 I_31721 (I541962,I2683,I541676,I541662,);
nand I_31722 (I541993,I672850,I672853);
and I_31723 (I542010,I541993,I672856);
DFFARX1 I_31724 (I542010,I2683,I541676,I542036,);
nor I_31725 (I542044,I542036,I541903);
DFFARX1 I_31726 (I542044,I2683,I541676,I541644,);
nand I_31727 (I542075,I542036,I541945);
nand I_31728 (I541653,I541928,I542075);
not I_31729 (I542106,I542036);
nor I_31730 (I542123,I542106,I541846);
DFFARX1 I_31731 (I542123,I2683,I541676,I541665,);
nor I_31732 (I542154,I672862,I672853);
or I_31733 (I541656,I541903,I542154);
nor I_31734 (I541647,I542036,I542154);
or I_31735 (I541650,I541770,I542154);
DFFARX1 I_31736 (I542154,I2683,I541676,I541668,);
not I_31737 (I542254,I2690);
DFFARX1 I_31738 (I22170,I2683,I542254,I542280,);
not I_31739 (I542288,I542280);
nand I_31740 (I542305,I22167,I22158);
and I_31741 (I542322,I542305,I22158);
DFFARX1 I_31742 (I542322,I2683,I542254,I542348,);
not I_31743 (I542356,I22161);
DFFARX1 I_31744 (I22176,I2683,I542254,I542382,);
not I_31745 (I542390,I542382);
nor I_31746 (I542407,I542390,I542288);
and I_31747 (I542424,I542407,I22161);
nor I_31748 (I542441,I542390,I542356);
nor I_31749 (I542237,I542348,I542441);
DFFARX1 I_31750 (I22161,I2683,I542254,I542481,);
nor I_31751 (I542489,I542481,I542348);
not I_31752 (I542506,I542489);
not I_31753 (I542523,I542481);
nor I_31754 (I542540,I542523,I542424);
DFFARX1 I_31755 (I542540,I2683,I542254,I542240,);
nand I_31756 (I542571,I22179,I22164);
and I_31757 (I542588,I542571,I22182);
DFFARX1 I_31758 (I542588,I2683,I542254,I542614,);
nor I_31759 (I542622,I542614,I542481);
DFFARX1 I_31760 (I542622,I2683,I542254,I542222,);
nand I_31761 (I542653,I542614,I542523);
nand I_31762 (I542231,I542506,I542653);
not I_31763 (I542684,I542614);
nor I_31764 (I542701,I542684,I542424);
DFFARX1 I_31765 (I542701,I2683,I542254,I542243,);
nor I_31766 (I542732,I22173,I22164);
or I_31767 (I542234,I542481,I542732);
nor I_31768 (I542225,I542614,I542732);
or I_31769 (I542228,I542348,I542732);
DFFARX1 I_31770 (I542732,I2683,I542254,I542246,);
not I_31771 (I542832,I2690);
DFFARX1 I_31772 (I1039431,I2683,I542832,I542858,);
not I_31773 (I542866,I542858);
nand I_31774 (I542883,I1039416,I1039404);
and I_31775 (I542900,I542883,I1039419);
DFFARX1 I_31776 (I542900,I2683,I542832,I542926,);
not I_31777 (I542934,I1039404);
DFFARX1 I_31778 (I1039422,I2683,I542832,I542960,);
not I_31779 (I542968,I542960);
nor I_31780 (I542985,I542968,I542866);
and I_31781 (I543002,I542985,I1039404);
nor I_31782 (I543019,I542968,I542934);
nor I_31783 (I542815,I542926,I543019);
DFFARX1 I_31784 (I1039410,I2683,I542832,I543059,);
nor I_31785 (I543067,I543059,I542926);
not I_31786 (I543084,I543067);
not I_31787 (I543101,I543059);
nor I_31788 (I543118,I543101,I543002);
DFFARX1 I_31789 (I543118,I2683,I542832,I542818,);
nand I_31790 (I543149,I1039407,I1039413);
and I_31791 (I543166,I543149,I1039428);
DFFARX1 I_31792 (I543166,I2683,I542832,I543192,);
nor I_31793 (I543200,I543192,I543059);
DFFARX1 I_31794 (I543200,I2683,I542832,I542800,);
nand I_31795 (I543231,I543192,I543101);
nand I_31796 (I542809,I543084,I543231);
not I_31797 (I543262,I543192);
nor I_31798 (I543279,I543262,I543002);
DFFARX1 I_31799 (I543279,I2683,I542832,I542821,);
nor I_31800 (I543310,I1039425,I1039413);
or I_31801 (I542812,I543059,I543310);
nor I_31802 (I542803,I543192,I543310);
or I_31803 (I542806,I542926,I543310);
DFFARX1 I_31804 (I543310,I2683,I542832,I542824,);
not I_31805 (I543410,I2690);
DFFARX1 I_31806 (I112287,I2683,I543410,I543436,);
not I_31807 (I543444,I543436);
nand I_31808 (I543461,I112302,I112275);
and I_31809 (I543478,I543461,I112290);
DFFARX1 I_31810 (I543478,I2683,I543410,I543504,);
not I_31811 (I543512,I112293);
DFFARX1 I_31812 (I112278,I2683,I543410,I543538,);
not I_31813 (I543546,I543538);
nor I_31814 (I543563,I543546,I543444);
and I_31815 (I543580,I543563,I112293);
nor I_31816 (I543597,I543546,I543512);
nor I_31817 (I543393,I543504,I543597);
DFFARX1 I_31818 (I112284,I2683,I543410,I543637,);
nor I_31819 (I543645,I543637,I543504);
not I_31820 (I543662,I543645);
not I_31821 (I543679,I543637);
nor I_31822 (I543696,I543679,I543580);
DFFARX1 I_31823 (I543696,I2683,I543410,I543396,);
nand I_31824 (I543727,I112299,I112281);
and I_31825 (I543744,I543727,I112296);
DFFARX1 I_31826 (I543744,I2683,I543410,I543770,);
nor I_31827 (I543778,I543770,I543637);
DFFARX1 I_31828 (I543778,I2683,I543410,I543378,);
nand I_31829 (I543809,I543770,I543679);
nand I_31830 (I543387,I543662,I543809);
not I_31831 (I543840,I543770);
nor I_31832 (I543857,I543840,I543580);
DFFARX1 I_31833 (I543857,I2683,I543410,I543399,);
nor I_31834 (I543888,I112275,I112281);
or I_31835 (I543390,I543637,I543888);
nor I_31836 (I543381,I543770,I543888);
or I_31837 (I543384,I543504,I543888);
DFFARX1 I_31838 (I543888,I2683,I543410,I543402,);
not I_31839 (I543988,I2690);
DFFARX1 I_31840 (I633867,I2683,I543988,I544014,);
not I_31841 (I544022,I544014);
nand I_31842 (I544039,I633855,I633873);
and I_31843 (I544056,I544039,I633870);
DFFARX1 I_31844 (I544056,I2683,I543988,I544082,);
not I_31845 (I544090,I633861);
DFFARX1 I_31846 (I633858,I2683,I543988,I544116,);
not I_31847 (I544124,I544116);
nor I_31848 (I544141,I544124,I544022);
and I_31849 (I544158,I544141,I633861);
nor I_31850 (I544175,I544124,I544090);
nor I_31851 (I543971,I544082,I544175);
DFFARX1 I_31852 (I633852,I2683,I543988,I544215,);
nor I_31853 (I544223,I544215,I544082);
not I_31854 (I544240,I544223);
not I_31855 (I544257,I544215);
nor I_31856 (I544274,I544257,I544158);
DFFARX1 I_31857 (I544274,I2683,I543988,I543974,);
nand I_31858 (I544305,I633852,I633855);
and I_31859 (I544322,I544305,I633858);
DFFARX1 I_31860 (I544322,I2683,I543988,I544348,);
nor I_31861 (I544356,I544348,I544215);
DFFARX1 I_31862 (I544356,I2683,I543988,I543956,);
nand I_31863 (I544387,I544348,I544257);
nand I_31864 (I543965,I544240,I544387);
not I_31865 (I544418,I544348);
nor I_31866 (I544435,I544418,I544158);
DFFARX1 I_31867 (I544435,I2683,I543988,I543977,);
nor I_31868 (I544466,I633864,I633855);
or I_31869 (I543968,I544215,I544466);
nor I_31870 (I543959,I544348,I544466);
or I_31871 (I543962,I544082,I544466);
DFFARX1 I_31872 (I544466,I2683,I543988,I543980,);
not I_31873 (I544566,I2690);
DFFARX1 I_31874 (I1011116,I2683,I544566,I544592,);
not I_31875 (I544600,I544592);
nand I_31876 (I544617,I1011140,I1011122);
and I_31877 (I544634,I544617,I1011128);
DFFARX1 I_31878 (I544634,I2683,I544566,I544660,);
not I_31879 (I544668,I1011134);
DFFARX1 I_31880 (I1011119,I2683,I544566,I544694,);
not I_31881 (I544702,I544694);
nor I_31882 (I544719,I544702,I544600);
and I_31883 (I544736,I544719,I1011134);
nor I_31884 (I544753,I544702,I544668);
nor I_31885 (I544549,I544660,I544753);
DFFARX1 I_31886 (I1011131,I2683,I544566,I544793,);
nor I_31887 (I544801,I544793,I544660);
not I_31888 (I544818,I544801);
not I_31889 (I544835,I544793);
nor I_31890 (I544852,I544835,I544736);
DFFARX1 I_31891 (I544852,I2683,I544566,I544552,);
nand I_31892 (I544883,I1011137,I1011125);
and I_31893 (I544900,I544883,I1011119);
DFFARX1 I_31894 (I544900,I2683,I544566,I544926,);
nor I_31895 (I544934,I544926,I544793);
DFFARX1 I_31896 (I544934,I2683,I544566,I544534,);
nand I_31897 (I544965,I544926,I544835);
nand I_31898 (I544543,I544818,I544965);
not I_31899 (I544996,I544926);
nor I_31900 (I545013,I544996,I544736);
DFFARX1 I_31901 (I545013,I2683,I544566,I544555,);
nor I_31902 (I545044,I1011116,I1011125);
or I_31903 (I544546,I544793,I545044);
nor I_31904 (I544537,I544926,I545044);
or I_31905 (I544540,I544660,I545044);
DFFARX1 I_31906 (I545044,I2683,I544566,I544558,);
not I_31907 (I545144,I2690);
DFFARX1 I_31908 (I1084056,I2683,I545144,I545170,);
not I_31909 (I545178,I545170);
nand I_31910 (I545195,I1084041,I1084029);
and I_31911 (I545212,I545195,I1084044);
DFFARX1 I_31912 (I545212,I2683,I545144,I545238,);
not I_31913 (I545246,I1084029);
DFFARX1 I_31914 (I1084047,I2683,I545144,I545272,);
not I_31915 (I545280,I545272);
nor I_31916 (I545297,I545280,I545178);
and I_31917 (I545314,I545297,I1084029);
nor I_31918 (I545331,I545280,I545246);
nor I_31919 (I545127,I545238,I545331);
DFFARX1 I_31920 (I1084035,I2683,I545144,I545371,);
nor I_31921 (I545379,I545371,I545238);
not I_31922 (I545396,I545379);
not I_31923 (I545413,I545371);
nor I_31924 (I545430,I545413,I545314);
DFFARX1 I_31925 (I545430,I2683,I545144,I545130,);
nand I_31926 (I545461,I1084032,I1084038);
and I_31927 (I545478,I545461,I1084053);
DFFARX1 I_31928 (I545478,I2683,I545144,I545504,);
nor I_31929 (I545512,I545504,I545371);
DFFARX1 I_31930 (I545512,I2683,I545144,I545112,);
nand I_31931 (I545543,I545504,I545413);
nand I_31932 (I545121,I545396,I545543);
not I_31933 (I545574,I545504);
nor I_31934 (I545591,I545574,I545314);
DFFARX1 I_31935 (I545591,I2683,I545144,I545133,);
nor I_31936 (I545622,I1084050,I1084038);
or I_31937 (I545124,I545371,I545622);
nor I_31938 (I545115,I545504,I545622);
or I_31939 (I545118,I545238,I545622);
DFFARX1 I_31940 (I545622,I2683,I545144,I545136,);
not I_31941 (I545722,I2690);
DFFARX1 I_31942 (I290714,I2683,I545722,I545748,);
not I_31943 (I545756,I545748);
nand I_31944 (I545773,I290717,I290693);
and I_31945 (I545790,I545773,I290690);
DFFARX1 I_31946 (I545790,I2683,I545722,I545816,);
not I_31947 (I545824,I290696);
DFFARX1 I_31948 (I290690,I2683,I545722,I545850,);
not I_31949 (I545858,I545850);
nor I_31950 (I545875,I545858,I545756);
and I_31951 (I545892,I545875,I290696);
nor I_31952 (I545909,I545858,I545824);
nor I_31953 (I545705,I545816,I545909);
DFFARX1 I_31954 (I290699,I2683,I545722,I545949,);
nor I_31955 (I545957,I545949,I545816);
not I_31956 (I545974,I545957);
not I_31957 (I545991,I545949);
nor I_31958 (I546008,I545991,I545892);
DFFARX1 I_31959 (I546008,I2683,I545722,I545708,);
nand I_31960 (I546039,I290702,I290711);
and I_31961 (I546056,I546039,I290708);
DFFARX1 I_31962 (I546056,I2683,I545722,I546082,);
nor I_31963 (I546090,I546082,I545949);
DFFARX1 I_31964 (I546090,I2683,I545722,I545690,);
nand I_31965 (I546121,I546082,I545991);
nand I_31966 (I545699,I545974,I546121);
not I_31967 (I546152,I546082);
nor I_31968 (I546169,I546152,I545892);
DFFARX1 I_31969 (I546169,I2683,I545722,I545711,);
nor I_31970 (I546200,I290705,I290711);
or I_31971 (I545702,I545949,I546200);
nor I_31972 (I545693,I546082,I546200);
or I_31973 (I545696,I545816,I546200);
DFFARX1 I_31974 (I546200,I2683,I545722,I545714,);
not I_31975 (I546300,I2690);
DFFARX1 I_31976 (I446274,I2683,I546300,I546326,);
not I_31977 (I546334,I546326);
nand I_31978 (I546351,I446283,I446292);
and I_31979 (I546368,I546351,I446298);
DFFARX1 I_31980 (I546368,I2683,I546300,I546394,);
not I_31981 (I546402,I446295);
DFFARX1 I_31982 (I446280,I2683,I546300,I546428,);
not I_31983 (I546436,I546428);
nor I_31984 (I546453,I546436,I546334);
and I_31985 (I546470,I546453,I446295);
nor I_31986 (I546487,I546436,I546402);
nor I_31987 (I546283,I546394,I546487);
DFFARX1 I_31988 (I446289,I2683,I546300,I546527,);
nor I_31989 (I546535,I546527,I546394);
not I_31990 (I546552,I546535);
not I_31991 (I546569,I546527);
nor I_31992 (I546586,I546569,I546470);
DFFARX1 I_31993 (I546586,I2683,I546300,I546286,);
nand I_31994 (I546617,I446286,I446277);
and I_31995 (I546634,I546617,I446274);
DFFARX1 I_31996 (I546634,I2683,I546300,I546660,);
nor I_31997 (I546668,I546660,I546527);
DFFARX1 I_31998 (I546668,I2683,I546300,I546268,);
nand I_31999 (I546699,I546660,I546569);
nand I_32000 (I546277,I546552,I546699);
not I_32001 (I546730,I546660);
nor I_32002 (I546747,I546730,I546470);
DFFARX1 I_32003 (I546747,I2683,I546300,I546289,);
nor I_32004 (I546778,I446277,I446277);
or I_32005 (I546280,I546527,I546778);
nor I_32006 (I546271,I546660,I546778);
or I_32007 (I546274,I546394,I546778);
DFFARX1 I_32008 (I546778,I2683,I546300,I546292,);
not I_32009 (I546878,I2690);
DFFARX1 I_32010 (I445696,I2683,I546878,I546904,);
not I_32011 (I546912,I546904);
nand I_32012 (I546929,I445705,I445714);
and I_32013 (I546946,I546929,I445720);
DFFARX1 I_32014 (I546946,I2683,I546878,I546972,);
not I_32015 (I546980,I445717);
DFFARX1 I_32016 (I445702,I2683,I546878,I547006,);
not I_32017 (I547014,I547006);
nor I_32018 (I547031,I547014,I546912);
and I_32019 (I547048,I547031,I445717);
nor I_32020 (I547065,I547014,I546980);
nor I_32021 (I546861,I546972,I547065);
DFFARX1 I_32022 (I445711,I2683,I546878,I547105,);
nor I_32023 (I547113,I547105,I546972);
not I_32024 (I547130,I547113);
not I_32025 (I547147,I547105);
nor I_32026 (I547164,I547147,I547048);
DFFARX1 I_32027 (I547164,I2683,I546878,I546864,);
nand I_32028 (I547195,I445708,I445699);
and I_32029 (I547212,I547195,I445696);
DFFARX1 I_32030 (I547212,I2683,I546878,I547238,);
nor I_32031 (I547246,I547238,I547105);
DFFARX1 I_32032 (I547246,I2683,I546878,I546846,);
nand I_32033 (I547277,I547238,I547147);
nand I_32034 (I546855,I547130,I547277);
not I_32035 (I547308,I547238);
nor I_32036 (I547325,I547308,I547048);
DFFARX1 I_32037 (I547325,I2683,I546878,I546867,);
nor I_32038 (I547356,I445699,I445699);
or I_32039 (I546858,I547105,I547356);
nor I_32040 (I546849,I547238,I547356);
or I_32041 (I546852,I546972,I547356);
DFFARX1 I_32042 (I547356,I2683,I546878,I546870,);
not I_32043 (I547456,I2690);
DFFARX1 I_32044 (I131315,I2683,I547456,I547482,);
not I_32045 (I547490,I547482);
nand I_32046 (I547507,I131318,I131339);
and I_32047 (I547524,I547507,I131327);
DFFARX1 I_32048 (I547524,I2683,I547456,I547550,);
not I_32049 (I547558,I131324);
DFFARX1 I_32050 (I131315,I2683,I547456,I547584,);
not I_32051 (I547592,I547584);
nor I_32052 (I547609,I547592,I547490);
and I_32053 (I547626,I547609,I131324);
nor I_32054 (I547643,I547592,I547558);
nor I_32055 (I547439,I547550,I547643);
DFFARX1 I_32056 (I131333,I2683,I547456,I547683,);
nor I_32057 (I547691,I547683,I547550);
not I_32058 (I547708,I547691);
not I_32059 (I547725,I547683);
nor I_32060 (I547742,I547725,I547626);
DFFARX1 I_32061 (I547742,I2683,I547456,I547442,);
nand I_32062 (I547773,I131318,I131321);
and I_32063 (I547790,I547773,I131330);
DFFARX1 I_32064 (I547790,I2683,I547456,I547816,);
nor I_32065 (I547824,I547816,I547683);
DFFARX1 I_32066 (I547824,I2683,I547456,I547424,);
nand I_32067 (I547855,I547816,I547725);
nand I_32068 (I547433,I547708,I547855);
not I_32069 (I547886,I547816);
nor I_32070 (I547903,I547886,I547626);
DFFARX1 I_32071 (I547903,I2683,I547456,I547445,);
nor I_32072 (I547934,I131336,I131321);
or I_32073 (I547436,I547683,I547934);
nor I_32074 (I547427,I547816,I547934);
or I_32075 (I547430,I547550,I547934);
DFFARX1 I_32076 (I547934,I2683,I547456,I547448,);
not I_32077 (I548034,I2690);
DFFARX1 I_32078 (I341563,I2683,I548034,I548060,);
not I_32079 (I548068,I548060);
nand I_32080 (I548085,I341554,I341572);
and I_32081 (I548102,I548085,I341575);
DFFARX1 I_32082 (I548102,I2683,I548034,I548128,);
not I_32083 (I548136,I341569);
DFFARX1 I_32084 (I341557,I2683,I548034,I548162,);
not I_32085 (I548170,I548162);
nor I_32086 (I548187,I548170,I548068);
and I_32087 (I548204,I548187,I341569);
nor I_32088 (I548221,I548170,I548136);
nor I_32089 (I548017,I548128,I548221);
DFFARX1 I_32090 (I341566,I2683,I548034,I548261,);
nor I_32091 (I548269,I548261,I548128);
not I_32092 (I548286,I548269);
not I_32093 (I548303,I548261);
nor I_32094 (I548320,I548303,I548204);
DFFARX1 I_32095 (I548320,I2683,I548034,I548020,);
nand I_32096 (I548351,I341581,I341578);
and I_32097 (I548368,I548351,I341560);
DFFARX1 I_32098 (I548368,I2683,I548034,I548394,);
nor I_32099 (I548402,I548394,I548261);
DFFARX1 I_32100 (I548402,I2683,I548034,I548002,);
nand I_32101 (I548433,I548394,I548303);
nand I_32102 (I548011,I548286,I548433);
not I_32103 (I548464,I548394);
nor I_32104 (I548481,I548464,I548204);
DFFARX1 I_32105 (I548481,I2683,I548034,I548023,);
nor I_32106 (I548512,I341554,I341578);
or I_32107 (I548014,I548261,I548512);
nor I_32108 (I548005,I548394,I548512);
or I_32109 (I548008,I548128,I548512);
DFFARX1 I_32110 (I548512,I2683,I548034,I548026,);
not I_32111 (I548612,I2690);
DFFARX1 I_32112 (I374747,I2683,I548612,I548638,);
not I_32113 (I548646,I548638);
nand I_32114 (I548663,I374738,I374756);
and I_32115 (I548680,I548663,I374759);
DFFARX1 I_32116 (I548680,I2683,I548612,I548706,);
not I_32117 (I548714,I374753);
DFFARX1 I_32118 (I374741,I2683,I548612,I548740,);
not I_32119 (I548748,I548740);
nor I_32120 (I548765,I548748,I548646);
and I_32121 (I548782,I548765,I374753);
nor I_32122 (I548799,I548748,I548714);
nor I_32123 (I548595,I548706,I548799);
DFFARX1 I_32124 (I374750,I2683,I548612,I548839,);
nor I_32125 (I548847,I548839,I548706);
not I_32126 (I548864,I548847);
not I_32127 (I548881,I548839);
nor I_32128 (I548898,I548881,I548782);
DFFARX1 I_32129 (I548898,I2683,I548612,I548598,);
nand I_32130 (I548929,I374765,I374762);
and I_32131 (I548946,I548929,I374744);
DFFARX1 I_32132 (I548946,I2683,I548612,I548972,);
nor I_32133 (I548980,I548972,I548839);
DFFARX1 I_32134 (I548980,I2683,I548612,I548580,);
nand I_32135 (I549011,I548972,I548881);
nand I_32136 (I548589,I548864,I549011);
not I_32137 (I549042,I548972);
nor I_32138 (I549059,I549042,I548782);
DFFARX1 I_32139 (I549059,I2683,I548612,I548601,);
nor I_32140 (I549090,I374738,I374762);
or I_32141 (I548592,I548839,I549090);
nor I_32142 (I548583,I548972,I549090);
or I_32143 (I548586,I548706,I549090);
DFFARX1 I_32144 (I549090,I2683,I548612,I548604,);
not I_32145 (I549190,I2690);
DFFARX1 I_32146 (I343739,I2683,I549190,I549216,);
not I_32147 (I549224,I549216);
nand I_32148 (I549241,I343730,I343748);
and I_32149 (I549258,I549241,I343751);
DFFARX1 I_32150 (I549258,I2683,I549190,I549284,);
not I_32151 (I549292,I343745);
DFFARX1 I_32152 (I343733,I2683,I549190,I549318,);
not I_32153 (I549326,I549318);
nor I_32154 (I549343,I549326,I549224);
and I_32155 (I549360,I549343,I343745);
nor I_32156 (I549377,I549326,I549292);
nor I_32157 (I549173,I549284,I549377);
DFFARX1 I_32158 (I343742,I2683,I549190,I549417,);
nor I_32159 (I549425,I549417,I549284);
not I_32160 (I549442,I549425);
not I_32161 (I549459,I549417);
nor I_32162 (I549476,I549459,I549360);
DFFARX1 I_32163 (I549476,I2683,I549190,I549176,);
nand I_32164 (I549507,I343757,I343754);
and I_32165 (I549524,I549507,I343736);
DFFARX1 I_32166 (I549524,I2683,I549190,I549550,);
nor I_32167 (I549558,I549550,I549417);
DFFARX1 I_32168 (I549558,I2683,I549190,I549158,);
nand I_32169 (I549589,I549550,I549459);
nand I_32170 (I549167,I549442,I549589);
not I_32171 (I549620,I549550);
nor I_32172 (I549637,I549620,I549360);
DFFARX1 I_32173 (I549637,I2683,I549190,I549179,);
nor I_32174 (I549668,I343730,I343754);
or I_32175 (I549170,I549417,I549668);
nor I_32176 (I549161,I549550,I549668);
or I_32177 (I549164,I549284,I549668);
DFFARX1 I_32178 (I549668,I2683,I549190,I549182,);
not I_32179 (I549768,I2690);
DFFARX1 I_32180 (I924162,I2683,I549768,I549794,);
not I_32181 (I549802,I549794);
nand I_32182 (I549819,I924144,I924156);
and I_32183 (I549836,I549819,I924159);
DFFARX1 I_32184 (I549836,I2683,I549768,I549862,);
not I_32185 (I549870,I924153);
DFFARX1 I_32186 (I924150,I2683,I549768,I549896,);
not I_32187 (I549904,I549896);
nor I_32188 (I549921,I549904,I549802);
and I_32189 (I549938,I549921,I924153);
nor I_32190 (I549955,I549904,I549870);
nor I_32191 (I549751,I549862,I549955);
DFFARX1 I_32192 (I924168,I2683,I549768,I549995,);
nor I_32193 (I550003,I549995,I549862);
not I_32194 (I550020,I550003);
not I_32195 (I550037,I549995);
nor I_32196 (I550054,I550037,I549938);
DFFARX1 I_32197 (I550054,I2683,I549768,I549754,);
nand I_32198 (I550085,I924147,I924147);
and I_32199 (I550102,I550085,I924144);
DFFARX1 I_32200 (I550102,I2683,I549768,I550128,);
nor I_32201 (I550136,I550128,I549995);
DFFARX1 I_32202 (I550136,I2683,I549768,I549736,);
nand I_32203 (I550167,I550128,I550037);
nand I_32204 (I549745,I550020,I550167);
not I_32205 (I550198,I550128);
nor I_32206 (I550215,I550198,I549938);
DFFARX1 I_32207 (I550215,I2683,I549768,I549757,);
nor I_32208 (I550246,I924165,I924147);
or I_32209 (I549748,I549995,I550246);
nor I_32210 (I549739,I550128,I550246);
or I_32211 (I549742,I549862,I550246);
DFFARX1 I_32212 (I550246,I2683,I549768,I549760,);
not I_32213 (I550346,I2690);
DFFARX1 I_32214 (I190815,I2683,I550346,I550372,);
not I_32215 (I550380,I550372);
nand I_32216 (I550397,I190818,I190839);
and I_32217 (I550414,I550397,I190827);
DFFARX1 I_32218 (I550414,I2683,I550346,I550440,);
not I_32219 (I550448,I190824);
DFFARX1 I_32220 (I190815,I2683,I550346,I550474,);
not I_32221 (I550482,I550474);
nor I_32222 (I550499,I550482,I550380);
and I_32223 (I550516,I550499,I190824);
nor I_32224 (I550533,I550482,I550448);
nor I_32225 (I550329,I550440,I550533);
DFFARX1 I_32226 (I190833,I2683,I550346,I550573,);
nor I_32227 (I550581,I550573,I550440);
not I_32228 (I550598,I550581);
not I_32229 (I550615,I550573);
nor I_32230 (I550632,I550615,I550516);
DFFARX1 I_32231 (I550632,I2683,I550346,I550332,);
nand I_32232 (I550663,I190818,I190821);
and I_32233 (I550680,I550663,I190830);
DFFARX1 I_32234 (I550680,I2683,I550346,I550706,);
nor I_32235 (I550714,I550706,I550573);
DFFARX1 I_32236 (I550714,I2683,I550346,I550314,);
nand I_32237 (I550745,I550706,I550615);
nand I_32238 (I550323,I550598,I550745);
not I_32239 (I550776,I550706);
nor I_32240 (I550793,I550776,I550516);
DFFARX1 I_32241 (I550793,I2683,I550346,I550335,);
nor I_32242 (I550824,I190836,I190821);
or I_32243 (I550326,I550573,I550824);
nor I_32244 (I550317,I550706,I550824);
or I_32245 (I550320,I550440,I550824);
DFFARX1 I_32246 (I550824,I2683,I550346,I550338,);
not I_32247 (I550924,I2690);
DFFARX1 I_32248 (I904510,I2683,I550924,I550950,);
not I_32249 (I550958,I550950);
nand I_32250 (I550975,I904492,I904504);
and I_32251 (I550992,I550975,I904507);
DFFARX1 I_32252 (I550992,I2683,I550924,I551018,);
not I_32253 (I551026,I904501);
DFFARX1 I_32254 (I904498,I2683,I550924,I551052,);
not I_32255 (I551060,I551052);
nor I_32256 (I551077,I551060,I550958);
and I_32257 (I551094,I551077,I904501);
nor I_32258 (I551111,I551060,I551026);
nor I_32259 (I550907,I551018,I551111);
DFFARX1 I_32260 (I904516,I2683,I550924,I551151,);
nor I_32261 (I551159,I551151,I551018);
not I_32262 (I551176,I551159);
not I_32263 (I551193,I551151);
nor I_32264 (I551210,I551193,I551094);
DFFARX1 I_32265 (I551210,I2683,I550924,I550910,);
nand I_32266 (I551241,I904495,I904495);
and I_32267 (I551258,I551241,I904492);
DFFARX1 I_32268 (I551258,I2683,I550924,I551284,);
nor I_32269 (I551292,I551284,I551151);
DFFARX1 I_32270 (I551292,I2683,I550924,I550892,);
nand I_32271 (I551323,I551284,I551193);
nand I_32272 (I550901,I551176,I551323);
not I_32273 (I551354,I551284);
nor I_32274 (I551371,I551354,I551094);
DFFARX1 I_32275 (I551371,I2683,I550924,I550913,);
nor I_32276 (I551402,I904513,I904495);
or I_32277 (I550904,I551151,I551402);
nor I_32278 (I550895,I551284,I551402);
or I_32279 (I550898,I551018,I551402);
DFFARX1 I_32280 (I551402,I2683,I550924,I550916,);
not I_32281 (I551502,I2690);
DFFARX1 I_32282 (I184865,I2683,I551502,I551528,);
not I_32283 (I551536,I551528);
nand I_32284 (I551553,I184868,I184889);
and I_32285 (I551570,I551553,I184877);
DFFARX1 I_32286 (I551570,I2683,I551502,I551596,);
not I_32287 (I551604,I184874);
DFFARX1 I_32288 (I184865,I2683,I551502,I551630,);
not I_32289 (I551638,I551630);
nor I_32290 (I551655,I551638,I551536);
and I_32291 (I551672,I551655,I184874);
nor I_32292 (I551689,I551638,I551604);
nor I_32293 (I551485,I551596,I551689);
DFFARX1 I_32294 (I184883,I2683,I551502,I551729,);
nor I_32295 (I551737,I551729,I551596);
not I_32296 (I551754,I551737);
not I_32297 (I551771,I551729);
nor I_32298 (I551788,I551771,I551672);
DFFARX1 I_32299 (I551788,I2683,I551502,I551488,);
nand I_32300 (I551819,I184868,I184871);
and I_32301 (I551836,I551819,I184880);
DFFARX1 I_32302 (I551836,I2683,I551502,I551862,);
nor I_32303 (I551870,I551862,I551729);
DFFARX1 I_32304 (I551870,I2683,I551502,I551470,);
nand I_32305 (I551901,I551862,I551771);
nand I_32306 (I551479,I551754,I551901);
not I_32307 (I551932,I551862);
nor I_32308 (I551949,I551932,I551672);
DFFARX1 I_32309 (I551949,I2683,I551502,I551491,);
nor I_32310 (I551980,I184886,I184871);
or I_32311 (I551482,I551729,I551980);
nor I_32312 (I551473,I551862,I551980);
or I_32313 (I551476,I551596,I551980);
DFFARX1 I_32314 (I551980,I2683,I551502,I551494,);
not I_32315 (I552080,I2690);
DFFARX1 I_32316 (I323067,I2683,I552080,I552106,);
not I_32317 (I552114,I552106);
nand I_32318 (I552131,I323058,I323076);
and I_32319 (I552148,I552131,I323079);
DFFARX1 I_32320 (I552148,I2683,I552080,I552174,);
not I_32321 (I552182,I323073);
DFFARX1 I_32322 (I323061,I2683,I552080,I552208,);
not I_32323 (I552216,I552208);
nor I_32324 (I552233,I552216,I552114);
and I_32325 (I552250,I552233,I323073);
nor I_32326 (I552267,I552216,I552182);
nor I_32327 (I552063,I552174,I552267);
DFFARX1 I_32328 (I323070,I2683,I552080,I552307,);
nor I_32329 (I552315,I552307,I552174);
not I_32330 (I552332,I552315);
not I_32331 (I552349,I552307);
nor I_32332 (I552366,I552349,I552250);
DFFARX1 I_32333 (I552366,I2683,I552080,I552066,);
nand I_32334 (I552397,I323085,I323082);
and I_32335 (I552414,I552397,I323064);
DFFARX1 I_32336 (I552414,I2683,I552080,I552440,);
nor I_32337 (I552448,I552440,I552307);
DFFARX1 I_32338 (I552448,I2683,I552080,I552048,);
nand I_32339 (I552479,I552440,I552349);
nand I_32340 (I552057,I552332,I552479);
not I_32341 (I552510,I552440);
nor I_32342 (I552527,I552510,I552250);
DFFARX1 I_32343 (I552527,I2683,I552080,I552069,);
nor I_32344 (I552558,I323058,I323082);
or I_32345 (I552060,I552307,I552558);
nor I_32346 (I552051,I552440,I552558);
or I_32347 (I552054,I552174,I552558);
DFFARX1 I_32348 (I552558,I2683,I552080,I552072,);
not I_32349 (I552658,I2690);
DFFARX1 I_32350 (I104900,I2683,I552658,I552684,);
not I_32351 (I552692,I552684);
nand I_32352 (I552709,I104909,I104918);
and I_32353 (I552726,I552709,I104897);
DFFARX1 I_32354 (I552726,I2683,I552658,I552752,);
not I_32355 (I552760,I104900);
DFFARX1 I_32356 (I104915,I2683,I552658,I552786,);
not I_32357 (I552794,I552786);
nor I_32358 (I552811,I552794,I552692);
and I_32359 (I552828,I552811,I104900);
nor I_32360 (I552845,I552794,I552760);
nor I_32361 (I552641,I552752,I552845);
DFFARX1 I_32362 (I104906,I2683,I552658,I552885,);
nor I_32363 (I552893,I552885,I552752);
not I_32364 (I552910,I552893);
not I_32365 (I552927,I552885);
nor I_32366 (I552944,I552927,I552828);
DFFARX1 I_32367 (I552944,I2683,I552658,I552644,);
nand I_32368 (I552975,I104921,I104897);
and I_32369 (I552992,I552975,I104903);
DFFARX1 I_32370 (I552992,I2683,I552658,I553018,);
nor I_32371 (I553026,I553018,I552885);
DFFARX1 I_32372 (I553026,I2683,I552658,I552626,);
nand I_32373 (I553057,I553018,I552927);
nand I_32374 (I552635,I552910,I553057);
not I_32375 (I553088,I553018);
nor I_32376 (I553105,I553088,I552828);
DFFARX1 I_32377 (I553105,I2683,I552658,I552647,);
nor I_32378 (I553136,I104912,I104897);
or I_32379 (I552638,I552885,I553136);
nor I_32380 (I552629,I553018,I553136);
or I_32381 (I552632,I552752,I553136);
DFFARX1 I_32382 (I553136,I2683,I552658,I552650,);
not I_32383 (I553236,I2690);
DFFARX1 I_32384 (I309686,I2683,I553236,I553262,);
not I_32385 (I553270,I553262);
nand I_32386 (I553287,I309689,I309665);
and I_32387 (I553304,I553287,I309662);
DFFARX1 I_32388 (I553304,I2683,I553236,I553330,);
not I_32389 (I553338,I309668);
DFFARX1 I_32390 (I309662,I2683,I553236,I553364,);
not I_32391 (I553372,I553364);
nor I_32392 (I553389,I553372,I553270);
and I_32393 (I553406,I553389,I309668);
nor I_32394 (I553423,I553372,I553338);
nor I_32395 (I553219,I553330,I553423);
DFFARX1 I_32396 (I309671,I2683,I553236,I553463,);
nor I_32397 (I553471,I553463,I553330);
not I_32398 (I553488,I553471);
not I_32399 (I553505,I553463);
nor I_32400 (I553522,I553505,I553406);
DFFARX1 I_32401 (I553522,I2683,I553236,I553222,);
nand I_32402 (I553553,I309674,I309683);
and I_32403 (I553570,I553553,I309680);
DFFARX1 I_32404 (I553570,I2683,I553236,I553596,);
nor I_32405 (I553604,I553596,I553463);
DFFARX1 I_32406 (I553604,I2683,I553236,I553204,);
nand I_32407 (I553635,I553596,I553505);
nand I_32408 (I553213,I553488,I553635);
not I_32409 (I553666,I553596);
nor I_32410 (I553683,I553666,I553406);
DFFARX1 I_32411 (I553683,I2683,I553236,I553225,);
nor I_32412 (I553714,I309677,I309683);
or I_32413 (I553216,I553463,I553714);
nor I_32414 (I553207,I553596,I553714);
or I_32415 (I553210,I553330,I553714);
DFFARX1 I_32416 (I553714,I2683,I553236,I553228,);
not I_32417 (I553814,I2690);
DFFARX1 I_32418 (I859426,I2683,I553814,I553840,);
not I_32419 (I553848,I553840);
nand I_32420 (I553865,I859408,I859420);
and I_32421 (I553882,I553865,I859423);
DFFARX1 I_32422 (I553882,I2683,I553814,I553908,);
not I_32423 (I553916,I859417);
DFFARX1 I_32424 (I859414,I2683,I553814,I553942,);
not I_32425 (I553950,I553942);
nor I_32426 (I553967,I553950,I553848);
and I_32427 (I553984,I553967,I859417);
nor I_32428 (I554001,I553950,I553916);
nor I_32429 (I553797,I553908,I554001);
DFFARX1 I_32430 (I859432,I2683,I553814,I554041,);
nor I_32431 (I554049,I554041,I553908);
not I_32432 (I554066,I554049);
not I_32433 (I554083,I554041);
nor I_32434 (I554100,I554083,I553984);
DFFARX1 I_32435 (I554100,I2683,I553814,I553800,);
nand I_32436 (I554131,I859411,I859411);
and I_32437 (I554148,I554131,I859408);
DFFARX1 I_32438 (I554148,I2683,I553814,I554174,);
nor I_32439 (I554182,I554174,I554041);
DFFARX1 I_32440 (I554182,I2683,I553814,I553782,);
nand I_32441 (I554213,I554174,I554083);
nand I_32442 (I553791,I554066,I554213);
not I_32443 (I554244,I554174);
nor I_32444 (I554261,I554244,I553984);
DFFARX1 I_32445 (I554261,I2683,I553814,I553803,);
nor I_32446 (I554292,I859429,I859411);
or I_32447 (I553794,I554041,I554292);
nor I_32448 (I553785,I554174,I554292);
or I_32449 (I553788,I553908,I554292);
DFFARX1 I_32450 (I554292,I2683,I553814,I553806,);
not I_32451 (I554392,I2690);
DFFARX1 I_32452 (I984222,I2683,I554392,I554418,);
not I_32453 (I554426,I554418);
nand I_32454 (I554443,I984225,I984234);
and I_32455 (I554460,I554443,I984237);
DFFARX1 I_32456 (I554460,I2683,I554392,I554486,);
not I_32457 (I554494,I984246);
DFFARX1 I_32458 (I984228,I2683,I554392,I554520,);
not I_32459 (I554528,I554520);
nor I_32460 (I554545,I554528,I554426);
and I_32461 (I554562,I554545,I984246);
nor I_32462 (I554579,I554528,I554494);
nor I_32463 (I554375,I554486,I554579);
DFFARX1 I_32464 (I984225,I2683,I554392,I554619,);
nor I_32465 (I554627,I554619,I554486);
not I_32466 (I554644,I554627);
not I_32467 (I554661,I554619);
nor I_32468 (I554678,I554661,I554562);
DFFARX1 I_32469 (I554678,I2683,I554392,I554378,);
nand I_32470 (I554709,I984243,I984222);
and I_32471 (I554726,I554709,I984240);
DFFARX1 I_32472 (I554726,I2683,I554392,I554752,);
nor I_32473 (I554760,I554752,I554619);
DFFARX1 I_32474 (I554760,I2683,I554392,I554360,);
nand I_32475 (I554791,I554752,I554661);
nand I_32476 (I554369,I554644,I554791);
not I_32477 (I554822,I554752);
nor I_32478 (I554839,I554822,I554562);
DFFARX1 I_32479 (I554839,I2683,I554392,I554381,);
nor I_32480 (I554870,I984231,I984222);
or I_32481 (I554372,I554619,I554870);
nor I_32482 (I554363,I554752,I554870);
or I_32483 (I554366,I554486,I554870);
DFFARX1 I_32484 (I554870,I2683,I554392,I554384,);
not I_32485 (I554970,I2690);
DFFARX1 I_32486 (I913180,I2683,I554970,I554996,);
not I_32487 (I555004,I554996);
nand I_32488 (I555021,I913162,I913174);
and I_32489 (I555038,I555021,I913177);
DFFARX1 I_32490 (I555038,I2683,I554970,I555064,);
not I_32491 (I555072,I913171);
DFFARX1 I_32492 (I913168,I2683,I554970,I555098,);
not I_32493 (I555106,I555098);
nor I_32494 (I555123,I555106,I555004);
and I_32495 (I555140,I555123,I913171);
nor I_32496 (I555157,I555106,I555072);
nor I_32497 (I554953,I555064,I555157);
DFFARX1 I_32498 (I913186,I2683,I554970,I555197,);
nor I_32499 (I555205,I555197,I555064);
not I_32500 (I555222,I555205);
not I_32501 (I555239,I555197);
nor I_32502 (I555256,I555239,I555140);
DFFARX1 I_32503 (I555256,I2683,I554970,I554956,);
nand I_32504 (I555287,I913165,I913165);
and I_32505 (I555304,I555287,I913162);
DFFARX1 I_32506 (I555304,I2683,I554970,I555330,);
nor I_32507 (I555338,I555330,I555197);
DFFARX1 I_32508 (I555338,I2683,I554970,I554938,);
nand I_32509 (I555369,I555330,I555239);
nand I_32510 (I554947,I555222,I555369);
not I_32511 (I555400,I555330);
nor I_32512 (I555417,I555400,I555140);
DFFARX1 I_32513 (I555417,I2683,I554970,I554959,);
nor I_32514 (I555448,I913183,I913165);
or I_32515 (I554950,I555197,I555448);
nor I_32516 (I554941,I555330,I555448);
or I_32517 (I554944,I555064,I555448);
DFFARX1 I_32518 (I555448,I2683,I554970,I554962,);
not I_32519 (I555548,I2690);
DFFARX1 I_32520 (I406817,I2683,I555548,I555574,);
not I_32521 (I555582,I555574);
nand I_32522 (I555599,I406832,I406817);
and I_32523 (I555616,I555599,I406820);
DFFARX1 I_32524 (I555616,I2683,I555548,I555642,);
not I_32525 (I555650,I406820);
DFFARX1 I_32526 (I406829,I2683,I555548,I555676,);
not I_32527 (I555684,I555676);
nor I_32528 (I555701,I555684,I555582);
and I_32529 (I555718,I555701,I406820);
nor I_32530 (I555735,I555684,I555650);
nor I_32531 (I555531,I555642,I555735);
DFFARX1 I_32532 (I406823,I2683,I555548,I555775,);
nor I_32533 (I555783,I555775,I555642);
not I_32534 (I555800,I555783);
not I_32535 (I555817,I555775);
nor I_32536 (I555834,I555817,I555718);
DFFARX1 I_32537 (I555834,I2683,I555548,I555534,);
nand I_32538 (I555865,I406826,I406835);
and I_32539 (I555882,I555865,I406841);
DFFARX1 I_32540 (I555882,I2683,I555548,I555908,);
nor I_32541 (I555916,I555908,I555775);
DFFARX1 I_32542 (I555916,I2683,I555548,I555516,);
nand I_32543 (I555947,I555908,I555817);
nand I_32544 (I555525,I555800,I555947);
not I_32545 (I555978,I555908);
nor I_32546 (I555995,I555978,I555718);
DFFARX1 I_32547 (I555995,I2683,I555548,I555537,);
nor I_32548 (I556026,I406838,I406835);
or I_32549 (I555528,I555775,I556026);
nor I_32550 (I555519,I555908,I556026);
or I_32551 (I555522,I555642,I556026);
DFFARX1 I_32552 (I556026,I2683,I555548,I555540,);
not I_32553 (I556126,I2690);
DFFARX1 I_32554 (I652839,I2683,I556126,I556152,);
not I_32555 (I556160,I556152);
nand I_32556 (I556177,I652827,I652845);
and I_32557 (I556194,I556177,I652842);
DFFARX1 I_32558 (I556194,I2683,I556126,I556220,);
not I_32559 (I556228,I652833);
DFFARX1 I_32560 (I652830,I2683,I556126,I556254,);
not I_32561 (I556262,I556254);
nor I_32562 (I556279,I556262,I556160);
and I_32563 (I556296,I556279,I652833);
nor I_32564 (I556313,I556262,I556228);
nor I_32565 (I556109,I556220,I556313);
DFFARX1 I_32566 (I652824,I2683,I556126,I556353,);
nor I_32567 (I556361,I556353,I556220);
not I_32568 (I556378,I556361);
not I_32569 (I556395,I556353);
nor I_32570 (I556412,I556395,I556296);
DFFARX1 I_32571 (I556412,I2683,I556126,I556112,);
nand I_32572 (I556443,I652824,I652827);
and I_32573 (I556460,I556443,I652830);
DFFARX1 I_32574 (I556460,I2683,I556126,I556486,);
nor I_32575 (I556494,I556486,I556353);
DFFARX1 I_32576 (I556494,I2683,I556126,I556094,);
nand I_32577 (I556525,I556486,I556395);
nand I_32578 (I556103,I556378,I556525);
not I_32579 (I556556,I556486);
nor I_32580 (I556573,I556556,I556296);
DFFARX1 I_32581 (I556573,I2683,I556126,I556115,);
nor I_32582 (I556604,I652836,I652827);
or I_32583 (I556106,I556353,I556604);
nor I_32584 (I556097,I556486,I556604);
or I_32585 (I556100,I556220,I556604);
DFFARX1 I_32586 (I556604,I2683,I556126,I556118,);
not I_32587 (I556704,I2690);
DFFARX1 I_32588 (I184270,I2683,I556704,I556730,);
not I_32589 (I556738,I556730);
nand I_32590 (I556755,I184273,I184294);
and I_32591 (I556772,I556755,I184282);
DFFARX1 I_32592 (I556772,I2683,I556704,I556798,);
not I_32593 (I556806,I184279);
DFFARX1 I_32594 (I184270,I2683,I556704,I556832,);
not I_32595 (I556840,I556832);
nor I_32596 (I556857,I556840,I556738);
and I_32597 (I556874,I556857,I184279);
nor I_32598 (I556891,I556840,I556806);
nor I_32599 (I556687,I556798,I556891);
DFFARX1 I_32600 (I184288,I2683,I556704,I556931,);
nor I_32601 (I556939,I556931,I556798);
not I_32602 (I556956,I556939);
not I_32603 (I556973,I556931);
nor I_32604 (I556990,I556973,I556874);
DFFARX1 I_32605 (I556990,I2683,I556704,I556690,);
nand I_32606 (I557021,I184273,I184276);
and I_32607 (I557038,I557021,I184285);
DFFARX1 I_32608 (I557038,I2683,I556704,I557064,);
nor I_32609 (I557072,I557064,I556931);
DFFARX1 I_32610 (I557072,I2683,I556704,I556672,);
nand I_32611 (I557103,I557064,I556973);
nand I_32612 (I556681,I556956,I557103);
not I_32613 (I557134,I557064);
nor I_32614 (I557151,I557134,I556874);
DFFARX1 I_32615 (I557151,I2683,I556704,I556693,);
nor I_32616 (I557182,I184291,I184276);
or I_32617 (I556684,I556931,I557182);
nor I_32618 (I556675,I557064,I557182);
or I_32619 (I556678,I556798,I557182);
DFFARX1 I_32620 (I557182,I2683,I556704,I556696,);
not I_32621 (I557282,I2690);
DFFARX1 I_32622 (I389435,I2683,I557282,I557308,);
not I_32623 (I557316,I557308);
nand I_32624 (I557333,I389426,I389444);
and I_32625 (I557350,I557333,I389447);
DFFARX1 I_32626 (I557350,I2683,I557282,I557376,);
not I_32627 (I557384,I389441);
DFFARX1 I_32628 (I389429,I2683,I557282,I557410,);
not I_32629 (I557418,I557410);
nor I_32630 (I557435,I557418,I557316);
and I_32631 (I557452,I557435,I389441);
nor I_32632 (I557469,I557418,I557384);
nor I_32633 (I557265,I557376,I557469);
DFFARX1 I_32634 (I389438,I2683,I557282,I557509,);
nor I_32635 (I557517,I557509,I557376);
not I_32636 (I557534,I557517);
not I_32637 (I557551,I557509);
nor I_32638 (I557568,I557551,I557452);
DFFARX1 I_32639 (I557568,I2683,I557282,I557268,);
nand I_32640 (I557599,I389453,I389450);
and I_32641 (I557616,I557599,I389432);
DFFARX1 I_32642 (I557616,I2683,I557282,I557642,);
nor I_32643 (I557650,I557642,I557509);
DFFARX1 I_32644 (I557650,I2683,I557282,I557250,);
nand I_32645 (I557681,I557642,I557551);
nand I_32646 (I557259,I557534,I557681);
not I_32647 (I557712,I557642);
nor I_32648 (I557729,I557712,I557452);
DFFARX1 I_32649 (I557729,I2683,I557282,I557271,);
nor I_32650 (I557760,I389426,I389450);
or I_32651 (I557262,I557509,I557760);
nor I_32652 (I557253,I557642,I557760);
or I_32653 (I557256,I557376,I557760);
DFFARX1 I_32654 (I557760,I2683,I557282,I557274,);
not I_32655 (I557860,I2690);
DFFARX1 I_32656 (I972798,I2683,I557860,I557886,);
not I_32657 (I557894,I557886);
nand I_32658 (I557911,I972801,I972810);
and I_32659 (I557928,I557911,I972813);
DFFARX1 I_32660 (I557928,I2683,I557860,I557954,);
not I_32661 (I557962,I972822);
DFFARX1 I_32662 (I972804,I2683,I557860,I557988,);
not I_32663 (I557996,I557988);
nor I_32664 (I558013,I557996,I557894);
and I_32665 (I558030,I558013,I972822);
nor I_32666 (I558047,I557996,I557962);
nor I_32667 (I557843,I557954,I558047);
DFFARX1 I_32668 (I972801,I2683,I557860,I558087,);
nor I_32669 (I558095,I558087,I557954);
not I_32670 (I558112,I558095);
not I_32671 (I558129,I558087);
nor I_32672 (I558146,I558129,I558030);
DFFARX1 I_32673 (I558146,I2683,I557860,I557846,);
nand I_32674 (I558177,I972819,I972798);
and I_32675 (I558194,I558177,I972816);
DFFARX1 I_32676 (I558194,I2683,I557860,I558220,);
nor I_32677 (I558228,I558220,I558087);
DFFARX1 I_32678 (I558228,I2683,I557860,I557828,);
nand I_32679 (I558259,I558220,I558129);
nand I_32680 (I557837,I558112,I558259);
not I_32681 (I558290,I558220);
nor I_32682 (I558307,I558290,I558030);
DFFARX1 I_32683 (I558307,I2683,I557860,I557849,);
nor I_32684 (I558338,I972807,I972798);
or I_32685 (I557840,I558087,I558338);
nor I_32686 (I557831,I558220,I558338);
or I_32687 (I557834,I557954,I558338);
DFFARX1 I_32688 (I558338,I2683,I557860,I557852,);
not I_32689 (I558438,I2690);
DFFARX1 I_32690 (I311794,I2683,I558438,I558464,);
not I_32691 (I558472,I558464);
nand I_32692 (I558489,I311797,I311773);
and I_32693 (I558506,I558489,I311770);
DFFARX1 I_32694 (I558506,I2683,I558438,I558532,);
not I_32695 (I558540,I311776);
DFFARX1 I_32696 (I311770,I2683,I558438,I558566,);
not I_32697 (I558574,I558566);
nor I_32698 (I558591,I558574,I558472);
and I_32699 (I558608,I558591,I311776);
nor I_32700 (I558625,I558574,I558540);
nor I_32701 (I558421,I558532,I558625);
DFFARX1 I_32702 (I311779,I2683,I558438,I558665,);
nor I_32703 (I558673,I558665,I558532);
not I_32704 (I558690,I558673);
not I_32705 (I558707,I558665);
nor I_32706 (I558724,I558707,I558608);
DFFARX1 I_32707 (I558724,I2683,I558438,I558424,);
nand I_32708 (I558755,I311782,I311791);
and I_32709 (I558772,I558755,I311788);
DFFARX1 I_32710 (I558772,I2683,I558438,I558798,);
nor I_32711 (I558806,I558798,I558665);
DFFARX1 I_32712 (I558806,I2683,I558438,I558406,);
nand I_32713 (I558837,I558798,I558707);
nand I_32714 (I558415,I558690,I558837);
not I_32715 (I558868,I558798);
nor I_32716 (I558885,I558868,I558608);
DFFARX1 I_32717 (I558885,I2683,I558438,I558427,);
nor I_32718 (I558916,I311785,I311791);
or I_32719 (I558418,I558665,I558916);
nor I_32720 (I558409,I558798,I558916);
or I_32721 (I558412,I558532,I558916);
DFFARX1 I_32722 (I558916,I2683,I558438,I558430,);
not I_32723 (I559016,I2690);
DFFARX1 I_32724 (I773633,I2683,I559016,I559042,);
not I_32725 (I559050,I559042);
nand I_32726 (I559067,I773609,I773624);
and I_32727 (I559084,I559067,I773636);
DFFARX1 I_32728 (I559084,I2683,I559016,I559110,);
not I_32729 (I559118,I773621);
DFFARX1 I_32730 (I773612,I2683,I559016,I559144,);
not I_32731 (I559152,I559144);
nor I_32732 (I559169,I559152,I559050);
and I_32733 (I559186,I559169,I773621);
nor I_32734 (I559203,I559152,I559118);
nor I_32735 (I558999,I559110,I559203);
DFFARX1 I_32736 (I773609,I2683,I559016,I559243,);
nor I_32737 (I559251,I559243,I559110);
not I_32738 (I559268,I559251);
not I_32739 (I559285,I559243);
nor I_32740 (I559302,I559285,I559186);
DFFARX1 I_32741 (I559302,I2683,I559016,I559002,);
nand I_32742 (I559333,I773627,I773618);
and I_32743 (I559350,I559333,I773630);
DFFARX1 I_32744 (I559350,I2683,I559016,I559376,);
nor I_32745 (I559384,I559376,I559243);
DFFARX1 I_32746 (I559384,I2683,I559016,I558984,);
nand I_32747 (I559415,I559376,I559285);
nand I_32748 (I558993,I559268,I559415);
not I_32749 (I559446,I559376);
nor I_32750 (I559463,I559446,I559186);
DFFARX1 I_32751 (I559463,I2683,I559016,I559005,);
nor I_32752 (I559494,I773615,I773618);
or I_32753 (I558996,I559243,I559494);
nor I_32754 (I558987,I559376,I559494);
or I_32755 (I558990,I559110,I559494);
DFFARX1 I_32756 (I559494,I2683,I559016,I559008,);
not I_32757 (I559594,I2690);
DFFARX1 I_32758 (I255932,I2683,I559594,I559620,);
not I_32759 (I559628,I559620);
nand I_32760 (I559645,I255935,I255911);
and I_32761 (I559662,I559645,I255908);
DFFARX1 I_32762 (I559662,I2683,I559594,I559688,);
not I_32763 (I559696,I255914);
DFFARX1 I_32764 (I255908,I2683,I559594,I559722,);
not I_32765 (I559730,I559722);
nor I_32766 (I559747,I559730,I559628);
and I_32767 (I559764,I559747,I255914);
nor I_32768 (I559781,I559730,I559696);
nor I_32769 (I559577,I559688,I559781);
DFFARX1 I_32770 (I255917,I2683,I559594,I559821,);
nor I_32771 (I559829,I559821,I559688);
not I_32772 (I559846,I559829);
not I_32773 (I559863,I559821);
nor I_32774 (I559880,I559863,I559764);
DFFARX1 I_32775 (I559880,I2683,I559594,I559580,);
nand I_32776 (I559911,I255920,I255929);
and I_32777 (I559928,I559911,I255926);
DFFARX1 I_32778 (I559928,I2683,I559594,I559954,);
nor I_32779 (I559962,I559954,I559821);
DFFARX1 I_32780 (I559962,I2683,I559594,I559562,);
nand I_32781 (I559993,I559954,I559863);
nand I_32782 (I559571,I559846,I559993);
not I_32783 (I560024,I559954);
nor I_32784 (I560041,I560024,I559764);
DFFARX1 I_32785 (I560041,I2683,I559594,I559583,);
nor I_32786 (I560072,I255923,I255929);
or I_32787 (I559574,I559821,I560072);
nor I_32788 (I559565,I559954,I560072);
or I_32789 (I559568,I559688,I560072);
DFFARX1 I_32790 (I560072,I2683,I559594,I559586,);
not I_32791 (I560172,I2690);
DFFARX1 I_32792 (I182485,I2683,I560172,I560198,);
not I_32793 (I560206,I560198);
nand I_32794 (I560223,I182488,I182509);
and I_32795 (I560240,I560223,I182497);
DFFARX1 I_32796 (I560240,I2683,I560172,I560266,);
not I_32797 (I560274,I182494);
DFFARX1 I_32798 (I182485,I2683,I560172,I560300,);
not I_32799 (I560308,I560300);
nor I_32800 (I560325,I560308,I560206);
and I_32801 (I560342,I560325,I182494);
nor I_32802 (I560359,I560308,I560274);
nor I_32803 (I560155,I560266,I560359);
DFFARX1 I_32804 (I182503,I2683,I560172,I560399,);
nor I_32805 (I560407,I560399,I560266);
not I_32806 (I560424,I560407);
not I_32807 (I560441,I560399);
nor I_32808 (I560458,I560441,I560342);
DFFARX1 I_32809 (I560458,I2683,I560172,I560158,);
nand I_32810 (I560489,I182488,I182491);
and I_32811 (I560506,I560489,I182500);
DFFARX1 I_32812 (I560506,I2683,I560172,I560532,);
nor I_32813 (I560540,I560532,I560399);
DFFARX1 I_32814 (I560540,I2683,I560172,I560140,);
nand I_32815 (I560571,I560532,I560441);
nand I_32816 (I560149,I560424,I560571);
not I_32817 (I560602,I560532);
nor I_32818 (I560619,I560602,I560342);
DFFARX1 I_32819 (I560619,I2683,I560172,I560161,);
nor I_32820 (I560650,I182506,I182491);
or I_32821 (I560152,I560399,I560650);
nor I_32822 (I560143,I560532,I560650);
or I_32823 (I560146,I560266,I560650);
DFFARX1 I_32824 (I560650,I2683,I560172,I560164,);
not I_32825 (I560750,I2690);
DFFARX1 I_32826 (I688675,I2683,I560750,I560776,);
not I_32827 (I560784,I560776);
nand I_32828 (I560801,I688663,I688681);
and I_32829 (I560818,I560801,I688678);
DFFARX1 I_32830 (I560818,I2683,I560750,I560844,);
not I_32831 (I560852,I688669);
DFFARX1 I_32832 (I688666,I2683,I560750,I560878,);
not I_32833 (I560886,I560878);
nor I_32834 (I560903,I560886,I560784);
and I_32835 (I560920,I560903,I688669);
nor I_32836 (I560937,I560886,I560852);
nor I_32837 (I560733,I560844,I560937);
DFFARX1 I_32838 (I688660,I2683,I560750,I560977,);
nor I_32839 (I560985,I560977,I560844);
not I_32840 (I561002,I560985);
not I_32841 (I561019,I560977);
nor I_32842 (I561036,I561019,I560920);
DFFARX1 I_32843 (I561036,I2683,I560750,I560736,);
nand I_32844 (I561067,I688660,I688663);
and I_32845 (I561084,I561067,I688666);
DFFARX1 I_32846 (I561084,I2683,I560750,I561110,);
nor I_32847 (I561118,I561110,I560977);
DFFARX1 I_32848 (I561118,I2683,I560750,I560718,);
nand I_32849 (I561149,I561110,I561019);
nand I_32850 (I560727,I561002,I561149);
not I_32851 (I561180,I561110);
nor I_32852 (I561197,I561180,I560920);
DFFARX1 I_32853 (I561197,I2683,I560750,I560739,);
nor I_32854 (I561228,I688672,I688663);
or I_32855 (I560730,I560977,I561228);
nor I_32856 (I560721,I561110,I561228);
or I_32857 (I560724,I560844,I561228);
DFFARX1 I_32858 (I561228,I2683,I560750,I560742,);
not I_32859 (I561328,I2690);
DFFARX1 I_32860 (I120617,I2683,I561328,I561354,);
not I_32861 (I561362,I561354);
nand I_32862 (I561379,I120632,I120605);
and I_32863 (I561396,I561379,I120620);
DFFARX1 I_32864 (I561396,I2683,I561328,I561422,);
not I_32865 (I561430,I120623);
DFFARX1 I_32866 (I120608,I2683,I561328,I561456,);
not I_32867 (I561464,I561456);
nor I_32868 (I561481,I561464,I561362);
and I_32869 (I561498,I561481,I120623);
nor I_32870 (I561515,I561464,I561430);
nor I_32871 (I561311,I561422,I561515);
DFFARX1 I_32872 (I120614,I2683,I561328,I561555,);
nor I_32873 (I561563,I561555,I561422);
not I_32874 (I561580,I561563);
not I_32875 (I561597,I561555);
nor I_32876 (I561614,I561597,I561498);
DFFARX1 I_32877 (I561614,I2683,I561328,I561314,);
nand I_32878 (I561645,I120629,I120611);
and I_32879 (I561662,I561645,I120626);
DFFARX1 I_32880 (I561662,I2683,I561328,I561688,);
nor I_32881 (I561696,I561688,I561555);
DFFARX1 I_32882 (I561696,I2683,I561328,I561296,);
nand I_32883 (I561727,I561688,I561597);
nand I_32884 (I561305,I561580,I561727);
not I_32885 (I561758,I561688);
nor I_32886 (I561775,I561758,I561498);
DFFARX1 I_32887 (I561775,I2683,I561328,I561317,);
nor I_32888 (I561806,I120605,I120611);
or I_32889 (I561308,I561555,I561806);
nor I_32890 (I561299,I561688,I561806);
or I_32891 (I561302,I561422,I561806);
DFFARX1 I_32892 (I561806,I2683,I561328,I561320,);
not I_32893 (I561906,I2690);
DFFARX1 I_32894 (I55362,I2683,I561906,I561932,);
not I_32895 (I561940,I561932);
nand I_32896 (I561957,I55371,I55380);
and I_32897 (I561974,I561957,I55359);
DFFARX1 I_32898 (I561974,I2683,I561906,I562000,);
not I_32899 (I562008,I55362);
DFFARX1 I_32900 (I55377,I2683,I561906,I562034,);
not I_32901 (I562042,I562034);
nor I_32902 (I562059,I562042,I561940);
and I_32903 (I562076,I562059,I55362);
nor I_32904 (I562093,I562042,I562008);
nor I_32905 (I561889,I562000,I562093);
DFFARX1 I_32906 (I55368,I2683,I561906,I562133,);
nor I_32907 (I562141,I562133,I562000);
not I_32908 (I562158,I562141);
not I_32909 (I562175,I562133);
nor I_32910 (I562192,I562175,I562076);
DFFARX1 I_32911 (I562192,I2683,I561906,I561892,);
nand I_32912 (I562223,I55383,I55359);
and I_32913 (I562240,I562223,I55365);
DFFARX1 I_32914 (I562240,I2683,I561906,I562266,);
nor I_32915 (I562274,I562266,I562133);
DFFARX1 I_32916 (I562274,I2683,I561906,I561874,);
nand I_32917 (I562305,I562266,I562175);
nand I_32918 (I561883,I562158,I562305);
not I_32919 (I562336,I562266);
nor I_32920 (I562353,I562336,I562076);
DFFARX1 I_32921 (I562353,I2683,I561906,I561895,);
nor I_32922 (I562384,I55374,I55359);
or I_32923 (I561886,I562133,I562384);
nor I_32924 (I561877,I562266,I562384);
or I_32925 (I561880,I562000,I562384);
DFFARX1 I_32926 (I562384,I2683,I561906,I561898,);
not I_32927 (I562484,I2690);
DFFARX1 I_32928 (I125365,I2683,I562484,I562510,);
not I_32929 (I562518,I562510);
nand I_32930 (I562535,I125368,I125389);
and I_32931 (I562552,I562535,I125377);
DFFARX1 I_32932 (I562552,I2683,I562484,I562578,);
not I_32933 (I562586,I125374);
DFFARX1 I_32934 (I125365,I2683,I562484,I562612,);
not I_32935 (I562620,I562612);
nor I_32936 (I562637,I562620,I562518);
and I_32937 (I562654,I562637,I125374);
nor I_32938 (I562671,I562620,I562586);
nor I_32939 (I562467,I562578,I562671);
DFFARX1 I_32940 (I125383,I2683,I562484,I562711,);
nor I_32941 (I562719,I562711,I562578);
not I_32942 (I562736,I562719);
not I_32943 (I562753,I562711);
nor I_32944 (I562770,I562753,I562654);
DFFARX1 I_32945 (I562770,I2683,I562484,I562470,);
nand I_32946 (I562801,I125368,I125371);
and I_32947 (I562818,I562801,I125380);
DFFARX1 I_32948 (I562818,I2683,I562484,I562844,);
nor I_32949 (I562852,I562844,I562711);
DFFARX1 I_32950 (I562852,I2683,I562484,I562452,);
nand I_32951 (I562883,I562844,I562753);
nand I_32952 (I562461,I562736,I562883);
not I_32953 (I562914,I562844);
nor I_32954 (I562931,I562914,I562654);
DFFARX1 I_32955 (I562931,I2683,I562484,I562473,);
nor I_32956 (I562962,I125386,I125371);
or I_32957 (I562464,I562711,I562962);
nor I_32958 (I562455,I562844,I562962);
or I_32959 (I562458,I562578,I562962);
DFFARX1 I_32960 (I562962,I2683,I562484,I562476,);
not I_32961 (I563062,I2690);
DFFARX1 I_32962 (I896996,I2683,I563062,I563088,);
not I_32963 (I563096,I563088);
nand I_32964 (I563113,I896978,I896990);
and I_32965 (I563130,I563113,I896993);
DFFARX1 I_32966 (I563130,I2683,I563062,I563156,);
not I_32967 (I563164,I896987);
DFFARX1 I_32968 (I896984,I2683,I563062,I563190,);
not I_32969 (I563198,I563190);
nor I_32970 (I563215,I563198,I563096);
and I_32971 (I563232,I563215,I896987);
nor I_32972 (I563249,I563198,I563164);
nor I_32973 (I563045,I563156,I563249);
DFFARX1 I_32974 (I897002,I2683,I563062,I563289,);
nor I_32975 (I563297,I563289,I563156);
not I_32976 (I563314,I563297);
not I_32977 (I563331,I563289);
nor I_32978 (I563348,I563331,I563232);
DFFARX1 I_32979 (I563348,I2683,I563062,I563048,);
nand I_32980 (I563379,I896981,I896981);
and I_32981 (I563396,I563379,I896978);
DFFARX1 I_32982 (I563396,I2683,I563062,I563422,);
nor I_32983 (I563430,I563422,I563289);
DFFARX1 I_32984 (I563430,I2683,I563062,I563030,);
nand I_32985 (I563461,I563422,I563331);
nand I_32986 (I563039,I563314,I563461);
not I_32987 (I563492,I563422);
nor I_32988 (I563509,I563492,I563232);
DFFARX1 I_32989 (I563509,I2683,I563062,I563051,);
nor I_32990 (I563540,I896999,I896981);
or I_32991 (I563042,I563289,I563540);
nor I_32992 (I563033,I563422,I563540);
or I_32993 (I563036,I563156,I563540);
DFFARX1 I_32994 (I563540,I2683,I563062,I563054,);
not I_32995 (I563640,I2690);
DFFARX1 I_32996 (I1017474,I2683,I563640,I563666,);
not I_32997 (I563674,I563666);
nand I_32998 (I563691,I1017498,I1017480);
and I_32999 (I563708,I563691,I1017486);
DFFARX1 I_33000 (I563708,I2683,I563640,I563734,);
not I_33001 (I563742,I1017492);
DFFARX1 I_33002 (I1017477,I2683,I563640,I563768,);
not I_33003 (I563776,I563768);
nor I_33004 (I563793,I563776,I563674);
and I_33005 (I563810,I563793,I1017492);
nor I_33006 (I563827,I563776,I563742);
nor I_33007 (I563623,I563734,I563827);
DFFARX1 I_33008 (I1017489,I2683,I563640,I563867,);
nor I_33009 (I563875,I563867,I563734);
not I_33010 (I563892,I563875);
not I_33011 (I563909,I563867);
nor I_33012 (I563926,I563909,I563810);
DFFARX1 I_33013 (I563926,I2683,I563640,I563626,);
nand I_33014 (I563957,I1017495,I1017483);
and I_33015 (I563974,I563957,I1017477);
DFFARX1 I_33016 (I563974,I2683,I563640,I564000,);
nor I_33017 (I564008,I564000,I563867);
DFFARX1 I_33018 (I564008,I2683,I563640,I563608,);
nand I_33019 (I564039,I564000,I563909);
nand I_33020 (I563617,I563892,I564039);
not I_33021 (I564070,I564000);
nor I_33022 (I564087,I564070,I563810);
DFFARX1 I_33023 (I564087,I2683,I563640,I563629,);
nor I_33024 (I564118,I1017474,I1017483);
or I_33025 (I563620,I563867,I564118);
nor I_33026 (I563611,I564000,I564118);
or I_33027 (I563614,I563734,I564118);
DFFARX1 I_33028 (I564118,I2683,I563640,I563632,);
not I_33029 (I564218,I2690);
DFFARX1 I_33030 (I819787,I2683,I564218,I564244,);
not I_33031 (I564252,I564244);
nand I_33032 (I564269,I819784,I819802);
and I_33033 (I564286,I564269,I819799);
DFFARX1 I_33034 (I564286,I2683,I564218,I564312,);
not I_33035 (I564320,I819781);
DFFARX1 I_33036 (I819784,I2683,I564218,I564346,);
not I_33037 (I564354,I564346);
nor I_33038 (I564371,I564354,I564252);
and I_33039 (I564388,I564371,I819781);
nor I_33040 (I564405,I564354,I564320);
nor I_33041 (I564201,I564312,I564405);
DFFARX1 I_33042 (I819793,I2683,I564218,I564445,);
nor I_33043 (I564453,I564445,I564312);
not I_33044 (I564470,I564453);
not I_33045 (I564487,I564445);
nor I_33046 (I564504,I564487,I564388);
DFFARX1 I_33047 (I564504,I2683,I564218,I564204,);
nand I_33048 (I564535,I819796,I819781);
and I_33049 (I564552,I564535,I819787);
DFFARX1 I_33050 (I564552,I2683,I564218,I564578,);
nor I_33051 (I564586,I564578,I564445);
DFFARX1 I_33052 (I564586,I2683,I564218,I564186,);
nand I_33053 (I564617,I564578,I564487);
nand I_33054 (I564195,I564470,I564617);
not I_33055 (I564648,I564578);
nor I_33056 (I564665,I564648,I564388);
DFFARX1 I_33057 (I564665,I2683,I564218,I564207,);
nor I_33058 (I564696,I819790,I819781);
or I_33059 (I564198,I564445,I564696);
nor I_33060 (I564189,I564578,I564696);
or I_33061 (I564192,I564312,I564696);
DFFARX1 I_33062 (I564696,I2683,I564218,I564210,);
not I_33063 (I564796,I2690);
DFFARX1 I_33064 (I95941,I2683,I564796,I564822,);
not I_33065 (I564830,I564822);
nand I_33066 (I564847,I95950,I95959);
and I_33067 (I564864,I564847,I95938);
DFFARX1 I_33068 (I564864,I2683,I564796,I564890,);
not I_33069 (I564898,I95941);
DFFARX1 I_33070 (I95956,I2683,I564796,I564924,);
not I_33071 (I564932,I564924);
nor I_33072 (I564949,I564932,I564830);
and I_33073 (I564966,I564949,I95941);
nor I_33074 (I564983,I564932,I564898);
nor I_33075 (I564779,I564890,I564983);
DFFARX1 I_33076 (I95947,I2683,I564796,I565023,);
nor I_33077 (I565031,I565023,I564890);
not I_33078 (I565048,I565031);
not I_33079 (I565065,I565023);
nor I_33080 (I565082,I565065,I564966);
DFFARX1 I_33081 (I565082,I2683,I564796,I564782,);
nand I_33082 (I565113,I95962,I95938);
and I_33083 (I565130,I565113,I95944);
DFFARX1 I_33084 (I565130,I2683,I564796,I565156,);
nor I_33085 (I565164,I565156,I565023);
DFFARX1 I_33086 (I565164,I2683,I564796,I564764,);
nand I_33087 (I565195,I565156,I565065);
nand I_33088 (I564773,I565048,I565195);
not I_33089 (I565226,I565156);
nor I_33090 (I565243,I565226,I564966);
DFFARX1 I_33091 (I565243,I2683,I564796,I564785,);
nor I_33092 (I565274,I95953,I95938);
or I_33093 (I564776,I565023,I565274);
nor I_33094 (I564767,I565156,I565274);
or I_33095 (I564770,I564890,I565274);
DFFARX1 I_33096 (I565274,I2683,I564796,I564788,);
not I_33097 (I565374,I2690);
DFFARX1 I_33098 (I306524,I2683,I565374,I565400,);
not I_33099 (I565408,I565400);
nand I_33100 (I565425,I306527,I306503);
and I_33101 (I565442,I565425,I306500);
DFFARX1 I_33102 (I565442,I2683,I565374,I565468,);
not I_33103 (I565476,I306506);
DFFARX1 I_33104 (I306500,I2683,I565374,I565502,);
not I_33105 (I565510,I565502);
nor I_33106 (I565527,I565510,I565408);
and I_33107 (I565544,I565527,I306506);
nor I_33108 (I565561,I565510,I565476);
nor I_33109 (I565357,I565468,I565561);
DFFARX1 I_33110 (I306509,I2683,I565374,I565601,);
nor I_33111 (I565609,I565601,I565468);
not I_33112 (I565626,I565609);
not I_33113 (I565643,I565601);
nor I_33114 (I565660,I565643,I565544);
DFFARX1 I_33115 (I565660,I2683,I565374,I565360,);
nand I_33116 (I565691,I306512,I306521);
and I_33117 (I565708,I565691,I306518);
DFFARX1 I_33118 (I565708,I2683,I565374,I565734,);
nor I_33119 (I565742,I565734,I565601);
DFFARX1 I_33120 (I565742,I2683,I565374,I565342,);
nand I_33121 (I565773,I565734,I565643);
nand I_33122 (I565351,I565626,I565773);
not I_33123 (I565804,I565734);
nor I_33124 (I565821,I565804,I565544);
DFFARX1 I_33125 (I565821,I2683,I565374,I565363,);
nor I_33126 (I565852,I306515,I306521);
or I_33127 (I565354,I565601,I565852);
nor I_33128 (I565345,I565734,I565852);
or I_33129 (I565348,I565468,I565852);
DFFARX1 I_33130 (I565852,I2683,I565374,I565366,);
not I_33131 (I565952,I2690);
DFFARX1 I_33132 (I666541,I2683,I565952,I565978,);
not I_33133 (I565986,I565978);
nand I_33134 (I566003,I666529,I666547);
and I_33135 (I566020,I566003,I666544);
DFFARX1 I_33136 (I566020,I2683,I565952,I566046,);
not I_33137 (I566054,I666535);
DFFARX1 I_33138 (I666532,I2683,I565952,I566080,);
not I_33139 (I566088,I566080);
nor I_33140 (I566105,I566088,I565986);
and I_33141 (I566122,I566105,I666535);
nor I_33142 (I566139,I566088,I566054);
nor I_33143 (I565935,I566046,I566139);
DFFARX1 I_33144 (I666526,I2683,I565952,I566179,);
nor I_33145 (I566187,I566179,I566046);
not I_33146 (I566204,I566187);
not I_33147 (I566221,I566179);
nor I_33148 (I566238,I566221,I566122);
DFFARX1 I_33149 (I566238,I2683,I565952,I565938,);
nand I_33150 (I566269,I666526,I666529);
and I_33151 (I566286,I566269,I666532);
DFFARX1 I_33152 (I566286,I2683,I565952,I566312,);
nor I_33153 (I566320,I566312,I566179);
DFFARX1 I_33154 (I566320,I2683,I565952,I565920,);
nand I_33155 (I566351,I566312,I566221);
nand I_33156 (I565929,I566204,I566351);
not I_33157 (I566382,I566312);
nor I_33158 (I566399,I566382,I566122);
DFFARX1 I_33159 (I566399,I2683,I565952,I565941,);
nor I_33160 (I566430,I666538,I666529);
or I_33161 (I565932,I566179,I566430);
nor I_33162 (I565923,I566312,I566430);
or I_33163 (I565926,I566046,I566430);
DFFARX1 I_33164 (I566430,I2683,I565952,I565944,);
not I_33165 (I566530,I2690);
DFFARX1 I_33166 (I470550,I2683,I566530,I566556,);
not I_33167 (I566564,I566556);
nand I_33168 (I566581,I470559,I470568);
and I_33169 (I566598,I566581,I470574);
DFFARX1 I_33170 (I566598,I2683,I566530,I566624,);
not I_33171 (I566632,I470571);
DFFARX1 I_33172 (I470556,I2683,I566530,I566658,);
not I_33173 (I566666,I566658);
nor I_33174 (I566683,I566666,I566564);
and I_33175 (I566700,I566683,I470571);
nor I_33176 (I566717,I566666,I566632);
nor I_33177 (I566513,I566624,I566717);
DFFARX1 I_33178 (I470565,I2683,I566530,I566757,);
nor I_33179 (I566765,I566757,I566624);
not I_33180 (I566782,I566765);
not I_33181 (I566799,I566757);
nor I_33182 (I566816,I566799,I566700);
DFFARX1 I_33183 (I566816,I2683,I566530,I566516,);
nand I_33184 (I566847,I470562,I470553);
and I_33185 (I566864,I566847,I470550);
DFFARX1 I_33186 (I566864,I2683,I566530,I566890,);
nor I_33187 (I566898,I566890,I566757);
DFFARX1 I_33188 (I566898,I2683,I566530,I566498,);
nand I_33189 (I566929,I566890,I566799);
nand I_33190 (I566507,I566782,I566929);
not I_33191 (I566960,I566890);
nor I_33192 (I566977,I566960,I566700);
DFFARX1 I_33193 (I566977,I2683,I566530,I566519,);
nor I_33194 (I567008,I470553,I470553);
or I_33195 (I566510,I566757,I567008);
nor I_33196 (I566501,I566890,I567008);
or I_33197 (I566504,I566624,I567008);
DFFARX1 I_33198 (I567008,I2683,I566530,I566522,);
not I_33199 (I567108,I2690);
DFFARX1 I_33200 (I41142,I2683,I567108,I567134,);
not I_33201 (I567142,I567134);
nand I_33202 (I567159,I41139,I41130);
and I_33203 (I567176,I567159,I41130);
DFFARX1 I_33204 (I567176,I2683,I567108,I567202,);
not I_33205 (I567210,I41133);
DFFARX1 I_33206 (I41148,I2683,I567108,I567236,);
not I_33207 (I567244,I567236);
nor I_33208 (I567261,I567244,I567142);
and I_33209 (I567278,I567261,I41133);
nor I_33210 (I567295,I567244,I567210);
nor I_33211 (I567091,I567202,I567295);
DFFARX1 I_33212 (I41133,I2683,I567108,I567335,);
nor I_33213 (I567343,I567335,I567202);
not I_33214 (I567360,I567343);
not I_33215 (I567377,I567335);
nor I_33216 (I567394,I567377,I567278);
DFFARX1 I_33217 (I567394,I2683,I567108,I567094,);
nand I_33218 (I567425,I41151,I41136);
and I_33219 (I567442,I567425,I41154);
DFFARX1 I_33220 (I567442,I2683,I567108,I567468,);
nor I_33221 (I567476,I567468,I567335);
DFFARX1 I_33222 (I567476,I2683,I567108,I567076,);
nand I_33223 (I567507,I567468,I567377);
nand I_33224 (I567085,I567360,I567507);
not I_33225 (I567538,I567468);
nor I_33226 (I567555,I567538,I567278);
DFFARX1 I_33227 (I567555,I2683,I567108,I567097,);
nor I_33228 (I567586,I41145,I41136);
or I_33229 (I567088,I567335,I567586);
nor I_33230 (I567079,I567468,I567586);
or I_33231 (I567082,I567202,I567586);
DFFARX1 I_33232 (I567586,I2683,I567108,I567100,);
not I_33233 (I567686,I2690);
DFFARX1 I_33234 (I989730,I2683,I567686,I567712,);
not I_33235 (I567720,I567712);
nand I_33236 (I567737,I989754,I989736);
and I_33237 (I567754,I567737,I989742);
DFFARX1 I_33238 (I567754,I2683,I567686,I567780,);
not I_33239 (I567788,I989748);
DFFARX1 I_33240 (I989733,I2683,I567686,I567814,);
not I_33241 (I567822,I567814);
nor I_33242 (I567839,I567822,I567720);
and I_33243 (I567856,I567839,I989748);
nor I_33244 (I567873,I567822,I567788);
nor I_33245 (I567669,I567780,I567873);
DFFARX1 I_33246 (I989745,I2683,I567686,I567913,);
nor I_33247 (I567921,I567913,I567780);
not I_33248 (I567938,I567921);
not I_33249 (I567955,I567913);
nor I_33250 (I567972,I567955,I567856);
DFFARX1 I_33251 (I567972,I2683,I567686,I567672,);
nand I_33252 (I568003,I989751,I989739);
and I_33253 (I568020,I568003,I989733);
DFFARX1 I_33254 (I568020,I2683,I567686,I568046,);
nor I_33255 (I568054,I568046,I567913);
DFFARX1 I_33256 (I568054,I2683,I567686,I567654,);
nand I_33257 (I568085,I568046,I567955);
nand I_33258 (I567663,I567938,I568085);
not I_33259 (I568116,I568046);
nor I_33260 (I568133,I568116,I567856);
DFFARX1 I_33261 (I568133,I2683,I567686,I567675,);
nor I_33262 (I568164,I989730,I989739);
or I_33263 (I567666,I567913,I568164);
nor I_33264 (I567657,I568046,I568164);
or I_33265 (I567660,I567780,I568164);
DFFARX1 I_33266 (I568164,I2683,I567686,I567678,);
not I_33267 (I568264,I2690);
DFFARX1 I_33268 (I716139,I2683,I568264,I568290,);
not I_33269 (I568298,I568290);
nand I_33270 (I568315,I716115,I716130);
and I_33271 (I568332,I568315,I716142);
DFFARX1 I_33272 (I568332,I2683,I568264,I568358,);
not I_33273 (I568366,I716127);
DFFARX1 I_33274 (I716118,I2683,I568264,I568392,);
not I_33275 (I568400,I568392);
nor I_33276 (I568417,I568400,I568298);
and I_33277 (I568434,I568417,I716127);
nor I_33278 (I568451,I568400,I568366);
nor I_33279 (I568247,I568358,I568451);
DFFARX1 I_33280 (I716115,I2683,I568264,I568491,);
nor I_33281 (I568499,I568491,I568358);
not I_33282 (I568516,I568499);
not I_33283 (I568533,I568491);
nor I_33284 (I568550,I568533,I568434);
DFFARX1 I_33285 (I568550,I2683,I568264,I568250,);
nand I_33286 (I568581,I716133,I716124);
and I_33287 (I568598,I568581,I716136);
DFFARX1 I_33288 (I568598,I2683,I568264,I568624,);
nor I_33289 (I568632,I568624,I568491);
DFFARX1 I_33290 (I568632,I2683,I568264,I568232,);
nand I_33291 (I568663,I568624,I568533);
nand I_33292 (I568241,I568516,I568663);
not I_33293 (I568694,I568624);
nor I_33294 (I568711,I568694,I568434);
DFFARX1 I_33295 (I568711,I2683,I568264,I568253,);
nor I_33296 (I568742,I716121,I716124);
or I_33297 (I568244,I568491,I568742);
nor I_33298 (I568235,I568624,I568742);
or I_33299 (I568238,I568358,I568742);
DFFARX1 I_33300 (I568742,I2683,I568264,I568256,);
not I_33301 (I568842,I2690);
DFFARX1 I_33302 (I43250,I2683,I568842,I568868,);
not I_33303 (I568876,I568868);
nand I_33304 (I568893,I43247,I43238);
and I_33305 (I568910,I568893,I43238);
DFFARX1 I_33306 (I568910,I2683,I568842,I568936,);
not I_33307 (I568944,I43241);
DFFARX1 I_33308 (I43256,I2683,I568842,I568970,);
not I_33309 (I568978,I568970);
nor I_33310 (I568995,I568978,I568876);
and I_33311 (I569012,I568995,I43241);
nor I_33312 (I569029,I568978,I568944);
nor I_33313 (I568825,I568936,I569029);
DFFARX1 I_33314 (I43241,I2683,I568842,I569069,);
nor I_33315 (I569077,I569069,I568936);
not I_33316 (I569094,I569077);
not I_33317 (I569111,I569069);
nor I_33318 (I569128,I569111,I569012);
DFFARX1 I_33319 (I569128,I2683,I568842,I568828,);
nand I_33320 (I569159,I43259,I43244);
and I_33321 (I569176,I569159,I43262);
DFFARX1 I_33322 (I569176,I2683,I568842,I569202,);
nor I_33323 (I569210,I569202,I569069);
DFFARX1 I_33324 (I569210,I2683,I568842,I568810,);
nand I_33325 (I569241,I569202,I569111);
nand I_33326 (I568819,I569094,I569241);
not I_33327 (I569272,I569202);
nor I_33328 (I569289,I569272,I569012);
DFFARX1 I_33329 (I569289,I2683,I568842,I568831,);
nor I_33330 (I569320,I43253,I43244);
or I_33331 (I568822,I569069,I569320);
nor I_33332 (I568813,I569202,I569320);
or I_33333 (I568816,I568936,I569320);
DFFARX1 I_33334 (I569320,I2683,I568842,I568834,);
not I_33335 (I569420,I2690);
DFFARX1 I_33336 (I361147,I2683,I569420,I569446,);
not I_33337 (I569454,I569446);
nand I_33338 (I569471,I361138,I361156);
and I_33339 (I569488,I569471,I361159);
DFFARX1 I_33340 (I569488,I2683,I569420,I569514,);
not I_33341 (I569522,I361153);
DFFARX1 I_33342 (I361141,I2683,I569420,I569548,);
not I_33343 (I569556,I569548);
nor I_33344 (I569573,I569556,I569454);
and I_33345 (I569590,I569573,I361153);
nor I_33346 (I569607,I569556,I569522);
nor I_33347 (I569403,I569514,I569607);
DFFARX1 I_33348 (I361150,I2683,I569420,I569647,);
nor I_33349 (I569655,I569647,I569514);
not I_33350 (I569672,I569655);
not I_33351 (I569689,I569647);
nor I_33352 (I569706,I569689,I569590);
DFFARX1 I_33353 (I569706,I2683,I569420,I569406,);
nand I_33354 (I569737,I361165,I361162);
and I_33355 (I569754,I569737,I361144);
DFFARX1 I_33356 (I569754,I2683,I569420,I569780,);
nor I_33357 (I569788,I569780,I569647);
DFFARX1 I_33358 (I569788,I2683,I569420,I569388,);
nand I_33359 (I569819,I569780,I569689);
nand I_33360 (I569397,I569672,I569819);
not I_33361 (I569850,I569780);
nor I_33362 (I569867,I569850,I569590);
DFFARX1 I_33363 (I569867,I2683,I569420,I569409,);
nor I_33364 (I569898,I361138,I361162);
or I_33365 (I569400,I569647,I569898);
nor I_33366 (I569391,I569780,I569898);
or I_33367 (I569394,I569514,I569898);
DFFARX1 I_33368 (I569898,I2683,I569420,I569412,);
not I_33369 (I569998,I2690);
DFFARX1 I_33370 (I485578,I2683,I569998,I570024,);
not I_33371 (I570032,I570024);
nand I_33372 (I570049,I485587,I485596);
and I_33373 (I570066,I570049,I485602);
DFFARX1 I_33374 (I570066,I2683,I569998,I570092,);
not I_33375 (I570100,I485599);
DFFARX1 I_33376 (I485584,I2683,I569998,I570126,);
not I_33377 (I570134,I570126);
nor I_33378 (I570151,I570134,I570032);
and I_33379 (I570168,I570151,I485599);
nor I_33380 (I570185,I570134,I570100);
nor I_33381 (I569981,I570092,I570185);
DFFARX1 I_33382 (I485593,I2683,I569998,I570225,);
nor I_33383 (I570233,I570225,I570092);
not I_33384 (I570250,I570233);
not I_33385 (I570267,I570225);
nor I_33386 (I570284,I570267,I570168);
DFFARX1 I_33387 (I570284,I2683,I569998,I569984,);
nand I_33388 (I570315,I485590,I485581);
and I_33389 (I570332,I570315,I485578);
DFFARX1 I_33390 (I570332,I2683,I569998,I570358,);
nor I_33391 (I570366,I570358,I570225);
DFFARX1 I_33392 (I570366,I2683,I569998,I569966,);
nand I_33393 (I570397,I570358,I570267);
nand I_33394 (I569975,I570250,I570397);
not I_33395 (I570428,I570358);
nor I_33396 (I570445,I570428,I570168);
DFFARX1 I_33397 (I570445,I2683,I569998,I569987,);
nor I_33398 (I570476,I485581,I485581);
or I_33399 (I569978,I570225,I570476);
nor I_33400 (I569969,I570358,I570476);
or I_33401 (I569972,I570092,I570476);
DFFARX1 I_33402 (I570476,I2683,I569998,I569990,);
not I_33403 (I570576,I2690);
DFFARX1 I_33404 (I431807,I2683,I570576,I570602,);
not I_33405 (I570610,I570602);
nand I_33406 (I570627,I431822,I431807);
and I_33407 (I570644,I570627,I431810);
DFFARX1 I_33408 (I570644,I2683,I570576,I570670,);
not I_33409 (I570678,I431810);
DFFARX1 I_33410 (I431819,I2683,I570576,I570704,);
not I_33411 (I570712,I570704);
nor I_33412 (I570729,I570712,I570610);
and I_33413 (I570746,I570729,I431810);
nor I_33414 (I570763,I570712,I570678);
nor I_33415 (I570559,I570670,I570763);
DFFARX1 I_33416 (I431813,I2683,I570576,I570803,);
nor I_33417 (I570811,I570803,I570670);
not I_33418 (I570828,I570811);
not I_33419 (I570845,I570803);
nor I_33420 (I570862,I570845,I570746);
DFFARX1 I_33421 (I570862,I2683,I570576,I570562,);
nand I_33422 (I570893,I431816,I431825);
and I_33423 (I570910,I570893,I431831);
DFFARX1 I_33424 (I570910,I2683,I570576,I570936,);
nor I_33425 (I570944,I570936,I570803);
DFFARX1 I_33426 (I570944,I2683,I570576,I570544,);
nand I_33427 (I570975,I570936,I570845);
nand I_33428 (I570553,I570828,I570975);
not I_33429 (I571006,I570936);
nor I_33430 (I571023,I571006,I570746);
DFFARX1 I_33431 (I571023,I2683,I570576,I570565,);
nor I_33432 (I571054,I431828,I431825);
or I_33433 (I570556,I570803,I571054);
nor I_33434 (I570547,I570936,I571054);
or I_33435 (I570550,I570670,I571054);
DFFARX1 I_33436 (I571054,I2683,I570576,I570568,);
not I_33437 (I571154,I2690);
DFFARX1 I_33438 (I630705,I2683,I571154,I571180,);
not I_33439 (I571188,I571180);
nand I_33440 (I571205,I630693,I630711);
and I_33441 (I571222,I571205,I630708);
DFFARX1 I_33442 (I571222,I2683,I571154,I571248,);
not I_33443 (I571256,I630699);
DFFARX1 I_33444 (I630696,I2683,I571154,I571282,);
not I_33445 (I571290,I571282);
nor I_33446 (I571307,I571290,I571188);
and I_33447 (I571324,I571307,I630699);
nor I_33448 (I571341,I571290,I571256);
nor I_33449 (I571137,I571248,I571341);
DFFARX1 I_33450 (I630690,I2683,I571154,I571381,);
nor I_33451 (I571389,I571381,I571248);
not I_33452 (I571406,I571389);
not I_33453 (I571423,I571381);
nor I_33454 (I571440,I571423,I571324);
DFFARX1 I_33455 (I571440,I2683,I571154,I571140,);
nand I_33456 (I571471,I630690,I630693);
and I_33457 (I571488,I571471,I630696);
DFFARX1 I_33458 (I571488,I2683,I571154,I571514,);
nor I_33459 (I571522,I571514,I571381);
DFFARX1 I_33460 (I571522,I2683,I571154,I571122,);
nand I_33461 (I571553,I571514,I571423);
nand I_33462 (I571131,I571406,I571553);
not I_33463 (I571584,I571514);
nor I_33464 (I571601,I571584,I571324);
DFFARX1 I_33465 (I571601,I2683,I571154,I571143,);
nor I_33466 (I571632,I630702,I630693);
or I_33467 (I571134,I571381,I571632);
nor I_33468 (I571125,I571514,I571632);
or I_33469 (I571128,I571248,I571632);
DFFARX1 I_33470 (I571632,I2683,I571154,I571146,);
not I_33471 (I571732,I2690);
DFFARX1 I_33472 (I1038836,I2683,I571732,I571758,);
not I_33473 (I571766,I571758);
nand I_33474 (I571783,I1038821,I1038809);
and I_33475 (I571800,I571783,I1038824);
DFFARX1 I_33476 (I571800,I2683,I571732,I571826,);
not I_33477 (I571834,I1038809);
DFFARX1 I_33478 (I1038827,I2683,I571732,I571860,);
not I_33479 (I571868,I571860);
nor I_33480 (I571885,I571868,I571766);
and I_33481 (I571902,I571885,I1038809);
nor I_33482 (I571919,I571868,I571834);
nor I_33483 (I571715,I571826,I571919);
DFFARX1 I_33484 (I1038815,I2683,I571732,I571959,);
nor I_33485 (I571967,I571959,I571826);
not I_33486 (I571984,I571967);
not I_33487 (I572001,I571959);
nor I_33488 (I572018,I572001,I571902);
DFFARX1 I_33489 (I572018,I2683,I571732,I571718,);
nand I_33490 (I572049,I1038812,I1038818);
and I_33491 (I572066,I572049,I1038833);
DFFARX1 I_33492 (I572066,I2683,I571732,I572092,);
nor I_33493 (I572100,I572092,I571959);
DFFARX1 I_33494 (I572100,I2683,I571732,I571700,);
nand I_33495 (I572131,I572092,I572001);
nand I_33496 (I571709,I571984,I572131);
not I_33497 (I572162,I572092);
nor I_33498 (I572179,I572162,I571902);
DFFARX1 I_33499 (I572179,I2683,I571732,I571721,);
nor I_33500 (I572210,I1038830,I1038818);
or I_33501 (I571712,I571959,I572210);
nor I_33502 (I571703,I572092,I572210);
or I_33503 (I571706,I571826,I572210);
DFFARX1 I_33504 (I572210,I2683,I571732,I571724,);
not I_33505 (I572310,I2690);
DFFARX1 I_33506 (I881390,I2683,I572310,I572336,);
not I_33507 (I572344,I572336);
nand I_33508 (I572361,I881372,I881384);
and I_33509 (I572378,I572361,I881387);
DFFARX1 I_33510 (I572378,I2683,I572310,I572404,);
not I_33511 (I572412,I881381);
DFFARX1 I_33512 (I881378,I2683,I572310,I572438,);
not I_33513 (I572446,I572438);
nor I_33514 (I572463,I572446,I572344);
and I_33515 (I572480,I572463,I881381);
nor I_33516 (I572497,I572446,I572412);
nor I_33517 (I572293,I572404,I572497);
DFFARX1 I_33518 (I881396,I2683,I572310,I572537,);
nor I_33519 (I572545,I572537,I572404);
not I_33520 (I572562,I572545);
not I_33521 (I572579,I572537);
nor I_33522 (I572596,I572579,I572480);
DFFARX1 I_33523 (I572596,I2683,I572310,I572296,);
nand I_33524 (I572627,I881375,I881375);
and I_33525 (I572644,I572627,I881372);
DFFARX1 I_33526 (I572644,I2683,I572310,I572670,);
nor I_33527 (I572678,I572670,I572537);
DFFARX1 I_33528 (I572678,I2683,I572310,I572278,);
nand I_33529 (I572709,I572670,I572579);
nand I_33530 (I572287,I572562,I572709);
not I_33531 (I572740,I572670);
nor I_33532 (I572757,I572740,I572480);
DFFARX1 I_33533 (I572757,I2683,I572310,I572299,);
nor I_33534 (I572788,I881393,I881375);
or I_33535 (I572290,I572537,I572788);
nor I_33536 (I572281,I572670,I572788);
or I_33537 (I572284,I572404,I572788);
DFFARX1 I_33538 (I572788,I2683,I572310,I572302,);
not I_33539 (I572888,I2690);
DFFARX1 I_33540 (I187245,I2683,I572888,I572914,);
not I_33541 (I572922,I572914);
nand I_33542 (I572939,I187248,I187269);
and I_33543 (I572956,I572939,I187257);
DFFARX1 I_33544 (I572956,I2683,I572888,I572982,);
not I_33545 (I572990,I187254);
DFFARX1 I_33546 (I187245,I2683,I572888,I573016,);
not I_33547 (I573024,I573016);
nor I_33548 (I573041,I573024,I572922);
and I_33549 (I573058,I573041,I187254);
nor I_33550 (I573075,I573024,I572990);
nor I_33551 (I572871,I572982,I573075);
DFFARX1 I_33552 (I187263,I2683,I572888,I573115,);
nor I_33553 (I573123,I573115,I572982);
not I_33554 (I573140,I573123);
not I_33555 (I573157,I573115);
nor I_33556 (I573174,I573157,I573058);
DFFARX1 I_33557 (I573174,I2683,I572888,I572874,);
nand I_33558 (I573205,I187248,I187251);
and I_33559 (I573222,I573205,I187260);
DFFARX1 I_33560 (I573222,I2683,I572888,I573248,);
nor I_33561 (I573256,I573248,I573115);
DFFARX1 I_33562 (I573256,I2683,I572888,I572856,);
nand I_33563 (I573287,I573248,I573157);
nand I_33564 (I572865,I573140,I573287);
not I_33565 (I573318,I573248);
nor I_33566 (I573335,I573318,I573058);
DFFARX1 I_33567 (I573335,I2683,I572888,I572877,);
nor I_33568 (I573366,I187266,I187251);
or I_33569 (I572868,I573115,I573366);
nor I_33570 (I572859,I573248,I573366);
or I_33571 (I572862,I572982,I573366);
DFFARX1 I_33572 (I573366,I2683,I572888,I572880,);
not I_33573 (I573466,I2690);
DFFARX1 I_33574 (I466504,I2683,I573466,I573492,);
not I_33575 (I573500,I573492);
nand I_33576 (I573517,I466513,I466522);
and I_33577 (I573534,I573517,I466528);
DFFARX1 I_33578 (I573534,I2683,I573466,I573560,);
not I_33579 (I573568,I466525);
DFFARX1 I_33580 (I466510,I2683,I573466,I573594,);
not I_33581 (I573602,I573594);
nor I_33582 (I573619,I573602,I573500);
and I_33583 (I573636,I573619,I466525);
nor I_33584 (I573653,I573602,I573568);
nor I_33585 (I573449,I573560,I573653);
DFFARX1 I_33586 (I466519,I2683,I573466,I573693,);
nor I_33587 (I573701,I573693,I573560);
not I_33588 (I573718,I573701);
not I_33589 (I573735,I573693);
nor I_33590 (I573752,I573735,I573636);
DFFARX1 I_33591 (I573752,I2683,I573466,I573452,);
nand I_33592 (I573783,I466516,I466507);
and I_33593 (I573800,I573783,I466504);
DFFARX1 I_33594 (I573800,I2683,I573466,I573826,);
nor I_33595 (I573834,I573826,I573693);
DFFARX1 I_33596 (I573834,I2683,I573466,I573434,);
nand I_33597 (I573865,I573826,I573735);
nand I_33598 (I573443,I573718,I573865);
not I_33599 (I573896,I573826);
nor I_33600 (I573913,I573896,I573636);
DFFARX1 I_33601 (I573913,I2683,I573466,I573455,);
nor I_33602 (I573944,I466507,I466507);
or I_33603 (I573446,I573693,I573944);
nor I_33604 (I573437,I573826,I573944);
or I_33605 (I573440,I573560,I573944);
DFFARX1 I_33606 (I573944,I2683,I573466,I573458,);
not I_33607 (I574044,I2690);
DFFARX1 I_33608 (I686040,I2683,I574044,I574070,);
not I_33609 (I574078,I574070);
nand I_33610 (I574095,I686028,I686046);
and I_33611 (I574112,I574095,I686043);
DFFARX1 I_33612 (I574112,I2683,I574044,I574138,);
not I_33613 (I574146,I686034);
DFFARX1 I_33614 (I686031,I2683,I574044,I574172,);
not I_33615 (I574180,I574172);
nor I_33616 (I574197,I574180,I574078);
and I_33617 (I574214,I574197,I686034);
nor I_33618 (I574231,I574180,I574146);
nor I_33619 (I574027,I574138,I574231);
DFFARX1 I_33620 (I686025,I2683,I574044,I574271,);
nor I_33621 (I574279,I574271,I574138);
not I_33622 (I574296,I574279);
not I_33623 (I574313,I574271);
nor I_33624 (I574330,I574313,I574214);
DFFARX1 I_33625 (I574330,I2683,I574044,I574030,);
nand I_33626 (I574361,I686025,I686028);
and I_33627 (I574378,I574361,I686031);
DFFARX1 I_33628 (I574378,I2683,I574044,I574404,);
nor I_33629 (I574412,I574404,I574271);
DFFARX1 I_33630 (I574412,I2683,I574044,I574012,);
nand I_33631 (I574443,I574404,I574313);
nand I_33632 (I574021,I574296,I574443);
not I_33633 (I574474,I574404);
nor I_33634 (I574491,I574474,I574214);
DFFARX1 I_33635 (I574491,I2683,I574044,I574033,);
nor I_33636 (I574522,I686037,I686028);
or I_33637 (I574024,I574271,I574522);
nor I_33638 (I574015,I574404,I574522);
or I_33639 (I574018,I574138,I574522);
DFFARX1 I_33640 (I574522,I2683,I574044,I574036,);
not I_33641 (I574622,I2690);
DFFARX1 I_33642 (I716785,I2683,I574622,I574648,);
not I_33643 (I574656,I574648);
nand I_33644 (I574673,I716761,I716776);
and I_33645 (I574690,I574673,I716788);
DFFARX1 I_33646 (I574690,I2683,I574622,I574716,);
not I_33647 (I574724,I716773);
DFFARX1 I_33648 (I716764,I2683,I574622,I574750,);
not I_33649 (I574758,I574750);
nor I_33650 (I574775,I574758,I574656);
and I_33651 (I574792,I574775,I716773);
nor I_33652 (I574809,I574758,I574724);
nor I_33653 (I574605,I574716,I574809);
DFFARX1 I_33654 (I716761,I2683,I574622,I574849,);
nor I_33655 (I574857,I574849,I574716);
not I_33656 (I574874,I574857);
not I_33657 (I574891,I574849);
nor I_33658 (I574908,I574891,I574792);
DFFARX1 I_33659 (I574908,I2683,I574622,I574608,);
nand I_33660 (I574939,I716779,I716770);
and I_33661 (I574956,I574939,I716782);
DFFARX1 I_33662 (I574956,I2683,I574622,I574982,);
nor I_33663 (I574990,I574982,I574849);
DFFARX1 I_33664 (I574990,I2683,I574622,I574590,);
nand I_33665 (I575021,I574982,I574891);
nand I_33666 (I574599,I574874,I575021);
not I_33667 (I575052,I574982);
nor I_33668 (I575069,I575052,I574792);
DFFARX1 I_33669 (I575069,I2683,I574622,I574611,);
nor I_33670 (I575100,I716767,I716770);
or I_33671 (I574602,I574849,I575100);
nor I_33672 (I574593,I574982,I575100);
or I_33673 (I574596,I574716,I575100);
DFFARX1 I_33674 (I575100,I2683,I574622,I574614,);
not I_33675 (I575200,I2690);
DFFARX1 I_33676 (I223785,I2683,I575200,I575226,);
not I_33677 (I575234,I575226);
nand I_33678 (I575251,I223788,I223764);
and I_33679 (I575268,I575251,I223761);
DFFARX1 I_33680 (I575268,I2683,I575200,I575294,);
not I_33681 (I575302,I223767);
DFFARX1 I_33682 (I223761,I2683,I575200,I575328,);
not I_33683 (I575336,I575328);
nor I_33684 (I575353,I575336,I575234);
and I_33685 (I575370,I575353,I223767);
nor I_33686 (I575387,I575336,I575302);
nor I_33687 (I575183,I575294,I575387);
DFFARX1 I_33688 (I223770,I2683,I575200,I575427,);
nor I_33689 (I575435,I575427,I575294);
not I_33690 (I575452,I575435);
not I_33691 (I575469,I575427);
nor I_33692 (I575486,I575469,I575370);
DFFARX1 I_33693 (I575486,I2683,I575200,I575186,);
nand I_33694 (I575517,I223773,I223782);
and I_33695 (I575534,I575517,I223779);
DFFARX1 I_33696 (I575534,I2683,I575200,I575560,);
nor I_33697 (I575568,I575560,I575427);
DFFARX1 I_33698 (I575568,I2683,I575200,I575168,);
nand I_33699 (I575599,I575560,I575469);
nand I_33700 (I575177,I575452,I575599);
not I_33701 (I575630,I575560);
nor I_33702 (I575647,I575630,I575370);
DFFARX1 I_33703 (I575647,I2683,I575200,I575189,);
nor I_33704 (I575678,I223776,I223782);
or I_33705 (I575180,I575427,I575678);
nor I_33706 (I575171,I575560,I575678);
or I_33707 (I575174,I575294,I575678);
DFFARX1 I_33708 (I575678,I2683,I575200,I575192,);
not I_33709 (I575778,I2690);
DFFARX1 I_33710 (I883124,I2683,I575778,I575804,);
not I_33711 (I575812,I575804);
nand I_33712 (I575829,I883106,I883118);
and I_33713 (I575846,I575829,I883121);
DFFARX1 I_33714 (I575846,I2683,I575778,I575872,);
not I_33715 (I575880,I883115);
DFFARX1 I_33716 (I883112,I2683,I575778,I575906,);
not I_33717 (I575914,I575906);
nor I_33718 (I575931,I575914,I575812);
and I_33719 (I575948,I575931,I883115);
nor I_33720 (I575965,I575914,I575880);
nor I_33721 (I575761,I575872,I575965);
DFFARX1 I_33722 (I883130,I2683,I575778,I576005,);
nor I_33723 (I576013,I576005,I575872);
not I_33724 (I576030,I576013);
not I_33725 (I576047,I576005);
nor I_33726 (I576064,I576047,I575948);
DFFARX1 I_33727 (I576064,I2683,I575778,I575764,);
nand I_33728 (I576095,I883109,I883109);
and I_33729 (I576112,I576095,I883106);
DFFARX1 I_33730 (I576112,I2683,I575778,I576138,);
nor I_33731 (I576146,I576138,I576005);
DFFARX1 I_33732 (I576146,I2683,I575778,I575746,);
nand I_33733 (I576177,I576138,I576047);
nand I_33734 (I575755,I576030,I576177);
not I_33735 (I576208,I576138);
nor I_33736 (I576225,I576208,I575948);
DFFARX1 I_33737 (I576225,I2683,I575778,I575767,);
nor I_33738 (I576256,I883127,I883109);
or I_33739 (I575758,I576005,I576256);
nor I_33740 (I575749,I576138,I576256);
or I_33741 (I575752,I575872,I576256);
DFFARX1 I_33742 (I576256,I2683,I575778,I575770,);
not I_33743 (I576356,I2690);
DFFARX1 I_33744 (I1012850,I2683,I576356,I576382,);
not I_33745 (I576390,I576382);
nand I_33746 (I576407,I1012874,I1012856);
and I_33747 (I576424,I576407,I1012862);
DFFARX1 I_33748 (I576424,I2683,I576356,I576450,);
not I_33749 (I576458,I1012868);
DFFARX1 I_33750 (I1012853,I2683,I576356,I576484,);
not I_33751 (I576492,I576484);
nor I_33752 (I576509,I576492,I576390);
and I_33753 (I576526,I576509,I1012868);
nor I_33754 (I576543,I576492,I576458);
nor I_33755 (I576339,I576450,I576543);
DFFARX1 I_33756 (I1012865,I2683,I576356,I576583,);
nor I_33757 (I576591,I576583,I576450);
not I_33758 (I576608,I576591);
not I_33759 (I576625,I576583);
nor I_33760 (I576642,I576625,I576526);
DFFARX1 I_33761 (I576642,I2683,I576356,I576342,);
nand I_33762 (I576673,I1012871,I1012859);
and I_33763 (I576690,I576673,I1012853);
DFFARX1 I_33764 (I576690,I2683,I576356,I576716,);
nor I_33765 (I576724,I576716,I576583);
DFFARX1 I_33766 (I576724,I2683,I576356,I576324,);
nand I_33767 (I576755,I576716,I576625);
nand I_33768 (I576333,I576608,I576755);
not I_33769 (I576786,I576716);
nor I_33770 (I576803,I576786,I576526);
DFFARX1 I_33771 (I576803,I2683,I576356,I576345,);
nor I_33772 (I576834,I1012850,I1012859);
or I_33773 (I576336,I576583,I576834);
nor I_33774 (I576327,I576716,I576834);
or I_33775 (I576330,I576450,I576834);
DFFARX1 I_33776 (I576834,I2683,I576356,I576348,);
not I_33777 (I576934,I2690);
DFFARX1 I_33778 (I1072156,I2683,I576934,I576960,);
not I_33779 (I576968,I576960);
nand I_33780 (I576985,I1072141,I1072129);
and I_33781 (I577002,I576985,I1072144);
DFFARX1 I_33782 (I577002,I2683,I576934,I577028,);
not I_33783 (I577036,I1072129);
DFFARX1 I_33784 (I1072147,I2683,I576934,I577062,);
not I_33785 (I577070,I577062);
nor I_33786 (I577087,I577070,I576968);
and I_33787 (I577104,I577087,I1072129);
nor I_33788 (I577121,I577070,I577036);
nor I_33789 (I576917,I577028,I577121);
DFFARX1 I_33790 (I1072135,I2683,I576934,I577161,);
nor I_33791 (I577169,I577161,I577028);
not I_33792 (I577186,I577169);
not I_33793 (I577203,I577161);
nor I_33794 (I577220,I577203,I577104);
DFFARX1 I_33795 (I577220,I2683,I576934,I576920,);
nand I_33796 (I577251,I1072132,I1072138);
and I_33797 (I577268,I577251,I1072153);
DFFARX1 I_33798 (I577268,I2683,I576934,I577294,);
nor I_33799 (I577302,I577294,I577161);
DFFARX1 I_33800 (I577302,I2683,I576934,I576902,);
nand I_33801 (I577333,I577294,I577203);
nand I_33802 (I576911,I577186,I577333);
not I_33803 (I577364,I577294);
nor I_33804 (I577381,I577364,I577104);
DFFARX1 I_33805 (I577381,I2683,I576934,I576923,);
nor I_33806 (I577412,I1072150,I1072138);
or I_33807 (I576914,I577161,I577412);
nor I_33808 (I576905,I577294,I577412);
or I_33809 (I576908,I577028,I577412);
DFFARX1 I_33810 (I577412,I2683,I576934,I576926,);
not I_33811 (I577512,I2690);
DFFARX1 I_33812 (I433558,I2683,I577512,I577538,);
not I_33813 (I577546,I577538);
nand I_33814 (I577563,I433567,I433576);
and I_33815 (I577580,I577563,I433582);
DFFARX1 I_33816 (I577580,I2683,I577512,I577606,);
not I_33817 (I577614,I433579);
DFFARX1 I_33818 (I433564,I2683,I577512,I577640,);
not I_33819 (I577648,I577640);
nor I_33820 (I577665,I577648,I577546);
and I_33821 (I577682,I577665,I433579);
nor I_33822 (I577699,I577648,I577614);
nor I_33823 (I577495,I577606,I577699);
DFFARX1 I_33824 (I433573,I2683,I577512,I577739,);
nor I_33825 (I577747,I577739,I577606);
not I_33826 (I577764,I577747);
not I_33827 (I577781,I577739);
nor I_33828 (I577798,I577781,I577682);
DFFARX1 I_33829 (I577798,I2683,I577512,I577498,);
nand I_33830 (I577829,I433570,I433561);
and I_33831 (I577846,I577829,I433558);
DFFARX1 I_33832 (I577846,I2683,I577512,I577872,);
nor I_33833 (I577880,I577872,I577739);
DFFARX1 I_33834 (I577880,I2683,I577512,I577480,);
nand I_33835 (I577911,I577872,I577781);
nand I_33836 (I577489,I577764,I577911);
not I_33837 (I577942,I577872);
nor I_33838 (I577959,I577942,I577682);
DFFARX1 I_33839 (I577959,I2683,I577512,I577501,);
nor I_33840 (I577990,I433561,I433561);
or I_33841 (I577492,I577739,I577990);
nor I_33842 (I577483,I577872,I577990);
or I_33843 (I577486,I577606,I577990);
DFFARX1 I_33844 (I577990,I2683,I577512,I577504,);
not I_33845 (I578090,I2690);
DFFARX1 I_33846 (I491936,I2683,I578090,I578116,);
not I_33847 (I578124,I578116);
nand I_33848 (I578141,I491945,I491954);
and I_33849 (I578158,I578141,I491960);
DFFARX1 I_33850 (I578158,I2683,I578090,I578184,);
not I_33851 (I578192,I491957);
DFFARX1 I_33852 (I491942,I2683,I578090,I578218,);
not I_33853 (I578226,I578218);
nor I_33854 (I578243,I578226,I578124);
and I_33855 (I578260,I578243,I491957);
nor I_33856 (I578277,I578226,I578192);
nor I_33857 (I578073,I578184,I578277);
DFFARX1 I_33858 (I491951,I2683,I578090,I578317,);
nor I_33859 (I578325,I578317,I578184);
not I_33860 (I578342,I578325);
not I_33861 (I578359,I578317);
nor I_33862 (I578376,I578359,I578260);
DFFARX1 I_33863 (I578376,I2683,I578090,I578076,);
nand I_33864 (I578407,I491948,I491939);
and I_33865 (I578424,I578407,I491936);
DFFARX1 I_33866 (I578424,I2683,I578090,I578450,);
nor I_33867 (I578458,I578450,I578317);
DFFARX1 I_33868 (I578458,I2683,I578090,I578058,);
nand I_33869 (I578489,I578450,I578359);
nand I_33870 (I578067,I578342,I578489);
not I_33871 (I578520,I578450);
nor I_33872 (I578537,I578520,I578260);
DFFARX1 I_33873 (I578537,I2683,I578090,I578079,);
nor I_33874 (I578568,I491939,I491939);
or I_33875 (I578070,I578317,I578568);
nor I_33876 (I578061,I578450,I578568);
or I_33877 (I578064,I578184,I578568);
DFFARX1 I_33878 (I578568,I2683,I578090,I578082,);
not I_33879 (I578668,I2690);
DFFARX1 I_33880 (I153925,I2683,I578668,I578694,);
not I_33881 (I578702,I578694);
nand I_33882 (I578719,I153928,I153949);
and I_33883 (I578736,I578719,I153937);
DFFARX1 I_33884 (I578736,I2683,I578668,I578762,);
not I_33885 (I578770,I153934);
DFFARX1 I_33886 (I153925,I2683,I578668,I578796,);
not I_33887 (I578804,I578796);
nor I_33888 (I578821,I578804,I578702);
and I_33889 (I578838,I578821,I153934);
nor I_33890 (I578855,I578804,I578770);
nor I_33891 (I578651,I578762,I578855);
DFFARX1 I_33892 (I153943,I2683,I578668,I578895,);
nor I_33893 (I578903,I578895,I578762);
not I_33894 (I578920,I578903);
not I_33895 (I578937,I578895);
nor I_33896 (I578954,I578937,I578838);
DFFARX1 I_33897 (I578954,I2683,I578668,I578654,);
nand I_33898 (I578985,I153928,I153931);
and I_33899 (I579002,I578985,I153940);
DFFARX1 I_33900 (I579002,I2683,I578668,I579028,);
nor I_33901 (I579036,I579028,I578895);
DFFARX1 I_33902 (I579036,I2683,I578668,I578636,);
nand I_33903 (I579067,I579028,I578937);
nand I_33904 (I578645,I578920,I579067);
not I_33905 (I579098,I579028);
nor I_33906 (I579115,I579098,I578838);
DFFARX1 I_33907 (I579115,I2683,I578668,I578657,);
nor I_33908 (I579146,I153946,I153931);
or I_33909 (I578648,I578895,I579146);
nor I_33910 (I578639,I579028,I579146);
or I_33911 (I578642,I578762,I579146);
DFFARX1 I_33912 (I579146,I2683,I578668,I578660,);
not I_33913 (I579246,I2690);
DFFARX1 I_33914 (I957566,I2683,I579246,I579272,);
not I_33915 (I579280,I579272);
nand I_33916 (I579297,I957569,I957578);
and I_33917 (I579314,I579297,I957581);
DFFARX1 I_33918 (I579314,I2683,I579246,I579340,);
not I_33919 (I579348,I957590);
DFFARX1 I_33920 (I957572,I2683,I579246,I579374,);
not I_33921 (I579382,I579374);
nor I_33922 (I579399,I579382,I579280);
and I_33923 (I579416,I579399,I957590);
nor I_33924 (I579433,I579382,I579348);
nor I_33925 (I579229,I579340,I579433);
DFFARX1 I_33926 (I957569,I2683,I579246,I579473,);
nor I_33927 (I579481,I579473,I579340);
not I_33928 (I579498,I579481);
not I_33929 (I579515,I579473);
nor I_33930 (I579532,I579515,I579416);
DFFARX1 I_33931 (I579532,I2683,I579246,I579232,);
nand I_33932 (I579563,I957587,I957566);
and I_33933 (I579580,I579563,I957584);
DFFARX1 I_33934 (I579580,I2683,I579246,I579606,);
nor I_33935 (I579614,I579606,I579473);
DFFARX1 I_33936 (I579614,I2683,I579246,I579214,);
nand I_33937 (I579645,I579606,I579515);
nand I_33938 (I579223,I579498,I579645);
not I_33939 (I579676,I579606);
nor I_33940 (I579693,I579676,I579416);
DFFARX1 I_33941 (I579693,I2683,I579246,I579235,);
nor I_33942 (I579724,I957575,I957566);
or I_33943 (I579226,I579473,I579724);
nor I_33944 (I579217,I579606,I579724);
or I_33945 (I579220,I579340,I579724);
DFFARX1 I_33946 (I579724,I2683,I579246,I579238,);
not I_33947 (I579824,I2690);
DFFARX1 I_33948 (I934566,I2683,I579824,I579850,);
not I_33949 (I579858,I579850);
nand I_33950 (I579875,I934548,I934560);
and I_33951 (I579892,I579875,I934563);
DFFARX1 I_33952 (I579892,I2683,I579824,I579918,);
not I_33953 (I579926,I934557);
DFFARX1 I_33954 (I934554,I2683,I579824,I579952,);
not I_33955 (I579960,I579952);
nor I_33956 (I579977,I579960,I579858);
and I_33957 (I579994,I579977,I934557);
nor I_33958 (I580011,I579960,I579926);
nor I_33959 (I579807,I579918,I580011);
DFFARX1 I_33960 (I934572,I2683,I579824,I580051,);
nor I_33961 (I580059,I580051,I579918);
not I_33962 (I580076,I580059);
not I_33963 (I580093,I580051);
nor I_33964 (I580110,I580093,I579994);
DFFARX1 I_33965 (I580110,I2683,I579824,I579810,);
nand I_33966 (I580141,I934551,I934551);
and I_33967 (I580158,I580141,I934548);
DFFARX1 I_33968 (I580158,I2683,I579824,I580184,);
nor I_33969 (I580192,I580184,I580051);
DFFARX1 I_33970 (I580192,I2683,I579824,I579792,);
nand I_33971 (I580223,I580184,I580093);
nand I_33972 (I579801,I580076,I580223);
not I_33973 (I580254,I580184);
nor I_33974 (I580271,I580254,I579994);
DFFARX1 I_33975 (I580271,I2683,I579824,I579813,);
nor I_33976 (I580302,I934569,I934551);
or I_33977 (I579804,I580051,I580302);
nor I_33978 (I579795,I580184,I580302);
or I_33979 (I579798,I579918,I580302);
DFFARX1 I_33980 (I580302,I2683,I579824,I579816,);
not I_33981 (I580402,I2690);
DFFARX1 I_33982 (I5674,I2683,I580402,I580428,);
not I_33983 (I580436,I580428);
nand I_33984 (I580453,I5677,I5689);
and I_33985 (I580470,I580453,I5668);
DFFARX1 I_33986 (I580470,I2683,I580402,I580496,);
not I_33987 (I580504,I5668);
DFFARX1 I_33988 (I5671,I2683,I580402,I580530,);
not I_33989 (I580538,I580530);
nor I_33990 (I580555,I580538,I580436);
and I_33991 (I580572,I580555,I5668);
nor I_33992 (I580589,I580538,I580504);
nor I_33993 (I580385,I580496,I580589);
DFFARX1 I_33994 (I5683,I2683,I580402,I580629,);
nor I_33995 (I580637,I580629,I580496);
not I_33996 (I580654,I580637);
not I_33997 (I580671,I580629);
nor I_33998 (I580688,I580671,I580572);
DFFARX1 I_33999 (I580688,I2683,I580402,I580388,);
nand I_34000 (I580719,I5686,I5671);
and I_34001 (I580736,I580719,I5680);
DFFARX1 I_34002 (I580736,I2683,I580402,I580762,);
nor I_34003 (I580770,I580762,I580629);
DFFARX1 I_34004 (I580770,I2683,I580402,I580370,);
nand I_34005 (I580801,I580762,I580671);
nand I_34006 (I580379,I580654,I580801);
not I_34007 (I580832,I580762);
nor I_34008 (I580849,I580832,I580572);
DFFARX1 I_34009 (I580849,I2683,I580402,I580391,);
nor I_34010 (I580880,I5674,I5671);
or I_34011 (I580382,I580629,I580880);
nor I_34012 (I580373,I580762,I580880);
or I_34013 (I580376,I580496,I580880);
DFFARX1 I_34014 (I580880,I2683,I580402,I580394,);
not I_34015 (I580980,I2690);
DFFARX1 I_34016 (I629651,I2683,I580980,I581006,);
not I_34017 (I581014,I581006);
nand I_34018 (I581031,I629639,I629657);
and I_34019 (I581048,I581031,I629654);
DFFARX1 I_34020 (I581048,I2683,I580980,I581074,);
not I_34021 (I581082,I629645);
DFFARX1 I_34022 (I629642,I2683,I580980,I581108,);
not I_34023 (I581116,I581108);
nor I_34024 (I581133,I581116,I581014);
and I_34025 (I581150,I581133,I629645);
nor I_34026 (I581167,I581116,I581082);
nor I_34027 (I580963,I581074,I581167);
DFFARX1 I_34028 (I629636,I2683,I580980,I581207,);
nor I_34029 (I581215,I581207,I581074);
not I_34030 (I581232,I581215);
not I_34031 (I581249,I581207);
nor I_34032 (I581266,I581249,I581150);
DFFARX1 I_34033 (I581266,I2683,I580980,I580966,);
nand I_34034 (I581297,I629636,I629639);
and I_34035 (I581314,I581297,I629642);
DFFARX1 I_34036 (I581314,I2683,I580980,I581340,);
nor I_34037 (I581348,I581340,I581207);
DFFARX1 I_34038 (I581348,I2683,I580980,I580948,);
nand I_34039 (I581379,I581340,I581249);
nand I_34040 (I580957,I581232,I581379);
not I_34041 (I581410,I581340);
nor I_34042 (I581427,I581410,I581150);
DFFARX1 I_34043 (I581427,I2683,I580980,I580969,);
nor I_34044 (I581458,I629648,I629639);
or I_34045 (I580960,I581207,I581458);
nor I_34046 (I580951,I581340,I581458);
or I_34047 (I580954,I581074,I581458);
DFFARX1 I_34048 (I581458,I2683,I580980,I580972,);
not I_34049 (I581558,I2690);
DFFARX1 I_34050 (I371483,I2683,I581558,I581584,);
not I_34051 (I581592,I581584);
nand I_34052 (I581609,I371474,I371492);
and I_34053 (I581626,I581609,I371495);
DFFARX1 I_34054 (I581626,I2683,I581558,I581652,);
not I_34055 (I581660,I371489);
DFFARX1 I_34056 (I371477,I2683,I581558,I581686,);
not I_34057 (I581694,I581686);
nor I_34058 (I581711,I581694,I581592);
and I_34059 (I581728,I581711,I371489);
nor I_34060 (I581745,I581694,I581660);
nor I_34061 (I581541,I581652,I581745);
DFFARX1 I_34062 (I371486,I2683,I581558,I581785,);
nor I_34063 (I581793,I581785,I581652);
not I_34064 (I581810,I581793);
not I_34065 (I581827,I581785);
nor I_34066 (I581844,I581827,I581728);
DFFARX1 I_34067 (I581844,I2683,I581558,I581544,);
nand I_34068 (I581875,I371501,I371498);
and I_34069 (I581892,I581875,I371480);
DFFARX1 I_34070 (I581892,I2683,I581558,I581918,);
nor I_34071 (I581926,I581918,I581785);
DFFARX1 I_34072 (I581926,I2683,I581558,I581526,);
nand I_34073 (I581957,I581918,I581827);
nand I_34074 (I581535,I581810,I581957);
not I_34075 (I581988,I581918);
nor I_34076 (I582005,I581988,I581728);
DFFARX1 I_34077 (I582005,I2683,I581558,I581547,);
nor I_34078 (I582036,I371474,I371498);
or I_34079 (I581538,I581785,I582036);
nor I_34080 (I581529,I581918,I582036);
or I_34081 (I581532,I581652,I582036);
DFFARX1 I_34082 (I582036,I2683,I581558,I581550,);
not I_34083 (I582136,I2690);
DFFARX1 I_34084 (I301781,I2683,I582136,I582162,);
not I_34085 (I582170,I582162);
nand I_34086 (I582187,I301784,I301760);
and I_34087 (I582204,I582187,I301757);
DFFARX1 I_34088 (I582204,I2683,I582136,I582230,);
not I_34089 (I582238,I301763);
DFFARX1 I_34090 (I301757,I2683,I582136,I582264,);
not I_34091 (I582272,I582264);
nor I_34092 (I582289,I582272,I582170);
and I_34093 (I582306,I582289,I301763);
nor I_34094 (I582323,I582272,I582238);
nor I_34095 (I582119,I582230,I582323);
DFFARX1 I_34096 (I301766,I2683,I582136,I582363,);
nor I_34097 (I582371,I582363,I582230);
not I_34098 (I582388,I582371);
not I_34099 (I582405,I582363);
nor I_34100 (I582422,I582405,I582306);
DFFARX1 I_34101 (I582422,I2683,I582136,I582122,);
nand I_34102 (I582453,I301769,I301778);
and I_34103 (I582470,I582453,I301775);
DFFARX1 I_34104 (I582470,I2683,I582136,I582496,);
nor I_34105 (I582504,I582496,I582363);
DFFARX1 I_34106 (I582504,I2683,I582136,I582104,);
nand I_34107 (I582535,I582496,I582405);
nand I_34108 (I582113,I582388,I582535);
not I_34109 (I582566,I582496);
nor I_34110 (I582583,I582566,I582306);
DFFARX1 I_34111 (I582583,I2683,I582136,I582125,);
nor I_34112 (I582614,I301772,I301778);
or I_34113 (I582116,I582363,I582614);
nor I_34114 (I582107,I582496,I582614);
or I_34115 (I582110,I582230,I582614);
DFFARX1 I_34116 (I582614,I2683,I582136,I582128,);
not I_34117 (I582714,I2690);
DFFARX1 I_34118 (I177725,I2683,I582714,I582740,);
not I_34119 (I582748,I582740);
nand I_34120 (I582765,I177728,I177749);
and I_34121 (I582782,I582765,I177737);
DFFARX1 I_34122 (I582782,I2683,I582714,I582808,);
not I_34123 (I582816,I177734);
DFFARX1 I_34124 (I177725,I2683,I582714,I582842,);
not I_34125 (I582850,I582842);
nor I_34126 (I582867,I582850,I582748);
and I_34127 (I582884,I582867,I177734);
nor I_34128 (I582901,I582850,I582816);
nor I_34129 (I582697,I582808,I582901);
DFFARX1 I_34130 (I177743,I2683,I582714,I582941,);
nor I_34131 (I582949,I582941,I582808);
not I_34132 (I582966,I582949);
not I_34133 (I582983,I582941);
nor I_34134 (I583000,I582983,I582884);
DFFARX1 I_34135 (I583000,I2683,I582714,I582700,);
nand I_34136 (I583031,I177728,I177731);
and I_34137 (I583048,I583031,I177740);
DFFARX1 I_34138 (I583048,I2683,I582714,I583074,);
nor I_34139 (I583082,I583074,I582941);
DFFARX1 I_34140 (I583082,I2683,I582714,I582682,);
nand I_34141 (I583113,I583074,I582983);
nand I_34142 (I582691,I582966,I583113);
not I_34143 (I583144,I583074);
nor I_34144 (I583161,I583144,I582884);
DFFARX1 I_34145 (I583161,I2683,I582714,I582703,);
nor I_34146 (I583192,I177746,I177731);
or I_34147 (I582694,I582941,I583192);
nor I_34148 (I582685,I583074,I583192);
or I_34149 (I582688,I582808,I583192);
DFFARX1 I_34150 (I583192,I2683,I582714,I582706,);
not I_34151 (I583292,I2690);
DFFARX1 I_34152 (I145000,I2683,I583292,I583318,);
not I_34153 (I583326,I583318);
nand I_34154 (I583343,I145003,I145024);
and I_34155 (I583360,I583343,I145012);
DFFARX1 I_34156 (I583360,I2683,I583292,I583386,);
not I_34157 (I583394,I145009);
DFFARX1 I_34158 (I145000,I2683,I583292,I583420,);
not I_34159 (I583428,I583420);
nor I_34160 (I583445,I583428,I583326);
and I_34161 (I583462,I583445,I145009);
nor I_34162 (I583479,I583428,I583394);
nor I_34163 (I583275,I583386,I583479);
DFFARX1 I_34164 (I145018,I2683,I583292,I583519,);
nor I_34165 (I583527,I583519,I583386);
not I_34166 (I583544,I583527);
not I_34167 (I583561,I583519);
nor I_34168 (I583578,I583561,I583462);
DFFARX1 I_34169 (I583578,I2683,I583292,I583278,);
nand I_34170 (I583609,I145003,I145006);
and I_34171 (I583626,I583609,I145015);
DFFARX1 I_34172 (I583626,I2683,I583292,I583652,);
nor I_34173 (I583660,I583652,I583519);
DFFARX1 I_34174 (I583660,I2683,I583292,I583260,);
nand I_34175 (I583691,I583652,I583561);
nand I_34176 (I583269,I583544,I583691);
not I_34177 (I583722,I583652);
nor I_34178 (I583739,I583722,I583462);
DFFARX1 I_34179 (I583739,I2683,I583292,I583281,);
nor I_34180 (I583770,I145021,I145006);
or I_34181 (I583272,I583519,I583770);
nor I_34182 (I583263,I583652,I583770);
or I_34183 (I583266,I583386,I583770);
DFFARX1 I_34184 (I583770,I2683,I583292,I583284,);
not I_34185 (I583870,I2690);
DFFARX1 I_34186 (I230109,I2683,I583870,I583896,);
not I_34187 (I583904,I583896);
nand I_34188 (I583921,I230112,I230088);
and I_34189 (I583938,I583921,I230085);
DFFARX1 I_34190 (I583938,I2683,I583870,I583964,);
not I_34191 (I583972,I230091);
DFFARX1 I_34192 (I230085,I2683,I583870,I583998,);
not I_34193 (I584006,I583998);
nor I_34194 (I584023,I584006,I583904);
and I_34195 (I584040,I584023,I230091);
nor I_34196 (I584057,I584006,I583972);
nor I_34197 (I583853,I583964,I584057);
DFFARX1 I_34198 (I230094,I2683,I583870,I584097,);
nor I_34199 (I584105,I584097,I583964);
not I_34200 (I584122,I584105);
not I_34201 (I584139,I584097);
nor I_34202 (I584156,I584139,I584040);
DFFARX1 I_34203 (I584156,I2683,I583870,I583856,);
nand I_34204 (I584187,I230097,I230106);
and I_34205 (I584204,I584187,I230103);
DFFARX1 I_34206 (I584204,I2683,I583870,I584230,);
nor I_34207 (I584238,I584230,I584097);
DFFARX1 I_34208 (I584238,I2683,I583870,I583838,);
nand I_34209 (I584269,I584230,I584139);
nand I_34210 (I583847,I584122,I584269);
not I_34211 (I584300,I584230);
nor I_34212 (I584317,I584300,I584040);
DFFARX1 I_34213 (I584317,I2683,I583870,I583859,);
nor I_34214 (I584348,I230100,I230106);
or I_34215 (I583850,I584097,I584348);
nor I_34216 (I583841,I584230,I584348);
or I_34217 (I583844,I583964,I584348);
DFFARX1 I_34218 (I584348,I2683,I583870,I583862,);
not I_34219 (I584448,I2690);
DFFARX1 I_34220 (I627543,I2683,I584448,I584474,);
not I_34221 (I584482,I584474);
nand I_34222 (I584499,I627531,I627549);
and I_34223 (I584516,I584499,I627546);
DFFARX1 I_34224 (I584516,I2683,I584448,I584542,);
not I_34225 (I584550,I627537);
DFFARX1 I_34226 (I627534,I2683,I584448,I584576,);
not I_34227 (I584584,I584576);
nor I_34228 (I584601,I584584,I584482);
and I_34229 (I584618,I584601,I627537);
nor I_34230 (I584635,I584584,I584550);
nor I_34231 (I584431,I584542,I584635);
DFFARX1 I_34232 (I627528,I2683,I584448,I584675,);
nor I_34233 (I584683,I584675,I584542);
not I_34234 (I584700,I584683);
not I_34235 (I584717,I584675);
nor I_34236 (I584734,I584717,I584618);
DFFARX1 I_34237 (I584734,I2683,I584448,I584434,);
nand I_34238 (I584765,I627528,I627531);
and I_34239 (I584782,I584765,I627534);
DFFARX1 I_34240 (I584782,I2683,I584448,I584808,);
nor I_34241 (I584816,I584808,I584675);
DFFARX1 I_34242 (I584816,I2683,I584448,I584416,);
nand I_34243 (I584847,I584808,I584717);
nand I_34244 (I584425,I584700,I584847);
not I_34245 (I584878,I584808);
nor I_34246 (I584895,I584878,I584618);
DFFARX1 I_34247 (I584895,I2683,I584448,I584437,);
nor I_34248 (I584926,I627540,I627531);
or I_34249 (I584428,I584675,I584926);
nor I_34250 (I584419,I584808,I584926);
or I_34251 (I584422,I584542,I584926);
DFFARX1 I_34252 (I584926,I2683,I584448,I584440,);
not I_34253 (I585026,I2690);
DFFARX1 I_34254 (I316539,I2683,I585026,I585052,);
not I_34255 (I585060,I585052);
nand I_34256 (I585077,I316530,I316548);
and I_34257 (I585094,I585077,I316551);
DFFARX1 I_34258 (I585094,I2683,I585026,I585120,);
not I_34259 (I585128,I316545);
DFFARX1 I_34260 (I316533,I2683,I585026,I585154,);
not I_34261 (I585162,I585154);
nor I_34262 (I585179,I585162,I585060);
and I_34263 (I585196,I585179,I316545);
nor I_34264 (I585213,I585162,I585128);
nor I_34265 (I585009,I585120,I585213);
DFFARX1 I_34266 (I316542,I2683,I585026,I585253,);
nor I_34267 (I585261,I585253,I585120);
not I_34268 (I585278,I585261);
not I_34269 (I585295,I585253);
nor I_34270 (I585312,I585295,I585196);
DFFARX1 I_34271 (I585312,I2683,I585026,I585012,);
nand I_34272 (I585343,I316557,I316554);
and I_34273 (I585360,I585343,I316536);
DFFARX1 I_34274 (I585360,I2683,I585026,I585386,);
nor I_34275 (I585394,I585386,I585253);
DFFARX1 I_34276 (I585394,I2683,I585026,I584994,);
nand I_34277 (I585425,I585386,I585295);
nand I_34278 (I585003,I585278,I585425);
not I_34279 (I585456,I585386);
nor I_34280 (I585473,I585456,I585196);
DFFARX1 I_34281 (I585473,I2683,I585026,I585015,);
nor I_34282 (I585504,I316530,I316554);
or I_34283 (I585006,I585253,I585504);
nor I_34284 (I584997,I585386,I585504);
or I_34285 (I585000,I585120,I585504);
DFFARX1 I_34286 (I585504,I2683,I585026,I585018,);
not I_34287 (I585604,I2690);
DFFARX1 I_34288 (I136075,I2683,I585604,I585630,);
not I_34289 (I585638,I585630);
nand I_34290 (I585655,I136078,I136099);
and I_34291 (I585672,I585655,I136087);
DFFARX1 I_34292 (I585672,I2683,I585604,I585698,);
not I_34293 (I585706,I136084);
DFFARX1 I_34294 (I136075,I2683,I585604,I585732,);
not I_34295 (I585740,I585732);
nor I_34296 (I585757,I585740,I585638);
and I_34297 (I585774,I585757,I136084);
nor I_34298 (I585791,I585740,I585706);
nor I_34299 (I585587,I585698,I585791);
DFFARX1 I_34300 (I136093,I2683,I585604,I585831,);
nor I_34301 (I585839,I585831,I585698);
not I_34302 (I585856,I585839);
not I_34303 (I585873,I585831);
nor I_34304 (I585890,I585873,I585774);
DFFARX1 I_34305 (I585890,I2683,I585604,I585590,);
nand I_34306 (I585921,I136078,I136081);
and I_34307 (I585938,I585921,I136090);
DFFARX1 I_34308 (I585938,I2683,I585604,I585964,);
nor I_34309 (I585972,I585964,I585831);
DFFARX1 I_34310 (I585972,I2683,I585604,I585572,);
nand I_34311 (I586003,I585964,I585873);
nand I_34312 (I585581,I585856,I586003);
not I_34313 (I586034,I585964);
nor I_34314 (I586051,I586034,I585774);
DFFARX1 I_34315 (I586051,I2683,I585604,I585593,);
nor I_34316 (I586082,I136096,I136081);
or I_34317 (I585584,I585831,I586082);
nor I_34318 (I585575,I585964,I586082);
or I_34319 (I585578,I585698,I586082);
DFFARX1 I_34320 (I586082,I2683,I585604,I585596,);
not I_34321 (I586182,I2690);
DFFARX1 I_34322 (I623854,I2683,I586182,I586208,);
not I_34323 (I586216,I586208);
nand I_34324 (I586233,I623842,I623860);
and I_34325 (I586250,I586233,I623857);
DFFARX1 I_34326 (I586250,I2683,I586182,I586276,);
not I_34327 (I586284,I623848);
DFFARX1 I_34328 (I623845,I2683,I586182,I586310,);
not I_34329 (I586318,I586310);
nor I_34330 (I586335,I586318,I586216);
and I_34331 (I586352,I586335,I623848);
nor I_34332 (I586369,I586318,I586284);
nor I_34333 (I586165,I586276,I586369);
DFFARX1 I_34334 (I623839,I2683,I586182,I586409,);
nor I_34335 (I586417,I586409,I586276);
not I_34336 (I586434,I586417);
not I_34337 (I586451,I586409);
nor I_34338 (I586468,I586451,I586352);
DFFARX1 I_34339 (I586468,I2683,I586182,I586168,);
nand I_34340 (I586499,I623839,I623842);
and I_34341 (I586516,I586499,I623845);
DFFARX1 I_34342 (I586516,I2683,I586182,I586542,);
nor I_34343 (I586550,I586542,I586409);
DFFARX1 I_34344 (I586550,I2683,I586182,I586150,);
nand I_34345 (I586581,I586542,I586451);
nand I_34346 (I586159,I586434,I586581);
not I_34347 (I586612,I586542);
nor I_34348 (I586629,I586612,I586352);
DFFARX1 I_34349 (I586629,I2683,I586182,I586171,);
nor I_34350 (I586660,I623851,I623842);
or I_34351 (I586162,I586409,I586660);
nor I_34352 (I586153,I586542,I586660);
or I_34353 (I586156,I586276,I586660);
DFFARX1 I_34354 (I586660,I2683,I586182,I586174,);
not I_34355 (I586760,I2690);
DFFARX1 I_34356 (I759421,I2683,I586760,I586786,);
not I_34357 (I586794,I586786);
nand I_34358 (I586811,I759397,I759412);
and I_34359 (I586828,I586811,I759424);
DFFARX1 I_34360 (I586828,I2683,I586760,I586854,);
not I_34361 (I586862,I759409);
DFFARX1 I_34362 (I759400,I2683,I586760,I586888,);
not I_34363 (I586896,I586888);
nor I_34364 (I586913,I586896,I586794);
and I_34365 (I586930,I586913,I759409);
nor I_34366 (I586947,I586896,I586862);
nor I_34367 (I586743,I586854,I586947);
DFFARX1 I_34368 (I759397,I2683,I586760,I586987,);
nor I_34369 (I586995,I586987,I586854);
not I_34370 (I587012,I586995);
not I_34371 (I587029,I586987);
nor I_34372 (I587046,I587029,I586930);
DFFARX1 I_34373 (I587046,I2683,I586760,I586746,);
nand I_34374 (I587077,I759415,I759406);
and I_34375 (I587094,I587077,I759418);
DFFARX1 I_34376 (I587094,I2683,I586760,I587120,);
nor I_34377 (I587128,I587120,I586987);
DFFARX1 I_34378 (I587128,I2683,I586760,I586728,);
nand I_34379 (I587159,I587120,I587029);
nand I_34380 (I586737,I587012,I587159);
not I_34381 (I587190,I587120);
nor I_34382 (I587207,I587190,I586930);
DFFARX1 I_34383 (I587207,I2683,I586760,I586749,);
nor I_34384 (I587238,I759403,I759406);
or I_34385 (I586740,I586987,I587238);
nor I_34386 (I586731,I587120,I587238);
or I_34387 (I586734,I586854,I587238);
DFFARX1 I_34388 (I587238,I2683,I586760,I586752,);
not I_34389 (I587338,I2690);
DFFARX1 I_34390 (I13211,I2683,I587338,I587364,);
not I_34391 (I587372,I587364);
nand I_34392 (I587389,I13208,I13199);
and I_34393 (I587406,I587389,I13199);
DFFARX1 I_34394 (I587406,I2683,I587338,I587432,);
not I_34395 (I587440,I13202);
DFFARX1 I_34396 (I13217,I2683,I587338,I587466,);
not I_34397 (I587474,I587466);
nor I_34398 (I587491,I587474,I587372);
and I_34399 (I587508,I587491,I13202);
nor I_34400 (I587525,I587474,I587440);
nor I_34401 (I587321,I587432,I587525);
DFFARX1 I_34402 (I13202,I2683,I587338,I587565,);
nor I_34403 (I587573,I587565,I587432);
not I_34404 (I587590,I587573);
not I_34405 (I587607,I587565);
nor I_34406 (I587624,I587607,I587508);
DFFARX1 I_34407 (I587624,I2683,I587338,I587324,);
nand I_34408 (I587655,I13220,I13205);
and I_34409 (I587672,I587655,I13223);
DFFARX1 I_34410 (I587672,I2683,I587338,I587698,);
nor I_34411 (I587706,I587698,I587565);
DFFARX1 I_34412 (I587706,I2683,I587338,I587306,);
nand I_34413 (I587737,I587698,I587607);
nand I_34414 (I587315,I587590,I587737);
not I_34415 (I587768,I587698);
nor I_34416 (I587785,I587768,I587508);
DFFARX1 I_34417 (I587785,I2683,I587338,I587327,);
nor I_34418 (I587816,I13214,I13205);
or I_34419 (I587318,I587565,I587816);
nor I_34420 (I587309,I587698,I587816);
or I_34421 (I587312,I587432,I587816);
DFFARX1 I_34422 (I587816,I2683,I587338,I587330,);
not I_34423 (I587916,I2690);
DFFARX1 I_34424 (I328507,I2683,I587916,I587942,);
not I_34425 (I587950,I587942);
nand I_34426 (I587967,I328498,I328516);
and I_34427 (I587984,I587967,I328519);
DFFARX1 I_34428 (I587984,I2683,I587916,I588010,);
not I_34429 (I588018,I328513);
DFFARX1 I_34430 (I328501,I2683,I587916,I588044,);
not I_34431 (I588052,I588044);
nor I_34432 (I588069,I588052,I587950);
and I_34433 (I588086,I588069,I328513);
nor I_34434 (I588103,I588052,I588018);
nor I_34435 (I587899,I588010,I588103);
DFFARX1 I_34436 (I328510,I2683,I587916,I588143,);
nor I_34437 (I588151,I588143,I588010);
not I_34438 (I588168,I588151);
not I_34439 (I588185,I588143);
nor I_34440 (I588202,I588185,I588086);
DFFARX1 I_34441 (I588202,I2683,I587916,I587902,);
nand I_34442 (I588233,I328525,I328522);
and I_34443 (I588250,I588233,I328504);
DFFARX1 I_34444 (I588250,I2683,I587916,I588276,);
nor I_34445 (I588284,I588276,I588143);
DFFARX1 I_34446 (I588284,I2683,I587916,I587884,);
nand I_34447 (I588315,I588276,I588185);
nand I_34448 (I587893,I588168,I588315);
not I_34449 (I588346,I588276);
nor I_34450 (I588363,I588346,I588086);
DFFARX1 I_34451 (I588363,I2683,I587916,I587905,);
nor I_34452 (I588394,I328498,I328522);
or I_34453 (I587896,I588143,I588394);
nor I_34454 (I587887,I588276,I588394);
or I_34455 (I587890,I588010,I588394);
DFFARX1 I_34456 (I588394,I2683,I587916,I587908,);
not I_34457 (I588494,I2690);
DFFARX1 I_34458 (I211045,I2683,I588494,I588520,);
not I_34459 (I588528,I588520);
nand I_34460 (I588545,I211048,I211069);
and I_34461 (I588562,I588545,I211057);
DFFARX1 I_34462 (I588562,I2683,I588494,I588588,);
not I_34463 (I588596,I211054);
DFFARX1 I_34464 (I211045,I2683,I588494,I588622,);
not I_34465 (I588630,I588622);
nor I_34466 (I588647,I588630,I588528);
and I_34467 (I588664,I588647,I211054);
nor I_34468 (I588681,I588630,I588596);
nor I_34469 (I588477,I588588,I588681);
DFFARX1 I_34470 (I211063,I2683,I588494,I588721,);
nor I_34471 (I588729,I588721,I588588);
not I_34472 (I588746,I588729);
not I_34473 (I588763,I588721);
nor I_34474 (I588780,I588763,I588664);
DFFARX1 I_34475 (I588780,I2683,I588494,I588480,);
nand I_34476 (I588811,I211048,I211051);
and I_34477 (I588828,I588811,I211060);
DFFARX1 I_34478 (I588828,I2683,I588494,I588854,);
nor I_34479 (I588862,I588854,I588721);
DFFARX1 I_34480 (I588862,I2683,I588494,I588462,);
nand I_34481 (I588893,I588854,I588763);
nand I_34482 (I588471,I588746,I588893);
not I_34483 (I588924,I588854);
nor I_34484 (I588941,I588924,I588664);
DFFARX1 I_34485 (I588941,I2683,I588494,I588483,);
nor I_34486 (I588972,I211066,I211051);
or I_34487 (I588474,I588721,I588972);
nor I_34488 (I588465,I588854,I588972);
or I_34489 (I588468,I588588,I588972);
DFFARX1 I_34490 (I588972,I2683,I588494,I588486,);
not I_34491 (I589072,I2690);
DFFARX1 I_34492 (I883702,I2683,I589072,I589098,);
not I_34493 (I589106,I589098);
nand I_34494 (I589123,I883684,I883696);
and I_34495 (I589140,I589123,I883699);
DFFARX1 I_34496 (I589140,I2683,I589072,I589166,);
not I_34497 (I589174,I883693);
DFFARX1 I_34498 (I883690,I2683,I589072,I589200,);
not I_34499 (I589208,I589200);
nor I_34500 (I589225,I589208,I589106);
and I_34501 (I589242,I589225,I883693);
nor I_34502 (I589259,I589208,I589174);
nor I_34503 (I589055,I589166,I589259);
DFFARX1 I_34504 (I883708,I2683,I589072,I589299,);
nor I_34505 (I589307,I589299,I589166);
not I_34506 (I589324,I589307);
not I_34507 (I589341,I589299);
nor I_34508 (I589358,I589341,I589242);
DFFARX1 I_34509 (I589358,I2683,I589072,I589058,);
nand I_34510 (I589389,I883687,I883687);
and I_34511 (I589406,I589389,I883684);
DFFARX1 I_34512 (I589406,I2683,I589072,I589432,);
nor I_34513 (I589440,I589432,I589299);
DFFARX1 I_34514 (I589440,I2683,I589072,I589040,);
nand I_34515 (I589471,I589432,I589341);
nand I_34516 (I589049,I589324,I589471);
not I_34517 (I589502,I589432);
nor I_34518 (I589519,I589502,I589242);
DFFARX1 I_34519 (I589519,I2683,I589072,I589061,);
nor I_34520 (I589550,I883705,I883687);
or I_34521 (I589052,I589299,I589550);
nor I_34522 (I589043,I589432,I589550);
or I_34523 (I589046,I589166,I589550);
DFFARX1 I_34524 (I589550,I2683,I589072,I589064,);
not I_34525 (I589650,I2690);
DFFARX1 I_34526 (I746501,I2683,I589650,I589676,);
not I_34527 (I589684,I589676);
nand I_34528 (I589701,I746477,I746492);
and I_34529 (I589718,I589701,I746504);
DFFARX1 I_34530 (I589718,I2683,I589650,I589744,);
not I_34531 (I589752,I746489);
DFFARX1 I_34532 (I746480,I2683,I589650,I589778,);
not I_34533 (I589786,I589778);
nor I_34534 (I589803,I589786,I589684);
and I_34535 (I589820,I589803,I746489);
nor I_34536 (I589837,I589786,I589752);
nor I_34537 (I589633,I589744,I589837);
DFFARX1 I_34538 (I746477,I2683,I589650,I589877,);
nor I_34539 (I589885,I589877,I589744);
not I_34540 (I589902,I589885);
not I_34541 (I589919,I589877);
nor I_34542 (I589936,I589919,I589820);
DFFARX1 I_34543 (I589936,I2683,I589650,I589636,);
nand I_34544 (I589967,I746495,I746486);
and I_34545 (I589984,I589967,I746498);
DFFARX1 I_34546 (I589984,I2683,I589650,I590010,);
nor I_34547 (I590018,I590010,I589877);
DFFARX1 I_34548 (I590018,I2683,I589650,I589618,);
nand I_34549 (I590049,I590010,I589919);
nand I_34550 (I589627,I589902,I590049);
not I_34551 (I590080,I590010);
nor I_34552 (I590097,I590080,I589820);
DFFARX1 I_34553 (I590097,I2683,I589650,I589639,);
nor I_34554 (I590128,I746483,I746486);
or I_34555 (I589630,I589877,I590128);
nor I_34556 (I589621,I590010,I590128);
or I_34557 (I589624,I589744,I590128);
DFFARX1 I_34558 (I590128,I2683,I589650,I589642,);
not I_34559 (I590228,I2690);
DFFARX1 I_34560 (I266472,I2683,I590228,I590254,);
not I_34561 (I590262,I590254);
nand I_34562 (I590279,I266475,I266451);
and I_34563 (I590296,I590279,I266448);
DFFARX1 I_34564 (I590296,I2683,I590228,I590322,);
not I_34565 (I590330,I266454);
DFFARX1 I_34566 (I266448,I2683,I590228,I590356,);
not I_34567 (I590364,I590356);
nor I_34568 (I590381,I590364,I590262);
and I_34569 (I590398,I590381,I266454);
nor I_34570 (I590415,I590364,I590330);
nor I_34571 (I590211,I590322,I590415);
DFFARX1 I_34572 (I266457,I2683,I590228,I590455,);
nor I_34573 (I590463,I590455,I590322);
not I_34574 (I590480,I590463);
not I_34575 (I590497,I590455);
nor I_34576 (I590514,I590497,I590398);
DFFARX1 I_34577 (I590514,I2683,I590228,I590214,);
nand I_34578 (I590545,I266460,I266469);
and I_34579 (I590562,I590545,I266466);
DFFARX1 I_34580 (I590562,I2683,I590228,I590588,);
nor I_34581 (I590596,I590588,I590455);
DFFARX1 I_34582 (I590596,I2683,I590228,I590196,);
nand I_34583 (I590627,I590588,I590497);
nand I_34584 (I590205,I590480,I590627);
not I_34585 (I590658,I590588);
nor I_34586 (I590675,I590658,I590398);
DFFARX1 I_34587 (I590675,I2683,I590228,I590217,);
nor I_34588 (I590706,I266463,I266469);
or I_34589 (I590208,I590455,I590706);
nor I_34590 (I590199,I590588,I590706);
or I_34591 (I590202,I590322,I590706);
DFFARX1 I_34592 (I590706,I2683,I590228,I590220,);
not I_34593 (I590806,I2690);
DFFARX1 I_34594 (I849022,I2683,I590806,I590832,);
not I_34595 (I590840,I590832);
nand I_34596 (I590857,I849004,I849016);
and I_34597 (I590874,I590857,I849019);
DFFARX1 I_34598 (I590874,I2683,I590806,I590900,);
not I_34599 (I590908,I849013);
DFFARX1 I_34600 (I849010,I2683,I590806,I590934,);
not I_34601 (I590942,I590934);
nor I_34602 (I590959,I590942,I590840);
and I_34603 (I590976,I590959,I849013);
nor I_34604 (I590993,I590942,I590908);
nor I_34605 (I590789,I590900,I590993);
DFFARX1 I_34606 (I849028,I2683,I590806,I591033,);
nor I_34607 (I591041,I591033,I590900);
not I_34608 (I591058,I591041);
not I_34609 (I591075,I591033);
nor I_34610 (I591092,I591075,I590976);
DFFARX1 I_34611 (I591092,I2683,I590806,I590792,);
nand I_34612 (I591123,I849007,I849007);
and I_34613 (I591140,I591123,I849004);
DFFARX1 I_34614 (I591140,I2683,I590806,I591166,);
nor I_34615 (I591174,I591166,I591033);
DFFARX1 I_34616 (I591174,I2683,I590806,I590774,);
nand I_34617 (I591205,I591166,I591075);
nand I_34618 (I590783,I591058,I591205);
not I_34619 (I591236,I591166);
nor I_34620 (I591253,I591236,I590976);
DFFARX1 I_34621 (I591253,I2683,I590806,I590795,);
nor I_34622 (I591284,I849025,I849007);
or I_34623 (I590786,I591033,I591284);
nor I_34624 (I590777,I591166,I591284);
or I_34625 (I590780,I590900,I591284);
DFFARX1 I_34626 (I591284,I2683,I590806,I590798,);
not I_34627 (I591384,I2690);
DFFARX1 I_34628 (I993198,I2683,I591384,I591410,);
not I_34629 (I591418,I591410);
nand I_34630 (I591435,I993222,I993204);
and I_34631 (I591452,I591435,I993210);
DFFARX1 I_34632 (I591452,I2683,I591384,I591478,);
not I_34633 (I591486,I993216);
DFFARX1 I_34634 (I993201,I2683,I591384,I591512,);
not I_34635 (I591520,I591512);
nor I_34636 (I591537,I591520,I591418);
and I_34637 (I591554,I591537,I993216);
nor I_34638 (I591571,I591520,I591486);
nor I_34639 (I591367,I591478,I591571);
DFFARX1 I_34640 (I993213,I2683,I591384,I591611,);
nor I_34641 (I591619,I591611,I591478);
not I_34642 (I591636,I591619);
not I_34643 (I591653,I591611);
nor I_34644 (I591670,I591653,I591554);
DFFARX1 I_34645 (I591670,I2683,I591384,I591370,);
nand I_34646 (I591701,I993219,I993207);
and I_34647 (I591718,I591701,I993201);
DFFARX1 I_34648 (I591718,I2683,I591384,I591744,);
nor I_34649 (I591752,I591744,I591611);
DFFARX1 I_34650 (I591752,I2683,I591384,I591352,);
nand I_34651 (I591783,I591744,I591653);
nand I_34652 (I591361,I591636,I591783);
not I_34653 (I591814,I591744);
nor I_34654 (I591831,I591814,I591554);
DFFARX1 I_34655 (I591831,I2683,I591384,I591373,);
nor I_34656 (I591862,I993198,I993207);
or I_34657 (I591364,I591611,I591862);
nor I_34658 (I591355,I591744,I591862);
or I_34659 (I591358,I591478,I591862);
DFFARX1 I_34660 (I591862,I2683,I591384,I591376,);
not I_34661 (I591962,I2690);
DFFARX1 I_34662 (I879078,I2683,I591962,I591988,);
not I_34663 (I591996,I591988);
nand I_34664 (I592013,I879060,I879072);
and I_34665 (I592030,I592013,I879075);
DFFARX1 I_34666 (I592030,I2683,I591962,I592056,);
not I_34667 (I592064,I879069);
DFFARX1 I_34668 (I879066,I2683,I591962,I592090,);
not I_34669 (I592098,I592090);
nor I_34670 (I592115,I592098,I591996);
and I_34671 (I592132,I592115,I879069);
nor I_34672 (I592149,I592098,I592064);
nor I_34673 (I591945,I592056,I592149);
DFFARX1 I_34674 (I879084,I2683,I591962,I592189,);
nor I_34675 (I592197,I592189,I592056);
not I_34676 (I592214,I592197);
not I_34677 (I592231,I592189);
nor I_34678 (I592248,I592231,I592132);
DFFARX1 I_34679 (I592248,I2683,I591962,I591948,);
nand I_34680 (I592279,I879063,I879063);
and I_34681 (I592296,I592279,I879060);
DFFARX1 I_34682 (I592296,I2683,I591962,I592322,);
nor I_34683 (I592330,I592322,I592189);
DFFARX1 I_34684 (I592330,I2683,I591962,I591930,);
nand I_34685 (I592361,I592322,I592231);
nand I_34686 (I591939,I592214,I592361);
not I_34687 (I592392,I592322);
nor I_34688 (I592409,I592392,I592132);
DFFARX1 I_34689 (I592409,I2683,I591962,I591951,);
nor I_34690 (I592440,I879081,I879063);
or I_34691 (I591942,I592189,I592440);
nor I_34692 (I591933,I592322,I592440);
or I_34693 (I591936,I592056,I592440);
DFFARX1 I_34694 (I592440,I2683,I591962,I591954,);
not I_34695 (I592540,I2690);
DFFARX1 I_34696 (I282809,I2683,I592540,I592566,);
not I_34697 (I592574,I592566);
nand I_34698 (I592591,I282812,I282788);
and I_34699 (I592608,I592591,I282785);
DFFARX1 I_34700 (I592608,I2683,I592540,I592634,);
not I_34701 (I592642,I282791);
DFFARX1 I_34702 (I282785,I2683,I592540,I592668,);
not I_34703 (I592676,I592668);
nor I_34704 (I592693,I592676,I592574);
and I_34705 (I592710,I592693,I282791);
nor I_34706 (I592727,I592676,I592642);
nor I_34707 (I592523,I592634,I592727);
DFFARX1 I_34708 (I282794,I2683,I592540,I592767,);
nor I_34709 (I592775,I592767,I592634);
not I_34710 (I592792,I592775);
not I_34711 (I592809,I592767);
nor I_34712 (I592826,I592809,I592710);
DFFARX1 I_34713 (I592826,I2683,I592540,I592526,);
nand I_34714 (I592857,I282797,I282806);
and I_34715 (I592874,I592857,I282803);
DFFARX1 I_34716 (I592874,I2683,I592540,I592900,);
nor I_34717 (I592908,I592900,I592767);
DFFARX1 I_34718 (I592908,I2683,I592540,I592508,);
nand I_34719 (I592939,I592900,I592809);
nand I_34720 (I592517,I592792,I592939);
not I_34721 (I592970,I592900);
nor I_34722 (I592987,I592970,I592710);
DFFARX1 I_34723 (I592987,I2683,I592540,I592529,);
nor I_34724 (I593018,I282800,I282806);
or I_34725 (I592520,I592767,I593018);
nor I_34726 (I592511,I592900,I593018);
or I_34727 (I592514,I592634,I593018);
DFFARX1 I_34728 (I593018,I2683,I592540,I592532,);
not I_34729 (I593118,I2690);
DFFARX1 I_34730 (I441650,I2683,I593118,I593144,);
not I_34731 (I593152,I593144);
nand I_34732 (I593169,I441659,I441668);
and I_34733 (I593186,I593169,I441674);
DFFARX1 I_34734 (I593186,I2683,I593118,I593212,);
not I_34735 (I593220,I441671);
DFFARX1 I_34736 (I441656,I2683,I593118,I593246,);
not I_34737 (I593254,I593246);
nor I_34738 (I593271,I593254,I593152);
and I_34739 (I593288,I593271,I441671);
nor I_34740 (I593305,I593254,I593220);
nor I_34741 (I593101,I593212,I593305);
DFFARX1 I_34742 (I441665,I2683,I593118,I593345,);
nor I_34743 (I593353,I593345,I593212);
not I_34744 (I593370,I593353);
not I_34745 (I593387,I593345);
nor I_34746 (I593404,I593387,I593288);
DFFARX1 I_34747 (I593404,I2683,I593118,I593104,);
nand I_34748 (I593435,I441662,I441653);
and I_34749 (I593452,I593435,I441650);
DFFARX1 I_34750 (I593452,I2683,I593118,I593478,);
nor I_34751 (I593486,I593478,I593345);
DFFARX1 I_34752 (I593486,I2683,I593118,I593086,);
nand I_34753 (I593517,I593478,I593387);
nand I_34754 (I593095,I593370,I593517);
not I_34755 (I593548,I593478);
nor I_34756 (I593565,I593548,I593288);
DFFARX1 I_34757 (I593565,I2683,I593118,I593107,);
nor I_34758 (I593596,I441653,I441653);
or I_34759 (I593098,I593345,I593596);
nor I_34760 (I593089,I593478,I593596);
or I_34761 (I593092,I593212,I593596);
DFFARX1 I_34762 (I593596,I2683,I593118,I593110,);
not I_34763 (I593696,I2690);
DFFARX1 I_34764 (I990308,I2683,I593696,I593722,);
not I_34765 (I593730,I593722);
nand I_34766 (I593747,I990332,I990314);
and I_34767 (I593764,I593747,I990320);
DFFARX1 I_34768 (I593764,I2683,I593696,I593790,);
not I_34769 (I593798,I990326);
DFFARX1 I_34770 (I990311,I2683,I593696,I593824,);
not I_34771 (I593832,I593824);
nor I_34772 (I593849,I593832,I593730);
and I_34773 (I593866,I593849,I990326);
nor I_34774 (I593883,I593832,I593798);
nor I_34775 (I593679,I593790,I593883);
DFFARX1 I_34776 (I990323,I2683,I593696,I593923,);
nor I_34777 (I593931,I593923,I593790);
not I_34778 (I593948,I593931);
not I_34779 (I593965,I593923);
nor I_34780 (I593982,I593965,I593866);
DFFARX1 I_34781 (I593982,I2683,I593696,I593682,);
nand I_34782 (I594013,I990329,I990317);
and I_34783 (I594030,I594013,I990311);
DFFARX1 I_34784 (I594030,I2683,I593696,I594056,);
nor I_34785 (I594064,I594056,I593923);
DFFARX1 I_34786 (I594064,I2683,I593696,I593664,);
nand I_34787 (I594095,I594056,I593965);
nand I_34788 (I593673,I593948,I594095);
not I_34789 (I594126,I594056);
nor I_34790 (I594143,I594126,I593866);
DFFARX1 I_34791 (I594143,I2683,I593696,I593685,);
nor I_34792 (I594174,I990308,I990317);
or I_34793 (I593676,I593923,I594174);
nor I_34794 (I593667,I594056,I594174);
or I_34795 (I593670,I593790,I594174);
DFFARX1 I_34796 (I594174,I2683,I593696,I593688,);
not I_34797 (I594274,I2690);
DFFARX1 I_34798 (I40615,I2683,I594274,I594300,);
not I_34799 (I594308,I594300);
nand I_34800 (I594325,I40612,I40603);
and I_34801 (I594342,I594325,I40603);
DFFARX1 I_34802 (I594342,I2683,I594274,I594368,);
not I_34803 (I594376,I40606);
DFFARX1 I_34804 (I40621,I2683,I594274,I594402,);
not I_34805 (I594410,I594402);
nor I_34806 (I594427,I594410,I594308);
and I_34807 (I594444,I594427,I40606);
nor I_34808 (I594461,I594410,I594376);
nor I_34809 (I594257,I594368,I594461);
DFFARX1 I_34810 (I40606,I2683,I594274,I594501,);
nor I_34811 (I594509,I594501,I594368);
not I_34812 (I594526,I594509);
not I_34813 (I594543,I594501);
nor I_34814 (I594560,I594543,I594444);
DFFARX1 I_34815 (I594560,I2683,I594274,I594260,);
nand I_34816 (I594591,I40624,I40609);
and I_34817 (I594608,I594591,I40627);
DFFARX1 I_34818 (I594608,I2683,I594274,I594634,);
nor I_34819 (I594642,I594634,I594501);
DFFARX1 I_34820 (I594642,I2683,I594274,I594242,);
nand I_34821 (I594673,I594634,I594543);
nand I_34822 (I594251,I594526,I594673);
not I_34823 (I594704,I594634);
nor I_34824 (I594721,I594704,I594444);
DFFARX1 I_34825 (I594721,I2683,I594274,I594263,);
nor I_34826 (I594752,I40618,I40609);
or I_34827 (I594254,I594501,I594752);
nor I_34828 (I594245,I594634,I594752);
or I_34829 (I594248,I594368,I594752);
DFFARX1 I_34830 (I594752,I2683,I594274,I594266,);
not I_34831 (I594852,I2690);
DFFARX1 I_34832 (I272269,I2683,I594852,I594878,);
not I_34833 (I594886,I594878);
nand I_34834 (I594903,I272272,I272248);
and I_34835 (I594920,I594903,I272245);
DFFARX1 I_34836 (I594920,I2683,I594852,I594946,);
not I_34837 (I594954,I272251);
DFFARX1 I_34838 (I272245,I2683,I594852,I594980,);
not I_34839 (I594988,I594980);
nor I_34840 (I595005,I594988,I594886);
and I_34841 (I595022,I595005,I272251);
nor I_34842 (I595039,I594988,I594954);
nor I_34843 (I594835,I594946,I595039);
DFFARX1 I_34844 (I272254,I2683,I594852,I595079,);
nor I_34845 (I595087,I595079,I594946);
not I_34846 (I595104,I595087);
not I_34847 (I595121,I595079);
nor I_34848 (I595138,I595121,I595022);
DFFARX1 I_34849 (I595138,I2683,I594852,I594838,);
nand I_34850 (I595169,I272257,I272266);
and I_34851 (I595186,I595169,I272263);
DFFARX1 I_34852 (I595186,I2683,I594852,I595212,);
nor I_34853 (I595220,I595212,I595079);
DFFARX1 I_34854 (I595220,I2683,I594852,I594820,);
nand I_34855 (I595251,I595212,I595121);
nand I_34856 (I594829,I595104,I595251);
not I_34857 (I595282,I595212);
nor I_34858 (I595299,I595282,I595022);
DFFARX1 I_34859 (I595299,I2683,I594852,I594841,);
nor I_34860 (I595330,I272260,I272266);
or I_34861 (I594832,I595079,I595330);
nor I_34862 (I594823,I595212,I595330);
or I_34863 (I594826,I594946,I595330);
DFFARX1 I_34864 (I595330,I2683,I594852,I594844,);
not I_34865 (I595430,I2690);
DFFARX1 I_34866 (I384539,I2683,I595430,I595456,);
not I_34867 (I595464,I595456);
nand I_34868 (I595481,I384530,I384548);
and I_34869 (I595498,I595481,I384551);
DFFARX1 I_34870 (I595498,I2683,I595430,I595524,);
not I_34871 (I595532,I384545);
DFFARX1 I_34872 (I384533,I2683,I595430,I595558,);
not I_34873 (I595566,I595558);
nor I_34874 (I595583,I595566,I595464);
and I_34875 (I595600,I595583,I384545);
nor I_34876 (I595617,I595566,I595532);
nor I_34877 (I595413,I595524,I595617);
DFFARX1 I_34878 (I384542,I2683,I595430,I595657,);
nor I_34879 (I595665,I595657,I595524);
not I_34880 (I595682,I595665);
not I_34881 (I595699,I595657);
nor I_34882 (I595716,I595699,I595600);
DFFARX1 I_34883 (I595716,I2683,I595430,I595416,);
nand I_34884 (I595747,I384557,I384554);
and I_34885 (I595764,I595747,I384536);
DFFARX1 I_34886 (I595764,I2683,I595430,I595790,);
nor I_34887 (I595798,I595790,I595657);
DFFARX1 I_34888 (I595798,I2683,I595430,I595398,);
nand I_34889 (I595829,I595790,I595699);
nand I_34890 (I595407,I595682,I595829);
not I_34891 (I595860,I595790);
nor I_34892 (I595877,I595860,I595600);
DFFARX1 I_34893 (I595877,I2683,I595430,I595419,);
nor I_34894 (I595908,I384530,I384554);
or I_34895 (I595410,I595657,I595908);
nor I_34896 (I595401,I595790,I595908);
or I_34897 (I595404,I595524,I595908);
DFFARX1 I_34898 (I595908,I2683,I595430,I595422,);
not I_34899 (I596008,I2690);
DFFARX1 I_34900 (I648623,I2683,I596008,I596034,);
not I_34901 (I596042,I596034);
nand I_34902 (I596059,I648611,I648629);
and I_34903 (I596076,I596059,I648626);
DFFARX1 I_34904 (I596076,I2683,I596008,I596102,);
not I_34905 (I596110,I648617);
DFFARX1 I_34906 (I648614,I2683,I596008,I596136,);
not I_34907 (I596144,I596136);
nor I_34908 (I596161,I596144,I596042);
and I_34909 (I596178,I596161,I648617);
nor I_34910 (I596195,I596144,I596110);
nor I_34911 (I595991,I596102,I596195);
DFFARX1 I_34912 (I648608,I2683,I596008,I596235,);
nor I_34913 (I596243,I596235,I596102);
not I_34914 (I596260,I596243);
not I_34915 (I596277,I596235);
nor I_34916 (I596294,I596277,I596178);
DFFARX1 I_34917 (I596294,I2683,I596008,I595994,);
nand I_34918 (I596325,I648608,I648611);
and I_34919 (I596342,I596325,I648614);
DFFARX1 I_34920 (I596342,I2683,I596008,I596368,);
nor I_34921 (I596376,I596368,I596235);
DFFARX1 I_34922 (I596376,I2683,I596008,I595976,);
nand I_34923 (I596407,I596368,I596277);
nand I_34924 (I595985,I596260,I596407);
not I_34925 (I596438,I596368);
nor I_34926 (I596455,I596438,I596178);
DFFARX1 I_34927 (I596455,I2683,I596008,I595997,);
nor I_34928 (I596486,I648620,I648611);
or I_34929 (I595988,I596235,I596486);
nor I_34930 (I595979,I596368,I596486);
or I_34931 (I595982,I596102,I596486);
DFFARX1 I_34932 (I596486,I2683,I596008,I596000,);
not I_34933 (I596586,I2690);
DFFARX1 I_34934 (I70118,I2683,I596586,I596612,);
not I_34935 (I596620,I596612);
nand I_34936 (I596637,I70127,I70136);
and I_34937 (I596654,I596637,I70115);
DFFARX1 I_34938 (I596654,I2683,I596586,I596680,);
not I_34939 (I596688,I70118);
DFFARX1 I_34940 (I70133,I2683,I596586,I596714,);
not I_34941 (I596722,I596714);
nor I_34942 (I596739,I596722,I596620);
and I_34943 (I596756,I596739,I70118);
nor I_34944 (I596773,I596722,I596688);
nor I_34945 (I596569,I596680,I596773);
DFFARX1 I_34946 (I70124,I2683,I596586,I596813,);
nor I_34947 (I596821,I596813,I596680);
not I_34948 (I596838,I596821);
not I_34949 (I596855,I596813);
nor I_34950 (I596872,I596855,I596756);
DFFARX1 I_34951 (I596872,I2683,I596586,I596572,);
nand I_34952 (I596903,I70139,I70115);
and I_34953 (I596920,I596903,I70121);
DFFARX1 I_34954 (I596920,I2683,I596586,I596946,);
nor I_34955 (I596954,I596946,I596813);
DFFARX1 I_34956 (I596954,I2683,I596586,I596554,);
nand I_34957 (I596985,I596946,I596855);
nand I_34958 (I596563,I596838,I596985);
not I_34959 (I597016,I596946);
nor I_34960 (I597033,I597016,I596756);
DFFARX1 I_34961 (I597033,I2683,I596586,I596575,);
nor I_34962 (I597064,I70130,I70115);
or I_34963 (I596566,I596813,I597064);
nor I_34964 (I596557,I596946,I597064);
or I_34965 (I596560,I596680,I597064);
DFFARX1 I_34966 (I597064,I2683,I596586,I596578,);
not I_34967 (I597164,I2690);
DFFARX1 I_34968 (I683932,I2683,I597164,I597190,);
not I_34969 (I597198,I597190);
nand I_34970 (I597215,I683920,I683938);
and I_34971 (I597232,I597215,I683935);
DFFARX1 I_34972 (I597232,I2683,I597164,I597258,);
not I_34973 (I597266,I683926);
DFFARX1 I_34974 (I683923,I2683,I597164,I597292,);
not I_34975 (I597300,I597292);
nor I_34976 (I597317,I597300,I597198);
and I_34977 (I597334,I597317,I683926);
nor I_34978 (I597351,I597300,I597266);
nor I_34979 (I597147,I597258,I597351);
DFFARX1 I_34980 (I683917,I2683,I597164,I597391,);
nor I_34981 (I597399,I597391,I597258);
not I_34982 (I597416,I597399);
not I_34983 (I597433,I597391);
nor I_34984 (I597450,I597433,I597334);
DFFARX1 I_34985 (I597450,I2683,I597164,I597150,);
nand I_34986 (I597481,I683917,I683920);
and I_34987 (I597498,I597481,I683923);
DFFARX1 I_34988 (I597498,I2683,I597164,I597524,);
nor I_34989 (I597532,I597524,I597391);
DFFARX1 I_34990 (I597532,I2683,I597164,I597132,);
nand I_34991 (I597563,I597524,I597433);
nand I_34992 (I597141,I597416,I597563);
not I_34993 (I597594,I597524);
nor I_34994 (I597611,I597594,I597334);
DFFARX1 I_34995 (I597611,I2683,I597164,I597153,);
nor I_34996 (I597642,I683929,I683920);
or I_34997 (I597144,I597391,I597642);
nor I_34998 (I597135,I597524,I597642);
or I_34999 (I597138,I597258,I597642);
DFFARX1 I_35000 (I597642,I2683,I597164,I597156,);
not I_35001 (I597742,I2690);
DFFARX1 I_35002 (I835728,I2683,I597742,I597768,);
not I_35003 (I597776,I597768);
nand I_35004 (I597793,I835710,I835722);
and I_35005 (I597810,I597793,I835725);
DFFARX1 I_35006 (I597810,I2683,I597742,I597836,);
not I_35007 (I597844,I835719);
DFFARX1 I_35008 (I835716,I2683,I597742,I597870,);
not I_35009 (I597878,I597870);
nor I_35010 (I597895,I597878,I597776);
and I_35011 (I597912,I597895,I835719);
nor I_35012 (I597929,I597878,I597844);
nor I_35013 (I597725,I597836,I597929);
DFFARX1 I_35014 (I835734,I2683,I597742,I597969,);
nor I_35015 (I597977,I597969,I597836);
not I_35016 (I597994,I597977);
not I_35017 (I598011,I597969);
nor I_35018 (I598028,I598011,I597912);
DFFARX1 I_35019 (I598028,I2683,I597742,I597728,);
nand I_35020 (I598059,I835713,I835713);
and I_35021 (I598076,I598059,I835710);
DFFARX1 I_35022 (I598076,I2683,I597742,I598102,);
nor I_35023 (I598110,I598102,I597969);
DFFARX1 I_35024 (I598110,I2683,I597742,I597710,);
nand I_35025 (I598141,I598102,I598011);
nand I_35026 (I597719,I597994,I598141);
not I_35027 (I598172,I598102);
nor I_35028 (I598189,I598172,I597912);
DFFARX1 I_35029 (I598189,I2683,I597742,I597731,);
nor I_35030 (I598220,I835731,I835713);
or I_35031 (I597722,I597969,I598220);
nor I_35032 (I597713,I598102,I598220);
or I_35033 (I597716,I597836,I598220);
DFFARX1 I_35034 (I598220,I2683,I597742,I597734,);
not I_35035 (I598320,I2690);
DFFARX1 I_35036 (I358427,I2683,I598320,I598346,);
not I_35037 (I598354,I598346);
nand I_35038 (I598371,I358418,I358436);
and I_35039 (I598388,I598371,I358439);
DFFARX1 I_35040 (I598388,I2683,I598320,I598414,);
not I_35041 (I598422,I358433);
DFFARX1 I_35042 (I358421,I2683,I598320,I598448,);
not I_35043 (I598456,I598448);
nor I_35044 (I598473,I598456,I598354);
and I_35045 (I598490,I598473,I358433);
nor I_35046 (I598507,I598456,I598422);
nor I_35047 (I598303,I598414,I598507);
DFFARX1 I_35048 (I358430,I2683,I598320,I598547,);
nor I_35049 (I598555,I598547,I598414);
not I_35050 (I598572,I598555);
not I_35051 (I598589,I598547);
nor I_35052 (I598606,I598589,I598490);
DFFARX1 I_35053 (I598606,I2683,I598320,I598306,);
nand I_35054 (I598637,I358445,I358442);
and I_35055 (I598654,I598637,I358424);
DFFARX1 I_35056 (I598654,I2683,I598320,I598680,);
nor I_35057 (I598688,I598680,I598547);
DFFARX1 I_35058 (I598688,I2683,I598320,I598288,);
nand I_35059 (I598719,I598680,I598589);
nand I_35060 (I598297,I598572,I598719);
not I_35061 (I598750,I598680);
nor I_35062 (I598767,I598750,I598490);
DFFARX1 I_35063 (I598767,I2683,I598320,I598309,);
nor I_35064 (I598798,I358418,I358442);
or I_35065 (I598300,I598547,I598798);
nor I_35066 (I598291,I598680,I598798);
or I_35067 (I598294,I598414,I598798);
DFFARX1 I_35068 (I598798,I2683,I598320,I598312,);
not I_35069 (I598898,I2690);
DFFARX1 I_35070 (I50092,I2683,I598898,I598924,);
not I_35071 (I598932,I598924);
nand I_35072 (I598949,I50101,I50110);
and I_35073 (I598966,I598949,I50089);
DFFARX1 I_35074 (I598966,I2683,I598898,I598992,);
not I_35075 (I599000,I50092);
DFFARX1 I_35076 (I50107,I2683,I598898,I599026,);
not I_35077 (I599034,I599026);
nor I_35078 (I599051,I599034,I598932);
and I_35079 (I599068,I599051,I50092);
nor I_35080 (I599085,I599034,I599000);
nor I_35081 (I598881,I598992,I599085);
DFFARX1 I_35082 (I50098,I2683,I598898,I599125,);
nor I_35083 (I599133,I599125,I598992);
not I_35084 (I599150,I599133);
not I_35085 (I599167,I599125);
nor I_35086 (I599184,I599167,I599068);
DFFARX1 I_35087 (I599184,I2683,I598898,I598884,);
nand I_35088 (I599215,I50113,I50089);
and I_35089 (I599232,I599215,I50095);
DFFARX1 I_35090 (I599232,I2683,I598898,I599258,);
nor I_35091 (I599266,I599258,I599125);
DFFARX1 I_35092 (I599266,I2683,I598898,I598866,);
nand I_35093 (I599297,I599258,I599167);
nand I_35094 (I598875,I599150,I599297);
not I_35095 (I599328,I599258);
nor I_35096 (I599345,I599328,I599068);
DFFARX1 I_35097 (I599345,I2683,I598898,I598887,);
nor I_35098 (I599376,I50104,I50089);
or I_35099 (I598878,I599125,I599376);
nor I_35100 (I598869,I599258,I599376);
or I_35101 (I598872,I598992,I599376);
DFFARX1 I_35102 (I599376,I2683,I598898,I598890,);
not I_35103 (I599476,I2690);
DFFARX1 I_35104 (I107008,I2683,I599476,I599502,);
not I_35105 (I599510,I599502);
nand I_35106 (I599527,I107017,I107026);
and I_35107 (I599544,I599527,I107005);
DFFARX1 I_35108 (I599544,I2683,I599476,I599570,);
not I_35109 (I599578,I107008);
DFFARX1 I_35110 (I107023,I2683,I599476,I599604,);
not I_35111 (I599612,I599604);
nor I_35112 (I599629,I599612,I599510);
and I_35113 (I599646,I599629,I107008);
nor I_35114 (I599663,I599612,I599578);
nor I_35115 (I599459,I599570,I599663);
DFFARX1 I_35116 (I107014,I2683,I599476,I599703,);
nor I_35117 (I599711,I599703,I599570);
not I_35118 (I599728,I599711);
not I_35119 (I599745,I599703);
nor I_35120 (I599762,I599745,I599646);
DFFARX1 I_35121 (I599762,I2683,I599476,I599462,);
nand I_35122 (I599793,I107029,I107005);
and I_35123 (I599810,I599793,I107011);
DFFARX1 I_35124 (I599810,I2683,I599476,I599836,);
nor I_35125 (I599844,I599836,I599703);
DFFARX1 I_35126 (I599844,I2683,I599476,I599444,);
nand I_35127 (I599875,I599836,I599745);
nand I_35128 (I599453,I599728,I599875);
not I_35129 (I599906,I599836);
nor I_35130 (I599923,I599906,I599646);
DFFARX1 I_35131 (I599923,I2683,I599476,I599465,);
nor I_35132 (I599954,I107020,I107005);
or I_35133 (I599456,I599703,I599954);
nor I_35134 (I599447,I599836,I599954);
or I_35135 (I599450,I599570,I599954);
DFFARX1 I_35136 (I599954,I2683,I599476,I599468,);
not I_35137 (I600054,I2690);
DFFARX1 I_35138 (I242757,I2683,I600054,I600080,);
not I_35139 (I600088,I600080);
nand I_35140 (I600105,I242760,I242736);
and I_35141 (I600122,I600105,I242733);
DFFARX1 I_35142 (I600122,I2683,I600054,I600148,);
not I_35143 (I600156,I242739);
DFFARX1 I_35144 (I242733,I2683,I600054,I600182,);
not I_35145 (I600190,I600182);
nor I_35146 (I600207,I600190,I600088);
and I_35147 (I600224,I600207,I242739);
nor I_35148 (I600241,I600190,I600156);
nor I_35149 (I600037,I600148,I600241);
DFFARX1 I_35150 (I242742,I2683,I600054,I600281,);
nor I_35151 (I600289,I600281,I600148);
not I_35152 (I600306,I600289);
not I_35153 (I600323,I600281);
nor I_35154 (I600340,I600323,I600224);
DFFARX1 I_35155 (I600340,I2683,I600054,I600040,);
nand I_35156 (I600371,I242745,I242754);
and I_35157 (I600388,I600371,I242751);
DFFARX1 I_35158 (I600388,I2683,I600054,I600414,);
nor I_35159 (I600422,I600414,I600281);
DFFARX1 I_35160 (I600422,I2683,I600054,I600022,);
nand I_35161 (I600453,I600414,I600323);
nand I_35162 (I600031,I600306,I600453);
not I_35163 (I600484,I600414);
nor I_35164 (I600501,I600484,I600224);
DFFARX1 I_35165 (I600501,I2683,I600054,I600043,);
nor I_35166 (I600532,I242748,I242754);
or I_35167 (I600034,I600281,I600532);
nor I_35168 (I600025,I600414,I600532);
or I_35169 (I600028,I600148,I600532);
DFFARX1 I_35170 (I600532,I2683,I600054,I600046,);
not I_35171 (I600632,I2690);
DFFARX1 I_35172 (I731643,I2683,I600632,I600658,);
not I_35173 (I600666,I600658);
nand I_35174 (I600683,I731619,I731634);
and I_35175 (I600700,I600683,I731646);
DFFARX1 I_35176 (I600700,I2683,I600632,I600726,);
not I_35177 (I600734,I731631);
DFFARX1 I_35178 (I731622,I2683,I600632,I600760,);
not I_35179 (I600768,I600760);
nor I_35180 (I600785,I600768,I600666);
and I_35181 (I600802,I600785,I731631);
nor I_35182 (I600819,I600768,I600734);
nor I_35183 (I600615,I600726,I600819);
DFFARX1 I_35184 (I731619,I2683,I600632,I600859,);
nor I_35185 (I600867,I600859,I600726);
not I_35186 (I600884,I600867);
not I_35187 (I600901,I600859);
nor I_35188 (I600918,I600901,I600802);
DFFARX1 I_35189 (I600918,I2683,I600632,I600618,);
nand I_35190 (I600949,I731637,I731628);
and I_35191 (I600966,I600949,I731640);
DFFARX1 I_35192 (I600966,I2683,I600632,I600992,);
nor I_35193 (I601000,I600992,I600859);
DFFARX1 I_35194 (I601000,I2683,I600632,I600600,);
nand I_35195 (I601031,I600992,I600901);
nand I_35196 (I600609,I600884,I601031);
not I_35197 (I601062,I600992);
nor I_35198 (I601079,I601062,I600802);
DFFARX1 I_35199 (I601079,I2683,I600632,I600621,);
nor I_35200 (I601110,I731625,I731628);
or I_35201 (I600612,I600859,I601110);
nor I_35202 (I600603,I600992,I601110);
or I_35203 (I600606,I600726,I601110);
DFFARX1 I_35204 (I601110,I2683,I600632,I600624,);
not I_35205 (I601210,I2690);
DFFARX1 I_35206 (I453210,I2683,I601210,I601236,);
not I_35207 (I601244,I601236);
nand I_35208 (I601261,I453219,I453228);
and I_35209 (I601278,I601261,I453234);
DFFARX1 I_35210 (I601278,I2683,I601210,I601304,);
not I_35211 (I601312,I453231);
DFFARX1 I_35212 (I453216,I2683,I601210,I601338,);
not I_35213 (I601346,I601338);
nor I_35214 (I601363,I601346,I601244);
and I_35215 (I601380,I601363,I453231);
nor I_35216 (I601397,I601346,I601312);
nor I_35217 (I601193,I601304,I601397);
DFFARX1 I_35218 (I453225,I2683,I601210,I601437,);
nor I_35219 (I601445,I601437,I601304);
not I_35220 (I601462,I601445);
not I_35221 (I601479,I601437);
nor I_35222 (I601496,I601479,I601380);
DFFARX1 I_35223 (I601496,I2683,I601210,I601196,);
nand I_35224 (I601527,I453222,I453213);
and I_35225 (I601544,I601527,I453210);
DFFARX1 I_35226 (I601544,I2683,I601210,I601570,);
nor I_35227 (I601578,I601570,I601437);
DFFARX1 I_35228 (I601578,I2683,I601210,I601178,);
nand I_35229 (I601609,I601570,I601479);
nand I_35230 (I601187,I601462,I601609);
not I_35231 (I601640,I601570);
nor I_35232 (I601657,I601640,I601380);
DFFARX1 I_35233 (I601657,I2683,I601210,I601199,);
nor I_35234 (I601688,I453213,I453213);
or I_35235 (I601190,I601437,I601688);
nor I_35236 (I601181,I601570,I601688);
or I_35237 (I601184,I601304,I601688);
DFFARX1 I_35238 (I601688,I2683,I601210,I601202,);
not I_35239 (I601788,I2690);
DFFARX1 I_35240 (I419907,I2683,I601788,I601814,);
not I_35241 (I601822,I601814);
nand I_35242 (I601839,I419922,I419907);
and I_35243 (I601856,I601839,I419910);
DFFARX1 I_35244 (I601856,I2683,I601788,I601882,);
not I_35245 (I601890,I419910);
DFFARX1 I_35246 (I419919,I2683,I601788,I601916,);
not I_35247 (I601924,I601916);
nor I_35248 (I601941,I601924,I601822);
and I_35249 (I601958,I601941,I419910);
nor I_35250 (I601975,I601924,I601890);
nor I_35251 (I601771,I601882,I601975);
DFFARX1 I_35252 (I419913,I2683,I601788,I602015,);
nor I_35253 (I602023,I602015,I601882);
not I_35254 (I602040,I602023);
not I_35255 (I602057,I602015);
nor I_35256 (I602074,I602057,I601958);
DFFARX1 I_35257 (I602074,I2683,I601788,I601774,);
nand I_35258 (I602105,I419916,I419925);
and I_35259 (I602122,I602105,I419931);
DFFARX1 I_35260 (I602122,I2683,I601788,I602148,);
nor I_35261 (I602156,I602148,I602015);
DFFARX1 I_35262 (I602156,I2683,I601788,I601756,);
nand I_35263 (I602187,I602148,I602057);
nand I_35264 (I601765,I602040,I602187);
not I_35265 (I602218,I602148);
nor I_35266 (I602235,I602218,I601958);
DFFARX1 I_35267 (I602235,I2683,I601788,I601777,);
nor I_35268 (I602266,I419928,I419925);
or I_35269 (I601768,I602015,I602266);
nor I_35270 (I601759,I602148,I602266);
or I_35271 (I601762,I601882,I602266);
DFFARX1 I_35272 (I602266,I2683,I601788,I601780,);
not I_35273 (I602366,I2690);
DFFARX1 I_35274 (I374203,I2683,I602366,I602392,);
not I_35275 (I602400,I602392);
nand I_35276 (I602417,I374194,I374212);
and I_35277 (I602434,I602417,I374215);
DFFARX1 I_35278 (I602434,I2683,I602366,I602460,);
not I_35279 (I602468,I374209);
DFFARX1 I_35280 (I374197,I2683,I602366,I602494,);
not I_35281 (I602502,I602494);
nor I_35282 (I602519,I602502,I602400);
and I_35283 (I602536,I602519,I374209);
nor I_35284 (I602553,I602502,I602468);
nor I_35285 (I602349,I602460,I602553);
DFFARX1 I_35286 (I374206,I2683,I602366,I602593,);
nor I_35287 (I602601,I602593,I602460);
not I_35288 (I602618,I602601);
not I_35289 (I602635,I602593);
nor I_35290 (I602652,I602635,I602536);
DFFARX1 I_35291 (I602652,I2683,I602366,I602352,);
nand I_35292 (I602683,I374221,I374218);
and I_35293 (I602700,I602683,I374200);
DFFARX1 I_35294 (I602700,I2683,I602366,I602726,);
nor I_35295 (I602734,I602726,I602593);
DFFARX1 I_35296 (I602734,I2683,I602366,I602334,);
nand I_35297 (I602765,I602726,I602635);
nand I_35298 (I602343,I602618,I602765);
not I_35299 (I602796,I602726);
nor I_35300 (I602813,I602796,I602536);
DFFARX1 I_35301 (I602813,I2683,I602366,I602355,);
nor I_35302 (I602844,I374194,I374218);
or I_35303 (I602346,I602593,I602844);
nor I_35304 (I602337,I602726,I602844);
or I_35305 (I602340,I602460,I602844);
DFFARX1 I_35306 (I602844,I2683,I602366,I602358,);
not I_35307 (I602944,I2690);
DFFARX1 I_35308 (I783323,I2683,I602944,I602970,);
not I_35309 (I602978,I602970);
nand I_35310 (I602995,I783299,I783314);
and I_35311 (I603012,I602995,I783326);
DFFARX1 I_35312 (I603012,I2683,I602944,I603038,);
not I_35313 (I603046,I783311);
DFFARX1 I_35314 (I783302,I2683,I602944,I603072,);
not I_35315 (I603080,I603072);
nor I_35316 (I603097,I603080,I602978);
and I_35317 (I603114,I603097,I783311);
nor I_35318 (I603131,I603080,I603046);
nor I_35319 (I602927,I603038,I603131);
DFFARX1 I_35320 (I783299,I2683,I602944,I603171,);
nor I_35321 (I603179,I603171,I603038);
not I_35322 (I603196,I603179);
not I_35323 (I603213,I603171);
nor I_35324 (I603230,I603213,I603114);
DFFARX1 I_35325 (I603230,I2683,I602944,I602930,);
nand I_35326 (I603261,I783317,I783308);
and I_35327 (I603278,I603261,I783320);
DFFARX1 I_35328 (I603278,I2683,I602944,I603304,);
nor I_35329 (I603312,I603304,I603171);
DFFARX1 I_35330 (I603312,I2683,I602944,I602912,);
nand I_35331 (I603343,I603304,I603213);
nand I_35332 (I602921,I603196,I603343);
not I_35333 (I603374,I603304);
nor I_35334 (I603391,I603374,I603114);
DFFARX1 I_35335 (I603391,I2683,I602944,I602933,);
nor I_35336 (I603422,I783305,I783308);
or I_35337 (I602924,I603171,I603422);
nor I_35338 (I602915,I603304,I603422);
or I_35339 (I602918,I603038,I603422);
DFFARX1 I_35340 (I603422,I2683,I602944,I602936,);
not I_35341 (I603522,I2690);
DFFARX1 I_35342 (I81185,I2683,I603522,I603548,);
not I_35343 (I603556,I603548);
nand I_35344 (I603573,I81194,I81203);
and I_35345 (I603590,I603573,I81182);
DFFARX1 I_35346 (I603590,I2683,I603522,I603616,);
not I_35347 (I603624,I81185);
DFFARX1 I_35348 (I81200,I2683,I603522,I603650,);
not I_35349 (I603658,I603650);
nor I_35350 (I603675,I603658,I603556);
and I_35351 (I603692,I603675,I81185);
nor I_35352 (I603709,I603658,I603624);
nor I_35353 (I603505,I603616,I603709);
DFFARX1 I_35354 (I81191,I2683,I603522,I603749,);
nor I_35355 (I603757,I603749,I603616);
not I_35356 (I603774,I603757);
not I_35357 (I603791,I603749);
nor I_35358 (I603808,I603791,I603692);
DFFARX1 I_35359 (I603808,I2683,I603522,I603508,);
nand I_35360 (I603839,I81206,I81182);
and I_35361 (I603856,I603839,I81188);
DFFARX1 I_35362 (I603856,I2683,I603522,I603882,);
nor I_35363 (I603890,I603882,I603749);
DFFARX1 I_35364 (I603890,I2683,I603522,I603490,);
nand I_35365 (I603921,I603882,I603791);
nand I_35366 (I603499,I603774,I603921);
not I_35367 (I603952,I603882);
nor I_35368 (I603969,I603952,I603692);
DFFARX1 I_35369 (I603969,I2683,I603522,I603511,);
nor I_35370 (I604000,I81197,I81182);
or I_35371 (I603502,I603749,I604000);
nor I_35372 (I603493,I603882,I604000);
or I_35373 (I603496,I603616,I604000);
DFFARX1 I_35374 (I604000,I2683,I603522,I603514,);
not I_35375 (I604100,I2690);
DFFARX1 I_35376 (I747147,I2683,I604100,I604126,);
not I_35377 (I604134,I604126);
nand I_35378 (I604151,I747123,I747138);
and I_35379 (I604168,I604151,I747150);
DFFARX1 I_35380 (I604168,I2683,I604100,I604194,);
not I_35381 (I604202,I747135);
DFFARX1 I_35382 (I747126,I2683,I604100,I604228,);
not I_35383 (I604236,I604228);
nor I_35384 (I604253,I604236,I604134);
and I_35385 (I604270,I604253,I747135);
nor I_35386 (I604287,I604236,I604202);
nor I_35387 (I604083,I604194,I604287);
DFFARX1 I_35388 (I747123,I2683,I604100,I604327,);
nor I_35389 (I604335,I604327,I604194);
not I_35390 (I604352,I604335);
not I_35391 (I604369,I604327);
nor I_35392 (I604386,I604369,I604270);
DFFARX1 I_35393 (I604386,I2683,I604100,I604086,);
nand I_35394 (I604417,I747141,I747132);
and I_35395 (I604434,I604417,I747144);
DFFARX1 I_35396 (I604434,I2683,I604100,I604460,);
nor I_35397 (I604468,I604460,I604327);
DFFARX1 I_35398 (I604468,I2683,I604100,I604068,);
nand I_35399 (I604499,I604460,I604369);
nand I_35400 (I604077,I604352,I604499);
not I_35401 (I604530,I604460);
nor I_35402 (I604547,I604530,I604270);
DFFARX1 I_35403 (I604547,I2683,I604100,I604089,);
nor I_35404 (I604578,I747129,I747132);
or I_35405 (I604080,I604327,I604578);
nor I_35406 (I604071,I604460,I604578);
or I_35407 (I604074,I604194,I604578);
DFFARX1 I_35408 (I604578,I2683,I604100,I604092,);
not I_35409 (I604678,I2690);
DFFARX1 I_35410 (I457256,I2683,I604678,I604704,);
not I_35411 (I604712,I604704);
nand I_35412 (I604729,I457265,I457274);
and I_35413 (I604746,I604729,I457280);
DFFARX1 I_35414 (I604746,I2683,I604678,I604772,);
not I_35415 (I604780,I457277);
DFFARX1 I_35416 (I457262,I2683,I604678,I604806,);
not I_35417 (I604814,I604806);
nor I_35418 (I604831,I604814,I604712);
and I_35419 (I604848,I604831,I457277);
nor I_35420 (I604865,I604814,I604780);
nor I_35421 (I604661,I604772,I604865);
DFFARX1 I_35422 (I457271,I2683,I604678,I604905,);
nor I_35423 (I604913,I604905,I604772);
not I_35424 (I604930,I604913);
not I_35425 (I604947,I604905);
nor I_35426 (I604964,I604947,I604848);
DFFARX1 I_35427 (I604964,I2683,I604678,I604664,);
nand I_35428 (I604995,I457268,I457259);
and I_35429 (I605012,I604995,I457256);
DFFARX1 I_35430 (I605012,I2683,I604678,I605038,);
nor I_35431 (I605046,I605038,I604905);
DFFARX1 I_35432 (I605046,I2683,I604678,I604646,);
nand I_35433 (I605077,I605038,I604947);
nand I_35434 (I604655,I604930,I605077);
not I_35435 (I605108,I605038);
nor I_35436 (I605125,I605108,I604848);
DFFARX1 I_35437 (I605125,I2683,I604678,I604667,);
nor I_35438 (I605156,I457259,I457259);
or I_35439 (I604658,I604905,I605156);
nor I_35440 (I604649,I605038,I605156);
or I_35441 (I604652,I604772,I605156);
DFFARX1 I_35442 (I605156,I2683,I604678,I604670,);
not I_35443 (I605256,I2690);
DFFARX1 I_35444 (I694472,I2683,I605256,I605282,);
not I_35445 (I605290,I605282);
nand I_35446 (I605307,I694460,I694478);
and I_35447 (I605324,I605307,I694475);
DFFARX1 I_35448 (I605324,I2683,I605256,I605350,);
not I_35449 (I605358,I694466);
DFFARX1 I_35450 (I694463,I2683,I605256,I605384,);
not I_35451 (I605392,I605384);
nor I_35452 (I605409,I605392,I605290);
and I_35453 (I605426,I605409,I694466);
nor I_35454 (I605443,I605392,I605358);
nor I_35455 (I605239,I605350,I605443);
DFFARX1 I_35456 (I694457,I2683,I605256,I605483,);
nor I_35457 (I605491,I605483,I605350);
not I_35458 (I605508,I605491);
not I_35459 (I605525,I605483);
nor I_35460 (I605542,I605525,I605426);
DFFARX1 I_35461 (I605542,I2683,I605256,I605242,);
nand I_35462 (I605573,I694457,I694460);
and I_35463 (I605590,I605573,I694463);
DFFARX1 I_35464 (I605590,I2683,I605256,I605616,);
nor I_35465 (I605624,I605616,I605483);
DFFARX1 I_35466 (I605624,I2683,I605256,I605224,);
nand I_35467 (I605655,I605616,I605525);
nand I_35468 (I605233,I605508,I605655);
not I_35469 (I605686,I605616);
nor I_35470 (I605703,I605686,I605426);
DFFARX1 I_35471 (I605703,I2683,I605256,I605245,);
nor I_35472 (I605734,I694469,I694460);
or I_35473 (I605236,I605483,I605734);
nor I_35474 (I605227,I605616,I605734);
or I_35475 (I605230,I605350,I605734);
DFFARX1 I_35476 (I605734,I2683,I605256,I605248,);
not I_35477 (I605834,I2690);
DFFARX1 I_35478 (I194385,I2683,I605834,I605860,);
not I_35479 (I605868,I605860);
nand I_35480 (I605885,I194388,I194409);
and I_35481 (I605902,I605885,I194397);
DFFARX1 I_35482 (I605902,I2683,I605834,I605928,);
not I_35483 (I605936,I194394);
DFFARX1 I_35484 (I194385,I2683,I605834,I605962,);
not I_35485 (I605970,I605962);
nor I_35486 (I605987,I605970,I605868);
and I_35487 (I606004,I605987,I194394);
nor I_35488 (I606021,I605970,I605936);
nor I_35489 (I605817,I605928,I606021);
DFFARX1 I_35490 (I194403,I2683,I605834,I606061,);
nor I_35491 (I606069,I606061,I605928);
not I_35492 (I606086,I606069);
not I_35493 (I606103,I606061);
nor I_35494 (I606120,I606103,I606004);
DFFARX1 I_35495 (I606120,I2683,I605834,I605820,);
nand I_35496 (I606151,I194388,I194391);
and I_35497 (I606168,I606151,I194400);
DFFARX1 I_35498 (I606168,I2683,I605834,I606194,);
nor I_35499 (I606202,I606194,I606061);
DFFARX1 I_35500 (I606202,I2683,I605834,I605802,);
nand I_35501 (I606233,I606194,I606103);
nand I_35502 (I605811,I606086,I606233);
not I_35503 (I606264,I606194);
nor I_35504 (I606281,I606264,I606004);
DFFARX1 I_35505 (I606281,I2683,I605834,I605823,);
nor I_35506 (I606312,I194406,I194391);
or I_35507 (I605814,I606061,I606312);
nor I_35508 (I605805,I606194,I606312);
or I_35509 (I605808,I605928,I606312);
DFFARX1 I_35510 (I606312,I2683,I605834,I605826,);
not I_35511 (I606412,I2690);
DFFARX1 I_35512 (I313902,I2683,I606412,I606438,);
not I_35513 (I606446,I606438);
nand I_35514 (I606463,I313905,I313881);
and I_35515 (I606480,I606463,I313878);
DFFARX1 I_35516 (I606480,I2683,I606412,I606506,);
not I_35517 (I606514,I313884);
DFFARX1 I_35518 (I313878,I2683,I606412,I606540,);
not I_35519 (I606548,I606540);
nor I_35520 (I606565,I606548,I606446);
and I_35521 (I606582,I606565,I313884);
nor I_35522 (I606599,I606548,I606514);
nor I_35523 (I606395,I606506,I606599);
DFFARX1 I_35524 (I313887,I2683,I606412,I606639,);
nor I_35525 (I606647,I606639,I606506);
not I_35526 (I606664,I606647);
not I_35527 (I606681,I606639);
nor I_35528 (I606698,I606681,I606582);
DFFARX1 I_35529 (I606698,I2683,I606412,I606398,);
nand I_35530 (I606729,I313890,I313899);
and I_35531 (I606746,I606729,I313896);
DFFARX1 I_35532 (I606746,I2683,I606412,I606772,);
nor I_35533 (I606780,I606772,I606639);
DFFARX1 I_35534 (I606780,I2683,I606412,I606380,);
nand I_35535 (I606811,I606772,I606681);
nand I_35536 (I606389,I606664,I606811);
not I_35537 (I606842,I606772);
nor I_35538 (I606859,I606842,I606582);
DFFARX1 I_35539 (I606859,I2683,I606412,I606401,);
nor I_35540 (I606890,I313893,I313899);
or I_35541 (I606392,I606639,I606890);
nor I_35542 (I606383,I606772,I606890);
or I_35543 (I606386,I606506,I606890);
DFFARX1 I_35544 (I606890,I2683,I606412,I606404,);
not I_35545 (I606990,I2690);
DFFARX1 I_35546 (I813055,I2683,I606990,I607016,);
not I_35547 (I607024,I607016);
nand I_35548 (I607041,I813052,I813070);
and I_35549 (I607058,I607041,I813067);
DFFARX1 I_35550 (I607058,I2683,I606990,I607084,);
not I_35551 (I607092,I813049);
DFFARX1 I_35552 (I813052,I2683,I606990,I607118,);
not I_35553 (I607126,I607118);
nor I_35554 (I607143,I607126,I607024);
and I_35555 (I607160,I607143,I813049);
nor I_35556 (I607177,I607126,I607092);
nor I_35557 (I606973,I607084,I607177);
DFFARX1 I_35558 (I813061,I2683,I606990,I607217,);
nor I_35559 (I607225,I607217,I607084);
not I_35560 (I607242,I607225);
not I_35561 (I607259,I607217);
nor I_35562 (I607276,I607259,I607160);
DFFARX1 I_35563 (I607276,I2683,I606990,I606976,);
nand I_35564 (I607307,I813064,I813049);
and I_35565 (I607324,I607307,I813055);
DFFARX1 I_35566 (I607324,I2683,I606990,I607350,);
nor I_35567 (I607358,I607350,I607217);
DFFARX1 I_35568 (I607358,I2683,I606990,I606958,);
nand I_35569 (I607389,I607350,I607259);
nand I_35570 (I606967,I607242,I607389);
not I_35571 (I607420,I607350);
nor I_35572 (I607437,I607420,I607160);
DFFARX1 I_35573 (I607437,I2683,I606990,I606979,);
nor I_35574 (I607468,I813058,I813049);
or I_35575 (I606970,I607217,I607468);
nor I_35576 (I606961,I607350,I607468);
or I_35577 (I606964,I607084,I607468);
DFFARX1 I_35578 (I607468,I2683,I606990,I606982,);
not I_35579 (I607568,I2690);
DFFARX1 I_35580 (I3294,I2683,I607568,I607594,);
not I_35581 (I607602,I607594);
nand I_35582 (I607619,I3297,I3309);
and I_35583 (I607636,I607619,I3288);
DFFARX1 I_35584 (I607636,I2683,I607568,I607662,);
not I_35585 (I607670,I3288);
DFFARX1 I_35586 (I3291,I2683,I607568,I607696,);
not I_35587 (I607704,I607696);
nor I_35588 (I607721,I607704,I607602);
and I_35589 (I607738,I607721,I3288);
nor I_35590 (I607755,I607704,I607670);
nor I_35591 (I607551,I607662,I607755);
DFFARX1 I_35592 (I3303,I2683,I607568,I607795,);
nor I_35593 (I607803,I607795,I607662);
not I_35594 (I607820,I607803);
not I_35595 (I607837,I607795);
nor I_35596 (I607854,I607837,I607738);
DFFARX1 I_35597 (I607854,I2683,I607568,I607554,);
nand I_35598 (I607885,I3306,I3291);
and I_35599 (I607902,I607885,I3300);
DFFARX1 I_35600 (I607902,I2683,I607568,I607928,);
nor I_35601 (I607936,I607928,I607795);
DFFARX1 I_35602 (I607936,I2683,I607568,I607536,);
nand I_35603 (I607967,I607928,I607837);
nand I_35604 (I607545,I607820,I607967);
not I_35605 (I607998,I607928);
nor I_35606 (I608015,I607998,I607738);
DFFARX1 I_35607 (I608015,I2683,I607568,I607557,);
nor I_35608 (I608046,I3294,I3291);
or I_35609 (I607548,I607795,I608046);
nor I_35610 (I607539,I607928,I608046);
or I_35611 (I607542,I607662,I608046);
DFFARX1 I_35612 (I608046,I2683,I607568,I607560,);
not I_35613 (I608146,I2690);
DFFARX1 I_35614 (I712909,I2683,I608146,I608172,);
not I_35615 (I608180,I608172);
nand I_35616 (I608197,I712885,I712900);
and I_35617 (I608214,I608197,I712912);
DFFARX1 I_35618 (I608214,I2683,I608146,I608240,);
not I_35619 (I608248,I712897);
DFFARX1 I_35620 (I712888,I2683,I608146,I608274,);
not I_35621 (I608282,I608274);
nor I_35622 (I608299,I608282,I608180);
and I_35623 (I608316,I608299,I712897);
nor I_35624 (I608333,I608282,I608248);
nor I_35625 (I608129,I608240,I608333);
DFFARX1 I_35626 (I712885,I2683,I608146,I608373,);
nor I_35627 (I608381,I608373,I608240);
not I_35628 (I608398,I608381);
not I_35629 (I608415,I608373);
nor I_35630 (I608432,I608415,I608316);
DFFARX1 I_35631 (I608432,I2683,I608146,I608132,);
nand I_35632 (I608463,I712903,I712894);
and I_35633 (I608480,I608463,I712906);
DFFARX1 I_35634 (I608480,I2683,I608146,I608506,);
nor I_35635 (I608514,I608506,I608373);
DFFARX1 I_35636 (I608514,I2683,I608146,I608114,);
nand I_35637 (I608545,I608506,I608415);
nand I_35638 (I608123,I608398,I608545);
not I_35639 (I608576,I608506);
nor I_35640 (I608593,I608576,I608316);
DFFARX1 I_35641 (I608593,I2683,I608146,I608135,);
nor I_35642 (I608624,I712891,I712894);
or I_35643 (I608126,I608373,I608624);
nor I_35644 (I608117,I608506,I608624);
or I_35645 (I608120,I608240,I608624);
DFFARX1 I_35646 (I608624,I2683,I608146,I608138,);
not I_35647 (I608724,I2690);
DFFARX1 I_35648 (I139645,I2683,I608724,I608750,);
not I_35649 (I608758,I608750);
nand I_35650 (I608775,I139648,I139669);
and I_35651 (I608792,I608775,I139657);
DFFARX1 I_35652 (I608792,I2683,I608724,I608818,);
not I_35653 (I608826,I139654);
DFFARX1 I_35654 (I139645,I2683,I608724,I608852,);
not I_35655 (I608860,I608852);
nor I_35656 (I608877,I608860,I608758);
and I_35657 (I608894,I608877,I139654);
nor I_35658 (I608911,I608860,I608826);
nor I_35659 (I608707,I608818,I608911);
DFFARX1 I_35660 (I139663,I2683,I608724,I608951,);
nor I_35661 (I608959,I608951,I608818);
not I_35662 (I608976,I608959);
not I_35663 (I608993,I608951);
nor I_35664 (I609010,I608993,I608894);
DFFARX1 I_35665 (I609010,I2683,I608724,I608710,);
nand I_35666 (I609041,I139648,I139651);
and I_35667 (I609058,I609041,I139660);
DFFARX1 I_35668 (I609058,I2683,I608724,I609084,);
nor I_35669 (I609092,I609084,I608951);
DFFARX1 I_35670 (I609092,I2683,I608724,I608692,);
nand I_35671 (I609123,I609084,I608993);
nand I_35672 (I608701,I608976,I609123);
not I_35673 (I609154,I609084);
nor I_35674 (I609171,I609154,I608894);
DFFARX1 I_35675 (I609171,I2683,I608724,I608713,);
nor I_35676 (I609202,I139666,I139651);
or I_35677 (I608704,I608951,I609202);
nor I_35678 (I608695,I609084,I609202);
or I_35679 (I608698,I608818,I609202);
DFFARX1 I_35680 (I609202,I2683,I608724,I608716,);
not I_35681 (I609302,I2690);
DFFARX1 I_35682 (I1059066,I2683,I609302,I609328,);
not I_35683 (I609336,I609328);
nand I_35684 (I609353,I1059051,I1059039);
and I_35685 (I609370,I609353,I1059054);
DFFARX1 I_35686 (I609370,I2683,I609302,I609396,);
not I_35687 (I609404,I1059039);
DFFARX1 I_35688 (I1059057,I2683,I609302,I609430,);
not I_35689 (I609438,I609430);
nor I_35690 (I609455,I609438,I609336);
and I_35691 (I609472,I609455,I1059039);
nor I_35692 (I609489,I609438,I609404);
nor I_35693 (I609285,I609396,I609489);
DFFARX1 I_35694 (I1059045,I2683,I609302,I609529,);
nor I_35695 (I609537,I609529,I609396);
not I_35696 (I609554,I609537);
not I_35697 (I609571,I609529);
nor I_35698 (I609588,I609571,I609472);
DFFARX1 I_35699 (I609588,I2683,I609302,I609288,);
nand I_35700 (I609619,I1059042,I1059048);
and I_35701 (I609636,I609619,I1059063);
DFFARX1 I_35702 (I609636,I2683,I609302,I609662,);
nor I_35703 (I609670,I609662,I609529);
DFFARX1 I_35704 (I609670,I2683,I609302,I609270,);
nand I_35705 (I609701,I609662,I609571);
nand I_35706 (I609279,I609554,I609701);
not I_35707 (I609732,I609662);
nor I_35708 (I609749,I609732,I609472);
DFFARX1 I_35709 (I609749,I2683,I609302,I609291,);
nor I_35710 (I609780,I1059060,I1059048);
or I_35711 (I609282,I609529,I609780);
nor I_35712 (I609273,I609662,I609780);
or I_35713 (I609276,I609396,I609780);
DFFARX1 I_35714 (I609780,I2683,I609302,I609294,);
not I_35715 (I609880,I2690);
DFFARX1 I_35716 (I1082866,I2683,I609880,I609906,);
not I_35717 (I609914,I609906);
nand I_35718 (I609931,I1082851,I1082839);
and I_35719 (I609948,I609931,I1082854);
DFFARX1 I_35720 (I609948,I2683,I609880,I609974,);
not I_35721 (I609982,I1082839);
DFFARX1 I_35722 (I1082857,I2683,I609880,I610008,);
not I_35723 (I610016,I610008);
nor I_35724 (I610033,I610016,I609914);
and I_35725 (I610050,I610033,I1082839);
nor I_35726 (I610067,I610016,I609982);
nor I_35727 (I609863,I609974,I610067);
DFFARX1 I_35728 (I1082845,I2683,I609880,I610107,);
nor I_35729 (I610115,I610107,I609974);
not I_35730 (I610132,I610115);
not I_35731 (I610149,I610107);
nor I_35732 (I610166,I610149,I610050);
DFFARX1 I_35733 (I610166,I2683,I609880,I609866,);
nand I_35734 (I610197,I1082842,I1082848);
and I_35735 (I610214,I610197,I1082863);
DFFARX1 I_35736 (I610214,I2683,I609880,I610240,);
nor I_35737 (I610248,I610240,I610107);
DFFARX1 I_35738 (I610248,I2683,I609880,I609848,);
nand I_35739 (I610279,I610240,I610149);
nand I_35740 (I609857,I610132,I610279);
not I_35741 (I610310,I610240);
nor I_35742 (I610327,I610310,I610050);
DFFARX1 I_35743 (I610327,I2683,I609880,I609869,);
nor I_35744 (I610358,I1082860,I1082848);
or I_35745 (I609860,I610107,I610358);
nor I_35746 (I609851,I610240,I610358);
or I_35747 (I609854,I609974,I610358);
DFFARX1 I_35748 (I610358,I2683,I609880,I609872,);
not I_35749 (I610458,I2690);
DFFARX1 I_35750 (I725183,I2683,I610458,I610484,);
not I_35751 (I610492,I610484);
nand I_35752 (I610509,I725159,I725174);
and I_35753 (I610526,I610509,I725186);
DFFARX1 I_35754 (I610526,I2683,I610458,I610552,);
not I_35755 (I610560,I725171);
DFFARX1 I_35756 (I725162,I2683,I610458,I610586,);
not I_35757 (I610594,I610586);
nor I_35758 (I610611,I610594,I610492);
and I_35759 (I610628,I610611,I725171);
nor I_35760 (I610645,I610594,I610560);
nor I_35761 (I610441,I610552,I610645);
DFFARX1 I_35762 (I725159,I2683,I610458,I610685,);
nor I_35763 (I610693,I610685,I610552);
not I_35764 (I610710,I610693);
not I_35765 (I610727,I610685);
nor I_35766 (I610744,I610727,I610628);
DFFARX1 I_35767 (I610744,I2683,I610458,I610444,);
nand I_35768 (I610775,I725177,I725168);
and I_35769 (I610792,I610775,I725180);
DFFARX1 I_35770 (I610792,I2683,I610458,I610818,);
nor I_35771 (I610826,I610818,I610685);
DFFARX1 I_35772 (I610826,I2683,I610458,I610426,);
nand I_35773 (I610857,I610818,I610727);
nand I_35774 (I610435,I610710,I610857);
not I_35775 (I610888,I610818);
nor I_35776 (I610905,I610888,I610628);
DFFARX1 I_35777 (I610905,I2683,I610458,I610447,);
nor I_35778 (I610936,I725165,I725168);
or I_35779 (I610438,I610685,I610936);
nor I_35780 (I610429,I610818,I610936);
or I_35781 (I610432,I610552,I610936);
DFFARX1 I_35782 (I610936,I2683,I610458,I610450,);
not I_35783 (I611036,I2690);
DFFARX1 I_35784 (I464192,I2683,I611036,I611062,);
not I_35785 (I611070,I611062);
nand I_35786 (I611087,I464201,I464210);
and I_35787 (I611104,I611087,I464216);
DFFARX1 I_35788 (I611104,I2683,I611036,I611130,);
not I_35789 (I611138,I464213);
DFFARX1 I_35790 (I464198,I2683,I611036,I611164,);
not I_35791 (I611172,I611164);
nor I_35792 (I611189,I611172,I611070);
and I_35793 (I611206,I611189,I464213);
nor I_35794 (I611223,I611172,I611138);
nor I_35795 (I611019,I611130,I611223);
DFFARX1 I_35796 (I464207,I2683,I611036,I611263,);
nor I_35797 (I611271,I611263,I611130);
not I_35798 (I611288,I611271);
not I_35799 (I611305,I611263);
nor I_35800 (I611322,I611305,I611206);
DFFARX1 I_35801 (I611322,I2683,I611036,I611022,);
nand I_35802 (I611353,I464204,I464195);
and I_35803 (I611370,I611353,I464192);
DFFARX1 I_35804 (I611370,I2683,I611036,I611396,);
nor I_35805 (I611404,I611396,I611263);
DFFARX1 I_35806 (I611404,I2683,I611036,I611004,);
nand I_35807 (I611435,I611396,I611305);
nand I_35808 (I611013,I611288,I611435);
not I_35809 (I611466,I611396);
nor I_35810 (I611483,I611466,I611206);
DFFARX1 I_35811 (I611483,I2683,I611036,I611025,);
nor I_35812 (I611514,I464195,I464195);
or I_35813 (I611016,I611263,I611514);
nor I_35814 (I611007,I611396,I611514);
or I_35815 (I611010,I611130,I611514);
DFFARX1 I_35816 (I611514,I2683,I611036,I611028,);
not I_35817 (I611614,I2690);
DFFARX1 I_35818 (I855958,I2683,I611614,I611640,);
not I_35819 (I611648,I611640);
nand I_35820 (I611665,I855940,I855952);
and I_35821 (I611682,I611665,I855955);
DFFARX1 I_35822 (I611682,I2683,I611614,I611708,);
not I_35823 (I611716,I855949);
DFFARX1 I_35824 (I855946,I2683,I611614,I611742,);
not I_35825 (I611750,I611742);
nor I_35826 (I611767,I611750,I611648);
and I_35827 (I611784,I611767,I855949);
nor I_35828 (I611801,I611750,I611716);
nor I_35829 (I611597,I611708,I611801);
DFFARX1 I_35830 (I855964,I2683,I611614,I611841,);
nor I_35831 (I611849,I611841,I611708);
not I_35832 (I611866,I611849);
not I_35833 (I611883,I611841);
nor I_35834 (I611900,I611883,I611784);
DFFARX1 I_35835 (I611900,I2683,I611614,I611600,);
nand I_35836 (I611931,I855943,I855943);
and I_35837 (I611948,I611931,I855940);
DFFARX1 I_35838 (I611948,I2683,I611614,I611974,);
nor I_35839 (I611982,I611974,I611841);
DFFARX1 I_35840 (I611982,I2683,I611614,I611582,);
nand I_35841 (I612013,I611974,I611883);
nand I_35842 (I611591,I611866,I612013);
not I_35843 (I612044,I611974);
nor I_35844 (I612061,I612044,I611784);
DFFARX1 I_35845 (I612061,I2683,I611614,I611603,);
nor I_35846 (I612092,I855961,I855943);
or I_35847 (I611594,I611841,I612092);
nor I_35848 (I611585,I611974,I612092);
or I_35849 (I611588,I611708,I612092);
DFFARX1 I_35850 (I612092,I2683,I611614,I611606,);
not I_35851 (I612192,I2690);
DFFARX1 I_35852 (I402057,I2683,I612192,I612218,);
not I_35853 (I612226,I612218);
nand I_35854 (I612243,I402072,I402057);
and I_35855 (I612260,I612243,I402060);
DFFARX1 I_35856 (I612260,I2683,I612192,I612286,);
not I_35857 (I612294,I402060);
DFFARX1 I_35858 (I402069,I2683,I612192,I612320,);
not I_35859 (I612328,I612320);
nor I_35860 (I612345,I612328,I612226);
and I_35861 (I612362,I612345,I402060);
nor I_35862 (I612379,I612328,I612294);
nor I_35863 (I612175,I612286,I612379);
DFFARX1 I_35864 (I402063,I2683,I612192,I612419,);
nor I_35865 (I612427,I612419,I612286);
not I_35866 (I612444,I612427);
not I_35867 (I612461,I612419);
nor I_35868 (I612478,I612461,I612362);
DFFARX1 I_35869 (I612478,I2683,I612192,I612178,);
nand I_35870 (I612509,I402066,I402075);
and I_35871 (I612526,I612509,I402081);
DFFARX1 I_35872 (I612526,I2683,I612192,I612552,);
nor I_35873 (I612560,I612552,I612419);
DFFARX1 I_35874 (I612560,I2683,I612192,I612160,);
nand I_35875 (I612591,I612552,I612461);
nand I_35876 (I612169,I612444,I612591);
not I_35877 (I612622,I612552);
nor I_35878 (I612639,I612622,I612362);
DFFARX1 I_35879 (I612639,I2683,I612192,I612181,);
nor I_35880 (I612670,I402078,I402075);
or I_35881 (I612172,I612419,I612670);
nor I_35882 (I612163,I612552,I612670);
or I_35883 (I612166,I612286,I612670);
DFFARX1 I_35884 (I612670,I2683,I612192,I612184,);
not I_35885 (I612770,I2690);
DFFARX1 I_35886 (I453788,I2683,I612770,I612796,);
not I_35887 (I612804,I612796);
nand I_35888 (I612821,I453797,I453806);
and I_35889 (I612838,I612821,I453812);
DFFARX1 I_35890 (I612838,I2683,I612770,I612864,);
not I_35891 (I612872,I453809);
DFFARX1 I_35892 (I453794,I2683,I612770,I612898,);
not I_35893 (I612906,I612898);
nor I_35894 (I612923,I612906,I612804);
and I_35895 (I612940,I612923,I453809);
nor I_35896 (I612957,I612906,I612872);
nor I_35897 (I612753,I612864,I612957);
DFFARX1 I_35898 (I453803,I2683,I612770,I612997,);
nor I_35899 (I613005,I612997,I612864);
not I_35900 (I613022,I613005);
not I_35901 (I613039,I612997);
nor I_35902 (I613056,I613039,I612940);
DFFARX1 I_35903 (I613056,I2683,I612770,I612756,);
nand I_35904 (I613087,I453800,I453791);
and I_35905 (I613104,I613087,I453788);
DFFARX1 I_35906 (I613104,I2683,I612770,I613130,);
nor I_35907 (I613138,I613130,I612997);
DFFARX1 I_35908 (I613138,I2683,I612770,I612738,);
nand I_35909 (I613169,I613130,I613039);
nand I_35910 (I612747,I613022,I613169);
not I_35911 (I613200,I613130);
nor I_35912 (I613217,I613200,I612940);
DFFARX1 I_35913 (I613217,I2683,I612770,I612759,);
nor I_35914 (I613248,I453791,I453791);
or I_35915 (I612750,I612997,I613248);
nor I_35916 (I612741,I613130,I613248);
or I_35917 (I612744,I612864,I613248);
DFFARX1 I_35918 (I613248,I2683,I612770,I612762,);
not I_35919 (I613348,I2690);
DFFARX1 I_35920 (I691310,I2683,I613348,I613374,);
not I_35921 (I613382,I613374);
nand I_35922 (I613399,I691298,I691316);
and I_35923 (I613416,I613399,I691313);
DFFARX1 I_35924 (I613416,I2683,I613348,I613442,);
not I_35925 (I613450,I691304);
DFFARX1 I_35926 (I691301,I2683,I613348,I613476,);
not I_35927 (I613484,I613476);
nor I_35928 (I613501,I613484,I613382);
and I_35929 (I613518,I613501,I691304);
nor I_35930 (I613535,I613484,I613450);
nor I_35931 (I613331,I613442,I613535);
DFFARX1 I_35932 (I691295,I2683,I613348,I613575,);
nor I_35933 (I613583,I613575,I613442);
not I_35934 (I613600,I613583);
not I_35935 (I613617,I613575);
nor I_35936 (I613634,I613617,I613518);
DFFARX1 I_35937 (I613634,I2683,I613348,I613334,);
nand I_35938 (I613665,I691295,I691298);
and I_35939 (I613682,I613665,I691301);
DFFARX1 I_35940 (I613682,I2683,I613348,I613708,);
nor I_35941 (I613716,I613708,I613575);
DFFARX1 I_35942 (I613716,I2683,I613348,I613316,);
nand I_35943 (I613747,I613708,I613617);
nand I_35944 (I613325,I613600,I613747);
not I_35945 (I613778,I613708);
nor I_35946 (I613795,I613778,I613518);
DFFARX1 I_35947 (I613795,I2683,I613348,I613337,);
nor I_35948 (I613826,I691307,I691298);
or I_35949 (I613328,I613575,I613826);
nor I_35950 (I613319,I613708,I613826);
or I_35951 (I613322,I613442,I613826);
DFFARX1 I_35952 (I613826,I2683,I613348,I613340,);
not I_35953 (I613926,I2690);
DFFARX1 I_35954 (I854802,I2683,I613926,I613952,);
not I_35955 (I613960,I613952);
nand I_35956 (I613977,I854784,I854796);
and I_35957 (I613994,I613977,I854799);
DFFARX1 I_35958 (I613994,I2683,I613926,I614020,);
not I_35959 (I614028,I854793);
DFFARX1 I_35960 (I854790,I2683,I613926,I614054,);
not I_35961 (I614062,I614054);
nor I_35962 (I614079,I614062,I613960);
and I_35963 (I614096,I614079,I854793);
nor I_35964 (I614113,I614062,I614028);
nor I_35965 (I613909,I614020,I614113);
DFFARX1 I_35966 (I854808,I2683,I613926,I614153,);
nor I_35967 (I614161,I614153,I614020);
not I_35968 (I614178,I614161);
not I_35969 (I614195,I614153);
nor I_35970 (I614212,I614195,I614096);
DFFARX1 I_35971 (I614212,I2683,I613926,I613912,);
nand I_35972 (I614243,I854787,I854787);
and I_35973 (I614260,I614243,I854784);
DFFARX1 I_35974 (I614260,I2683,I613926,I614286,);
nor I_35975 (I614294,I614286,I614153);
DFFARX1 I_35976 (I614294,I2683,I613926,I613894,);
nand I_35977 (I614325,I614286,I614195);
nand I_35978 (I613903,I614178,I614325);
not I_35979 (I614356,I614286);
nor I_35980 (I614373,I614356,I614096);
DFFARX1 I_35981 (I614373,I2683,I613926,I613915,);
nor I_35982 (I614404,I854805,I854787);
or I_35983 (I613906,I614153,I614404);
nor I_35984 (I613897,I614286,I614404);
or I_35985 (I613900,I614020,I614404);
DFFARX1 I_35986 (I614404,I2683,I613926,I613918,);
not I_35987 (I614504,I2690);
DFFARX1 I_35988 (I1076321,I2683,I614504,I614530,);
not I_35989 (I614538,I614530);
nand I_35990 (I614555,I1076306,I1076294);
and I_35991 (I614572,I614555,I1076309);
DFFARX1 I_35992 (I614572,I2683,I614504,I614598,);
not I_35993 (I614606,I1076294);
DFFARX1 I_35994 (I1076312,I2683,I614504,I614632,);
not I_35995 (I614640,I614632);
nor I_35996 (I614657,I614640,I614538);
and I_35997 (I614674,I614657,I1076294);
nor I_35998 (I614691,I614640,I614606);
nor I_35999 (I614487,I614598,I614691);
DFFARX1 I_36000 (I1076300,I2683,I614504,I614731,);
nor I_36001 (I614739,I614731,I614598);
not I_36002 (I614756,I614739);
not I_36003 (I614773,I614731);
nor I_36004 (I614790,I614773,I614674);
DFFARX1 I_36005 (I614790,I2683,I614504,I614490,);
nand I_36006 (I614821,I1076297,I1076303);
and I_36007 (I614838,I614821,I1076318);
DFFARX1 I_36008 (I614838,I2683,I614504,I614864,);
nor I_36009 (I614872,I614864,I614731);
DFFARX1 I_36010 (I614872,I2683,I614504,I614472,);
nand I_36011 (I614903,I614864,I614773);
nand I_36012 (I614481,I614756,I614903);
not I_36013 (I614934,I614864);
nor I_36014 (I614951,I614934,I614674);
DFFARX1 I_36015 (I614951,I2683,I614504,I614493,);
nor I_36016 (I614982,I1076315,I1076303);
or I_36017 (I614484,I614731,I614982);
nor I_36018 (I614475,I614864,I614982);
or I_36019 (I614478,I614598,I614982);
DFFARX1 I_36020 (I614982,I2683,I614504,I614496,);
not I_36021 (I615082,I2690);
DFFARX1 I_36022 (I165825,I2683,I615082,I615108,);
not I_36023 (I615116,I615108);
nand I_36024 (I615133,I165828,I165849);
and I_36025 (I615150,I615133,I165837);
DFFARX1 I_36026 (I615150,I2683,I615082,I615176,);
not I_36027 (I615184,I165834);
DFFARX1 I_36028 (I165825,I2683,I615082,I615210,);
not I_36029 (I615218,I615210);
nor I_36030 (I615235,I615218,I615116);
and I_36031 (I615252,I615235,I165834);
nor I_36032 (I615269,I615218,I615184);
nor I_36033 (I615065,I615176,I615269);
DFFARX1 I_36034 (I165843,I2683,I615082,I615309,);
nor I_36035 (I615317,I615309,I615176);
not I_36036 (I615334,I615317);
not I_36037 (I615351,I615309);
nor I_36038 (I615368,I615351,I615252);
DFFARX1 I_36039 (I615368,I2683,I615082,I615068,);
nand I_36040 (I615399,I165828,I165831);
and I_36041 (I615416,I615399,I165840);
DFFARX1 I_36042 (I615416,I2683,I615082,I615442,);
nor I_36043 (I615450,I615442,I615309);
DFFARX1 I_36044 (I615450,I2683,I615082,I615050,);
nand I_36045 (I615481,I615442,I615351);
nand I_36046 (I615059,I615334,I615481);
not I_36047 (I615512,I615442);
nor I_36048 (I615529,I615512,I615252);
DFFARX1 I_36049 (I615529,I2683,I615082,I615071,);
nor I_36050 (I615560,I165846,I165831);
or I_36051 (I615062,I615309,I615560);
nor I_36052 (I615053,I615442,I615560);
or I_36053 (I615056,I615176,I615560);
DFFARX1 I_36054 (I615560,I2683,I615082,I615074,);
not I_36055 (I615660,I2690);
DFFARX1 I_36056 (I472284,I2683,I615660,I615686,);
not I_36057 (I615694,I615686);
nand I_36058 (I615711,I472293,I472302);
and I_36059 (I615728,I615711,I472308);
DFFARX1 I_36060 (I615728,I2683,I615660,I615754,);
not I_36061 (I615762,I472305);
DFFARX1 I_36062 (I472290,I2683,I615660,I615788,);
not I_36063 (I615796,I615788);
nor I_36064 (I615813,I615796,I615694);
and I_36065 (I615830,I615813,I472305);
nor I_36066 (I615847,I615796,I615762);
nor I_36067 (I615643,I615754,I615847);
DFFARX1 I_36068 (I472299,I2683,I615660,I615887,);
nor I_36069 (I615895,I615887,I615754);
not I_36070 (I615912,I615895);
not I_36071 (I615929,I615887);
nor I_36072 (I615946,I615929,I615830);
DFFARX1 I_36073 (I615946,I2683,I615660,I615646,);
nand I_36074 (I615977,I472296,I472287);
and I_36075 (I615994,I615977,I472284);
DFFARX1 I_36076 (I615994,I2683,I615660,I616020,);
nor I_36077 (I616028,I616020,I615887);
DFFARX1 I_36078 (I616028,I2683,I615660,I615628,);
nand I_36079 (I616059,I616020,I615929);
nand I_36080 (I615637,I615912,I616059);
not I_36081 (I616090,I616020);
nor I_36082 (I616107,I616090,I615830);
DFFARX1 I_36083 (I616107,I2683,I615660,I615649,);
nor I_36084 (I616138,I472287,I472287);
or I_36085 (I615640,I615887,I616138);
nor I_36086 (I615631,I616020,I616138);
or I_36087 (I615634,I615754,I616138);
DFFARX1 I_36088 (I616138,I2683,I615660,I615652,);
not I_36089 (I616238,I2690);
DFFARX1 I_36090 (I1098336,I2683,I616238,I616264,);
not I_36091 (I616272,I616264);
nand I_36092 (I616289,I1098321,I1098309);
and I_36093 (I616306,I616289,I1098324);
DFFARX1 I_36094 (I616306,I2683,I616238,I616332,);
not I_36095 (I616340,I1098309);
DFFARX1 I_36096 (I1098327,I2683,I616238,I616366,);
not I_36097 (I616374,I616366);
nor I_36098 (I616391,I616374,I616272);
and I_36099 (I616408,I616391,I1098309);
nor I_36100 (I616425,I616374,I616340);
nor I_36101 (I616221,I616332,I616425);
DFFARX1 I_36102 (I1098315,I2683,I616238,I616465,);
nor I_36103 (I616473,I616465,I616332);
not I_36104 (I616490,I616473);
not I_36105 (I616507,I616465);
nor I_36106 (I616524,I616507,I616408);
DFFARX1 I_36107 (I616524,I2683,I616238,I616224,);
nand I_36108 (I616555,I1098312,I1098318);
and I_36109 (I616572,I616555,I1098333);
DFFARX1 I_36110 (I616572,I2683,I616238,I616598,);
nor I_36111 (I616606,I616598,I616465);
DFFARX1 I_36112 (I616606,I2683,I616238,I616206,);
nand I_36113 (I616637,I616598,I616507);
nand I_36114 (I616215,I616490,I616637);
not I_36115 (I616668,I616598);
nor I_36116 (I616685,I616668,I616408);
DFFARX1 I_36117 (I616685,I2683,I616238,I616227,);
nor I_36118 (I616716,I1098330,I1098318);
or I_36119 (I616218,I616465,I616716);
nor I_36120 (I616209,I616598,I616716);
or I_36121 (I616212,I616332,I616716);
DFFARX1 I_36122 (I616716,I2683,I616238,I616230,);
not I_36123 (I616816,I2690);
DFFARX1 I_36124 (I54835,I2683,I616816,I616842,);
not I_36125 (I616850,I616842);
nand I_36126 (I616867,I54844,I54853);
and I_36127 (I616884,I616867,I54832);
DFFARX1 I_36128 (I616884,I2683,I616816,I616910,);
not I_36129 (I616918,I54835);
DFFARX1 I_36130 (I54850,I2683,I616816,I616944,);
not I_36131 (I616952,I616944);
nor I_36132 (I616969,I616952,I616850);
and I_36133 (I616986,I616969,I54835);
nor I_36134 (I617003,I616952,I616918);
nor I_36135 (I616799,I616910,I617003);
DFFARX1 I_36136 (I54841,I2683,I616816,I617043,);
nor I_36137 (I617051,I617043,I616910);
not I_36138 (I617068,I617051);
not I_36139 (I617085,I617043);
nor I_36140 (I617102,I617085,I616986);
DFFARX1 I_36141 (I617102,I2683,I616816,I616802,);
nand I_36142 (I617133,I54856,I54832);
and I_36143 (I617150,I617133,I54838);
DFFARX1 I_36144 (I617150,I2683,I616816,I617176,);
nor I_36145 (I617184,I617176,I617043);
DFFARX1 I_36146 (I617184,I2683,I616816,I616784,);
nand I_36147 (I617215,I617176,I617085);
nand I_36148 (I616793,I617068,I617215);
not I_36149 (I617246,I617176);
nor I_36150 (I617263,I617246,I616986);
DFFARX1 I_36151 (I617263,I2683,I616816,I616805,);
nor I_36152 (I617294,I54847,I54832);
or I_36153 (I616796,I617043,I617294);
nor I_36154 (I616787,I617176,I617294);
or I_36155 (I616790,I616910,I617294);
DFFARX1 I_36156 (I617294,I2683,I616816,I616808,);
not I_36157 (I617394,I2690);
DFFARX1 I_36158 (I832260,I2683,I617394,I617420,);
not I_36159 (I617428,I617420);
nand I_36160 (I617445,I832242,I832254);
and I_36161 (I617462,I617445,I832257);
DFFARX1 I_36162 (I617462,I2683,I617394,I617488,);
not I_36163 (I617496,I832251);
DFFARX1 I_36164 (I832248,I2683,I617394,I617522,);
not I_36165 (I617530,I617522);
nor I_36166 (I617547,I617530,I617428);
and I_36167 (I617564,I617547,I832251);
nor I_36168 (I617581,I617530,I617496);
nor I_36169 (I617377,I617488,I617581);
DFFARX1 I_36170 (I832266,I2683,I617394,I617621,);
nor I_36171 (I617629,I617621,I617488);
not I_36172 (I617646,I617629);
not I_36173 (I617663,I617621);
nor I_36174 (I617680,I617663,I617564);
DFFARX1 I_36175 (I617680,I2683,I617394,I617380,);
nand I_36176 (I617711,I832245,I832245);
and I_36177 (I617728,I617711,I832242);
DFFARX1 I_36178 (I617728,I2683,I617394,I617754,);
nor I_36179 (I617762,I617754,I617621);
DFFARX1 I_36180 (I617762,I2683,I617394,I617362,);
nand I_36181 (I617793,I617754,I617663);
nand I_36182 (I617371,I617646,I617793);
not I_36183 (I617824,I617754);
nor I_36184 (I617841,I617824,I617564);
DFFARX1 I_36185 (I617841,I2683,I617394,I617383,);
nor I_36186 (I617872,I832263,I832245);
or I_36187 (I617374,I617621,I617872);
nor I_36188 (I617365,I617754,I617872);
or I_36189 (I617368,I617488,I617872);
DFFARX1 I_36190 (I617872,I2683,I617394,I617386,);
not I_36191 (I617972,I2690);
DFFARX1 I_36192 (I198550,I2683,I617972,I617998,);
not I_36193 (I618006,I617998);
nand I_36194 (I618023,I198553,I198574);
and I_36195 (I618040,I618023,I198562);
DFFARX1 I_36196 (I618040,I2683,I617972,I618066,);
not I_36197 (I618074,I198559);
DFFARX1 I_36198 (I198550,I2683,I617972,I618100,);
not I_36199 (I618108,I618100);
nor I_36200 (I618125,I618108,I618006);
and I_36201 (I618142,I618125,I198559);
nor I_36202 (I618159,I618108,I618074);
nor I_36203 (I617955,I618066,I618159);
DFFARX1 I_36204 (I198568,I2683,I617972,I618199,);
nor I_36205 (I618207,I618199,I618066);
not I_36206 (I618224,I618207);
not I_36207 (I618241,I618199);
nor I_36208 (I618258,I618241,I618142);
DFFARX1 I_36209 (I618258,I2683,I617972,I617958,);
nand I_36210 (I618289,I198553,I198556);
and I_36211 (I618306,I618289,I198565);
DFFARX1 I_36212 (I618306,I2683,I617972,I618332,);
nor I_36213 (I618340,I618332,I618199);
DFFARX1 I_36214 (I618340,I2683,I617972,I617940,);
nand I_36215 (I618371,I618332,I618241);
nand I_36216 (I617949,I618224,I618371);
not I_36217 (I618402,I618332);
nor I_36218 (I618419,I618402,I618142);
DFFARX1 I_36219 (I618419,I2683,I617972,I617961,);
nor I_36220 (I618450,I198571,I198556);
or I_36221 (I617952,I618199,I618450);
nor I_36222 (I617943,I618332,I618450);
or I_36223 (I617946,I618066,I618450);
DFFARX1 I_36224 (I618450,I2683,I617972,I617964,);
not I_36225 (I618550,I2690);
DFFARX1 I_36226 (I985310,I2683,I618550,I618576,);
not I_36227 (I618584,I618576);
nand I_36228 (I618601,I985313,I985322);
and I_36229 (I618618,I618601,I985325);
DFFARX1 I_36230 (I618618,I2683,I618550,I618644,);
not I_36231 (I618652,I985334);
DFFARX1 I_36232 (I985316,I2683,I618550,I618678,);
not I_36233 (I618686,I618678);
nor I_36234 (I618703,I618686,I618584);
and I_36235 (I618720,I618703,I985334);
nor I_36236 (I618737,I618686,I618652);
nor I_36237 (I618533,I618644,I618737);
DFFARX1 I_36238 (I985313,I2683,I618550,I618777,);
nor I_36239 (I618785,I618777,I618644);
not I_36240 (I618802,I618785);
not I_36241 (I618819,I618777);
nor I_36242 (I618836,I618819,I618720);
DFFARX1 I_36243 (I618836,I2683,I618550,I618536,);
nand I_36244 (I618867,I985331,I985310);
and I_36245 (I618884,I618867,I985328);
DFFARX1 I_36246 (I618884,I2683,I618550,I618910,);
nor I_36247 (I618918,I618910,I618777);
DFFARX1 I_36248 (I618918,I2683,I618550,I618518,);
nand I_36249 (I618949,I618910,I618819);
nand I_36250 (I618527,I618802,I618949);
not I_36251 (I618980,I618910);
nor I_36252 (I618997,I618980,I618720);
DFFARX1 I_36253 (I618997,I2683,I618550,I618539,);
nor I_36254 (I619028,I985319,I985310);
or I_36255 (I618530,I618777,I619028);
nor I_36256 (I618521,I618910,I619028);
or I_36257 (I618524,I618644,I619028);
DFFARX1 I_36258 (I619028,I2683,I618550,I618542,);
not I_36259 (I619125,I2690);
DFFARX1 I_36260 (I1075714,I2683,I619125,I619151,);
not I_36261 (I619159,I619151);
nand I_36262 (I619176,I1075711,I1075720);
and I_36263 (I619193,I619176,I1075699);
DFFARX1 I_36264 (I619193,I2683,I619125,I619219,);
DFFARX1 I_36265 (I619219,I2683,I619125,I619114,);
DFFARX1 I_36266 (I1075702,I2683,I619125,I619250,);
nand I_36267 (I619258,I619250,I1075717);
not I_36268 (I619275,I619258);
DFFARX1 I_36269 (I619275,I2683,I619125,I619301,);
not I_36270 (I619309,I619301);
nor I_36271 (I619117,I619159,I619309);
DFFARX1 I_36272 (I1075723,I2683,I619125,I619349,);
nor I_36273 (I619108,I619349,I619219);
nor I_36274 (I619099,I619349,I619275);
nand I_36275 (I619385,I1075705,I1075726);
and I_36276 (I619402,I619385,I1075708);
DFFARX1 I_36277 (I619402,I2683,I619125,I619428,);
not I_36278 (I619436,I619428);
nand I_36279 (I619453,I619436,I619349);
nand I_36280 (I619102,I619436,I619258);
nor I_36281 (I619484,I1075699,I1075726);
and I_36282 (I619501,I619349,I619484);
nor I_36283 (I619518,I619436,I619501);
DFFARX1 I_36284 (I619518,I2683,I619125,I619111,);
nor I_36285 (I619549,I619151,I619484);
DFFARX1 I_36286 (I619549,I2683,I619125,I619096,);
nor I_36287 (I619580,I619428,I619484);
not I_36288 (I619597,I619580);
nand I_36289 (I619105,I619597,I619453);
not I_36290 (I619652,I2690);
DFFARX1 I_36291 (I199151,I2683,I619652,I619678,);
not I_36292 (I619686,I619678);
nand I_36293 (I619703,I199148,I199166);
and I_36294 (I619720,I619703,I199157);
DFFARX1 I_36295 (I619720,I2683,I619652,I619746,);
DFFARX1 I_36296 (I619746,I2683,I619652,I619641,);
DFFARX1 I_36297 (I199163,I2683,I619652,I619777,);
nand I_36298 (I619785,I619777,I199160);
not I_36299 (I619802,I619785);
DFFARX1 I_36300 (I619802,I2683,I619652,I619828,);
not I_36301 (I619836,I619828);
nor I_36302 (I619644,I619686,I619836);
DFFARX1 I_36303 (I199154,I2683,I619652,I619876,);
nor I_36304 (I619635,I619876,I619746);
nor I_36305 (I619626,I619876,I619802);
nand I_36306 (I619912,I199145,I199169);
and I_36307 (I619929,I619912,I199148);
DFFARX1 I_36308 (I619929,I2683,I619652,I619955,);
not I_36309 (I619963,I619955);
nand I_36310 (I619980,I619963,I619876);
nand I_36311 (I619629,I619963,I619785);
nor I_36312 (I620011,I199145,I199169);
and I_36313 (I620028,I619876,I620011);
nor I_36314 (I620045,I619963,I620028);
DFFARX1 I_36315 (I620045,I2683,I619652,I619638,);
nor I_36316 (I620076,I619678,I620011);
DFFARX1 I_36317 (I620076,I2683,I619652,I619623,);
nor I_36318 (I620107,I619955,I620011);
not I_36319 (I620124,I620107);
nand I_36320 (I619632,I620124,I619980);
not I_36321 (I620179,I2690);
DFFARX1 I_36322 (I1090589,I2683,I620179,I620205,);
not I_36323 (I620213,I620205);
nand I_36324 (I620230,I1090586,I1090595);
and I_36325 (I620247,I620230,I1090574);
DFFARX1 I_36326 (I620247,I2683,I620179,I620273,);
DFFARX1 I_36327 (I620273,I2683,I620179,I620168,);
DFFARX1 I_36328 (I1090577,I2683,I620179,I620304,);
nand I_36329 (I620312,I620304,I1090592);
not I_36330 (I620329,I620312);
DFFARX1 I_36331 (I620329,I2683,I620179,I620355,);
not I_36332 (I620363,I620355);
nor I_36333 (I620171,I620213,I620363);
DFFARX1 I_36334 (I1090598,I2683,I620179,I620403,);
nor I_36335 (I620162,I620403,I620273);
nor I_36336 (I620153,I620403,I620329);
nand I_36337 (I620439,I1090580,I1090601);
and I_36338 (I620456,I620439,I1090583);
DFFARX1 I_36339 (I620456,I2683,I620179,I620482,);
not I_36340 (I620490,I620482);
nand I_36341 (I620507,I620490,I620403);
nand I_36342 (I620156,I620490,I620312);
nor I_36343 (I620538,I1090574,I1090601);
and I_36344 (I620555,I620403,I620538);
nor I_36345 (I620572,I620490,I620555);
DFFARX1 I_36346 (I620572,I2683,I620179,I620165,);
nor I_36347 (I620603,I620205,I620538);
DFFARX1 I_36348 (I620603,I2683,I620179,I620150,);
nor I_36349 (I620634,I620482,I620538);
not I_36350 (I620651,I620634);
nand I_36351 (I620159,I620651,I620507);
not I_36352 (I620706,I2690);
DFFARX1 I_36353 (I1053699,I2683,I620706,I620732,);
not I_36354 (I620740,I620732);
nand I_36355 (I620757,I1053696,I1053705);
and I_36356 (I620774,I620757,I1053684);
DFFARX1 I_36357 (I620774,I2683,I620706,I620800,);
DFFARX1 I_36358 (I620800,I2683,I620706,I620695,);
DFFARX1 I_36359 (I1053687,I2683,I620706,I620831,);
nand I_36360 (I620839,I620831,I1053702);
not I_36361 (I620856,I620839);
DFFARX1 I_36362 (I620856,I2683,I620706,I620882,);
not I_36363 (I620890,I620882);
nor I_36364 (I620698,I620740,I620890);
DFFARX1 I_36365 (I1053708,I2683,I620706,I620930,);
nor I_36366 (I620689,I620930,I620800);
nor I_36367 (I620680,I620930,I620856);
nand I_36368 (I620966,I1053690,I1053711);
and I_36369 (I620983,I620966,I1053693);
DFFARX1 I_36370 (I620983,I2683,I620706,I621009,);
not I_36371 (I621017,I621009);
nand I_36372 (I621034,I621017,I620930);
nand I_36373 (I620683,I621017,I620839);
nor I_36374 (I621065,I1053684,I1053711);
and I_36375 (I621082,I620930,I621065);
nor I_36376 (I621099,I621017,I621082);
DFFARX1 I_36377 (I621099,I2683,I620706,I620692,);
nor I_36378 (I621130,I620732,I621065);
DFFARX1 I_36379 (I621130,I2683,I620706,I620677,);
nor I_36380 (I621161,I621009,I621065);
not I_36381 (I621178,I621161);
nand I_36382 (I620686,I621178,I621034);
not I_36383 (I621233,I2690);
DFFARX1 I_36384 (I76990,I2683,I621233,I621259,);
not I_36385 (I621267,I621259);
nand I_36386 (I621284,I76966,I76975);
and I_36387 (I621301,I621284,I76969);
DFFARX1 I_36388 (I621301,I2683,I621233,I621327,);
DFFARX1 I_36389 (I621327,I2683,I621233,I621222,);
DFFARX1 I_36390 (I76987,I2683,I621233,I621358,);
nand I_36391 (I621366,I621358,I76978);
not I_36392 (I621383,I621366);
DFFARX1 I_36393 (I621383,I2683,I621233,I621409,);
not I_36394 (I621417,I621409);
nor I_36395 (I621225,I621267,I621417);
DFFARX1 I_36396 (I76972,I2683,I621233,I621457,);
nor I_36397 (I621216,I621457,I621327);
nor I_36398 (I621207,I621457,I621383);
nand I_36399 (I621493,I76984,I76981);
and I_36400 (I621510,I621493,I76969);
DFFARX1 I_36401 (I621510,I2683,I621233,I621536,);
not I_36402 (I621544,I621536);
nand I_36403 (I621561,I621544,I621457);
nand I_36404 (I621210,I621544,I621366);
nor I_36405 (I621592,I76966,I76981);
and I_36406 (I621609,I621457,I621592);
nor I_36407 (I621626,I621544,I621609);
DFFARX1 I_36408 (I621626,I2683,I621233,I621219,);
nor I_36409 (I621657,I621259,I621592);
DFFARX1 I_36410 (I621657,I2683,I621233,I621204,);
nor I_36411 (I621688,I621536,I621592);
not I_36412 (I621705,I621688);
nand I_36413 (I621213,I621705,I621561);
not I_36414 (I621760,I2690);
DFFARX1 I_36415 (I917226,I2683,I621760,I621786,);
not I_36416 (I621794,I621786);
nand I_36417 (I621811,I917208,I917208);
and I_36418 (I621828,I621811,I917214);
DFFARX1 I_36419 (I621828,I2683,I621760,I621854,);
DFFARX1 I_36420 (I621854,I2683,I621760,I621749,);
DFFARX1 I_36421 (I917211,I2683,I621760,I621885,);
nand I_36422 (I621893,I621885,I917220);
not I_36423 (I621910,I621893);
DFFARX1 I_36424 (I621910,I2683,I621760,I621936,);
not I_36425 (I621944,I621936);
nor I_36426 (I621752,I621794,I621944);
DFFARX1 I_36427 (I917232,I2683,I621760,I621984,);
nor I_36428 (I621743,I621984,I621854);
nor I_36429 (I621734,I621984,I621910);
nand I_36430 (I622020,I917223,I917217);
and I_36431 (I622037,I622020,I917211);
DFFARX1 I_36432 (I622037,I2683,I621760,I622063,);
not I_36433 (I622071,I622063);
nand I_36434 (I622088,I622071,I621984);
nand I_36435 (I621737,I622071,I621893);
nor I_36436 (I622119,I917229,I917217);
and I_36437 (I622136,I621984,I622119);
nor I_36438 (I622153,I622071,I622136);
DFFARX1 I_36439 (I622153,I2683,I621760,I621746,);
nor I_36440 (I622184,I621786,I622119);
DFFARX1 I_36441 (I622184,I2683,I621760,I621731,);
nor I_36442 (I622215,I622063,I622119);
not I_36443 (I622232,I622215);
nand I_36444 (I621740,I622232,I622088);
not I_36445 (I622287,I2690);
DFFARX1 I_36446 (I912602,I2683,I622287,I622313,);
not I_36447 (I622321,I622313);
nand I_36448 (I622338,I912584,I912584);
and I_36449 (I622355,I622338,I912590);
DFFARX1 I_36450 (I622355,I2683,I622287,I622381,);
DFFARX1 I_36451 (I622381,I2683,I622287,I622276,);
DFFARX1 I_36452 (I912587,I2683,I622287,I622412,);
nand I_36453 (I622420,I622412,I912596);
not I_36454 (I622437,I622420);
DFFARX1 I_36455 (I622437,I2683,I622287,I622463,);
not I_36456 (I622471,I622463);
nor I_36457 (I622279,I622321,I622471);
DFFARX1 I_36458 (I912608,I2683,I622287,I622511,);
nor I_36459 (I622270,I622511,I622381);
nor I_36460 (I622261,I622511,I622437);
nand I_36461 (I622547,I912599,I912593);
and I_36462 (I622564,I622547,I912587);
DFFARX1 I_36463 (I622564,I2683,I622287,I622590,);
not I_36464 (I622598,I622590);
nand I_36465 (I622615,I622598,I622511);
nand I_36466 (I622264,I622598,I622420);
nor I_36467 (I622646,I912605,I912593);
and I_36468 (I622663,I622511,I622646);
nor I_36469 (I622680,I622598,I622663);
DFFARX1 I_36470 (I622680,I2683,I622287,I622273,);
nor I_36471 (I622711,I622313,I622646);
DFFARX1 I_36472 (I622711,I2683,I622287,I622258,);
nor I_36473 (I622742,I622590,I622646);
not I_36474 (I622759,I622742);
nand I_36475 (I622267,I622759,I622615);
not I_36476 (I622814,I2690);
DFFARX1 I_36477 (I982058,I2683,I622814,I622840,);
not I_36478 (I622848,I622840);
nand I_36479 (I622865,I982064,I982046);
and I_36480 (I622882,I622865,I982055);
DFFARX1 I_36481 (I622882,I2683,I622814,I622908,);
DFFARX1 I_36482 (I622908,I2683,I622814,I622803,);
DFFARX1 I_36483 (I982061,I2683,I622814,I622939,);
nand I_36484 (I622947,I622939,I982049);
not I_36485 (I622964,I622947);
DFFARX1 I_36486 (I622964,I2683,I622814,I622990,);
not I_36487 (I622998,I622990);
nor I_36488 (I622806,I622848,I622998);
DFFARX1 I_36489 (I982067,I2683,I622814,I623038,);
nor I_36490 (I622797,I623038,I622908);
nor I_36491 (I622788,I623038,I622964);
nand I_36492 (I623074,I982046,I982052);
and I_36493 (I623091,I623074,I982070);
DFFARX1 I_36494 (I623091,I2683,I622814,I623117,);
not I_36495 (I623125,I623117);
nand I_36496 (I623142,I623125,I623038);
nand I_36497 (I622791,I623125,I622947);
nor I_36498 (I623173,I982049,I982052);
and I_36499 (I623190,I623038,I623173);
nor I_36500 (I623207,I623125,I623190);
DFFARX1 I_36501 (I623207,I2683,I622814,I622800,);
nor I_36502 (I623238,I622840,I623173);
DFFARX1 I_36503 (I623238,I2683,I622814,I622785,);
nor I_36504 (I623269,I623117,I623173);
not I_36505 (I623286,I623269);
nand I_36506 (I622794,I623286,I623142);
not I_36507 (I623341,I2690);
DFFARX1 I_36508 (I454959,I2683,I623341,I623367,);
not I_36509 (I623375,I623367);
nand I_36510 (I623392,I454944,I454965);
and I_36511 (I623409,I623392,I454953);
DFFARX1 I_36512 (I623409,I2683,I623341,I623435,);
DFFARX1 I_36513 (I623435,I2683,I623341,I623330,);
DFFARX1 I_36514 (I454947,I2683,I623341,I623466,);
nand I_36515 (I623474,I623466,I454956);
not I_36516 (I623491,I623474);
DFFARX1 I_36517 (I623491,I2683,I623341,I623517,);
not I_36518 (I623525,I623517);
nor I_36519 (I623333,I623375,I623525);
DFFARX1 I_36520 (I454962,I2683,I623341,I623565,);
nor I_36521 (I623324,I623565,I623435);
nor I_36522 (I623315,I623565,I623491);
nand I_36523 (I623601,I454944,I454947);
and I_36524 (I623618,I623601,I454968);
DFFARX1 I_36525 (I623618,I2683,I623341,I623644,);
not I_36526 (I623652,I623644);
nand I_36527 (I623669,I623652,I623565);
nand I_36528 (I623318,I623652,I623474);
nor I_36529 (I623700,I454950,I454947);
and I_36530 (I623717,I623565,I623700);
nor I_36531 (I623734,I623652,I623717);
DFFARX1 I_36532 (I623734,I2683,I623341,I623327,);
nor I_36533 (I623765,I623367,I623700);
DFFARX1 I_36534 (I623765,I2683,I623341,I623312,);
nor I_36535 (I623796,I623644,I623700);
not I_36536 (I623813,I623796);
nand I_36537 (I623321,I623813,I623669);
not I_36538 (I623868,I2690);
DFFARX1 I_36539 (I232202,I2683,I623868,I623894,);
not I_36540 (I623902,I623894);
nand I_36541 (I623919,I232193,I232193);
and I_36542 (I623936,I623919,I232211);
DFFARX1 I_36543 (I623936,I2683,I623868,I623962,);
DFFARX1 I_36544 (I623962,I2683,I623868,I623857,);
DFFARX1 I_36545 (I232214,I2683,I623868,I623993,);
nand I_36546 (I624001,I623993,I232196);
not I_36547 (I624018,I624001);
DFFARX1 I_36548 (I624018,I2683,I623868,I624044,);
not I_36549 (I624052,I624044);
nor I_36550 (I623860,I623902,I624052);
DFFARX1 I_36551 (I232208,I2683,I623868,I624092,);
nor I_36552 (I623851,I624092,I623962);
nor I_36553 (I623842,I624092,I624018);
nand I_36554 (I624128,I232220,I232199);
and I_36555 (I624145,I624128,I232205);
DFFARX1 I_36556 (I624145,I2683,I623868,I624171,);
not I_36557 (I624179,I624171);
nand I_36558 (I624196,I624179,I624092);
nand I_36559 (I623845,I624179,I624001);
nor I_36560 (I624227,I232217,I232199);
and I_36561 (I624244,I624092,I624227);
nor I_36562 (I624261,I624179,I624244);
DFFARX1 I_36563 (I624261,I2683,I623868,I623854,);
nor I_36564 (I624292,I623894,I624227);
DFFARX1 I_36565 (I624292,I2683,I623868,I623839,);
nor I_36566 (I624323,I624171,I624227);
not I_36567 (I624340,I624323);
nand I_36568 (I623848,I624340,I624196);
not I_36569 (I624395,I2690);
DFFARX1 I_36570 (I474611,I2683,I624395,I624421,);
not I_36571 (I624429,I624421);
nand I_36572 (I624446,I474596,I474617);
and I_36573 (I624463,I624446,I474605);
DFFARX1 I_36574 (I624463,I2683,I624395,I624489,);
DFFARX1 I_36575 (I624489,I2683,I624395,I624384,);
DFFARX1 I_36576 (I474599,I2683,I624395,I624520,);
nand I_36577 (I624528,I624520,I474608);
not I_36578 (I624545,I624528);
DFFARX1 I_36579 (I624545,I2683,I624395,I624571,);
not I_36580 (I624579,I624571);
nor I_36581 (I624387,I624429,I624579);
DFFARX1 I_36582 (I474614,I2683,I624395,I624619,);
nor I_36583 (I624378,I624619,I624489);
nor I_36584 (I624369,I624619,I624545);
nand I_36585 (I624655,I474596,I474599);
and I_36586 (I624672,I624655,I474620);
DFFARX1 I_36587 (I624672,I2683,I624395,I624698,);
not I_36588 (I624706,I624698);
nand I_36589 (I624723,I624706,I624619);
nand I_36590 (I624372,I624706,I624528);
nor I_36591 (I624754,I474602,I474599);
and I_36592 (I624771,I624619,I624754);
nor I_36593 (I624788,I624706,I624771);
DFFARX1 I_36594 (I624788,I2683,I624395,I624381,);
nor I_36595 (I624819,I624421,I624754);
DFFARX1 I_36596 (I624819,I2683,I624395,I624366,);
nor I_36597 (I624850,I624698,I624754);
not I_36598 (I624867,I624850);
nand I_36599 (I624375,I624867,I624723);
not I_36600 (I624922,I2690);
DFFARX1 I_36601 (I483859,I2683,I624922,I624948,);
not I_36602 (I624956,I624948);
nand I_36603 (I624973,I483844,I483865);
and I_36604 (I624990,I624973,I483853);
DFFARX1 I_36605 (I624990,I2683,I624922,I625016,);
DFFARX1 I_36606 (I625016,I2683,I624922,I624911,);
DFFARX1 I_36607 (I483847,I2683,I624922,I625047,);
nand I_36608 (I625055,I625047,I483856);
not I_36609 (I625072,I625055);
DFFARX1 I_36610 (I625072,I2683,I624922,I625098,);
not I_36611 (I625106,I625098);
nor I_36612 (I624914,I624956,I625106);
DFFARX1 I_36613 (I483862,I2683,I624922,I625146,);
nor I_36614 (I624905,I625146,I625016);
nor I_36615 (I624896,I625146,I625072);
nand I_36616 (I625182,I483844,I483847);
and I_36617 (I625199,I625182,I483868);
DFFARX1 I_36618 (I625199,I2683,I624922,I625225,);
not I_36619 (I625233,I625225);
nand I_36620 (I625250,I625233,I625146);
nand I_36621 (I624899,I625233,I625055);
nor I_36622 (I625281,I483850,I483847);
and I_36623 (I625298,I625146,I625281);
nor I_36624 (I625315,I625233,I625298);
DFFARX1 I_36625 (I625315,I2683,I624922,I624908,);
nor I_36626 (I625346,I624948,I625281);
DFFARX1 I_36627 (I625346,I2683,I624922,I624893,);
nor I_36628 (I625377,I625225,I625281);
not I_36629 (I625394,I625377);
nand I_36630 (I624902,I625394,I625250);
not I_36631 (I625449,I2690);
DFFARX1 I_36632 (I209266,I2683,I625449,I625475,);
not I_36633 (I625483,I625475);
nand I_36634 (I625500,I209263,I209281);
and I_36635 (I625517,I625500,I209272);
DFFARX1 I_36636 (I625517,I2683,I625449,I625543,);
DFFARX1 I_36637 (I625543,I2683,I625449,I625438,);
DFFARX1 I_36638 (I209278,I2683,I625449,I625574,);
nand I_36639 (I625582,I625574,I209275);
not I_36640 (I625599,I625582);
DFFARX1 I_36641 (I625599,I2683,I625449,I625625,);
not I_36642 (I625633,I625625);
nor I_36643 (I625441,I625483,I625633);
DFFARX1 I_36644 (I209269,I2683,I625449,I625673,);
nor I_36645 (I625432,I625673,I625543);
nor I_36646 (I625423,I625673,I625599);
nand I_36647 (I625709,I209260,I209284);
and I_36648 (I625726,I625709,I209263);
DFFARX1 I_36649 (I625726,I2683,I625449,I625752,);
not I_36650 (I625760,I625752);
nand I_36651 (I625777,I625760,I625673);
nand I_36652 (I625426,I625760,I625582);
nor I_36653 (I625808,I209260,I209284);
and I_36654 (I625825,I625673,I625808);
nor I_36655 (I625842,I625760,I625825);
DFFARX1 I_36656 (I625842,I2683,I625449,I625435,);
nor I_36657 (I625873,I625475,I625808);
DFFARX1 I_36658 (I625873,I2683,I625449,I625420,);
nor I_36659 (I625904,I625752,I625808);
not I_36660 (I625921,I625904);
nand I_36661 (I625429,I625921,I625777);
not I_36662 (I625976,I2690);
DFFARX1 I_36663 (I486171,I2683,I625976,I626002,);
not I_36664 (I626010,I626002);
nand I_36665 (I626027,I486156,I486177);
and I_36666 (I626044,I626027,I486165);
DFFARX1 I_36667 (I626044,I2683,I625976,I626070,);
DFFARX1 I_36668 (I626070,I2683,I625976,I625965,);
DFFARX1 I_36669 (I486159,I2683,I625976,I626101,);
nand I_36670 (I626109,I626101,I486168);
not I_36671 (I626126,I626109);
DFFARX1 I_36672 (I626126,I2683,I625976,I626152,);
not I_36673 (I626160,I626152);
nor I_36674 (I625968,I626010,I626160);
DFFARX1 I_36675 (I486174,I2683,I625976,I626200,);
nor I_36676 (I625959,I626200,I626070);
nor I_36677 (I625950,I626200,I626126);
nand I_36678 (I626236,I486156,I486159);
and I_36679 (I626253,I626236,I486180);
DFFARX1 I_36680 (I626253,I2683,I625976,I626279,);
not I_36681 (I626287,I626279);
nand I_36682 (I626304,I626287,I626200);
nand I_36683 (I625953,I626287,I626109);
nor I_36684 (I626335,I486162,I486159);
and I_36685 (I626352,I626200,I626335);
nor I_36686 (I626369,I626287,I626352);
DFFARX1 I_36687 (I626369,I2683,I625976,I625962,);
nor I_36688 (I626400,I626002,I626335);
DFFARX1 I_36689 (I626400,I2683,I625976,I625947,);
nor I_36690 (I626431,I626279,I626335);
not I_36691 (I626448,I626431);
nand I_36692 (I625956,I626448,I626304);
not I_36693 (I626503,I2690);
DFFARX1 I_36694 (I437041,I2683,I626503,I626529,);
not I_36695 (I626537,I626529);
nand I_36696 (I626554,I437026,I437047);
and I_36697 (I626571,I626554,I437035);
DFFARX1 I_36698 (I626571,I2683,I626503,I626597,);
DFFARX1 I_36699 (I626597,I2683,I626503,I626492,);
DFFARX1 I_36700 (I437029,I2683,I626503,I626628,);
nand I_36701 (I626636,I626628,I437038);
not I_36702 (I626653,I626636);
DFFARX1 I_36703 (I626653,I2683,I626503,I626679,);
not I_36704 (I626687,I626679);
nor I_36705 (I626495,I626537,I626687);
DFFARX1 I_36706 (I437044,I2683,I626503,I626727,);
nor I_36707 (I626486,I626727,I626597);
nor I_36708 (I626477,I626727,I626653);
nand I_36709 (I626763,I437026,I437029);
and I_36710 (I626780,I626763,I437050);
DFFARX1 I_36711 (I626780,I2683,I626503,I626806,);
not I_36712 (I626814,I626806);
nand I_36713 (I626831,I626814,I626727);
nand I_36714 (I626480,I626814,I626636);
nor I_36715 (I626862,I437032,I437029);
and I_36716 (I626879,I626727,I626862);
nor I_36717 (I626896,I626814,I626879);
DFFARX1 I_36718 (I626896,I2683,I626503,I626489,);
nor I_36719 (I626927,I626529,I626862);
DFFARX1 I_36720 (I626927,I2683,I626503,I626474,);
nor I_36721 (I626958,I626806,I626862);
not I_36722 (I626975,I626958);
nand I_36723 (I626483,I626975,I626831);
not I_36724 (I627030,I2690);
DFFARX1 I_36725 (I1099514,I2683,I627030,I627056,);
not I_36726 (I627064,I627056);
nand I_36727 (I627081,I1099511,I1099520);
and I_36728 (I627098,I627081,I1099499);
DFFARX1 I_36729 (I627098,I2683,I627030,I627124,);
DFFARX1 I_36730 (I627124,I2683,I627030,I627019,);
DFFARX1 I_36731 (I1099502,I2683,I627030,I627155,);
nand I_36732 (I627163,I627155,I1099517);
not I_36733 (I627180,I627163);
DFFARX1 I_36734 (I627180,I2683,I627030,I627206,);
not I_36735 (I627214,I627206);
nor I_36736 (I627022,I627064,I627214);
DFFARX1 I_36737 (I1099523,I2683,I627030,I627254,);
nor I_36738 (I627013,I627254,I627124);
nor I_36739 (I627004,I627254,I627180);
nand I_36740 (I627290,I1099505,I1099526);
and I_36741 (I627307,I627290,I1099508);
DFFARX1 I_36742 (I627307,I2683,I627030,I627333,);
not I_36743 (I627341,I627333);
nand I_36744 (I627358,I627341,I627254);
nand I_36745 (I627007,I627341,I627163);
nor I_36746 (I627389,I1099499,I1099526);
and I_36747 (I627406,I627254,I627389);
nor I_36748 (I627423,I627341,I627406);
DFFARX1 I_36749 (I627423,I2683,I627030,I627016,);
nor I_36750 (I627454,I627056,I627389);
DFFARX1 I_36751 (I627454,I2683,I627030,I627001,);
nor I_36752 (I627485,I627333,I627389);
not I_36753 (I627502,I627485);
nand I_36754 (I627010,I627502,I627358);
not I_36755 (I627557,I2690);
DFFARX1 I_36756 (I953640,I2683,I627557,I627583,);
not I_36757 (I627591,I627583);
nand I_36758 (I627608,I953622,I953622);
and I_36759 (I627625,I627608,I953628);
DFFARX1 I_36760 (I627625,I2683,I627557,I627651,);
DFFARX1 I_36761 (I627651,I2683,I627557,I627546,);
DFFARX1 I_36762 (I953625,I2683,I627557,I627682,);
nand I_36763 (I627690,I627682,I953634);
not I_36764 (I627707,I627690);
DFFARX1 I_36765 (I627707,I2683,I627557,I627733,);
not I_36766 (I627741,I627733);
nor I_36767 (I627549,I627591,I627741);
DFFARX1 I_36768 (I953646,I2683,I627557,I627781,);
nor I_36769 (I627540,I627781,I627651);
nor I_36770 (I627531,I627781,I627707);
nand I_36771 (I627817,I953637,I953631);
and I_36772 (I627834,I627817,I953625);
DFFARX1 I_36773 (I627834,I2683,I627557,I627860,);
not I_36774 (I627868,I627860);
nand I_36775 (I627885,I627868,I627781);
nand I_36776 (I627534,I627868,I627690);
nor I_36777 (I627916,I953643,I953631);
and I_36778 (I627933,I627781,I627916);
nor I_36779 (I627950,I627868,I627933);
DFFARX1 I_36780 (I627950,I2683,I627557,I627543,);
nor I_36781 (I627981,I627583,I627916);
DFFARX1 I_36782 (I627981,I2683,I627557,I627528,);
nor I_36783 (I628012,I627860,I627916);
not I_36784 (I628029,I628012);
nand I_36785 (I627537,I628029,I627885);
not I_36786 (I628084,I2690);
DFFARX1 I_36787 (I92800,I2683,I628084,I628110,);
not I_36788 (I628118,I628110);
nand I_36789 (I628135,I92776,I92785);
and I_36790 (I628152,I628135,I92779);
DFFARX1 I_36791 (I628152,I2683,I628084,I628178,);
DFFARX1 I_36792 (I628178,I2683,I628084,I628073,);
DFFARX1 I_36793 (I92797,I2683,I628084,I628209,);
nand I_36794 (I628217,I628209,I92788);
not I_36795 (I628234,I628217);
DFFARX1 I_36796 (I628234,I2683,I628084,I628260,);
not I_36797 (I628268,I628260);
nor I_36798 (I628076,I628118,I628268);
DFFARX1 I_36799 (I92782,I2683,I628084,I628308,);
nor I_36800 (I628067,I628308,I628178);
nor I_36801 (I628058,I628308,I628234);
nand I_36802 (I628344,I92794,I92791);
and I_36803 (I628361,I628344,I92779);
DFFARX1 I_36804 (I628361,I2683,I628084,I628387,);
not I_36805 (I628395,I628387);
nand I_36806 (I628412,I628395,I628308);
nand I_36807 (I628061,I628395,I628217);
nor I_36808 (I628443,I92776,I92791);
and I_36809 (I628460,I628308,I628443);
nor I_36810 (I628477,I628395,I628460);
DFFARX1 I_36811 (I628477,I2683,I628084,I628070,);
nor I_36812 (I628508,I628110,I628443);
DFFARX1 I_36813 (I628508,I2683,I628084,I628055,);
nor I_36814 (I628539,I628387,I628443);
not I_36815 (I628556,I628539);
nand I_36816 (I628064,I628556,I628412);
not I_36817 (I628611,I2690);
DFFARX1 I_36818 (I448601,I2683,I628611,I628637,);
not I_36819 (I628645,I628637);
nand I_36820 (I628662,I448586,I448607);
and I_36821 (I628679,I628662,I448595);
DFFARX1 I_36822 (I628679,I2683,I628611,I628705,);
DFFARX1 I_36823 (I628705,I2683,I628611,I628600,);
DFFARX1 I_36824 (I448589,I2683,I628611,I628736,);
nand I_36825 (I628744,I628736,I448598);
not I_36826 (I628761,I628744);
DFFARX1 I_36827 (I628761,I2683,I628611,I628787,);
not I_36828 (I628795,I628787);
nor I_36829 (I628603,I628645,I628795);
DFFARX1 I_36830 (I448604,I2683,I628611,I628835,);
nor I_36831 (I628594,I628835,I628705);
nor I_36832 (I628585,I628835,I628761);
nand I_36833 (I628871,I448586,I448589);
and I_36834 (I628888,I628871,I448610);
DFFARX1 I_36835 (I628888,I2683,I628611,I628914,);
not I_36836 (I628922,I628914);
nand I_36837 (I628939,I628922,I628835);
nand I_36838 (I628588,I628922,I628744);
nor I_36839 (I628970,I448592,I448589);
and I_36840 (I628987,I628835,I628970);
nor I_36841 (I629004,I628922,I628987);
DFFARX1 I_36842 (I629004,I2683,I628611,I628597,);
nor I_36843 (I629035,I628637,I628970);
DFFARX1 I_36844 (I629035,I2683,I628611,I628582,);
nor I_36845 (I629066,I628914,I628970);
not I_36846 (I629083,I629066);
nand I_36847 (I628591,I629083,I628939);
not I_36848 (I629138,I2690);
DFFARX1 I_36849 (I275416,I2683,I629138,I629164,);
not I_36850 (I629172,I629164);
nand I_36851 (I629189,I275407,I275407);
and I_36852 (I629206,I629189,I275425);
DFFARX1 I_36853 (I629206,I2683,I629138,I629232,);
DFFARX1 I_36854 (I629232,I2683,I629138,I629127,);
DFFARX1 I_36855 (I275428,I2683,I629138,I629263,);
nand I_36856 (I629271,I629263,I275410);
not I_36857 (I629288,I629271);
DFFARX1 I_36858 (I629288,I2683,I629138,I629314,);
not I_36859 (I629322,I629314);
nor I_36860 (I629130,I629172,I629322);
DFFARX1 I_36861 (I275422,I2683,I629138,I629362,);
nor I_36862 (I629121,I629362,I629232);
nor I_36863 (I629112,I629362,I629288);
nand I_36864 (I629398,I275434,I275413);
and I_36865 (I629415,I629398,I275419);
DFFARX1 I_36866 (I629415,I2683,I629138,I629441,);
not I_36867 (I629449,I629441);
nand I_36868 (I629466,I629449,I629362);
nand I_36869 (I629115,I629449,I629271);
nor I_36870 (I629497,I275431,I275413);
and I_36871 (I629514,I629362,I629497);
nor I_36872 (I629531,I629449,I629514);
DFFARX1 I_36873 (I629531,I2683,I629138,I629124,);
nor I_36874 (I629562,I629164,I629497);
DFFARX1 I_36875 (I629562,I2683,I629138,I629109,);
nor I_36876 (I629593,I629441,I629497);
not I_36877 (I629610,I629593);
nand I_36878 (I629118,I629610,I629466);
not I_36879 (I629665,I2690);
DFFARX1 I_36880 (I270673,I2683,I629665,I629691,);
not I_36881 (I629699,I629691);
nand I_36882 (I629716,I270664,I270664);
and I_36883 (I629733,I629716,I270682);
DFFARX1 I_36884 (I629733,I2683,I629665,I629759,);
DFFARX1 I_36885 (I629759,I2683,I629665,I629654,);
DFFARX1 I_36886 (I270685,I2683,I629665,I629790,);
nand I_36887 (I629798,I629790,I270667);
not I_36888 (I629815,I629798);
DFFARX1 I_36889 (I629815,I2683,I629665,I629841,);
not I_36890 (I629849,I629841);
nor I_36891 (I629657,I629699,I629849);
DFFARX1 I_36892 (I270679,I2683,I629665,I629889,);
nor I_36893 (I629648,I629889,I629759);
nor I_36894 (I629639,I629889,I629815);
nand I_36895 (I629925,I270691,I270670);
and I_36896 (I629942,I629925,I270676);
DFFARX1 I_36897 (I629942,I2683,I629665,I629968,);
not I_36898 (I629976,I629968);
nand I_36899 (I629993,I629976,I629889);
nand I_36900 (I629642,I629976,I629798);
nor I_36901 (I630024,I270688,I270670);
and I_36902 (I630041,I629889,I630024);
nor I_36903 (I630058,I629976,I630041);
DFFARX1 I_36904 (I630058,I2683,I629665,I629651,);
nor I_36905 (I630089,I629691,I630024);
DFFARX1 I_36906 (I630089,I2683,I629665,I629636,);
nor I_36907 (I630120,I629968,I630024);
not I_36908 (I630137,I630120);
nand I_36909 (I629645,I630137,I629993);
not I_36910 (I630192,I2690);
DFFARX1 I_36911 (I978250,I2683,I630192,I630218,);
not I_36912 (I630226,I630218);
nand I_36913 (I630243,I978256,I978238);
and I_36914 (I630260,I630243,I978247);
DFFARX1 I_36915 (I630260,I2683,I630192,I630286,);
DFFARX1 I_36916 (I630286,I2683,I630192,I630181,);
DFFARX1 I_36917 (I978253,I2683,I630192,I630317,);
nand I_36918 (I630325,I630317,I978241);
not I_36919 (I630342,I630325);
DFFARX1 I_36920 (I630342,I2683,I630192,I630368,);
not I_36921 (I630376,I630368);
nor I_36922 (I630184,I630226,I630376);
DFFARX1 I_36923 (I978259,I2683,I630192,I630416,);
nor I_36924 (I630175,I630416,I630286);
nor I_36925 (I630166,I630416,I630342);
nand I_36926 (I630452,I978238,I978244);
and I_36927 (I630469,I630452,I978262);
DFFARX1 I_36928 (I630469,I2683,I630192,I630495,);
not I_36929 (I630503,I630495);
nand I_36930 (I630520,I630503,I630416);
nand I_36931 (I630169,I630503,I630325);
nor I_36932 (I630551,I978241,I978244);
and I_36933 (I630568,I630416,I630551);
nor I_36934 (I630585,I630503,I630568);
DFFARX1 I_36935 (I630585,I2683,I630192,I630178,);
nor I_36936 (I630616,I630218,I630551);
DFFARX1 I_36937 (I630616,I2683,I630192,I630163,);
nor I_36938 (I630647,I630495,I630551);
not I_36939 (I630664,I630647);
nand I_36940 (I630172,I630664,I630520);
not I_36941 (I630719,I2690);
DFFARX1 I_36942 (I1068574,I2683,I630719,I630745,);
not I_36943 (I630753,I630745);
nand I_36944 (I630770,I1068571,I1068580);
and I_36945 (I630787,I630770,I1068559);
DFFARX1 I_36946 (I630787,I2683,I630719,I630813,);
DFFARX1 I_36947 (I630813,I2683,I630719,I630708,);
DFFARX1 I_36948 (I1068562,I2683,I630719,I630844,);
nand I_36949 (I630852,I630844,I1068577);
not I_36950 (I630869,I630852);
DFFARX1 I_36951 (I630869,I2683,I630719,I630895,);
not I_36952 (I630903,I630895);
nor I_36953 (I630711,I630753,I630903);
DFFARX1 I_36954 (I1068583,I2683,I630719,I630943,);
nor I_36955 (I630702,I630943,I630813);
nor I_36956 (I630693,I630943,I630869);
nand I_36957 (I630979,I1068565,I1068586);
and I_36958 (I630996,I630979,I1068568);
DFFARX1 I_36959 (I630996,I2683,I630719,I631022,);
not I_36960 (I631030,I631022);
nand I_36961 (I631047,I631030,I630943);
nand I_36962 (I630696,I631030,I630852);
nor I_36963 (I631078,I1068559,I1068586);
and I_36964 (I631095,I630943,I631078);
nor I_36965 (I631112,I631030,I631095);
DFFARX1 I_36966 (I631112,I2683,I630719,I630705,);
nor I_36967 (I631143,I630745,I631078);
DFFARX1 I_36968 (I631143,I2683,I630719,I630690,);
nor I_36969 (I631174,I631022,I631078);
not I_36970 (I631191,I631174);
nand I_36971 (I630699,I631191,I631047);
not I_36972 (I631246,I2690);
DFFARX1 I_36973 (I2412,I2683,I631246,I631272,);
not I_36974 (I631280,I631272);
nand I_36975 (I631297,I1700,I1436);
and I_36976 (I631314,I631297,I1908);
DFFARX1 I_36977 (I631314,I2683,I631246,I631340,);
DFFARX1 I_36978 (I631340,I2683,I631246,I631235,);
DFFARX1 I_36979 (I1404,I2683,I631246,I631371,);
nand I_36980 (I631379,I631371,I1444);
not I_36981 (I631396,I631379);
DFFARX1 I_36982 (I631396,I2683,I631246,I631422,);
not I_36983 (I631430,I631422);
nor I_36984 (I631238,I631280,I631430);
DFFARX1 I_36985 (I2084,I2683,I631246,I631470,);
nor I_36986 (I631229,I631470,I631340);
nor I_36987 (I631220,I631470,I631396);
nand I_36988 (I631506,I2644,I2572);
and I_36989 (I631523,I631506,I2492);
DFFARX1 I_36990 (I631523,I2683,I631246,I631549,);
not I_36991 (I631557,I631549);
nand I_36992 (I631574,I631557,I631470);
nand I_36993 (I631223,I631557,I631379);
nor I_36994 (I631605,I2164,I2572);
and I_36995 (I631622,I631470,I631605);
nor I_36996 (I631639,I631557,I631622);
DFFARX1 I_36997 (I631639,I2683,I631246,I631232,);
nor I_36998 (I631670,I631272,I631605);
DFFARX1 I_36999 (I631670,I2683,I631246,I631217,);
nor I_37000 (I631701,I631549,I631605);
not I_37001 (I631718,I631701);
nand I_37002 (I631226,I631718,I631574);
not I_37003 (I631773,I2690);
DFFARX1 I_37004 (I249066,I2683,I631773,I631799,);
not I_37005 (I631807,I631799);
nand I_37006 (I631824,I249057,I249057);
and I_37007 (I631841,I631824,I249075);
DFFARX1 I_37008 (I631841,I2683,I631773,I631867,);
DFFARX1 I_37009 (I631867,I2683,I631773,I631762,);
DFFARX1 I_37010 (I249078,I2683,I631773,I631898,);
nand I_37011 (I631906,I631898,I249060);
not I_37012 (I631923,I631906);
DFFARX1 I_37013 (I631923,I2683,I631773,I631949,);
not I_37014 (I631957,I631949);
nor I_37015 (I631765,I631807,I631957);
DFFARX1 I_37016 (I249072,I2683,I631773,I631997,);
nor I_37017 (I631756,I631997,I631867);
nor I_37018 (I631747,I631997,I631923);
nand I_37019 (I632033,I249084,I249063);
and I_37020 (I632050,I632033,I249069);
DFFARX1 I_37021 (I632050,I2683,I631773,I632076,);
not I_37022 (I632084,I632076);
nand I_37023 (I632101,I632084,I631997);
nand I_37024 (I631750,I632084,I631906);
nor I_37025 (I632132,I249081,I249063);
and I_37026 (I632149,I631997,I632132);
nor I_37027 (I632166,I632084,I632149);
DFFARX1 I_37028 (I632166,I2683,I631773,I631759,);
nor I_37029 (I632197,I631799,I632132);
DFFARX1 I_37030 (I632197,I2683,I631773,I631744,);
nor I_37031 (I632228,I632076,I632132);
not I_37032 (I632245,I632228);
nand I_37033 (I631753,I632245,I632101);
not I_37034 (I632300,I2690);
DFFARX1 I_37035 (I244850,I2683,I632300,I632326,);
not I_37036 (I632334,I632326);
nand I_37037 (I632351,I244841,I244841);
and I_37038 (I632368,I632351,I244859);
DFFARX1 I_37039 (I632368,I2683,I632300,I632394,);
DFFARX1 I_37040 (I632394,I2683,I632300,I632289,);
DFFARX1 I_37041 (I244862,I2683,I632300,I632425,);
nand I_37042 (I632433,I632425,I244844);
not I_37043 (I632450,I632433);
DFFARX1 I_37044 (I632450,I2683,I632300,I632476,);
not I_37045 (I632484,I632476);
nor I_37046 (I632292,I632334,I632484);
DFFARX1 I_37047 (I244856,I2683,I632300,I632524,);
nor I_37048 (I632283,I632524,I632394);
nor I_37049 (I632274,I632524,I632450);
nand I_37050 (I632560,I244868,I244847);
and I_37051 (I632577,I632560,I244853);
DFFARX1 I_37052 (I632577,I2683,I632300,I632603,);
not I_37053 (I632611,I632603);
nand I_37054 (I632628,I632611,I632524);
nand I_37055 (I632277,I632611,I632433);
nor I_37056 (I632659,I244865,I244847);
and I_37057 (I632676,I632524,I632659);
nor I_37058 (I632693,I632611,I632676);
DFFARX1 I_37059 (I632693,I2683,I632300,I632286,);
nor I_37060 (I632724,I632326,I632659);
DFFARX1 I_37061 (I632724,I2683,I632300,I632271,);
nor I_37062 (I632755,I632603,I632659);
not I_37063 (I632772,I632755);
nand I_37064 (I632280,I632772,I632628);
not I_37065 (I632827,I2690);
DFFARX1 I_37066 (I413368,I2683,I632827,I632853,);
not I_37067 (I632861,I632853);
nand I_37068 (I632878,I413386,I413377);
and I_37069 (I632895,I632878,I413380);
DFFARX1 I_37070 (I632895,I2683,I632827,I632921,);
DFFARX1 I_37071 (I632921,I2683,I632827,I632816,);
DFFARX1 I_37072 (I413374,I2683,I632827,I632952,);
nand I_37073 (I632960,I632952,I413365);
not I_37074 (I632977,I632960);
DFFARX1 I_37075 (I632977,I2683,I632827,I633003,);
not I_37076 (I633011,I633003);
nor I_37077 (I632819,I632861,I633011);
DFFARX1 I_37078 (I413371,I2683,I632827,I633051,);
nor I_37079 (I632810,I633051,I632921);
nor I_37080 (I632801,I633051,I632977);
nand I_37081 (I633087,I413365,I413362);
and I_37082 (I633104,I633087,I413383);
DFFARX1 I_37083 (I633104,I2683,I632827,I633130,);
not I_37084 (I633138,I633130);
nand I_37085 (I633155,I633138,I633051);
nand I_37086 (I632804,I633138,I632960);
nor I_37087 (I633186,I413362,I413362);
and I_37088 (I633203,I633051,I633186);
nor I_37089 (I633220,I633138,I633203);
DFFARX1 I_37090 (I633220,I2683,I632827,I632813,);
nor I_37091 (I633251,I632853,I633186);
DFFARX1 I_37092 (I633251,I2683,I632827,I632798,);
nor I_37093 (I633282,I633130,I633186);
not I_37094 (I633299,I633282);
nand I_37095 (I632807,I633299,I633155);
not I_37096 (I633354,I2690);
DFFARX1 I_37097 (I1042989,I2683,I633354,I633380,);
not I_37098 (I633388,I633380);
nand I_37099 (I633405,I1042986,I1042995);
and I_37100 (I633422,I633405,I1042974);
DFFARX1 I_37101 (I633422,I2683,I633354,I633448,);
DFFARX1 I_37102 (I633448,I2683,I633354,I633343,);
DFFARX1 I_37103 (I1042977,I2683,I633354,I633479,);
nand I_37104 (I633487,I633479,I1042992);
not I_37105 (I633504,I633487);
DFFARX1 I_37106 (I633504,I2683,I633354,I633530,);
not I_37107 (I633538,I633530);
nor I_37108 (I633346,I633388,I633538);
DFFARX1 I_37109 (I1042998,I2683,I633354,I633578,);
nor I_37110 (I633337,I633578,I633448);
nor I_37111 (I633328,I633578,I633504);
nand I_37112 (I633614,I1042980,I1043001);
and I_37113 (I633631,I633614,I1042983);
DFFARX1 I_37114 (I633631,I2683,I633354,I633657,);
not I_37115 (I633665,I633657);
nand I_37116 (I633682,I633665,I633578);
nand I_37117 (I633331,I633665,I633487);
nor I_37118 (I633713,I1042974,I1043001);
and I_37119 (I633730,I633578,I633713);
nor I_37120 (I633747,I633665,I633730);
DFFARX1 I_37121 (I633747,I2683,I633354,I633340,);
nor I_37122 (I633778,I633380,I633713);
DFFARX1 I_37123 (I633778,I2683,I633354,I633325,);
nor I_37124 (I633809,I633657,I633713);
not I_37125 (I633826,I633809);
nand I_37126 (I633334,I633826,I633682);
not I_37127 (I633881,I2690);
DFFARX1 I_37128 (I823717,I2683,I633881,I633907,);
not I_37129 (I633915,I633907);
nand I_37130 (I633932,I823726,I823714);
and I_37131 (I633949,I633932,I823711);
DFFARX1 I_37132 (I633949,I2683,I633881,I633975,);
DFFARX1 I_37133 (I633975,I2683,I633881,I633870,);
DFFARX1 I_37134 (I823711,I2683,I633881,I634006,);
nand I_37135 (I634014,I634006,I823708);
not I_37136 (I634031,I634014);
DFFARX1 I_37137 (I634031,I2683,I633881,I634057,);
not I_37138 (I634065,I634057);
nor I_37139 (I633873,I633915,I634065);
DFFARX1 I_37140 (I823714,I2683,I633881,I634105,);
nor I_37141 (I633864,I634105,I633975);
nor I_37142 (I633855,I634105,I634031);
nand I_37143 (I634141,I823729,I823720);
and I_37144 (I634158,I634141,I823723);
DFFARX1 I_37145 (I634158,I2683,I633881,I634184,);
not I_37146 (I634192,I634184);
nand I_37147 (I634209,I634192,I634105);
nand I_37148 (I633858,I634192,I634014);
nor I_37149 (I634240,I823708,I823720);
and I_37150 (I634257,I634105,I634240);
nor I_37151 (I634274,I634192,I634257);
DFFARX1 I_37152 (I634274,I2683,I633881,I633867,);
nor I_37153 (I634305,I633907,I634240);
DFFARX1 I_37154 (I634305,I2683,I633881,I633852,);
nor I_37155 (I634336,I634184,I634240);
not I_37156 (I634353,I634336);
nand I_37157 (I633861,I634353,I634209);
not I_37158 (I634408,I2690);
DFFARX1 I_37159 (I166426,I2683,I634408,I634434,);
not I_37160 (I634442,I634434);
nand I_37161 (I634459,I166423,I166441);
and I_37162 (I634476,I634459,I166432);
DFFARX1 I_37163 (I634476,I2683,I634408,I634502,);
DFFARX1 I_37164 (I634502,I2683,I634408,I634397,);
DFFARX1 I_37165 (I166438,I2683,I634408,I634533,);
nand I_37166 (I634541,I634533,I166435);
not I_37167 (I634558,I634541);
DFFARX1 I_37168 (I634558,I2683,I634408,I634584,);
not I_37169 (I634592,I634584);
nor I_37170 (I634400,I634442,I634592);
DFFARX1 I_37171 (I166429,I2683,I634408,I634632,);
nor I_37172 (I634391,I634632,I634502);
nor I_37173 (I634382,I634632,I634558);
nand I_37174 (I634668,I166420,I166444);
and I_37175 (I634685,I634668,I166423);
DFFARX1 I_37176 (I634685,I2683,I634408,I634711,);
not I_37177 (I634719,I634711);
nand I_37178 (I634736,I634719,I634632);
nand I_37179 (I634385,I634719,I634541);
nor I_37180 (I634767,I166420,I166444);
and I_37181 (I634784,I634632,I634767);
nor I_37182 (I634801,I634719,I634784);
DFFARX1 I_37183 (I634801,I2683,I634408,I634394,);
nor I_37184 (I634832,I634434,I634767);
DFFARX1 I_37185 (I634832,I2683,I634408,I634379,);
nor I_37186 (I634863,I634711,I634767);
not I_37187 (I634880,I634863);
nand I_37188 (I634388,I634880,I634736);
not I_37189 (I634935,I2690);
DFFARX1 I_37190 (I822595,I2683,I634935,I634961,);
not I_37191 (I634969,I634961);
nand I_37192 (I634986,I822604,I822592);
and I_37193 (I635003,I634986,I822589);
DFFARX1 I_37194 (I635003,I2683,I634935,I635029,);
DFFARX1 I_37195 (I635029,I2683,I634935,I634924,);
DFFARX1 I_37196 (I822589,I2683,I634935,I635060,);
nand I_37197 (I635068,I635060,I822586);
not I_37198 (I635085,I635068);
DFFARX1 I_37199 (I635085,I2683,I634935,I635111,);
not I_37200 (I635119,I635111);
nor I_37201 (I634927,I634969,I635119);
DFFARX1 I_37202 (I822592,I2683,I634935,I635159,);
nor I_37203 (I634918,I635159,I635029);
nor I_37204 (I634909,I635159,I635085);
nand I_37205 (I635195,I822607,I822598);
and I_37206 (I635212,I635195,I822601);
DFFARX1 I_37207 (I635212,I2683,I634935,I635238,);
not I_37208 (I635246,I635238);
nand I_37209 (I635263,I635246,I635159);
nand I_37210 (I634912,I635246,I635068);
nor I_37211 (I635294,I822586,I822598);
and I_37212 (I635311,I635159,I635294);
nor I_37213 (I635328,I635246,I635311);
DFFARX1 I_37214 (I635328,I2683,I634935,I634921,);
nor I_37215 (I635359,I634961,I635294);
DFFARX1 I_37216 (I635359,I2683,I634935,I634906,);
nor I_37217 (I635390,I635238,I635294);
not I_37218 (I635407,I635390);
nand I_37219 (I634915,I635407,I635263);
not I_37220 (I635462,I2690);
DFFARX1 I_37221 (I423483,I2683,I635462,I635488,);
not I_37222 (I635496,I635488);
nand I_37223 (I635513,I423501,I423492);
and I_37224 (I635530,I635513,I423495);
DFFARX1 I_37225 (I635530,I2683,I635462,I635556,);
DFFARX1 I_37226 (I635556,I2683,I635462,I635451,);
DFFARX1 I_37227 (I423489,I2683,I635462,I635587,);
nand I_37228 (I635595,I635587,I423480);
not I_37229 (I635612,I635595);
DFFARX1 I_37230 (I635612,I2683,I635462,I635638,);
not I_37231 (I635646,I635638);
nor I_37232 (I635454,I635496,I635646);
DFFARX1 I_37233 (I423486,I2683,I635462,I635686,);
nor I_37234 (I635445,I635686,I635556);
nor I_37235 (I635436,I635686,I635612);
nand I_37236 (I635722,I423480,I423477);
and I_37237 (I635739,I635722,I423498);
DFFARX1 I_37238 (I635739,I2683,I635462,I635765,);
not I_37239 (I635773,I635765);
nand I_37240 (I635790,I635773,I635686);
nand I_37241 (I635439,I635773,I635595);
nor I_37242 (I635821,I423477,I423477);
and I_37243 (I635838,I635686,I635821);
nor I_37244 (I635855,I635773,I635838);
DFFARX1 I_37245 (I635855,I2683,I635462,I635448,);
nor I_37246 (I635886,I635488,I635821);
DFFARX1 I_37247 (I635886,I2683,I635462,I635433,);
nor I_37248 (I635917,I635765,I635821);
not I_37249 (I635934,I635917);
nand I_37250 (I635442,I635934,I635790);
not I_37251 (I635989,I2690);
DFFARX1 I_37252 (I585572,I2683,I635989,I636015,);
not I_37253 (I636023,I636015);
nand I_37254 (I636040,I585575,I585572);
and I_37255 (I636057,I636040,I585584);
DFFARX1 I_37256 (I636057,I2683,I635989,I636083,);
DFFARX1 I_37257 (I636083,I2683,I635989,I635978,);
DFFARX1 I_37258 (I585581,I2683,I635989,I636114,);
nand I_37259 (I636122,I636114,I585587);
not I_37260 (I636139,I636122);
DFFARX1 I_37261 (I636139,I2683,I635989,I636165,);
not I_37262 (I636173,I636165);
nor I_37263 (I635981,I636023,I636173);
DFFARX1 I_37264 (I585596,I2683,I635989,I636213,);
nor I_37265 (I635972,I636213,I636083);
nor I_37266 (I635963,I636213,I636139);
nand I_37267 (I636249,I585590,I585578);
and I_37268 (I636266,I636249,I585575);
DFFARX1 I_37269 (I636266,I2683,I635989,I636292,);
not I_37270 (I636300,I636292);
nand I_37271 (I636317,I636300,I636213);
nand I_37272 (I635966,I636300,I636122);
nor I_37273 (I636348,I585593,I585578);
and I_37274 (I636365,I636213,I636348);
nor I_37275 (I636382,I636300,I636365);
DFFARX1 I_37276 (I636382,I2683,I635989,I635975,);
nor I_37277 (I636413,I636015,I636348);
DFFARX1 I_37278 (I636413,I2683,I635989,I635960,);
nor I_37279 (I636444,I636292,I636348);
not I_37280 (I636461,I636444);
nand I_37281 (I635969,I636461,I636317);
not I_37282 (I636516,I2690);
DFFARX1 I_37283 (I269619,I2683,I636516,I636542,);
not I_37284 (I636550,I636542);
nand I_37285 (I636567,I269610,I269610);
and I_37286 (I636584,I636567,I269628);
DFFARX1 I_37287 (I636584,I2683,I636516,I636610,);
DFFARX1 I_37288 (I636610,I2683,I636516,I636505,);
DFFARX1 I_37289 (I269631,I2683,I636516,I636641,);
nand I_37290 (I636649,I636641,I269613);
not I_37291 (I636666,I636649);
DFFARX1 I_37292 (I636666,I2683,I636516,I636692,);
not I_37293 (I636700,I636692);
nor I_37294 (I636508,I636550,I636700);
DFFARX1 I_37295 (I269625,I2683,I636516,I636740,);
nor I_37296 (I636499,I636740,I636610);
nor I_37297 (I636490,I636740,I636666);
nand I_37298 (I636776,I269637,I269616);
and I_37299 (I636793,I636776,I269622);
DFFARX1 I_37300 (I636793,I2683,I636516,I636819,);
not I_37301 (I636827,I636819);
nand I_37302 (I636844,I636827,I636740);
nand I_37303 (I636493,I636827,I636649);
nor I_37304 (I636875,I269634,I269616);
and I_37305 (I636892,I636740,I636875);
nor I_37306 (I636909,I636827,I636892);
DFFARX1 I_37307 (I636909,I2683,I636516,I636502,);
nor I_37308 (I636940,I636542,I636875);
DFFARX1 I_37309 (I636940,I2683,I636516,I636487,);
nor I_37310 (I636971,I636819,I636875);
not I_37311 (I636988,I636971);
nand I_37312 (I636496,I636988,I636844);
not I_37313 (I637043,I2690);
DFFARX1 I_37314 (I535286,I2683,I637043,I637069,);
not I_37315 (I637077,I637069);
nand I_37316 (I637094,I535289,I535286);
and I_37317 (I637111,I637094,I535298);
DFFARX1 I_37318 (I637111,I2683,I637043,I637137,);
DFFARX1 I_37319 (I637137,I2683,I637043,I637032,);
DFFARX1 I_37320 (I535295,I2683,I637043,I637168,);
nand I_37321 (I637176,I637168,I535301);
not I_37322 (I637193,I637176);
DFFARX1 I_37323 (I637193,I2683,I637043,I637219,);
not I_37324 (I637227,I637219);
nor I_37325 (I637035,I637077,I637227);
DFFARX1 I_37326 (I535310,I2683,I637043,I637267,);
nor I_37327 (I637026,I637267,I637137);
nor I_37328 (I637017,I637267,I637193);
nand I_37329 (I637303,I535304,I535292);
and I_37330 (I637320,I637303,I535289);
DFFARX1 I_37331 (I637320,I2683,I637043,I637346,);
not I_37332 (I637354,I637346);
nand I_37333 (I637371,I637354,I637267);
nand I_37334 (I637020,I637354,I637176);
nor I_37335 (I637402,I535307,I535292);
and I_37336 (I637419,I637267,I637402);
nor I_37337 (I637436,I637354,I637419);
DFFARX1 I_37338 (I637436,I2683,I637043,I637029,);
nor I_37339 (I637467,I637069,I637402);
DFFARX1 I_37340 (I637467,I2683,I637043,I637014,);
nor I_37341 (I637498,I637346,I637402);
not I_37342 (I637515,I637498);
nand I_37343 (I637023,I637515,I637371);
not I_37344 (I637570,I2690);
DFFARX1 I_37345 (I17951,I2683,I637570,I637596,);
not I_37346 (I637604,I637596);
nand I_37347 (I637621,I17963,I17966);
and I_37348 (I637638,I637621,I17942);
DFFARX1 I_37349 (I637638,I2683,I637570,I637664,);
DFFARX1 I_37350 (I637664,I2683,I637570,I637559,);
DFFARX1 I_37351 (I17960,I2683,I637570,I637695,);
nand I_37352 (I637703,I637695,I17948);
not I_37353 (I637720,I637703);
DFFARX1 I_37354 (I637720,I2683,I637570,I637746,);
not I_37355 (I637754,I637746);
nor I_37356 (I637562,I637604,I637754);
DFFARX1 I_37357 (I17945,I2683,I637570,I637794,);
nor I_37358 (I637553,I637794,I637664);
nor I_37359 (I637544,I637794,I637720);
nand I_37360 (I637830,I17954,I17945);
and I_37361 (I637847,I637830,I17942);
DFFARX1 I_37362 (I637847,I2683,I637570,I637873,);
not I_37363 (I637881,I637873);
nand I_37364 (I637898,I637881,I637794);
nand I_37365 (I637547,I637881,I637703);
nor I_37366 (I637929,I17957,I17945);
and I_37367 (I637946,I637794,I637929);
nor I_37368 (I637963,I637881,I637946);
DFFARX1 I_37369 (I637963,I2683,I637570,I637556,);
nor I_37370 (I637994,I637596,I637929);
DFFARX1 I_37371 (I637994,I2683,I637570,I637541,);
nor I_37372 (I638025,I637873,I637929);
not I_37373 (I638042,I638025);
nand I_37374 (I637550,I638042,I637898);
not I_37375 (I638097,I2690);
DFFARX1 I_37376 (I943236,I2683,I638097,I638123,);
not I_37377 (I638131,I638123);
nand I_37378 (I638148,I943218,I943218);
and I_37379 (I638165,I638148,I943224);
DFFARX1 I_37380 (I638165,I2683,I638097,I638191,);
DFFARX1 I_37381 (I638191,I2683,I638097,I638086,);
DFFARX1 I_37382 (I943221,I2683,I638097,I638222,);
nand I_37383 (I638230,I638222,I943230);
not I_37384 (I638247,I638230);
DFFARX1 I_37385 (I638247,I2683,I638097,I638273,);
not I_37386 (I638281,I638273);
nor I_37387 (I638089,I638131,I638281);
DFFARX1 I_37388 (I943242,I2683,I638097,I638321,);
nor I_37389 (I638080,I638321,I638191);
nor I_37390 (I638071,I638321,I638247);
nand I_37391 (I638357,I943233,I943227);
and I_37392 (I638374,I638357,I943221);
DFFARX1 I_37393 (I638374,I2683,I638097,I638400,);
not I_37394 (I638408,I638400);
nand I_37395 (I638425,I638408,I638321);
nand I_37396 (I638074,I638408,I638230);
nor I_37397 (I638456,I943239,I943227);
and I_37398 (I638473,I638321,I638456);
nor I_37399 (I638490,I638408,I638473);
DFFARX1 I_37400 (I638490,I2683,I638097,I638083,);
nor I_37401 (I638521,I638123,I638456);
DFFARX1 I_37402 (I638521,I2683,I638097,I638068,);
nor I_37403 (I638552,I638400,I638456);
not I_37404 (I638569,I638552);
nand I_37405 (I638077,I638569,I638425);
not I_37406 (I638624,I2690);
DFFARX1 I_37407 (I733560,I2683,I638624,I638650,);
not I_37408 (I638658,I638650);
nand I_37409 (I638675,I733575,I733557);
and I_37410 (I638692,I638675,I733557);
DFFARX1 I_37411 (I638692,I2683,I638624,I638718,);
DFFARX1 I_37412 (I638718,I2683,I638624,I638613,);
DFFARX1 I_37413 (I733566,I2683,I638624,I638749,);
nand I_37414 (I638757,I638749,I733584);
not I_37415 (I638774,I638757);
DFFARX1 I_37416 (I638774,I2683,I638624,I638800,);
not I_37417 (I638808,I638800);
nor I_37418 (I638616,I638658,I638808);
DFFARX1 I_37419 (I733581,I2683,I638624,I638848,);
nor I_37420 (I638607,I638848,I638718);
nor I_37421 (I638598,I638848,I638774);
nand I_37422 (I638884,I733578,I733569);
and I_37423 (I638901,I638884,I733563);
DFFARX1 I_37424 (I638901,I2683,I638624,I638927,);
not I_37425 (I638935,I638927);
nand I_37426 (I638952,I638935,I638848);
nand I_37427 (I638601,I638935,I638757);
nor I_37428 (I638983,I733572,I733569);
and I_37429 (I639000,I638848,I638983);
nor I_37430 (I639017,I638935,I639000);
DFFARX1 I_37431 (I639017,I2683,I638624,I638610,);
nor I_37432 (I639048,I638650,I638983);
DFFARX1 I_37433 (I639048,I2683,I638624,I638595,);
nor I_37434 (I639079,I638927,I638983);
not I_37435 (I639096,I639079);
nand I_37436 (I638604,I639096,I638952);
not I_37437 (I639151,I2690);
DFFARX1 I_37438 (I986954,I2683,I639151,I639177,);
not I_37439 (I639185,I639177);
nand I_37440 (I639202,I986960,I986942);
and I_37441 (I639219,I639202,I986951);
DFFARX1 I_37442 (I639219,I2683,I639151,I639245,);
DFFARX1 I_37443 (I639245,I2683,I639151,I639140,);
DFFARX1 I_37444 (I986957,I2683,I639151,I639276,);
nand I_37445 (I639284,I639276,I986945);
not I_37446 (I639301,I639284);
DFFARX1 I_37447 (I639301,I2683,I639151,I639327,);
not I_37448 (I639335,I639327);
nor I_37449 (I639143,I639185,I639335);
DFFARX1 I_37450 (I986963,I2683,I639151,I639375,);
nor I_37451 (I639134,I639375,I639245);
nor I_37452 (I639125,I639375,I639301);
nand I_37453 (I639411,I986942,I986948);
and I_37454 (I639428,I639411,I986966);
DFFARX1 I_37455 (I639428,I2683,I639151,I639454,);
not I_37456 (I639462,I639454);
nand I_37457 (I639479,I639462,I639375);
nand I_37458 (I639128,I639462,I639284);
nor I_37459 (I639510,I986945,I986948);
and I_37460 (I639527,I639375,I639510);
nor I_37461 (I639544,I639462,I639527);
DFFARX1 I_37462 (I639544,I2683,I639151,I639137,);
nor I_37463 (I639575,I639177,I639510);
DFFARX1 I_37464 (I639575,I2683,I639151,I639122,);
nor I_37465 (I639606,I639454,I639510);
not I_37466 (I639623,I639606);
nand I_37467 (I639131,I639623,I639479);
not I_37468 (I639678,I2690);
DFFARX1 I_37469 (I769090,I2683,I639678,I639704,);
not I_37470 (I639712,I639704);
nand I_37471 (I639729,I769105,I769087);
and I_37472 (I639746,I639729,I769087);
DFFARX1 I_37473 (I639746,I2683,I639678,I639772,);
DFFARX1 I_37474 (I639772,I2683,I639678,I639667,);
DFFARX1 I_37475 (I769096,I2683,I639678,I639803,);
nand I_37476 (I639811,I639803,I769114);
not I_37477 (I639828,I639811);
DFFARX1 I_37478 (I639828,I2683,I639678,I639854,);
not I_37479 (I639862,I639854);
nor I_37480 (I639670,I639712,I639862);
DFFARX1 I_37481 (I769111,I2683,I639678,I639902,);
nor I_37482 (I639661,I639902,I639772);
nor I_37483 (I639652,I639902,I639828);
nand I_37484 (I639938,I769108,I769099);
and I_37485 (I639955,I639938,I769093);
DFFARX1 I_37486 (I639955,I2683,I639678,I639981,);
not I_37487 (I639989,I639981);
nand I_37488 (I640006,I639989,I639902);
nand I_37489 (I639655,I639989,I639811);
nor I_37490 (I640037,I769102,I769099);
and I_37491 (I640054,I639902,I640037);
nor I_37492 (I640071,I639989,I640054);
DFFARX1 I_37493 (I640071,I2683,I639678,I639664,);
nor I_37494 (I640102,I639704,I640037);
DFFARX1 I_37495 (I640102,I2683,I639678,I639649,);
nor I_37496 (I640133,I639981,I640037);
not I_37497 (I640150,I640133);
nand I_37498 (I639658,I640150,I640006);
not I_37499 (I640205,I2690);
DFFARX1 I_37500 (I173566,I2683,I640205,I640231,);
not I_37501 (I640239,I640231);
nand I_37502 (I640256,I173563,I173581);
and I_37503 (I640273,I640256,I173572);
DFFARX1 I_37504 (I640273,I2683,I640205,I640299,);
DFFARX1 I_37505 (I640299,I2683,I640205,I640194,);
DFFARX1 I_37506 (I173578,I2683,I640205,I640330,);
nand I_37507 (I640338,I640330,I173575);
not I_37508 (I640355,I640338);
DFFARX1 I_37509 (I640355,I2683,I640205,I640381,);
not I_37510 (I640389,I640381);
nor I_37511 (I640197,I640239,I640389);
DFFARX1 I_37512 (I173569,I2683,I640205,I640429,);
nor I_37513 (I640188,I640429,I640299);
nor I_37514 (I640179,I640429,I640355);
nand I_37515 (I640465,I173560,I173584);
and I_37516 (I640482,I640465,I173563);
DFFARX1 I_37517 (I640482,I2683,I640205,I640508,);
not I_37518 (I640516,I640508);
nand I_37519 (I640533,I640516,I640429);
nand I_37520 (I640182,I640516,I640338);
nor I_37521 (I640564,I173560,I173584);
and I_37522 (I640581,I640429,I640564);
nor I_37523 (I640598,I640516,I640581);
DFFARX1 I_37524 (I640598,I2683,I640205,I640191,);
nor I_37525 (I640629,I640231,I640564);
DFFARX1 I_37526 (I640629,I2683,I640205,I640176,);
nor I_37527 (I640660,I640508,I640564);
not I_37528 (I640677,I640660);
nand I_37529 (I640185,I640677,I640533);
not I_37530 (I640732,I2690);
DFFARX1 I_37531 (I2004,I2683,I640732,I640758,);
not I_37532 (I640766,I640758);
nand I_37533 (I640783,I2524,I1836);
and I_37534 (I640800,I640783,I2076);
DFFARX1 I_37535 (I640800,I2683,I640732,I640826,);
DFFARX1 I_37536 (I640826,I2683,I640732,I640721,);
DFFARX1 I_37537 (I2596,I2683,I640732,I640857,);
nand I_37538 (I640865,I640857,I1884);
not I_37539 (I640882,I640865);
DFFARX1 I_37540 (I640882,I2683,I640732,I640908,);
not I_37541 (I640916,I640908);
nor I_37542 (I640724,I640766,I640916);
DFFARX1 I_37543 (I2228,I2683,I640732,I640956,);
nor I_37544 (I640715,I640956,I640826);
nor I_37545 (I640706,I640956,I640882);
nand I_37546 (I640992,I1804,I2100);
and I_37547 (I641009,I640992,I2348);
DFFARX1 I_37548 (I641009,I2683,I640732,I641035,);
not I_37549 (I641043,I641035);
nand I_37550 (I641060,I641043,I640956);
nand I_37551 (I640709,I641043,I640865);
nor I_37552 (I641091,I2308,I2100);
and I_37553 (I641108,I640956,I641091);
nor I_37554 (I641125,I641043,I641108);
DFFARX1 I_37555 (I641125,I2683,I640732,I640718,);
nor I_37556 (I641156,I640758,I641091);
DFFARX1 I_37557 (I641156,I2683,I640732,I640703,);
nor I_37558 (I641187,I641035,I641091);
not I_37559 (I641204,I641187);
nand I_37560 (I640712,I641204,I641060);
not I_37561 (I641259,I2690);
DFFARX1 I_37562 (I239053,I2683,I641259,I641285,);
not I_37563 (I641293,I641285);
nand I_37564 (I641310,I239044,I239044);
and I_37565 (I641327,I641310,I239062);
DFFARX1 I_37566 (I641327,I2683,I641259,I641353,);
DFFARX1 I_37567 (I641353,I2683,I641259,I641248,);
DFFARX1 I_37568 (I239065,I2683,I641259,I641384,);
nand I_37569 (I641392,I641384,I239047);
not I_37570 (I641409,I641392);
DFFARX1 I_37571 (I641409,I2683,I641259,I641435,);
not I_37572 (I641443,I641435);
nor I_37573 (I641251,I641293,I641443);
DFFARX1 I_37574 (I239059,I2683,I641259,I641483,);
nor I_37575 (I641242,I641483,I641353);
nor I_37576 (I641233,I641483,I641409);
nand I_37577 (I641519,I239071,I239050);
and I_37578 (I641536,I641519,I239056);
DFFARX1 I_37579 (I641536,I2683,I641259,I641562,);
not I_37580 (I641570,I641562);
nand I_37581 (I641587,I641570,I641483);
nand I_37582 (I641236,I641570,I641392);
nor I_37583 (I641618,I239068,I239050);
and I_37584 (I641635,I641483,I641618);
nor I_37585 (I641652,I641570,I641635);
DFFARX1 I_37586 (I641652,I2683,I641259,I641245,);
nor I_37587 (I641683,I641285,I641618);
DFFARX1 I_37588 (I641683,I2683,I641259,I641230,);
nor I_37589 (I641714,I641562,I641618);
not I_37590 (I641731,I641714);
nand I_37591 (I641239,I641731,I641587);
not I_37592 (I641786,I2690);
DFFARX1 I_37593 (I2404,I2683,I641786,I641812,);
not I_37594 (I641820,I641812);
nand I_37595 (I641837,I2292,I1748);
and I_37596 (I641854,I641837,I2652);
DFFARX1 I_37597 (I641854,I2683,I641786,I641880,);
DFFARX1 I_37598 (I641880,I2683,I641786,I641775,);
DFFARX1 I_37599 (I1500,I2683,I641786,I641911,);
nand I_37600 (I641919,I641911,I2476);
not I_37601 (I641936,I641919);
DFFARX1 I_37602 (I641936,I2683,I641786,I641962,);
not I_37603 (I641970,I641962);
nor I_37604 (I641778,I641820,I641970);
DFFARX1 I_37605 (I1780,I2683,I641786,I642010,);
nor I_37606 (I641769,I642010,I641880);
nor I_37607 (I641760,I642010,I641936);
nand I_37608 (I642046,I2260,I2052);
and I_37609 (I642063,I642046,I2564);
DFFARX1 I_37610 (I642063,I2683,I641786,I642089,);
not I_37611 (I642097,I642089);
nand I_37612 (I642114,I642097,I642010);
nand I_37613 (I641763,I642097,I641919);
nor I_37614 (I642145,I1420,I2052);
and I_37615 (I642162,I642010,I642145);
nor I_37616 (I642179,I642097,I642162);
DFFARX1 I_37617 (I642179,I2683,I641786,I641772,);
nor I_37618 (I642210,I641812,I642145);
DFFARX1 I_37619 (I642210,I2683,I641786,I641757,);
nor I_37620 (I642241,I642089,I642145);
not I_37621 (I642258,I642241);
nand I_37622 (I641766,I642258,I642114);
not I_37623 (I642313,I2690);
DFFARX1 I_37624 (I946126,I2683,I642313,I642339,);
not I_37625 (I642347,I642339);
nand I_37626 (I642364,I946108,I946108);
and I_37627 (I642381,I642364,I946114);
DFFARX1 I_37628 (I642381,I2683,I642313,I642407,);
DFFARX1 I_37629 (I642407,I2683,I642313,I642302,);
DFFARX1 I_37630 (I946111,I2683,I642313,I642438,);
nand I_37631 (I642446,I642438,I946120);
not I_37632 (I642463,I642446);
DFFARX1 I_37633 (I642463,I2683,I642313,I642489,);
not I_37634 (I642497,I642489);
nor I_37635 (I642305,I642347,I642497);
DFFARX1 I_37636 (I946132,I2683,I642313,I642537,);
nor I_37637 (I642296,I642537,I642407);
nor I_37638 (I642287,I642537,I642463);
nand I_37639 (I642573,I946123,I946117);
and I_37640 (I642590,I642573,I946111);
DFFARX1 I_37641 (I642590,I2683,I642313,I642616,);
not I_37642 (I642624,I642616);
nand I_37643 (I642641,I642624,I642537);
nand I_37644 (I642290,I642624,I642446);
nor I_37645 (I642672,I946129,I946117);
and I_37646 (I642689,I642537,I642672);
nor I_37647 (I642706,I642624,I642689);
DFFARX1 I_37648 (I642706,I2683,I642313,I642299,);
nor I_37649 (I642737,I642339,I642672);
DFFARX1 I_37650 (I642737,I2683,I642313,I642284,);
nor I_37651 (I642768,I642616,I642672);
not I_37652 (I642785,I642768);
nand I_37653 (I642293,I642785,I642641);
not I_37654 (I642840,I2690);
DFFARX1 I_37655 (I810253,I2683,I642840,I642866,);
not I_37656 (I642874,I642866);
nand I_37657 (I642891,I810262,I810250);
and I_37658 (I642908,I642891,I810247);
DFFARX1 I_37659 (I642908,I2683,I642840,I642934,);
DFFARX1 I_37660 (I642934,I2683,I642840,I642829,);
DFFARX1 I_37661 (I810247,I2683,I642840,I642965,);
nand I_37662 (I642973,I642965,I810244);
not I_37663 (I642990,I642973);
DFFARX1 I_37664 (I642990,I2683,I642840,I643016,);
not I_37665 (I643024,I643016);
nor I_37666 (I642832,I642874,I643024);
DFFARX1 I_37667 (I810250,I2683,I642840,I643064,);
nor I_37668 (I642823,I643064,I642934);
nor I_37669 (I642814,I643064,I642990);
nand I_37670 (I643100,I810265,I810256);
and I_37671 (I643117,I643100,I810259);
DFFARX1 I_37672 (I643117,I2683,I642840,I643143,);
not I_37673 (I643151,I643143);
nand I_37674 (I643168,I643151,I643064);
nand I_37675 (I642817,I643151,I642973);
nor I_37676 (I643199,I810244,I810256);
and I_37677 (I643216,I643064,I643199);
nor I_37678 (I643233,I643151,I643216);
DFFARX1 I_37679 (I643233,I2683,I642840,I642826,);
nor I_37680 (I643264,I642866,I643199);
DFFARX1 I_37681 (I643264,I2683,I642840,I642811,);
nor I_37682 (I643295,I643143,I643199);
not I_37683 (I643312,I643295);
nand I_37684 (I642820,I643312,I643168);
not I_37685 (I643367,I2690);
DFFARX1 I_37686 (I345912,I2683,I643367,I643393,);
not I_37687 (I643401,I643393);
nand I_37688 (I643418,I345909,I345918);
and I_37689 (I643435,I643418,I345927);
DFFARX1 I_37690 (I643435,I2683,I643367,I643461,);
DFFARX1 I_37691 (I643461,I2683,I643367,I643356,);
DFFARX1 I_37692 (I345930,I2683,I643367,I643492,);
nand I_37693 (I643500,I643492,I345933);
not I_37694 (I643517,I643500);
DFFARX1 I_37695 (I643517,I2683,I643367,I643543,);
not I_37696 (I643551,I643543);
nor I_37697 (I643359,I643401,I643551);
DFFARX1 I_37698 (I345906,I2683,I643367,I643591,);
nor I_37699 (I643350,I643591,I643461);
nor I_37700 (I643341,I643591,I643517);
nand I_37701 (I643627,I345921,I345924);
and I_37702 (I643644,I643627,I345915);
DFFARX1 I_37703 (I643644,I2683,I643367,I643670,);
not I_37704 (I643678,I643670);
nand I_37705 (I643695,I643678,I643591);
nand I_37706 (I643344,I643678,I643500);
nor I_37707 (I643726,I345906,I345924);
and I_37708 (I643743,I643591,I643726);
nor I_37709 (I643760,I643678,I643743);
DFFARX1 I_37710 (I643760,I2683,I643367,I643353,);
nor I_37711 (I643791,I643393,I643726);
DFFARX1 I_37712 (I643791,I2683,I643367,I643338,);
nor I_37713 (I643822,I643670,I643726);
not I_37714 (I643839,I643822);
nand I_37715 (I643347,I643839,I643695);
not I_37716 (I643894,I2690);
DFFARX1 I_37717 (I483281,I2683,I643894,I643920,);
not I_37718 (I643928,I643920);
nand I_37719 (I643945,I483266,I483287);
and I_37720 (I643962,I643945,I483275);
DFFARX1 I_37721 (I643962,I2683,I643894,I643988,);
DFFARX1 I_37722 (I643988,I2683,I643894,I643883,);
DFFARX1 I_37723 (I483269,I2683,I643894,I644019,);
nand I_37724 (I644027,I644019,I483278);
not I_37725 (I644044,I644027);
DFFARX1 I_37726 (I644044,I2683,I643894,I644070,);
not I_37727 (I644078,I644070);
nor I_37728 (I643886,I643928,I644078);
DFFARX1 I_37729 (I483284,I2683,I643894,I644118,);
nor I_37730 (I643877,I644118,I643988);
nor I_37731 (I643868,I644118,I644044);
nand I_37732 (I644154,I483266,I483269);
and I_37733 (I644171,I644154,I483290);
DFFARX1 I_37734 (I644171,I2683,I643894,I644197,);
not I_37735 (I644205,I644197);
nand I_37736 (I644222,I644205,I644118);
nand I_37737 (I643871,I644205,I644027);
nor I_37738 (I644253,I483272,I483269);
and I_37739 (I644270,I644118,I644253);
nor I_37740 (I644287,I644205,I644270);
DFFARX1 I_37741 (I644287,I2683,I643894,I643880,);
nor I_37742 (I644318,I643920,I644253);
DFFARX1 I_37743 (I644318,I2683,I643894,I643865,);
nor I_37744 (I644349,I644197,I644253);
not I_37745 (I644366,I644349);
nand I_37746 (I643874,I644366,I644222);
not I_37747 (I644421,I2690);
DFFARX1 I_37748 (I1508,I2683,I644421,I644447,);
not I_37749 (I644455,I644447);
nand I_37750 (I644472,I1796,I1716);
and I_37751 (I644489,I644472,I2612);
DFFARX1 I_37752 (I644489,I2683,I644421,I644515,);
DFFARX1 I_37753 (I644515,I2683,I644421,I644410,);
DFFARX1 I_37754 (I2276,I2683,I644421,I644546,);
nand I_37755 (I644554,I644546,I1492);
not I_37756 (I644571,I644554);
DFFARX1 I_37757 (I644571,I2683,I644421,I644597,);
not I_37758 (I644605,I644597);
nor I_37759 (I644413,I644455,I644605);
DFFARX1 I_37760 (I1988,I2683,I644421,I644645,);
nor I_37761 (I644404,I644645,I644515);
nor I_37762 (I644395,I644645,I644571);
nand I_37763 (I644681,I1996,I1636);
and I_37764 (I644698,I644681,I2380);
DFFARX1 I_37765 (I644698,I2683,I644421,I644724,);
not I_37766 (I644732,I644724);
nand I_37767 (I644749,I644732,I644645);
nand I_37768 (I644398,I644732,I644554);
nor I_37769 (I644780,I2044,I1636);
and I_37770 (I644797,I644645,I644780);
nor I_37771 (I644814,I644732,I644797);
DFFARX1 I_37772 (I644814,I2683,I644421,I644407,);
nor I_37773 (I644845,I644447,I644780);
DFFARX1 I_37774 (I644845,I2683,I644421,I644392,);
nor I_37775 (I644876,I644724,I644780);
not I_37776 (I644893,I644876);
nand I_37777 (I644401,I644893,I644749);
not I_37778 (I644948,I2690);
DFFARX1 I_37779 (I783948,I2683,I644948,I644974,);
not I_37780 (I644982,I644974);
nand I_37781 (I644999,I783963,I783945);
and I_37782 (I645016,I644999,I783945);
DFFARX1 I_37783 (I645016,I2683,I644948,I645042,);
DFFARX1 I_37784 (I645042,I2683,I644948,I644937,);
DFFARX1 I_37785 (I783954,I2683,I644948,I645073,);
nand I_37786 (I645081,I645073,I783972);
not I_37787 (I645098,I645081);
DFFARX1 I_37788 (I645098,I2683,I644948,I645124,);
not I_37789 (I645132,I645124);
nor I_37790 (I644940,I644982,I645132);
DFFARX1 I_37791 (I783969,I2683,I644948,I645172,);
nor I_37792 (I644931,I645172,I645042);
nor I_37793 (I644922,I645172,I645098);
nand I_37794 (I645208,I783966,I783957);
and I_37795 (I645225,I645208,I783951);
DFFARX1 I_37796 (I645225,I2683,I644948,I645251,);
not I_37797 (I645259,I645251);
nand I_37798 (I645276,I645259,I645172);
nand I_37799 (I644925,I645259,I645081);
nor I_37800 (I645307,I783960,I783957);
and I_37801 (I645324,I645172,I645307);
nor I_37802 (I645341,I645259,I645324);
DFFARX1 I_37803 (I645341,I2683,I644948,I644934,);
nor I_37804 (I645372,I644974,I645307);
DFFARX1 I_37805 (I645372,I2683,I644948,I644919,);
nor I_37806 (I645403,I645251,I645307);
not I_37807 (I645420,I645403);
nand I_37808 (I644928,I645420,I645276);
not I_37809 (I645475,I2690);
DFFARX1 I_37810 (I1079284,I2683,I645475,I645501,);
not I_37811 (I645509,I645501);
nand I_37812 (I645526,I1079281,I1079290);
and I_37813 (I645543,I645526,I1079269);
DFFARX1 I_37814 (I645543,I2683,I645475,I645569,);
DFFARX1 I_37815 (I645569,I2683,I645475,I645464,);
DFFARX1 I_37816 (I1079272,I2683,I645475,I645600,);
nand I_37817 (I645608,I645600,I1079287);
not I_37818 (I645625,I645608);
DFFARX1 I_37819 (I645625,I2683,I645475,I645651,);
not I_37820 (I645659,I645651);
nor I_37821 (I645467,I645509,I645659);
DFFARX1 I_37822 (I1079293,I2683,I645475,I645699,);
nor I_37823 (I645458,I645699,I645569);
nor I_37824 (I645449,I645699,I645625);
nand I_37825 (I645735,I1079275,I1079296);
and I_37826 (I645752,I645735,I1079278);
DFFARX1 I_37827 (I645752,I2683,I645475,I645778,);
not I_37828 (I645786,I645778);
nand I_37829 (I645803,I645786,I645699);
nand I_37830 (I645452,I645786,I645608);
nor I_37831 (I645834,I1079269,I1079296);
and I_37832 (I645851,I645699,I645834);
nor I_37833 (I645868,I645786,I645851);
DFFARX1 I_37834 (I645868,I2683,I645475,I645461,);
nor I_37835 (I645899,I645501,I645834);
DFFARX1 I_37836 (I645899,I2683,I645475,I645446,);
nor I_37837 (I645930,I645778,I645834);
not I_37838 (I645947,I645930);
nand I_37839 (I645455,I645947,I645803);
not I_37840 (I646002,I2690);
DFFARX1 I_37841 (I375832,I2683,I646002,I646028,);
not I_37842 (I646036,I646028);
nand I_37843 (I646053,I375829,I375838);
and I_37844 (I646070,I646053,I375847);
DFFARX1 I_37845 (I646070,I2683,I646002,I646096,);
DFFARX1 I_37846 (I646096,I2683,I646002,I645991,);
DFFARX1 I_37847 (I375850,I2683,I646002,I646127,);
nand I_37848 (I646135,I646127,I375853);
not I_37849 (I646152,I646135);
DFFARX1 I_37850 (I646152,I2683,I646002,I646178,);
not I_37851 (I646186,I646178);
nor I_37852 (I645994,I646036,I646186);
DFFARX1 I_37853 (I375826,I2683,I646002,I646226,);
nor I_37854 (I645985,I646226,I646096);
nor I_37855 (I645976,I646226,I646152);
nand I_37856 (I646262,I375841,I375844);
and I_37857 (I646279,I646262,I375835);
DFFARX1 I_37858 (I646279,I2683,I646002,I646305,);
not I_37859 (I646313,I646305);
nand I_37860 (I646330,I646313,I646226);
nand I_37861 (I645979,I646313,I646135);
nor I_37862 (I646361,I375826,I375844);
and I_37863 (I646378,I646226,I646361);
nor I_37864 (I646395,I646313,I646378);
DFFARX1 I_37865 (I646395,I2683,I646002,I645988,);
nor I_37866 (I646426,I646028,I646361);
DFFARX1 I_37867 (I646426,I2683,I646002,I645973,);
nor I_37868 (I646457,I646305,I646361);
not I_37869 (I646474,I646457);
nand I_37870 (I645982,I646474,I646330);
not I_37871 (I646529,I2690);
DFFARX1 I_37872 (I481547,I2683,I646529,I646555,);
not I_37873 (I646563,I646555);
nand I_37874 (I646580,I481532,I481553);
and I_37875 (I646597,I646580,I481541);
DFFARX1 I_37876 (I646597,I2683,I646529,I646623,);
DFFARX1 I_37877 (I646623,I2683,I646529,I646518,);
DFFARX1 I_37878 (I481535,I2683,I646529,I646654,);
nand I_37879 (I646662,I646654,I481544);
not I_37880 (I646679,I646662);
DFFARX1 I_37881 (I646679,I2683,I646529,I646705,);
not I_37882 (I646713,I646705);
nor I_37883 (I646521,I646563,I646713);
DFFARX1 I_37884 (I481550,I2683,I646529,I646753,);
nor I_37885 (I646512,I646753,I646623);
nor I_37886 (I646503,I646753,I646679);
nand I_37887 (I646789,I481532,I481535);
and I_37888 (I646806,I646789,I481556);
DFFARX1 I_37889 (I646806,I2683,I646529,I646832,);
not I_37890 (I646840,I646832);
nand I_37891 (I646857,I646840,I646753);
nand I_37892 (I646506,I646840,I646662);
nor I_37893 (I646888,I481538,I481535);
and I_37894 (I646905,I646753,I646888);
nor I_37895 (I646922,I646840,I646905);
DFFARX1 I_37896 (I646922,I2683,I646529,I646515,);
nor I_37897 (I646953,I646555,I646888);
DFFARX1 I_37898 (I646953,I2683,I646529,I646500,);
nor I_37899 (I646984,I646832,I646888);
not I_37900 (I647001,I646984);
nand I_37901 (I646509,I647001,I646857);
not I_37902 (I647056,I2690);
DFFARX1 I_37903 (I497716,I2683,I647056,I647082,);
not I_37904 (I647090,I647082);
nand I_37905 (I647107,I497719,I497716);
and I_37906 (I647124,I647107,I497728);
DFFARX1 I_37907 (I647124,I2683,I647056,I647150,);
DFFARX1 I_37908 (I647150,I2683,I647056,I647045,);
DFFARX1 I_37909 (I497725,I2683,I647056,I647181,);
nand I_37910 (I647189,I647181,I497731);
not I_37911 (I647206,I647189);
DFFARX1 I_37912 (I647206,I2683,I647056,I647232,);
not I_37913 (I647240,I647232);
nor I_37914 (I647048,I647090,I647240);
DFFARX1 I_37915 (I497740,I2683,I647056,I647280,);
nor I_37916 (I647039,I647280,I647150);
nor I_37917 (I647030,I647280,I647206);
nand I_37918 (I647316,I497734,I497722);
and I_37919 (I647333,I647316,I497719);
DFFARX1 I_37920 (I647333,I2683,I647056,I647359,);
not I_37921 (I647367,I647359);
nand I_37922 (I647384,I647367,I647280);
nand I_37923 (I647033,I647367,I647189);
nor I_37924 (I647415,I497737,I497722);
and I_37925 (I647432,I647280,I647415);
nor I_37926 (I647449,I647367,I647432);
DFFARX1 I_37927 (I647449,I2683,I647056,I647042,);
nor I_37928 (I647480,I647082,I647415);
DFFARX1 I_37929 (I647480,I2683,I647056,I647027,);
nor I_37930 (I647511,I647359,I647415);
not I_37931 (I647528,I647511);
nand I_37932 (I647036,I647528,I647384);
not I_37933 (I647583,I2690);
DFFARX1 I_37934 (I612738,I2683,I647583,I647609,);
not I_37935 (I647617,I647609);
nand I_37936 (I647634,I612741,I612738);
and I_37937 (I647651,I647634,I612750);
DFFARX1 I_37938 (I647651,I2683,I647583,I647677,);
DFFARX1 I_37939 (I647677,I2683,I647583,I647572,);
DFFARX1 I_37940 (I612747,I2683,I647583,I647708,);
nand I_37941 (I647716,I647708,I612753);
not I_37942 (I647733,I647716);
DFFARX1 I_37943 (I647733,I2683,I647583,I647759,);
not I_37944 (I647767,I647759);
nor I_37945 (I647575,I647617,I647767);
DFFARX1 I_37946 (I612762,I2683,I647583,I647807,);
nor I_37947 (I647566,I647807,I647677);
nor I_37948 (I647557,I647807,I647733);
nand I_37949 (I647843,I612756,I612744);
and I_37950 (I647860,I647843,I612741);
DFFARX1 I_37951 (I647860,I2683,I647583,I647886,);
not I_37952 (I647894,I647886);
nand I_37953 (I647911,I647894,I647807);
nand I_37954 (I647560,I647894,I647716);
nor I_37955 (I647942,I612759,I612744);
and I_37956 (I647959,I647807,I647942);
nor I_37957 (I647976,I647894,I647959);
DFFARX1 I_37958 (I647976,I2683,I647583,I647569,);
nor I_37959 (I648007,I647609,I647942);
DFFARX1 I_37960 (I648007,I2683,I647583,I647554,);
nor I_37961 (I648038,I647886,I647942);
not I_37962 (I648055,I648038);
nand I_37963 (I647563,I648055,I647911);
not I_37964 (I648110,I2690);
DFFARX1 I_37965 (I317080,I2683,I648110,I648136,);
not I_37966 (I648144,I648136);
nand I_37967 (I648161,I317077,I317086);
and I_37968 (I648178,I648161,I317095);
DFFARX1 I_37969 (I648178,I2683,I648110,I648204,);
DFFARX1 I_37970 (I648204,I2683,I648110,I648099,);
DFFARX1 I_37971 (I317098,I2683,I648110,I648235,);
nand I_37972 (I648243,I648235,I317101);
not I_37973 (I648260,I648243);
DFFARX1 I_37974 (I648260,I2683,I648110,I648286,);
not I_37975 (I648294,I648286);
nor I_37976 (I648102,I648144,I648294);
DFFARX1 I_37977 (I317074,I2683,I648110,I648334,);
nor I_37978 (I648093,I648334,I648204);
nor I_37979 (I648084,I648334,I648260);
nand I_37980 (I648370,I317089,I317092);
and I_37981 (I648387,I648370,I317083);
DFFARX1 I_37982 (I648387,I2683,I648110,I648413,);
not I_37983 (I648421,I648413);
nand I_37984 (I648438,I648421,I648334);
nand I_37985 (I648087,I648421,I648243);
nor I_37986 (I648469,I317074,I317092);
and I_37987 (I648486,I648334,I648469);
nor I_37988 (I648503,I648421,I648486);
DFFARX1 I_37989 (I648503,I2683,I648110,I648096,);
nor I_37990 (I648534,I648136,I648469);
DFFARX1 I_37991 (I648534,I2683,I648110,I648081,);
nor I_37992 (I648565,I648413,I648469);
not I_37993 (I648582,I648565);
nand I_37994 (I648090,I648582,I648438);
not I_37995 (I648637,I2690);
DFFARX1 I_37996 (I1028241,I2683,I648637,I648663,);
not I_37997 (I648671,I648663);
nand I_37998 (I648688,I1028235,I1028253);
and I_37999 (I648705,I648688,I1028238);
DFFARX1 I_38000 (I648705,I2683,I648637,I648731,);
DFFARX1 I_38001 (I648731,I2683,I648637,I648626,);
DFFARX1 I_38002 (I1028259,I2683,I648637,I648762,);
nand I_38003 (I648770,I648762,I1028244);
not I_38004 (I648787,I648770);
DFFARX1 I_38005 (I648787,I2683,I648637,I648813,);
not I_38006 (I648821,I648813);
nor I_38007 (I648629,I648671,I648821);
DFFARX1 I_38008 (I1028256,I2683,I648637,I648861,);
nor I_38009 (I648620,I648861,I648731);
nor I_38010 (I648611,I648861,I648787);
nand I_38011 (I648897,I1028247,I1028262);
and I_38012 (I648914,I648897,I1028250);
DFFARX1 I_38013 (I648914,I2683,I648637,I648940,);
not I_38014 (I648948,I648940);
nand I_38015 (I648965,I648948,I648861);
nand I_38016 (I648614,I648948,I648770);
nor I_38017 (I648996,I1028235,I1028262);
and I_38018 (I649013,I648861,I648996);
nor I_38019 (I649030,I648948,I649013);
DFFARX1 I_38020 (I649030,I2683,I648637,I648623,);
nor I_38021 (I649061,I648663,I648996);
DFFARX1 I_38022 (I649061,I2683,I648637,I648608,);
nor I_38023 (I649092,I648940,I648996);
not I_38024 (I649109,I649092);
nand I_38025 (I648617,I649109,I648965);
not I_38026 (I649164,I2690);
DFFARX1 I_38027 (I185466,I2683,I649164,I649190,);
not I_38028 (I649198,I649190);
nand I_38029 (I649215,I185463,I185481);
and I_38030 (I649232,I649215,I185472);
DFFARX1 I_38031 (I649232,I2683,I649164,I649258,);
DFFARX1 I_38032 (I649258,I2683,I649164,I649153,);
DFFARX1 I_38033 (I185478,I2683,I649164,I649289,);
nand I_38034 (I649297,I649289,I185475);
not I_38035 (I649314,I649297);
DFFARX1 I_38036 (I649314,I2683,I649164,I649340,);
not I_38037 (I649348,I649340);
nor I_38038 (I649156,I649198,I649348);
DFFARX1 I_38039 (I185469,I2683,I649164,I649388,);
nor I_38040 (I649147,I649388,I649258);
nor I_38041 (I649138,I649388,I649314);
nand I_38042 (I649424,I185460,I185484);
and I_38043 (I649441,I649424,I185463);
DFFARX1 I_38044 (I649441,I2683,I649164,I649467,);
not I_38045 (I649475,I649467);
nand I_38046 (I649492,I649475,I649388);
nand I_38047 (I649141,I649475,I649297);
nor I_38048 (I649523,I185460,I185484);
and I_38049 (I649540,I649388,I649523);
nor I_38050 (I649557,I649475,I649540);
DFFARX1 I_38051 (I649557,I2683,I649164,I649150,);
nor I_38052 (I649588,I649190,I649523);
DFFARX1 I_38053 (I649588,I2683,I649164,I649135,);
nor I_38054 (I649619,I649467,I649523);
not I_38055 (I649636,I649619);
nand I_38056 (I649144,I649636,I649492);
not I_38057 (I649691,I2690);
DFFARX1 I_38058 (I954796,I2683,I649691,I649717,);
not I_38059 (I649725,I649717);
nand I_38060 (I649742,I954778,I954778);
and I_38061 (I649759,I649742,I954784);
DFFARX1 I_38062 (I649759,I2683,I649691,I649785,);
DFFARX1 I_38063 (I649785,I2683,I649691,I649680,);
DFFARX1 I_38064 (I954781,I2683,I649691,I649816,);
nand I_38065 (I649824,I649816,I954790);
not I_38066 (I649841,I649824);
DFFARX1 I_38067 (I649841,I2683,I649691,I649867,);
not I_38068 (I649875,I649867);
nor I_38069 (I649683,I649725,I649875);
DFFARX1 I_38070 (I954802,I2683,I649691,I649915,);
nor I_38071 (I649674,I649915,I649785);
nor I_38072 (I649665,I649915,I649841);
nand I_38073 (I649951,I954793,I954787);
and I_38074 (I649968,I649951,I954781);
DFFARX1 I_38075 (I649968,I2683,I649691,I649994,);
not I_38076 (I650002,I649994);
nand I_38077 (I650019,I650002,I649915);
nand I_38078 (I649668,I650002,I649824);
nor I_38079 (I650050,I954799,I954787);
and I_38080 (I650067,I649915,I650050);
nor I_38081 (I650084,I650002,I650067);
DFFARX1 I_38082 (I650084,I2683,I649691,I649677,);
nor I_38083 (I650115,I649717,I650050);
DFFARX1 I_38084 (I650115,I2683,I649691,I649662,);
nor I_38085 (I650146,I649994,I650050);
not I_38086 (I650163,I650146);
nand I_38087 (I649671,I650163,I650019);
not I_38088 (I650218,I2690);
DFFARX1 I_38089 (I917804,I2683,I650218,I650244,);
not I_38090 (I650252,I650244);
nand I_38091 (I650269,I917786,I917786);
and I_38092 (I650286,I650269,I917792);
DFFARX1 I_38093 (I650286,I2683,I650218,I650312,);
DFFARX1 I_38094 (I650312,I2683,I650218,I650207,);
DFFARX1 I_38095 (I917789,I2683,I650218,I650343,);
nand I_38096 (I650351,I650343,I917798);
not I_38097 (I650368,I650351);
DFFARX1 I_38098 (I650368,I2683,I650218,I650394,);
not I_38099 (I650402,I650394);
nor I_38100 (I650210,I650252,I650402);
DFFARX1 I_38101 (I917810,I2683,I650218,I650442,);
nor I_38102 (I650201,I650442,I650312);
nor I_38103 (I650192,I650442,I650368);
nand I_38104 (I650478,I917801,I917795);
and I_38105 (I650495,I650478,I917789);
DFFARX1 I_38106 (I650495,I2683,I650218,I650521,);
not I_38107 (I650529,I650521);
nand I_38108 (I650546,I650529,I650442);
nand I_38109 (I650195,I650529,I650351);
nor I_38110 (I650577,I917807,I917795);
and I_38111 (I650594,I650442,I650577);
nor I_38112 (I650611,I650529,I650594);
DFFARX1 I_38113 (I650611,I2683,I650218,I650204,);
nor I_38114 (I650642,I650244,I650577);
DFFARX1 I_38115 (I650642,I2683,I650218,I650189,);
nor I_38116 (I650673,I650521,I650577);
not I_38117 (I650690,I650673);
nand I_38118 (I650198,I650690,I650546);
not I_38119 (I650745,I2690);
DFFARX1 I_38120 (I852490,I2683,I650745,I650771,);
not I_38121 (I650779,I650771);
nand I_38122 (I650796,I852472,I852472);
and I_38123 (I650813,I650796,I852478);
DFFARX1 I_38124 (I650813,I2683,I650745,I650839,);
DFFARX1 I_38125 (I650839,I2683,I650745,I650734,);
DFFARX1 I_38126 (I852475,I2683,I650745,I650870,);
nand I_38127 (I650878,I650870,I852484);
not I_38128 (I650895,I650878);
DFFARX1 I_38129 (I650895,I2683,I650745,I650921,);
not I_38130 (I650929,I650921);
nor I_38131 (I650737,I650779,I650929);
DFFARX1 I_38132 (I852496,I2683,I650745,I650969,);
nor I_38133 (I650728,I650969,I650839);
nor I_38134 (I650719,I650969,I650895);
nand I_38135 (I651005,I852487,I852481);
and I_38136 (I651022,I651005,I852475);
DFFARX1 I_38137 (I651022,I2683,I650745,I651048,);
not I_38138 (I651056,I651048);
nand I_38139 (I651073,I651056,I650969);
nand I_38140 (I650722,I651056,I650878);
nor I_38141 (I651104,I852493,I852481);
and I_38142 (I651121,I650969,I651104);
nor I_38143 (I651138,I651056,I651121);
DFFARX1 I_38144 (I651138,I2683,I650745,I650731,);
nor I_38145 (I651169,I650771,I651104);
DFFARX1 I_38146 (I651169,I2683,I650745,I650716,);
nor I_38147 (I651200,I651048,I651104);
not I_38148 (I651217,I651200);
nand I_38149 (I650725,I651217,I651073);
not I_38150 (I651272,I2690);
DFFARX1 I_38151 (I447445,I2683,I651272,I651298,);
not I_38152 (I651306,I651298);
nand I_38153 (I651323,I447430,I447451);
and I_38154 (I651340,I651323,I447439);
DFFARX1 I_38155 (I651340,I2683,I651272,I651366,);
DFFARX1 I_38156 (I651366,I2683,I651272,I651261,);
DFFARX1 I_38157 (I447433,I2683,I651272,I651397,);
nand I_38158 (I651405,I651397,I447442);
not I_38159 (I651422,I651405);
DFFARX1 I_38160 (I651422,I2683,I651272,I651448,);
not I_38161 (I651456,I651448);
nor I_38162 (I651264,I651306,I651456);
DFFARX1 I_38163 (I447448,I2683,I651272,I651496,);
nor I_38164 (I651255,I651496,I651366);
nor I_38165 (I651246,I651496,I651422);
nand I_38166 (I651532,I447430,I447433);
and I_38167 (I651549,I651532,I447454);
DFFARX1 I_38168 (I651549,I2683,I651272,I651575,);
not I_38169 (I651583,I651575);
nand I_38170 (I651600,I651583,I651496);
nand I_38171 (I651249,I651583,I651405);
nor I_38172 (I651631,I447436,I447433);
and I_38173 (I651648,I651496,I651631);
nor I_38174 (I651665,I651583,I651648);
DFFARX1 I_38175 (I651665,I2683,I651272,I651258,);
nor I_38176 (I651696,I651298,I651631);
DFFARX1 I_38177 (I651696,I2683,I651272,I651243,);
nor I_38178 (I651727,I651575,I651631);
not I_38179 (I651744,I651727);
nand I_38180 (I651252,I651744,I651600);
not I_38181 (I651799,I2690);
DFFARX1 I_38182 (I816424,I2683,I651799,I651825,);
not I_38183 (I651833,I651825);
nand I_38184 (I651850,I816433,I816421);
and I_38185 (I651867,I651850,I816418);
DFFARX1 I_38186 (I651867,I2683,I651799,I651893,);
DFFARX1 I_38187 (I651893,I2683,I651799,I651788,);
DFFARX1 I_38188 (I816418,I2683,I651799,I651924,);
nand I_38189 (I651932,I651924,I816415);
not I_38190 (I651949,I651932);
DFFARX1 I_38191 (I651949,I2683,I651799,I651975,);
not I_38192 (I651983,I651975);
nor I_38193 (I651791,I651833,I651983);
DFFARX1 I_38194 (I816421,I2683,I651799,I652023,);
nor I_38195 (I651782,I652023,I651893);
nor I_38196 (I651773,I652023,I651949);
nand I_38197 (I652059,I816436,I816427);
and I_38198 (I652076,I652059,I816430);
DFFARX1 I_38199 (I652076,I2683,I651799,I652102,);
not I_38200 (I652110,I652102);
nand I_38201 (I652127,I652110,I652023);
nand I_38202 (I651776,I652110,I651932);
nor I_38203 (I652158,I816415,I816427);
and I_38204 (I652175,I652023,I652158);
nor I_38205 (I652192,I652110,I652175);
DFFARX1 I_38206 (I652192,I2683,I651799,I651785,);
nor I_38207 (I652223,I651825,I652158);
DFFARX1 I_38208 (I652223,I2683,I651799,I651770,);
nor I_38209 (I652254,I652102,I652158);
not I_38210 (I652271,I652254);
nand I_38211 (I651779,I652271,I652127);
not I_38212 (I652326,I2690);
DFFARX1 I_38213 (I322520,I2683,I652326,I652352,);
not I_38214 (I652360,I652352);
nand I_38215 (I652377,I322517,I322526);
and I_38216 (I652394,I652377,I322535);
DFFARX1 I_38217 (I652394,I2683,I652326,I652420,);
DFFARX1 I_38218 (I652420,I2683,I652326,I652315,);
DFFARX1 I_38219 (I322538,I2683,I652326,I652451,);
nand I_38220 (I652459,I652451,I322541);
not I_38221 (I652476,I652459);
DFFARX1 I_38222 (I652476,I2683,I652326,I652502,);
not I_38223 (I652510,I652502);
nor I_38224 (I652318,I652360,I652510);
DFFARX1 I_38225 (I322514,I2683,I652326,I652550,);
nor I_38226 (I652309,I652550,I652420);
nor I_38227 (I652300,I652550,I652476);
nand I_38228 (I652586,I322529,I322532);
and I_38229 (I652603,I652586,I322523);
DFFARX1 I_38230 (I652603,I2683,I652326,I652629,);
not I_38231 (I652637,I652629);
nand I_38232 (I652654,I652637,I652550);
nand I_38233 (I652303,I652637,I652459);
nor I_38234 (I652685,I322514,I322532);
and I_38235 (I652702,I652550,I652685);
nor I_38236 (I652719,I652637,I652702);
DFFARX1 I_38237 (I652719,I2683,I652326,I652312,);
nor I_38238 (I652750,I652352,I652685);
DFFARX1 I_38239 (I652750,I2683,I652326,I652297,);
nor I_38240 (I652781,I652629,I652685);
not I_38241 (I652798,I652781);
nand I_38242 (I652306,I652798,I652654);
not I_38243 (I652853,I2690);
DFFARX1 I_38244 (I1050129,I2683,I652853,I652879,);
not I_38245 (I652887,I652879);
nand I_38246 (I652904,I1050126,I1050135);
and I_38247 (I652921,I652904,I1050114);
DFFARX1 I_38248 (I652921,I2683,I652853,I652947,);
DFFARX1 I_38249 (I652947,I2683,I652853,I652842,);
DFFARX1 I_38250 (I1050117,I2683,I652853,I652978,);
nand I_38251 (I652986,I652978,I1050132);
not I_38252 (I653003,I652986);
DFFARX1 I_38253 (I653003,I2683,I652853,I653029,);
not I_38254 (I653037,I653029);
nor I_38255 (I652845,I652887,I653037);
DFFARX1 I_38256 (I1050138,I2683,I652853,I653077,);
nor I_38257 (I652836,I653077,I652947);
nor I_38258 (I652827,I653077,I653003);
nand I_38259 (I653113,I1050120,I1050141);
and I_38260 (I653130,I653113,I1050123);
DFFARX1 I_38261 (I653130,I2683,I652853,I653156,);
not I_38262 (I653164,I653156);
nand I_38263 (I653181,I653164,I653077);
nand I_38264 (I652830,I653164,I652986);
nor I_38265 (I653212,I1050114,I1050141);
and I_38266 (I653229,I653077,I653212);
nor I_38267 (I653246,I653164,I653229);
DFFARX1 I_38268 (I653246,I2683,I652853,I652839,);
nor I_38269 (I653277,I652879,I653212);
DFFARX1 I_38270 (I653277,I2683,I652853,I652824,);
nor I_38271 (I653308,I653156,I653212);
not I_38272 (I653325,I653308);
nand I_38273 (I652833,I653325,I653181);
not I_38274 (I653380,I2690);
DFFARX1 I_38275 (I296496,I2683,I653380,I653406,);
not I_38276 (I653414,I653406);
nand I_38277 (I653431,I296487,I296487);
and I_38278 (I653448,I653431,I296505);
DFFARX1 I_38279 (I653448,I2683,I653380,I653474,);
DFFARX1 I_38280 (I653474,I2683,I653380,I653369,);
DFFARX1 I_38281 (I296508,I2683,I653380,I653505,);
nand I_38282 (I653513,I653505,I296490);
not I_38283 (I653530,I653513);
DFFARX1 I_38284 (I653530,I2683,I653380,I653556,);
not I_38285 (I653564,I653556);
nor I_38286 (I653372,I653414,I653564);
DFFARX1 I_38287 (I296502,I2683,I653380,I653604,);
nor I_38288 (I653363,I653604,I653474);
nor I_38289 (I653354,I653604,I653530);
nand I_38290 (I653640,I296514,I296493);
and I_38291 (I653657,I653640,I296499);
DFFARX1 I_38292 (I653657,I2683,I653380,I653683,);
not I_38293 (I653691,I653683);
nand I_38294 (I653708,I653691,I653604);
nand I_38295 (I653357,I653691,I653513);
nor I_38296 (I653739,I296511,I296493);
and I_38297 (I653756,I653604,I653739);
nor I_38298 (I653773,I653691,I653756);
DFFARX1 I_38299 (I653773,I2683,I653380,I653366,);
nor I_38300 (I653804,I653406,I653739);
DFFARX1 I_38301 (I653804,I2683,I653380,I653351,);
nor I_38302 (I653835,I653683,I653739);
not I_38303 (I653852,I653835);
nand I_38304 (I653360,I653852,I653708);
not I_38305 (I653907,I2690);
DFFARX1 I_38306 (I162261,I2683,I653907,I653933,);
not I_38307 (I653941,I653933);
nand I_38308 (I653958,I162258,I162276);
and I_38309 (I653975,I653958,I162267);
DFFARX1 I_38310 (I653975,I2683,I653907,I654001,);
DFFARX1 I_38311 (I654001,I2683,I653907,I653896,);
DFFARX1 I_38312 (I162273,I2683,I653907,I654032,);
nand I_38313 (I654040,I654032,I162270);
not I_38314 (I654057,I654040);
DFFARX1 I_38315 (I654057,I2683,I653907,I654083,);
not I_38316 (I654091,I654083);
nor I_38317 (I653899,I653941,I654091);
DFFARX1 I_38318 (I162264,I2683,I653907,I654131,);
nor I_38319 (I653890,I654131,I654001);
nor I_38320 (I653881,I654131,I654057);
nand I_38321 (I654167,I162255,I162279);
and I_38322 (I654184,I654167,I162258);
DFFARX1 I_38323 (I654184,I2683,I653907,I654210,);
not I_38324 (I654218,I654210);
nand I_38325 (I654235,I654218,I654131);
nand I_38326 (I653884,I654218,I654040);
nor I_38327 (I654266,I162255,I162279);
and I_38328 (I654283,I654131,I654266);
nor I_38329 (I654300,I654218,I654283);
DFFARX1 I_38330 (I654300,I2683,I653907,I653893,);
nor I_38331 (I654331,I653933,I654266);
DFFARX1 I_38332 (I654331,I2683,I653907,I653878,);
nor I_38333 (I654362,I654210,I654266);
not I_38334 (I654379,I654362);
nand I_38335 (I653887,I654379,I654235);
not I_38336 (I654434,I2690);
DFFARX1 I_38337 (I189631,I2683,I654434,I654460,);
not I_38338 (I654468,I654460);
nand I_38339 (I654485,I189628,I189646);
and I_38340 (I654502,I654485,I189637);
DFFARX1 I_38341 (I654502,I2683,I654434,I654528,);
DFFARX1 I_38342 (I654528,I2683,I654434,I654423,);
DFFARX1 I_38343 (I189643,I2683,I654434,I654559,);
nand I_38344 (I654567,I654559,I189640);
not I_38345 (I654584,I654567);
DFFARX1 I_38346 (I654584,I2683,I654434,I654610,);
not I_38347 (I654618,I654610);
nor I_38348 (I654426,I654468,I654618);
DFFARX1 I_38349 (I189634,I2683,I654434,I654658,);
nor I_38350 (I654417,I654658,I654528);
nor I_38351 (I654408,I654658,I654584);
nand I_38352 (I654694,I189625,I189649);
and I_38353 (I654711,I654694,I189628);
DFFARX1 I_38354 (I654711,I2683,I654434,I654737,);
not I_38355 (I654745,I654737);
nand I_38356 (I654762,I654745,I654658);
nand I_38357 (I654411,I654745,I654567);
nor I_38358 (I654793,I189625,I189649);
and I_38359 (I654810,I654658,I654793);
nor I_38360 (I654827,I654745,I654810);
DFFARX1 I_38361 (I654827,I2683,I654434,I654420,);
nor I_38362 (I654858,I654460,I654793);
DFFARX1 I_38363 (I654858,I2683,I654434,I654405,);
nor I_38364 (I654889,I654737,I654793);
not I_38365 (I654906,I654889);
nand I_38366 (I654414,I654906,I654762);
not I_38367 (I654961,I2690);
DFFARX1 I_38368 (I39558,I2683,I654961,I654987,);
not I_38369 (I654995,I654987);
nand I_38370 (I655012,I39570,I39573);
and I_38371 (I655029,I655012,I39549);
DFFARX1 I_38372 (I655029,I2683,I654961,I655055,);
DFFARX1 I_38373 (I655055,I2683,I654961,I654950,);
DFFARX1 I_38374 (I39567,I2683,I654961,I655086,);
nand I_38375 (I655094,I655086,I39555);
not I_38376 (I655111,I655094);
DFFARX1 I_38377 (I655111,I2683,I654961,I655137,);
not I_38378 (I655145,I655137);
nor I_38379 (I654953,I654995,I655145);
DFFARX1 I_38380 (I39552,I2683,I654961,I655185,);
nor I_38381 (I654944,I655185,I655055);
nor I_38382 (I654935,I655185,I655111);
nand I_38383 (I655221,I39561,I39552);
and I_38384 (I655238,I655221,I39549);
DFFARX1 I_38385 (I655238,I2683,I654961,I655264,);
not I_38386 (I655272,I655264);
nand I_38387 (I655289,I655272,I655185);
nand I_38388 (I654938,I655272,I655094);
nor I_38389 (I655320,I39564,I39552);
and I_38390 (I655337,I655185,I655320);
nor I_38391 (I655354,I655272,I655337);
DFFARX1 I_38392 (I655354,I2683,I654961,I654947,);
nor I_38393 (I655385,I654987,I655320);
DFFARX1 I_38394 (I655385,I2683,I654961,I654932,);
nor I_38395 (I655416,I655264,I655320);
not I_38396 (I655433,I655416);
nand I_38397 (I654941,I655433,I655289);
not I_38398 (I655488,I2690);
DFFARX1 I_38399 (I1011712,I2683,I655488,I655514,);
not I_38400 (I655522,I655514);
nand I_38401 (I655539,I1011694,I1011697);
and I_38402 (I655556,I655539,I1011709);
DFFARX1 I_38403 (I655556,I2683,I655488,I655582,);
DFFARX1 I_38404 (I655582,I2683,I655488,I655477,);
DFFARX1 I_38405 (I1011718,I2683,I655488,I655613,);
nand I_38406 (I655621,I655613,I1011703);
not I_38407 (I655638,I655621);
DFFARX1 I_38408 (I655638,I2683,I655488,I655664,);
not I_38409 (I655672,I655664);
nor I_38410 (I655480,I655522,I655672);
DFFARX1 I_38411 (I1011715,I2683,I655488,I655712,);
nor I_38412 (I655471,I655712,I655582);
nor I_38413 (I655462,I655712,I655638);
nand I_38414 (I655748,I1011706,I1011700);
and I_38415 (I655765,I655748,I1011694);
DFFARX1 I_38416 (I655765,I2683,I655488,I655791,);
not I_38417 (I655799,I655791);
nand I_38418 (I655816,I655799,I655712);
nand I_38419 (I655465,I655799,I655621);
nor I_38420 (I655847,I1011697,I1011700);
and I_38421 (I655864,I655712,I655847);
nor I_38422 (I655881,I655799,I655864);
DFFARX1 I_38423 (I655881,I2683,I655488,I655474,);
nor I_38424 (I655912,I655514,I655847);
DFFARX1 I_38425 (I655912,I2683,I655488,I655459,);
nor I_38426 (I655943,I655791,I655847);
not I_38427 (I655960,I655943);
nand I_38428 (I655468,I655960,I655816);
not I_38429 (I656015,I2690);
DFFARX1 I_38430 (I192011,I2683,I656015,I656041,);
not I_38431 (I656049,I656041);
nand I_38432 (I656066,I192008,I192026);
and I_38433 (I656083,I656066,I192017);
DFFARX1 I_38434 (I656083,I2683,I656015,I656109,);
DFFARX1 I_38435 (I656109,I2683,I656015,I656004,);
DFFARX1 I_38436 (I192023,I2683,I656015,I656140,);
nand I_38437 (I656148,I656140,I192020);
not I_38438 (I656165,I656148);
DFFARX1 I_38439 (I656165,I2683,I656015,I656191,);
not I_38440 (I656199,I656191);
nor I_38441 (I656007,I656049,I656199);
DFFARX1 I_38442 (I192014,I2683,I656015,I656239,);
nor I_38443 (I655998,I656239,I656109);
nor I_38444 (I655989,I656239,I656165);
nand I_38445 (I656275,I192005,I192029);
and I_38446 (I656292,I656275,I192008);
DFFARX1 I_38447 (I656292,I2683,I656015,I656318,);
not I_38448 (I656326,I656318);
nand I_38449 (I656343,I656326,I656239);
nand I_38450 (I655992,I656326,I656148);
nor I_38451 (I656374,I192005,I192029);
and I_38452 (I656391,I656239,I656374);
nor I_38453 (I656408,I656326,I656391);
DFFARX1 I_38454 (I656408,I2683,I656015,I656001,);
nor I_38455 (I656439,I656041,I656374);
DFFARX1 I_38456 (I656439,I2683,I656015,I655986,);
nor I_38457 (I656470,I656318,I656374);
not I_38458 (I656487,I656470);
nand I_38459 (I655995,I656487,I656343);
not I_38460 (I656542,I2690);
DFFARX1 I_38461 (I840930,I2683,I656542,I656568,);
not I_38462 (I656576,I656568);
nand I_38463 (I656593,I840912,I840912);
and I_38464 (I656610,I656593,I840918);
DFFARX1 I_38465 (I656610,I2683,I656542,I656636,);
DFFARX1 I_38466 (I656636,I2683,I656542,I656531,);
DFFARX1 I_38467 (I840915,I2683,I656542,I656667,);
nand I_38468 (I656675,I656667,I840924);
not I_38469 (I656692,I656675);
DFFARX1 I_38470 (I656692,I2683,I656542,I656718,);
not I_38471 (I656726,I656718);
nor I_38472 (I656534,I656576,I656726);
DFFARX1 I_38473 (I840936,I2683,I656542,I656766,);
nor I_38474 (I656525,I656766,I656636);
nor I_38475 (I656516,I656766,I656692);
nand I_38476 (I656802,I840927,I840921);
and I_38477 (I656819,I656802,I840915);
DFFARX1 I_38478 (I656819,I2683,I656542,I656845,);
not I_38479 (I656853,I656845);
nand I_38480 (I656870,I656853,I656766);
nand I_38481 (I656519,I656853,I656675);
nor I_38482 (I656901,I840933,I840921);
and I_38483 (I656918,I656766,I656901);
nor I_38484 (I656935,I656853,I656918);
DFFARX1 I_38485 (I656935,I2683,I656542,I656528,);
nor I_38486 (I656966,I656568,I656901);
DFFARX1 I_38487 (I656966,I2683,I656542,I656513,);
nor I_38488 (I656997,I656845,I656901);
not I_38489 (I657014,I656997);
nand I_38490 (I656522,I657014,I656870);
not I_38491 (I657069,I2690);
DFFARX1 I_38492 (I302820,I2683,I657069,I657095,);
not I_38493 (I657103,I657095);
nand I_38494 (I657120,I302811,I302811);
and I_38495 (I657137,I657120,I302829);
DFFARX1 I_38496 (I657137,I2683,I657069,I657163,);
DFFARX1 I_38497 (I657163,I2683,I657069,I657058,);
DFFARX1 I_38498 (I302832,I2683,I657069,I657194,);
nand I_38499 (I657202,I657194,I302814);
not I_38500 (I657219,I657202);
DFFARX1 I_38501 (I657219,I2683,I657069,I657245,);
not I_38502 (I657253,I657245);
nor I_38503 (I657061,I657103,I657253);
DFFARX1 I_38504 (I302826,I2683,I657069,I657293,);
nor I_38505 (I657052,I657293,I657163);
nor I_38506 (I657043,I657293,I657219);
nand I_38507 (I657329,I302838,I302817);
and I_38508 (I657346,I657329,I302823);
DFFARX1 I_38509 (I657346,I2683,I657069,I657372,);
not I_38510 (I657380,I657372);
nand I_38511 (I657397,I657380,I657293);
nand I_38512 (I657046,I657380,I657202);
nor I_38513 (I657428,I302835,I302817);
and I_38514 (I657445,I657293,I657428);
nor I_38515 (I657462,I657380,I657445);
DFFARX1 I_38516 (I657462,I2683,I657069,I657055,);
nor I_38517 (I657493,I657095,I657428);
DFFARX1 I_38518 (I657493,I2683,I657069,I657040,);
nor I_38519 (I657524,I657372,I657428);
not I_38520 (I657541,I657524);
nand I_38521 (I657049,I657541,I657397);
not I_38522 (I657596,I2690);
DFFARX1 I_38523 (I42720,I2683,I657596,I657622,);
not I_38524 (I657630,I657622);
nand I_38525 (I657647,I42732,I42735);
and I_38526 (I657664,I657647,I42711);
DFFARX1 I_38527 (I657664,I2683,I657596,I657690,);
DFFARX1 I_38528 (I657690,I2683,I657596,I657585,);
DFFARX1 I_38529 (I42729,I2683,I657596,I657721,);
nand I_38530 (I657729,I657721,I42717);
not I_38531 (I657746,I657729);
DFFARX1 I_38532 (I657746,I2683,I657596,I657772,);
not I_38533 (I657780,I657772);
nor I_38534 (I657588,I657630,I657780);
DFFARX1 I_38535 (I42714,I2683,I657596,I657820,);
nor I_38536 (I657579,I657820,I657690);
nor I_38537 (I657570,I657820,I657746);
nand I_38538 (I657856,I42723,I42714);
and I_38539 (I657873,I657856,I42711);
DFFARX1 I_38540 (I657873,I2683,I657596,I657899,);
not I_38541 (I657907,I657899);
nand I_38542 (I657924,I657907,I657820);
nand I_38543 (I657573,I657907,I657729);
nor I_38544 (I657955,I42726,I42714);
and I_38545 (I657972,I657820,I657955);
nor I_38546 (I657989,I657907,I657972);
DFFARX1 I_38547 (I657989,I2683,I657596,I657582,);
nor I_38548 (I658020,I657622,I657955);
DFFARX1 I_38549 (I658020,I2683,I657596,I657567,);
nor I_38550 (I658051,I657899,I657955);
not I_38551 (I658068,I658051);
nand I_38552 (I657576,I658068,I657924);
not I_38553 (I658123,I2690);
DFFARX1 I_38554 (I16370,I2683,I658123,I658149,);
not I_38555 (I658157,I658149);
nand I_38556 (I658174,I16382,I16385);
and I_38557 (I658191,I658174,I16361);
DFFARX1 I_38558 (I658191,I2683,I658123,I658217,);
DFFARX1 I_38559 (I658217,I2683,I658123,I658112,);
DFFARX1 I_38560 (I16379,I2683,I658123,I658248,);
nand I_38561 (I658256,I658248,I16367);
not I_38562 (I658273,I658256);
DFFARX1 I_38563 (I658273,I2683,I658123,I658299,);
not I_38564 (I658307,I658299);
nor I_38565 (I658115,I658157,I658307);
DFFARX1 I_38566 (I16364,I2683,I658123,I658347,);
nor I_38567 (I658106,I658347,I658217);
nor I_38568 (I658097,I658347,I658273);
nand I_38569 (I658383,I16373,I16364);
and I_38570 (I658400,I658383,I16361);
DFFARX1 I_38571 (I658400,I2683,I658123,I658426,);
not I_38572 (I658434,I658426);
nand I_38573 (I658451,I658434,I658347);
nand I_38574 (I658100,I658434,I658256);
nor I_38575 (I658482,I16376,I16364);
and I_38576 (I658499,I658347,I658482);
nor I_38577 (I658516,I658434,I658499);
DFFARX1 I_38578 (I658516,I2683,I658123,I658109,);
nor I_38579 (I658547,I658149,I658482);
DFFARX1 I_38580 (I658547,I2683,I658123,I658094,);
nor I_38581 (I658578,I658426,I658482);
not I_38582 (I658595,I658578);
nand I_38583 (I658103,I658595,I658451);
not I_38584 (I658650,I2690);
DFFARX1 I_38585 (I67504,I2683,I658650,I658676,);
not I_38586 (I658684,I658676);
nand I_38587 (I658701,I67480,I67489);
and I_38588 (I658718,I658701,I67483);
DFFARX1 I_38589 (I658718,I2683,I658650,I658744,);
DFFARX1 I_38590 (I658744,I2683,I658650,I658639,);
DFFARX1 I_38591 (I67501,I2683,I658650,I658775,);
nand I_38592 (I658783,I658775,I67492);
not I_38593 (I658800,I658783);
DFFARX1 I_38594 (I658800,I2683,I658650,I658826,);
not I_38595 (I658834,I658826);
nor I_38596 (I658642,I658684,I658834);
DFFARX1 I_38597 (I67486,I2683,I658650,I658874,);
nor I_38598 (I658633,I658874,I658744);
nor I_38599 (I658624,I658874,I658800);
nand I_38600 (I658910,I67498,I67495);
and I_38601 (I658927,I658910,I67483);
DFFARX1 I_38602 (I658927,I2683,I658650,I658953,);
not I_38603 (I658961,I658953);
nand I_38604 (I658978,I658961,I658874);
nand I_38605 (I658627,I658961,I658783);
nor I_38606 (I659009,I67480,I67495);
and I_38607 (I659026,I658874,I659009);
nor I_38608 (I659043,I658961,I659026);
DFFARX1 I_38609 (I659043,I2683,I658650,I658636,);
nor I_38610 (I659074,I658676,I659009);
DFFARX1 I_38611 (I659074,I2683,I658650,I658621,);
nor I_38612 (I659105,I658953,I659009);
not I_38613 (I659122,I659105);
nand I_38614 (I658630,I659122,I658978);
not I_38615 (I659177,I2690);
DFFARX1 I_38616 (I1051319,I2683,I659177,I659203,);
not I_38617 (I659211,I659203);
nand I_38618 (I659228,I1051316,I1051325);
and I_38619 (I659245,I659228,I1051304);
DFFARX1 I_38620 (I659245,I2683,I659177,I659271,);
DFFARX1 I_38621 (I659271,I2683,I659177,I659166,);
DFFARX1 I_38622 (I1051307,I2683,I659177,I659302,);
nand I_38623 (I659310,I659302,I1051322);
not I_38624 (I659327,I659310);
DFFARX1 I_38625 (I659327,I2683,I659177,I659353,);
not I_38626 (I659361,I659353);
nor I_38627 (I659169,I659211,I659361);
DFFARX1 I_38628 (I1051328,I2683,I659177,I659401,);
nor I_38629 (I659160,I659401,I659271);
nor I_38630 (I659151,I659401,I659327);
nand I_38631 (I659437,I1051310,I1051331);
and I_38632 (I659454,I659437,I1051313);
DFFARX1 I_38633 (I659454,I2683,I659177,I659480,);
not I_38634 (I659488,I659480);
nand I_38635 (I659505,I659488,I659401);
nand I_38636 (I659154,I659488,I659310);
nor I_38637 (I659536,I1051304,I1051331);
and I_38638 (I659553,I659401,I659536);
nor I_38639 (I659570,I659488,I659553);
DFFARX1 I_38640 (I659570,I2683,I659177,I659163,);
nor I_38641 (I659601,I659203,I659536);
DFFARX1 I_38642 (I659601,I2683,I659177,I659148,);
nor I_38643 (I659632,I659480,I659536);
not I_38644 (I659649,I659632);
nand I_38645 (I659157,I659649,I659505);
not I_38646 (I659704,I2690);
DFFARX1 I_38647 (I260660,I2683,I659704,I659730,);
not I_38648 (I659738,I659730);
nand I_38649 (I659755,I260651,I260651);
and I_38650 (I659772,I659755,I260669);
DFFARX1 I_38651 (I659772,I2683,I659704,I659798,);
DFFARX1 I_38652 (I659798,I2683,I659704,I659693,);
DFFARX1 I_38653 (I260672,I2683,I659704,I659829,);
nand I_38654 (I659837,I659829,I260654);
not I_38655 (I659854,I659837);
DFFARX1 I_38656 (I659854,I2683,I659704,I659880,);
not I_38657 (I659888,I659880);
nor I_38658 (I659696,I659738,I659888);
DFFARX1 I_38659 (I260666,I2683,I659704,I659928,);
nor I_38660 (I659687,I659928,I659798);
nor I_38661 (I659678,I659928,I659854);
nand I_38662 (I659964,I260678,I260657);
and I_38663 (I659981,I659964,I260663);
DFFARX1 I_38664 (I659981,I2683,I659704,I660007,);
not I_38665 (I660015,I660007);
nand I_38666 (I660032,I660015,I659928);
nand I_38667 (I659681,I660015,I659837);
nor I_38668 (I660063,I260675,I260657);
and I_38669 (I660080,I659928,I660063);
nor I_38670 (I660097,I660015,I660080);
DFFARX1 I_38671 (I660097,I2683,I659704,I659690,);
nor I_38672 (I660128,I659730,I660063);
DFFARX1 I_38673 (I660128,I2683,I659704,I659675,);
nor I_38674 (I660159,I660007,I660063);
not I_38675 (I660176,I660159);
nand I_38676 (I659684,I660176,I660032);
not I_38677 (I660231,I2690);
DFFARX1 I_38678 (I906822,I2683,I660231,I660257,);
not I_38679 (I660265,I660257);
nand I_38680 (I660282,I906804,I906804);
and I_38681 (I660299,I660282,I906810);
DFFARX1 I_38682 (I660299,I2683,I660231,I660325,);
DFFARX1 I_38683 (I660325,I2683,I660231,I660220,);
DFFARX1 I_38684 (I906807,I2683,I660231,I660356,);
nand I_38685 (I660364,I660356,I906816);
not I_38686 (I660381,I660364);
DFFARX1 I_38687 (I660381,I2683,I660231,I660407,);
not I_38688 (I660415,I660407);
nor I_38689 (I660223,I660265,I660415);
DFFARX1 I_38690 (I906828,I2683,I660231,I660455,);
nor I_38691 (I660214,I660455,I660325);
nor I_38692 (I660205,I660455,I660381);
nand I_38693 (I660491,I906819,I906813);
and I_38694 (I660508,I660491,I906807);
DFFARX1 I_38695 (I660508,I2683,I660231,I660534,);
not I_38696 (I660542,I660534);
nand I_38697 (I660559,I660542,I660455);
nand I_38698 (I660208,I660542,I660364);
nor I_38699 (I660590,I906825,I906813);
and I_38700 (I660607,I660455,I660590);
nor I_38701 (I660624,I660542,I660607);
DFFARX1 I_38702 (I660624,I2683,I660231,I660217,);
nor I_38703 (I660655,I660257,I660590);
DFFARX1 I_38704 (I660655,I2683,I660231,I660202,);
nor I_38705 (I660686,I660534,I660590);
not I_38706 (I660703,I660686);
nand I_38707 (I660211,I660703,I660559);
not I_38708 (I660758,I2690);
DFFARX1 I_38709 (I844398,I2683,I660758,I660784,);
not I_38710 (I660792,I660784);
nand I_38711 (I660809,I844380,I844380);
and I_38712 (I660826,I660809,I844386);
DFFARX1 I_38713 (I660826,I2683,I660758,I660852,);
DFFARX1 I_38714 (I660852,I2683,I660758,I660747,);
DFFARX1 I_38715 (I844383,I2683,I660758,I660883,);
nand I_38716 (I660891,I660883,I844392);
not I_38717 (I660908,I660891);
DFFARX1 I_38718 (I660908,I2683,I660758,I660934,);
not I_38719 (I660942,I660934);
nor I_38720 (I660750,I660792,I660942);
DFFARX1 I_38721 (I844404,I2683,I660758,I660982,);
nor I_38722 (I660741,I660982,I660852);
nor I_38723 (I660732,I660982,I660908);
nand I_38724 (I661018,I844395,I844389);
and I_38725 (I661035,I661018,I844383);
DFFARX1 I_38726 (I661035,I2683,I660758,I661061,);
not I_38727 (I661069,I661061);
nand I_38728 (I661086,I661069,I660982);
nand I_38729 (I660735,I661069,I660891);
nor I_38730 (I661117,I844401,I844389);
and I_38731 (I661134,I660982,I661117);
nor I_38732 (I661151,I661069,I661134);
DFFARX1 I_38733 (I661151,I2683,I660758,I660744,);
nor I_38734 (I661182,I660784,I661117);
DFFARX1 I_38735 (I661182,I2683,I660758,I660729,);
nor I_38736 (I661213,I661061,I661117);
not I_38737 (I661230,I661213);
nand I_38738 (I660738,I661230,I661086);
not I_38739 (I661285,I2690);
DFFARX1 I_38740 (I337752,I2683,I661285,I661311,);
not I_38741 (I661319,I661311);
nand I_38742 (I661336,I337749,I337758);
and I_38743 (I661353,I661336,I337767);
DFFARX1 I_38744 (I661353,I2683,I661285,I661379,);
DFFARX1 I_38745 (I661379,I2683,I661285,I661274,);
DFFARX1 I_38746 (I337770,I2683,I661285,I661410,);
nand I_38747 (I661418,I661410,I337773);
not I_38748 (I661435,I661418);
DFFARX1 I_38749 (I661435,I2683,I661285,I661461,);
not I_38750 (I661469,I661461);
nor I_38751 (I661277,I661319,I661469);
DFFARX1 I_38752 (I337746,I2683,I661285,I661509,);
nor I_38753 (I661268,I661509,I661379);
nor I_38754 (I661259,I661509,I661435);
nand I_38755 (I661545,I337761,I337764);
and I_38756 (I661562,I661545,I337755);
DFFARX1 I_38757 (I661562,I2683,I661285,I661588,);
not I_38758 (I661596,I661588);
nand I_38759 (I661613,I661596,I661509);
nand I_38760 (I661262,I661596,I661418);
nor I_38761 (I661644,I337746,I337764);
and I_38762 (I661661,I661509,I661644);
nor I_38763 (I661678,I661596,I661661);
DFFARX1 I_38764 (I661678,I2683,I661285,I661271,);
nor I_38765 (I661709,I661311,I661644);
DFFARX1 I_38766 (I661709,I2683,I661285,I661256,);
nor I_38767 (I661740,I661588,I661644);
not I_38768 (I661757,I661740);
nand I_38769 (I661265,I661757,I661613);
not I_38770 (I661812,I2690);
DFFARX1 I_38771 (I848444,I2683,I661812,I661838,);
not I_38772 (I661846,I661838);
nand I_38773 (I661863,I848426,I848426);
and I_38774 (I661880,I661863,I848432);
DFFARX1 I_38775 (I661880,I2683,I661812,I661906,);
DFFARX1 I_38776 (I661906,I2683,I661812,I661801,);
DFFARX1 I_38777 (I848429,I2683,I661812,I661937,);
nand I_38778 (I661945,I661937,I848438);
not I_38779 (I661962,I661945);
DFFARX1 I_38780 (I661962,I2683,I661812,I661988,);
not I_38781 (I661996,I661988);
nor I_38782 (I661804,I661846,I661996);
DFFARX1 I_38783 (I848450,I2683,I661812,I662036,);
nor I_38784 (I661795,I662036,I661906);
nor I_38785 (I661786,I662036,I661962);
nand I_38786 (I662072,I848441,I848435);
and I_38787 (I662089,I662072,I848429);
DFFARX1 I_38788 (I662089,I2683,I661812,I662115,);
not I_38789 (I662123,I662115);
nand I_38790 (I662140,I662123,I662036);
nand I_38791 (I661789,I662123,I661945);
nor I_38792 (I662171,I848447,I848435);
and I_38793 (I662188,I662036,I662171);
nor I_38794 (I662205,I662123,I662188);
DFFARX1 I_38795 (I662205,I2683,I661812,I661798,);
nor I_38796 (I662236,I661838,I662171);
DFFARX1 I_38797 (I662236,I2683,I661812,I661783,);
nor I_38798 (I662267,I662115,I662171);
not I_38799 (I662284,I662267);
nand I_38800 (I661792,I662284,I662140);
not I_38801 (I662339,I2690);
DFFARX1 I_38802 (I726454,I2683,I662339,I662365,);
not I_38803 (I662373,I662365);
nand I_38804 (I662390,I726469,I726451);
and I_38805 (I662407,I662390,I726451);
DFFARX1 I_38806 (I662407,I2683,I662339,I662433,);
DFFARX1 I_38807 (I662433,I2683,I662339,I662328,);
DFFARX1 I_38808 (I726460,I2683,I662339,I662464,);
nand I_38809 (I662472,I662464,I726478);
not I_38810 (I662489,I662472);
DFFARX1 I_38811 (I662489,I2683,I662339,I662515,);
not I_38812 (I662523,I662515);
nor I_38813 (I662331,I662373,I662523);
DFFARX1 I_38814 (I726475,I2683,I662339,I662563,);
nor I_38815 (I662322,I662563,I662433);
nor I_38816 (I662313,I662563,I662489);
nand I_38817 (I662599,I726472,I726463);
and I_38818 (I662616,I662599,I726457);
DFFARX1 I_38819 (I662616,I2683,I662339,I662642,);
not I_38820 (I662650,I662642);
nand I_38821 (I662667,I662650,I662563);
nand I_38822 (I662316,I662650,I662472);
nor I_38823 (I662698,I726466,I726463);
and I_38824 (I662715,I662563,I662698);
nor I_38825 (I662732,I662650,I662715);
DFFARX1 I_38826 (I662732,I2683,I662339,I662325,);
nor I_38827 (I662763,I662365,I662698);
DFFARX1 I_38828 (I662763,I2683,I662339,I662310,);
nor I_38829 (I662794,I662642,I662698);
not I_38830 (I662811,I662794);
nand I_38831 (I662319,I662811,I662667);
not I_38832 (I662866,I2690);
DFFARX1 I_38833 (I79625,I2683,I662866,I662892,);
not I_38834 (I662900,I662892);
nand I_38835 (I662917,I79601,I79610);
and I_38836 (I662934,I662917,I79604);
DFFARX1 I_38837 (I662934,I2683,I662866,I662960,);
DFFARX1 I_38838 (I662960,I2683,I662866,I662855,);
DFFARX1 I_38839 (I79622,I2683,I662866,I662991,);
nand I_38840 (I662999,I662991,I79613);
not I_38841 (I663016,I662999);
DFFARX1 I_38842 (I663016,I2683,I662866,I663042,);
not I_38843 (I663050,I663042);
nor I_38844 (I662858,I662900,I663050);
DFFARX1 I_38845 (I79607,I2683,I662866,I663090,);
nor I_38846 (I662849,I663090,I662960);
nor I_38847 (I662840,I663090,I663016);
nand I_38848 (I663126,I79619,I79616);
and I_38849 (I663143,I663126,I79604);
DFFARX1 I_38850 (I663143,I2683,I662866,I663169,);
not I_38851 (I663177,I663169);
nand I_38852 (I663194,I663177,I663090);
nand I_38853 (I662843,I663177,I662999);
nor I_38854 (I663225,I79601,I79616);
and I_38855 (I663242,I663090,I663225);
nor I_38856 (I663259,I663177,I663242);
DFFARX1 I_38857 (I663259,I2683,I662866,I662852,);
nor I_38858 (I663290,I662892,I663225);
DFFARX1 I_38859 (I663290,I2683,I662866,I662837,);
nor I_38860 (I663321,I663169,I663225);
not I_38861 (I663338,I663321);
nand I_38862 (I662846,I663338,I663194);
not I_38863 (I663393,I2690);
DFFARX1 I_38864 (I94381,I2683,I663393,I663419,);
not I_38865 (I663427,I663419);
nand I_38866 (I663444,I94357,I94366);
and I_38867 (I663461,I663444,I94360);
DFFARX1 I_38868 (I663461,I2683,I663393,I663487,);
DFFARX1 I_38869 (I663487,I2683,I663393,I663382,);
DFFARX1 I_38870 (I94378,I2683,I663393,I663518,);
nand I_38871 (I663526,I663518,I94369);
not I_38872 (I663543,I663526);
DFFARX1 I_38873 (I663543,I2683,I663393,I663569,);
not I_38874 (I663577,I663569);
nor I_38875 (I663385,I663427,I663577);
DFFARX1 I_38876 (I94363,I2683,I663393,I663617,);
nor I_38877 (I663376,I663617,I663487);
nor I_38878 (I663367,I663617,I663543);
nand I_38879 (I663653,I94375,I94372);
and I_38880 (I663670,I663653,I94360);
DFFARX1 I_38881 (I663670,I2683,I663393,I663696,);
not I_38882 (I663704,I663696);
nand I_38883 (I663721,I663704,I663617);
nand I_38884 (I663370,I663704,I663526);
nor I_38885 (I663752,I94357,I94372);
and I_38886 (I663769,I663617,I663752);
nor I_38887 (I663786,I663704,I663769);
DFFARX1 I_38888 (I663786,I2683,I663393,I663379,);
nor I_38889 (I663817,I663419,I663752);
DFFARX1 I_38890 (I663817,I2683,I663393,I663364,);
nor I_38891 (I663848,I663696,I663752);
not I_38892 (I663865,I663848);
nand I_38893 (I663373,I663865,I663721);
not I_38894 (I663920,I2690);
DFFARX1 I_38895 (I856536,I2683,I663920,I663946,);
not I_38896 (I663954,I663946);
nand I_38897 (I663971,I856518,I856518);
and I_38898 (I663988,I663971,I856524);
DFFARX1 I_38899 (I663988,I2683,I663920,I664014,);
DFFARX1 I_38900 (I664014,I2683,I663920,I663909,);
DFFARX1 I_38901 (I856521,I2683,I663920,I664045,);
nand I_38902 (I664053,I664045,I856530);
not I_38903 (I664070,I664053);
DFFARX1 I_38904 (I664070,I2683,I663920,I664096,);
not I_38905 (I664104,I664096);
nor I_38906 (I663912,I663954,I664104);
DFFARX1 I_38907 (I856542,I2683,I663920,I664144,);
nor I_38908 (I663903,I664144,I664014);
nor I_38909 (I663894,I664144,I664070);
nand I_38910 (I664180,I856533,I856527);
and I_38911 (I664197,I664180,I856521);
DFFARX1 I_38912 (I664197,I2683,I663920,I664223,);
not I_38913 (I664231,I664223);
nand I_38914 (I664248,I664231,I664144);
nand I_38915 (I663897,I664231,I664053);
nor I_38916 (I664279,I856539,I856527);
and I_38917 (I664296,I664144,I664279);
nor I_38918 (I664313,I664231,I664296);
DFFARX1 I_38919 (I664313,I2683,I663920,I663906,);
nor I_38920 (I664344,I663946,I664279);
DFFARX1 I_38921 (I664344,I2683,I663920,I663891,);
nor I_38922 (I664375,I664223,I664279);
not I_38923 (I664392,I664375);
nand I_38924 (I663900,I664392,I664248);
not I_38925 (I664447,I2690);
DFFARX1 I_38926 (I702552,I2683,I664447,I664473,);
not I_38927 (I664481,I664473);
nand I_38928 (I664498,I702567,I702549);
and I_38929 (I664515,I664498,I702549);
DFFARX1 I_38930 (I664515,I2683,I664447,I664541,);
DFFARX1 I_38931 (I664541,I2683,I664447,I664436,);
DFFARX1 I_38932 (I702558,I2683,I664447,I664572,);
nand I_38933 (I664580,I664572,I702576);
not I_38934 (I664597,I664580);
DFFARX1 I_38935 (I664597,I2683,I664447,I664623,);
not I_38936 (I664631,I664623);
nor I_38937 (I664439,I664481,I664631);
DFFARX1 I_38938 (I702573,I2683,I664447,I664671,);
nor I_38939 (I664430,I664671,I664541);
nor I_38940 (I664421,I664671,I664597);
nand I_38941 (I664707,I702570,I702561);
and I_38942 (I664724,I664707,I702555);
DFFARX1 I_38943 (I664724,I2683,I664447,I664750,);
not I_38944 (I664758,I664750);
nand I_38945 (I664775,I664758,I664671);
nand I_38946 (I664424,I664758,I664580);
nor I_38947 (I664806,I702564,I702561);
and I_38948 (I664823,I664671,I664806);
nor I_38949 (I664840,I664758,I664823);
DFFARX1 I_38950 (I664840,I2683,I664447,I664433,);
nor I_38951 (I664871,I664473,I664806);
DFFARX1 I_38952 (I664871,I2683,I664447,I664418,);
nor I_38953 (I664902,I664750,I664806);
not I_38954 (I664919,I664902);
nand I_38955 (I664427,I664919,I664775);
not I_38956 (I664974,I2690);
DFFARX1 I_38957 (I178326,I2683,I664974,I665000,);
not I_38958 (I665008,I665000);
nand I_38959 (I665025,I178323,I178341);
and I_38960 (I665042,I665025,I178332);
DFFARX1 I_38961 (I665042,I2683,I664974,I665068,);
DFFARX1 I_38962 (I665068,I2683,I664974,I664963,);
DFFARX1 I_38963 (I178338,I2683,I664974,I665099,);
nand I_38964 (I665107,I665099,I178335);
not I_38965 (I665124,I665107);
DFFARX1 I_38966 (I665124,I2683,I664974,I665150,);
not I_38967 (I665158,I665150);
nor I_38968 (I664966,I665008,I665158);
DFFARX1 I_38969 (I178329,I2683,I664974,I665198,);
nor I_38970 (I664957,I665198,I665068);
nor I_38971 (I664948,I665198,I665124);
nand I_38972 (I665234,I178320,I178344);
and I_38973 (I665251,I665234,I178323);
DFFARX1 I_38974 (I665251,I2683,I664974,I665277,);
not I_38975 (I665285,I665277);
nand I_38976 (I665302,I665285,I665198);
nand I_38977 (I664951,I665285,I665107);
nor I_38978 (I665333,I178320,I178344);
and I_38979 (I665350,I665198,I665333);
nor I_38980 (I665367,I665285,I665350);
DFFARX1 I_38981 (I665367,I2683,I664974,I664960,);
nor I_38982 (I665398,I665000,I665333);
DFFARX1 I_38983 (I665398,I2683,I664974,I664945,);
nor I_38984 (I665429,I665277,I665333);
not I_38985 (I665446,I665429);
nand I_38986 (I664954,I665446,I665302);
not I_38987 (I665501,I2690);
DFFARX1 I_38988 (I750356,I2683,I665501,I665527,);
not I_38989 (I665535,I665527);
nand I_38990 (I665552,I750371,I750353);
and I_38991 (I665569,I665552,I750353);
DFFARX1 I_38992 (I665569,I2683,I665501,I665595,);
DFFARX1 I_38993 (I665595,I2683,I665501,I665490,);
DFFARX1 I_38994 (I750362,I2683,I665501,I665626,);
nand I_38995 (I665634,I665626,I750380);
not I_38996 (I665651,I665634);
DFFARX1 I_38997 (I665651,I2683,I665501,I665677,);
not I_38998 (I665685,I665677);
nor I_38999 (I665493,I665535,I665685);
DFFARX1 I_39000 (I750377,I2683,I665501,I665725,);
nor I_39001 (I665484,I665725,I665595);
nor I_39002 (I665475,I665725,I665651);
nand I_39003 (I665761,I750374,I750365);
and I_39004 (I665778,I665761,I750359);
DFFARX1 I_39005 (I665778,I2683,I665501,I665804,);
not I_39006 (I665812,I665804);
nand I_39007 (I665829,I665812,I665725);
nand I_39008 (I665478,I665812,I665634);
nor I_39009 (I665860,I750368,I750365);
and I_39010 (I665877,I665725,I665860);
nor I_39011 (I665894,I665812,I665877);
DFFARX1 I_39012 (I665894,I2683,I665501,I665487,);
nor I_39013 (I665925,I665527,I665860);
DFFARX1 I_39014 (I665925,I2683,I665501,I665472,);
nor I_39015 (I665956,I665804,I665860);
not I_39016 (I665973,I665956);
nand I_39017 (I665481,I665973,I665829);
not I_39018 (I666028,I2690);
DFFARX1 I_39019 (I811375,I2683,I666028,I666054,);
not I_39020 (I666062,I666054);
nand I_39021 (I666079,I811384,I811372);
and I_39022 (I666096,I666079,I811369);
DFFARX1 I_39023 (I666096,I2683,I666028,I666122,);
DFFARX1 I_39024 (I666122,I2683,I666028,I666017,);
DFFARX1 I_39025 (I811369,I2683,I666028,I666153,);
nand I_39026 (I666161,I666153,I811366);
not I_39027 (I666178,I666161);
DFFARX1 I_39028 (I666178,I2683,I666028,I666204,);
not I_39029 (I666212,I666204);
nor I_39030 (I666020,I666062,I666212);
DFFARX1 I_39031 (I811372,I2683,I666028,I666252,);
nor I_39032 (I666011,I666252,I666122);
nor I_39033 (I666002,I666252,I666178);
nand I_39034 (I666288,I811387,I811378);
and I_39035 (I666305,I666288,I811381);
DFFARX1 I_39036 (I666305,I2683,I666028,I666331,);
not I_39037 (I666339,I666331);
nand I_39038 (I666356,I666339,I666252);
nand I_39039 (I666005,I666339,I666161);
nor I_39040 (I666387,I811366,I811378);
and I_39041 (I666404,I666252,I666387);
nor I_39042 (I666421,I666339,I666404);
DFFARX1 I_39043 (I666421,I2683,I666028,I666014,);
nor I_39044 (I666452,I666054,I666387);
DFFARX1 I_39045 (I666452,I2683,I666028,I665999,);
nor I_39046 (I666483,I666331,I666387);
not I_39047 (I666500,I666483);
nand I_39048 (I666008,I666500,I666356);
not I_39049 (I666555,I2690);
DFFARX1 I_39050 (I459005,I2683,I666555,I666581,);
not I_39051 (I666589,I666581);
nand I_39052 (I666606,I458990,I459011);
and I_39053 (I666623,I666606,I458999);
DFFARX1 I_39054 (I666623,I2683,I666555,I666649,);
DFFARX1 I_39055 (I666649,I2683,I666555,I666544,);
DFFARX1 I_39056 (I458993,I2683,I666555,I666680,);
nand I_39057 (I666688,I666680,I459002);
not I_39058 (I666705,I666688);
DFFARX1 I_39059 (I666705,I2683,I666555,I666731,);
not I_39060 (I666739,I666731);
nor I_39061 (I666547,I666589,I666739);
DFFARX1 I_39062 (I459008,I2683,I666555,I666779,);
nor I_39063 (I666538,I666779,I666649);
nor I_39064 (I666529,I666779,I666705);
nand I_39065 (I666815,I458990,I458993);
and I_39066 (I666832,I666815,I459014);
DFFARX1 I_39067 (I666832,I2683,I666555,I666858,);
not I_39068 (I666866,I666858);
nand I_39069 (I666883,I666866,I666779);
nand I_39070 (I666532,I666866,I666688);
nor I_39071 (I666914,I458996,I458993);
and I_39072 (I666931,I666779,I666914);
nor I_39073 (I666948,I666866,I666931);
DFFARX1 I_39074 (I666948,I2683,I666555,I666541,);
nor I_39075 (I666979,I666581,I666914);
DFFARX1 I_39076 (I666979,I2683,I666555,I666526,);
nor I_39077 (I667010,I666858,I666914);
not I_39078 (I667027,I667010);
nand I_39079 (I666535,I667027,I666883);
not I_39080 (I667082,I2690);
DFFARX1 I_39081 (I246431,I2683,I667082,I667108,);
not I_39082 (I667116,I667108);
nand I_39083 (I667133,I246422,I246422);
and I_39084 (I667150,I667133,I246440);
DFFARX1 I_39085 (I667150,I2683,I667082,I667176,);
DFFARX1 I_39086 (I667176,I2683,I667082,I667071,);
DFFARX1 I_39087 (I246443,I2683,I667082,I667207,);
nand I_39088 (I667215,I667207,I246425);
not I_39089 (I667232,I667215);
DFFARX1 I_39090 (I667232,I2683,I667082,I667258,);
not I_39091 (I667266,I667258);
nor I_39092 (I667074,I667116,I667266);
DFFARX1 I_39093 (I246437,I2683,I667082,I667306,);
nor I_39094 (I667065,I667306,I667176);
nor I_39095 (I667056,I667306,I667232);
nand I_39096 (I667342,I246449,I246428);
and I_39097 (I667359,I667342,I246434);
DFFARX1 I_39098 (I667359,I2683,I667082,I667385,);
not I_39099 (I667393,I667385);
nand I_39100 (I667410,I667393,I667306);
nand I_39101 (I667059,I667393,I667215);
nor I_39102 (I667441,I246446,I246428);
and I_39103 (I667458,I667306,I667441);
nor I_39104 (I667475,I667393,I667458);
DFFARX1 I_39105 (I667475,I2683,I667082,I667068,);
nor I_39106 (I667506,I667108,I667441);
DFFARX1 I_39107 (I667506,I2683,I667082,I667053,);
nor I_39108 (I667537,I667385,I667441);
not I_39109 (I667554,I667537);
nand I_39110 (I667062,I667554,I667410);
not I_39111 (I667609,I2690);
DFFARX1 I_39112 (I1055484,I2683,I667609,I667635,);
not I_39113 (I667643,I667635);
nand I_39114 (I667660,I1055481,I1055490);
and I_39115 (I667677,I667660,I1055469);
DFFARX1 I_39116 (I667677,I2683,I667609,I667703,);
DFFARX1 I_39117 (I667703,I2683,I667609,I667598,);
DFFARX1 I_39118 (I1055472,I2683,I667609,I667734,);
nand I_39119 (I667742,I667734,I1055487);
not I_39120 (I667759,I667742);
DFFARX1 I_39121 (I667759,I2683,I667609,I667785,);
not I_39122 (I667793,I667785);
nor I_39123 (I667601,I667643,I667793);
DFFARX1 I_39124 (I1055493,I2683,I667609,I667833,);
nor I_39125 (I667592,I667833,I667703);
nor I_39126 (I667583,I667833,I667759);
nand I_39127 (I667869,I1055475,I1055496);
and I_39128 (I667886,I667869,I1055478);
DFFARX1 I_39129 (I667886,I2683,I667609,I667912,);
not I_39130 (I667920,I667912);
nand I_39131 (I667937,I667920,I667833);
nand I_39132 (I667586,I667920,I667742);
nor I_39133 (I667968,I1055469,I1055496);
and I_39134 (I667985,I667833,I667968);
nor I_39135 (I668002,I667920,I667985);
DFFARX1 I_39136 (I668002,I2683,I667609,I667595,);
nor I_39137 (I668033,I667635,I667968);
DFFARX1 I_39138 (I668033,I2683,I667609,I667580,);
nor I_39139 (I668064,I667912,I667968);
not I_39140 (I668081,I668064);
nand I_39141 (I667589,I668081,I667937);
not I_39142 (I668136,I2690);
DFFARX1 I_39143 (I1074524,I2683,I668136,I668162,);
not I_39144 (I668170,I668162);
nand I_39145 (I668187,I1074521,I1074530);
and I_39146 (I668204,I668187,I1074509);
DFFARX1 I_39147 (I668204,I2683,I668136,I668230,);
DFFARX1 I_39148 (I668230,I2683,I668136,I668125,);
DFFARX1 I_39149 (I1074512,I2683,I668136,I668261,);
nand I_39150 (I668269,I668261,I1074527);
not I_39151 (I668286,I668269);
DFFARX1 I_39152 (I668286,I2683,I668136,I668312,);
not I_39153 (I668320,I668312);
nor I_39154 (I668128,I668170,I668320);
DFFARX1 I_39155 (I1074533,I2683,I668136,I668360,);
nor I_39156 (I668119,I668360,I668230);
nor I_39157 (I668110,I668360,I668286);
nand I_39158 (I668396,I1074515,I1074536);
and I_39159 (I668413,I668396,I1074518);
DFFARX1 I_39160 (I668413,I2683,I668136,I668439,);
not I_39161 (I668447,I668439);
nand I_39162 (I668464,I668447,I668360);
nand I_39163 (I668113,I668447,I668269);
nor I_39164 (I668495,I1074509,I1074536);
and I_39165 (I668512,I668360,I668495);
nor I_39166 (I668529,I668447,I668512);
DFFARX1 I_39167 (I668529,I2683,I668136,I668122,);
nor I_39168 (I668560,I668162,I668495);
DFFARX1 I_39169 (I668560,I2683,I668136,I668107,);
nor I_39170 (I668591,I668439,I668495);
not I_39171 (I668608,I668591);
nand I_39172 (I668116,I668608,I668464);
not I_39173 (I668663,I2690);
DFFARX1 I_39174 (I498294,I2683,I668663,I668689,);
not I_39175 (I668697,I668689);
nand I_39176 (I668714,I498297,I498294);
and I_39177 (I668731,I668714,I498306);
DFFARX1 I_39178 (I668731,I2683,I668663,I668757,);
DFFARX1 I_39179 (I668757,I2683,I668663,I668652,);
DFFARX1 I_39180 (I498303,I2683,I668663,I668788,);
nand I_39181 (I668796,I668788,I498309);
not I_39182 (I668813,I668796);
DFFARX1 I_39183 (I668813,I2683,I668663,I668839,);
not I_39184 (I668847,I668839);
nor I_39185 (I668655,I668697,I668847);
DFFARX1 I_39186 (I498318,I2683,I668663,I668887,);
nor I_39187 (I668646,I668887,I668757);
nor I_39188 (I668637,I668887,I668813);
nand I_39189 (I668923,I498312,I498300);
and I_39190 (I668940,I668923,I498297);
DFFARX1 I_39191 (I668940,I2683,I668663,I668966,);
not I_39192 (I668974,I668966);
nand I_39193 (I668991,I668974,I668887);
nand I_39194 (I668640,I668974,I668796);
nor I_39195 (I669022,I498315,I498300);
and I_39196 (I669039,I668887,I669022);
nor I_39197 (I669056,I668974,I669039);
DFFARX1 I_39198 (I669056,I2683,I668663,I668649,);
nor I_39199 (I669087,I668689,I669022);
DFFARX1 I_39200 (I669087,I2683,I668663,I668634,);
nor I_39201 (I669118,I668966,I669022);
not I_39202 (I669135,I669118);
nand I_39203 (I668643,I669135,I668991);
not I_39204 (I669190,I2690);
DFFARX1 I_39205 (I100178,I2683,I669190,I669216,);
not I_39206 (I669224,I669216);
nand I_39207 (I669241,I100154,I100163);
and I_39208 (I669258,I669241,I100157);
DFFARX1 I_39209 (I669258,I2683,I669190,I669284,);
DFFARX1 I_39210 (I669284,I2683,I669190,I669179,);
DFFARX1 I_39211 (I100175,I2683,I669190,I669315,);
nand I_39212 (I669323,I669315,I100166);
not I_39213 (I669340,I669323);
DFFARX1 I_39214 (I669340,I2683,I669190,I669366,);
not I_39215 (I669374,I669366);
nor I_39216 (I669182,I669224,I669374);
DFFARX1 I_39217 (I100160,I2683,I669190,I669414,);
nor I_39218 (I669173,I669414,I669284);
nor I_39219 (I669164,I669414,I669340);
nand I_39220 (I669450,I100172,I100169);
and I_39221 (I669467,I669450,I100157);
DFFARX1 I_39222 (I669467,I2683,I669190,I669493,);
not I_39223 (I669501,I669493);
nand I_39224 (I669518,I669501,I669414);
nand I_39225 (I669167,I669501,I669323);
nor I_39226 (I669549,I100154,I100169);
and I_39227 (I669566,I669414,I669549);
nor I_39228 (I669583,I669501,I669566);
DFFARX1 I_39229 (I669583,I2683,I669190,I669176,);
nor I_39230 (I669614,I669216,I669549);
DFFARX1 I_39231 (I669614,I2683,I669190,I669161,);
nor I_39232 (I669645,I669493,I669549);
not I_39233 (I669662,I669645);
nand I_39234 (I669170,I669662,I669518);
not I_39235 (I669717,I2690);
DFFARX1 I_39236 (I1073929,I2683,I669717,I669743,);
not I_39237 (I669751,I669743);
nand I_39238 (I669768,I1073926,I1073935);
and I_39239 (I669785,I669768,I1073914);
DFFARX1 I_39240 (I669785,I2683,I669717,I669811,);
DFFARX1 I_39241 (I669811,I2683,I669717,I669706,);
DFFARX1 I_39242 (I1073917,I2683,I669717,I669842,);
nand I_39243 (I669850,I669842,I1073932);
not I_39244 (I669867,I669850);
DFFARX1 I_39245 (I669867,I2683,I669717,I669893,);
not I_39246 (I669901,I669893);
nor I_39247 (I669709,I669751,I669901);
DFFARX1 I_39248 (I1073938,I2683,I669717,I669941,);
nor I_39249 (I669700,I669941,I669811);
nor I_39250 (I669691,I669941,I669867);
nand I_39251 (I669977,I1073920,I1073941);
and I_39252 (I669994,I669977,I1073923);
DFFARX1 I_39253 (I669994,I2683,I669717,I670020,);
not I_39254 (I670028,I670020);
nand I_39255 (I670045,I670028,I669941);
nand I_39256 (I669694,I670028,I669850);
nor I_39257 (I670076,I1073914,I1073941);
and I_39258 (I670093,I669941,I670076);
nor I_39259 (I670110,I670028,I670093);
DFFARX1 I_39260 (I670110,I2683,I669717,I669703,);
nor I_39261 (I670141,I669743,I670076);
DFFARX1 I_39262 (I670141,I2683,I669717,I669688,);
nor I_39263 (I670172,I670020,I670076);
not I_39264 (I670189,I670172);
nand I_39265 (I669697,I670189,I670045);
not I_39266 (I670244,I2690);
DFFARX1 I_39267 (I796228,I2683,I670244,I670270,);
not I_39268 (I670278,I670270);
nand I_39269 (I670295,I796237,I796225);
and I_39270 (I670312,I670295,I796222);
DFFARX1 I_39271 (I670312,I2683,I670244,I670338,);
DFFARX1 I_39272 (I670338,I2683,I670244,I670233,);
DFFARX1 I_39273 (I796222,I2683,I670244,I670369,);
nand I_39274 (I670377,I670369,I796219);
not I_39275 (I670394,I670377);
DFFARX1 I_39276 (I670394,I2683,I670244,I670420,);
not I_39277 (I670428,I670420);
nor I_39278 (I670236,I670278,I670428);
DFFARX1 I_39279 (I796225,I2683,I670244,I670468,);
nor I_39280 (I670227,I670468,I670338);
nor I_39281 (I670218,I670468,I670394);
nand I_39282 (I670504,I796240,I796231);
and I_39283 (I670521,I670504,I796234);
DFFARX1 I_39284 (I670521,I2683,I670244,I670547,);
not I_39285 (I670555,I670547);
nand I_39286 (I670572,I670555,I670468);
nand I_39287 (I670221,I670555,I670377);
nor I_39288 (I670603,I796219,I796231);
and I_39289 (I670620,I670468,I670603);
nor I_39290 (I670637,I670555,I670620);
DFFARX1 I_39291 (I670637,I2683,I670244,I670230,);
nor I_39292 (I670668,I670270,I670603);
DFFARX1 I_39293 (I670668,I2683,I670244,I670215,);
nor I_39294 (I670699,I670547,I670603);
not I_39295 (I670716,I670699);
nand I_39296 (I670224,I670716,I670572);
not I_39297 (I670771,I2690);
DFFARX1 I_39298 (I849600,I2683,I670771,I670797,);
not I_39299 (I670805,I670797);
nand I_39300 (I670822,I849582,I849582);
and I_39301 (I670839,I670822,I849588);
DFFARX1 I_39302 (I670839,I2683,I670771,I670865,);
DFFARX1 I_39303 (I670865,I2683,I670771,I670760,);
DFFARX1 I_39304 (I849585,I2683,I670771,I670896,);
nand I_39305 (I670904,I670896,I849594);
not I_39306 (I670921,I670904);
DFFARX1 I_39307 (I670921,I2683,I670771,I670947,);
not I_39308 (I670955,I670947);
nor I_39309 (I670763,I670805,I670955);
DFFARX1 I_39310 (I849606,I2683,I670771,I670995,);
nor I_39311 (I670754,I670995,I670865);
nor I_39312 (I670745,I670995,I670921);
nand I_39313 (I671031,I849597,I849591);
and I_39314 (I671048,I671031,I849585);
DFFARX1 I_39315 (I671048,I2683,I670771,I671074,);
not I_39316 (I671082,I671074);
nand I_39317 (I671099,I671082,I670995);
nand I_39318 (I670748,I671082,I670904);
nor I_39319 (I671130,I849603,I849591);
and I_39320 (I671147,I670995,I671130);
nor I_39321 (I671164,I671082,I671147);
DFFARX1 I_39322 (I671164,I2683,I670771,I670757,);
nor I_39323 (I671195,I670797,I671130);
DFFARX1 I_39324 (I671195,I2683,I670771,I670742,);
nor I_39325 (I671226,I671074,I671130);
not I_39326 (I671243,I671226);
nand I_39327 (I670751,I671243,I671099);
not I_39328 (I671298,I2690);
DFFARX1 I_39329 (I280159,I2683,I671298,I671324,);
not I_39330 (I671332,I671324);
nand I_39331 (I671349,I280150,I280150);
and I_39332 (I671366,I671349,I280168);
DFFARX1 I_39333 (I671366,I2683,I671298,I671392,);
DFFARX1 I_39334 (I671392,I2683,I671298,I671287,);
DFFARX1 I_39335 (I280171,I2683,I671298,I671423,);
nand I_39336 (I671431,I671423,I280153);
not I_39337 (I671448,I671431);
DFFARX1 I_39338 (I671448,I2683,I671298,I671474,);
not I_39339 (I671482,I671474);
nor I_39340 (I671290,I671332,I671482);
DFFARX1 I_39341 (I280165,I2683,I671298,I671522,);
nor I_39342 (I671281,I671522,I671392);
nor I_39343 (I671272,I671522,I671448);
nand I_39344 (I671558,I280177,I280156);
and I_39345 (I671575,I671558,I280162);
DFFARX1 I_39346 (I671575,I2683,I671298,I671601,);
not I_39347 (I671609,I671601);
nand I_39348 (I671626,I671609,I671522);
nand I_39349 (I671275,I671609,I671431);
nor I_39350 (I671657,I280174,I280156);
and I_39351 (I671674,I671522,I671657);
nor I_39352 (I671691,I671609,I671674);
DFFARX1 I_39353 (I671691,I2683,I671298,I671284,);
nor I_39354 (I671722,I671324,I671657);
DFFARX1 I_39355 (I671722,I2683,I671298,I671269,);
nor I_39356 (I671753,I671601,I671657);
not I_39357 (I671770,I671753);
nand I_39358 (I671278,I671770,I671626);
not I_39359 (I671825,I2690);
DFFARX1 I_39360 (I864050,I2683,I671825,I671851,);
not I_39361 (I671859,I671851);
nand I_39362 (I671876,I864032,I864032);
and I_39363 (I671893,I671876,I864038);
DFFARX1 I_39364 (I671893,I2683,I671825,I671919,);
DFFARX1 I_39365 (I671919,I2683,I671825,I671814,);
DFFARX1 I_39366 (I864035,I2683,I671825,I671950,);
nand I_39367 (I671958,I671950,I864044);
not I_39368 (I671975,I671958);
DFFARX1 I_39369 (I671975,I2683,I671825,I672001,);
not I_39370 (I672009,I672001);
nor I_39371 (I671817,I671859,I672009);
DFFARX1 I_39372 (I864056,I2683,I671825,I672049,);
nor I_39373 (I671808,I672049,I671919);
nor I_39374 (I671799,I672049,I671975);
nand I_39375 (I672085,I864047,I864041);
and I_39376 (I672102,I672085,I864035);
DFFARX1 I_39377 (I672102,I2683,I671825,I672128,);
not I_39378 (I672136,I672128);
nand I_39379 (I672153,I672136,I672049);
nand I_39380 (I671802,I672136,I671958);
nor I_39381 (I672184,I864053,I864041);
and I_39382 (I672201,I672049,I672184);
nor I_39383 (I672218,I672136,I672201);
DFFARX1 I_39384 (I672218,I2683,I671825,I671811,);
nor I_39385 (I672249,I671851,I672184);
DFFARX1 I_39386 (I672249,I2683,I671825,I671796,);
nor I_39387 (I672280,I672128,I672184);
not I_39388 (I672297,I672280);
nand I_39389 (I671805,I672297,I672153);
not I_39390 (I672352,I2690);
DFFARX1 I_39391 (I862316,I2683,I672352,I672378,);
not I_39392 (I672386,I672378);
nand I_39393 (I672403,I862298,I862298);
and I_39394 (I672420,I672403,I862304);
DFFARX1 I_39395 (I672420,I2683,I672352,I672446,);
DFFARX1 I_39396 (I672446,I2683,I672352,I672341,);
DFFARX1 I_39397 (I862301,I2683,I672352,I672477,);
nand I_39398 (I672485,I672477,I862310);
not I_39399 (I672502,I672485);
DFFARX1 I_39400 (I672502,I2683,I672352,I672528,);
not I_39401 (I672536,I672528);
nor I_39402 (I672344,I672386,I672536);
DFFARX1 I_39403 (I862322,I2683,I672352,I672576,);
nor I_39404 (I672335,I672576,I672446);
nor I_39405 (I672326,I672576,I672502);
nand I_39406 (I672612,I862313,I862307);
and I_39407 (I672629,I672612,I862301);
DFFARX1 I_39408 (I672629,I2683,I672352,I672655,);
not I_39409 (I672663,I672655);
nand I_39410 (I672680,I672663,I672576);
nand I_39411 (I672329,I672663,I672485);
nor I_39412 (I672711,I862319,I862307);
and I_39413 (I672728,I672576,I672711);
nor I_39414 (I672745,I672663,I672728);
DFFARX1 I_39415 (I672745,I2683,I672352,I672338,);
nor I_39416 (I672776,I672378,I672711);
DFFARX1 I_39417 (I672776,I2683,I672352,I672323,);
nor I_39418 (I672807,I672655,I672711);
not I_39419 (I672824,I672807);
nand I_39420 (I672332,I672824,I672680);
not I_39421 (I672879,I2690);
DFFARX1 I_39422 (I829370,I2683,I672879,I672905,);
not I_39423 (I672913,I672905);
nand I_39424 (I672930,I829352,I829352);
and I_39425 (I672947,I672930,I829358);
DFFARX1 I_39426 (I672947,I2683,I672879,I672973,);
DFFARX1 I_39427 (I672973,I2683,I672879,I672868,);
DFFARX1 I_39428 (I829355,I2683,I672879,I673004,);
nand I_39429 (I673012,I673004,I829364);
not I_39430 (I673029,I673012);
DFFARX1 I_39431 (I673029,I2683,I672879,I673055,);
not I_39432 (I673063,I673055);
nor I_39433 (I672871,I672913,I673063);
DFFARX1 I_39434 (I829376,I2683,I672879,I673103,);
nor I_39435 (I672862,I673103,I672973);
nor I_39436 (I672853,I673103,I673029);
nand I_39437 (I673139,I829367,I829361);
and I_39438 (I673156,I673139,I829355);
DFFARX1 I_39439 (I673156,I2683,I672879,I673182,);
not I_39440 (I673190,I673182);
nand I_39441 (I673207,I673190,I673103);
nand I_39442 (I672856,I673190,I673012);
nor I_39443 (I673238,I829373,I829361);
and I_39444 (I673255,I673103,I673238);
nor I_39445 (I673272,I673190,I673255);
DFFARX1 I_39446 (I673272,I2683,I672879,I672865,);
nor I_39447 (I673303,I672905,I673238);
DFFARX1 I_39448 (I673303,I2683,I672879,I672850,);
nor I_39449 (I673334,I673182,I673238);
not I_39450 (I673351,I673334);
nand I_39451 (I672859,I673351,I673207);
not I_39452 (I673406,I2690);
DFFARX1 I_39453 (I1097729,I2683,I673406,I673432,);
not I_39454 (I673440,I673432);
nand I_39455 (I673457,I1097726,I1097735);
and I_39456 (I673474,I673457,I1097714);
DFFARX1 I_39457 (I673474,I2683,I673406,I673500,);
DFFARX1 I_39458 (I673500,I2683,I673406,I673395,);
DFFARX1 I_39459 (I1097717,I2683,I673406,I673531,);
nand I_39460 (I673539,I673531,I1097732);
not I_39461 (I673556,I673539);
DFFARX1 I_39462 (I673556,I2683,I673406,I673582,);
not I_39463 (I673590,I673582);
nor I_39464 (I673398,I673440,I673590);
DFFARX1 I_39465 (I1097738,I2683,I673406,I673630,);
nor I_39466 (I673389,I673630,I673500);
nor I_39467 (I673380,I673630,I673556);
nand I_39468 (I673666,I1097720,I1097741);
and I_39469 (I673683,I673666,I1097723);
DFFARX1 I_39470 (I673683,I2683,I673406,I673709,);
not I_39471 (I673717,I673709);
nand I_39472 (I673734,I673717,I673630);
nand I_39473 (I673383,I673717,I673539);
nor I_39474 (I673765,I1097714,I1097741);
and I_39475 (I673782,I673630,I673765);
nor I_39476 (I673799,I673717,I673782);
DFFARX1 I_39477 (I673799,I2683,I673406,I673392,);
nor I_39478 (I673830,I673432,I673765);
DFFARX1 I_39479 (I673830,I2683,I673406,I673377,);
nor I_39480 (I673861,I673709,I673765);
not I_39481 (I673878,I673861);
nand I_39482 (I673386,I673878,I673734);
not I_39483 (I673933,I2690);
DFFARX1 I_39484 (I715472,I2683,I673933,I673959,);
not I_39485 (I673967,I673959);
nand I_39486 (I673984,I715487,I715469);
and I_39487 (I674001,I673984,I715469);
DFFARX1 I_39488 (I674001,I2683,I673933,I674027,);
DFFARX1 I_39489 (I674027,I2683,I673933,I673922,);
DFFARX1 I_39490 (I715478,I2683,I673933,I674058,);
nand I_39491 (I674066,I674058,I715496);
not I_39492 (I674083,I674066);
DFFARX1 I_39493 (I674083,I2683,I673933,I674109,);
not I_39494 (I674117,I674109);
nor I_39495 (I673925,I673967,I674117);
DFFARX1 I_39496 (I715493,I2683,I673933,I674157,);
nor I_39497 (I673916,I674157,I674027);
nor I_39498 (I673907,I674157,I674083);
nand I_39499 (I674193,I715490,I715481);
and I_39500 (I674210,I674193,I715475);
DFFARX1 I_39501 (I674210,I2683,I673933,I674236,);
not I_39502 (I674244,I674236);
nand I_39503 (I674261,I674244,I674157);
nand I_39504 (I673910,I674244,I674066);
nor I_39505 (I674292,I715484,I715481);
and I_39506 (I674309,I674157,I674292);
nor I_39507 (I674326,I674244,I674309);
DFFARX1 I_39508 (I674326,I2683,I673933,I673919,);
nor I_39509 (I674357,I673959,I674292);
DFFARX1 I_39510 (I674357,I2683,I673933,I673904,);
nor I_39511 (I674388,I674236,I674292);
not I_39512 (I674405,I674388);
nand I_39513 (I673913,I674405,I674261);
not I_39514 (I674460,I2690);
DFFARX1 I_39515 (I868096,I2683,I674460,I674486,);
not I_39516 (I674494,I674486);
nand I_39517 (I674511,I868078,I868078);
and I_39518 (I674528,I674511,I868084);
DFFARX1 I_39519 (I674528,I2683,I674460,I674554,);
DFFARX1 I_39520 (I674554,I2683,I674460,I674449,);
DFFARX1 I_39521 (I868081,I2683,I674460,I674585,);
nand I_39522 (I674593,I674585,I868090);
not I_39523 (I674610,I674593);
DFFARX1 I_39524 (I674610,I2683,I674460,I674636,);
not I_39525 (I674644,I674636);
nor I_39526 (I674452,I674494,I674644);
DFFARX1 I_39527 (I868102,I2683,I674460,I674684,);
nor I_39528 (I674443,I674684,I674554);
nor I_39529 (I674434,I674684,I674610);
nand I_39530 (I674720,I868093,I868087);
and I_39531 (I674737,I674720,I868081);
DFFARX1 I_39532 (I674737,I2683,I674460,I674763,);
not I_39533 (I674771,I674763);
nand I_39534 (I674788,I674771,I674684);
nand I_39535 (I674437,I674771,I674593);
nor I_39536 (I674819,I868099,I868087);
and I_39537 (I674836,I674684,I674819);
nor I_39538 (I674853,I674771,I674836);
DFFARX1 I_39539 (I674853,I2683,I674460,I674446,);
nor I_39540 (I674884,I674486,I674819);
DFFARX1 I_39541 (I674884,I2683,I674460,I674431,);
nor I_39542 (I674915,I674763,I674819);
not I_39543 (I674932,I674915);
nand I_39544 (I674440,I674932,I674788);
not I_39545 (I674987,I2690);
DFFARX1 I_39546 (I397303,I2683,I674987,I675013,);
not I_39547 (I675021,I675013);
nand I_39548 (I675038,I397321,I397312);
and I_39549 (I675055,I675038,I397315);
DFFARX1 I_39550 (I675055,I2683,I674987,I675081,);
DFFARX1 I_39551 (I675081,I2683,I674987,I674976,);
DFFARX1 I_39552 (I397309,I2683,I674987,I675112,);
nand I_39553 (I675120,I675112,I397300);
not I_39554 (I675137,I675120);
DFFARX1 I_39555 (I675137,I2683,I674987,I675163,);
not I_39556 (I675171,I675163);
nor I_39557 (I674979,I675021,I675171);
DFFARX1 I_39558 (I397306,I2683,I674987,I675211,);
nor I_39559 (I674970,I675211,I675081);
nor I_39560 (I674961,I675211,I675137);
nand I_39561 (I675247,I397300,I397297);
and I_39562 (I675264,I675247,I397318);
DFFARX1 I_39563 (I675264,I2683,I674987,I675290,);
not I_39564 (I675298,I675290);
nand I_39565 (I675315,I675298,I675211);
nand I_39566 (I674964,I675298,I675120);
nor I_39567 (I675346,I397297,I397297);
and I_39568 (I675363,I675211,I675346);
nor I_39569 (I675380,I675298,I675363);
DFFARX1 I_39570 (I675380,I2683,I674987,I674973,);
nor I_39571 (I675411,I675013,I675346);
DFFARX1 I_39572 (I675411,I2683,I674987,I674958,);
nor I_39573 (I675442,I675290,I675346);
not I_39574 (I675459,I675442);
nand I_39575 (I674967,I675459,I675315);
not I_39576 (I675514,I2690);
DFFARX1 I_39577 (I888904,I2683,I675514,I675540,);
not I_39578 (I675548,I675540);
nand I_39579 (I675565,I888886,I888886);
and I_39580 (I675582,I675565,I888892);
DFFARX1 I_39581 (I675582,I2683,I675514,I675608,);
DFFARX1 I_39582 (I675608,I2683,I675514,I675503,);
DFFARX1 I_39583 (I888889,I2683,I675514,I675639,);
nand I_39584 (I675647,I675639,I888898);
not I_39585 (I675664,I675647);
DFFARX1 I_39586 (I675664,I2683,I675514,I675690,);
not I_39587 (I675698,I675690);
nor I_39588 (I675506,I675548,I675698);
DFFARX1 I_39589 (I888910,I2683,I675514,I675738,);
nor I_39590 (I675497,I675738,I675608);
nor I_39591 (I675488,I675738,I675664);
nand I_39592 (I675774,I888901,I888895);
and I_39593 (I675791,I675774,I888889);
DFFARX1 I_39594 (I675791,I2683,I675514,I675817,);
not I_39595 (I675825,I675817);
nand I_39596 (I675842,I675825,I675738);
nand I_39597 (I675491,I675825,I675647);
nor I_39598 (I675873,I888907,I888895);
and I_39599 (I675890,I675738,I675873);
nor I_39600 (I675907,I675825,I675890);
DFFARX1 I_39601 (I675907,I2683,I675514,I675500,);
nor I_39602 (I675938,I675540,I675873);
DFFARX1 I_39603 (I675938,I2683,I675514,I675485,);
nor I_39604 (I675969,I675817,I675873);
not I_39605 (I675986,I675969);
nand I_39606 (I675494,I675986,I675842);
not I_39607 (I676041,I2690);
DFFARX1 I_39608 (I898152,I2683,I676041,I676067,);
not I_39609 (I676075,I676067);
nand I_39610 (I676092,I898134,I898134);
and I_39611 (I676109,I676092,I898140);
DFFARX1 I_39612 (I676109,I2683,I676041,I676135,);
DFFARX1 I_39613 (I676135,I2683,I676041,I676030,);
DFFARX1 I_39614 (I898137,I2683,I676041,I676166,);
nand I_39615 (I676174,I676166,I898146);
not I_39616 (I676191,I676174);
DFFARX1 I_39617 (I676191,I2683,I676041,I676217,);
not I_39618 (I676225,I676217);
nor I_39619 (I676033,I676075,I676225);
DFFARX1 I_39620 (I898158,I2683,I676041,I676265,);
nor I_39621 (I676024,I676265,I676135);
nor I_39622 (I676015,I676265,I676191);
nand I_39623 (I676301,I898149,I898143);
and I_39624 (I676318,I676301,I898137);
DFFARX1 I_39625 (I676318,I2683,I676041,I676344,);
not I_39626 (I676352,I676344);
nand I_39627 (I676369,I676352,I676265);
nand I_39628 (I676018,I676352,I676174);
nor I_39629 (I676400,I898155,I898143);
and I_39630 (I676417,I676265,I676400);
nor I_39631 (I676434,I676352,I676417);
DFFARX1 I_39632 (I676434,I2683,I676041,I676027,);
nor I_39633 (I676465,I676067,I676400);
DFFARX1 I_39634 (I676465,I2683,I676041,I676012,);
nor I_39635 (I676496,I676344,I676400);
not I_39636 (I676513,I676496);
nand I_39637 (I676021,I676513,I676369);
not I_39638 (I676568,I2690);
DFFARX1 I_39639 (I26383,I2683,I676568,I676594,);
not I_39640 (I676602,I676594);
nand I_39641 (I676619,I26395,I26398);
and I_39642 (I676636,I676619,I26374);
DFFARX1 I_39643 (I676636,I2683,I676568,I676662,);
DFFARX1 I_39644 (I676662,I2683,I676568,I676557,);
DFFARX1 I_39645 (I26392,I2683,I676568,I676693,);
nand I_39646 (I676701,I676693,I26380);
not I_39647 (I676718,I676701);
DFFARX1 I_39648 (I676718,I2683,I676568,I676744,);
not I_39649 (I676752,I676744);
nor I_39650 (I676560,I676602,I676752);
DFFARX1 I_39651 (I26377,I2683,I676568,I676792,);
nor I_39652 (I676551,I676792,I676662);
nor I_39653 (I676542,I676792,I676718);
nand I_39654 (I676828,I26386,I26377);
and I_39655 (I676845,I676828,I26374);
DFFARX1 I_39656 (I676845,I2683,I676568,I676871,);
not I_39657 (I676879,I676871);
nand I_39658 (I676896,I676879,I676792);
nand I_39659 (I676545,I676879,I676701);
nor I_39660 (I676927,I26389,I26377);
and I_39661 (I676944,I676792,I676927);
nor I_39662 (I676961,I676879,I676944);
DFFARX1 I_39663 (I676961,I2683,I676568,I676554,);
nor I_39664 (I676992,I676594,I676927);
DFFARX1 I_39665 (I676992,I2683,I676568,I676539,);
nor I_39666 (I677023,I676871,I676927);
not I_39667 (I677040,I677023);
nand I_39668 (I676548,I677040,I676896);
not I_39669 (I677095,I2690);
DFFARX1 I_39670 (I101759,I2683,I677095,I677121,);
not I_39671 (I677129,I677121);
nand I_39672 (I677146,I101735,I101744);
and I_39673 (I677163,I677146,I101738);
DFFARX1 I_39674 (I677163,I2683,I677095,I677189,);
DFFARX1 I_39675 (I677189,I2683,I677095,I677084,);
DFFARX1 I_39676 (I101756,I2683,I677095,I677220,);
nand I_39677 (I677228,I677220,I101747);
not I_39678 (I677245,I677228);
DFFARX1 I_39679 (I677245,I2683,I677095,I677271,);
not I_39680 (I677279,I677271);
nor I_39681 (I677087,I677129,I677279);
DFFARX1 I_39682 (I101741,I2683,I677095,I677319,);
nor I_39683 (I677078,I677319,I677189);
nor I_39684 (I677069,I677319,I677245);
nand I_39685 (I677355,I101753,I101750);
and I_39686 (I677372,I677355,I101738);
DFFARX1 I_39687 (I677372,I2683,I677095,I677398,);
not I_39688 (I677406,I677398);
nand I_39689 (I677423,I677406,I677319);
nand I_39690 (I677072,I677406,I677228);
nor I_39691 (I677454,I101735,I101750);
and I_39692 (I677471,I677319,I677454);
nor I_39693 (I677488,I677406,I677471);
DFFARX1 I_39694 (I677488,I2683,I677095,I677081,);
nor I_39695 (I677519,I677121,I677454);
DFFARX1 I_39696 (I677519,I2683,I677095,I677066,);
nor I_39697 (I677550,I677398,I677454);
not I_39698 (I677567,I677550);
nand I_39699 (I677075,I677567,I677423);
not I_39700 (I677622,I2690);
DFFARX1 I_39701 (I378552,I2683,I677622,I677648,);
not I_39702 (I677656,I677648);
nand I_39703 (I677673,I378549,I378558);
and I_39704 (I677690,I677673,I378567);
DFFARX1 I_39705 (I677690,I2683,I677622,I677716,);
DFFARX1 I_39706 (I677716,I2683,I677622,I677611,);
DFFARX1 I_39707 (I378570,I2683,I677622,I677747,);
nand I_39708 (I677755,I677747,I378573);
not I_39709 (I677772,I677755);
DFFARX1 I_39710 (I677772,I2683,I677622,I677798,);
not I_39711 (I677806,I677798);
nor I_39712 (I677614,I677656,I677806);
DFFARX1 I_39713 (I378546,I2683,I677622,I677846,);
nor I_39714 (I677605,I677846,I677716);
nor I_39715 (I677596,I677846,I677772);
nand I_39716 (I677882,I378561,I378564);
and I_39717 (I677899,I677882,I378555);
DFFARX1 I_39718 (I677899,I2683,I677622,I677925,);
not I_39719 (I677933,I677925);
nand I_39720 (I677950,I677933,I677846);
nand I_39721 (I677599,I677933,I677755);
nor I_39722 (I677981,I378546,I378564);
and I_39723 (I677998,I677846,I677981);
nor I_39724 (I678015,I677933,I677998);
DFFARX1 I_39725 (I678015,I2683,I677622,I677608,);
nor I_39726 (I678046,I677648,I677981);
DFFARX1 I_39727 (I678046,I2683,I677622,I677593,);
nor I_39728 (I678077,I677925,I677981);
not I_39729 (I678094,I678077);
nand I_39730 (I677602,I678094,I677950);
not I_39731 (I678149,I2690);
DFFARX1 I_39732 (I1041204,I2683,I678149,I678175,);
not I_39733 (I678183,I678175);
nand I_39734 (I678200,I1041201,I1041210);
and I_39735 (I678217,I678200,I1041189);
DFFARX1 I_39736 (I678217,I2683,I678149,I678243,);
DFFARX1 I_39737 (I678243,I2683,I678149,I678138,);
DFFARX1 I_39738 (I1041192,I2683,I678149,I678274,);
nand I_39739 (I678282,I678274,I1041207);
not I_39740 (I678299,I678282);
DFFARX1 I_39741 (I678299,I2683,I678149,I678325,);
not I_39742 (I678333,I678325);
nor I_39743 (I678141,I678183,I678333);
DFFARX1 I_39744 (I1041213,I2683,I678149,I678373,);
nor I_39745 (I678132,I678373,I678243);
nor I_39746 (I678123,I678373,I678299);
nand I_39747 (I678409,I1041195,I1041216);
and I_39748 (I678426,I678409,I1041198);
DFFARX1 I_39749 (I678426,I2683,I678149,I678452,);
not I_39750 (I678460,I678452);
nand I_39751 (I678477,I678460,I678373);
nand I_39752 (I678126,I678460,I678282);
nor I_39753 (I678508,I1041189,I1041216);
and I_39754 (I678525,I678373,I678508);
nor I_39755 (I678542,I678460,I678525);
DFFARX1 I_39756 (I678542,I2683,I678149,I678135,);
nor I_39757 (I678573,I678175,I678508);
DFFARX1 I_39758 (I678573,I2683,I678149,I678120,);
nor I_39759 (I678604,I678452,I678508);
not I_39760 (I678621,I678604);
nand I_39761 (I678129,I678621,I678477);
not I_39762 (I678676,I2690);
DFFARX1 I_39763 (I302293,I2683,I678676,I678702,);
not I_39764 (I678710,I678702);
nand I_39765 (I678727,I302284,I302284);
and I_39766 (I678744,I678727,I302302);
DFFARX1 I_39767 (I678744,I2683,I678676,I678770,);
DFFARX1 I_39768 (I678770,I2683,I678676,I678665,);
DFFARX1 I_39769 (I302305,I2683,I678676,I678801,);
nand I_39770 (I678809,I678801,I302287);
not I_39771 (I678826,I678809);
DFFARX1 I_39772 (I678826,I2683,I678676,I678852,);
not I_39773 (I678860,I678852);
nor I_39774 (I678668,I678710,I678860);
DFFARX1 I_39775 (I302299,I2683,I678676,I678900,);
nor I_39776 (I678659,I678900,I678770);
nor I_39777 (I678650,I678900,I678826);
nand I_39778 (I678936,I302311,I302290);
and I_39779 (I678953,I678936,I302296);
DFFARX1 I_39780 (I678953,I2683,I678676,I678979,);
not I_39781 (I678987,I678979);
nand I_39782 (I679004,I678987,I678900);
nand I_39783 (I678653,I678987,I678809);
nor I_39784 (I679035,I302308,I302290);
and I_39785 (I679052,I678900,I679035);
nor I_39786 (I679069,I678987,I679052);
DFFARX1 I_39787 (I679069,I2683,I678676,I678662,);
nor I_39788 (I679100,I678702,I679035);
DFFARX1 I_39789 (I679100,I2683,I678676,I678647,);
nor I_39790 (I679131,I678979,I679035);
not I_39791 (I679148,I679131);
nand I_39792 (I678656,I679148,I679004);
not I_39793 (I679203,I2690);
DFFARX1 I_39794 (I776842,I2683,I679203,I679229,);
not I_39795 (I679237,I679229);
nand I_39796 (I679254,I776857,I776839);
and I_39797 (I679271,I679254,I776839);
DFFARX1 I_39798 (I679271,I2683,I679203,I679297,);
DFFARX1 I_39799 (I679297,I2683,I679203,I679192,);
DFFARX1 I_39800 (I776848,I2683,I679203,I679328,);
nand I_39801 (I679336,I679328,I776866);
not I_39802 (I679353,I679336);
DFFARX1 I_39803 (I679353,I2683,I679203,I679379,);
not I_39804 (I679387,I679379);
nor I_39805 (I679195,I679237,I679387);
DFFARX1 I_39806 (I776863,I2683,I679203,I679427,);
nor I_39807 (I679186,I679427,I679297);
nor I_39808 (I679177,I679427,I679353);
nand I_39809 (I679463,I776860,I776851);
and I_39810 (I679480,I679463,I776845);
DFFARX1 I_39811 (I679480,I2683,I679203,I679506,);
not I_39812 (I679514,I679506);
nand I_39813 (I679531,I679514,I679427);
nand I_39814 (I679180,I679514,I679336);
nor I_39815 (I679562,I776854,I776851);
and I_39816 (I679579,I679427,I679562);
nor I_39817 (I679596,I679514,I679579);
DFFARX1 I_39818 (I679596,I2683,I679203,I679189,);
nor I_39819 (I679627,I679229,I679562);
DFFARX1 I_39820 (I679627,I2683,I679203,I679174,);
nor I_39821 (I679658,I679506,I679562);
not I_39822 (I679675,I679658);
nand I_39823 (I679183,I679675,I679531);
not I_39824 (I679730,I2690);
DFFARX1 I_39825 (I528350,I2683,I679730,I679756,);
not I_39826 (I679764,I679756);
nand I_39827 (I679781,I528353,I528350);
and I_39828 (I679798,I679781,I528362);
DFFARX1 I_39829 (I679798,I2683,I679730,I679824,);
DFFARX1 I_39830 (I679824,I2683,I679730,I679719,);
DFFARX1 I_39831 (I528359,I2683,I679730,I679855,);
nand I_39832 (I679863,I679855,I528365);
not I_39833 (I679880,I679863);
DFFARX1 I_39834 (I679880,I2683,I679730,I679906,);
not I_39835 (I679914,I679906);
nor I_39836 (I679722,I679764,I679914);
DFFARX1 I_39837 (I528374,I2683,I679730,I679954,);
nor I_39838 (I679713,I679954,I679824);
nor I_39839 (I679704,I679954,I679880);
nand I_39840 (I679990,I528368,I528356);
and I_39841 (I680007,I679990,I528353);
DFFARX1 I_39842 (I680007,I2683,I679730,I680033,);
not I_39843 (I680041,I680033);
nand I_39844 (I680058,I680041,I679954);
nand I_39845 (I679707,I680041,I679863);
nor I_39846 (I680089,I528371,I528356);
and I_39847 (I680106,I679954,I680089);
nor I_39848 (I680123,I680041,I680106);
DFFARX1 I_39849 (I680123,I2683,I679730,I679716,);
nor I_39850 (I680154,I679756,I680089);
DFFARX1 I_39851 (I680154,I2683,I679730,I679701,);
nor I_39852 (I680185,I680033,I680089);
not I_39853 (I680202,I680185);
nand I_39854 (I679710,I680202,I680058);
not I_39855 (I680257,I2690);
DFFARX1 I_39856 (I850756,I2683,I680257,I680283,);
not I_39857 (I680291,I680283);
nand I_39858 (I680308,I850738,I850738);
and I_39859 (I680325,I680308,I850744);
DFFARX1 I_39860 (I680325,I2683,I680257,I680351,);
DFFARX1 I_39861 (I680351,I2683,I680257,I680246,);
DFFARX1 I_39862 (I850741,I2683,I680257,I680382,);
nand I_39863 (I680390,I680382,I850750);
not I_39864 (I680407,I680390);
DFFARX1 I_39865 (I680407,I2683,I680257,I680433,);
not I_39866 (I680441,I680433);
nor I_39867 (I680249,I680291,I680441);
DFFARX1 I_39868 (I850762,I2683,I680257,I680481,);
nor I_39869 (I680240,I680481,I680351);
nor I_39870 (I680231,I680481,I680407);
nand I_39871 (I680517,I850753,I850747);
and I_39872 (I680534,I680517,I850741);
DFFARX1 I_39873 (I680534,I2683,I680257,I680560,);
not I_39874 (I680568,I680560);
nand I_39875 (I680585,I680568,I680481);
nand I_39876 (I680234,I680568,I680390);
nor I_39877 (I680616,I850759,I850747);
and I_39878 (I680633,I680481,I680616);
nor I_39879 (I680650,I680568,I680633);
DFFARX1 I_39880 (I680650,I2683,I680257,I680243,);
nor I_39881 (I680681,I680283,I680616);
DFFARX1 I_39882 (I680681,I2683,I680257,I680228,);
nor I_39883 (I680712,I680560,I680616);
not I_39884 (I680729,I680712);
nand I_39885 (I680237,I680729,I680585);
not I_39886 (I680784,I2690);
DFFARX1 I_39887 (I1080474,I2683,I680784,I680810,);
not I_39888 (I680818,I680810);
nand I_39889 (I680835,I1080471,I1080480);
and I_39890 (I680852,I680835,I1080459);
DFFARX1 I_39891 (I680852,I2683,I680784,I680878,);
DFFARX1 I_39892 (I680878,I2683,I680784,I680773,);
DFFARX1 I_39893 (I1080462,I2683,I680784,I680909,);
nand I_39894 (I680917,I680909,I1080477);
not I_39895 (I680934,I680917);
DFFARX1 I_39896 (I680934,I2683,I680784,I680960,);
not I_39897 (I680968,I680960);
nor I_39898 (I680776,I680818,I680968);
DFFARX1 I_39899 (I1080483,I2683,I680784,I681008,);
nor I_39900 (I680767,I681008,I680878);
nor I_39901 (I680758,I681008,I680934);
nand I_39902 (I681044,I1080465,I1080486);
and I_39903 (I681061,I681044,I1080468);
DFFARX1 I_39904 (I681061,I2683,I680784,I681087,);
not I_39905 (I681095,I681087);
nand I_39906 (I681112,I681095,I681008);
nand I_39907 (I680761,I681095,I680917);
nor I_39908 (I681143,I1080459,I1080486);
and I_39909 (I681160,I681008,I681143);
nor I_39910 (I681177,I681095,I681160);
DFFARX1 I_39911 (I681177,I2683,I680784,I680770,);
nor I_39912 (I681208,I680810,I681143);
DFFARX1 I_39913 (I681208,I2683,I680784,I680755,);
nor I_39914 (I681239,I681087,I681143);
not I_39915 (I681256,I681239);
nand I_39916 (I680764,I681256,I681112);
not I_39917 (I681311,I2690);
DFFARX1 I_39918 (I303874,I2683,I681311,I681337,);
not I_39919 (I681345,I681337);
nand I_39920 (I681362,I303865,I303865);
and I_39921 (I681379,I681362,I303883);
DFFARX1 I_39922 (I681379,I2683,I681311,I681405,);
DFFARX1 I_39923 (I681405,I2683,I681311,I681300,);
DFFARX1 I_39924 (I303886,I2683,I681311,I681436,);
nand I_39925 (I681444,I681436,I303868);
not I_39926 (I681461,I681444);
DFFARX1 I_39927 (I681461,I2683,I681311,I681487,);
not I_39928 (I681495,I681487);
nor I_39929 (I681303,I681345,I681495);
DFFARX1 I_39930 (I303880,I2683,I681311,I681535,);
nor I_39931 (I681294,I681535,I681405);
nor I_39932 (I681285,I681535,I681461);
nand I_39933 (I681571,I303892,I303871);
and I_39934 (I681588,I681571,I303877);
DFFARX1 I_39935 (I681588,I2683,I681311,I681614,);
not I_39936 (I681622,I681614);
nand I_39937 (I681639,I681622,I681535);
nand I_39938 (I681288,I681622,I681444);
nor I_39939 (I681670,I303889,I303871);
and I_39940 (I681687,I681535,I681670);
nor I_39941 (I681704,I681622,I681687);
DFFARX1 I_39942 (I681704,I2683,I681311,I681297,);
nor I_39943 (I681735,I681337,I681670);
DFFARX1 I_39944 (I681735,I2683,I681311,I681282,);
nor I_39945 (I681766,I681614,I681670);
not I_39946 (I681783,I681766);
nand I_39947 (I681291,I681783,I681639);
not I_39948 (I681838,I2690);
DFFARX1 I_39949 (I792992,I2683,I681838,I681864,);
not I_39950 (I681872,I681864);
nand I_39951 (I681889,I793007,I792989);
and I_39952 (I681906,I681889,I792989);
DFFARX1 I_39953 (I681906,I2683,I681838,I681932,);
DFFARX1 I_39954 (I681932,I2683,I681838,I681827,);
DFFARX1 I_39955 (I792998,I2683,I681838,I681963,);
nand I_39956 (I681971,I681963,I793016);
not I_39957 (I681988,I681971);
DFFARX1 I_39958 (I681988,I2683,I681838,I682014,);
not I_39959 (I682022,I682014);
nor I_39960 (I681830,I681872,I682022);
DFFARX1 I_39961 (I793013,I2683,I681838,I682062,);
nor I_39962 (I681821,I682062,I681932);
nor I_39963 (I681812,I682062,I681988);
nand I_39964 (I682098,I793010,I793001);
and I_39965 (I682115,I682098,I792995);
DFFARX1 I_39966 (I682115,I2683,I681838,I682141,);
not I_39967 (I682149,I682141);
nand I_39968 (I682166,I682149,I682062);
nand I_39969 (I681815,I682149,I681971);
nor I_39970 (I682197,I793004,I793001);
and I_39971 (I682214,I682062,I682197);
nor I_39972 (I682231,I682149,I682214);
DFFARX1 I_39973 (I682231,I2683,I681838,I681824,);
nor I_39974 (I682262,I681864,I682197);
DFFARX1 I_39975 (I682262,I2683,I681838,I681809,);
nor I_39976 (I682293,I682141,I682197);
not I_39977 (I682310,I682293);
nand I_39978 (I681818,I682310,I682166);
not I_39979 (I682365,I2690);
DFFARX1 I_39980 (I1029363,I2683,I682365,I682391,);
not I_39981 (I682399,I682391);
nand I_39982 (I682416,I1029357,I1029375);
and I_39983 (I682433,I682416,I1029360);
DFFARX1 I_39984 (I682433,I2683,I682365,I682459,);
DFFARX1 I_39985 (I682459,I2683,I682365,I682354,);
DFFARX1 I_39986 (I1029381,I2683,I682365,I682490,);
nand I_39987 (I682498,I682490,I1029366);
not I_39988 (I682515,I682498);
DFFARX1 I_39989 (I682515,I2683,I682365,I682541,);
not I_39990 (I682549,I682541);
nor I_39991 (I682357,I682399,I682549);
DFFARX1 I_39992 (I1029378,I2683,I682365,I682589,);
nor I_39993 (I682348,I682589,I682459);
nor I_39994 (I682339,I682589,I682515);
nand I_39995 (I682625,I1029369,I1029384);
and I_39996 (I682642,I682625,I1029372);
DFFARX1 I_39997 (I682642,I2683,I682365,I682668,);
not I_39998 (I682676,I682668);
nand I_39999 (I682693,I682676,I682589);
nand I_40000 (I682342,I682676,I682498);
nor I_40001 (I682724,I1029357,I1029384);
and I_40002 (I682741,I682589,I682724);
nor I_40003 (I682758,I682676,I682741);
DFFARX1 I_40004 (I682758,I2683,I682365,I682351,);
nor I_40005 (I682789,I682391,I682724);
DFFARX1 I_40006 (I682789,I2683,I682365,I682336,);
nor I_40007 (I682820,I682668,I682724);
not I_40008 (I682837,I682820);
nand I_40009 (I682345,I682837,I682693);
not I_40010 (I682892,I2690);
DFFARX1 I_40011 (I160476,I2683,I682892,I682918,);
not I_40012 (I682926,I682918);
nand I_40013 (I682943,I160473,I160491);
and I_40014 (I682960,I682943,I160482);
DFFARX1 I_40015 (I682960,I2683,I682892,I682986,);
DFFARX1 I_40016 (I682986,I2683,I682892,I682881,);
DFFARX1 I_40017 (I160488,I2683,I682892,I683017,);
nand I_40018 (I683025,I683017,I160485);
not I_40019 (I683042,I683025);
DFFARX1 I_40020 (I683042,I2683,I682892,I683068,);
not I_40021 (I683076,I683068);
nor I_40022 (I682884,I682926,I683076);
DFFARX1 I_40023 (I160479,I2683,I682892,I683116,);
nor I_40024 (I682875,I683116,I682986);
nor I_40025 (I682866,I683116,I683042);
nand I_40026 (I683152,I160470,I160494);
and I_40027 (I683169,I683152,I160473);
DFFARX1 I_40028 (I683169,I2683,I682892,I683195,);
not I_40029 (I683203,I683195);
nand I_40030 (I683220,I683203,I683116);
nand I_40031 (I682869,I683203,I683025);
nor I_40032 (I683251,I160470,I160494);
and I_40033 (I683268,I683116,I683251);
nor I_40034 (I683285,I683203,I683268);
DFFARX1 I_40035 (I683285,I2683,I682892,I682878,);
nor I_40036 (I683316,I682918,I683251);
DFFARX1 I_40037 (I683316,I2683,I682892,I682863,);
nor I_40038 (I683347,I683195,I683251);
not I_40039 (I683364,I683347);
nand I_40040 (I682872,I683364,I683220);
not I_40041 (I683419,I2690);
DFFARX1 I_40042 (I937456,I2683,I683419,I683445,);
not I_40043 (I683453,I683445);
nand I_40044 (I683470,I937438,I937438);
and I_40045 (I683487,I683470,I937444);
DFFARX1 I_40046 (I683487,I2683,I683419,I683513,);
DFFARX1 I_40047 (I683513,I2683,I683419,I683408,);
DFFARX1 I_40048 (I937441,I2683,I683419,I683544,);
nand I_40049 (I683552,I683544,I937450);
not I_40050 (I683569,I683552);
DFFARX1 I_40051 (I683569,I2683,I683419,I683595,);
not I_40052 (I683603,I683595);
nor I_40053 (I683411,I683453,I683603);
DFFARX1 I_40054 (I937462,I2683,I683419,I683643,);
nor I_40055 (I683402,I683643,I683513);
nor I_40056 (I683393,I683643,I683569);
nand I_40057 (I683679,I937453,I937447);
and I_40058 (I683696,I683679,I937441);
DFFARX1 I_40059 (I683696,I2683,I683419,I683722,);
not I_40060 (I683730,I683722);
nand I_40061 (I683747,I683730,I683643);
nand I_40062 (I683396,I683730,I683552);
nor I_40063 (I683778,I937459,I937447);
and I_40064 (I683795,I683643,I683778);
nor I_40065 (I683812,I683730,I683795);
DFFARX1 I_40066 (I683812,I2683,I683419,I683405,);
nor I_40067 (I683843,I683445,I683778);
DFFARX1 I_40068 (I683843,I2683,I683419,I683390,);
nor I_40069 (I683874,I683722,I683778);
not I_40070 (I683891,I683874);
nand I_40071 (I683399,I683891,I683747);
not I_40072 (I683946,I2690);
DFFARX1 I_40073 (I217446,I2683,I683946,I683972,);
not I_40074 (I683980,I683972);
nand I_40075 (I683997,I217437,I217437);
and I_40076 (I684014,I683997,I217455);
DFFARX1 I_40077 (I684014,I2683,I683946,I684040,);
DFFARX1 I_40078 (I684040,I2683,I683946,I683935,);
DFFARX1 I_40079 (I217458,I2683,I683946,I684071,);
nand I_40080 (I684079,I684071,I217440);
not I_40081 (I684096,I684079);
DFFARX1 I_40082 (I684096,I2683,I683946,I684122,);
not I_40083 (I684130,I684122);
nor I_40084 (I683938,I683980,I684130);
DFFARX1 I_40085 (I217452,I2683,I683946,I684170,);
nor I_40086 (I683929,I684170,I684040);
nor I_40087 (I683920,I684170,I684096);
nand I_40088 (I684206,I217464,I217443);
and I_40089 (I684223,I684206,I217449);
DFFARX1 I_40090 (I684223,I2683,I683946,I684249,);
not I_40091 (I684257,I684249);
nand I_40092 (I684274,I684257,I684170);
nand I_40093 (I683923,I684257,I684079);
nor I_40094 (I684305,I217461,I217443);
and I_40095 (I684322,I684170,I684305);
nor I_40096 (I684339,I684257,I684322);
DFFARX1 I_40097 (I684339,I2683,I683946,I683932,);
nor I_40098 (I684370,I683972,I684305);
DFFARX1 I_40099 (I684370,I2683,I683946,I683917,);
nor I_40100 (I684401,I684249,I684305);
not I_40101 (I684418,I684401);
nand I_40102 (I683926,I684418,I684274);
not I_40103 (I684473,I2690);
DFFARX1 I_40104 (I598288,I2683,I684473,I684499,);
not I_40105 (I684507,I684499);
nand I_40106 (I684524,I598291,I598288);
and I_40107 (I684541,I684524,I598300);
DFFARX1 I_40108 (I684541,I2683,I684473,I684567,);
DFFARX1 I_40109 (I684567,I2683,I684473,I684462,);
DFFARX1 I_40110 (I598297,I2683,I684473,I684598,);
nand I_40111 (I684606,I684598,I598303);
not I_40112 (I684623,I684606);
DFFARX1 I_40113 (I684623,I2683,I684473,I684649,);
not I_40114 (I684657,I684649);
nor I_40115 (I684465,I684507,I684657);
DFFARX1 I_40116 (I598312,I2683,I684473,I684697,);
nor I_40117 (I684456,I684697,I684567);
nor I_40118 (I684447,I684697,I684623);
nand I_40119 (I684733,I598306,I598294);
and I_40120 (I684750,I684733,I598291);
DFFARX1 I_40121 (I684750,I2683,I684473,I684776,);
not I_40122 (I684784,I684776);
nand I_40123 (I684801,I684784,I684697);
nand I_40124 (I684450,I684784,I684606);
nor I_40125 (I684832,I598309,I598294);
and I_40126 (I684849,I684697,I684832);
nor I_40127 (I684866,I684784,I684849);
DFFARX1 I_40128 (I684866,I2683,I684473,I684459,);
nor I_40129 (I684897,I684499,I684832);
DFFARX1 I_40130 (I684897,I2683,I684473,I684444,);
nor I_40131 (I684928,I684776,I684832);
not I_40132 (I684945,I684928);
nand I_40133 (I684453,I684945,I684801);
not I_40134 (I685000,I2690);
DFFARX1 I_40135 (I970090,I2683,I685000,I685026,);
not I_40136 (I685034,I685026);
nand I_40137 (I685051,I970096,I970078);
and I_40138 (I685068,I685051,I970087);
DFFARX1 I_40139 (I685068,I2683,I685000,I685094,);
DFFARX1 I_40140 (I685094,I2683,I685000,I684989,);
DFFARX1 I_40141 (I970093,I2683,I685000,I685125,);
nand I_40142 (I685133,I685125,I970081);
not I_40143 (I685150,I685133);
DFFARX1 I_40144 (I685150,I2683,I685000,I685176,);
not I_40145 (I685184,I685176);
nor I_40146 (I684992,I685034,I685184);
DFFARX1 I_40147 (I970099,I2683,I685000,I685224,);
nor I_40148 (I684983,I685224,I685094);
nor I_40149 (I684974,I685224,I685150);
nand I_40150 (I685260,I970078,I970084);
and I_40151 (I685277,I685260,I970102);
DFFARX1 I_40152 (I685277,I2683,I685000,I685303,);
not I_40153 (I685311,I685303);
nand I_40154 (I685328,I685311,I685224);
nand I_40155 (I684977,I685311,I685133);
nor I_40156 (I685359,I970081,I970084);
and I_40157 (I685376,I685224,I685359);
nor I_40158 (I685393,I685311,I685376);
DFFARX1 I_40159 (I685393,I2683,I685000,I684986,);
nor I_40160 (I685424,I685026,I685359);
DFFARX1 I_40161 (I685424,I2683,I685000,I684971,);
nor I_40162 (I685455,I685303,I685359);
not I_40163 (I685472,I685455);
nand I_40164 (I684980,I685472,I685328);
not I_40165 (I685527,I2690);
DFFARX1 I_40166 (I1004776,I2683,I685527,I685553,);
not I_40167 (I685561,I685553);
nand I_40168 (I685578,I1004758,I1004761);
and I_40169 (I685595,I685578,I1004773);
DFFARX1 I_40170 (I685595,I2683,I685527,I685621,);
DFFARX1 I_40171 (I685621,I2683,I685527,I685516,);
DFFARX1 I_40172 (I1004782,I2683,I685527,I685652,);
nand I_40173 (I685660,I685652,I1004767);
not I_40174 (I685677,I685660);
DFFARX1 I_40175 (I685677,I2683,I685527,I685703,);
not I_40176 (I685711,I685703);
nor I_40177 (I685519,I685561,I685711);
DFFARX1 I_40178 (I1004779,I2683,I685527,I685751,);
nor I_40179 (I685510,I685751,I685621);
nor I_40180 (I685501,I685751,I685677);
nand I_40181 (I685787,I1004770,I1004764);
and I_40182 (I685804,I685787,I1004758);
DFFARX1 I_40183 (I685804,I2683,I685527,I685830,);
not I_40184 (I685838,I685830);
nand I_40185 (I685855,I685838,I685751);
nand I_40186 (I685504,I685838,I685660);
nor I_40187 (I685886,I1004761,I1004764);
and I_40188 (I685903,I685751,I685886);
nor I_40189 (I685920,I685838,I685903);
DFFARX1 I_40190 (I685920,I2683,I685527,I685513,);
nor I_40191 (I685951,I685553,I685886);
DFFARX1 I_40192 (I685951,I2683,I685527,I685498,);
nor I_40193 (I685982,I685830,I685886);
not I_40194 (I685999,I685982);
nand I_40195 (I685507,I685999,I685855);
not I_40196 (I686054,I2690);
DFFARX1 I_40197 (I203911,I2683,I686054,I686080,);
not I_40198 (I686088,I686080);
nand I_40199 (I686105,I203908,I203926);
and I_40200 (I686122,I686105,I203917);
DFFARX1 I_40201 (I686122,I2683,I686054,I686148,);
DFFARX1 I_40202 (I686148,I2683,I686054,I686043,);
DFFARX1 I_40203 (I203923,I2683,I686054,I686179,);
nand I_40204 (I686187,I686179,I203920);
not I_40205 (I686204,I686187);
DFFARX1 I_40206 (I686204,I2683,I686054,I686230,);
not I_40207 (I686238,I686230);
nor I_40208 (I686046,I686088,I686238);
DFFARX1 I_40209 (I203914,I2683,I686054,I686278,);
nor I_40210 (I686037,I686278,I686148);
nor I_40211 (I686028,I686278,I686204);
nand I_40212 (I686314,I203905,I203929);
and I_40213 (I686331,I686314,I203908);
DFFARX1 I_40214 (I686331,I2683,I686054,I686357,);
not I_40215 (I686365,I686357);
nand I_40216 (I686382,I686365,I686278);
nand I_40217 (I686031,I686365,I686187);
nor I_40218 (I686413,I203905,I203929);
and I_40219 (I686430,I686278,I686413);
nor I_40220 (I686447,I686365,I686430);
DFFARX1 I_40221 (I686447,I2683,I686054,I686040,);
nor I_40222 (I686478,I686080,I686413);
DFFARX1 I_40223 (I686478,I2683,I686054,I686025,);
nor I_40224 (I686509,I686357,I686413);
not I_40225 (I686526,I686509);
nand I_40226 (I686034,I686526,I686382);
not I_40227 (I686581,I2690);
DFFARX1 I_40228 (I509854,I2683,I686581,I686607,);
not I_40229 (I686615,I686607);
nand I_40230 (I686632,I509857,I509854);
and I_40231 (I686649,I686632,I509866);
DFFARX1 I_40232 (I686649,I2683,I686581,I686675,);
DFFARX1 I_40233 (I686675,I2683,I686581,I686570,);
DFFARX1 I_40234 (I509863,I2683,I686581,I686706,);
nand I_40235 (I686714,I686706,I509869);
not I_40236 (I686731,I686714);
DFFARX1 I_40237 (I686731,I2683,I686581,I686757,);
not I_40238 (I686765,I686757);
nor I_40239 (I686573,I686615,I686765);
DFFARX1 I_40240 (I509878,I2683,I686581,I686805,);
nor I_40241 (I686564,I686805,I686675);
nor I_40242 (I686555,I686805,I686731);
nand I_40243 (I686841,I509872,I509860);
and I_40244 (I686858,I686841,I509857);
DFFARX1 I_40245 (I686858,I2683,I686581,I686884,);
not I_40246 (I686892,I686884);
nand I_40247 (I686909,I686892,I686805);
nand I_40248 (I686558,I686892,I686714);
nor I_40249 (I686940,I509875,I509860);
and I_40250 (I686957,I686805,I686940);
nor I_40251 (I686974,I686892,I686957);
DFFARX1 I_40252 (I686974,I2683,I686581,I686567,);
nor I_40253 (I687005,I686607,I686940);
DFFARX1 I_40254 (I687005,I2683,I686581,I686552,);
nor I_40255 (I687036,I686884,I686940);
not I_40256 (I687053,I687036);
nand I_40257 (I686561,I687053,I686909);
not I_40258 (I687108,I2690);
DFFARX1 I_40259 (I180706,I2683,I687108,I687134,);
not I_40260 (I687142,I687134);
nand I_40261 (I687159,I180703,I180721);
and I_40262 (I687176,I687159,I180712);
DFFARX1 I_40263 (I687176,I2683,I687108,I687202,);
DFFARX1 I_40264 (I687202,I2683,I687108,I687097,);
DFFARX1 I_40265 (I180718,I2683,I687108,I687233,);
nand I_40266 (I687241,I687233,I180715);
not I_40267 (I687258,I687241);
DFFARX1 I_40268 (I687258,I2683,I687108,I687284,);
not I_40269 (I687292,I687284);
nor I_40270 (I687100,I687142,I687292);
DFFARX1 I_40271 (I180709,I2683,I687108,I687332,);
nor I_40272 (I687091,I687332,I687202);
nor I_40273 (I687082,I687332,I687258);
nand I_40274 (I687368,I180700,I180724);
and I_40275 (I687385,I687368,I180703);
DFFARX1 I_40276 (I687385,I2683,I687108,I687411,);
not I_40277 (I687419,I687411);
nand I_40278 (I687436,I687419,I687332);
nand I_40279 (I687085,I687419,I687241);
nor I_40280 (I687467,I180700,I180724);
and I_40281 (I687484,I687332,I687467);
nor I_40282 (I687501,I687419,I687484);
DFFARX1 I_40283 (I687501,I2683,I687108,I687094,);
nor I_40284 (I687532,I687134,I687467);
DFFARX1 I_40285 (I687532,I2683,I687108,I687079,);
nor I_40286 (I687563,I687411,I687467);
not I_40287 (I687580,I687563);
nand I_40288 (I687088,I687580,I687436);
not I_40289 (I687635,I2690);
DFFARX1 I_40290 (I208671,I2683,I687635,I687661,);
not I_40291 (I687669,I687661);
nand I_40292 (I687686,I208668,I208686);
and I_40293 (I687703,I687686,I208677);
DFFARX1 I_40294 (I687703,I2683,I687635,I687729,);
DFFARX1 I_40295 (I687729,I2683,I687635,I687624,);
DFFARX1 I_40296 (I208683,I2683,I687635,I687760,);
nand I_40297 (I687768,I687760,I208680);
not I_40298 (I687785,I687768);
DFFARX1 I_40299 (I687785,I2683,I687635,I687811,);
not I_40300 (I687819,I687811);
nor I_40301 (I687627,I687669,I687819);
DFFARX1 I_40302 (I208674,I2683,I687635,I687859,);
nor I_40303 (I687618,I687859,I687729);
nor I_40304 (I687609,I687859,I687785);
nand I_40305 (I687895,I208665,I208689);
and I_40306 (I687912,I687895,I208668);
DFFARX1 I_40307 (I687912,I2683,I687635,I687938,);
not I_40308 (I687946,I687938);
nand I_40309 (I687963,I687946,I687859);
nand I_40310 (I687612,I687946,I687768);
nor I_40311 (I687994,I208665,I208689);
and I_40312 (I688011,I687859,I687994);
nor I_40313 (I688028,I687946,I688011);
DFFARX1 I_40314 (I688028,I2683,I687635,I687621,);
nor I_40315 (I688059,I687661,I687994);
DFFARX1 I_40316 (I688059,I2683,I687635,I687606,);
nor I_40317 (I688090,I687938,I687994);
not I_40318 (I688107,I688090);
nand I_40319 (I687615,I688107,I687963);
not I_40320 (I688162,I2690);
DFFARX1 I_40321 (I430623,I2683,I688162,I688188,);
not I_40322 (I688196,I688188);
nand I_40323 (I688213,I430641,I430632);
and I_40324 (I688230,I688213,I430635);
DFFARX1 I_40325 (I688230,I2683,I688162,I688256,);
DFFARX1 I_40326 (I688256,I2683,I688162,I688151,);
DFFARX1 I_40327 (I430629,I2683,I688162,I688287,);
nand I_40328 (I688295,I688287,I430620);
not I_40329 (I688312,I688295);
DFFARX1 I_40330 (I688312,I2683,I688162,I688338,);
not I_40331 (I688346,I688338);
nor I_40332 (I688154,I688196,I688346);
DFFARX1 I_40333 (I430626,I2683,I688162,I688386,);
nor I_40334 (I688145,I688386,I688256);
nor I_40335 (I688136,I688386,I688312);
nand I_40336 (I688422,I430620,I430617);
and I_40337 (I688439,I688422,I430638);
DFFARX1 I_40338 (I688439,I2683,I688162,I688465,);
not I_40339 (I688473,I688465);
nand I_40340 (I688490,I688473,I688386);
nand I_40341 (I688139,I688473,I688295);
nor I_40342 (I688521,I430617,I430617);
and I_40343 (I688538,I688386,I688521);
nor I_40344 (I688555,I688473,I688538);
DFFARX1 I_40345 (I688555,I2683,I688162,I688148,);
nor I_40346 (I688586,I688188,I688521);
DFFARX1 I_40347 (I688586,I2683,I688162,I688133,);
nor I_40348 (I688617,I688465,I688521);
not I_40349 (I688634,I688617);
nand I_40350 (I688142,I688634,I688490);
not I_40351 (I688689,I2690);
DFFARX1 I_40352 (I782010,I2683,I688689,I688715,);
not I_40353 (I688723,I688715);
nand I_40354 (I688740,I782025,I782007);
and I_40355 (I688757,I688740,I782007);
DFFARX1 I_40356 (I688757,I2683,I688689,I688783,);
DFFARX1 I_40357 (I688783,I2683,I688689,I688678,);
DFFARX1 I_40358 (I782016,I2683,I688689,I688814,);
nand I_40359 (I688822,I688814,I782034);
not I_40360 (I688839,I688822);
DFFARX1 I_40361 (I688839,I2683,I688689,I688865,);
not I_40362 (I688873,I688865);
nor I_40363 (I688681,I688723,I688873);
DFFARX1 I_40364 (I782031,I2683,I688689,I688913,);
nor I_40365 (I688672,I688913,I688783);
nor I_40366 (I688663,I688913,I688839);
nand I_40367 (I688949,I782028,I782019);
and I_40368 (I688966,I688949,I782013);
DFFARX1 I_40369 (I688966,I2683,I688689,I688992,);
not I_40370 (I689000,I688992);
nand I_40371 (I689017,I689000,I688913);
nand I_40372 (I688666,I689000,I688822);
nor I_40373 (I689048,I782022,I782019);
and I_40374 (I689065,I688913,I689048);
nor I_40375 (I689082,I689000,I689065);
DFFARX1 I_40376 (I689082,I2683,I688689,I688675,);
nor I_40377 (I689113,I688715,I689048);
DFFARX1 I_40378 (I689113,I2683,I688689,I688660,);
nor I_40379 (I689144,I688992,I689048);
not I_40380 (I689161,I689144);
nand I_40381 (I688669,I689161,I689017);
not I_40382 (I689216,I2690);
DFFARX1 I_40383 (I54329,I2683,I689216,I689242,);
not I_40384 (I689250,I689242);
nand I_40385 (I689267,I54305,I54314);
and I_40386 (I689284,I689267,I54308);
DFFARX1 I_40387 (I689284,I2683,I689216,I689310,);
DFFARX1 I_40388 (I689310,I2683,I689216,I689205,);
DFFARX1 I_40389 (I54326,I2683,I689216,I689341,);
nand I_40390 (I689349,I689341,I54317);
not I_40391 (I689366,I689349);
DFFARX1 I_40392 (I689366,I2683,I689216,I689392,);
not I_40393 (I689400,I689392);
nor I_40394 (I689208,I689250,I689400);
DFFARX1 I_40395 (I54311,I2683,I689216,I689440,);
nor I_40396 (I689199,I689440,I689310);
nor I_40397 (I689190,I689440,I689366);
nand I_40398 (I689476,I54323,I54320);
and I_40399 (I689493,I689476,I54308);
DFFARX1 I_40400 (I689493,I2683,I689216,I689519,);
not I_40401 (I689527,I689519);
nand I_40402 (I689544,I689527,I689440);
nand I_40403 (I689193,I689527,I689349);
nor I_40404 (I689575,I54305,I54320);
and I_40405 (I689592,I689440,I689575);
nor I_40406 (I689609,I689527,I689592);
DFFARX1 I_40407 (I689609,I2683,I689216,I689202,);
nor I_40408 (I689640,I689242,I689575);
DFFARX1 I_40409 (I689640,I2683,I689216,I689187,);
nor I_40410 (I689671,I689519,I689575);
not I_40411 (I689688,I689671);
nand I_40412 (I689196,I689688,I689544);
not I_40413 (I689743,I2690);
DFFARX1 I_40414 (I576324,I2683,I689743,I689769,);
not I_40415 (I689777,I689769);
nand I_40416 (I689794,I576327,I576324);
and I_40417 (I689811,I689794,I576336);
DFFARX1 I_40418 (I689811,I2683,I689743,I689837,);
DFFARX1 I_40419 (I689837,I2683,I689743,I689732,);
DFFARX1 I_40420 (I576333,I2683,I689743,I689868,);
nand I_40421 (I689876,I689868,I576339);
not I_40422 (I689893,I689876);
DFFARX1 I_40423 (I689893,I2683,I689743,I689919,);
not I_40424 (I689927,I689919);
nor I_40425 (I689735,I689777,I689927);
DFFARX1 I_40426 (I576348,I2683,I689743,I689967,);
nor I_40427 (I689726,I689967,I689837);
nor I_40428 (I689717,I689967,I689893);
nand I_40429 (I690003,I576342,I576330);
and I_40430 (I690020,I690003,I576327);
DFFARX1 I_40431 (I690020,I2683,I689743,I690046,);
not I_40432 (I690054,I690046);
nand I_40433 (I690071,I690054,I689967);
nand I_40434 (I689720,I690054,I689876);
nor I_40435 (I690102,I576345,I576330);
and I_40436 (I690119,I689967,I690102);
nor I_40437 (I690136,I690054,I690119);
DFFARX1 I_40438 (I690136,I2683,I689743,I689729,);
nor I_40439 (I690167,I689769,I690102);
DFFARX1 I_40440 (I690167,I2683,I689743,I689714,);
nor I_40441 (I690198,I690046,I690102);
not I_40442 (I690215,I690198);
nand I_40443 (I689723,I690215,I690071);
not I_40444 (I690270,I2690);
DFFARX1 I_40445 (I422888,I2683,I690270,I690296,);
not I_40446 (I690304,I690296);
nand I_40447 (I690321,I422906,I422897);
and I_40448 (I690338,I690321,I422900);
DFFARX1 I_40449 (I690338,I2683,I690270,I690364,);
DFFARX1 I_40450 (I690364,I2683,I690270,I690259,);
DFFARX1 I_40451 (I422894,I2683,I690270,I690395,);
nand I_40452 (I690403,I690395,I422885);
not I_40453 (I690420,I690403);
DFFARX1 I_40454 (I690420,I2683,I690270,I690446,);
not I_40455 (I690454,I690446);
nor I_40456 (I690262,I690304,I690454);
DFFARX1 I_40457 (I422891,I2683,I690270,I690494,);
nor I_40458 (I690253,I690494,I690364);
nor I_40459 (I690244,I690494,I690420);
nand I_40460 (I690530,I422885,I422882);
and I_40461 (I690547,I690530,I422903);
DFFARX1 I_40462 (I690547,I2683,I690270,I690573,);
not I_40463 (I690581,I690573);
nand I_40464 (I690598,I690581,I690494);
nand I_40465 (I690247,I690581,I690403);
nor I_40466 (I690629,I422882,I422882);
and I_40467 (I690646,I690494,I690629);
nor I_40468 (I690663,I690581,I690646);
DFFARX1 I_40469 (I690663,I2683,I690270,I690256,);
nor I_40470 (I690694,I690296,I690629);
DFFARX1 I_40471 (I690694,I2683,I690270,I690241,);
nor I_40472 (I690725,I690573,I690629);
not I_40473 (I690742,I690725);
nand I_40474 (I690250,I690742,I690598);
not I_40475 (I690797,I2690);
DFFARX1 I_40476 (I1100109,I2683,I690797,I690823,);
not I_40477 (I690831,I690823);
nand I_40478 (I690848,I1100106,I1100115);
and I_40479 (I690865,I690848,I1100094);
DFFARX1 I_40480 (I690865,I2683,I690797,I690891,);
DFFARX1 I_40481 (I690891,I2683,I690797,I690786,);
DFFARX1 I_40482 (I1100097,I2683,I690797,I690922,);
nand I_40483 (I690930,I690922,I1100112);
not I_40484 (I690947,I690930);
DFFARX1 I_40485 (I690947,I2683,I690797,I690973,);
not I_40486 (I690981,I690973);
nor I_40487 (I690789,I690831,I690981);
DFFARX1 I_40488 (I1100118,I2683,I690797,I691021,);
nor I_40489 (I690780,I691021,I690891);
nor I_40490 (I690771,I691021,I690947);
nand I_40491 (I691057,I1100100,I1100121);
and I_40492 (I691074,I691057,I1100103);
DFFARX1 I_40493 (I691074,I2683,I690797,I691100,);
not I_40494 (I691108,I691100);
nand I_40495 (I691125,I691108,I691021);
nand I_40496 (I690774,I691108,I690930);
nor I_40497 (I691156,I1100094,I1100121);
and I_40498 (I691173,I691021,I691156);
nor I_40499 (I691190,I691108,I691173);
DFFARX1 I_40500 (I691190,I2683,I690797,I690783,);
nor I_40501 (I691221,I690823,I691156);
DFFARX1 I_40502 (I691221,I2683,I690797,I690768,);
nor I_40503 (I691252,I691100,I691156);
not I_40504 (I691269,I691252);
nand I_40505 (I690777,I691269,I691125);
not I_40506 (I691324,I2690);
DFFARX1 I_40507 (I405633,I2683,I691324,I691350,);
not I_40508 (I691358,I691350);
nand I_40509 (I691375,I405651,I405642);
and I_40510 (I691392,I691375,I405645);
DFFARX1 I_40511 (I691392,I2683,I691324,I691418,);
DFFARX1 I_40512 (I691418,I2683,I691324,I691313,);
DFFARX1 I_40513 (I405639,I2683,I691324,I691449,);
nand I_40514 (I691457,I691449,I405630);
not I_40515 (I691474,I691457);
DFFARX1 I_40516 (I691474,I2683,I691324,I691500,);
not I_40517 (I691508,I691500);
nor I_40518 (I691316,I691358,I691508);
DFFARX1 I_40519 (I405636,I2683,I691324,I691548,);
nor I_40520 (I691307,I691548,I691418);
nor I_40521 (I691298,I691548,I691474);
nand I_40522 (I691584,I405630,I405627);
and I_40523 (I691601,I691584,I405648);
DFFARX1 I_40524 (I691601,I2683,I691324,I691627,);
not I_40525 (I691635,I691627);
nand I_40526 (I691652,I691635,I691548);
nand I_40527 (I691301,I691635,I691457);
nor I_40528 (I691683,I405627,I405627);
and I_40529 (I691700,I691548,I691683);
nor I_40530 (I691717,I691635,I691700);
DFFARX1 I_40531 (I691717,I2683,I691324,I691310,);
nor I_40532 (I691748,I691350,I691683);
DFFARX1 I_40533 (I691748,I2683,I691324,I691295,);
nor I_40534 (I691779,I691627,I691683);
not I_40535 (I691796,I691779);
nand I_40536 (I691304,I691796,I691652);
not I_40537 (I691851,I2690);
DFFARX1 I_40538 (I220608,I2683,I691851,I691877,);
not I_40539 (I691885,I691877);
nand I_40540 (I691902,I220599,I220599);
and I_40541 (I691919,I691902,I220617);
DFFARX1 I_40542 (I691919,I2683,I691851,I691945,);
DFFARX1 I_40543 (I691945,I2683,I691851,I691840,);
DFFARX1 I_40544 (I220620,I2683,I691851,I691976,);
nand I_40545 (I691984,I691976,I220602);
not I_40546 (I692001,I691984);
DFFARX1 I_40547 (I692001,I2683,I691851,I692027,);
not I_40548 (I692035,I692027);
nor I_40549 (I691843,I691885,I692035);
DFFARX1 I_40550 (I220614,I2683,I691851,I692075,);
nor I_40551 (I691834,I692075,I691945);
nor I_40552 (I691825,I692075,I692001);
nand I_40553 (I692111,I220626,I220605);
and I_40554 (I692128,I692111,I220611);
DFFARX1 I_40555 (I692128,I2683,I691851,I692154,);
not I_40556 (I692162,I692154);
nand I_40557 (I692179,I692162,I692075);
nand I_40558 (I691828,I692162,I691984);
nor I_40559 (I692210,I220623,I220605);
and I_40560 (I692227,I692075,I692210);
nor I_40561 (I692244,I692162,I692227);
DFFARX1 I_40562 (I692244,I2683,I691851,I691837,);
nor I_40563 (I692275,I691877,I692210);
DFFARX1 I_40564 (I692275,I2683,I691851,I691822,);
nor I_40565 (I692306,I692154,I692210);
not I_40566 (I692323,I692306);
nand I_40567 (I691831,I692323,I692179);
not I_40568 (I692378,I2690);
DFFARX1 I_40569 (I519102,I2683,I692378,I692404,);
not I_40570 (I692412,I692404);
nand I_40571 (I692429,I519105,I519102);
and I_40572 (I692446,I692429,I519114);
DFFARX1 I_40573 (I692446,I2683,I692378,I692472,);
DFFARX1 I_40574 (I692472,I2683,I692378,I692367,);
DFFARX1 I_40575 (I519111,I2683,I692378,I692503,);
nand I_40576 (I692511,I692503,I519117);
not I_40577 (I692528,I692511);
DFFARX1 I_40578 (I692528,I2683,I692378,I692554,);
not I_40579 (I692562,I692554);
nor I_40580 (I692370,I692412,I692562);
DFFARX1 I_40581 (I519126,I2683,I692378,I692602,);
nor I_40582 (I692361,I692602,I692472);
nor I_40583 (I692352,I692602,I692528);
nand I_40584 (I692638,I519120,I519108);
and I_40585 (I692655,I692638,I519105);
DFFARX1 I_40586 (I692655,I2683,I692378,I692681,);
not I_40587 (I692689,I692681);
nand I_40588 (I692706,I692689,I692602);
nand I_40589 (I692355,I692689,I692511);
nor I_40590 (I692737,I519123,I519108);
and I_40591 (I692754,I692602,I692737);
nor I_40592 (I692771,I692689,I692754);
DFFARX1 I_40593 (I692771,I2683,I692378,I692364,);
nor I_40594 (I692802,I692404,I692737);
DFFARX1 I_40595 (I692802,I2683,I692378,I692349,);
nor I_40596 (I692833,I692681,I692737);
not I_40597 (I692850,I692833);
nand I_40598 (I692358,I692850,I692706);
not I_40599 (I692905,I2690);
DFFARX1 I_40600 (I1088209,I2683,I692905,I692931,);
not I_40601 (I692939,I692931);
nand I_40602 (I692956,I1088206,I1088215);
and I_40603 (I692973,I692956,I1088194);
DFFARX1 I_40604 (I692973,I2683,I692905,I692999,);
DFFARX1 I_40605 (I692999,I2683,I692905,I692894,);
DFFARX1 I_40606 (I1088197,I2683,I692905,I693030,);
nand I_40607 (I693038,I693030,I1088212);
not I_40608 (I693055,I693038);
DFFARX1 I_40609 (I693055,I2683,I692905,I693081,);
not I_40610 (I693089,I693081);
nor I_40611 (I692897,I692939,I693089);
DFFARX1 I_40612 (I1088218,I2683,I692905,I693129,);
nor I_40613 (I692888,I693129,I692999);
nor I_40614 (I692879,I693129,I693055);
nand I_40615 (I693165,I1088200,I1088221);
and I_40616 (I693182,I693165,I1088203);
DFFARX1 I_40617 (I693182,I2683,I692905,I693208,);
not I_40618 (I693216,I693208);
nand I_40619 (I693233,I693216,I693129);
nand I_40620 (I692882,I693216,I693038);
nor I_40621 (I693264,I1088194,I1088221);
and I_40622 (I693281,I693129,I693264);
nor I_40623 (I693298,I693216,I693281);
DFFARX1 I_40624 (I693298,I2683,I692905,I692891,);
nor I_40625 (I693329,I692931,I693264);
DFFARX1 I_40626 (I693329,I2683,I692905,I692876,);
nor I_40627 (I693360,I693208,I693264);
not I_40628 (I693377,I693360);
nand I_40629 (I692885,I693377,I693233);
not I_40630 (I693432,I2690);
DFFARX1 I_40631 (I717410,I2683,I693432,I693458,);
not I_40632 (I693466,I693458);
nand I_40633 (I693483,I717425,I717407);
and I_40634 (I693500,I693483,I717407);
DFFARX1 I_40635 (I693500,I2683,I693432,I693526,);
DFFARX1 I_40636 (I693526,I2683,I693432,I693421,);
DFFARX1 I_40637 (I717416,I2683,I693432,I693557,);
nand I_40638 (I693565,I693557,I717434);
not I_40639 (I693582,I693565);
DFFARX1 I_40640 (I693582,I2683,I693432,I693608,);
not I_40641 (I693616,I693608);
nor I_40642 (I693424,I693466,I693616);
DFFARX1 I_40643 (I717431,I2683,I693432,I693656,);
nor I_40644 (I693415,I693656,I693526);
nor I_40645 (I693406,I693656,I693582);
nand I_40646 (I693692,I717428,I717419);
and I_40647 (I693709,I693692,I717413);
DFFARX1 I_40648 (I693709,I2683,I693432,I693735,);
not I_40649 (I693743,I693735);
nand I_40650 (I693760,I693743,I693656);
nand I_40651 (I693409,I693743,I693565);
nor I_40652 (I693791,I717422,I717419);
and I_40653 (I693808,I693656,I693791);
nor I_40654 (I693825,I693743,I693808);
DFFARX1 I_40655 (I693825,I2683,I693432,I693418,);
nor I_40656 (I693856,I693458,I693791);
DFFARX1 I_40657 (I693856,I2683,I693432,I693403,);
nor I_40658 (I693887,I693735,I693791);
not I_40659 (I693904,I693887);
nand I_40660 (I693412,I693904,I693760);
not I_40661 (I693959,I2690);
DFFARX1 I_40662 (I879656,I2683,I693959,I693985,);
not I_40663 (I693993,I693985);
nand I_40664 (I694010,I879638,I879638);
and I_40665 (I694027,I694010,I879644);
DFFARX1 I_40666 (I694027,I2683,I693959,I694053,);
DFFARX1 I_40667 (I694053,I2683,I693959,I693948,);
DFFARX1 I_40668 (I879641,I2683,I693959,I694084,);
nand I_40669 (I694092,I694084,I879650);
not I_40670 (I694109,I694092);
DFFARX1 I_40671 (I694109,I2683,I693959,I694135,);
not I_40672 (I694143,I694135);
nor I_40673 (I693951,I693993,I694143);
DFFARX1 I_40674 (I879662,I2683,I693959,I694183,);
nor I_40675 (I693942,I694183,I694053);
nor I_40676 (I693933,I694183,I694109);
nand I_40677 (I694219,I879653,I879647);
and I_40678 (I694236,I694219,I879641);
DFFARX1 I_40679 (I694236,I2683,I693959,I694262,);
not I_40680 (I694270,I694262);
nand I_40681 (I694287,I694270,I694183);
nand I_40682 (I693936,I694270,I694092);
nor I_40683 (I694318,I879659,I879647);
and I_40684 (I694335,I694183,I694318);
nor I_40685 (I694352,I694270,I694335);
DFFARX1 I_40686 (I694352,I2683,I693959,I693945,);
nor I_40687 (I694383,I693985,I694318);
DFFARX1 I_40688 (I694383,I2683,I693959,I693930,);
nor I_40689 (I694414,I694262,I694318);
not I_40690 (I694431,I694414);
nand I_40691 (I693939,I694431,I694287);
not I_40692 (I694486,I2690);
DFFARX1 I_40693 (I66977,I2683,I694486,I694512,);
not I_40694 (I694520,I694512);
nand I_40695 (I694537,I66953,I66962);
and I_40696 (I694554,I694537,I66956);
DFFARX1 I_40697 (I694554,I2683,I694486,I694580,);
DFFARX1 I_40698 (I694580,I2683,I694486,I694475,);
DFFARX1 I_40699 (I66974,I2683,I694486,I694611,);
nand I_40700 (I694619,I694611,I66965);
not I_40701 (I694636,I694619);
DFFARX1 I_40702 (I694636,I2683,I694486,I694662,);
not I_40703 (I694670,I694662);
nor I_40704 (I694478,I694520,I694670);
DFFARX1 I_40705 (I66959,I2683,I694486,I694710,);
nor I_40706 (I694469,I694710,I694580);
nor I_40707 (I694460,I694710,I694636);
nand I_40708 (I694746,I66971,I66968);
and I_40709 (I694763,I694746,I66956);
DFFARX1 I_40710 (I694763,I2683,I694486,I694789,);
not I_40711 (I694797,I694789);
nand I_40712 (I694814,I694797,I694710);
nand I_40713 (I694463,I694797,I694619);
nor I_40714 (I694845,I66953,I66968);
and I_40715 (I694862,I694710,I694845);
nor I_40716 (I694879,I694797,I694862);
DFFARX1 I_40717 (I694879,I2683,I694486,I694472,);
nor I_40718 (I694910,I694512,I694845);
DFFARX1 I_40719 (I694910,I2683,I694486,I694457,);
nor I_40720 (I694941,I694789,I694845);
not I_40721 (I694958,I694941);
nand I_40722 (I694466,I694958,I694814);
not I_40723 (I695013,I2690);
DFFARX1 I_40724 (I850178,I2683,I695013,I695039,);
not I_40725 (I695047,I695039);
nand I_40726 (I695064,I850160,I850160);
and I_40727 (I695081,I695064,I850166);
DFFARX1 I_40728 (I695081,I2683,I695013,I695107,);
DFFARX1 I_40729 (I695107,I2683,I695013,I695002,);
DFFARX1 I_40730 (I850163,I2683,I695013,I695138,);
nand I_40731 (I695146,I695138,I850172);
not I_40732 (I695163,I695146);
DFFARX1 I_40733 (I695163,I2683,I695013,I695189,);
not I_40734 (I695197,I695189);
nor I_40735 (I695005,I695047,I695197);
DFFARX1 I_40736 (I850184,I2683,I695013,I695237,);
nor I_40737 (I694996,I695237,I695107);
nor I_40738 (I694987,I695237,I695163);
nand I_40739 (I695273,I850175,I850169);
and I_40740 (I695290,I695273,I850163);
DFFARX1 I_40741 (I695290,I2683,I695013,I695316,);
not I_40742 (I695324,I695316);
nand I_40743 (I695341,I695324,I695237);
nand I_40744 (I694990,I695324,I695146);
nor I_40745 (I695372,I850181,I850169);
and I_40746 (I695389,I695237,I695372);
nor I_40747 (I695406,I695324,I695389);
DFFARX1 I_40748 (I695406,I2683,I695013,I694999,);
nor I_40749 (I695437,I695039,I695372);
DFFARX1 I_40750 (I695437,I2683,I695013,I694984,);
nor I_40751 (I695468,I695316,I695372);
not I_40752 (I695485,I695468);
nand I_40753 (I694993,I695485,I695341);
not I_40754 (I695540,I2690);
DFFARX1 I_40755 (I20059,I2683,I695540,I695566,);
not I_40756 (I695574,I695566);
nand I_40757 (I695591,I20071,I20074);
and I_40758 (I695608,I695591,I20050);
DFFARX1 I_40759 (I695608,I2683,I695540,I695634,);
DFFARX1 I_40760 (I695634,I2683,I695540,I695529,);
DFFARX1 I_40761 (I20068,I2683,I695540,I695665,);
nand I_40762 (I695673,I695665,I20056);
not I_40763 (I695690,I695673);
DFFARX1 I_40764 (I695690,I2683,I695540,I695716,);
not I_40765 (I695724,I695716);
nor I_40766 (I695532,I695574,I695724);
DFFARX1 I_40767 (I20053,I2683,I695540,I695764,);
nor I_40768 (I695523,I695764,I695634);
nor I_40769 (I695514,I695764,I695690);
nand I_40770 (I695800,I20062,I20053);
and I_40771 (I695817,I695800,I20050);
DFFARX1 I_40772 (I695817,I2683,I695540,I695843,);
not I_40773 (I695851,I695843);
nand I_40774 (I695868,I695851,I695764);
nand I_40775 (I695517,I695851,I695673);
nor I_40776 (I695899,I20065,I20053);
and I_40777 (I695916,I695764,I695899);
nor I_40778 (I695933,I695851,I695916);
DFFARX1 I_40779 (I695933,I2683,I695540,I695526,);
nor I_40780 (I695964,I695566,I695899);
DFFARX1 I_40781 (I695964,I2683,I695540,I695511,);
nor I_40782 (I695995,I695843,I695899);
not I_40783 (I696012,I695995);
nand I_40784 (I695520,I696012,I695868);
not I_40785 (I696067,I2690);
DFFARX1 I_40786 (I835150,I2683,I696067,I696093,);
not I_40787 (I696101,I696093);
nand I_40788 (I696118,I835132,I835132);
and I_40789 (I696135,I696118,I835138);
DFFARX1 I_40790 (I696135,I2683,I696067,I696161,);
DFFARX1 I_40791 (I696161,I2683,I696067,I696056,);
DFFARX1 I_40792 (I835135,I2683,I696067,I696192,);
nand I_40793 (I696200,I696192,I835144);
not I_40794 (I696217,I696200);
DFFARX1 I_40795 (I696217,I2683,I696067,I696243,);
not I_40796 (I696251,I696243);
nor I_40797 (I696059,I696101,I696251);
DFFARX1 I_40798 (I835156,I2683,I696067,I696291,);
nor I_40799 (I696050,I696291,I696161);
nor I_40800 (I696041,I696291,I696217);
nand I_40801 (I696327,I835147,I835141);
and I_40802 (I696344,I696327,I835135);
DFFARX1 I_40803 (I696344,I2683,I696067,I696370,);
not I_40804 (I696378,I696370);
nand I_40805 (I696395,I696378,I696291);
nand I_40806 (I696044,I696378,I696200);
nor I_40807 (I696426,I835153,I835141);
and I_40808 (I696443,I696291,I696426);
nor I_40809 (I696460,I696378,I696443);
DFFARX1 I_40810 (I696460,I2683,I696067,I696053,);
nor I_40811 (I696491,I696093,I696426);
DFFARX1 I_40812 (I696491,I2683,I696067,I696038,);
nor I_40813 (I696522,I696370,I696426);
not I_40814 (I696539,I696522);
nand I_40815 (I696047,I696539,I696395);
not I_40816 (I696594,I2690);
DFFARX1 I_40817 (I612160,I2683,I696594,I696620,);
not I_40818 (I696628,I696620);
nand I_40819 (I696645,I612163,I612160);
and I_40820 (I696662,I696645,I612172);
DFFARX1 I_40821 (I696662,I2683,I696594,I696688,);
DFFARX1 I_40822 (I696688,I2683,I696594,I696583,);
DFFARX1 I_40823 (I612169,I2683,I696594,I696719,);
nand I_40824 (I696727,I696719,I612175);
not I_40825 (I696744,I696727);
DFFARX1 I_40826 (I696744,I2683,I696594,I696770,);
not I_40827 (I696778,I696770);
nor I_40828 (I696586,I696628,I696778);
DFFARX1 I_40829 (I612184,I2683,I696594,I696818,);
nor I_40830 (I696577,I696818,I696688);
nor I_40831 (I696568,I696818,I696744);
nand I_40832 (I696854,I612178,I612166);
and I_40833 (I696871,I696854,I612163);
DFFARX1 I_40834 (I696871,I2683,I696594,I696897,);
not I_40835 (I696905,I696897);
nand I_40836 (I696922,I696905,I696818);
nand I_40837 (I696571,I696905,I696727);
nor I_40838 (I696953,I612181,I612166);
and I_40839 (I696970,I696818,I696953);
nor I_40840 (I696987,I696905,I696970);
DFFARX1 I_40841 (I696987,I2683,I696594,I696580,);
nor I_40842 (I697018,I696620,I696953);
DFFARX1 I_40843 (I697018,I2683,I696594,I696565,);
nor I_40844 (I697049,I696897,I696953);
not I_40845 (I697066,I697049);
nand I_40846 (I696574,I697066,I696922);
not I_40847 (I697121,I2690);
DFFARX1 I_40848 (I789116,I2683,I697121,I697147,);
not I_40849 (I697155,I697147);
nand I_40850 (I697172,I789131,I789113);
and I_40851 (I697189,I697172,I789113);
DFFARX1 I_40852 (I697189,I2683,I697121,I697215,);
DFFARX1 I_40853 (I697215,I2683,I697121,I697110,);
DFFARX1 I_40854 (I789122,I2683,I697121,I697246,);
nand I_40855 (I697254,I697246,I789140);
not I_40856 (I697271,I697254);
DFFARX1 I_40857 (I697271,I2683,I697121,I697297,);
not I_40858 (I697305,I697297);
nor I_40859 (I697113,I697155,I697305);
DFFARX1 I_40860 (I789137,I2683,I697121,I697345,);
nor I_40861 (I697104,I697345,I697215);
nor I_40862 (I697095,I697345,I697271);
nand I_40863 (I697381,I789134,I789125);
and I_40864 (I697398,I697381,I789119);
DFFARX1 I_40865 (I697398,I2683,I697121,I697424,);
not I_40866 (I697432,I697424);
nand I_40867 (I697449,I697432,I697345);
nand I_40868 (I697098,I697432,I697254);
nor I_40869 (I697480,I789128,I789125);
and I_40870 (I697497,I697345,I697480);
nor I_40871 (I697514,I697432,I697497);
DFFARX1 I_40872 (I697514,I2683,I697121,I697107,);
nor I_40873 (I697545,I697147,I697480);
DFFARX1 I_40874 (I697545,I2683,I697121,I697092,);
nor I_40875 (I697576,I697424,I697480);
not I_40876 (I697593,I697576);
nand I_40877 (I697101,I697593,I697449);
not I_40878 (I697648,I2690);
DFFARX1 I_40879 (I422293,I2683,I697648,I697674,);
not I_40880 (I697682,I697674);
nand I_40881 (I697699,I422311,I422302);
and I_40882 (I697716,I697699,I422305);
DFFARX1 I_40883 (I697716,I2683,I697648,I697742,);
DFFARX1 I_40884 (I697742,I2683,I697648,I697637,);
DFFARX1 I_40885 (I422299,I2683,I697648,I697773,);
nand I_40886 (I697781,I697773,I422290);
not I_40887 (I697798,I697781);
DFFARX1 I_40888 (I697798,I2683,I697648,I697824,);
not I_40889 (I697832,I697824);
nor I_40890 (I697640,I697682,I697832);
DFFARX1 I_40891 (I422296,I2683,I697648,I697872,);
nor I_40892 (I697631,I697872,I697742);
nor I_40893 (I697622,I697872,I697798);
nand I_40894 (I697908,I422290,I422287);
and I_40895 (I697925,I697908,I422308);
DFFARX1 I_40896 (I697925,I2683,I697648,I697951,);
not I_40897 (I697959,I697951);
nand I_40898 (I697976,I697959,I697872);
nand I_40899 (I697625,I697959,I697781);
nor I_40900 (I698007,I422287,I422287);
and I_40901 (I698024,I697872,I698007);
nor I_40902 (I698041,I697959,I698024);
DFFARX1 I_40903 (I698041,I2683,I697648,I697634,);
nor I_40904 (I698072,I697674,I698007);
DFFARX1 I_40905 (I698072,I2683,I697648,I697619,);
nor I_40906 (I698103,I697951,I698007);
not I_40907 (I698120,I698103);
nand I_40908 (I697628,I698120,I697976);
not I_40909 (I698175,I2690);
DFFARX1 I_40910 (I764568,I2683,I698175,I698201,);
not I_40911 (I698209,I698201);
nand I_40912 (I698226,I764583,I764565);
and I_40913 (I698243,I698226,I764565);
DFFARX1 I_40914 (I698243,I2683,I698175,I698269,);
DFFARX1 I_40915 (I698269,I2683,I698175,I698164,);
DFFARX1 I_40916 (I764574,I2683,I698175,I698300,);
nand I_40917 (I698308,I698300,I764592);
not I_40918 (I698325,I698308);
DFFARX1 I_40919 (I698325,I2683,I698175,I698351,);
not I_40920 (I698359,I698351);
nor I_40921 (I698167,I698209,I698359);
DFFARX1 I_40922 (I764589,I2683,I698175,I698399,);
nor I_40923 (I698158,I698399,I698269);
nor I_40924 (I698149,I698399,I698325);
nand I_40925 (I698435,I764586,I764577);
and I_40926 (I698452,I698435,I764571);
DFFARX1 I_40927 (I698452,I2683,I698175,I698478,);
not I_40928 (I698486,I698478);
nand I_40929 (I698503,I698486,I698399);
nand I_40930 (I698152,I698486,I698308);
nor I_40931 (I698534,I764580,I764577);
and I_40932 (I698551,I698399,I698534);
nor I_40933 (I698568,I698486,I698551);
DFFARX1 I_40934 (I698568,I2683,I698175,I698161,);
nor I_40935 (I698599,I698201,I698534);
DFFARX1 I_40936 (I698599,I2683,I698175,I698146,);
nor I_40937 (I698630,I698478,I698534);
not I_40938 (I698647,I698630);
nand I_40939 (I698155,I698647,I698503);
not I_40940 (I698708,I2690);
DFFARX1 I_40941 (I333944,I2683,I698708,I698734,);
DFFARX1 I_40942 (I333941,I2683,I698708,I698751,);
not I_40943 (I698759,I698751);
not I_40944 (I698776,I333956);
nor I_40945 (I698793,I698776,I333959);
not I_40946 (I698810,I333947);
nor I_40947 (I698827,I698793,I333953);
nor I_40948 (I698844,I698751,I698827);
DFFARX1 I_40949 (I698844,I2683,I698708,I698694,);
nor I_40950 (I698875,I333953,I333959);
nand I_40951 (I698892,I698875,I333956);
DFFARX1 I_40952 (I698892,I2683,I698708,I698697,);
nor I_40953 (I698923,I698810,I333953);
nand I_40954 (I698940,I698923,I333965);
nor I_40955 (I698957,I698734,I698940);
DFFARX1 I_40956 (I698957,I2683,I698708,I698673,);
not I_40957 (I698988,I698940);
nand I_40958 (I698685,I698751,I698988);
DFFARX1 I_40959 (I698940,I2683,I698708,I699028,);
not I_40960 (I699036,I699028);
not I_40961 (I699053,I333953);
not I_40962 (I699070,I333938);
nor I_40963 (I699087,I699070,I333947);
nor I_40964 (I698700,I699036,I699087);
nor I_40965 (I699118,I699070,I333950);
and I_40966 (I699135,I699118,I333938);
or I_40967 (I699152,I699135,I333962);
DFFARX1 I_40968 (I699152,I2683,I698708,I699178,);
nor I_40969 (I698688,I699178,I698734);
not I_40970 (I699200,I699178);
and I_40971 (I699217,I699200,I698734);
nor I_40972 (I698682,I698759,I699217);
nand I_40973 (I699248,I699200,I698810);
nor I_40974 (I698676,I699070,I699248);
nand I_40975 (I698679,I699200,I698988);
nand I_40976 (I699293,I698810,I333938);
nor I_40977 (I698691,I699053,I699293);
not I_40978 (I699354,I2690);
DFFARX1 I_40979 (I252746,I2683,I699354,I699380,);
DFFARX1 I_40980 (I252752,I2683,I699354,I699397,);
not I_40981 (I699405,I699397);
not I_40982 (I699422,I252773);
nor I_40983 (I699439,I699422,I252761);
not I_40984 (I699456,I252770);
nor I_40985 (I699473,I699439,I252755);
nor I_40986 (I699490,I699397,I699473);
DFFARX1 I_40987 (I699490,I2683,I699354,I699340,);
nor I_40988 (I699521,I252755,I252761);
nand I_40989 (I699538,I699521,I252773);
DFFARX1 I_40990 (I699538,I2683,I699354,I699343,);
nor I_40991 (I699569,I699456,I252755);
nand I_40992 (I699586,I699569,I252746);
nor I_40993 (I699603,I699380,I699586);
DFFARX1 I_40994 (I699603,I2683,I699354,I699319,);
not I_40995 (I699634,I699586);
nand I_40996 (I699331,I699397,I699634);
DFFARX1 I_40997 (I699586,I2683,I699354,I699674,);
not I_40998 (I699682,I699674);
not I_40999 (I699699,I252755);
not I_41000 (I699716,I252758);
nor I_41001 (I699733,I699716,I252770);
nor I_41002 (I699346,I699682,I699733);
nor I_41003 (I699764,I699716,I252767);
and I_41004 (I699781,I699764,I252749);
or I_41005 (I699798,I699781,I252764);
DFFARX1 I_41006 (I699798,I2683,I699354,I699824,);
nor I_41007 (I699334,I699824,I699380);
not I_41008 (I699846,I699824);
and I_41009 (I699863,I699846,I699380);
nor I_41010 (I699328,I699405,I699863);
nand I_41011 (I699894,I699846,I699456);
nor I_41012 (I699322,I699716,I699894);
nand I_41013 (I699325,I699846,I699634);
nand I_41014 (I699939,I699456,I252758);
nor I_41015 (I699337,I699699,I699939);
not I_41016 (I700000,I2690);
DFFARX1 I_41017 (I606964,I2683,I700000,I700026,);
DFFARX1 I_41018 (I606958,I2683,I700000,I700043,);
not I_41019 (I700051,I700043);
not I_41020 (I700068,I606973);
nor I_41021 (I700085,I700068,I606958);
not I_41022 (I700102,I606967);
nor I_41023 (I700119,I700085,I606976);
nor I_41024 (I700136,I700043,I700119);
DFFARX1 I_41025 (I700136,I2683,I700000,I699986,);
nor I_41026 (I700167,I606976,I606958);
nand I_41027 (I700184,I700167,I606973);
DFFARX1 I_41028 (I700184,I2683,I700000,I699989,);
nor I_41029 (I700215,I700102,I606976);
nand I_41030 (I700232,I700215,I606961);
nor I_41031 (I700249,I700026,I700232);
DFFARX1 I_41032 (I700249,I2683,I700000,I699965,);
not I_41033 (I700280,I700232);
nand I_41034 (I699977,I700043,I700280);
DFFARX1 I_41035 (I700232,I2683,I700000,I700320,);
not I_41036 (I700328,I700320);
not I_41037 (I700345,I606976);
not I_41038 (I700362,I606970);
nor I_41039 (I700379,I700362,I606967);
nor I_41040 (I699992,I700328,I700379);
nor I_41041 (I700410,I700362,I606979);
and I_41042 (I700427,I700410,I606982);
or I_41043 (I700444,I700427,I606961);
DFFARX1 I_41044 (I700444,I2683,I700000,I700470,);
nor I_41045 (I699980,I700470,I700026);
not I_41046 (I700492,I700470);
and I_41047 (I700509,I700492,I700026);
nor I_41048 (I699974,I700051,I700509);
nand I_41049 (I700540,I700492,I700102);
nor I_41050 (I699968,I700362,I700540);
nand I_41051 (I699971,I700492,I700280);
nand I_41052 (I700585,I700102,I606970);
nor I_41053 (I699983,I700345,I700585);
not I_41054 (I700646,I2690);
DFFARX1 I_41055 (I681288,I2683,I700646,I700672,);
DFFARX1 I_41056 (I681285,I2683,I700646,I700689,);
not I_41057 (I700697,I700689);
not I_41058 (I700714,I681285);
nor I_41059 (I700731,I700714,I681288);
not I_41060 (I700748,I681300);
nor I_41061 (I700765,I700731,I681294);
nor I_41062 (I700782,I700689,I700765);
DFFARX1 I_41063 (I700782,I2683,I700646,I700632,);
nor I_41064 (I700813,I681294,I681288);
nand I_41065 (I700830,I700813,I681285);
DFFARX1 I_41066 (I700830,I2683,I700646,I700635,);
nor I_41067 (I700861,I700748,I681294);
nand I_41068 (I700878,I700861,I681282);
nor I_41069 (I700895,I700672,I700878);
DFFARX1 I_41070 (I700895,I2683,I700646,I700611,);
not I_41071 (I700926,I700878);
nand I_41072 (I700623,I700689,I700926);
DFFARX1 I_41073 (I700878,I2683,I700646,I700966,);
not I_41074 (I700974,I700966);
not I_41075 (I700991,I681294);
not I_41076 (I701008,I681291);
nor I_41077 (I701025,I701008,I681300);
nor I_41078 (I700638,I700974,I701025);
nor I_41079 (I701056,I701008,I681297);
and I_41080 (I701073,I701056,I681303);
or I_41081 (I701090,I701073,I681282);
DFFARX1 I_41082 (I701090,I2683,I700646,I701116,);
nor I_41083 (I700626,I701116,I700672);
not I_41084 (I701138,I701116);
and I_41085 (I701155,I701138,I700672);
nor I_41086 (I700620,I700697,I701155);
nand I_41087 (I701186,I701138,I700748);
nor I_41088 (I700614,I701008,I701186);
nand I_41089 (I700617,I701138,I700926);
nand I_41090 (I701231,I700748,I681291);
nor I_41091 (I700629,I700991,I701231);
not I_41092 (I701292,I2690);
DFFARX1 I_41093 (I223234,I2683,I701292,I701318,);
DFFARX1 I_41094 (I223240,I2683,I701292,I701335,);
not I_41095 (I701343,I701335);
not I_41096 (I701360,I223261);
nor I_41097 (I701377,I701360,I223249);
not I_41098 (I701394,I223258);
nor I_41099 (I701411,I701377,I223243);
nor I_41100 (I701428,I701335,I701411);
DFFARX1 I_41101 (I701428,I2683,I701292,I701278,);
nor I_41102 (I701459,I223243,I223249);
nand I_41103 (I701476,I701459,I223261);
DFFARX1 I_41104 (I701476,I2683,I701292,I701281,);
nor I_41105 (I701507,I701394,I223243);
nand I_41106 (I701524,I701507,I223234);
nor I_41107 (I701541,I701318,I701524);
DFFARX1 I_41108 (I701541,I2683,I701292,I701257,);
not I_41109 (I701572,I701524);
nand I_41110 (I701269,I701335,I701572);
DFFARX1 I_41111 (I701524,I2683,I701292,I701612,);
not I_41112 (I701620,I701612);
not I_41113 (I701637,I223243);
not I_41114 (I701654,I223246);
nor I_41115 (I701671,I701654,I223258);
nor I_41116 (I701284,I701620,I701671);
nor I_41117 (I701702,I701654,I223255);
and I_41118 (I701719,I701702,I223237);
or I_41119 (I701736,I701719,I223252);
DFFARX1 I_41120 (I701736,I2683,I701292,I701762,);
nor I_41121 (I701272,I701762,I701318);
not I_41122 (I701784,I701762);
and I_41123 (I701801,I701784,I701318);
nor I_41124 (I701266,I701343,I701801);
nand I_41125 (I701832,I701784,I701394);
nor I_41126 (I701260,I701654,I701832);
nand I_41127 (I701263,I701784,I701572);
nand I_41128 (I701877,I701394,I223246);
nor I_41129 (I701275,I701637,I701877);
not I_41130 (I701938,I2690);
DFFARX1 I_41131 (I939768,I2683,I701938,I701964,);
DFFARX1 I_41132 (I939750,I2683,I701938,I701981,);
not I_41133 (I701989,I701981);
not I_41134 (I702006,I939759);
nor I_41135 (I702023,I702006,I939771);
not I_41136 (I702040,I939753);
nor I_41137 (I702057,I702023,I939762);
nor I_41138 (I702074,I701981,I702057);
DFFARX1 I_41139 (I702074,I2683,I701938,I701924,);
nor I_41140 (I702105,I939762,I939771);
nand I_41141 (I702122,I702105,I939759);
DFFARX1 I_41142 (I702122,I2683,I701938,I701927,);
nor I_41143 (I702153,I702040,I939762);
nand I_41144 (I702170,I702153,I939774);
nor I_41145 (I702187,I701964,I702170);
DFFARX1 I_41146 (I702187,I2683,I701938,I701903,);
not I_41147 (I702218,I702170);
nand I_41148 (I701915,I701981,I702218);
DFFARX1 I_41149 (I702170,I2683,I701938,I702258,);
not I_41150 (I702266,I702258);
not I_41151 (I702283,I939762);
not I_41152 (I702300,I939750);
nor I_41153 (I702317,I702300,I939753);
nor I_41154 (I701930,I702266,I702317);
nor I_41155 (I702348,I702300,I939756);
and I_41156 (I702365,I702348,I939765);
or I_41157 (I702382,I702365,I939753);
DFFARX1 I_41158 (I702382,I2683,I701938,I702408,);
nor I_41159 (I701918,I702408,I701964);
not I_41160 (I702430,I702408);
and I_41161 (I702447,I702430,I701964);
nor I_41162 (I701912,I701989,I702447);
nand I_41163 (I702478,I702430,I702040);
nor I_41164 (I701906,I702300,I702478);
nand I_41165 (I701909,I702430,I702218);
nand I_41166 (I702523,I702040,I939750);
nor I_41167 (I701921,I702283,I702523);
not I_41168 (I702584,I2690);
DFFARX1 I_41169 (I201531,I2683,I702584,I702610,);
DFFARX1 I_41170 (I201543,I2683,I702584,I702627,);
not I_41171 (I702635,I702627);
not I_41172 (I702652,I201549);
nor I_41173 (I702669,I702652,I201534);
not I_41174 (I702686,I201525);
nor I_41175 (I702703,I702669,I201546);
nor I_41176 (I702720,I702627,I702703);
DFFARX1 I_41177 (I702720,I2683,I702584,I702570,);
nor I_41178 (I702751,I201546,I201534);
nand I_41179 (I702768,I702751,I201549);
DFFARX1 I_41180 (I702768,I2683,I702584,I702573,);
nor I_41181 (I702799,I702686,I201546);
nand I_41182 (I702816,I702799,I201528);
nor I_41183 (I702833,I702610,I702816);
DFFARX1 I_41184 (I702833,I2683,I702584,I702549,);
not I_41185 (I702864,I702816);
nand I_41186 (I702561,I702627,I702864);
DFFARX1 I_41187 (I702816,I2683,I702584,I702904,);
not I_41188 (I702912,I702904);
not I_41189 (I702929,I201546);
not I_41190 (I702946,I201537);
nor I_41191 (I702963,I702946,I201525);
nor I_41192 (I702576,I702912,I702963);
nor I_41193 (I702994,I702946,I201540);
and I_41194 (I703011,I702994,I201528);
or I_41195 (I703028,I703011,I201525);
DFFARX1 I_41196 (I703028,I2683,I702584,I703054,);
nor I_41197 (I702564,I703054,I702610);
not I_41198 (I703076,I703054);
and I_41199 (I703093,I703076,I702610);
nor I_41200 (I702558,I702635,I703093);
nand I_41201 (I703124,I703076,I702686);
nor I_41202 (I702552,I702946,I703124);
nand I_41203 (I702555,I703076,I702864);
nand I_41204 (I703169,I702686,I201537);
nor I_41205 (I702567,I702929,I703169);
not I_41206 (I703230,I2690);
DFFARX1 I_41207 (I314405,I2683,I703230,I703256,);
DFFARX1 I_41208 (I314411,I2683,I703230,I703273,);
not I_41209 (I703281,I703273);
not I_41210 (I703298,I314432);
nor I_41211 (I703315,I703298,I314420);
not I_41212 (I703332,I314429);
nor I_41213 (I703349,I703315,I314414);
nor I_41214 (I703366,I703273,I703349);
DFFARX1 I_41215 (I703366,I2683,I703230,I703216,);
nor I_41216 (I703397,I314414,I314420);
nand I_41217 (I703414,I703397,I314432);
DFFARX1 I_41218 (I703414,I2683,I703230,I703219,);
nor I_41219 (I703445,I703332,I314414);
nand I_41220 (I703462,I703445,I314405);
nor I_41221 (I703479,I703256,I703462);
DFFARX1 I_41222 (I703479,I2683,I703230,I703195,);
not I_41223 (I703510,I703462);
nand I_41224 (I703207,I703273,I703510);
DFFARX1 I_41225 (I703462,I2683,I703230,I703550,);
not I_41226 (I703558,I703550);
not I_41227 (I703575,I314414);
not I_41228 (I703592,I314417);
nor I_41229 (I703609,I703592,I314429);
nor I_41230 (I703222,I703558,I703609);
nor I_41231 (I703640,I703592,I314426);
and I_41232 (I703657,I703640,I314408);
or I_41233 (I703674,I703657,I314423);
DFFARX1 I_41234 (I703674,I2683,I703230,I703700,);
nor I_41235 (I703210,I703700,I703256);
not I_41236 (I703722,I703700);
and I_41237 (I703739,I703722,I703256);
nor I_41238 (I703204,I703281,I703739);
nand I_41239 (I703770,I703722,I703332);
nor I_41240 (I703198,I703592,I703770);
nand I_41241 (I703201,I703722,I703510);
nand I_41242 (I703815,I703332,I314417);
nor I_41243 (I703213,I703575,I703815);
not I_41244 (I703876,I2690);
DFFARX1 I_41245 (I866362,I2683,I703876,I703902,);
DFFARX1 I_41246 (I866344,I2683,I703876,I703919,);
not I_41247 (I703927,I703919);
not I_41248 (I703944,I866353);
nor I_41249 (I703961,I703944,I866365);
not I_41250 (I703978,I866347);
nor I_41251 (I703995,I703961,I866356);
nor I_41252 (I704012,I703919,I703995);
DFFARX1 I_41253 (I704012,I2683,I703876,I703862,);
nor I_41254 (I704043,I866356,I866365);
nand I_41255 (I704060,I704043,I866353);
DFFARX1 I_41256 (I704060,I2683,I703876,I703865,);
nor I_41257 (I704091,I703978,I866356);
nand I_41258 (I704108,I704091,I866368);
nor I_41259 (I704125,I703902,I704108);
DFFARX1 I_41260 (I704125,I2683,I703876,I703841,);
not I_41261 (I704156,I704108);
nand I_41262 (I703853,I703919,I704156);
DFFARX1 I_41263 (I704108,I2683,I703876,I704196,);
not I_41264 (I704204,I704196);
not I_41265 (I704221,I866356);
not I_41266 (I704238,I866344);
nor I_41267 (I704255,I704238,I866347);
nor I_41268 (I703868,I704204,I704255);
nor I_41269 (I704286,I704238,I866350);
and I_41270 (I704303,I704286,I866359);
or I_41271 (I704320,I704303,I866347);
DFFARX1 I_41272 (I704320,I2683,I703876,I704346,);
nor I_41273 (I703856,I704346,I703902);
not I_41274 (I704368,I704346);
and I_41275 (I704385,I704368,I703902);
nor I_41276 (I703850,I703927,I704385);
nand I_41277 (I704416,I704368,I703978);
nor I_41278 (I703844,I704238,I704416);
nand I_41279 (I703847,I704368,I704156);
nand I_41280 (I704461,I703978,I866344);
nor I_41281 (I703859,I704221,I704461);
not I_41282 (I704522,I2690);
DFFARX1 I_41283 (I9836,I2683,I704522,I704548,);
DFFARX1 I_41284 (I9833,I2683,I704522,I704565,);
not I_41285 (I704573,I704565);
not I_41286 (I704590,I9845);
nor I_41287 (I704607,I704590,I9842);
not I_41288 (I704624,I9851);
nor I_41289 (I704641,I704607,I9848);
nor I_41290 (I704658,I704565,I704641);
DFFARX1 I_41291 (I704658,I2683,I704522,I704508,);
nor I_41292 (I704689,I9848,I9842);
nand I_41293 (I704706,I704689,I9845);
DFFARX1 I_41294 (I704706,I2683,I704522,I704511,);
nor I_41295 (I704737,I704624,I9848);
nand I_41296 (I704754,I704737,I9839);
nor I_41297 (I704771,I704548,I704754);
DFFARX1 I_41298 (I704771,I2683,I704522,I704487,);
not I_41299 (I704802,I704754);
nand I_41300 (I704499,I704565,I704802);
DFFARX1 I_41301 (I704754,I2683,I704522,I704842,);
not I_41302 (I704850,I704842);
not I_41303 (I704867,I9848);
not I_41304 (I704884,I9839);
nor I_41305 (I704901,I704884,I9851);
nor I_41306 (I704514,I704850,I704901);
nor I_41307 (I704932,I704884,I9833);
and I_41308 (I704949,I704932,I9854);
or I_41309 (I704966,I704949,I9836);
DFFARX1 I_41310 (I704966,I2683,I704522,I704992,);
nor I_41311 (I704502,I704992,I704548);
not I_41312 (I705014,I704992);
and I_41313 (I705031,I705014,I704548);
nor I_41314 (I704496,I704573,I705031);
nand I_41315 (I705062,I705014,I704624);
nor I_41316 (I704490,I704884,I705062);
nand I_41317 (I704493,I705014,I704802);
nand I_41318 (I705107,I704624,I9839);
nor I_41319 (I704505,I704867,I705107);
not I_41320 (I705168,I2690);
DFFARX1 I_41321 (I357880,I2683,I705168,I705194,);
DFFARX1 I_41322 (I357877,I2683,I705168,I705211,);
not I_41323 (I705219,I705211);
not I_41324 (I705236,I357892);
nor I_41325 (I705253,I705236,I357895);
not I_41326 (I705270,I357883);
nor I_41327 (I705287,I705253,I357889);
nor I_41328 (I705304,I705211,I705287);
DFFARX1 I_41329 (I705304,I2683,I705168,I705154,);
nor I_41330 (I705335,I357889,I357895);
nand I_41331 (I705352,I705335,I357892);
DFFARX1 I_41332 (I705352,I2683,I705168,I705157,);
nor I_41333 (I705383,I705270,I357889);
nand I_41334 (I705400,I705383,I357901);
nor I_41335 (I705417,I705194,I705400);
DFFARX1 I_41336 (I705417,I2683,I705168,I705133,);
not I_41337 (I705448,I705400);
nand I_41338 (I705145,I705211,I705448);
DFFARX1 I_41339 (I705400,I2683,I705168,I705488,);
not I_41340 (I705496,I705488);
not I_41341 (I705513,I357889);
not I_41342 (I705530,I357874);
nor I_41343 (I705547,I705530,I357883);
nor I_41344 (I705160,I705496,I705547);
nor I_41345 (I705578,I705530,I357886);
and I_41346 (I705595,I705578,I357874);
or I_41347 (I705612,I705595,I357898);
DFFARX1 I_41348 (I705612,I2683,I705168,I705638,);
nor I_41349 (I705148,I705638,I705194);
not I_41350 (I705660,I705638);
and I_41351 (I705677,I705660,I705194);
nor I_41352 (I705142,I705219,I705677);
nand I_41353 (I705708,I705660,I705270);
nor I_41354 (I705136,I705530,I705708);
nand I_41355 (I705139,I705660,I705448);
nand I_41356 (I705753,I705270,I357874);
nor I_41357 (I705151,I705513,I705753);
not I_41358 (I705814,I2690);
DFFARX1 I_41359 (I404440,I2683,I705814,I705840,);
DFFARX1 I_41360 (I404452,I2683,I705814,I705857,);
not I_41361 (I705865,I705857);
not I_41362 (I705882,I404437);
nor I_41363 (I705899,I705882,I404455);
not I_41364 (I705916,I404461);
nor I_41365 (I705933,I705899,I404443);
nor I_41366 (I705950,I705857,I705933);
DFFARX1 I_41367 (I705950,I2683,I705814,I705800,);
nor I_41368 (I705981,I404443,I404455);
nand I_41369 (I705998,I705981,I404437);
DFFARX1 I_41370 (I705998,I2683,I705814,I705803,);
nor I_41371 (I706029,I705916,I404443);
nand I_41372 (I706046,I706029,I404446);
nor I_41373 (I706063,I705840,I706046);
DFFARX1 I_41374 (I706063,I2683,I705814,I705779,);
not I_41375 (I706094,I706046);
nand I_41376 (I705791,I705857,I706094);
DFFARX1 I_41377 (I706046,I2683,I705814,I706134,);
not I_41378 (I706142,I706134);
not I_41379 (I706159,I404443);
not I_41380 (I706176,I404449);
nor I_41381 (I706193,I706176,I404461);
nor I_41382 (I705806,I706142,I706193);
nor I_41383 (I706224,I706176,I404458);
and I_41384 (I706241,I706224,I404437);
or I_41385 (I706258,I706241,I404440);
DFFARX1 I_41386 (I706258,I2683,I705814,I706284,);
nor I_41387 (I705794,I706284,I705840);
not I_41388 (I706306,I706284);
and I_41389 (I706323,I706306,I705840);
nor I_41390 (I705788,I705865,I706323);
nand I_41391 (I706354,I706306,I705916);
nor I_41392 (I705782,I706176,I706354);
nand I_41393 (I705785,I706306,I706094);
nand I_41394 (I706399,I705916,I404449);
nor I_41395 (I705797,I706159,I706399);
not I_41396 (I706460,I2690);
DFFARX1 I_41397 (I180111,I2683,I706460,I706486,);
DFFARX1 I_41398 (I180123,I2683,I706460,I706503,);
not I_41399 (I706511,I706503);
not I_41400 (I706528,I180129);
nor I_41401 (I706545,I706528,I180114);
not I_41402 (I706562,I180105);
nor I_41403 (I706579,I706545,I180126);
nor I_41404 (I706596,I706503,I706579);
DFFARX1 I_41405 (I706596,I2683,I706460,I706446,);
nor I_41406 (I706627,I180126,I180114);
nand I_41407 (I706644,I706627,I180129);
DFFARX1 I_41408 (I706644,I2683,I706460,I706449,);
nor I_41409 (I706675,I706562,I180126);
nand I_41410 (I706692,I706675,I180108);
nor I_41411 (I706709,I706486,I706692);
DFFARX1 I_41412 (I706709,I2683,I706460,I706425,);
not I_41413 (I706740,I706692);
nand I_41414 (I706437,I706503,I706740);
DFFARX1 I_41415 (I706692,I2683,I706460,I706780,);
not I_41416 (I706788,I706780);
not I_41417 (I706805,I180126);
not I_41418 (I706822,I180117);
nor I_41419 (I706839,I706822,I180105);
nor I_41420 (I706452,I706788,I706839);
nor I_41421 (I706870,I706822,I180120);
and I_41422 (I706887,I706870,I180108);
or I_41423 (I706904,I706887,I180105);
DFFARX1 I_41424 (I706904,I2683,I706460,I706930,);
nor I_41425 (I706440,I706930,I706486);
not I_41426 (I706952,I706930);
and I_41427 (I706969,I706952,I706486);
nor I_41428 (I706434,I706511,I706969);
nand I_41429 (I707000,I706952,I706562);
nor I_41430 (I706428,I706822,I707000);
nand I_41431 (I706431,I706952,I706740);
nand I_41432 (I707045,I706562,I180117);
nor I_41433 (I706443,I706805,I707045);
not I_41434 (I707106,I2690);
DFFARX1 I_41435 (I172376,I2683,I707106,I707132,);
DFFARX1 I_41436 (I172388,I2683,I707106,I707149,);
not I_41437 (I707157,I707149);
not I_41438 (I707174,I172394);
nor I_41439 (I707191,I707174,I172379);
not I_41440 (I707208,I172370);
nor I_41441 (I707225,I707191,I172391);
nor I_41442 (I707242,I707149,I707225);
DFFARX1 I_41443 (I707242,I2683,I707106,I707092,);
nor I_41444 (I707273,I172391,I172379);
nand I_41445 (I707290,I707273,I172394);
DFFARX1 I_41446 (I707290,I2683,I707106,I707095,);
nor I_41447 (I707321,I707208,I172391);
nand I_41448 (I707338,I707321,I172373);
nor I_41449 (I707355,I707132,I707338);
DFFARX1 I_41450 (I707355,I2683,I707106,I707071,);
not I_41451 (I707386,I707338);
nand I_41452 (I707083,I707149,I707386);
DFFARX1 I_41453 (I707338,I2683,I707106,I707426,);
not I_41454 (I707434,I707426);
not I_41455 (I707451,I172391);
not I_41456 (I707468,I172382);
nor I_41457 (I707485,I707468,I172370);
nor I_41458 (I707098,I707434,I707485);
nor I_41459 (I707516,I707468,I172385);
and I_41460 (I707533,I707516,I172373);
or I_41461 (I707550,I707533,I172370);
DFFARX1 I_41462 (I707550,I2683,I707106,I707576,);
nor I_41463 (I707086,I707576,I707132);
not I_41464 (I707598,I707576);
and I_41465 (I707615,I707598,I707132);
nor I_41466 (I707080,I707157,I707615);
nand I_41467 (I707646,I707598,I707208);
nor I_41468 (I707074,I707468,I707646);
nand I_41469 (I707077,I707598,I707386);
nand I_41470 (I707691,I707208,I172382);
nor I_41471 (I707089,I707451,I707691);
not I_41472 (I707752,I2690);
DFFARX1 I_41473 (I267502,I2683,I707752,I707778,);
DFFARX1 I_41474 (I267508,I2683,I707752,I707795,);
not I_41475 (I707803,I707795);
not I_41476 (I707820,I267529);
nor I_41477 (I707837,I707820,I267517);
not I_41478 (I707854,I267526);
nor I_41479 (I707871,I707837,I267511);
nor I_41480 (I707888,I707795,I707871);
DFFARX1 I_41481 (I707888,I2683,I707752,I707738,);
nor I_41482 (I707919,I267511,I267517);
nand I_41483 (I707936,I707919,I267529);
DFFARX1 I_41484 (I707936,I2683,I707752,I707741,);
nor I_41485 (I707967,I707854,I267511);
nand I_41486 (I707984,I707967,I267502);
nor I_41487 (I708001,I707778,I707984);
DFFARX1 I_41488 (I708001,I2683,I707752,I707717,);
not I_41489 (I708032,I707984);
nand I_41490 (I707729,I707795,I708032);
DFFARX1 I_41491 (I707984,I2683,I707752,I708072,);
not I_41492 (I708080,I708072);
not I_41493 (I708097,I267511);
not I_41494 (I708114,I267514);
nor I_41495 (I708131,I708114,I267526);
nor I_41496 (I707744,I708080,I708131);
nor I_41497 (I708162,I708114,I267523);
and I_41498 (I708179,I708162,I267505);
or I_41499 (I708196,I708179,I267520);
DFFARX1 I_41500 (I708196,I2683,I707752,I708222,);
nor I_41501 (I707732,I708222,I707778);
not I_41502 (I708244,I708222);
and I_41503 (I708261,I708244,I707778);
nor I_41504 (I707726,I707803,I708261);
nand I_41505 (I708292,I708244,I707854);
nor I_41506 (I707720,I708114,I708292);
nand I_41507 (I707723,I708244,I708032);
nand I_41508 (I708337,I707854,I267514);
nor I_41509 (I707735,I708097,I708337);
not I_41510 (I708398,I2690);
DFFARX1 I_41511 (I596560,I2683,I708398,I708424,);
DFFARX1 I_41512 (I596554,I2683,I708398,I708441,);
not I_41513 (I708449,I708441);
not I_41514 (I708466,I596569);
nor I_41515 (I708483,I708466,I596554);
not I_41516 (I708500,I596563);
nor I_41517 (I708517,I708483,I596572);
nor I_41518 (I708534,I708441,I708517);
DFFARX1 I_41519 (I708534,I2683,I708398,I708384,);
nor I_41520 (I708565,I596572,I596554);
nand I_41521 (I708582,I708565,I596569);
DFFARX1 I_41522 (I708582,I2683,I708398,I708387,);
nor I_41523 (I708613,I708500,I596572);
nand I_41524 (I708630,I708613,I596557);
nor I_41525 (I708647,I708424,I708630);
DFFARX1 I_41526 (I708647,I2683,I708398,I708363,);
not I_41527 (I708678,I708630);
nand I_41528 (I708375,I708441,I708678);
DFFARX1 I_41529 (I708630,I2683,I708398,I708718,);
not I_41530 (I708726,I708718);
not I_41531 (I708743,I596572);
not I_41532 (I708760,I596566);
nor I_41533 (I708777,I708760,I596563);
nor I_41534 (I708390,I708726,I708777);
nor I_41535 (I708808,I708760,I596575);
and I_41536 (I708825,I708808,I596578);
or I_41537 (I708842,I708825,I596557);
DFFARX1 I_41538 (I708842,I2683,I708398,I708868,);
nor I_41539 (I708378,I708868,I708424);
not I_41540 (I708890,I708868);
and I_41541 (I708907,I708890,I708424);
nor I_41542 (I708372,I708449,I708907);
nand I_41543 (I708938,I708890,I708500);
nor I_41544 (I708366,I708760,I708938);
nand I_41545 (I708369,I708890,I708678);
nand I_41546 (I708983,I708500,I596566);
nor I_41547 (I708381,I708743,I708983);
not I_41548 (I709044,I2690);
DFFARX1 I_41549 (I549164,I2683,I709044,I709070,);
DFFARX1 I_41550 (I549158,I2683,I709044,I709087,);
not I_41551 (I709095,I709087);
not I_41552 (I709112,I549173);
nor I_41553 (I709129,I709112,I549158);
not I_41554 (I709146,I549167);
nor I_41555 (I709163,I709129,I549176);
nor I_41556 (I709180,I709087,I709163);
DFFARX1 I_41557 (I709180,I2683,I709044,I709030,);
nor I_41558 (I709211,I549176,I549158);
nand I_41559 (I709228,I709211,I549173);
DFFARX1 I_41560 (I709228,I2683,I709044,I709033,);
nor I_41561 (I709259,I709146,I549176);
nand I_41562 (I709276,I709259,I549161);
nor I_41563 (I709293,I709070,I709276);
DFFARX1 I_41564 (I709293,I2683,I709044,I709009,);
not I_41565 (I709324,I709276);
nand I_41566 (I709021,I709087,I709324);
DFFARX1 I_41567 (I709276,I2683,I709044,I709364,);
not I_41568 (I709372,I709364);
not I_41569 (I709389,I549176);
not I_41570 (I709406,I549170);
nor I_41571 (I709423,I709406,I549167);
nor I_41572 (I709036,I709372,I709423);
nor I_41573 (I709454,I709406,I549179);
and I_41574 (I709471,I709454,I549182);
or I_41575 (I709488,I709471,I549161);
DFFARX1 I_41576 (I709488,I2683,I709044,I709514,);
nor I_41577 (I709024,I709514,I709070);
not I_41578 (I709536,I709514);
and I_41579 (I709553,I709536,I709070);
nor I_41580 (I709018,I709095,I709553);
nand I_41581 (I709584,I709536,I709146);
nor I_41582 (I709012,I709406,I709584);
nand I_41583 (I709015,I709536,I709324);
nand I_41584 (I709629,I709146,I549170);
nor I_41585 (I709027,I709389,I709629);
not I_41586 (I709690,I2690);
DFFARX1 I_41587 (I480379,I2683,I709690,I709716,);
DFFARX1 I_41588 (I480391,I2683,I709690,I709733,);
not I_41589 (I709741,I709733);
not I_41590 (I709758,I480400);
nor I_41591 (I709775,I709758,I480376);
not I_41592 (I709792,I480394);
nor I_41593 (I709809,I709775,I480388);
nor I_41594 (I709826,I709733,I709809);
DFFARX1 I_41595 (I709826,I2683,I709690,I709676,);
nor I_41596 (I709857,I480388,I480376);
nand I_41597 (I709874,I709857,I480400);
DFFARX1 I_41598 (I709874,I2683,I709690,I709679,);
nor I_41599 (I709905,I709792,I480388);
nand I_41600 (I709922,I709905,I480382);
nor I_41601 (I709939,I709716,I709922);
DFFARX1 I_41602 (I709939,I2683,I709690,I709655,);
not I_41603 (I709970,I709922);
nand I_41604 (I709667,I709733,I709970);
DFFARX1 I_41605 (I709922,I2683,I709690,I710010,);
not I_41606 (I710018,I710010);
not I_41607 (I710035,I480388);
not I_41608 (I710052,I480397);
nor I_41609 (I710069,I710052,I480394);
nor I_41610 (I709682,I710018,I710069);
nor I_41611 (I710100,I710052,I480379);
and I_41612 (I710117,I710100,I480376);
or I_41613 (I710134,I710117,I480385);
DFFARX1 I_41614 (I710134,I2683,I709690,I710160,);
nor I_41615 (I709670,I710160,I709716);
not I_41616 (I710182,I710160);
and I_41617 (I710199,I710182,I709716);
nor I_41618 (I709664,I709741,I710199);
nand I_41619 (I710230,I710182,I709792);
nor I_41620 (I709658,I710052,I710230);
nand I_41621 (I709661,I710182,I709970);
nand I_41622 (I710275,I709792,I480397);
nor I_41623 (I709673,I710035,I710275);
not I_41624 (I710336,I2690);
DFFARX1 I_41625 (I513906,I2683,I710336,I710362,);
DFFARX1 I_41626 (I513900,I2683,I710336,I710379,);
not I_41627 (I710387,I710379);
not I_41628 (I710404,I513915);
nor I_41629 (I710421,I710404,I513900);
not I_41630 (I710438,I513909);
nor I_41631 (I710455,I710421,I513918);
nor I_41632 (I710472,I710379,I710455);
DFFARX1 I_41633 (I710472,I2683,I710336,I710322,);
nor I_41634 (I710503,I513918,I513900);
nand I_41635 (I710520,I710503,I513915);
DFFARX1 I_41636 (I710520,I2683,I710336,I710325,);
nor I_41637 (I710551,I710438,I513918);
nand I_41638 (I710568,I710551,I513903);
nor I_41639 (I710585,I710362,I710568);
DFFARX1 I_41640 (I710585,I2683,I710336,I710301,);
not I_41641 (I710616,I710568);
nand I_41642 (I710313,I710379,I710616);
DFFARX1 I_41643 (I710568,I2683,I710336,I710656,);
not I_41644 (I710664,I710656);
not I_41645 (I710681,I513918);
not I_41646 (I710698,I513912);
nor I_41647 (I710715,I710698,I513909);
nor I_41648 (I710328,I710664,I710715);
nor I_41649 (I710746,I710698,I513921);
and I_41650 (I710763,I710746,I513924);
or I_41651 (I710780,I710763,I513903);
DFFARX1 I_41652 (I710780,I2683,I710336,I710806,);
nor I_41653 (I710316,I710806,I710362);
not I_41654 (I710828,I710806);
and I_41655 (I710845,I710828,I710362);
nor I_41656 (I710310,I710387,I710845);
nand I_41657 (I710876,I710828,I710438);
nor I_41658 (I710304,I710698,I710876);
nand I_41659 (I710307,I710828,I710616);
nand I_41660 (I710921,I710438,I513912);
nor I_41661 (I710319,I710681,I710921);
not I_41662 (I710982,I2690);
DFFARX1 I_41663 (I525466,I2683,I710982,I711008,);
DFFARX1 I_41664 (I525460,I2683,I710982,I711025,);
not I_41665 (I711033,I711025);
not I_41666 (I711050,I525475);
nor I_41667 (I711067,I711050,I525460);
not I_41668 (I711084,I525469);
nor I_41669 (I711101,I711067,I525478);
nor I_41670 (I711118,I711025,I711101);
DFFARX1 I_41671 (I711118,I2683,I710982,I710968,);
nor I_41672 (I711149,I525478,I525460);
nand I_41673 (I711166,I711149,I525475);
DFFARX1 I_41674 (I711166,I2683,I710982,I710971,);
nor I_41675 (I711197,I711084,I525478);
nand I_41676 (I711214,I711197,I525463);
nor I_41677 (I711231,I711008,I711214);
DFFARX1 I_41678 (I711231,I2683,I710982,I710947,);
not I_41679 (I711262,I711214);
nand I_41680 (I710959,I711025,I711262);
DFFARX1 I_41681 (I711214,I2683,I710982,I711302,);
not I_41682 (I711310,I711302);
not I_41683 (I711327,I525478);
not I_41684 (I711344,I525472);
nor I_41685 (I711361,I711344,I525469);
nor I_41686 (I710974,I711310,I711361);
nor I_41687 (I711392,I711344,I525481);
and I_41688 (I711409,I711392,I525484);
or I_41689 (I711426,I711409,I525463);
DFFARX1 I_41690 (I711426,I2683,I710982,I711452,);
nor I_41691 (I710962,I711452,I711008);
not I_41692 (I711474,I711452);
and I_41693 (I711491,I711474,I711008);
nor I_41694 (I710956,I711033,I711491);
nand I_41695 (I711522,I711474,I711084);
nor I_41696 (I710950,I711344,I711522);
nand I_41697 (I710953,I711474,I711262);
nand I_41698 (I711567,I711084,I525472);
nor I_41699 (I710965,I711327,I711567);
not I_41700 (I711628,I2690);
DFFARX1 I_41701 (I165236,I2683,I711628,I711654,);
DFFARX1 I_41702 (I165248,I2683,I711628,I711671,);
not I_41703 (I711679,I711671);
not I_41704 (I711696,I165254);
nor I_41705 (I711713,I711696,I165239);
not I_41706 (I711730,I165230);
nor I_41707 (I711747,I711713,I165251);
nor I_41708 (I711764,I711671,I711747);
DFFARX1 I_41709 (I711764,I2683,I711628,I711614,);
nor I_41710 (I711795,I165251,I165239);
nand I_41711 (I711812,I711795,I165254);
DFFARX1 I_41712 (I711812,I2683,I711628,I711617,);
nor I_41713 (I711843,I711730,I165251);
nand I_41714 (I711860,I711843,I165233);
nor I_41715 (I711877,I711654,I711860);
DFFARX1 I_41716 (I711877,I2683,I711628,I711593,);
not I_41717 (I711908,I711860);
nand I_41718 (I711605,I711671,I711908);
DFFARX1 I_41719 (I711860,I2683,I711628,I711948,);
not I_41720 (I711956,I711948);
not I_41721 (I711973,I165251);
not I_41722 (I711990,I165242);
nor I_41723 (I712007,I711990,I165230);
nor I_41724 (I711620,I711956,I712007);
nor I_41725 (I712038,I711990,I165245);
and I_41726 (I712055,I712038,I165233);
or I_41727 (I712072,I712055,I165230);
DFFARX1 I_41728 (I712072,I2683,I711628,I712098,);
nor I_41729 (I711608,I712098,I711654);
not I_41730 (I712120,I712098);
and I_41731 (I712137,I712120,I711654);
nor I_41732 (I711602,I711679,I712137);
nand I_41733 (I712168,I712120,I711730);
nor I_41734 (I711596,I711990,I712168);
nand I_41735 (I711599,I712120,I711908);
nand I_41736 (I712213,I711730,I165242);
nor I_41737 (I711611,I711973,I712213);
not I_41738 (I712274,I2690);
DFFARX1 I_41739 (I1077484,I2683,I712274,I712300,);
DFFARX1 I_41740 (I1077508,I2683,I712274,I712317,);
not I_41741 (I712325,I712317);
not I_41742 (I712342,I1077490);
nor I_41743 (I712359,I712342,I1077499);
not I_41744 (I712376,I1077484);
nor I_41745 (I712393,I712359,I1077505);
nor I_41746 (I712410,I712317,I712393);
DFFARX1 I_41747 (I712410,I2683,I712274,I712260,);
nor I_41748 (I712441,I1077505,I1077499);
nand I_41749 (I712458,I712441,I1077490);
DFFARX1 I_41750 (I712458,I2683,I712274,I712263,);
nor I_41751 (I712489,I712376,I1077505);
nand I_41752 (I712506,I712489,I1077502);
nor I_41753 (I712523,I712300,I712506);
DFFARX1 I_41754 (I712523,I2683,I712274,I712239,);
not I_41755 (I712554,I712506);
nand I_41756 (I712251,I712317,I712554);
DFFARX1 I_41757 (I712506,I2683,I712274,I712594,);
not I_41758 (I712602,I712594);
not I_41759 (I712619,I1077505);
not I_41760 (I712636,I1077496);
nor I_41761 (I712653,I712636,I1077484);
nor I_41762 (I712266,I712602,I712653);
nor I_41763 (I712684,I712636,I1077487);
and I_41764 (I712701,I712684,I1077511);
or I_41765 (I712718,I712701,I1077493);
DFFARX1 I_41766 (I712718,I2683,I712274,I712744,);
nor I_41767 (I712254,I712744,I712300);
not I_41768 (I712766,I712744);
and I_41769 (I712783,I712766,I712300);
nor I_41770 (I712248,I712325,I712783);
nand I_41771 (I712814,I712766,I712376);
nor I_41772 (I712242,I712636,I712814);
nand I_41773 (I712245,I712766,I712554);
nand I_41774 (I712859,I712376,I1077496);
nor I_41775 (I712257,I712619,I712859);
not I_41776 (I712920,I2690);
DFFARX1 I_41777 (I1070344,I2683,I712920,I712946,);
DFFARX1 I_41778 (I1070368,I2683,I712920,I712963,);
not I_41779 (I712971,I712963);
not I_41780 (I712988,I1070350);
nor I_41781 (I713005,I712988,I1070359);
not I_41782 (I713022,I1070344);
nor I_41783 (I713039,I713005,I1070365);
nor I_41784 (I713056,I712963,I713039);
DFFARX1 I_41785 (I713056,I2683,I712920,I712906,);
nor I_41786 (I713087,I1070365,I1070359);
nand I_41787 (I713104,I713087,I1070350);
DFFARX1 I_41788 (I713104,I2683,I712920,I712909,);
nor I_41789 (I713135,I713022,I1070365);
nand I_41790 (I713152,I713135,I1070362);
nor I_41791 (I713169,I712946,I713152);
DFFARX1 I_41792 (I713169,I2683,I712920,I712885,);
not I_41793 (I713200,I713152);
nand I_41794 (I712897,I712963,I713200);
DFFARX1 I_41795 (I713152,I2683,I712920,I713240,);
not I_41796 (I713248,I713240);
not I_41797 (I713265,I1070365);
not I_41798 (I713282,I1070356);
nor I_41799 (I713299,I713282,I1070344);
nor I_41800 (I712912,I713248,I713299);
nor I_41801 (I713330,I713282,I1070347);
and I_41802 (I713347,I713330,I1070371);
or I_41803 (I713364,I713347,I1070353);
DFFARX1 I_41804 (I713364,I2683,I712920,I713390,);
nor I_41805 (I712900,I713390,I712946);
not I_41806 (I713412,I713390);
and I_41807 (I713429,I713412,I712946);
nor I_41808 (I712894,I712971,I713429);
nand I_41809 (I713460,I713412,I713022);
nor I_41810 (I712888,I713282,I713460);
nand I_41811 (I712891,I713412,I713200);
nand I_41812 (I713505,I713022,I1070356);
nor I_41813 (I712903,I713265,I713505);
not I_41814 (I713566,I2690);
DFFARX1 I_41815 (I988048,I2683,I713566,I713592,);
DFFARX1 I_41816 (I988054,I2683,I713566,I713609,);
not I_41817 (I713617,I713609);
not I_41818 (I713634,I988051);
nor I_41819 (I713651,I713634,I988030);
not I_41820 (I713668,I988033);
nor I_41821 (I713685,I713651,I988039);
nor I_41822 (I713702,I713609,I713685);
DFFARX1 I_41823 (I713702,I2683,I713566,I713552,);
nor I_41824 (I713733,I988039,I988030);
nand I_41825 (I713750,I713733,I988051);
DFFARX1 I_41826 (I713750,I2683,I713566,I713555,);
nor I_41827 (I713781,I713668,I988039);
nand I_41828 (I713798,I713781,I988033);
nor I_41829 (I713815,I713592,I713798);
DFFARX1 I_41830 (I713815,I2683,I713566,I713531,);
not I_41831 (I713846,I713798);
nand I_41832 (I713543,I713609,I713846);
DFFARX1 I_41833 (I713798,I2683,I713566,I713886,);
not I_41834 (I713894,I713886);
not I_41835 (I713911,I988039);
not I_41836 (I713928,I988042);
nor I_41837 (I713945,I713928,I988033);
nor I_41838 (I713558,I713894,I713945);
nor I_41839 (I713976,I713928,I988030);
and I_41840 (I713993,I713976,I988036);
or I_41841 (I714010,I713993,I988045);
DFFARX1 I_41842 (I714010,I2683,I713566,I714036,);
nor I_41843 (I713546,I714036,I713592);
not I_41844 (I714058,I714036);
and I_41845 (I714075,I714058,I713592);
nor I_41846 (I713540,I713617,I714075);
nand I_41847 (I714106,I714058,I713668);
nor I_41848 (I713534,I713928,I714106);
nand I_41849 (I713537,I714058,I713846);
nand I_41850 (I714151,I713668,I988042);
nor I_41851 (I713549,I713911,I714151);
not I_41852 (I714212,I2690);
DFFARX1 I_41853 (I48508,I2683,I714212,I714238,);
DFFARX1 I_41854 (I48514,I2683,I714212,I714255,);
not I_41855 (I714263,I714255);
not I_41856 (I714280,I48532);
nor I_41857 (I714297,I714280,I48511);
not I_41858 (I714314,I48517);
nor I_41859 (I714331,I714297,I48523);
nor I_41860 (I714348,I714255,I714331);
DFFARX1 I_41861 (I714348,I2683,I714212,I714198,);
nor I_41862 (I714379,I48523,I48511);
nand I_41863 (I714396,I714379,I48532);
DFFARX1 I_41864 (I714396,I2683,I714212,I714201,);
nor I_41865 (I714427,I714314,I48523);
nand I_41866 (I714444,I714427,I48529);
nor I_41867 (I714461,I714238,I714444);
DFFARX1 I_41868 (I714461,I2683,I714212,I714177,);
not I_41869 (I714492,I714444);
nand I_41870 (I714189,I714255,I714492);
DFFARX1 I_41871 (I714444,I2683,I714212,I714532,);
not I_41872 (I714540,I714532);
not I_41873 (I714557,I48523);
not I_41874 (I714574,I48511);
nor I_41875 (I714591,I714574,I48517);
nor I_41876 (I714204,I714540,I714591);
nor I_41877 (I714622,I714574,I48520);
and I_41878 (I714639,I714622,I48508);
or I_41879 (I714656,I714639,I48526);
DFFARX1 I_41880 (I714656,I2683,I714212,I714682,);
nor I_41881 (I714192,I714682,I714238);
not I_41882 (I714704,I714682);
and I_41883 (I714721,I714704,I714238);
nor I_41884 (I714186,I714263,I714721);
nand I_41885 (I714752,I714704,I714314);
nor I_41886 (I714180,I714574,I714752);
nand I_41887 (I714183,I714704,I714492);
nand I_41888 (I714797,I714314,I48511);
nor I_41889 (I714195,I714557,I714797);
not I_41890 (I714858,I2690);
DFFARX1 I_41891 (I278042,I2683,I714858,I714884,);
DFFARX1 I_41892 (I278048,I2683,I714858,I714901,);
not I_41893 (I714909,I714901);
not I_41894 (I714926,I278069);
nor I_41895 (I714943,I714926,I278057);
not I_41896 (I714960,I278066);
nor I_41897 (I714977,I714943,I278051);
nor I_41898 (I714994,I714901,I714977);
DFFARX1 I_41899 (I714994,I2683,I714858,I714844,);
nor I_41900 (I715025,I278051,I278057);
nand I_41901 (I715042,I715025,I278069);
DFFARX1 I_41902 (I715042,I2683,I714858,I714847,);
nor I_41903 (I715073,I714960,I278051);
nand I_41904 (I715090,I715073,I278042);
nor I_41905 (I715107,I714884,I715090);
DFFARX1 I_41906 (I715107,I2683,I714858,I714823,);
not I_41907 (I715138,I715090);
nand I_41908 (I714835,I714901,I715138);
DFFARX1 I_41909 (I715090,I2683,I714858,I715178,);
not I_41910 (I715186,I715178);
not I_41911 (I715203,I278051);
not I_41912 (I715220,I278054);
nor I_41913 (I715237,I715220,I278066);
nor I_41914 (I714850,I715186,I715237);
nor I_41915 (I715268,I715220,I278063);
and I_41916 (I715285,I715268,I278045);
or I_41917 (I715302,I715285,I278060);
DFFARX1 I_41918 (I715302,I2683,I714858,I715328,);
nor I_41919 (I714838,I715328,I714884);
not I_41920 (I715350,I715328);
and I_41921 (I715367,I715350,I714884);
nor I_41922 (I714832,I714909,I715367);
nand I_41923 (I715398,I715350,I714960);
nor I_41924 (I714826,I715220,I715398);
nand I_41925 (I714829,I715350,I715138);
nand I_41926 (I715443,I714960,I278054);
nor I_41927 (I714841,I715203,I715443);
not I_41928 (I715504,I2690);
DFFARX1 I_41929 (I308608,I2683,I715504,I715530,);
DFFARX1 I_41930 (I308614,I2683,I715504,I715547,);
not I_41931 (I715555,I715547);
not I_41932 (I715572,I308635);
nor I_41933 (I715589,I715572,I308623);
not I_41934 (I715606,I308632);
nor I_41935 (I715623,I715589,I308617);
nor I_41936 (I715640,I715547,I715623);
DFFARX1 I_41937 (I715640,I2683,I715504,I715490,);
nor I_41938 (I715671,I308617,I308623);
nand I_41939 (I715688,I715671,I308635);
DFFARX1 I_41940 (I715688,I2683,I715504,I715493,);
nor I_41941 (I715719,I715606,I308617);
nand I_41942 (I715736,I715719,I308608);
nor I_41943 (I715753,I715530,I715736);
DFFARX1 I_41944 (I715753,I2683,I715504,I715469,);
not I_41945 (I715784,I715736);
nand I_41946 (I715481,I715547,I715784);
DFFARX1 I_41947 (I715736,I2683,I715504,I715824,);
not I_41948 (I715832,I715824);
not I_41949 (I715849,I308617);
not I_41950 (I715866,I308620);
nor I_41951 (I715883,I715866,I308632);
nor I_41952 (I715496,I715832,I715883);
nor I_41953 (I715914,I715866,I308629);
and I_41954 (I715931,I715914,I308611);
or I_41955 (I715948,I715931,I308626);
DFFARX1 I_41956 (I715948,I2683,I715504,I715974,);
nor I_41957 (I715484,I715974,I715530);
not I_41958 (I715996,I715974);
and I_41959 (I716013,I715996,I715530);
nor I_41960 (I715478,I715555,I716013);
nand I_41961 (I716044,I715996,I715606);
nor I_41962 (I715472,I715866,I716044);
nand I_41963 (I715475,I715996,I715784);
nand I_41964 (I716089,I715606,I308620);
nor I_41965 (I715487,I715849,I716089);
not I_41966 (I716150,I2690);
DFFARX1 I_41967 (I654938,I2683,I716150,I716176,);
DFFARX1 I_41968 (I654935,I2683,I716150,I716193,);
not I_41969 (I716201,I716193);
not I_41970 (I716218,I654935);
nor I_41971 (I716235,I716218,I654938);
not I_41972 (I716252,I654950);
nor I_41973 (I716269,I716235,I654944);
nor I_41974 (I716286,I716193,I716269);
DFFARX1 I_41975 (I716286,I2683,I716150,I716136,);
nor I_41976 (I716317,I654944,I654938);
nand I_41977 (I716334,I716317,I654935);
DFFARX1 I_41978 (I716334,I2683,I716150,I716139,);
nor I_41979 (I716365,I716252,I654944);
nand I_41980 (I716382,I716365,I654932);
nor I_41981 (I716399,I716176,I716382);
DFFARX1 I_41982 (I716399,I2683,I716150,I716115,);
not I_41983 (I716430,I716382);
nand I_41984 (I716127,I716193,I716430);
DFFARX1 I_41985 (I716382,I2683,I716150,I716470,);
not I_41986 (I716478,I716470);
not I_41987 (I716495,I654944);
not I_41988 (I716512,I654941);
nor I_41989 (I716529,I716512,I654950);
nor I_41990 (I716142,I716478,I716529);
nor I_41991 (I716560,I716512,I654947);
and I_41992 (I716577,I716560,I654953);
or I_41993 (I716594,I716577,I654932);
DFFARX1 I_41994 (I716594,I2683,I716150,I716620,);
nor I_41995 (I716130,I716620,I716176);
not I_41996 (I716642,I716620);
and I_41997 (I716659,I716642,I716176);
nor I_41998 (I716124,I716201,I716659);
nand I_41999 (I716690,I716642,I716252);
nor I_42000 (I716118,I716512,I716690);
nand I_42001 (I716121,I716642,I716430);
nand I_42002 (I716735,I716252,I654941);
nor I_42003 (I716133,I716495,I716735);
not I_42004 (I716796,I2690);
DFFARX1 I_42005 (I345368,I2683,I716796,I716822,);
DFFARX1 I_42006 (I345365,I2683,I716796,I716839,);
not I_42007 (I716847,I716839);
not I_42008 (I716864,I345380);
nor I_42009 (I716881,I716864,I345383);
not I_42010 (I716898,I345371);
nor I_42011 (I716915,I716881,I345377);
nor I_42012 (I716932,I716839,I716915);
DFFARX1 I_42013 (I716932,I2683,I716796,I716782,);
nor I_42014 (I716963,I345377,I345383);
nand I_42015 (I716980,I716963,I345380);
DFFARX1 I_42016 (I716980,I2683,I716796,I716785,);
nor I_42017 (I717011,I716898,I345377);
nand I_42018 (I717028,I717011,I345389);
nor I_42019 (I717045,I716822,I717028);
DFFARX1 I_42020 (I717045,I2683,I716796,I716761,);
not I_42021 (I717076,I717028);
nand I_42022 (I716773,I716839,I717076);
DFFARX1 I_42023 (I717028,I2683,I716796,I717116,);
not I_42024 (I717124,I717116);
not I_42025 (I717141,I345377);
not I_42026 (I717158,I345362);
nor I_42027 (I717175,I717158,I345371);
nor I_42028 (I716788,I717124,I717175);
nor I_42029 (I717206,I717158,I345374);
and I_42030 (I717223,I717206,I345362);
or I_42031 (I717240,I717223,I345386);
DFFARX1 I_42032 (I717240,I2683,I716796,I717266,);
nor I_42033 (I716776,I717266,I716822);
not I_42034 (I717288,I717266);
and I_42035 (I717305,I717288,I716822);
nor I_42036 (I716770,I716847,I717305);
nand I_42037 (I717336,I717288,I716898);
nor I_42038 (I716764,I717158,I717336);
nand I_42039 (I716767,I717288,I717076);
nand I_42040 (I717381,I716898,I345362);
nor I_42041 (I716779,I717141,I717381);
not I_42042 (I717442,I2690);
DFFARX1 I_42043 (I1067964,I2683,I717442,I717468,);
DFFARX1 I_42044 (I1067988,I2683,I717442,I717485,);
not I_42045 (I717493,I717485);
not I_42046 (I717510,I1067970);
nor I_42047 (I717527,I717510,I1067979);
not I_42048 (I717544,I1067964);
nor I_42049 (I717561,I717527,I1067985);
nor I_42050 (I717578,I717485,I717561);
DFFARX1 I_42051 (I717578,I2683,I717442,I717428,);
nor I_42052 (I717609,I1067985,I1067979);
nand I_42053 (I717626,I717609,I1067970);
DFFARX1 I_42054 (I717626,I2683,I717442,I717431,);
nor I_42055 (I717657,I717544,I1067985);
nand I_42056 (I717674,I717657,I1067982);
nor I_42057 (I717691,I717468,I717674);
DFFARX1 I_42058 (I717691,I2683,I717442,I717407,);
not I_42059 (I717722,I717674);
nand I_42060 (I717419,I717485,I717722);
DFFARX1 I_42061 (I717674,I2683,I717442,I717762,);
not I_42062 (I717770,I717762);
not I_42063 (I717787,I1067985);
not I_42064 (I717804,I1067976);
nor I_42065 (I717821,I717804,I1067964);
nor I_42066 (I717434,I717770,I717821);
nor I_42067 (I717852,I717804,I1067967);
and I_42068 (I717869,I717852,I1067991);
or I_42069 (I717886,I717869,I1067973);
DFFARX1 I_42070 (I717886,I2683,I717442,I717912,);
nor I_42071 (I717422,I717912,I717468);
not I_42072 (I717934,I717912);
and I_42073 (I717951,I717934,I717468);
nor I_42074 (I717416,I717493,I717951);
nand I_42075 (I717982,I717934,I717544);
nor I_42076 (I717410,I717804,I717982);
nand I_42077 (I717413,I717934,I717722);
nand I_42078 (I718027,I717544,I1067976);
nor I_42079 (I717425,I717787,I718027);
not I_42080 (I718088,I2690);
DFFARX1 I_42081 (I71696,I2683,I718088,I718114,);
DFFARX1 I_42082 (I71702,I2683,I718088,I718131,);
not I_42083 (I718139,I718131);
not I_42084 (I718156,I71720);
nor I_42085 (I718173,I718156,I71699);
not I_42086 (I718190,I71705);
nor I_42087 (I718207,I718173,I71711);
nor I_42088 (I718224,I718131,I718207);
DFFARX1 I_42089 (I718224,I2683,I718088,I718074,);
nor I_42090 (I718255,I71711,I71699);
nand I_42091 (I718272,I718255,I71720);
DFFARX1 I_42092 (I718272,I2683,I718088,I718077,);
nor I_42093 (I718303,I718190,I71711);
nand I_42094 (I718320,I718303,I71717);
nor I_42095 (I718337,I718114,I718320);
DFFARX1 I_42096 (I718337,I2683,I718088,I718053,);
not I_42097 (I718368,I718320);
nand I_42098 (I718065,I718131,I718368);
DFFARX1 I_42099 (I718320,I2683,I718088,I718408,);
not I_42100 (I718416,I718408);
not I_42101 (I718433,I71711);
not I_42102 (I718450,I71699);
nor I_42103 (I718467,I718450,I71705);
nor I_42104 (I718080,I718416,I718467);
nor I_42105 (I718498,I718450,I71708);
and I_42106 (I718515,I718498,I71696);
or I_42107 (I718532,I718515,I71714);
DFFARX1 I_42108 (I718532,I2683,I718088,I718558,);
nor I_42109 (I718068,I718558,I718114);
not I_42110 (I718580,I718558);
and I_42111 (I718597,I718580,I718114);
nor I_42112 (I718062,I718139,I718597);
nand I_42113 (I718628,I718580,I718190);
nor I_42114 (I718056,I718450,I718628);
nand I_42115 (I718059,I718580,I718368);
nand I_42116 (I718673,I718190,I71699);
nor I_42117 (I718071,I718433,I718673);
not I_42118 (I718734,I2690);
DFFARX1 I_42119 (I45873,I2683,I718734,I718760,);
DFFARX1 I_42120 (I45879,I2683,I718734,I718777,);
not I_42121 (I718785,I718777);
not I_42122 (I718802,I45873);
nor I_42123 (I718819,I718802,I45885);
not I_42124 (I718836,I45897);
nor I_42125 (I718853,I718819,I45891);
nor I_42126 (I718870,I718777,I718853);
DFFARX1 I_42127 (I718870,I2683,I718734,I718720,);
nor I_42128 (I718901,I45891,I45885);
nand I_42129 (I718918,I718901,I45873);
DFFARX1 I_42130 (I718918,I2683,I718734,I718723,);
nor I_42131 (I718949,I718836,I45891);
nand I_42132 (I718966,I718949,I45876);
nor I_42133 (I718983,I718760,I718966);
DFFARX1 I_42134 (I718983,I2683,I718734,I718699,);
not I_42135 (I719014,I718966);
nand I_42136 (I718711,I718777,I719014);
DFFARX1 I_42137 (I718966,I2683,I718734,I719054,);
not I_42138 (I719062,I719054);
not I_42139 (I719079,I45891);
not I_42140 (I719096,I45876);
nor I_42141 (I719113,I719096,I45897);
nor I_42142 (I718726,I719062,I719113);
nor I_42143 (I719144,I719096,I45894);
and I_42144 (I719161,I719144,I45888);
or I_42145 (I719178,I719161,I45882);
DFFARX1 I_42146 (I719178,I2683,I718734,I719204,);
nor I_42147 (I718714,I719204,I718760);
not I_42148 (I719226,I719204);
and I_42149 (I719243,I719226,I718760);
nor I_42150 (I718708,I718785,I719243);
nand I_42151 (I719274,I719226,I718836);
nor I_42152 (I718702,I719096,I719274);
nand I_42153 (I718705,I719226,I719014);
nand I_42154 (I719319,I718836,I45876);
nor I_42155 (I718717,I719079,I719319);
not I_42156 (I719380,I2690);
DFFARX1 I_42157 (I140246,I2683,I719380,I719406,);
DFFARX1 I_42158 (I140258,I2683,I719380,I719423,);
not I_42159 (I719431,I719423);
not I_42160 (I719448,I140264);
nor I_42161 (I719465,I719448,I140249);
not I_42162 (I719482,I140240);
nor I_42163 (I719499,I719465,I140261);
nor I_42164 (I719516,I719423,I719499);
DFFARX1 I_42165 (I719516,I2683,I719380,I719366,);
nor I_42166 (I719547,I140261,I140249);
nand I_42167 (I719564,I719547,I140264);
DFFARX1 I_42168 (I719564,I2683,I719380,I719369,);
nor I_42169 (I719595,I719482,I140261);
nand I_42170 (I719612,I719595,I140243);
nor I_42171 (I719629,I719406,I719612);
DFFARX1 I_42172 (I719629,I2683,I719380,I719345,);
not I_42173 (I719660,I719612);
nand I_42174 (I719357,I719423,I719660);
DFFARX1 I_42175 (I719612,I2683,I719380,I719700,);
not I_42176 (I719708,I719700);
not I_42177 (I719725,I140261);
not I_42178 (I719742,I140252);
nor I_42179 (I719759,I719742,I140240);
nor I_42180 (I719372,I719708,I719759);
nor I_42181 (I719790,I719742,I140255);
and I_42182 (I719807,I719790,I140243);
or I_42183 (I719824,I719807,I140240);
DFFARX1 I_42184 (I719824,I2683,I719380,I719850,);
nor I_42185 (I719360,I719850,I719406);
not I_42186 (I719872,I719850);
and I_42187 (I719889,I719872,I719406);
nor I_42188 (I719354,I719431,I719889);
nand I_42189 (I719920,I719872,I719482);
nor I_42190 (I719348,I719742,I719920);
nand I_42191 (I719351,I719872,I719660);
nand I_42192 (I719965,I719482,I140252);
nor I_42193 (I719363,I719725,I719965);
not I_42194 (I720026,I2690);
DFFARX1 I_42195 (I593670,I2683,I720026,I720052,);
DFFARX1 I_42196 (I593664,I2683,I720026,I720069,);
not I_42197 (I720077,I720069);
not I_42198 (I720094,I593679);
nor I_42199 (I720111,I720094,I593664);
not I_42200 (I720128,I593673);
nor I_42201 (I720145,I720111,I593682);
nor I_42202 (I720162,I720069,I720145);
DFFARX1 I_42203 (I720162,I2683,I720026,I720012,);
nor I_42204 (I720193,I593682,I593664);
nand I_42205 (I720210,I720193,I593679);
DFFARX1 I_42206 (I720210,I2683,I720026,I720015,);
nor I_42207 (I720241,I720128,I593682);
nand I_42208 (I720258,I720241,I593667);
nor I_42209 (I720275,I720052,I720258);
DFFARX1 I_42210 (I720275,I2683,I720026,I719991,);
not I_42211 (I720306,I720258);
nand I_42212 (I720003,I720069,I720306);
DFFARX1 I_42213 (I720258,I2683,I720026,I720346,);
not I_42214 (I720354,I720346);
not I_42215 (I720371,I593682);
not I_42216 (I720388,I593676);
nor I_42217 (I720405,I720388,I593673);
nor I_42218 (I720018,I720354,I720405);
nor I_42219 (I720436,I720388,I593685);
and I_42220 (I720453,I720436,I593688);
or I_42221 (I720470,I720453,I593667);
DFFARX1 I_42222 (I720470,I2683,I720026,I720496,);
nor I_42223 (I720006,I720496,I720052);
not I_42224 (I720518,I720496);
and I_42225 (I720535,I720518,I720052);
nor I_42226 (I720000,I720077,I720535);
nand I_42227 (I720566,I720518,I720128);
nor I_42228 (I719994,I720388,I720566);
nand I_42229 (I719997,I720518,I720306);
nand I_42230 (I720611,I720128,I593676);
nor I_42231 (I720009,I720371,I720611);
not I_42232 (I720672,I2690);
DFFARX1 I_42233 (I530668,I2683,I720672,I720698,);
DFFARX1 I_42234 (I530662,I2683,I720672,I720715,);
not I_42235 (I720723,I720715);
not I_42236 (I720740,I530677);
nor I_42237 (I720757,I720740,I530662);
not I_42238 (I720774,I530671);
nor I_42239 (I720791,I720757,I530680);
nor I_42240 (I720808,I720715,I720791);
DFFARX1 I_42241 (I720808,I2683,I720672,I720658,);
nor I_42242 (I720839,I530680,I530662);
nand I_42243 (I720856,I720839,I530677);
DFFARX1 I_42244 (I720856,I2683,I720672,I720661,);
nor I_42245 (I720887,I720774,I530680);
nand I_42246 (I720904,I720887,I530665);
nor I_42247 (I720921,I720698,I720904);
DFFARX1 I_42248 (I720921,I2683,I720672,I720637,);
not I_42249 (I720952,I720904);
nand I_42250 (I720649,I720715,I720952);
DFFARX1 I_42251 (I720904,I2683,I720672,I720992,);
not I_42252 (I721000,I720992);
not I_42253 (I721017,I530680);
not I_42254 (I721034,I530674);
nor I_42255 (I721051,I721034,I530671);
nor I_42256 (I720664,I721000,I721051);
nor I_42257 (I721082,I721034,I530683);
and I_42258 (I721099,I721082,I530686);
or I_42259 (I721116,I721099,I530665);
DFFARX1 I_42260 (I721116,I2683,I720672,I721142,);
nor I_42261 (I720652,I721142,I720698);
not I_42262 (I721164,I721142);
and I_42263 (I721181,I721164,I720698);
nor I_42264 (I720646,I720723,I721181);
nand I_42265 (I721212,I721164,I720774);
nor I_42266 (I720640,I721034,I721212);
nand I_42267 (I720643,I721164,I720952);
nand I_42268 (I721257,I720774,I530674);
nor I_42269 (I720655,I721017,I721257);
not I_42270 (I721318,I2690);
DFFARX1 I_42271 (I64318,I2683,I721318,I721344,);
DFFARX1 I_42272 (I64324,I2683,I721318,I721361,);
not I_42273 (I721369,I721361);
not I_42274 (I721386,I64342);
nor I_42275 (I721403,I721386,I64321);
not I_42276 (I721420,I64327);
nor I_42277 (I721437,I721403,I64333);
nor I_42278 (I721454,I721361,I721437);
DFFARX1 I_42279 (I721454,I2683,I721318,I721304,);
nor I_42280 (I721485,I64333,I64321);
nand I_42281 (I721502,I721485,I64342);
DFFARX1 I_42282 (I721502,I2683,I721318,I721307,);
nor I_42283 (I721533,I721420,I64333);
nand I_42284 (I721550,I721533,I64339);
nor I_42285 (I721567,I721344,I721550);
DFFARX1 I_42286 (I721567,I2683,I721318,I721283,);
not I_42287 (I721598,I721550);
nand I_42288 (I721295,I721361,I721598);
DFFARX1 I_42289 (I721550,I2683,I721318,I721638,);
not I_42290 (I721646,I721638);
not I_42291 (I721663,I64333);
not I_42292 (I721680,I64321);
nor I_42293 (I721697,I721680,I64327);
nor I_42294 (I721310,I721646,I721697);
nor I_42295 (I721728,I721680,I64330);
and I_42296 (I721745,I721728,I64318);
or I_42297 (I721762,I721745,I64336);
DFFARX1 I_42298 (I721762,I2683,I721318,I721788,);
nor I_42299 (I721298,I721788,I721344);
not I_42300 (I721810,I721788);
and I_42301 (I721827,I721810,I721344);
nor I_42302 (I721292,I721369,I721827);
nand I_42303 (I721858,I721810,I721420);
nor I_42304 (I721286,I721680,I721858);
nand I_42305 (I721289,I721810,I721598);
nand I_42306 (I721903,I721420,I64321);
nor I_42307 (I721301,I721663,I721903);
not I_42308 (I721964,I2690);
DFFARX1 I_42309 (I1063204,I2683,I721964,I721990,);
DFFARX1 I_42310 (I1063228,I2683,I721964,I722007,);
not I_42311 (I722015,I722007);
not I_42312 (I722032,I1063210);
nor I_42313 (I722049,I722032,I1063219);
not I_42314 (I722066,I1063204);
nor I_42315 (I722083,I722049,I1063225);
nor I_42316 (I722100,I722007,I722083);
DFFARX1 I_42317 (I722100,I2683,I721964,I721950,);
nor I_42318 (I722131,I1063225,I1063219);
nand I_42319 (I722148,I722131,I1063210);
DFFARX1 I_42320 (I722148,I2683,I721964,I721953,);
nor I_42321 (I722179,I722066,I1063225);
nand I_42322 (I722196,I722179,I1063222);
nor I_42323 (I722213,I721990,I722196);
DFFARX1 I_42324 (I722213,I2683,I721964,I721929,);
not I_42325 (I722244,I722196);
nand I_42326 (I721941,I722007,I722244);
DFFARX1 I_42327 (I722196,I2683,I721964,I722284,);
not I_42328 (I722292,I722284);
not I_42329 (I722309,I1063225);
not I_42330 (I722326,I1063216);
nor I_42331 (I722343,I722326,I1063204);
nor I_42332 (I721956,I722292,I722343);
nor I_42333 (I722374,I722326,I1063207);
and I_42334 (I722391,I722374,I1063231);
or I_42335 (I722408,I722391,I1063213);
DFFARX1 I_42336 (I722408,I2683,I721964,I722434,);
nor I_42337 (I721944,I722434,I721990);
not I_42338 (I722456,I722434);
and I_42339 (I722473,I722456,I721990);
nor I_42340 (I721938,I722015,I722473);
nand I_42341 (I722504,I722456,I722066);
nor I_42342 (I721932,I722326,I722504);
nand I_42343 (I721935,I722456,I722244);
nand I_42344 (I722549,I722066,I1063216);
nor I_42345 (I721947,I722309,I722549);
not I_42346 (I722610,I2690);
DFFARX1 I_42347 (I119433,I2683,I722610,I722636,);
DFFARX1 I_42348 (I119436,I2683,I722610,I722653,);
not I_42349 (I722661,I722653);
not I_42350 (I722678,I119421);
nor I_42351 (I722695,I722678,I119415);
not I_42352 (I722712,I119424);
nor I_42353 (I722729,I722695,I119439);
nor I_42354 (I722746,I722653,I722729);
DFFARX1 I_42355 (I722746,I2683,I722610,I722596,);
nor I_42356 (I722777,I119439,I119415);
nand I_42357 (I722794,I722777,I119421);
DFFARX1 I_42358 (I722794,I2683,I722610,I722599,);
nor I_42359 (I722825,I722712,I119439);
nand I_42360 (I722842,I722825,I119442);
nor I_42361 (I722859,I722636,I722842);
DFFARX1 I_42362 (I722859,I2683,I722610,I722575,);
not I_42363 (I722890,I722842);
nand I_42364 (I722587,I722653,I722890);
DFFARX1 I_42365 (I722842,I2683,I722610,I722930,);
not I_42366 (I722938,I722930);
not I_42367 (I722955,I119439);
not I_42368 (I722972,I119418);
nor I_42369 (I722989,I722972,I119424);
nor I_42370 (I722602,I722938,I722989);
nor I_42371 (I723020,I722972,I119427);
and I_42372 (I723037,I723020,I119415);
or I_42373 (I723054,I723037,I119430);
DFFARX1 I_42374 (I723054,I2683,I722610,I723080,);
nor I_42375 (I722590,I723080,I722636);
not I_42376 (I723102,I723080);
and I_42377 (I723119,I723102,I722636);
nor I_42378 (I722584,I722661,I723119);
nand I_42379 (I723150,I723102,I722712);
nor I_42380 (I722578,I722972,I723150);
nand I_42381 (I722581,I723102,I722890);
nand I_42382 (I723195,I722712,I119418);
nor I_42383 (I722593,I722955,I723195);
not I_42384 (I723256,I2690);
DFFARX1 I_42385 (I488471,I2683,I723256,I723282,);
DFFARX1 I_42386 (I488483,I2683,I723256,I723299,);
not I_42387 (I723307,I723299);
not I_42388 (I723324,I488492);
nor I_42389 (I723341,I723324,I488468);
not I_42390 (I723358,I488486);
nor I_42391 (I723375,I723341,I488480);
nor I_42392 (I723392,I723299,I723375);
DFFARX1 I_42393 (I723392,I2683,I723256,I723242,);
nor I_42394 (I723423,I488480,I488468);
nand I_42395 (I723440,I723423,I488492);
DFFARX1 I_42396 (I723440,I2683,I723256,I723245,);
nor I_42397 (I723471,I723358,I488480);
nand I_42398 (I723488,I723471,I488474);
nor I_42399 (I723505,I723282,I723488);
DFFARX1 I_42400 (I723505,I2683,I723256,I723221,);
not I_42401 (I723536,I723488);
nand I_42402 (I723233,I723299,I723536);
DFFARX1 I_42403 (I723488,I2683,I723256,I723576,);
not I_42404 (I723584,I723576);
not I_42405 (I723601,I488480);
not I_42406 (I723618,I488489);
nor I_42407 (I723635,I723618,I488486);
nor I_42408 (I723248,I723584,I723635);
nor I_42409 (I723666,I723618,I488471);
and I_42410 (I723683,I723666,I488468);
or I_42411 (I723700,I723683,I488477);
DFFARX1 I_42412 (I723700,I2683,I723256,I723726,);
nor I_42413 (I723236,I723726,I723282);
not I_42414 (I723748,I723726);
and I_42415 (I723765,I723748,I723282);
nor I_42416 (I723230,I723307,I723765);
nand I_42417 (I723796,I723748,I723358);
nor I_42418 (I723224,I723618,I723796);
nand I_42419 (I723227,I723748,I723536);
nand I_42420 (I723841,I723358,I488489);
nor I_42421 (I723239,I723601,I723841);
not I_42422 (I723902,I2690);
DFFARX1 I_42423 (I1095334,I2683,I723902,I723928,);
DFFARX1 I_42424 (I1095358,I2683,I723902,I723945,);
not I_42425 (I723953,I723945);
not I_42426 (I723970,I1095340);
nor I_42427 (I723987,I723970,I1095349);
not I_42428 (I724004,I1095334);
nor I_42429 (I724021,I723987,I1095355);
nor I_42430 (I724038,I723945,I724021);
DFFARX1 I_42431 (I724038,I2683,I723902,I723888,);
nor I_42432 (I724069,I1095355,I1095349);
nand I_42433 (I724086,I724069,I1095340);
DFFARX1 I_42434 (I724086,I2683,I723902,I723891,);
nor I_42435 (I724117,I724004,I1095355);
nand I_42436 (I724134,I724117,I1095352);
nor I_42437 (I724151,I723928,I724134);
DFFARX1 I_42438 (I724151,I2683,I723902,I723867,);
not I_42439 (I724182,I724134);
nand I_42440 (I723879,I723945,I724182);
DFFARX1 I_42441 (I724134,I2683,I723902,I724222,);
not I_42442 (I724230,I724222);
not I_42443 (I724247,I1095355);
not I_42444 (I724264,I1095346);
nor I_42445 (I724281,I724264,I1095334);
nor I_42446 (I723894,I724230,I724281);
nor I_42447 (I724312,I724264,I1095337);
and I_42448 (I724329,I724312,I1095361);
or I_42449 (I724346,I724329,I1095343);
DFFARX1 I_42450 (I724346,I2683,I723902,I724372,);
nor I_42451 (I723882,I724372,I723928);
not I_42452 (I724394,I724372);
and I_42453 (I724411,I724394,I723928);
nor I_42454 (I723876,I723953,I724411);
nand I_42455 (I724442,I724394,I724004);
nor I_42456 (I723870,I724264,I724442);
nand I_42457 (I723873,I724394,I724182);
nand I_42458 (I724487,I724004,I1095346);
nor I_42459 (I723885,I724247,I724487);
not I_42460 (I724548,I2690);
DFFARX1 I_42461 (I530090,I2683,I724548,I724574,);
DFFARX1 I_42462 (I530084,I2683,I724548,I724591,);
not I_42463 (I724599,I724591);
not I_42464 (I724616,I530099);
nor I_42465 (I724633,I724616,I530084);
not I_42466 (I724650,I530093);
nor I_42467 (I724667,I724633,I530102);
nor I_42468 (I724684,I724591,I724667);
DFFARX1 I_42469 (I724684,I2683,I724548,I724534,);
nor I_42470 (I724715,I530102,I530084);
nand I_42471 (I724732,I724715,I530099);
DFFARX1 I_42472 (I724732,I2683,I724548,I724537,);
nor I_42473 (I724763,I724650,I530102);
nand I_42474 (I724780,I724763,I530087);
nor I_42475 (I724797,I724574,I724780);
DFFARX1 I_42476 (I724797,I2683,I724548,I724513,);
not I_42477 (I724828,I724780);
nand I_42478 (I724525,I724591,I724828);
DFFARX1 I_42479 (I724780,I2683,I724548,I724868,);
not I_42480 (I724876,I724868);
not I_42481 (I724893,I530102);
not I_42482 (I724910,I530096);
nor I_42483 (I724927,I724910,I530093);
nor I_42484 (I724540,I724876,I724927);
nor I_42485 (I724958,I724910,I530105);
and I_42486 (I724975,I724958,I530108);
or I_42487 (I724992,I724975,I530087);
DFFARX1 I_42488 (I724992,I2683,I724548,I725018,);
nor I_42489 (I724528,I725018,I724574);
not I_42490 (I725040,I725018);
and I_42491 (I725057,I725040,I724574);
nor I_42492 (I724522,I724599,I725057);
nand I_42493 (I725088,I725040,I724650);
nor I_42494 (I724516,I724910,I725088);
nand I_42495 (I724519,I725040,I724828);
nand I_42496 (I725133,I724650,I530096);
nor I_42497 (I724531,I724893,I725133);
not I_42498 (I725194,I2690);
DFFARX1 I_42499 (I864628,I2683,I725194,I725220,);
DFFARX1 I_42500 (I864610,I2683,I725194,I725237,);
not I_42501 (I725245,I725237);
not I_42502 (I725262,I864619);
nor I_42503 (I725279,I725262,I864631);
not I_42504 (I725296,I864613);
nor I_42505 (I725313,I725279,I864622);
nor I_42506 (I725330,I725237,I725313);
DFFARX1 I_42507 (I725330,I2683,I725194,I725180,);
nor I_42508 (I725361,I864622,I864631);
nand I_42509 (I725378,I725361,I864619);
DFFARX1 I_42510 (I725378,I2683,I725194,I725183,);
nor I_42511 (I725409,I725296,I864622);
nand I_42512 (I725426,I725409,I864634);
nor I_42513 (I725443,I725220,I725426);
DFFARX1 I_42514 (I725443,I2683,I725194,I725159,);
not I_42515 (I725474,I725426);
nand I_42516 (I725171,I725237,I725474);
DFFARX1 I_42517 (I725426,I2683,I725194,I725514,);
not I_42518 (I725522,I725514);
not I_42519 (I725539,I864622);
not I_42520 (I725556,I864610);
nor I_42521 (I725573,I725556,I864613);
nor I_42522 (I725186,I725522,I725573);
nor I_42523 (I725604,I725556,I864616);
and I_42524 (I725621,I725604,I864625);
or I_42525 (I725638,I725621,I864613);
DFFARX1 I_42526 (I725638,I2683,I725194,I725664,);
nor I_42527 (I725174,I725664,I725220);
not I_42528 (I725686,I725664);
and I_42529 (I725703,I725686,I725220);
nor I_42530 (I725168,I725245,I725703);
nand I_42531 (I725734,I725686,I725296);
nor I_42532 (I725162,I725556,I725734);
nand I_42533 (I725165,I725686,I725474);
nand I_42534 (I725779,I725296,I864610);
nor I_42535 (I725177,I725539,I725779);
not I_42536 (I725840,I2690);
DFFARX1 I_42537 (I992051,I2683,I725840,I725866,);
DFFARX1 I_42538 (I992045,I2683,I725840,I725883,);
not I_42539 (I725891,I725883);
not I_42540 (I725908,I992054);
nor I_42541 (I725925,I725908,I992066);
not I_42542 (I725942,I992048);
nor I_42543 (I725959,I725925,I992045);
nor I_42544 (I725976,I725883,I725959);
DFFARX1 I_42545 (I725976,I2683,I725840,I725826,);
nor I_42546 (I726007,I992045,I992066);
nand I_42547 (I726024,I726007,I992054);
DFFARX1 I_42548 (I726024,I2683,I725840,I725829,);
nor I_42549 (I726055,I725942,I992045);
nand I_42550 (I726072,I726055,I992042);
nor I_42551 (I726089,I725866,I726072);
DFFARX1 I_42552 (I726089,I2683,I725840,I725805,);
not I_42553 (I726120,I726072);
nand I_42554 (I725817,I725883,I726120);
DFFARX1 I_42555 (I726072,I2683,I725840,I726160,);
not I_42556 (I726168,I726160);
not I_42557 (I726185,I992045);
not I_42558 (I726202,I992063);
nor I_42559 (I726219,I726202,I992048);
nor I_42560 (I725832,I726168,I726219);
nor I_42561 (I726250,I726202,I992057);
and I_42562 (I726267,I726250,I992042);
or I_42563 (I726284,I726267,I992060);
DFFARX1 I_42564 (I726284,I2683,I725840,I726310,);
nor I_42565 (I725820,I726310,I725866);
not I_42566 (I726332,I726310);
and I_42567 (I726349,I726332,I725866);
nor I_42568 (I725814,I725891,I726349);
nand I_42569 (I726380,I726332,I725942);
nor I_42570 (I725808,I726202,I726380);
nand I_42571 (I725811,I726332,I726120);
nand I_42572 (I726425,I725942,I992063);
nor I_42573 (I725823,I726185,I726425);
not I_42574 (I726486,I2690);
DFFARX1 I_42575 (I157501,I2683,I726486,I726512,);
DFFARX1 I_42576 (I157513,I2683,I726486,I726529,);
not I_42577 (I726537,I726529);
not I_42578 (I726554,I157519);
nor I_42579 (I726571,I726554,I157504);
not I_42580 (I726588,I157495);
nor I_42581 (I726605,I726571,I157516);
nor I_42582 (I726622,I726529,I726605);
DFFARX1 I_42583 (I726622,I2683,I726486,I726472,);
nor I_42584 (I726653,I157516,I157504);
nand I_42585 (I726670,I726653,I157519);
DFFARX1 I_42586 (I726670,I2683,I726486,I726475,);
nor I_42587 (I726701,I726588,I157516);
nand I_42588 (I726718,I726701,I157498);
nor I_42589 (I726735,I726512,I726718);
DFFARX1 I_42590 (I726735,I2683,I726486,I726451,);
not I_42591 (I726766,I726718);
nand I_42592 (I726463,I726529,I726766);
DFFARX1 I_42593 (I726718,I2683,I726486,I726806,);
not I_42594 (I726814,I726806);
not I_42595 (I726831,I157516);
not I_42596 (I726848,I157507);
nor I_42597 (I726865,I726848,I157495);
nor I_42598 (I726478,I726814,I726865);
nor I_42599 (I726896,I726848,I157510);
and I_42600 (I726913,I726896,I157498);
or I_42601 (I726930,I726913,I157495);
DFFARX1 I_42602 (I726930,I2683,I726486,I726956,);
nor I_42603 (I726466,I726956,I726512);
not I_42604 (I726978,I726956);
and I_42605 (I726995,I726978,I726512);
nor I_42606 (I726460,I726537,I726995);
nand I_42607 (I727026,I726978,I726588);
nor I_42608 (I726454,I726848,I727026);
nand I_42609 (I726457,I726978,I726766);
nand I_42610 (I727071,I726588,I157507);
nor I_42611 (I726469,I726831,I727071);
not I_42612 (I727132,I2690);
DFFARX1 I_42613 (I197366,I2683,I727132,I727158,);
DFFARX1 I_42614 (I197378,I2683,I727132,I727175,);
not I_42615 (I727183,I727175);
not I_42616 (I727200,I197384);
nor I_42617 (I727217,I727200,I197369);
not I_42618 (I727234,I197360);
nor I_42619 (I727251,I727217,I197381);
nor I_42620 (I727268,I727175,I727251);
DFFARX1 I_42621 (I727268,I2683,I727132,I727118,);
nor I_42622 (I727299,I197381,I197369);
nand I_42623 (I727316,I727299,I197384);
DFFARX1 I_42624 (I727316,I2683,I727132,I727121,);
nor I_42625 (I727347,I727234,I197381);
nand I_42626 (I727364,I727347,I197363);
nor I_42627 (I727381,I727158,I727364);
DFFARX1 I_42628 (I727381,I2683,I727132,I727097,);
not I_42629 (I727412,I727364);
nand I_42630 (I727109,I727175,I727412);
DFFARX1 I_42631 (I727364,I2683,I727132,I727452,);
not I_42632 (I727460,I727452);
not I_42633 (I727477,I197381);
not I_42634 (I727494,I197372);
nor I_42635 (I727511,I727494,I197360);
nor I_42636 (I727124,I727460,I727511);
nor I_42637 (I727542,I727494,I197375);
and I_42638 (I727559,I727542,I197363);
or I_42639 (I727576,I727559,I197360);
DFFARX1 I_42640 (I727576,I2683,I727132,I727602,);
nor I_42641 (I727112,I727602,I727158);
not I_42642 (I727624,I727602);
and I_42643 (I727641,I727624,I727158);
nor I_42644 (I727106,I727183,I727641);
nand I_42645 (I727672,I727624,I727234);
nor I_42646 (I727100,I727494,I727672);
nand I_42647 (I727103,I727624,I727412);
nand I_42648 (I727717,I727234,I197372);
nor I_42649 (I727115,I727477,I727717);
not I_42650 (I727778,I2690);
DFFARX1 I_42651 (I46927,I2683,I727778,I727804,);
DFFARX1 I_42652 (I46933,I2683,I727778,I727821,);
not I_42653 (I727829,I727821);
not I_42654 (I727846,I46951);
nor I_42655 (I727863,I727846,I46930);
not I_42656 (I727880,I46936);
nor I_42657 (I727897,I727863,I46942);
nor I_42658 (I727914,I727821,I727897);
DFFARX1 I_42659 (I727914,I2683,I727778,I727764,);
nor I_42660 (I727945,I46942,I46930);
nand I_42661 (I727962,I727945,I46951);
DFFARX1 I_42662 (I727962,I2683,I727778,I727767,);
nor I_42663 (I727993,I727880,I46942);
nand I_42664 (I728010,I727993,I46948);
nor I_42665 (I728027,I727804,I728010);
DFFARX1 I_42666 (I728027,I2683,I727778,I727743,);
not I_42667 (I728058,I728010);
nand I_42668 (I727755,I727821,I728058);
DFFARX1 I_42669 (I728010,I2683,I727778,I728098,);
not I_42670 (I728106,I728098);
not I_42671 (I728123,I46942);
not I_42672 (I728140,I46930);
nor I_42673 (I728157,I728140,I46936);
nor I_42674 (I727770,I728106,I728157);
nor I_42675 (I728188,I728140,I46939);
and I_42676 (I728205,I728188,I46927);
or I_42677 (I728222,I728205,I46945);
DFFARX1 I_42678 (I728222,I2683,I727778,I728248,);
nor I_42679 (I727758,I728248,I727804);
not I_42680 (I728270,I728248);
and I_42681 (I728287,I728270,I727804);
nor I_42682 (I727752,I727829,I728287);
nand I_42683 (I728318,I728270,I727880);
nor I_42684 (I727746,I728140,I728318);
nand I_42685 (I727749,I728270,I728058);
nand I_42686 (I728363,I727880,I46930);
nor I_42687 (I727761,I728123,I728363);
not I_42688 (I728424,I2690);
DFFARX1 I_42689 (I81709,I2683,I728424,I728450,);
DFFARX1 I_42690 (I81715,I2683,I728424,I728467,);
not I_42691 (I728475,I728467);
not I_42692 (I728492,I81733);
nor I_42693 (I728509,I728492,I81712);
not I_42694 (I728526,I81718);
nor I_42695 (I728543,I728509,I81724);
nor I_42696 (I728560,I728467,I728543);
DFFARX1 I_42697 (I728560,I2683,I728424,I728410,);
nor I_42698 (I728591,I81724,I81712);
nand I_42699 (I728608,I728591,I81733);
DFFARX1 I_42700 (I728608,I2683,I728424,I728413,);
nor I_42701 (I728639,I728526,I81724);
nand I_42702 (I728656,I728639,I81730);
nor I_42703 (I728673,I728450,I728656);
DFFARX1 I_42704 (I728673,I2683,I728424,I728389,);
not I_42705 (I728704,I728656);
nand I_42706 (I728401,I728467,I728704);
DFFARX1 I_42707 (I728656,I2683,I728424,I728744,);
not I_42708 (I728752,I728744);
not I_42709 (I728769,I81724);
not I_42710 (I728786,I81712);
nor I_42711 (I728803,I728786,I81718);
nor I_42712 (I728416,I728752,I728803);
nor I_42713 (I728834,I728786,I81721);
and I_42714 (I728851,I728834,I81709);
or I_42715 (I728868,I728851,I81727);
DFFARX1 I_42716 (I728868,I2683,I728424,I728894,);
nor I_42717 (I728404,I728894,I728450);
not I_42718 (I728916,I728894);
and I_42719 (I728933,I728916,I728450);
nor I_42720 (I728398,I728475,I728933);
nand I_42721 (I728964,I728916,I728526);
nor I_42722 (I728392,I728786,I728964);
nand I_42723 (I728395,I728916,I728704);
nand I_42724 (I729009,I728526,I81712);
nor I_42725 (I728407,I728769,I729009);
not I_42726 (I729070,I2690);
DFFARX1 I_42727 (I132511,I2683,I729070,I729096,);
DFFARX1 I_42728 (I132523,I2683,I729070,I729113,);
not I_42729 (I729121,I729113);
not I_42730 (I729138,I132529);
nor I_42731 (I729155,I729138,I132514);
not I_42732 (I729172,I132505);
nor I_42733 (I729189,I729155,I132526);
nor I_42734 (I729206,I729113,I729189);
DFFARX1 I_42735 (I729206,I2683,I729070,I729056,);
nor I_42736 (I729237,I132526,I132514);
nand I_42737 (I729254,I729237,I132529);
DFFARX1 I_42738 (I729254,I2683,I729070,I729059,);
nor I_42739 (I729285,I729172,I132526);
nand I_42740 (I729302,I729285,I132508);
nor I_42741 (I729319,I729096,I729302);
DFFARX1 I_42742 (I729319,I2683,I729070,I729035,);
not I_42743 (I729350,I729302);
nand I_42744 (I729047,I729113,I729350);
DFFARX1 I_42745 (I729302,I2683,I729070,I729390,);
not I_42746 (I729398,I729390);
not I_42747 (I729415,I132526);
not I_42748 (I729432,I132517);
nor I_42749 (I729449,I729432,I132505);
nor I_42750 (I729062,I729398,I729449);
nor I_42751 (I729480,I729432,I132520);
and I_42752 (I729497,I729480,I132508);
or I_42753 (I729514,I729497,I132505);
DFFARX1 I_42754 (I729514,I2683,I729070,I729540,);
nor I_42755 (I729050,I729540,I729096);
not I_42756 (I729562,I729540);
and I_42757 (I729579,I729562,I729096);
nor I_42758 (I729044,I729121,I729579);
nand I_42759 (I729610,I729562,I729172);
nor I_42760 (I729038,I729432,I729610);
nand I_42761 (I729041,I729562,I729350);
nand I_42762 (I729655,I729172,I132517);
nor I_42763 (I729053,I729415,I729655);
not I_42764 (I729716,I2690);
DFFARX1 I_42765 (I412770,I2683,I729716,I729742,);
DFFARX1 I_42766 (I412782,I2683,I729716,I729759,);
not I_42767 (I729767,I729759);
not I_42768 (I729784,I412767);
nor I_42769 (I729801,I729784,I412785);
not I_42770 (I729818,I412791);
nor I_42771 (I729835,I729801,I412773);
nor I_42772 (I729852,I729759,I729835);
DFFARX1 I_42773 (I729852,I2683,I729716,I729702,);
nor I_42774 (I729883,I412773,I412785);
nand I_42775 (I729900,I729883,I412767);
DFFARX1 I_42776 (I729900,I2683,I729716,I729705,);
nor I_42777 (I729931,I729818,I412773);
nand I_42778 (I729948,I729931,I412776);
nor I_42779 (I729965,I729742,I729948);
DFFARX1 I_42780 (I729965,I2683,I729716,I729681,);
not I_42781 (I729996,I729948);
nand I_42782 (I729693,I729759,I729996);
DFFARX1 I_42783 (I729948,I2683,I729716,I730036,);
not I_42784 (I730044,I730036);
not I_42785 (I730061,I412773);
not I_42786 (I730078,I412779);
nor I_42787 (I730095,I730078,I412791);
nor I_42788 (I729708,I730044,I730095);
nor I_42789 (I730126,I730078,I412788);
and I_42790 (I730143,I730126,I412767);
or I_42791 (I730160,I730143,I412770);
DFFARX1 I_42792 (I730160,I2683,I729716,I730186,);
nor I_42793 (I729696,I730186,I729742);
not I_42794 (I730208,I730186);
and I_42795 (I730225,I730208,I729742);
nor I_42796 (I729690,I729767,I730225);
nand I_42797 (I730256,I730208,I729818);
nor I_42798 (I729684,I730078,I730256);
nand I_42799 (I729687,I730208,I729996);
nand I_42800 (I730301,I729818,I412779);
nor I_42801 (I729699,I730061,I730301);
not I_42802 (I730362,I2690);
DFFARX1 I_42803 (I221126,I2683,I730362,I730388,);
DFFARX1 I_42804 (I221132,I2683,I730362,I730405,);
not I_42805 (I730413,I730405);
not I_42806 (I730430,I221153);
nor I_42807 (I730447,I730430,I221141);
not I_42808 (I730464,I221150);
nor I_42809 (I730481,I730447,I221135);
nor I_42810 (I730498,I730405,I730481);
DFFARX1 I_42811 (I730498,I2683,I730362,I730348,);
nor I_42812 (I730529,I221135,I221141);
nand I_42813 (I730546,I730529,I221153);
DFFARX1 I_42814 (I730546,I2683,I730362,I730351,);
nor I_42815 (I730577,I730464,I221135);
nand I_42816 (I730594,I730577,I221126);
nor I_42817 (I730611,I730388,I730594);
DFFARX1 I_42818 (I730611,I2683,I730362,I730327,);
not I_42819 (I730642,I730594);
nand I_42820 (I730339,I730405,I730642);
DFFARX1 I_42821 (I730594,I2683,I730362,I730682,);
not I_42822 (I730690,I730682);
not I_42823 (I730707,I221135);
not I_42824 (I730724,I221138);
nor I_42825 (I730741,I730724,I221150);
nor I_42826 (I730354,I730690,I730741);
nor I_42827 (I730772,I730724,I221147);
and I_42828 (I730789,I730772,I221129);
or I_42829 (I730806,I730789,I221144);
DFFARX1 I_42830 (I730806,I2683,I730362,I730832,);
nor I_42831 (I730342,I730832,I730388);
not I_42832 (I730854,I730832);
and I_42833 (I730871,I730854,I730388);
nor I_42834 (I730336,I730413,I730871);
nand I_42835 (I730902,I730854,I730464);
nor I_42836 (I730330,I730724,I730902);
nand I_42837 (I730333,I730854,I730642);
nand I_42838 (I730947,I730464,I221138);
nor I_42839 (I730345,I730707,I730947);
not I_42840 (I731008,I2690);
DFFARX1 I_42841 (I317624,I2683,I731008,I731034,);
DFFARX1 I_42842 (I317621,I2683,I731008,I731051,);
not I_42843 (I731059,I731051);
not I_42844 (I731076,I317636);
nor I_42845 (I731093,I731076,I317639);
not I_42846 (I731110,I317627);
nor I_42847 (I731127,I731093,I317633);
nor I_42848 (I731144,I731051,I731127);
DFFARX1 I_42849 (I731144,I2683,I731008,I730994,);
nor I_42850 (I731175,I317633,I317639);
nand I_42851 (I731192,I731175,I317636);
DFFARX1 I_42852 (I731192,I2683,I731008,I730997,);
nor I_42853 (I731223,I731110,I317633);
nand I_42854 (I731240,I731223,I317645);
nor I_42855 (I731257,I731034,I731240);
DFFARX1 I_42856 (I731257,I2683,I731008,I730973,);
not I_42857 (I731288,I731240);
nand I_42858 (I730985,I731051,I731288);
DFFARX1 I_42859 (I731240,I2683,I731008,I731328,);
not I_42860 (I731336,I731328);
not I_42861 (I731353,I317633);
not I_42862 (I731370,I317618);
nor I_42863 (I731387,I731370,I317627);
nor I_42864 (I731000,I731336,I731387);
nor I_42865 (I731418,I731370,I317630);
and I_42866 (I731435,I731418,I317618);
or I_42867 (I731452,I731435,I317642);
DFFARX1 I_42868 (I731452,I2683,I731008,I731478,);
nor I_42869 (I730988,I731478,I731034);
not I_42870 (I731500,I731478);
and I_42871 (I731517,I731500,I731034);
nor I_42872 (I730982,I731059,I731517);
nand I_42873 (I731548,I731500,I731110);
nor I_42874 (I730976,I731370,I731548);
nand I_42875 (I730979,I731500,I731288);
nand I_42876 (I731593,I731110,I317618);
nor I_42877 (I730991,I731353,I731593);
not I_42878 (I731654,I2690);
DFFARX1 I_42879 (I843820,I2683,I731654,I731680,);
DFFARX1 I_42880 (I843802,I2683,I731654,I731697,);
not I_42881 (I731705,I731697);
not I_42882 (I731722,I843811);
nor I_42883 (I731739,I731722,I843823);
not I_42884 (I731756,I843805);
nor I_42885 (I731773,I731739,I843814);
nor I_42886 (I731790,I731697,I731773);
DFFARX1 I_42887 (I731790,I2683,I731654,I731640,);
nor I_42888 (I731821,I843814,I843823);
nand I_42889 (I731838,I731821,I843811);
DFFARX1 I_42890 (I731838,I2683,I731654,I731643,);
nor I_42891 (I731869,I731756,I843814);
nand I_42892 (I731886,I731869,I843826);
nor I_42893 (I731903,I731680,I731886);
DFFARX1 I_42894 (I731903,I2683,I731654,I731619,);
not I_42895 (I731934,I731886);
nand I_42896 (I731631,I731697,I731934);
DFFARX1 I_42897 (I731886,I2683,I731654,I731974,);
not I_42898 (I731982,I731974);
not I_42899 (I731999,I843814);
not I_42900 (I732016,I843802);
nor I_42901 (I732033,I732016,I843805);
nor I_42902 (I731646,I731982,I732033);
nor I_42903 (I732064,I732016,I843808);
and I_42904 (I732081,I732064,I843817);
or I_42905 (I732098,I732081,I843805);
DFFARX1 I_42906 (I732098,I2683,I731654,I732124,);
nor I_42907 (I731634,I732124,I731680);
not I_42908 (I732146,I732124);
and I_42909 (I732163,I732146,I731680);
nor I_42910 (I731628,I731705,I732163);
nand I_42911 (I732194,I732146,I731756);
nor I_42912 (I731622,I732016,I732194);
nand I_42913 (I731625,I732146,I731934);
nand I_42914 (I732239,I731756,I843802);
nor I_42915 (I731637,I731999,I732239);
not I_42916 (I732300,I2690);
DFFARX1 I_42917 (I591358,I2683,I732300,I732326,);
DFFARX1 I_42918 (I591352,I2683,I732300,I732343,);
not I_42919 (I732351,I732343);
not I_42920 (I732368,I591367);
nor I_42921 (I732385,I732368,I591352);
not I_42922 (I732402,I591361);
nor I_42923 (I732419,I732385,I591370);
nor I_42924 (I732436,I732343,I732419);
DFFARX1 I_42925 (I732436,I2683,I732300,I732286,);
nor I_42926 (I732467,I591370,I591352);
nand I_42927 (I732484,I732467,I591367);
DFFARX1 I_42928 (I732484,I2683,I732300,I732289,);
nor I_42929 (I732515,I732402,I591370);
nand I_42930 (I732532,I732515,I591355);
nor I_42931 (I732549,I732326,I732532);
DFFARX1 I_42932 (I732549,I2683,I732300,I732265,);
not I_42933 (I732580,I732532);
nand I_42934 (I732277,I732343,I732580);
DFFARX1 I_42935 (I732532,I2683,I732300,I732620,);
not I_42936 (I732628,I732620);
not I_42937 (I732645,I591370);
not I_42938 (I732662,I591364);
nor I_42939 (I732679,I732662,I591361);
nor I_42940 (I732292,I732628,I732679);
nor I_42941 (I732710,I732662,I591373);
and I_42942 (I732727,I732710,I591376);
or I_42943 (I732744,I732727,I591355);
DFFARX1 I_42944 (I732744,I2683,I732300,I732770,);
nor I_42945 (I732280,I732770,I732326);
not I_42946 (I732792,I732770);
and I_42947 (I732809,I732792,I732326);
nor I_42948 (I732274,I732351,I732809);
nand I_42949 (I732840,I732792,I732402);
nor I_42950 (I732268,I732662,I732840);
nand I_42951 (I732271,I732792,I732580);
nand I_42952 (I732885,I732402,I591364);
nor I_42953 (I732283,I732645,I732885);
not I_42954 (I732946,I2690);
DFFARX1 I_42955 (I298595,I2683,I732946,I732972,);
DFFARX1 I_42956 (I298601,I2683,I732946,I732989,);
not I_42957 (I732997,I732989);
not I_42958 (I733014,I298622);
nor I_42959 (I733031,I733014,I298610);
not I_42960 (I733048,I298619);
nor I_42961 (I733065,I733031,I298604);
nor I_42962 (I733082,I732989,I733065);
DFFARX1 I_42963 (I733082,I2683,I732946,I732932,);
nor I_42964 (I733113,I298604,I298610);
nand I_42965 (I733130,I733113,I298622);
DFFARX1 I_42966 (I733130,I2683,I732946,I732935,);
nor I_42967 (I733161,I733048,I298604);
nand I_42968 (I733178,I733161,I298595);
nor I_42969 (I733195,I732972,I733178);
DFFARX1 I_42970 (I733195,I2683,I732946,I732911,);
not I_42971 (I733226,I733178);
nand I_42972 (I732923,I732989,I733226);
DFFARX1 I_42973 (I733178,I2683,I732946,I733266,);
not I_42974 (I733274,I733266);
not I_42975 (I733291,I298604);
not I_42976 (I733308,I298607);
nor I_42977 (I733325,I733308,I298619);
nor I_42978 (I732938,I733274,I733325);
nor I_42979 (I733356,I733308,I298616);
and I_42980 (I733373,I733356,I298598);
or I_42981 (I733390,I733373,I298613);
DFFARX1 I_42982 (I733390,I2683,I732946,I733416,);
nor I_42983 (I732926,I733416,I732972);
not I_42984 (I733438,I733416);
and I_42985 (I733455,I733438,I732972);
nor I_42986 (I732920,I732997,I733455);
nand I_42987 (I733486,I733438,I733048);
nor I_42988 (I732914,I733308,I733486);
nand I_42989 (I732917,I733438,I733226);
nand I_42990 (I733531,I733048,I298607);
nor I_42991 (I732929,I733291,I733531);
not I_42992 (I733592,I2690);
DFFARX1 I_42993 (I973360,I2683,I733592,I733618,);
DFFARX1 I_42994 (I973366,I2683,I733592,I733635,);
not I_42995 (I733643,I733635);
not I_42996 (I733660,I973363);
nor I_42997 (I733677,I733660,I973342);
not I_42998 (I733694,I973345);
nor I_42999 (I733711,I733677,I973351);
nor I_43000 (I733728,I733635,I733711);
DFFARX1 I_43001 (I733728,I2683,I733592,I733578,);
nor I_43002 (I733759,I973351,I973342);
nand I_43003 (I733776,I733759,I973363);
DFFARX1 I_43004 (I733776,I2683,I733592,I733581,);
nor I_43005 (I733807,I733694,I973351);
nand I_43006 (I733824,I733807,I973345);
nor I_43007 (I733841,I733618,I733824);
DFFARX1 I_43008 (I733841,I2683,I733592,I733557,);
not I_43009 (I733872,I733824);
nand I_43010 (I733569,I733635,I733872);
DFFARX1 I_43011 (I733824,I2683,I733592,I733912,);
not I_43012 (I733920,I733912);
not I_43013 (I733937,I973351);
not I_43014 (I733954,I973354);
nor I_43015 (I733971,I733954,I973345);
nor I_43016 (I733584,I733920,I733971);
nor I_43017 (I734002,I733954,I973342);
and I_43018 (I734019,I734002,I973348);
or I_43019 (I734036,I734019,I973357);
DFFARX1 I_43020 (I734036,I2683,I733592,I734062,);
nor I_43021 (I733572,I734062,I733618);
not I_43022 (I734084,I734062);
and I_43023 (I734101,I734084,I733618);
nor I_43024 (I733566,I733643,I734101);
nand I_43025 (I734132,I734084,I733694);
nor I_43026 (I733560,I733954,I734132);
nand I_43027 (I733563,I734084,I733872);
nand I_43028 (I734177,I733694,I973354);
nor I_43029 (I733575,I733937,I734177);
not I_43030 (I734238,I2690);
DFFARX1 I_43031 (I539916,I2683,I734238,I734264,);
DFFARX1 I_43032 (I539910,I2683,I734238,I734281,);
not I_43033 (I734289,I734281);
not I_43034 (I734306,I539925);
nor I_43035 (I734323,I734306,I539910);
not I_43036 (I734340,I539919);
nor I_43037 (I734357,I734323,I539928);
nor I_43038 (I734374,I734281,I734357);
DFFARX1 I_43039 (I734374,I2683,I734238,I734224,);
nor I_43040 (I734405,I539928,I539910);
nand I_43041 (I734422,I734405,I539925);
DFFARX1 I_43042 (I734422,I2683,I734238,I734227,);
nor I_43043 (I734453,I734340,I539928);
nand I_43044 (I734470,I734453,I539913);
nor I_43045 (I734487,I734264,I734470);
DFFARX1 I_43046 (I734487,I2683,I734238,I734203,);
not I_43047 (I734518,I734470);
nand I_43048 (I734215,I734281,I734518);
DFFARX1 I_43049 (I734470,I2683,I734238,I734558,);
not I_43050 (I734566,I734558);
not I_43051 (I734583,I539928);
not I_43052 (I734600,I539922);
nor I_43053 (I734617,I734600,I539919);
nor I_43054 (I734230,I734566,I734617);
nor I_43055 (I734648,I734600,I539931);
and I_43056 (I734665,I734648,I539934);
or I_43057 (I734682,I734665,I539913);
DFFARX1 I_43058 (I734682,I2683,I734238,I734708,);
nor I_43059 (I734218,I734708,I734264);
not I_43060 (I734730,I734708);
and I_43061 (I734747,I734730,I734264);
nor I_43062 (I734212,I734289,I734747);
nand I_43063 (I734778,I734730,I734340);
nor I_43064 (I734206,I734600,I734778);
nand I_43065 (I734209,I734730,I734518);
nand I_43066 (I734823,I734340,I539922);
nor I_43067 (I734221,I734583,I734823);
not I_43068 (I734884,I2690);
DFFARX1 I_43069 (I415150,I2683,I734884,I734910,);
DFFARX1 I_43070 (I415162,I2683,I734884,I734927,);
not I_43071 (I734935,I734927);
not I_43072 (I734952,I415147);
nor I_43073 (I734969,I734952,I415165);
not I_43074 (I734986,I415171);
nor I_43075 (I735003,I734969,I415153);
nor I_43076 (I735020,I734927,I735003);
DFFARX1 I_43077 (I735020,I2683,I734884,I734870,);
nor I_43078 (I735051,I415153,I415165);
nand I_43079 (I735068,I735051,I415147);
DFFARX1 I_43080 (I735068,I2683,I734884,I734873,);
nor I_43081 (I735099,I734986,I415153);
nand I_43082 (I735116,I735099,I415156);
nor I_43083 (I735133,I734910,I735116);
DFFARX1 I_43084 (I735133,I2683,I734884,I734849,);
not I_43085 (I735164,I735116);
nand I_43086 (I734861,I734927,I735164);
DFFARX1 I_43087 (I735116,I2683,I734884,I735204,);
not I_43088 (I735212,I735204);
not I_43089 (I735229,I415153);
not I_43090 (I735246,I415159);
nor I_43091 (I735263,I735246,I415171);
nor I_43092 (I734876,I735212,I735263);
nor I_43093 (I735294,I735246,I415168);
and I_43094 (I735311,I735294,I415147);
or I_43095 (I735328,I735311,I415150);
DFFARX1 I_43096 (I735328,I2683,I734884,I735354,);
nor I_43097 (I734864,I735354,I734910);
not I_43098 (I735376,I735354);
and I_43099 (I735393,I735376,I734910);
nor I_43100 (I734858,I734935,I735393);
nand I_43101 (I735424,I735376,I734986);
nor I_43102 (I734852,I735246,I735424);
nand I_43103 (I734855,I735376,I735164);
nand I_43104 (I735469,I734986,I415159);
nor I_43105 (I734867,I735229,I735469);
not I_43106 (I735530,I2690);
DFFARX1 I_43107 (I240098,I2683,I735530,I735556,);
DFFARX1 I_43108 (I240104,I2683,I735530,I735573,);
not I_43109 (I735581,I735573);
not I_43110 (I735598,I240125);
nor I_43111 (I735615,I735598,I240113);
not I_43112 (I735632,I240122);
nor I_43113 (I735649,I735615,I240107);
nor I_43114 (I735666,I735573,I735649);
DFFARX1 I_43115 (I735666,I2683,I735530,I735516,);
nor I_43116 (I735697,I240107,I240113);
nand I_43117 (I735714,I735697,I240125);
DFFARX1 I_43118 (I735714,I2683,I735530,I735519,);
nor I_43119 (I735745,I735632,I240107);
nand I_43120 (I735762,I735745,I240098);
nor I_43121 (I735779,I735556,I735762);
DFFARX1 I_43122 (I735779,I2683,I735530,I735495,);
not I_43123 (I735810,I735762);
nand I_43124 (I735507,I735573,I735810);
DFFARX1 I_43125 (I735762,I2683,I735530,I735850,);
not I_43126 (I735858,I735850);
not I_43127 (I735875,I240107);
not I_43128 (I735892,I240110);
nor I_43129 (I735909,I735892,I240122);
nor I_43130 (I735522,I735858,I735909);
nor I_43131 (I735940,I735892,I240119);
and I_43132 (I735957,I735940,I240101);
or I_43133 (I735974,I735957,I240116);
DFFARX1 I_43134 (I735974,I2683,I735530,I736000,);
nor I_43135 (I735510,I736000,I735556);
not I_43136 (I736022,I736000);
and I_43137 (I736039,I736022,I735556);
nor I_43138 (I735504,I735581,I736039);
nand I_43139 (I736070,I736022,I735632);
nor I_43140 (I735498,I735892,I736070);
nand I_43141 (I735501,I736022,I735810);
nand I_43142 (I736115,I735632,I240110);
nor I_43143 (I735513,I735875,I736115);
not I_43144 (I736176,I2690);
DFFARX1 I_43145 (I1054874,I2683,I736176,I736202,);
DFFARX1 I_43146 (I1054898,I2683,I736176,I736219,);
not I_43147 (I736227,I736219);
not I_43148 (I736244,I1054880);
nor I_43149 (I736261,I736244,I1054889);
not I_43150 (I736278,I1054874);
nor I_43151 (I736295,I736261,I1054895);
nor I_43152 (I736312,I736219,I736295);
DFFARX1 I_43153 (I736312,I2683,I736176,I736162,);
nor I_43154 (I736343,I1054895,I1054889);
nand I_43155 (I736360,I736343,I1054880);
DFFARX1 I_43156 (I736360,I2683,I736176,I736165,);
nor I_43157 (I736391,I736278,I1054895);
nand I_43158 (I736408,I736391,I1054892);
nor I_43159 (I736425,I736202,I736408);
DFFARX1 I_43160 (I736425,I2683,I736176,I736141,);
not I_43161 (I736456,I736408);
nand I_43162 (I736153,I736219,I736456);
DFFARX1 I_43163 (I736408,I2683,I736176,I736496,);
not I_43164 (I736504,I736496);
not I_43165 (I736521,I1054895);
not I_43166 (I736538,I1054886);
nor I_43167 (I736555,I736538,I1054874);
nor I_43168 (I736168,I736504,I736555);
nor I_43169 (I736586,I736538,I1054877);
and I_43170 (I736603,I736586,I1054901);
or I_43171 (I736620,I736603,I1054883);
DFFARX1 I_43172 (I736620,I2683,I736176,I736646,);
nor I_43173 (I736156,I736646,I736202);
not I_43174 (I736668,I736646);
and I_43175 (I736685,I736668,I736202);
nor I_43176 (I736150,I736227,I736685);
nand I_43177 (I736716,I736668,I736278);
nor I_43178 (I736144,I736538,I736716);
nand I_43179 (I736147,I736668,I736456);
nand I_43180 (I736761,I736278,I1054886);
nor I_43181 (I736159,I736521,I736761);
not I_43182 (I736822,I2690);
DFFARX1 I_43183 (I622264,I2683,I736822,I736848,);
DFFARX1 I_43184 (I622261,I2683,I736822,I736865,);
not I_43185 (I736873,I736865);
not I_43186 (I736890,I622261);
nor I_43187 (I736907,I736890,I622264);
not I_43188 (I736924,I622276);
nor I_43189 (I736941,I736907,I622270);
nor I_43190 (I736958,I736865,I736941);
DFFARX1 I_43191 (I736958,I2683,I736822,I736808,);
nor I_43192 (I736989,I622270,I622264);
nand I_43193 (I737006,I736989,I622261);
DFFARX1 I_43194 (I737006,I2683,I736822,I736811,);
nor I_43195 (I737037,I736924,I622270);
nand I_43196 (I737054,I737037,I622258);
nor I_43197 (I737071,I736848,I737054);
DFFARX1 I_43198 (I737071,I2683,I736822,I736787,);
not I_43199 (I737102,I737054);
nand I_43200 (I736799,I736865,I737102);
DFFARX1 I_43201 (I737054,I2683,I736822,I737142,);
not I_43202 (I737150,I737142);
not I_43203 (I737167,I622270);
not I_43204 (I737184,I622267);
nor I_43205 (I737201,I737184,I622276);
nor I_43206 (I736814,I737150,I737201);
nor I_43207 (I737232,I737184,I622273);
and I_43208 (I737249,I737232,I622279);
or I_43209 (I737266,I737249,I622258);
DFFARX1 I_43210 (I737266,I2683,I736822,I737292,);
nor I_43211 (I736802,I737292,I736848);
not I_43212 (I737314,I737292);
and I_43213 (I737331,I737314,I736848);
nor I_43214 (I736796,I736873,I737331);
nand I_43215 (I737362,I737314,I736924);
nor I_43216 (I736790,I737184,I737362);
nand I_43217 (I736793,I737314,I737102);
nand I_43218 (I737407,I736924,I622267);
nor I_43219 (I736805,I737167,I737407);
not I_43220 (I737468,I2690);
DFFARX1 I_43221 (I91195,I2683,I737468,I737494,);
DFFARX1 I_43222 (I91201,I2683,I737468,I737511,);
not I_43223 (I737519,I737511);
not I_43224 (I737536,I91219);
nor I_43225 (I737553,I737536,I91198);
not I_43226 (I737570,I91204);
nor I_43227 (I737587,I737553,I91210);
nor I_43228 (I737604,I737511,I737587);
DFFARX1 I_43229 (I737604,I2683,I737468,I737454,);
nor I_43230 (I737635,I91210,I91198);
nand I_43231 (I737652,I737635,I91219);
DFFARX1 I_43232 (I737652,I2683,I737468,I737457,);
nor I_43233 (I737683,I737570,I91210);
nand I_43234 (I737700,I737683,I91216);
nor I_43235 (I737717,I737494,I737700);
DFFARX1 I_43236 (I737717,I2683,I737468,I737433,);
not I_43237 (I737748,I737700);
nand I_43238 (I737445,I737511,I737748);
DFFARX1 I_43239 (I737700,I2683,I737468,I737788,);
not I_43240 (I737796,I737788);
not I_43241 (I737813,I91210);
not I_43242 (I737830,I91198);
nor I_43243 (I737847,I737830,I91204);
nor I_43244 (I737460,I737796,I737847);
nor I_43245 (I737878,I737830,I91207);
and I_43246 (I737895,I737878,I91195);
or I_43247 (I737912,I737895,I91213);
DFFARX1 I_43248 (I737912,I2683,I737468,I737938,);
nor I_43249 (I737448,I737938,I737494);
not I_43250 (I737960,I737938);
and I_43251 (I737977,I737960,I737494);
nor I_43252 (I737442,I737519,I737977);
nand I_43253 (I738008,I737960,I737570);
nor I_43254 (I737436,I737830,I738008);
nand I_43255 (I737439,I737960,I737748);
nand I_43256 (I738053,I737570,I91198);
nor I_43257 (I737451,I737813,I738053);
not I_43258 (I738114,I2690);
DFFARX1 I_43259 (I803512,I2683,I738114,I738140,);
DFFARX1 I_43260 (I803515,I2683,I738114,I738157,);
not I_43261 (I738165,I738157);
not I_43262 (I738182,I803512);
nor I_43263 (I738199,I738182,I803524);
not I_43264 (I738216,I803533);
nor I_43265 (I738233,I738199,I803521);
nor I_43266 (I738250,I738157,I738233);
DFFARX1 I_43267 (I738250,I2683,I738114,I738100,);
nor I_43268 (I738281,I803521,I803524);
nand I_43269 (I738298,I738281,I803512);
DFFARX1 I_43270 (I738298,I2683,I738114,I738103,);
nor I_43271 (I738329,I738216,I803521);
nand I_43272 (I738346,I738329,I803527);
nor I_43273 (I738363,I738140,I738346);
DFFARX1 I_43274 (I738363,I2683,I738114,I738079,);
not I_43275 (I738394,I738346);
nand I_43276 (I738091,I738157,I738394);
DFFARX1 I_43277 (I738346,I2683,I738114,I738434,);
not I_43278 (I738442,I738434);
not I_43279 (I738459,I803521);
not I_43280 (I738476,I803518);
nor I_43281 (I738493,I738476,I803533);
nor I_43282 (I738106,I738442,I738493);
nor I_43283 (I738524,I738476,I803530);
and I_43284 (I738541,I738524,I803518);
or I_43285 (I738558,I738541,I803515);
DFFARX1 I_43286 (I738558,I2683,I738114,I738584,);
nor I_43287 (I738094,I738584,I738140);
not I_43288 (I738606,I738584);
and I_43289 (I738623,I738606,I738140);
nor I_43290 (I738088,I738165,I738623);
nand I_43291 (I738654,I738606,I738216);
nor I_43292 (I738082,I738476,I738654);
nand I_43293 (I738085,I738606,I738394);
nand I_43294 (I738699,I738216,I803518);
nor I_43295 (I738097,I738459,I738699);
not I_43296 (I738760,I2690);
DFFARX1 I_43297 (I645979,I2683,I738760,I738786,);
DFFARX1 I_43298 (I645976,I2683,I738760,I738803,);
not I_43299 (I738811,I738803);
not I_43300 (I738828,I645976);
nor I_43301 (I738845,I738828,I645979);
not I_43302 (I738862,I645991);
nor I_43303 (I738879,I738845,I645985);
nor I_43304 (I738896,I738803,I738879);
DFFARX1 I_43305 (I738896,I2683,I738760,I738746,);
nor I_43306 (I738927,I645985,I645979);
nand I_43307 (I738944,I738927,I645976);
DFFARX1 I_43308 (I738944,I2683,I738760,I738749,);
nor I_43309 (I738975,I738862,I645985);
nand I_43310 (I738992,I738975,I645973);
nor I_43311 (I739009,I738786,I738992);
DFFARX1 I_43312 (I739009,I2683,I738760,I738725,);
not I_43313 (I739040,I738992);
nand I_43314 (I738737,I738803,I739040);
DFFARX1 I_43315 (I738992,I2683,I738760,I739080,);
not I_43316 (I739088,I739080);
not I_43317 (I739105,I645985);
not I_43318 (I739122,I645982);
nor I_43319 (I739139,I739122,I645991);
nor I_43320 (I738752,I739088,I739139);
nor I_43321 (I739170,I739122,I645988);
and I_43322 (I739187,I739170,I645994);
or I_43323 (I739204,I739187,I645973);
DFFARX1 I_43324 (I739204,I2683,I738760,I739230,);
nor I_43325 (I738740,I739230,I738786);
not I_43326 (I739252,I739230);
and I_43327 (I739269,I739252,I738786);
nor I_43328 (I738734,I738811,I739269);
nand I_43329 (I739300,I739252,I738862);
nor I_43330 (I738728,I739122,I739300);
nand I_43331 (I738731,I739252,I739040);
nand I_43332 (I739345,I738862,I645982);
nor I_43333 (I738743,I739105,I739345);
not I_43334 (I739406,I2690);
DFFARX1 I_43335 (I70642,I2683,I739406,I739432,);
DFFARX1 I_43336 (I70648,I2683,I739406,I739449,);
not I_43337 (I739457,I739449);
not I_43338 (I739474,I70666);
nor I_43339 (I739491,I739474,I70645);
not I_43340 (I739508,I70651);
nor I_43341 (I739525,I739491,I70657);
nor I_43342 (I739542,I739449,I739525);
DFFARX1 I_43343 (I739542,I2683,I739406,I739392,);
nor I_43344 (I739573,I70657,I70645);
nand I_43345 (I739590,I739573,I70666);
DFFARX1 I_43346 (I739590,I2683,I739406,I739395,);
nor I_43347 (I739621,I739508,I70657);
nand I_43348 (I739638,I739621,I70663);
nor I_43349 (I739655,I739432,I739638);
DFFARX1 I_43350 (I739655,I2683,I739406,I739371,);
not I_43351 (I739686,I739638);
nand I_43352 (I739383,I739449,I739686);
DFFARX1 I_43353 (I739638,I2683,I739406,I739726,);
not I_43354 (I739734,I739726);
not I_43355 (I739751,I70657);
not I_43356 (I739768,I70645);
nor I_43357 (I739785,I739768,I70651);
nor I_43358 (I739398,I739734,I739785);
nor I_43359 (I739816,I739768,I70654);
and I_43360 (I739833,I739816,I70642);
or I_43361 (I739850,I739833,I70660);
DFFARX1 I_43362 (I739850,I2683,I739406,I739876,);
nor I_43363 (I739386,I739876,I739432);
not I_43364 (I739898,I739876);
and I_43365 (I739915,I739898,I739432);
nor I_43366 (I739380,I739457,I739915);
nand I_43367 (I739946,I739898,I739508);
nor I_43368 (I739374,I739768,I739946);
nand I_43369 (I739377,I739898,I739686);
nand I_43370 (I739991,I739508,I70645);
nor I_43371 (I739389,I739751,I739991);
not I_43372 (I740052,I2690);
DFFARX1 I_43373 (I288055,I2683,I740052,I740078,);
DFFARX1 I_43374 (I288061,I2683,I740052,I740095,);
not I_43375 (I740103,I740095);
not I_43376 (I740120,I288082);
nor I_43377 (I740137,I740120,I288070);
not I_43378 (I740154,I288079);
nor I_43379 (I740171,I740137,I288064);
nor I_43380 (I740188,I740095,I740171);
DFFARX1 I_43381 (I740188,I2683,I740052,I740038,);
nor I_43382 (I740219,I288064,I288070);
nand I_43383 (I740236,I740219,I288082);
DFFARX1 I_43384 (I740236,I2683,I740052,I740041,);
nor I_43385 (I740267,I740154,I288064);
nand I_43386 (I740284,I740267,I288055);
nor I_43387 (I740301,I740078,I740284);
DFFARX1 I_43388 (I740301,I2683,I740052,I740017,);
not I_43389 (I740332,I740284);
nand I_43390 (I740029,I740095,I740332);
DFFARX1 I_43391 (I740284,I2683,I740052,I740372,);
not I_43392 (I740380,I740372);
not I_43393 (I740397,I288064);
not I_43394 (I740414,I288067);
nor I_43395 (I740431,I740414,I288079);
nor I_43396 (I740044,I740380,I740431);
nor I_43397 (I740462,I740414,I288076);
and I_43398 (I740479,I740462,I288058);
or I_43399 (I740496,I740479,I288073);
DFFARX1 I_43400 (I740496,I2683,I740052,I740522,);
nor I_43401 (I740032,I740522,I740078);
not I_43402 (I740544,I740522);
and I_43403 (I740561,I740544,I740078);
nor I_43404 (I740026,I740103,I740561);
nand I_43405 (I740592,I740544,I740154);
nor I_43406 (I740020,I740414,I740592);
nand I_43407 (I740023,I740544,I740332);
nand I_43408 (I740637,I740154,I288067);
nor I_43409 (I740035,I740397,I740637);
not I_43410 (I740698,I2690);
DFFARX1 I_43411 (I236409,I2683,I740698,I740724,);
DFFARX1 I_43412 (I236415,I2683,I740698,I740741,);
not I_43413 (I740749,I740741);
not I_43414 (I740766,I236436);
nor I_43415 (I740783,I740766,I236424);
not I_43416 (I740800,I236433);
nor I_43417 (I740817,I740783,I236418);
nor I_43418 (I740834,I740741,I740817);
DFFARX1 I_43419 (I740834,I2683,I740698,I740684,);
nor I_43420 (I740865,I236418,I236424);
nand I_43421 (I740882,I740865,I236436);
DFFARX1 I_43422 (I740882,I2683,I740698,I740687,);
nor I_43423 (I740913,I740800,I236418);
nand I_43424 (I740930,I740913,I236409);
nor I_43425 (I740947,I740724,I740930);
DFFARX1 I_43426 (I740947,I2683,I740698,I740663,);
not I_43427 (I740978,I740930);
nand I_43428 (I740675,I740741,I740978);
DFFARX1 I_43429 (I740930,I2683,I740698,I741018,);
not I_43430 (I741026,I741018);
not I_43431 (I741043,I236418);
not I_43432 (I741060,I236421);
nor I_43433 (I741077,I741060,I236433);
nor I_43434 (I740690,I741026,I741077);
nor I_43435 (I741108,I741060,I236430);
and I_43436 (I741125,I741108,I236412);
or I_43437 (I741142,I741125,I236427);
DFFARX1 I_43438 (I741142,I2683,I740698,I741168,);
nor I_43439 (I740678,I741168,I740724);
not I_43440 (I741190,I741168);
and I_43441 (I741207,I741190,I740724);
nor I_43442 (I740672,I740749,I741207);
nand I_43443 (I741238,I741190,I740800);
nor I_43444 (I740666,I741060,I741238);
nand I_43445 (I740669,I741190,I740978);
nand I_43446 (I741283,I740800,I236421);
nor I_43447 (I740681,I741043,I741283);
not I_43448 (I741344,I2690);
DFFARX1 I_43449 (I277515,I2683,I741344,I741370,);
DFFARX1 I_43450 (I277521,I2683,I741344,I741387,);
not I_43451 (I741395,I741387);
not I_43452 (I741412,I277542);
nor I_43453 (I741429,I741412,I277530);
not I_43454 (I741446,I277539);
nor I_43455 (I741463,I741429,I277524);
nor I_43456 (I741480,I741387,I741463);
DFFARX1 I_43457 (I741480,I2683,I741344,I741330,);
nor I_43458 (I741511,I277524,I277530);
nand I_43459 (I741528,I741511,I277542);
DFFARX1 I_43460 (I741528,I2683,I741344,I741333,);
nor I_43461 (I741559,I741446,I277524);
nand I_43462 (I741576,I741559,I277515);
nor I_43463 (I741593,I741370,I741576);
DFFARX1 I_43464 (I741593,I2683,I741344,I741309,);
not I_43465 (I741624,I741576);
nand I_43466 (I741321,I741387,I741624);
DFFARX1 I_43467 (I741576,I2683,I741344,I741664,);
not I_43468 (I741672,I741664);
not I_43469 (I741689,I277524);
not I_43470 (I741706,I277527);
nor I_43471 (I741723,I741706,I277539);
nor I_43472 (I741336,I741672,I741723);
nor I_43473 (I741754,I741706,I277536);
and I_43474 (I741771,I741754,I277518);
or I_43475 (I741788,I741771,I277533);
DFFARX1 I_43476 (I741788,I2683,I741344,I741814,);
nor I_43477 (I741324,I741814,I741370);
not I_43478 (I741836,I741814);
and I_43479 (I741853,I741836,I741370);
nor I_43480 (I741318,I741395,I741853);
nand I_43481 (I741884,I741836,I741446);
nor I_43482 (I741312,I741706,I741884);
nand I_43483 (I741315,I741836,I741624);
nand I_43484 (I741929,I741446,I277527);
nor I_43485 (I741327,I741689,I741929);
not I_43486 (I741990,I2690);
DFFARX1 I_43487 (I358968,I2683,I741990,I742016,);
DFFARX1 I_43488 (I358965,I2683,I741990,I742033,);
not I_43489 (I742041,I742033);
not I_43490 (I742058,I358980);
nor I_43491 (I742075,I742058,I358983);
not I_43492 (I742092,I358971);
nor I_43493 (I742109,I742075,I358977);
nor I_43494 (I742126,I742033,I742109);
DFFARX1 I_43495 (I742126,I2683,I741990,I741976,);
nor I_43496 (I742157,I358977,I358983);
nand I_43497 (I742174,I742157,I358980);
DFFARX1 I_43498 (I742174,I2683,I741990,I741979,);
nor I_43499 (I742205,I742092,I358977);
nand I_43500 (I742222,I742205,I358989);
nor I_43501 (I742239,I742016,I742222);
DFFARX1 I_43502 (I742239,I2683,I741990,I741955,);
not I_43503 (I742270,I742222);
nand I_43504 (I741967,I742033,I742270);
DFFARX1 I_43505 (I742222,I2683,I741990,I742310,);
not I_43506 (I742318,I742310);
not I_43507 (I742335,I358977);
not I_43508 (I742352,I358962);
nor I_43509 (I742369,I742352,I358971);
nor I_43510 (I741982,I742318,I742369);
nor I_43511 (I742400,I742352,I358974);
and I_43512 (I742417,I742400,I358962);
or I_43513 (I742434,I742417,I358986);
DFFARX1 I_43514 (I742434,I2683,I741990,I742460,);
nor I_43515 (I741970,I742460,I742016);
not I_43516 (I742482,I742460);
and I_43517 (I742499,I742482,I742016);
nor I_43518 (I741964,I742041,I742499);
nand I_43519 (I742530,I742482,I742092);
nor I_43520 (I741958,I742352,I742530);
nand I_43521 (I741961,I742482,I742270);
nand I_43522 (I742575,I742092,I358962);
nor I_43523 (I741973,I742335,I742575);
not I_43524 (I742636,I2690);
DFFARX1 I_43525 (I262232,I2683,I742636,I742662,);
DFFARX1 I_43526 (I262238,I2683,I742636,I742679,);
not I_43527 (I742687,I742679);
not I_43528 (I742704,I262259);
nor I_43529 (I742721,I742704,I262247);
not I_43530 (I742738,I262256);
nor I_43531 (I742755,I742721,I262241);
nor I_43532 (I742772,I742679,I742755);
DFFARX1 I_43533 (I742772,I2683,I742636,I742622,);
nor I_43534 (I742803,I262241,I262247);
nand I_43535 (I742820,I742803,I262259);
DFFARX1 I_43536 (I742820,I2683,I742636,I742625,);
nor I_43537 (I742851,I742738,I262241);
nand I_43538 (I742868,I742851,I262232);
nor I_43539 (I742885,I742662,I742868);
DFFARX1 I_43540 (I742885,I2683,I742636,I742601,);
not I_43541 (I742916,I742868);
nand I_43542 (I742613,I742679,I742916);
DFFARX1 I_43543 (I742868,I2683,I742636,I742956,);
not I_43544 (I742964,I742956);
not I_43545 (I742981,I262241);
not I_43546 (I742998,I262244);
nor I_43547 (I743015,I742998,I262256);
nor I_43548 (I742628,I742964,I743015);
nor I_43549 (I743046,I742998,I262253);
and I_43550 (I743063,I743046,I262235);
or I_43551 (I743080,I743063,I262250);
DFFARX1 I_43552 (I743080,I2683,I742636,I743106,);
nor I_43553 (I742616,I743106,I742662);
not I_43554 (I743128,I743106);
and I_43555 (I743145,I743128,I742662);
nor I_43556 (I742610,I742687,I743145);
nand I_43557 (I743176,I743128,I742738);
nor I_43558 (I742604,I742998,I743176);
nand I_43559 (I742607,I743128,I742916);
nand I_43560 (I743221,I742738,I262244);
nor I_43561 (I742619,I742981,I743221);
not I_43562 (I743282,I2690);
DFFARX1 I_43563 (I595982,I2683,I743282,I743308,);
DFFARX1 I_43564 (I595976,I2683,I743282,I743325,);
not I_43565 (I743333,I743325);
not I_43566 (I743350,I595991);
nor I_43567 (I743367,I743350,I595976);
not I_43568 (I743384,I595985);
nor I_43569 (I743401,I743367,I595994);
nor I_43570 (I743418,I743325,I743401);
DFFARX1 I_43571 (I743418,I2683,I743282,I743268,);
nor I_43572 (I743449,I595994,I595976);
nand I_43573 (I743466,I743449,I595991);
DFFARX1 I_43574 (I743466,I2683,I743282,I743271,);
nor I_43575 (I743497,I743384,I595994);
nand I_43576 (I743514,I743497,I595979);
nor I_43577 (I743531,I743308,I743514);
DFFARX1 I_43578 (I743531,I2683,I743282,I743247,);
not I_43579 (I743562,I743514);
nand I_43580 (I743259,I743325,I743562);
DFFARX1 I_43581 (I743514,I2683,I743282,I743602,);
not I_43582 (I743610,I743602);
not I_43583 (I743627,I595994);
not I_43584 (I743644,I595988);
nor I_43585 (I743661,I743644,I595985);
nor I_43586 (I743274,I743610,I743661);
nor I_43587 (I743692,I743644,I595997);
and I_43588 (I743709,I743692,I596000);
or I_43589 (I743726,I743709,I595979);
DFFARX1 I_43590 (I743726,I2683,I743282,I743752,);
nor I_43591 (I743262,I743752,I743308);
not I_43592 (I743774,I743752);
and I_43593 (I743791,I743774,I743308);
nor I_43594 (I743256,I743333,I743791);
nand I_43595 (I743822,I743774,I743384);
nor I_43596 (I743250,I743644,I743822);
nand I_43597 (I743253,I743774,I743562);
nand I_43598 (I743867,I743384,I595988);
nor I_43599 (I743265,I743627,I743867);
not I_43600 (I743928,I2690);
DFFARX1 I_43601 (I84871,I2683,I743928,I743954,);
DFFARX1 I_43602 (I84877,I2683,I743928,I743971,);
not I_43603 (I743979,I743971);
not I_43604 (I743996,I84895);
nor I_43605 (I744013,I743996,I84874);
not I_43606 (I744030,I84880);
nor I_43607 (I744047,I744013,I84886);
nor I_43608 (I744064,I743971,I744047);
DFFARX1 I_43609 (I744064,I2683,I743928,I743914,);
nor I_43610 (I744095,I84886,I84874);
nand I_43611 (I744112,I744095,I84895);
DFFARX1 I_43612 (I744112,I2683,I743928,I743917,);
nor I_43613 (I744143,I744030,I84886);
nand I_43614 (I744160,I744143,I84892);
nor I_43615 (I744177,I743954,I744160);
DFFARX1 I_43616 (I744177,I2683,I743928,I743893,);
not I_43617 (I744208,I744160);
nand I_43618 (I743905,I743971,I744208);
DFFARX1 I_43619 (I744160,I2683,I743928,I744248,);
not I_43620 (I744256,I744248);
not I_43621 (I744273,I84886);
not I_43622 (I744290,I84874);
nor I_43623 (I744307,I744290,I84880);
nor I_43624 (I743920,I744256,I744307);
nor I_43625 (I744338,I744290,I84883);
and I_43626 (I744355,I744338,I84871);
or I_43627 (I744372,I744355,I84889);
DFFARX1 I_43628 (I744372,I2683,I743928,I744398,);
nor I_43629 (I743908,I744398,I743954);
not I_43630 (I744420,I744398);
and I_43631 (I744437,I744420,I743954);
nor I_43632 (I743902,I743979,I744437);
nand I_43633 (I744468,I744420,I744030);
nor I_43634 (I743896,I744290,I744468);
nand I_43635 (I743899,I744420,I744208);
nand I_43636 (I744513,I744030,I84874);
nor I_43637 (I743911,I744273,I744513);
not I_43638 (I744574,I2690);
DFFARX1 I_43639 (I1061419,I2683,I744574,I744600,);
DFFARX1 I_43640 (I1061443,I2683,I744574,I744617,);
not I_43641 (I744625,I744617);
not I_43642 (I744642,I1061425);
nor I_43643 (I744659,I744642,I1061434);
not I_43644 (I744676,I1061419);
nor I_43645 (I744693,I744659,I1061440);
nor I_43646 (I744710,I744617,I744693);
DFFARX1 I_43647 (I744710,I2683,I744574,I744560,);
nor I_43648 (I744741,I1061440,I1061434);
nand I_43649 (I744758,I744741,I1061425);
DFFARX1 I_43650 (I744758,I2683,I744574,I744563,);
nor I_43651 (I744789,I744676,I1061440);
nand I_43652 (I744806,I744789,I1061437);
nor I_43653 (I744823,I744600,I744806);
DFFARX1 I_43654 (I744823,I2683,I744574,I744539,);
not I_43655 (I744854,I744806);
nand I_43656 (I744551,I744617,I744854);
DFFARX1 I_43657 (I744806,I2683,I744574,I744894,);
not I_43658 (I744902,I744894);
not I_43659 (I744919,I1061440);
not I_43660 (I744936,I1061431);
nor I_43661 (I744953,I744936,I1061419);
nor I_43662 (I744566,I744902,I744953);
nor I_43663 (I744984,I744936,I1061422);
and I_43664 (I745001,I744984,I1061446);
or I_43665 (I745018,I745001,I1061428);
DFFARX1 I_43666 (I745018,I2683,I744574,I745044,);
nor I_43667 (I744554,I745044,I744600);
not I_43668 (I745066,I745044);
and I_43669 (I745083,I745066,I744600);
nor I_43670 (I744548,I744625,I745083);
nand I_43671 (I745114,I745066,I744676);
nor I_43672 (I744542,I744936,I745114);
nand I_43673 (I744545,I745066,I744854);
nand I_43674 (I745159,I744676,I1061431);
nor I_43675 (I744557,I744919,I745159);
not I_43676 (I745220,I2690);
DFFARX1 I_43677 (I63264,I2683,I745220,I745246,);
DFFARX1 I_43678 (I63270,I2683,I745220,I745263,);
not I_43679 (I745271,I745263);
not I_43680 (I745288,I63288);
nor I_43681 (I745305,I745288,I63267);
not I_43682 (I745322,I63273);
nor I_43683 (I745339,I745305,I63279);
nor I_43684 (I745356,I745263,I745339);
DFFARX1 I_43685 (I745356,I2683,I745220,I745206,);
nor I_43686 (I745387,I63279,I63267);
nand I_43687 (I745404,I745387,I63288);
DFFARX1 I_43688 (I745404,I2683,I745220,I745209,);
nor I_43689 (I745435,I745322,I63279);
nand I_43690 (I745452,I745435,I63285);
nor I_43691 (I745469,I745246,I745452);
DFFARX1 I_43692 (I745469,I2683,I745220,I745185,);
not I_43693 (I745500,I745452);
nand I_43694 (I745197,I745263,I745500);
DFFARX1 I_43695 (I745452,I2683,I745220,I745540,);
not I_43696 (I745548,I745540);
not I_43697 (I745565,I63279);
not I_43698 (I745582,I63267);
nor I_43699 (I745599,I745582,I63273);
nor I_43700 (I745212,I745548,I745599);
nor I_43701 (I745630,I745582,I63276);
and I_43702 (I745647,I745630,I63264);
or I_43703 (I745664,I745647,I63282);
DFFARX1 I_43704 (I745664,I2683,I745220,I745690,);
nor I_43705 (I745200,I745690,I745246);
not I_43706 (I745712,I745690);
and I_43707 (I745729,I745712,I745246);
nor I_43708 (I745194,I745271,I745729);
nand I_43709 (I745760,I745712,I745322);
nor I_43710 (I745188,I745582,I745760);
nand I_43711 (I745191,I745712,I745500);
nand I_43712 (I745805,I745322,I63267);
nor I_43713 (I745203,I745565,I745805);
not I_43714 (I745866,I2690);
DFFARX1 I_43715 (I884858,I2683,I745866,I745892,);
DFFARX1 I_43716 (I884840,I2683,I745866,I745909,);
not I_43717 (I745917,I745909);
not I_43718 (I745934,I884849);
nor I_43719 (I745951,I745934,I884861);
not I_43720 (I745968,I884843);
nor I_43721 (I745985,I745951,I884852);
nor I_43722 (I746002,I745909,I745985);
DFFARX1 I_43723 (I746002,I2683,I745866,I745852,);
nor I_43724 (I746033,I884852,I884861);
nand I_43725 (I746050,I746033,I884849);
DFFARX1 I_43726 (I746050,I2683,I745866,I745855,);
nor I_43727 (I746081,I745968,I884852);
nand I_43728 (I746098,I746081,I884864);
nor I_43729 (I746115,I745892,I746098);
DFFARX1 I_43730 (I746115,I2683,I745866,I745831,);
not I_43731 (I746146,I746098);
nand I_43732 (I745843,I745909,I746146);
DFFARX1 I_43733 (I746098,I2683,I745866,I746186,);
not I_43734 (I746194,I746186);
not I_43735 (I746211,I884852);
not I_43736 (I746228,I884840);
nor I_43737 (I746245,I746228,I884843);
nor I_43738 (I745858,I746194,I746245);
nor I_43739 (I746276,I746228,I884846);
and I_43740 (I746293,I746276,I884855);
or I_43741 (I746310,I746293,I884843);
DFFARX1 I_43742 (I746310,I2683,I745866,I746336,);
nor I_43743 (I745846,I746336,I745892);
not I_43744 (I746358,I746336);
and I_43745 (I746375,I746358,I745892);
nor I_43746 (I745840,I745917,I746375);
nand I_43747 (I746406,I746358,I745968);
nor I_43748 (I745834,I746228,I746406);
nand I_43749 (I745837,I746358,I746146);
nand I_43750 (I746451,I745968,I884840);
nor I_43751 (I745849,I746211,I746451);
not I_43752 (I746512,I2690);
DFFARX1 I_43753 (I382904,I2683,I746512,I746538,);
DFFARX1 I_43754 (I382901,I2683,I746512,I746555,);
not I_43755 (I746563,I746555);
not I_43756 (I746580,I382916);
nor I_43757 (I746597,I746580,I382919);
not I_43758 (I746614,I382907);
nor I_43759 (I746631,I746597,I382913);
nor I_43760 (I746648,I746555,I746631);
DFFARX1 I_43761 (I746648,I2683,I746512,I746498,);
nor I_43762 (I746679,I382913,I382919);
nand I_43763 (I746696,I746679,I382916);
DFFARX1 I_43764 (I746696,I2683,I746512,I746501,);
nor I_43765 (I746727,I746614,I382913);
nand I_43766 (I746744,I746727,I382925);
nor I_43767 (I746761,I746538,I746744);
DFFARX1 I_43768 (I746761,I2683,I746512,I746477,);
not I_43769 (I746792,I746744);
nand I_43770 (I746489,I746555,I746792);
DFFARX1 I_43771 (I746744,I2683,I746512,I746832,);
not I_43772 (I746840,I746832);
not I_43773 (I746857,I382913);
not I_43774 (I746874,I382898);
nor I_43775 (I746891,I746874,I382907);
nor I_43776 (I746504,I746840,I746891);
nor I_43777 (I746922,I746874,I382910);
and I_43778 (I746939,I746922,I382898);
or I_43779 (I746956,I746939,I382922);
DFFARX1 I_43780 (I746956,I2683,I746512,I746982,);
nor I_43781 (I746492,I746982,I746538);
not I_43782 (I747004,I746982);
and I_43783 (I747021,I747004,I746538);
nor I_43784 (I746486,I746563,I747021);
nand I_43785 (I747052,I747004,I746614);
nor I_43786 (I746480,I746874,I747052);
nand I_43787 (I746483,I747004,I746792);
nand I_43788 (I747097,I746614,I382898);
nor I_43789 (I746495,I746857,I747097);
not I_43790 (I747158,I2690);
DFFARX1 I_43791 (I420505,I2683,I747158,I747184,);
DFFARX1 I_43792 (I420517,I2683,I747158,I747201,);
not I_43793 (I747209,I747201);
not I_43794 (I747226,I420502);
nor I_43795 (I747243,I747226,I420520);
not I_43796 (I747260,I420526);
nor I_43797 (I747277,I747243,I420508);
nor I_43798 (I747294,I747201,I747277);
DFFARX1 I_43799 (I747294,I2683,I747158,I747144,);
nor I_43800 (I747325,I420508,I420520);
nand I_43801 (I747342,I747325,I420502);
DFFARX1 I_43802 (I747342,I2683,I747158,I747147,);
nor I_43803 (I747373,I747260,I420508);
nand I_43804 (I747390,I747373,I420511);
nor I_43805 (I747407,I747184,I747390);
DFFARX1 I_43806 (I747407,I2683,I747158,I747123,);
not I_43807 (I747438,I747390);
nand I_43808 (I747135,I747201,I747438);
DFFARX1 I_43809 (I747390,I2683,I747158,I747478,);
not I_43810 (I747486,I747478);
not I_43811 (I747503,I420508);
not I_43812 (I747520,I420514);
nor I_43813 (I747537,I747520,I420526);
nor I_43814 (I747150,I747486,I747537);
nor I_43815 (I747568,I747520,I420523);
and I_43816 (I747585,I747568,I420502);
or I_43817 (I747602,I747585,I420505);
DFFARX1 I_43818 (I747602,I2683,I747158,I747628,);
nor I_43819 (I747138,I747628,I747184);
not I_43820 (I747650,I747628);
and I_43821 (I747667,I747650,I747184);
nor I_43822 (I747132,I747209,I747667);
nand I_43823 (I747698,I747650,I747260);
nor I_43824 (I747126,I747520,I747698);
nand I_43825 (I747129,I747650,I747438);
nand I_43826 (I747743,I747260,I420514);
nor I_43827 (I747141,I747503,I747743);
not I_43828 (I747804,I2690);
DFFARX1 I_43829 (I355704,I2683,I747804,I747830,);
DFFARX1 I_43830 (I355701,I2683,I747804,I747847,);
not I_43831 (I747855,I747847);
not I_43832 (I747872,I355716);
nor I_43833 (I747889,I747872,I355719);
not I_43834 (I747906,I355707);
nor I_43835 (I747923,I747889,I355713);
nor I_43836 (I747940,I747847,I747923);
DFFARX1 I_43837 (I747940,I2683,I747804,I747790,);
nor I_43838 (I747971,I355713,I355719);
nand I_43839 (I747988,I747971,I355716);
DFFARX1 I_43840 (I747988,I2683,I747804,I747793,);
nor I_43841 (I748019,I747906,I355713);
nand I_43842 (I748036,I748019,I355725);
nor I_43843 (I748053,I747830,I748036);
DFFARX1 I_43844 (I748053,I2683,I747804,I747769,);
not I_43845 (I748084,I748036);
nand I_43846 (I747781,I747847,I748084);
DFFARX1 I_43847 (I748036,I2683,I747804,I748124,);
not I_43848 (I748132,I748124);
not I_43849 (I748149,I355713);
not I_43850 (I748166,I355698);
nor I_43851 (I748183,I748166,I355707);
nor I_43852 (I747796,I748132,I748183);
nor I_43853 (I748214,I748166,I355710);
and I_43854 (I748231,I748214,I355698);
or I_43855 (I748248,I748231,I355722);
DFFARX1 I_43856 (I748248,I2683,I747804,I748274,);
nor I_43857 (I747784,I748274,I747830);
not I_43858 (I748296,I748274);
and I_43859 (I748313,I748296,I747830);
nor I_43860 (I747778,I747855,I748313);
nand I_43861 (I748344,I748296,I747906);
nor I_43862 (I747772,I748166,I748344);
nand I_43863 (I747775,I748296,I748084);
nand I_43864 (I748389,I747906,I355698);
nor I_43865 (I747787,I748149,I748389);
not I_43866 (I748450,I2690);
DFFARX1 I_43867 (I641236,I2683,I748450,I748476,);
DFFARX1 I_43868 (I641233,I2683,I748450,I748493,);
not I_43869 (I748501,I748493);
not I_43870 (I748518,I641233);
nor I_43871 (I748535,I748518,I641236);
not I_43872 (I748552,I641248);
nor I_43873 (I748569,I748535,I641242);
nor I_43874 (I748586,I748493,I748569);
DFFARX1 I_43875 (I748586,I2683,I748450,I748436,);
nor I_43876 (I748617,I641242,I641236);
nand I_43877 (I748634,I748617,I641233);
DFFARX1 I_43878 (I748634,I2683,I748450,I748439,);
nor I_43879 (I748665,I748552,I641242);
nand I_43880 (I748682,I748665,I641230);
nor I_43881 (I748699,I748476,I748682);
DFFARX1 I_43882 (I748699,I2683,I748450,I748415,);
not I_43883 (I748730,I748682);
nand I_43884 (I748427,I748493,I748730);
DFFARX1 I_43885 (I748682,I2683,I748450,I748770,);
not I_43886 (I748778,I748770);
not I_43887 (I748795,I641242);
not I_43888 (I748812,I641239);
nor I_43889 (I748829,I748812,I641248);
nor I_43890 (I748442,I748778,I748829);
nor I_43891 (I748860,I748812,I641245);
and I_43892 (I748877,I748860,I641251);
or I_43893 (I748894,I748877,I641230);
DFFARX1 I_43894 (I748894,I2683,I748450,I748920,);
nor I_43895 (I748430,I748920,I748476);
not I_43896 (I748942,I748920);
and I_43897 (I748959,I748942,I748476);
nor I_43898 (I748424,I748501,I748959);
nand I_43899 (I748990,I748942,I748552);
nor I_43900 (I748418,I748812,I748990);
nand I_43901 (I748421,I748942,I748730);
nand I_43902 (I749035,I748552,I641239);
nor I_43903 (I748433,I748795,I749035);
not I_43904 (I749096,I2690);
DFFARX1 I_43905 (I555522,I2683,I749096,I749122,);
DFFARX1 I_43906 (I555516,I2683,I749096,I749139,);
not I_43907 (I749147,I749139);
not I_43908 (I749164,I555531);
nor I_43909 (I749181,I749164,I555516);
not I_43910 (I749198,I555525);
nor I_43911 (I749215,I749181,I555534);
nor I_43912 (I749232,I749139,I749215);
DFFARX1 I_43913 (I749232,I2683,I749096,I749082,);
nor I_43914 (I749263,I555534,I555516);
nand I_43915 (I749280,I749263,I555531);
DFFARX1 I_43916 (I749280,I2683,I749096,I749085,);
nor I_43917 (I749311,I749198,I555534);
nand I_43918 (I749328,I749311,I555519);
nor I_43919 (I749345,I749122,I749328);
DFFARX1 I_43920 (I749345,I2683,I749096,I749061,);
not I_43921 (I749376,I749328);
nand I_43922 (I749073,I749139,I749376);
DFFARX1 I_43923 (I749328,I2683,I749096,I749416,);
not I_43924 (I749424,I749416);
not I_43925 (I749441,I555534);
not I_43926 (I749458,I555528);
nor I_43927 (I749475,I749458,I555525);
nor I_43928 (I749088,I749424,I749475);
nor I_43929 (I749506,I749458,I555537);
and I_43930 (I749523,I749506,I555540);
or I_43931 (I749540,I749523,I555519);
DFFARX1 I_43932 (I749540,I2683,I749096,I749566,);
nor I_43933 (I749076,I749566,I749122);
not I_43934 (I749588,I749566);
and I_43935 (I749605,I749588,I749122);
nor I_43936 (I749070,I749147,I749605);
nand I_43937 (I749636,I749588,I749198);
nor I_43938 (I749064,I749458,I749636);
nand I_43939 (I749067,I749588,I749376);
nand I_43940 (I749681,I749198,I555528);
nor I_43941 (I749079,I749441,I749681);
not I_43942 (I749742,I2690);
DFFARX1 I_43943 (I682342,I2683,I749742,I749768,);
DFFARX1 I_43944 (I682339,I2683,I749742,I749785,);
not I_43945 (I749793,I749785);
not I_43946 (I749810,I682339);
nor I_43947 (I749827,I749810,I682342);
not I_43948 (I749844,I682354);
nor I_43949 (I749861,I749827,I682348);
nor I_43950 (I749878,I749785,I749861);
DFFARX1 I_43951 (I749878,I2683,I749742,I749728,);
nor I_43952 (I749909,I682348,I682342);
nand I_43953 (I749926,I749909,I682339);
DFFARX1 I_43954 (I749926,I2683,I749742,I749731,);
nor I_43955 (I749957,I749844,I682348);
nand I_43956 (I749974,I749957,I682336);
nor I_43957 (I749991,I749768,I749974);
DFFARX1 I_43958 (I749991,I2683,I749742,I749707,);
not I_43959 (I750022,I749974);
nand I_43960 (I749719,I749785,I750022);
DFFARX1 I_43961 (I749974,I2683,I749742,I750062,);
not I_43962 (I750070,I750062);
not I_43963 (I750087,I682348);
not I_43964 (I750104,I682345);
nor I_43965 (I750121,I750104,I682354);
nor I_43966 (I749734,I750070,I750121);
nor I_43967 (I750152,I750104,I682351);
and I_43968 (I750169,I750152,I682357);
or I_43969 (I750186,I750169,I682336);
DFFARX1 I_43970 (I750186,I2683,I749742,I750212,);
nor I_43971 (I749722,I750212,I749768);
not I_43972 (I750234,I750212);
and I_43973 (I750251,I750234,I749768);
nor I_43974 (I749716,I749793,I750251);
nand I_43975 (I750282,I750234,I749844);
nor I_43976 (I749710,I750104,I750282);
nand I_43977 (I749713,I750234,I750022);
nand I_43978 (I750327,I749844,I682345);
nor I_43979 (I749725,I750087,I750327);
not I_43980 (I750388,I2690);
DFFARX1 I_43981 (I663897,I2683,I750388,I750414,);
DFFARX1 I_43982 (I663894,I2683,I750388,I750431,);
not I_43983 (I750439,I750431);
not I_43984 (I750456,I663894);
nor I_43985 (I750473,I750456,I663897);
not I_43986 (I750490,I663909);
nor I_43987 (I750507,I750473,I663903);
nor I_43988 (I750524,I750431,I750507);
DFFARX1 I_43989 (I750524,I2683,I750388,I750374,);
nor I_43990 (I750555,I663903,I663897);
nand I_43991 (I750572,I750555,I663894);
DFFARX1 I_43992 (I750572,I2683,I750388,I750377,);
nor I_43993 (I750603,I750490,I663903);
nand I_43994 (I750620,I750603,I663891);
nor I_43995 (I750637,I750414,I750620);
DFFARX1 I_43996 (I750637,I2683,I750388,I750353,);
not I_43997 (I750668,I750620);
nand I_43998 (I750365,I750431,I750668);
DFFARX1 I_43999 (I750620,I2683,I750388,I750708,);
not I_44000 (I750716,I750708);
not I_44001 (I750733,I663903);
not I_44002 (I750750,I663900);
nor I_44003 (I750767,I750750,I663909);
nor I_44004 (I750380,I750716,I750767);
nor I_44005 (I750798,I750750,I663906);
and I_44006 (I750815,I750798,I663912);
or I_44007 (I750832,I750815,I663891);
DFFARX1 I_44008 (I750832,I2683,I750388,I750858,);
nor I_44009 (I750368,I750858,I750414);
not I_44010 (I750880,I750858);
and I_44011 (I750897,I750880,I750414);
nor I_44012 (I750362,I750439,I750897);
nand I_44013 (I750928,I750880,I750490);
nor I_44014 (I750356,I750750,I750928);
nand I_44015 (I750359,I750880,I750668);
nand I_44016 (I750973,I750490,I663900);
nor I_44017 (I750371,I750733,I750973);
not I_44018 (I751034,I2690);
DFFARX1 I_44019 (I190226,I2683,I751034,I751060,);
DFFARX1 I_44020 (I190238,I2683,I751034,I751077,);
not I_44021 (I751085,I751077);
not I_44022 (I751102,I190244);
nor I_44023 (I751119,I751102,I190229);
not I_44024 (I751136,I190220);
nor I_44025 (I751153,I751119,I190241);
nor I_44026 (I751170,I751077,I751153);
DFFARX1 I_44027 (I751170,I2683,I751034,I751020,);
nor I_44028 (I751201,I190241,I190229);
nand I_44029 (I751218,I751201,I190244);
DFFARX1 I_44030 (I751218,I2683,I751034,I751023,);
nor I_44031 (I751249,I751136,I190241);
nand I_44032 (I751266,I751249,I190223);
nor I_44033 (I751283,I751060,I751266);
DFFARX1 I_44034 (I751283,I2683,I751034,I750999,);
not I_44035 (I751314,I751266);
nand I_44036 (I751011,I751077,I751314);
DFFARX1 I_44037 (I751266,I2683,I751034,I751354,);
not I_44038 (I751362,I751354);
not I_44039 (I751379,I190241);
not I_44040 (I751396,I190232);
nor I_44041 (I751413,I751396,I190220);
nor I_44042 (I751026,I751362,I751413);
nor I_44043 (I751444,I751396,I190235);
and I_44044 (I751461,I751444,I190223);
or I_44045 (I751478,I751461,I190220);
DFFARX1 I_44046 (I751478,I2683,I751034,I751504,);
nor I_44047 (I751014,I751504,I751060);
not I_44048 (I751526,I751504);
and I_44049 (I751543,I751526,I751060);
nor I_44050 (I751008,I751085,I751543);
nand I_44051 (I751574,I751526,I751136);
nor I_44052 (I751002,I751396,I751574);
nand I_44053 (I751005,I751526,I751314);
nand I_44054 (I751619,I751136,I190232);
nor I_44055 (I751017,I751379,I751619);
not I_44056 (I751680,I2690);
DFFARX1 I_44057 (I933410,I2683,I751680,I751706,);
DFFARX1 I_44058 (I933392,I2683,I751680,I751723,);
not I_44059 (I751731,I751723);
not I_44060 (I751748,I933401);
nor I_44061 (I751765,I751748,I933413);
not I_44062 (I751782,I933395);
nor I_44063 (I751799,I751765,I933404);
nor I_44064 (I751816,I751723,I751799);
DFFARX1 I_44065 (I751816,I2683,I751680,I751666,);
nor I_44066 (I751847,I933404,I933413);
nand I_44067 (I751864,I751847,I933401);
DFFARX1 I_44068 (I751864,I2683,I751680,I751669,);
nor I_44069 (I751895,I751782,I933404);
nand I_44070 (I751912,I751895,I933416);
nor I_44071 (I751929,I751706,I751912);
DFFARX1 I_44072 (I751929,I2683,I751680,I751645,);
not I_44073 (I751960,I751912);
nand I_44074 (I751657,I751723,I751960);
DFFARX1 I_44075 (I751912,I2683,I751680,I752000,);
not I_44076 (I752008,I752000);
not I_44077 (I752025,I933404);
not I_44078 (I752042,I933392);
nor I_44079 (I752059,I752042,I933395);
nor I_44080 (I751672,I752008,I752059);
nor I_44081 (I752090,I752042,I933398);
and I_44082 (I752107,I752090,I933407);
or I_44083 (I752124,I752107,I933395);
DFFARX1 I_44084 (I752124,I2683,I751680,I752150,);
nor I_44085 (I751660,I752150,I751706);
not I_44086 (I752172,I752150);
and I_44087 (I752189,I752172,I751706);
nor I_44088 (I751654,I751731,I752189);
nand I_44089 (I752220,I752172,I751782);
nor I_44090 (I751648,I752042,I752220);
nand I_44091 (I751651,I752172,I751960);
nand I_44092 (I752265,I751782,I933392);
nor I_44093 (I751663,I752025,I752265);
not I_44094 (I752326,I2690);
DFFARX1 I_44095 (I683396,I2683,I752326,I752352,);
DFFARX1 I_44096 (I683393,I2683,I752326,I752369,);
not I_44097 (I752377,I752369);
not I_44098 (I752394,I683393);
nor I_44099 (I752411,I752394,I683396);
not I_44100 (I752428,I683408);
nor I_44101 (I752445,I752411,I683402);
nor I_44102 (I752462,I752369,I752445);
DFFARX1 I_44103 (I752462,I2683,I752326,I752312,);
nor I_44104 (I752493,I683402,I683396);
nand I_44105 (I752510,I752493,I683393);
DFFARX1 I_44106 (I752510,I2683,I752326,I752315,);
nor I_44107 (I752541,I752428,I683402);
nand I_44108 (I752558,I752541,I683390);
nor I_44109 (I752575,I752352,I752558);
DFFARX1 I_44110 (I752575,I2683,I752326,I752291,);
not I_44111 (I752606,I752558);
nand I_44112 (I752303,I752369,I752606);
DFFARX1 I_44113 (I752558,I2683,I752326,I752646,);
not I_44114 (I752654,I752646);
not I_44115 (I752671,I683402);
not I_44116 (I752688,I683399);
nor I_44117 (I752705,I752688,I683408);
nor I_44118 (I752318,I752654,I752705);
nor I_44119 (I752736,I752688,I683405);
and I_44120 (I752753,I752736,I683411);
or I_44121 (I752770,I752753,I683390);
DFFARX1 I_44122 (I752770,I2683,I752326,I752796,);
nor I_44123 (I752306,I752796,I752352);
not I_44124 (I752818,I752796);
and I_44125 (I752835,I752818,I752352);
nor I_44126 (I752300,I752377,I752835);
nand I_44127 (I752866,I752818,I752428);
nor I_44128 (I752294,I752688,I752866);
nand I_44129 (I752297,I752818,I752606);
nand I_44130 (I752911,I752428,I683399);
nor I_44131 (I752309,I752671,I752911);
not I_44132 (I752972,I2690);
DFFARX1 I_44133 (I416935,I2683,I752972,I752998,);
DFFARX1 I_44134 (I416947,I2683,I752972,I753015,);
not I_44135 (I753023,I753015);
not I_44136 (I753040,I416932);
nor I_44137 (I753057,I753040,I416950);
not I_44138 (I753074,I416956);
nor I_44139 (I753091,I753057,I416938);
nor I_44140 (I753108,I753015,I753091);
DFFARX1 I_44141 (I753108,I2683,I752972,I752958,);
nor I_44142 (I753139,I416938,I416950);
nand I_44143 (I753156,I753139,I416932);
DFFARX1 I_44144 (I753156,I2683,I752972,I752961,);
nor I_44145 (I753187,I753074,I416938);
nand I_44146 (I753204,I753187,I416941);
nor I_44147 (I753221,I752998,I753204);
DFFARX1 I_44148 (I753221,I2683,I752972,I752937,);
not I_44149 (I753252,I753204);
nand I_44150 (I752949,I753015,I753252);
DFFARX1 I_44151 (I753204,I2683,I752972,I753292,);
not I_44152 (I753300,I753292);
not I_44153 (I753317,I416938);
not I_44154 (I753334,I416944);
nor I_44155 (I753351,I753334,I416956);
nor I_44156 (I752964,I753300,I753351);
nor I_44157 (I753382,I753334,I416953);
and I_44158 (I753399,I753382,I416932);
or I_44159 (I753416,I753399,I416935);
DFFARX1 I_44160 (I753416,I2683,I752972,I753442,);
nor I_44161 (I752952,I753442,I752998);
not I_44162 (I753464,I753442);
and I_44163 (I753481,I753464,I752998);
nor I_44164 (I752946,I753023,I753481);
nand I_44165 (I753512,I753464,I753074);
nor I_44166 (I752940,I753334,I753512);
nand I_44167 (I752943,I753464,I753252);
nand I_44168 (I753557,I753074,I416944);
nor I_44169 (I752955,I753317,I753557);
not I_44170 (I753618,I2690);
DFFARX1 I_44171 (I299649,I2683,I753618,I753644,);
DFFARX1 I_44172 (I299655,I2683,I753618,I753661,);
not I_44173 (I753669,I753661);
not I_44174 (I753686,I299676);
nor I_44175 (I753703,I753686,I299664);
not I_44176 (I753720,I299673);
nor I_44177 (I753737,I753703,I299658);
nor I_44178 (I753754,I753661,I753737);
DFFARX1 I_44179 (I753754,I2683,I753618,I753604,);
nor I_44180 (I753785,I299658,I299664);
nand I_44181 (I753802,I753785,I299676);
DFFARX1 I_44182 (I753802,I2683,I753618,I753607,);
nor I_44183 (I753833,I753720,I299658);
nand I_44184 (I753850,I753833,I299649);
nor I_44185 (I753867,I753644,I753850);
DFFARX1 I_44186 (I753867,I2683,I753618,I753583,);
not I_44187 (I753898,I753850);
nand I_44188 (I753595,I753661,I753898);
DFFARX1 I_44189 (I753850,I2683,I753618,I753938,);
not I_44190 (I753946,I753938);
not I_44191 (I753963,I299658);
not I_44192 (I753980,I299661);
nor I_44193 (I753997,I753980,I299673);
nor I_44194 (I753610,I753946,I753997);
nor I_44195 (I754028,I753980,I299670);
and I_44196 (I754045,I754028,I299652);
or I_44197 (I754062,I754045,I299667);
DFFARX1 I_44198 (I754062,I2683,I753618,I754088,);
nor I_44199 (I753598,I754088,I753644);
not I_44200 (I754110,I754088);
and I_44201 (I754127,I754110,I753644);
nor I_44202 (I753592,I753669,I754127);
nand I_44203 (I754158,I754110,I753720);
nor I_44204 (I753586,I753980,I754158);
nand I_44205 (I753589,I754110,I753898);
nand I_44206 (I754203,I753720,I299661);
nor I_44207 (I753601,I753963,I754203);
not I_44208 (I754264,I2690);
DFFARX1 I_44209 (I451479,I2683,I754264,I754290,);
DFFARX1 I_44210 (I451491,I2683,I754264,I754307,);
not I_44211 (I754315,I754307);
not I_44212 (I754332,I451500);
nor I_44213 (I754349,I754332,I451476);
not I_44214 (I754366,I451494);
nor I_44215 (I754383,I754349,I451488);
nor I_44216 (I754400,I754307,I754383);
DFFARX1 I_44217 (I754400,I2683,I754264,I754250,);
nor I_44218 (I754431,I451488,I451476);
nand I_44219 (I754448,I754431,I451500);
DFFARX1 I_44220 (I754448,I2683,I754264,I754253,);
nor I_44221 (I754479,I754366,I451488);
nand I_44222 (I754496,I754479,I451482);
nor I_44223 (I754513,I754290,I754496);
DFFARX1 I_44224 (I754513,I2683,I754264,I754229,);
not I_44225 (I754544,I754496);
nand I_44226 (I754241,I754307,I754544);
DFFARX1 I_44227 (I754496,I2683,I754264,I754584,);
not I_44228 (I754592,I754584);
not I_44229 (I754609,I451488);
not I_44230 (I754626,I451497);
nor I_44231 (I754643,I754626,I451494);
nor I_44232 (I754256,I754592,I754643);
nor I_44233 (I754674,I754626,I451479);
and I_44234 (I754691,I754674,I451476);
or I_44235 (I754708,I754691,I451485);
DFFARX1 I_44236 (I754708,I2683,I754264,I754734,);
nor I_44237 (I754244,I754734,I754290);
not I_44238 (I754756,I754734);
and I_44239 (I754773,I754756,I754290);
nor I_44240 (I754238,I754315,I754773);
nand I_44241 (I754804,I754756,I754366);
nor I_44242 (I754232,I754626,I754804);
nand I_44243 (I754235,I754756,I754544);
nand I_44244 (I754849,I754366,I451497);
nor I_44245 (I754247,I754609,I754849);
not I_44246 (I754910,I2690);
DFFARX1 I_44247 (I642817,I2683,I754910,I754936,);
DFFARX1 I_44248 (I642814,I2683,I754910,I754953,);
not I_44249 (I754961,I754953);
not I_44250 (I754978,I642814);
nor I_44251 (I754995,I754978,I642817);
not I_44252 (I755012,I642829);
nor I_44253 (I755029,I754995,I642823);
nor I_44254 (I755046,I754953,I755029);
DFFARX1 I_44255 (I755046,I2683,I754910,I754896,);
nor I_44256 (I755077,I642823,I642817);
nand I_44257 (I755094,I755077,I642814);
DFFARX1 I_44258 (I755094,I2683,I754910,I754899,);
nor I_44259 (I755125,I755012,I642823);
nand I_44260 (I755142,I755125,I642811);
nor I_44261 (I755159,I754936,I755142);
DFFARX1 I_44262 (I755159,I2683,I754910,I754875,);
not I_44263 (I755190,I755142);
nand I_44264 (I754887,I754953,I755190);
DFFARX1 I_44265 (I755142,I2683,I754910,I755230,);
not I_44266 (I755238,I755230);
not I_44267 (I755255,I642823);
not I_44268 (I755272,I642820);
nor I_44269 (I755289,I755272,I642829);
nor I_44270 (I754902,I755238,I755289);
nor I_44271 (I755320,I755272,I642826);
and I_44272 (I755337,I755320,I642832);
or I_44273 (I755354,I755337,I642811);
DFFARX1 I_44274 (I755354,I2683,I754910,I755380,);
nor I_44275 (I754890,I755380,I754936);
not I_44276 (I755402,I755380);
and I_44277 (I755419,I755402,I754936);
nor I_44278 (I754884,I754961,I755419);
nand I_44279 (I755450,I755402,I755012);
nor I_44280 (I754878,I755272,I755450);
nand I_44281 (I754881,I755402,I755190);
nand I_44282 (I755495,I755012,I642820);
nor I_44283 (I754893,I755255,I755495);
not I_44284 (I755556,I2690);
DFFARX1 I_44285 (I646506,I2683,I755556,I755582,);
DFFARX1 I_44286 (I646503,I2683,I755556,I755599,);
not I_44287 (I755607,I755599);
not I_44288 (I755624,I646503);
nor I_44289 (I755641,I755624,I646506);
not I_44290 (I755658,I646518);
nor I_44291 (I755675,I755641,I646512);
nor I_44292 (I755692,I755599,I755675);
DFFARX1 I_44293 (I755692,I2683,I755556,I755542,);
nor I_44294 (I755723,I646512,I646506);
nand I_44295 (I755740,I755723,I646503);
DFFARX1 I_44296 (I755740,I2683,I755556,I755545,);
nor I_44297 (I755771,I755658,I646512);
nand I_44298 (I755788,I755771,I646500);
nor I_44299 (I755805,I755582,I755788);
DFFARX1 I_44300 (I755805,I2683,I755556,I755521,);
not I_44301 (I755836,I755788);
nand I_44302 (I755533,I755599,I755836);
DFFARX1 I_44303 (I755788,I2683,I755556,I755876,);
not I_44304 (I755884,I755876);
not I_44305 (I755901,I646512);
not I_44306 (I755918,I646509);
nor I_44307 (I755935,I755918,I646518);
nor I_44308 (I755548,I755884,I755935);
nor I_44309 (I755966,I755918,I646515);
and I_44310 (I755983,I755966,I646521);
or I_44311 (I756000,I755983,I646500);
DFFARX1 I_44312 (I756000,I2683,I755556,I756026,);
nor I_44313 (I755536,I756026,I755582);
not I_44314 (I756048,I756026);
and I_44315 (I756065,I756048,I755582);
nor I_44316 (I755530,I755607,I756065);
nand I_44317 (I756096,I756048,I755658);
nor I_44318 (I755524,I755918,I756096);
nand I_44319 (I755527,I756048,I755836);
nand I_44320 (I756141,I755658,I646509);
nor I_44321 (I755539,I755901,I756141);
not I_44322 (I756202,I2690);
DFFARX1 I_44323 (I842664,I2683,I756202,I756228,);
DFFARX1 I_44324 (I842646,I2683,I756202,I756245,);
not I_44325 (I756253,I756245);
not I_44326 (I756270,I842655);
nor I_44327 (I756287,I756270,I842667);
not I_44328 (I756304,I842649);
nor I_44329 (I756321,I756287,I842658);
nor I_44330 (I756338,I756245,I756321);
DFFARX1 I_44331 (I756338,I2683,I756202,I756188,);
nor I_44332 (I756369,I842658,I842667);
nand I_44333 (I756386,I756369,I842655);
DFFARX1 I_44334 (I756386,I2683,I756202,I756191,);
nor I_44335 (I756417,I756304,I842658);
nand I_44336 (I756434,I756417,I842670);
nor I_44337 (I756451,I756228,I756434);
DFFARX1 I_44338 (I756451,I2683,I756202,I756167,);
not I_44339 (I756482,I756434);
nand I_44340 (I756179,I756245,I756482);
DFFARX1 I_44341 (I756434,I2683,I756202,I756522,);
not I_44342 (I756530,I756522);
not I_44343 (I756547,I842658);
not I_44344 (I756564,I842646);
nor I_44345 (I756581,I756564,I842649);
nor I_44346 (I756194,I756530,I756581);
nor I_44347 (I756612,I756564,I842652);
and I_44348 (I756629,I756612,I842661);
or I_44349 (I756646,I756629,I842649);
DFFARX1 I_44350 (I756646,I2683,I756202,I756672,);
nor I_44351 (I756182,I756672,I756228);
not I_44352 (I756694,I756672);
and I_44353 (I756711,I756694,I756228);
nor I_44354 (I756176,I756253,I756711);
nand I_44355 (I756742,I756694,I756304);
nor I_44356 (I756170,I756564,I756742);
nand I_44357 (I756173,I756694,I756482);
nand I_44358 (I756787,I756304,I842646);
nor I_44359 (I756185,I756547,I756787);
not I_44360 (I756848,I2690);
DFFARX1 I_44361 (I551476,I2683,I756848,I756874,);
DFFARX1 I_44362 (I551470,I2683,I756848,I756891,);
not I_44363 (I756899,I756891);
not I_44364 (I756916,I551485);
nor I_44365 (I756933,I756916,I551470);
not I_44366 (I756950,I551479);
nor I_44367 (I756967,I756933,I551488);
nor I_44368 (I756984,I756891,I756967);
DFFARX1 I_44369 (I756984,I2683,I756848,I756834,);
nor I_44370 (I757015,I551488,I551470);
nand I_44371 (I757032,I757015,I551485);
DFFARX1 I_44372 (I757032,I2683,I756848,I756837,);
nor I_44373 (I757063,I756950,I551488);
nand I_44374 (I757080,I757063,I551473);
nor I_44375 (I757097,I756874,I757080);
DFFARX1 I_44376 (I757097,I2683,I756848,I756813,);
not I_44377 (I757128,I757080);
nand I_44378 (I756825,I756891,I757128);
DFFARX1 I_44379 (I757080,I2683,I756848,I757168,);
not I_44380 (I757176,I757168);
not I_44381 (I757193,I551488);
not I_44382 (I757210,I551482);
nor I_44383 (I757227,I757210,I551479);
nor I_44384 (I756840,I757176,I757227);
nor I_44385 (I757258,I757210,I551491);
and I_44386 (I757275,I757258,I551494);
or I_44387 (I757292,I757275,I551473);
DFFARX1 I_44388 (I757292,I2683,I756848,I757318,);
nor I_44389 (I756828,I757318,I756874);
not I_44390 (I757340,I757318);
and I_44391 (I757357,I757340,I756874);
nor I_44392 (I756822,I756899,I757357);
nand I_44393 (I757388,I757340,I756950);
nor I_44394 (I756816,I757210,I757388);
nand I_44395 (I756819,I757340,I757128);
nand I_44396 (I757433,I756950,I551482);
nor I_44397 (I756831,I757193,I757433);
not I_44398 (I757494,I2690);
DFFARX1 I_44399 (I450901,I2683,I757494,I757520,);
DFFARX1 I_44400 (I450913,I2683,I757494,I757537,);
not I_44401 (I757545,I757537);
not I_44402 (I757562,I450922);
nor I_44403 (I757579,I757562,I450898);
not I_44404 (I757596,I450916);
nor I_44405 (I757613,I757579,I450910);
nor I_44406 (I757630,I757537,I757613);
DFFARX1 I_44407 (I757630,I2683,I757494,I757480,);
nor I_44408 (I757661,I450910,I450898);
nand I_44409 (I757678,I757661,I450922);
DFFARX1 I_44410 (I757678,I2683,I757494,I757483,);
nor I_44411 (I757709,I757596,I450910);
nand I_44412 (I757726,I757709,I450904);
nor I_44413 (I757743,I757520,I757726);
DFFARX1 I_44414 (I757743,I2683,I757494,I757459,);
not I_44415 (I757774,I757726);
nand I_44416 (I757471,I757537,I757774);
DFFARX1 I_44417 (I757726,I2683,I757494,I757814,);
not I_44418 (I757822,I757814);
not I_44419 (I757839,I450910);
not I_44420 (I757856,I450919);
nor I_44421 (I757873,I757856,I450916);
nor I_44422 (I757486,I757822,I757873);
nor I_44423 (I757904,I757856,I450901);
and I_44424 (I757921,I757904,I450898);
or I_44425 (I757938,I757921,I450907);
DFFARX1 I_44426 (I757938,I2683,I757494,I757964,);
nor I_44427 (I757474,I757964,I757520);
not I_44428 (I757986,I757964);
and I_44429 (I758003,I757986,I757520);
nor I_44430 (I757468,I757545,I758003);
nand I_44431 (I758034,I757986,I757596);
nor I_44432 (I757462,I757856,I758034);
nand I_44433 (I757465,I757986,I757774);
nand I_44434 (I758079,I757596,I450919);
nor I_44435 (I757477,I757839,I758079);
not I_44436 (I758140,I2690);
DFFARX1 I_44437 (I644925,I2683,I758140,I758166,);
DFFARX1 I_44438 (I644922,I2683,I758140,I758183,);
not I_44439 (I758191,I758183);
not I_44440 (I758208,I644922);
nor I_44441 (I758225,I758208,I644925);
not I_44442 (I758242,I644937);
nor I_44443 (I758259,I758225,I644931);
nor I_44444 (I758276,I758183,I758259);
DFFARX1 I_44445 (I758276,I2683,I758140,I758126,);
nor I_44446 (I758307,I644931,I644925);
nand I_44447 (I758324,I758307,I644922);
DFFARX1 I_44448 (I758324,I2683,I758140,I758129,);
nor I_44449 (I758355,I758242,I644931);
nand I_44450 (I758372,I758355,I644919);
nor I_44451 (I758389,I758166,I758372);
DFFARX1 I_44452 (I758389,I2683,I758140,I758105,);
not I_44453 (I758420,I758372);
nand I_44454 (I758117,I758183,I758420);
DFFARX1 I_44455 (I758372,I2683,I758140,I758460,);
not I_44456 (I758468,I758460);
not I_44457 (I758485,I644931);
not I_44458 (I758502,I644928);
nor I_44459 (I758519,I758502,I644937);
nor I_44460 (I758132,I758468,I758519);
nor I_44461 (I758550,I758502,I644934);
and I_44462 (I758567,I758550,I644940);
or I_44463 (I758584,I758567,I644919);
DFFARX1 I_44464 (I758584,I2683,I758140,I758610,);
nor I_44465 (I758120,I758610,I758166);
not I_44466 (I758632,I758610);
and I_44467 (I758649,I758632,I758166);
nor I_44468 (I758114,I758191,I758649);
nand I_44469 (I758680,I758632,I758242);
nor I_44470 (I758108,I758502,I758680);
nand I_44471 (I758111,I758632,I758420);
nand I_44472 (I758725,I758242,I644928);
nor I_44473 (I758123,I758485,I758725);
not I_44474 (I758786,I2690);
DFFARX1 I_44475 (I416340,I2683,I758786,I758812,);
DFFARX1 I_44476 (I416352,I2683,I758786,I758829,);
not I_44477 (I758837,I758829);
not I_44478 (I758854,I416337);
nor I_44479 (I758871,I758854,I416355);
not I_44480 (I758888,I416361);
nor I_44481 (I758905,I758871,I416343);
nor I_44482 (I758922,I758829,I758905);
DFFARX1 I_44483 (I758922,I2683,I758786,I758772,);
nor I_44484 (I758953,I416343,I416355);
nand I_44485 (I758970,I758953,I416337);
DFFARX1 I_44486 (I758970,I2683,I758786,I758775,);
nor I_44487 (I759001,I758888,I416343);
nand I_44488 (I759018,I759001,I416346);
nor I_44489 (I759035,I758812,I759018);
DFFARX1 I_44490 (I759035,I2683,I758786,I758751,);
not I_44491 (I759066,I759018);
nand I_44492 (I758763,I758829,I759066);
DFFARX1 I_44493 (I759018,I2683,I758786,I759106,);
not I_44494 (I759114,I759106);
not I_44495 (I759131,I416343);
not I_44496 (I759148,I416349);
nor I_44497 (I759165,I759148,I416361);
nor I_44498 (I758778,I759114,I759165);
nor I_44499 (I759196,I759148,I416358);
and I_44500 (I759213,I759196,I416337);
or I_44501 (I759230,I759213,I416340);
DFFARX1 I_44502 (I759230,I2683,I758786,I759256,);
nor I_44503 (I758766,I759256,I758812);
not I_44504 (I759278,I759256);
and I_44505 (I759295,I759278,I758812);
nor I_44506 (I758760,I758837,I759295);
nand I_44507 (I759326,I759278,I758888);
nor I_44508 (I758754,I759148,I759326);
nand I_44509 (I758757,I759278,I759066);
nand I_44510 (I759371,I758888,I416349);
nor I_44511 (I758769,I759131,I759371);
not I_44512 (I759432,I2690);
DFFARX1 I_44513 (I1031669,I2683,I759432,I759458,);
DFFARX1 I_44514 (I1031693,I2683,I759432,I759475,);
not I_44515 (I759483,I759475);
not I_44516 (I759500,I1031675);
nor I_44517 (I759517,I759500,I1031684);
not I_44518 (I759534,I1031669);
nor I_44519 (I759551,I759517,I1031690);
nor I_44520 (I759568,I759475,I759551);
DFFARX1 I_44521 (I759568,I2683,I759432,I759418,);
nor I_44522 (I759599,I1031690,I1031684);
nand I_44523 (I759616,I759599,I1031675);
DFFARX1 I_44524 (I759616,I2683,I759432,I759421,);
nor I_44525 (I759647,I759534,I1031690);
nand I_44526 (I759664,I759647,I1031687);
nor I_44527 (I759681,I759458,I759664);
DFFARX1 I_44528 (I759681,I2683,I759432,I759397,);
not I_44529 (I759712,I759664);
nand I_44530 (I759409,I759475,I759712);
DFFARX1 I_44531 (I759664,I2683,I759432,I759752,);
not I_44532 (I759760,I759752);
not I_44533 (I759777,I1031690);
not I_44534 (I759794,I1031681);
nor I_44535 (I759811,I759794,I1031669);
nor I_44536 (I759424,I759760,I759811);
nor I_44537 (I759842,I759794,I1031672);
and I_44538 (I759859,I759842,I1031696);
or I_44539 (I759876,I759859,I1031678);
DFFARX1 I_44540 (I759876,I2683,I759432,I759902,);
nor I_44541 (I759412,I759902,I759458);
not I_44542 (I759924,I759902);
and I_44543 (I759941,I759924,I759458);
nor I_44544 (I759406,I759483,I759941);
nand I_44545 (I759972,I759924,I759534);
nor I_44546 (I759400,I759794,I759972);
nand I_44547 (I759403,I759924,I759712);
nand I_44548 (I760017,I759534,I1031681);
nor I_44549 (I759415,I759777,I760017);
not I_44550 (I760078,I2690);
DFFARX1 I_44551 (I853646,I2683,I760078,I760104,);
DFFARX1 I_44552 (I853628,I2683,I760078,I760121,);
not I_44553 (I760129,I760121);
not I_44554 (I760146,I853637);
nor I_44555 (I760163,I760146,I853649);
not I_44556 (I760180,I853631);
nor I_44557 (I760197,I760163,I853640);
nor I_44558 (I760214,I760121,I760197);
DFFARX1 I_44559 (I760214,I2683,I760078,I760064,);
nor I_44560 (I760245,I853640,I853649);
nand I_44561 (I760262,I760245,I853637);
DFFARX1 I_44562 (I760262,I2683,I760078,I760067,);
nor I_44563 (I760293,I760180,I853640);
nand I_44564 (I760310,I760293,I853652);
nor I_44565 (I760327,I760104,I760310);
DFFARX1 I_44566 (I760327,I2683,I760078,I760043,);
not I_44567 (I760358,I760310);
nand I_44568 (I760055,I760121,I760358);
DFFARX1 I_44569 (I760310,I2683,I760078,I760398,);
not I_44570 (I760406,I760398);
not I_44571 (I760423,I853640);
not I_44572 (I760440,I853628);
nor I_44573 (I760457,I760440,I853631);
nor I_44574 (I760070,I760406,I760457);
nor I_44575 (I760488,I760440,I853634);
and I_44576 (I760505,I760488,I853643);
or I_44577 (I760522,I760505,I853631);
DFFARX1 I_44578 (I760522,I2683,I760078,I760548,);
nor I_44579 (I760058,I760548,I760104);
not I_44580 (I760570,I760548);
and I_44581 (I760587,I760570,I760104);
nor I_44582 (I760052,I760129,I760587);
nand I_44583 (I760618,I760570,I760180);
nor I_44584 (I760046,I760440,I760618);
nand I_44585 (I760049,I760570,I760358);
nand I_44586 (I760663,I760180,I853628);
nor I_44587 (I760061,I760423,I760663);
not I_44588 (I760724,I2690);
DFFARX1 I_44589 (I872720,I2683,I760724,I760750,);
DFFARX1 I_44590 (I872702,I2683,I760724,I760767,);
not I_44591 (I760775,I760767);
not I_44592 (I760792,I872711);
nor I_44593 (I760809,I760792,I872723);
not I_44594 (I760826,I872705);
nor I_44595 (I760843,I760809,I872714);
nor I_44596 (I760860,I760767,I760843);
DFFARX1 I_44597 (I760860,I2683,I760724,I760710,);
nor I_44598 (I760891,I872714,I872723);
nand I_44599 (I760908,I760891,I872711);
DFFARX1 I_44600 (I760908,I2683,I760724,I760713,);
nor I_44601 (I760939,I760826,I872714);
nand I_44602 (I760956,I760939,I872726);
nor I_44603 (I760973,I760750,I760956);
DFFARX1 I_44604 (I760973,I2683,I760724,I760689,);
not I_44605 (I761004,I760956);
nand I_44606 (I760701,I760767,I761004);
DFFARX1 I_44607 (I760956,I2683,I760724,I761044,);
not I_44608 (I761052,I761044);
not I_44609 (I761069,I872714);
not I_44610 (I761086,I872702);
nor I_44611 (I761103,I761086,I872705);
nor I_44612 (I760716,I761052,I761103);
nor I_44613 (I761134,I761086,I872708);
and I_44614 (I761151,I761134,I872717);
or I_44615 (I761168,I761151,I872705);
DFFARX1 I_44616 (I761168,I2683,I760724,I761194,);
nor I_44617 (I760704,I761194,I760750);
not I_44618 (I761216,I761194);
and I_44619 (I761233,I761216,I760750);
nor I_44620 (I760698,I760775,I761233);
nand I_44621 (I761264,I761216,I760826);
nor I_44622 (I760692,I761086,I761264);
nand I_44623 (I760695,I761216,I761004);
nand I_44624 (I761309,I760826,I872702);
nor I_44625 (I760707,I761069,I761309);
not I_44626 (I761370,I2690);
DFFARX1 I_44627 (I808561,I2683,I761370,I761396,);
DFFARX1 I_44628 (I808564,I2683,I761370,I761413,);
not I_44629 (I761421,I761413);
not I_44630 (I761438,I808561);
nor I_44631 (I761455,I761438,I808573);
not I_44632 (I761472,I808582);
nor I_44633 (I761489,I761455,I808570);
nor I_44634 (I761506,I761413,I761489);
DFFARX1 I_44635 (I761506,I2683,I761370,I761356,);
nor I_44636 (I761537,I808570,I808573);
nand I_44637 (I761554,I761537,I808561);
DFFARX1 I_44638 (I761554,I2683,I761370,I761359,);
nor I_44639 (I761585,I761472,I808570);
nand I_44640 (I761602,I761585,I808576);
nor I_44641 (I761619,I761396,I761602);
DFFARX1 I_44642 (I761619,I2683,I761370,I761335,);
not I_44643 (I761650,I761602);
nand I_44644 (I761347,I761413,I761650);
DFFARX1 I_44645 (I761602,I2683,I761370,I761690,);
not I_44646 (I761698,I761690);
not I_44647 (I761715,I808570);
not I_44648 (I761732,I808567);
nor I_44649 (I761749,I761732,I808582);
nor I_44650 (I761362,I761698,I761749);
nor I_44651 (I761780,I761732,I808579);
and I_44652 (I761797,I761780,I808567);
or I_44653 (I761814,I761797,I808564);
DFFARX1 I_44654 (I761814,I2683,I761370,I761840,);
nor I_44655 (I761350,I761840,I761396);
not I_44656 (I761862,I761840);
and I_44657 (I761879,I761862,I761396);
nor I_44658 (I761344,I761421,I761879);
nand I_44659 (I761910,I761862,I761472);
nor I_44660 (I761338,I761732,I761910);
nand I_44661 (I761341,I761862,I761650);
nand I_44662 (I761955,I761472,I808567);
nor I_44663 (I761353,I761715,I761955);
not I_44664 (I762016,I2690);
DFFARX1 I_44665 (I673383,I2683,I762016,I762042,);
DFFARX1 I_44666 (I673380,I2683,I762016,I762059,);
not I_44667 (I762067,I762059);
not I_44668 (I762084,I673380);
nor I_44669 (I762101,I762084,I673383);
not I_44670 (I762118,I673395);
nor I_44671 (I762135,I762101,I673389);
nor I_44672 (I762152,I762059,I762135);
DFFARX1 I_44673 (I762152,I2683,I762016,I762002,);
nor I_44674 (I762183,I673389,I673383);
nand I_44675 (I762200,I762183,I673380);
DFFARX1 I_44676 (I762200,I2683,I762016,I762005,);
nor I_44677 (I762231,I762118,I673389);
nand I_44678 (I762248,I762231,I673377);
nor I_44679 (I762265,I762042,I762248);
DFFARX1 I_44680 (I762265,I2683,I762016,I761981,);
not I_44681 (I762296,I762248);
nand I_44682 (I761993,I762059,I762296);
DFFARX1 I_44683 (I762248,I2683,I762016,I762336,);
not I_44684 (I762344,I762336);
not I_44685 (I762361,I673389);
not I_44686 (I762378,I673386);
nor I_44687 (I762395,I762378,I673395);
nor I_44688 (I762008,I762344,I762395);
nor I_44689 (I762426,I762378,I673392);
and I_44690 (I762443,I762426,I673398);
or I_44691 (I762460,I762443,I673377);
DFFARX1 I_44692 (I762460,I2683,I762016,I762486,);
nor I_44693 (I761996,I762486,I762042);
not I_44694 (I762508,I762486);
and I_44695 (I762525,I762508,I762042);
nor I_44696 (I761990,I762067,I762525);
nand I_44697 (I762556,I762508,I762118);
nor I_44698 (I761984,I762378,I762556);
nand I_44699 (I761987,I762508,I762296);
nand I_44700 (I762601,I762118,I673386);
nor I_44701 (I761999,I762361,I762601);
not I_44702 (I762662,I2690);
DFFARX1 I_44703 (I1031074,I2683,I762662,I762688,);
DFFARX1 I_44704 (I1031098,I2683,I762662,I762705,);
not I_44705 (I762713,I762705);
not I_44706 (I762730,I1031080);
nor I_44707 (I762747,I762730,I1031089);
not I_44708 (I762764,I1031074);
nor I_44709 (I762781,I762747,I1031095);
nor I_44710 (I762798,I762705,I762781);
DFFARX1 I_44711 (I762798,I2683,I762662,I762648,);
nor I_44712 (I762829,I1031095,I1031089);
nand I_44713 (I762846,I762829,I1031080);
DFFARX1 I_44714 (I762846,I2683,I762662,I762651,);
nor I_44715 (I762877,I762764,I1031095);
nand I_44716 (I762894,I762877,I1031092);
nor I_44717 (I762911,I762688,I762894);
DFFARX1 I_44718 (I762911,I2683,I762662,I762627,);
not I_44719 (I762942,I762894);
nand I_44720 (I762639,I762705,I762942);
DFFARX1 I_44721 (I762894,I2683,I762662,I762982,);
not I_44722 (I762990,I762982);
not I_44723 (I763007,I1031095);
not I_44724 (I763024,I1031086);
nor I_44725 (I763041,I763024,I1031074);
nor I_44726 (I762654,I762990,I763041);
nor I_44727 (I763072,I763024,I1031077);
and I_44728 (I763089,I763072,I1031101);
or I_44729 (I763106,I763089,I1031083);
DFFARX1 I_44730 (I763106,I2683,I762662,I763132,);
nor I_44731 (I762642,I763132,I762688);
not I_44732 (I763154,I763132);
and I_44733 (I763171,I763154,I762688);
nor I_44734 (I762636,I762713,I763171);
nand I_44735 (I763202,I763154,I762764);
nor I_44736 (I762630,I763024,I763202);
nand I_44737 (I762633,I763154,I762942);
nand I_44738 (I763247,I762764,I1031086);
nor I_44739 (I762645,I763007,I763247);
not I_44740 (I763308,I2690);
DFFARX1 I_44741 (I242206,I2683,I763308,I763334,);
DFFARX1 I_44742 (I242212,I2683,I763308,I763351,);
not I_44743 (I763359,I763351);
not I_44744 (I763376,I242233);
nor I_44745 (I763393,I763376,I242221);
not I_44746 (I763410,I242230);
nor I_44747 (I763427,I763393,I242215);
nor I_44748 (I763444,I763351,I763427);
DFFARX1 I_44749 (I763444,I2683,I763308,I763294,);
nor I_44750 (I763475,I242215,I242221);
nand I_44751 (I763492,I763475,I242233);
DFFARX1 I_44752 (I763492,I2683,I763308,I763297,);
nor I_44753 (I763523,I763410,I242215);
nand I_44754 (I763540,I763523,I242206);
nor I_44755 (I763557,I763334,I763540);
DFFARX1 I_44756 (I763557,I2683,I763308,I763273,);
not I_44757 (I763588,I763540);
nand I_44758 (I763285,I763351,I763588);
DFFARX1 I_44759 (I763540,I2683,I763308,I763628,);
not I_44760 (I763636,I763628);
not I_44761 (I763653,I242215);
not I_44762 (I763670,I242218);
nor I_44763 (I763687,I763670,I242230);
nor I_44764 (I763300,I763636,I763687);
nor I_44765 (I763718,I763670,I242227);
and I_44766 (I763735,I763718,I242209);
or I_44767 (I763752,I763735,I242224);
DFFARX1 I_44768 (I763752,I2683,I763308,I763778,);
nor I_44769 (I763288,I763778,I763334);
not I_44770 (I763800,I763778);
and I_44771 (I763817,I763800,I763334);
nor I_44772 (I763282,I763359,I763817);
nand I_44773 (I763848,I763800,I763410);
nor I_44774 (I763276,I763670,I763848);
nand I_44775 (I763279,I763800,I763588);
nand I_44776 (I763893,I763410,I242218);
nor I_44777 (I763291,I763653,I763893);
not I_44778 (I763954,I2690);
DFFARX1 I_44779 (I215329,I2683,I763954,I763980,);
DFFARX1 I_44780 (I215335,I2683,I763954,I763997,);
not I_44781 (I764005,I763997);
not I_44782 (I764022,I215356);
nor I_44783 (I764039,I764022,I215344);
not I_44784 (I764056,I215353);
nor I_44785 (I764073,I764039,I215338);
nor I_44786 (I764090,I763997,I764073);
DFFARX1 I_44787 (I764090,I2683,I763954,I763940,);
nor I_44788 (I764121,I215338,I215344);
nand I_44789 (I764138,I764121,I215356);
DFFARX1 I_44790 (I764138,I2683,I763954,I763943,);
nor I_44791 (I764169,I764056,I215338);
nand I_44792 (I764186,I764169,I215329);
nor I_44793 (I764203,I763980,I764186);
DFFARX1 I_44794 (I764203,I2683,I763954,I763919,);
not I_44795 (I764234,I764186);
nand I_44796 (I763931,I763997,I764234);
DFFARX1 I_44797 (I764186,I2683,I763954,I764274,);
not I_44798 (I764282,I764274);
not I_44799 (I764299,I215338);
not I_44800 (I764316,I215341);
nor I_44801 (I764333,I764316,I215353);
nor I_44802 (I763946,I764282,I764333);
nor I_44803 (I764364,I764316,I215350);
and I_44804 (I764381,I764364,I215332);
or I_44805 (I764398,I764381,I215347);
DFFARX1 I_44806 (I764398,I2683,I763954,I764424,);
nor I_44807 (I763934,I764424,I763980);
not I_44808 (I764446,I764424);
and I_44809 (I764463,I764446,I763980);
nor I_44810 (I763928,I764005,I764463);
nand I_44811 (I764494,I764446,I764056);
nor I_44812 (I763922,I764316,I764494);
nand I_44813 (I763925,I764446,I764234);
nand I_44814 (I764539,I764056,I215341);
nor I_44815 (I763937,I764299,I764539);
not I_44816 (I764600,I2690);
DFFARX1 I_44817 (I63791,I2683,I764600,I764626,);
DFFARX1 I_44818 (I63797,I2683,I764600,I764643,);
not I_44819 (I764651,I764643);
not I_44820 (I764668,I63815);
nor I_44821 (I764685,I764668,I63794);
not I_44822 (I764702,I63800);
nor I_44823 (I764719,I764685,I63806);
nor I_44824 (I764736,I764643,I764719);
DFFARX1 I_44825 (I764736,I2683,I764600,I764586,);
nor I_44826 (I764767,I63806,I63794);
nand I_44827 (I764784,I764767,I63815);
DFFARX1 I_44828 (I764784,I2683,I764600,I764589,);
nor I_44829 (I764815,I764702,I63806);
nand I_44830 (I764832,I764815,I63812);
nor I_44831 (I764849,I764626,I764832);
DFFARX1 I_44832 (I764849,I2683,I764600,I764565,);
not I_44833 (I764880,I764832);
nand I_44834 (I764577,I764643,I764880);
DFFARX1 I_44835 (I764832,I2683,I764600,I764920,);
not I_44836 (I764928,I764920);
not I_44837 (I764945,I63806);
not I_44838 (I764962,I63794);
nor I_44839 (I764979,I764962,I63800);
nor I_44840 (I764592,I764928,I764979);
nor I_44841 (I765010,I764962,I63803);
and I_44842 (I765027,I765010,I63791);
or I_44843 (I765044,I765027,I63809);
DFFARX1 I_44844 (I765044,I2683,I764600,I765070,);
nor I_44845 (I764580,I765070,I764626);
not I_44846 (I765092,I765070);
and I_44847 (I765109,I765092,I764626);
nor I_44848 (I764574,I764651,I765109);
nand I_44849 (I765140,I765092,I764702);
nor I_44850 (I764568,I764962,I765140);
nand I_44851 (I764571,I765092,I764880);
nand I_44852 (I765185,I764702,I63794);
nor I_44853 (I764583,I764945,I765185);
not I_44854 (I765246,I2690);
DFFARX1 I_44855 (I342648,I2683,I765246,I765272,);
DFFARX1 I_44856 (I342645,I2683,I765246,I765289,);
not I_44857 (I765297,I765289);
not I_44858 (I765314,I342660);
nor I_44859 (I765331,I765314,I342663);
not I_44860 (I765348,I342651);
nor I_44861 (I765365,I765331,I342657);
nor I_44862 (I765382,I765289,I765365);
DFFARX1 I_44863 (I765382,I2683,I765246,I765232,);
nor I_44864 (I765413,I342657,I342663);
nand I_44865 (I765430,I765413,I342660);
DFFARX1 I_44866 (I765430,I2683,I765246,I765235,);
nor I_44867 (I765461,I765348,I342657);
nand I_44868 (I765478,I765461,I342669);
nor I_44869 (I765495,I765272,I765478);
DFFARX1 I_44870 (I765495,I2683,I765246,I765211,);
not I_44871 (I765526,I765478);
nand I_44872 (I765223,I765289,I765526);
DFFARX1 I_44873 (I765478,I2683,I765246,I765566,);
not I_44874 (I765574,I765566);
not I_44875 (I765591,I342657);
not I_44876 (I765608,I342642);
nor I_44877 (I765625,I765608,I342651);
nor I_44878 (I765238,I765574,I765625);
nor I_44879 (I765656,I765608,I342654);
and I_44880 (I765673,I765656,I342642);
or I_44881 (I765690,I765673,I342666);
DFFARX1 I_44882 (I765690,I2683,I765246,I765716,);
nor I_44883 (I765226,I765716,I765272);
not I_44884 (I765738,I765716);
and I_44885 (I765755,I765738,I765272);
nor I_44886 (I765220,I765297,I765755);
nand I_44887 (I765786,I765738,I765348);
nor I_44888 (I765214,I765608,I765786);
nand I_44889 (I765217,I765738,I765526);
nand I_44890 (I765831,I765348,I342642);
nor I_44891 (I765229,I765591,I765831);
not I_44892 (I765892,I2690);
DFFARX1 I_44893 (I575752,I2683,I765892,I765918,);
DFFARX1 I_44894 (I575746,I2683,I765892,I765935,);
not I_44895 (I765943,I765935);
not I_44896 (I765960,I575761);
nor I_44897 (I765977,I765960,I575746);
not I_44898 (I765994,I575755);
nor I_44899 (I766011,I765977,I575764);
nor I_44900 (I766028,I765935,I766011);
DFFARX1 I_44901 (I766028,I2683,I765892,I765878,);
nor I_44902 (I766059,I575764,I575746);
nand I_44903 (I766076,I766059,I575761);
DFFARX1 I_44904 (I766076,I2683,I765892,I765881,);
nor I_44905 (I766107,I765994,I575764);
nand I_44906 (I766124,I766107,I575749);
nor I_44907 (I766141,I765918,I766124);
DFFARX1 I_44908 (I766141,I2683,I765892,I765857,);
not I_44909 (I766172,I766124);
nand I_44910 (I765869,I765935,I766172);
DFFARX1 I_44911 (I766124,I2683,I765892,I766212,);
not I_44912 (I766220,I766212);
not I_44913 (I766237,I575764);
not I_44914 (I766254,I575758);
nor I_44915 (I766271,I766254,I575755);
nor I_44916 (I765884,I766220,I766271);
nor I_44917 (I766302,I766254,I575767);
and I_44918 (I766319,I766302,I575770);
or I_44919 (I766336,I766319,I575749);
DFFARX1 I_44920 (I766336,I2683,I765892,I766362,);
nor I_44921 (I765872,I766362,I765918);
not I_44922 (I766384,I766362);
and I_44923 (I766401,I766384,I765918);
nor I_44924 (I765866,I765943,I766401);
nand I_44925 (I766432,I766384,I765994);
nor I_44926 (I765860,I766254,I766432);
nand I_44927 (I765863,I766384,I766172);
nand I_44928 (I766477,I765994,I575758);
nor I_44929 (I765875,I766237,I766477);
not I_44930 (I766538,I2690);
DFFARX1 I_44931 (I893528,I2683,I766538,I766564,);
DFFARX1 I_44932 (I893510,I2683,I766538,I766581,);
not I_44933 (I766589,I766581);
not I_44934 (I766606,I893519);
nor I_44935 (I766623,I766606,I893531);
not I_44936 (I766640,I893513);
nor I_44937 (I766657,I766623,I893522);
nor I_44938 (I766674,I766581,I766657);
DFFARX1 I_44939 (I766674,I2683,I766538,I766524,);
nor I_44940 (I766705,I893522,I893531);
nand I_44941 (I766722,I766705,I893519);
DFFARX1 I_44942 (I766722,I2683,I766538,I766527,);
nor I_44943 (I766753,I766640,I893522);
nand I_44944 (I766770,I766753,I893534);
nor I_44945 (I766787,I766564,I766770);
DFFARX1 I_44946 (I766787,I2683,I766538,I766503,);
not I_44947 (I766818,I766770);
nand I_44948 (I766515,I766581,I766818);
DFFARX1 I_44949 (I766770,I2683,I766538,I766858,);
not I_44950 (I766866,I766858);
not I_44951 (I766883,I893522);
not I_44952 (I766900,I893510);
nor I_44953 (I766917,I766900,I893513);
nor I_44954 (I766530,I766866,I766917);
nor I_44955 (I766948,I766900,I893516);
and I_44956 (I766965,I766948,I893525);
or I_44957 (I766982,I766965,I893513);
DFFARX1 I_44958 (I766982,I2683,I766538,I767008,);
nor I_44959 (I766518,I767008,I766564);
not I_44960 (I767030,I767008);
and I_44961 (I767047,I767030,I766564);
nor I_44962 (I766512,I766589,I767047);
nand I_44963 (I767078,I767030,I766640);
nor I_44964 (I766506,I766900,I767078);
nand I_44965 (I766509,I767030,I766818);
nand I_44966 (I767123,I766640,I893510);
nor I_44967 (I766521,I766883,I767123);
not I_44968 (I767184,I2690);
DFFARX1 I_44969 (I1071534,I2683,I767184,I767210,);
DFFARX1 I_44970 (I1071558,I2683,I767184,I767227,);
not I_44971 (I767235,I767227);
not I_44972 (I767252,I1071540);
nor I_44973 (I767269,I767252,I1071549);
not I_44974 (I767286,I1071534);
nor I_44975 (I767303,I767269,I1071555);
nor I_44976 (I767320,I767227,I767303);
DFFARX1 I_44977 (I767320,I2683,I767184,I767170,);
nor I_44978 (I767351,I1071555,I1071549);
nand I_44979 (I767368,I767351,I1071540);
DFFARX1 I_44980 (I767368,I2683,I767184,I767173,);
nor I_44981 (I767399,I767286,I1071555);
nand I_44982 (I767416,I767399,I1071552);
nor I_44983 (I767433,I767210,I767416);
DFFARX1 I_44984 (I767433,I2683,I767184,I767149,);
not I_44985 (I767464,I767416);
nand I_44986 (I767161,I767227,I767464);
DFFARX1 I_44987 (I767416,I2683,I767184,I767504,);
not I_44988 (I767512,I767504);
not I_44989 (I767529,I1071555);
not I_44990 (I767546,I1071546);
nor I_44991 (I767563,I767546,I1071534);
nor I_44992 (I767176,I767512,I767563);
nor I_44993 (I767594,I767546,I1071537);
and I_44994 (I767611,I767594,I1071561);
or I_44995 (I767628,I767611,I1071543);
DFFARX1 I_44996 (I767628,I2683,I767184,I767654,);
nor I_44997 (I767164,I767654,I767210);
not I_44998 (I767676,I767654);
and I_44999 (I767693,I767676,I767210);
nor I_45000 (I767158,I767235,I767693);
nand I_45001 (I767724,I767676,I767286);
nor I_45002 (I767152,I767546,I767724);
nand I_45003 (I767155,I767676,I767464);
nand I_45004 (I767769,I767286,I1071546);
nor I_45005 (I767167,I767529,I767769);
not I_45006 (I767830,I2690);
DFFARX1 I_45007 (I810805,I2683,I767830,I767856,);
DFFARX1 I_45008 (I810808,I2683,I767830,I767873,);
not I_45009 (I767881,I767873);
not I_45010 (I767898,I810805);
nor I_45011 (I767915,I767898,I810817);
not I_45012 (I767932,I810826);
nor I_45013 (I767949,I767915,I810814);
nor I_45014 (I767966,I767873,I767949);
DFFARX1 I_45015 (I767966,I2683,I767830,I767816,);
nor I_45016 (I767997,I810814,I810817);
nand I_45017 (I768014,I767997,I810805);
DFFARX1 I_45018 (I768014,I2683,I767830,I767819,);
nor I_45019 (I768045,I767932,I810814);
nand I_45020 (I768062,I768045,I810820);
nor I_45021 (I768079,I767856,I768062);
DFFARX1 I_45022 (I768079,I2683,I767830,I767795,);
not I_45023 (I768110,I768062);
nand I_45024 (I767807,I767873,I768110);
DFFARX1 I_45025 (I768062,I2683,I767830,I768150,);
not I_45026 (I768158,I768150);
not I_45027 (I768175,I810814);
not I_45028 (I768192,I810811);
nor I_45029 (I768209,I768192,I810826);
nor I_45030 (I767822,I768158,I768209);
nor I_45031 (I768240,I768192,I810823);
and I_45032 (I768257,I768240,I810811);
or I_45033 (I768274,I768257,I810808);
DFFARX1 I_45034 (I768274,I2683,I767830,I768300,);
nor I_45035 (I767810,I768300,I767856);
not I_45036 (I768322,I768300);
and I_45037 (I768339,I768322,I767856);
nor I_45038 (I767804,I767881,I768339);
nand I_45039 (I768370,I768322,I767932);
nor I_45040 (I767798,I768192,I768370);
nand I_45041 (I767801,I768322,I768110);
nand I_45042 (I768415,I767932,I810811);
nor I_45043 (I767813,I768175,I768415);
not I_45044 (I768476,I2690);
DFFARX1 I_45045 (I216383,I2683,I768476,I768502,);
DFFARX1 I_45046 (I216389,I2683,I768476,I768519,);
not I_45047 (I768527,I768519);
not I_45048 (I768544,I216410);
nor I_45049 (I768561,I768544,I216398);
not I_45050 (I768578,I216407);
nor I_45051 (I768595,I768561,I216392);
nor I_45052 (I768612,I768519,I768595);
DFFARX1 I_45053 (I768612,I2683,I768476,I768462,);
nor I_45054 (I768643,I216392,I216398);
nand I_45055 (I768660,I768643,I216410);
DFFARX1 I_45056 (I768660,I2683,I768476,I768465,);
nor I_45057 (I768691,I768578,I216392);
nand I_45058 (I768708,I768691,I216383);
nor I_45059 (I768725,I768502,I768708);
DFFARX1 I_45060 (I768725,I2683,I768476,I768441,);
not I_45061 (I768756,I768708);
nand I_45062 (I768453,I768519,I768756);
DFFARX1 I_45063 (I768708,I2683,I768476,I768796,);
not I_45064 (I768804,I768796);
not I_45065 (I768821,I216392);
not I_45066 (I768838,I216395);
nor I_45067 (I768855,I768838,I216407);
nor I_45068 (I768468,I768804,I768855);
nor I_45069 (I768886,I768838,I216404);
and I_45070 (I768903,I768886,I216386);
or I_45071 (I768920,I768903,I216401);
DFFARX1 I_45072 (I768920,I2683,I768476,I768946,);
nor I_45073 (I768456,I768946,I768502);
not I_45074 (I768968,I768946);
and I_45075 (I768985,I768968,I768502);
nor I_45076 (I768450,I768527,I768985);
nand I_45077 (I769016,I768968,I768578);
nor I_45078 (I768444,I768838,I769016);
nand I_45079 (I768447,I768968,I768756);
nand I_45080 (I769061,I768578,I216395);
nor I_45081 (I768459,I768821,I769061);
not I_45082 (I769122,I2690);
DFFARX1 I_45083 (I644398,I2683,I769122,I769148,);
DFFARX1 I_45084 (I644395,I2683,I769122,I769165,);
not I_45085 (I769173,I769165);
not I_45086 (I769190,I644395);
nor I_45087 (I769207,I769190,I644398);
not I_45088 (I769224,I644410);
nor I_45089 (I769241,I769207,I644404);
nor I_45090 (I769258,I769165,I769241);
DFFARX1 I_45091 (I769258,I2683,I769122,I769108,);
nor I_45092 (I769289,I644404,I644398);
nand I_45093 (I769306,I769289,I644395);
DFFARX1 I_45094 (I769306,I2683,I769122,I769111,);
nor I_45095 (I769337,I769224,I644404);
nand I_45096 (I769354,I769337,I644392);
nor I_45097 (I769371,I769148,I769354);
DFFARX1 I_45098 (I769371,I2683,I769122,I769087,);
not I_45099 (I769402,I769354);
nand I_45100 (I769099,I769165,I769402);
DFFARX1 I_45101 (I769354,I2683,I769122,I769442,);
not I_45102 (I769450,I769442);
not I_45103 (I769467,I644404);
not I_45104 (I769484,I644401);
nor I_45105 (I769501,I769484,I644410);
nor I_45106 (I769114,I769450,I769501);
nor I_45107 (I769532,I769484,I644407);
and I_45108 (I769549,I769532,I644413);
or I_45109 (I769566,I769549,I644392);
DFFARX1 I_45110 (I769566,I2683,I769122,I769592,);
nor I_45111 (I769102,I769592,I769148);
not I_45112 (I769614,I769592);
and I_45113 (I769631,I769614,I769148);
nor I_45114 (I769096,I769173,I769631);
nand I_45115 (I769662,I769614,I769224);
nor I_45116 (I769090,I769484,I769662);
nand I_45117 (I769093,I769614,I769402);
nand I_45118 (I769707,I769224,I644401);
nor I_45119 (I769105,I769467,I769707);
not I_45120 (I769768,I2690);
DFFARX1 I_45121 (I467663,I2683,I769768,I769794,);
DFFARX1 I_45122 (I467675,I2683,I769768,I769811,);
not I_45123 (I769819,I769811);
not I_45124 (I769836,I467684);
nor I_45125 (I769853,I769836,I467660);
not I_45126 (I769870,I467678);
nor I_45127 (I769887,I769853,I467672);
nor I_45128 (I769904,I769811,I769887);
DFFARX1 I_45129 (I769904,I2683,I769768,I769754,);
nor I_45130 (I769935,I467672,I467660);
nand I_45131 (I769952,I769935,I467684);
DFFARX1 I_45132 (I769952,I2683,I769768,I769757,);
nor I_45133 (I769983,I769870,I467672);
nand I_45134 (I770000,I769983,I467666);
nor I_45135 (I770017,I769794,I770000);
DFFARX1 I_45136 (I770017,I2683,I769768,I769733,);
not I_45137 (I770048,I770000);
nand I_45138 (I769745,I769811,I770048);
DFFARX1 I_45139 (I770000,I2683,I769768,I770088,);
not I_45140 (I770096,I770088);
not I_45141 (I770113,I467672);
not I_45142 (I770130,I467681);
nor I_45143 (I770147,I770130,I467678);
nor I_45144 (I769760,I770096,I770147);
nor I_45145 (I770178,I770130,I467663);
and I_45146 (I770195,I770178,I467660);
or I_45147 (I770212,I770195,I467669);
DFFARX1 I_45148 (I770212,I2683,I769768,I770238,);
nor I_45149 (I769748,I770238,I769794);
not I_45150 (I770260,I770238);
and I_45151 (I770277,I770260,I769794);
nor I_45152 (I769742,I769819,I770277);
nand I_45153 (I770308,I770260,I769870);
nor I_45154 (I769736,I770130,I770308);
nand I_45155 (I769739,I770260,I770048);
nand I_45156 (I770353,I769870,I467681);
nor I_45157 (I769751,I770113,I770353);
not I_45158 (I770414,I2690);
DFFARX1 I_45159 (I1072724,I2683,I770414,I770440,);
DFFARX1 I_45160 (I1072748,I2683,I770414,I770457,);
not I_45161 (I770465,I770457);
not I_45162 (I770482,I1072730);
nor I_45163 (I770499,I770482,I1072739);
not I_45164 (I770516,I1072724);
nor I_45165 (I770533,I770499,I1072745);
nor I_45166 (I770550,I770457,I770533);
DFFARX1 I_45167 (I770550,I2683,I770414,I770400,);
nor I_45168 (I770581,I1072745,I1072739);
nand I_45169 (I770598,I770581,I1072730);
DFFARX1 I_45170 (I770598,I2683,I770414,I770403,);
nor I_45171 (I770629,I770516,I1072745);
nand I_45172 (I770646,I770629,I1072742);
nor I_45173 (I770663,I770440,I770646);
DFFARX1 I_45174 (I770663,I2683,I770414,I770379,);
not I_45175 (I770694,I770646);
nand I_45176 (I770391,I770457,I770694);
DFFARX1 I_45177 (I770646,I2683,I770414,I770734,);
not I_45178 (I770742,I770734);
not I_45179 (I770759,I1072745);
not I_45180 (I770776,I1072736);
nor I_45181 (I770793,I770776,I1072724);
nor I_45182 (I770406,I770742,I770793);
nor I_45183 (I770824,I770776,I1072727);
and I_45184 (I770841,I770824,I1072751);
or I_45185 (I770858,I770841,I1072733);
DFFARX1 I_45186 (I770858,I2683,I770414,I770884,);
nor I_45187 (I770394,I770884,I770440);
not I_45188 (I770906,I770884);
and I_45189 (I770923,I770906,I770440);
nor I_45190 (I770388,I770465,I770923);
nand I_45191 (I770954,I770906,I770516);
nor I_45192 (I770382,I770776,I770954);
nand I_45193 (I770385,I770906,I770694);
nand I_45194 (I770999,I770516,I1072736);
nor I_45195 (I770397,I770759,I770999);
not I_45196 (I771060,I2690);
DFFARX1 I_45197 (I1019217,I2683,I771060,I771086,);
DFFARX1 I_45198 (I1019211,I2683,I771060,I771103,);
not I_45199 (I771111,I771103);
not I_45200 (I771128,I1019220);
nor I_45201 (I771145,I771128,I1019232);
not I_45202 (I771162,I1019214);
nor I_45203 (I771179,I771145,I1019211);
nor I_45204 (I771196,I771103,I771179);
DFFARX1 I_45205 (I771196,I2683,I771060,I771046,);
nor I_45206 (I771227,I1019211,I1019232);
nand I_45207 (I771244,I771227,I1019220);
DFFARX1 I_45208 (I771244,I2683,I771060,I771049,);
nor I_45209 (I771275,I771162,I1019211);
nand I_45210 (I771292,I771275,I1019208);
nor I_45211 (I771309,I771086,I771292);
DFFARX1 I_45212 (I771309,I2683,I771060,I771025,);
not I_45213 (I771340,I771292);
nand I_45214 (I771037,I771103,I771340);
DFFARX1 I_45215 (I771292,I2683,I771060,I771380,);
not I_45216 (I771388,I771380);
not I_45217 (I771405,I1019211);
not I_45218 (I771422,I1019229);
nor I_45219 (I771439,I771422,I1019214);
nor I_45220 (I771052,I771388,I771439);
nor I_45221 (I771470,I771422,I1019223);
and I_45222 (I771487,I771470,I1019208);
or I_45223 (I771504,I771487,I1019226);
DFFARX1 I_45224 (I771504,I2683,I771060,I771530,);
nor I_45225 (I771040,I771530,I771086);
not I_45226 (I771552,I771530);
and I_45227 (I771569,I771552,I771086);
nor I_45228 (I771034,I771111,I771569);
nand I_45229 (I771600,I771552,I771162);
nor I_45230 (I771028,I771422,I771600);
nand I_45231 (I771031,I771552,I771340);
nand I_45232 (I771645,I771162,I1019229);
nor I_45233 (I771043,I771405,I771645);
not I_45234 (I771706,I2690);
DFFARX1 I_45235 (I457837,I2683,I771706,I771732,);
DFFARX1 I_45236 (I457849,I2683,I771706,I771749,);
not I_45237 (I771757,I771749);
not I_45238 (I771774,I457858);
nor I_45239 (I771791,I771774,I457834);
not I_45240 (I771808,I457852);
nor I_45241 (I771825,I771791,I457846);
nor I_45242 (I771842,I771749,I771825);
DFFARX1 I_45243 (I771842,I2683,I771706,I771692,);
nor I_45244 (I771873,I457846,I457834);
nand I_45245 (I771890,I771873,I457858);
DFFARX1 I_45246 (I771890,I2683,I771706,I771695,);
nor I_45247 (I771921,I771808,I457846);
nand I_45248 (I771938,I771921,I457840);
nor I_45249 (I771955,I771732,I771938);
DFFARX1 I_45250 (I771955,I2683,I771706,I771671,);
not I_45251 (I771986,I771938);
nand I_45252 (I771683,I771749,I771986);
DFFARX1 I_45253 (I771938,I2683,I771706,I772026,);
not I_45254 (I772034,I772026);
not I_45255 (I772051,I457846);
not I_45256 (I772068,I457855);
nor I_45257 (I772085,I772068,I457852);
nor I_45258 (I771698,I772034,I772085);
nor I_45259 (I772116,I772068,I457837);
and I_45260 (I772133,I772116,I457834);
or I_45261 (I772150,I772133,I457843);
DFFARX1 I_45262 (I772150,I2683,I771706,I772176,);
nor I_45263 (I771686,I772176,I771732);
not I_45264 (I772198,I772176);
and I_45265 (I772215,I772198,I771732);
nor I_45266 (I771680,I771757,I772215);
nand I_45267 (I772246,I772198,I771808);
nor I_45268 (I771674,I772068,I772246);
nand I_45269 (I771677,I772198,I771986);
nand I_45270 (I772291,I771808,I457855);
nor I_45271 (I771689,I772051,I772291);
not I_45272 (I772352,I2690);
DFFARX1 I_45273 (I327416,I2683,I772352,I772378,);
DFFARX1 I_45274 (I327413,I2683,I772352,I772395,);
not I_45275 (I772403,I772395);
not I_45276 (I772420,I327428);
nor I_45277 (I772437,I772420,I327431);
not I_45278 (I772454,I327419);
nor I_45279 (I772471,I772437,I327425);
nor I_45280 (I772488,I772395,I772471);
DFFARX1 I_45281 (I772488,I2683,I772352,I772338,);
nor I_45282 (I772519,I327425,I327431);
nand I_45283 (I772536,I772519,I327428);
DFFARX1 I_45284 (I772536,I2683,I772352,I772341,);
nor I_45285 (I772567,I772454,I327425);
nand I_45286 (I772584,I772567,I327437);
nor I_45287 (I772601,I772378,I772584);
DFFARX1 I_45288 (I772601,I2683,I772352,I772317,);
not I_45289 (I772632,I772584);
nand I_45290 (I772329,I772395,I772632);
DFFARX1 I_45291 (I772584,I2683,I772352,I772672,);
not I_45292 (I772680,I772672);
not I_45293 (I772697,I327425);
not I_45294 (I772714,I327410);
nor I_45295 (I772731,I772714,I327419);
nor I_45296 (I772344,I772680,I772731);
nor I_45297 (I772762,I772714,I327422);
and I_45298 (I772779,I772762,I327410);
or I_45299 (I772796,I772779,I327434);
DFFARX1 I_45300 (I772796,I2683,I772352,I772822,);
nor I_45301 (I772332,I772822,I772378);
not I_45302 (I772844,I772822);
and I_45303 (I772861,I772844,I772378);
nor I_45304 (I772326,I772403,I772861);
nand I_45305 (I772892,I772844,I772454);
nor I_45306 (I772320,I772714,I772892);
nand I_45307 (I772323,I772844,I772632);
nand I_45308 (I772937,I772454,I327410);
nor I_45309 (I772335,I772697,I772937);
not I_45310 (I772998,I2690);
DFFARX1 I_45311 (I1034049,I2683,I772998,I773024,);
DFFARX1 I_45312 (I1034073,I2683,I772998,I773041,);
not I_45313 (I773049,I773041);
not I_45314 (I773066,I1034055);
nor I_45315 (I773083,I773066,I1034064);
not I_45316 (I773100,I1034049);
nor I_45317 (I773117,I773083,I1034070);
nor I_45318 (I773134,I773041,I773117);
DFFARX1 I_45319 (I773134,I2683,I772998,I772984,);
nor I_45320 (I773165,I1034070,I1034064);
nand I_45321 (I773182,I773165,I1034055);
DFFARX1 I_45322 (I773182,I2683,I772998,I772987,);
nor I_45323 (I773213,I773100,I1034070);
nand I_45324 (I773230,I773213,I1034067);
nor I_45325 (I773247,I773024,I773230);
DFFARX1 I_45326 (I773247,I2683,I772998,I772963,);
not I_45327 (I773278,I773230);
nand I_45328 (I772975,I773041,I773278);
DFFARX1 I_45329 (I773230,I2683,I772998,I773318,);
not I_45330 (I773326,I773318);
not I_45331 (I773343,I1034070);
not I_45332 (I773360,I1034061);
nor I_45333 (I773377,I773360,I1034049);
nor I_45334 (I772990,I773326,I773377);
nor I_45335 (I773408,I773360,I1034052);
and I_45336 (I773425,I773408,I1034076);
or I_45337 (I773442,I773425,I1034058);
DFFARX1 I_45338 (I773442,I2683,I772998,I773468,);
nor I_45339 (I772978,I773468,I773024);
not I_45340 (I773490,I773468);
and I_45341 (I773507,I773490,I773024);
nor I_45342 (I772972,I773049,I773507);
nand I_45343 (I773538,I773490,I773100);
nor I_45344 (I772966,I773360,I773538);
nand I_45345 (I772969,I773490,I773278);
nand I_45346 (I773583,I773100,I1034061);
nor I_45347 (I772981,I773343,I773583);
not I_45348 (I773644,I2690);
DFFARX1 I_45349 (I616212,I2683,I773644,I773670,);
DFFARX1 I_45350 (I616206,I2683,I773644,I773687,);
not I_45351 (I773695,I773687);
not I_45352 (I773712,I616221);
nor I_45353 (I773729,I773712,I616206);
not I_45354 (I773746,I616215);
nor I_45355 (I773763,I773729,I616224);
nor I_45356 (I773780,I773687,I773763);
DFFARX1 I_45357 (I773780,I2683,I773644,I773630,);
nor I_45358 (I773811,I616224,I616206);
nand I_45359 (I773828,I773811,I616221);
DFFARX1 I_45360 (I773828,I2683,I773644,I773633,);
nor I_45361 (I773859,I773746,I616224);
nand I_45362 (I773876,I773859,I616209);
nor I_45363 (I773893,I773670,I773876);
DFFARX1 I_45364 (I773893,I2683,I773644,I773609,);
not I_45365 (I773924,I773876);
nand I_45366 (I773621,I773687,I773924);
DFFARX1 I_45367 (I773876,I2683,I773644,I773964,);
not I_45368 (I773972,I773964);
not I_45369 (I773989,I616224);
not I_45370 (I774006,I616218);
nor I_45371 (I774023,I774006,I616215);
nor I_45372 (I773636,I773972,I774023);
nor I_45373 (I774054,I774006,I616227);
and I_45374 (I774071,I774054,I616230);
or I_45375 (I774088,I774071,I616209);
DFFARX1 I_45376 (I774088,I2683,I773644,I774114,);
nor I_45377 (I773624,I774114,I773670);
not I_45378 (I774136,I774114);
and I_45379 (I774153,I774136,I773670);
nor I_45380 (I773618,I773695,I774153);
nand I_45381 (I774184,I774136,I773746);
nor I_45382 (I773612,I774006,I774184);
nand I_45383 (I773615,I774136,I773924);
nand I_45384 (I774229,I773746,I616218);
nor I_45385 (I773627,I773989,I774229);
not I_45386 (I774290,I2690);
DFFARX1 I_45387 (I656519,I2683,I774290,I774316,);
DFFARX1 I_45388 (I656516,I2683,I774290,I774333,);
not I_45389 (I774341,I774333);
not I_45390 (I774358,I656516);
nor I_45391 (I774375,I774358,I656519);
not I_45392 (I774392,I656531);
nor I_45393 (I774409,I774375,I656525);
nor I_45394 (I774426,I774333,I774409);
DFFARX1 I_45395 (I774426,I2683,I774290,I774276,);
nor I_45396 (I774457,I656525,I656519);
nand I_45397 (I774474,I774457,I656516);
DFFARX1 I_45398 (I774474,I2683,I774290,I774279,);
nor I_45399 (I774505,I774392,I656525);
nand I_45400 (I774522,I774505,I656513);
nor I_45401 (I774539,I774316,I774522);
DFFARX1 I_45402 (I774539,I2683,I774290,I774255,);
not I_45403 (I774570,I774522);
nand I_45404 (I774267,I774333,I774570);
DFFARX1 I_45405 (I774522,I2683,I774290,I774610,);
not I_45406 (I774618,I774610);
not I_45407 (I774635,I656525);
not I_45408 (I774652,I656522);
nor I_45409 (I774669,I774652,I656531);
nor I_45410 (I774282,I774618,I774669);
nor I_45411 (I774700,I774652,I656528);
and I_45412 (I774717,I774700,I656534);
or I_45413 (I774734,I774717,I656513);
DFFARX1 I_45414 (I774734,I2683,I774290,I774760,);
nor I_45415 (I774270,I774760,I774316);
not I_45416 (I774782,I774760);
and I_45417 (I774799,I774782,I774316);
nor I_45418 (I774264,I774341,I774799);
nand I_45419 (I774830,I774782,I774392);
nor I_45420 (I774258,I774652,I774830);
nand I_45421 (I774261,I774782,I774570);
nand I_45422 (I774875,I774392,I656522);
nor I_45423 (I774273,I774635,I774875);
not I_45424 (I774936,I2690);
DFFARX1 I_45425 (I1022079,I2683,I774936,I774962,);
DFFARX1 I_45426 (I1022076,I2683,I774936,I774979,);
not I_45427 (I774987,I774979);
not I_45428 (I775004,I1022073);
nor I_45429 (I775021,I775004,I1022064);
not I_45430 (I775038,I1022085);
nor I_45431 (I775055,I775021,I1022064);
nor I_45432 (I775072,I774979,I775055);
DFFARX1 I_45433 (I775072,I2683,I774936,I774922,);
nor I_45434 (I775103,I1022064,I1022064);
nand I_45435 (I775120,I775103,I1022073);
DFFARX1 I_45436 (I775120,I2683,I774936,I774925,);
nor I_45437 (I775151,I775038,I1022064);
nand I_45438 (I775168,I775151,I1022088);
nor I_45439 (I775185,I774962,I775168);
DFFARX1 I_45440 (I775185,I2683,I774936,I774901,);
not I_45441 (I775216,I775168);
nand I_45442 (I774913,I774979,I775216);
DFFARX1 I_45443 (I775168,I2683,I774936,I775256,);
not I_45444 (I775264,I775256);
not I_45445 (I775281,I1022064);
not I_45446 (I775298,I1022067);
nor I_45447 (I775315,I775298,I1022085);
nor I_45448 (I774928,I775264,I775315);
nor I_45449 (I775346,I775298,I1022070);
and I_45450 (I775363,I775346,I1022091);
or I_45451 (I775380,I775363,I1022082);
DFFARX1 I_45452 (I775380,I2683,I774936,I775406,);
nor I_45453 (I774916,I775406,I774962);
not I_45454 (I775428,I775406);
and I_45455 (I775445,I775428,I774962);
nor I_45456 (I774910,I774987,I775445);
nand I_45457 (I775476,I775428,I775038);
nor I_45458 (I774904,I775298,I775476);
nand I_45459 (I774907,I775428,I775216);
nand I_45460 (I775521,I775038,I1022067);
nor I_45461 (I774919,I775281,I775521);
not I_45462 (I775582,I2690);
DFFARX1 I_45463 (I929364,I2683,I775582,I775608,);
DFFARX1 I_45464 (I929346,I2683,I775582,I775625,);
not I_45465 (I775633,I775625);
not I_45466 (I775650,I929355);
nor I_45467 (I775667,I775650,I929367);
not I_45468 (I775684,I929349);
nor I_45469 (I775701,I775667,I929358);
nor I_45470 (I775718,I775625,I775701);
DFFARX1 I_45471 (I775718,I2683,I775582,I775568,);
nor I_45472 (I775749,I929358,I929367);
nand I_45473 (I775766,I775749,I929355);
DFFARX1 I_45474 (I775766,I2683,I775582,I775571,);
nor I_45475 (I775797,I775684,I929358);
nand I_45476 (I775814,I775797,I929370);
nor I_45477 (I775831,I775608,I775814);
DFFARX1 I_45478 (I775831,I2683,I775582,I775547,);
not I_45479 (I775862,I775814);
nand I_45480 (I775559,I775625,I775862);
DFFARX1 I_45481 (I775814,I2683,I775582,I775902,);
not I_45482 (I775910,I775902);
not I_45483 (I775927,I929358);
not I_45484 (I775944,I929346);
nor I_45485 (I775961,I775944,I929349);
nor I_45486 (I775574,I775910,I775961);
nor I_45487 (I775992,I775944,I929352);
and I_45488 (I776009,I775992,I929361);
or I_45489 (I776026,I776009,I929349);
DFFARX1 I_45490 (I776026,I2683,I775582,I776052,);
nor I_45491 (I775562,I776052,I775608);
not I_45492 (I776074,I776052);
and I_45493 (I776091,I776074,I775608);
nor I_45494 (I775556,I775633,I776091);
nand I_45495 (I776122,I776074,I775684);
nor I_45496 (I775550,I775944,I776122);
nand I_45497 (I775553,I776074,I775862);
nand I_45498 (I776167,I775684,I929346);
nor I_45499 (I775565,I775927,I776167);
not I_45500 (I776228,I2690);
DFFARX1 I_45501 (I590780,I2683,I776228,I776254,);
DFFARX1 I_45502 (I590774,I2683,I776228,I776271,);
not I_45503 (I776279,I776271);
not I_45504 (I776296,I590789);
nor I_45505 (I776313,I776296,I590774);
not I_45506 (I776330,I590783);
nor I_45507 (I776347,I776313,I590792);
nor I_45508 (I776364,I776271,I776347);
DFFARX1 I_45509 (I776364,I2683,I776228,I776214,);
nor I_45510 (I776395,I590792,I590774);
nand I_45511 (I776412,I776395,I590789);
DFFARX1 I_45512 (I776412,I2683,I776228,I776217,);
nor I_45513 (I776443,I776330,I590792);
nand I_45514 (I776460,I776443,I590777);
nor I_45515 (I776477,I776254,I776460);
DFFARX1 I_45516 (I776477,I2683,I776228,I776193,);
not I_45517 (I776508,I776460);
nand I_45518 (I776205,I776271,I776508);
DFFARX1 I_45519 (I776460,I2683,I776228,I776548,);
not I_45520 (I776556,I776548);
not I_45521 (I776573,I590792);
not I_45522 (I776590,I590786);
nor I_45523 (I776607,I776590,I590783);
nor I_45524 (I776220,I776556,I776607);
nor I_45525 (I776638,I776590,I590795);
and I_45526 (I776655,I776638,I590798);
or I_45527 (I776672,I776655,I590777);
DFFARX1 I_45528 (I776672,I2683,I776228,I776698,);
nor I_45529 (I776208,I776698,I776254);
not I_45530 (I776720,I776698);
and I_45531 (I776737,I776720,I776254);
nor I_45532 (I776202,I776279,I776737);
nand I_45533 (I776768,I776720,I776330);
nor I_45534 (I776196,I776590,I776768);
nand I_45535 (I776199,I776720,I776508);
nand I_45536 (I776813,I776330,I590786);
nor I_45537 (I776211,I776573,I776813);
not I_45538 (I776874,I2690);
DFFARX1 I_45539 (I609854,I2683,I776874,I776900,);
DFFARX1 I_45540 (I609848,I2683,I776874,I776917,);
not I_45541 (I776925,I776917);
not I_45542 (I776942,I609863);
nor I_45543 (I776959,I776942,I609848);
not I_45544 (I776976,I609857);
nor I_45545 (I776993,I776959,I609866);
nor I_45546 (I777010,I776917,I776993);
DFFARX1 I_45547 (I777010,I2683,I776874,I776860,);
nor I_45548 (I777041,I609866,I609848);
nand I_45549 (I777058,I777041,I609863);
DFFARX1 I_45550 (I777058,I2683,I776874,I776863,);
nor I_45551 (I777089,I776976,I609866);
nand I_45552 (I777106,I777089,I609851);
nor I_45553 (I777123,I776900,I777106);
DFFARX1 I_45554 (I777123,I2683,I776874,I776839,);
not I_45555 (I777154,I777106);
nand I_45556 (I776851,I776917,I777154);
DFFARX1 I_45557 (I777106,I2683,I776874,I777194,);
not I_45558 (I777202,I777194);
not I_45559 (I777219,I609866);
not I_45560 (I777236,I609860);
nor I_45561 (I777253,I777236,I609857);
nor I_45562 (I776866,I777202,I777253);
nor I_45563 (I777284,I777236,I609869);
and I_45564 (I777301,I777284,I609872);
or I_45565 (I777318,I777301,I609851);
DFFARX1 I_45566 (I777318,I2683,I776874,I777344,);
nor I_45567 (I776854,I777344,I776900);
not I_45568 (I777366,I777344);
and I_45569 (I777383,I777366,I776900);
nor I_45570 (I776848,I776925,I777383);
nand I_45571 (I777414,I777366,I776976);
nor I_45572 (I776842,I777236,I777414);
nand I_45573 (I776845,I777366,I777154);
nand I_45574 (I777459,I776976,I609860);
nor I_45575 (I776857,I777219,I777459);
not I_45576 (I777520,I2690);
DFFARX1 I_45577 (I251692,I2683,I777520,I777546,);
DFFARX1 I_45578 (I251698,I2683,I777520,I777563,);
not I_45579 (I777571,I777563);
not I_45580 (I777588,I251719);
nor I_45581 (I777605,I777588,I251707);
not I_45582 (I777622,I251716);
nor I_45583 (I777639,I777605,I251701);
nor I_45584 (I777656,I777563,I777639);
DFFARX1 I_45585 (I777656,I2683,I777520,I777506,);
nor I_45586 (I777687,I251701,I251707);
nand I_45587 (I777704,I777687,I251719);
DFFARX1 I_45588 (I777704,I2683,I777520,I777509,);
nor I_45589 (I777735,I777622,I251701);
nand I_45590 (I777752,I777735,I251692);
nor I_45591 (I777769,I777546,I777752);
DFFARX1 I_45592 (I777769,I2683,I777520,I777485,);
not I_45593 (I777800,I777752);
nand I_45594 (I777497,I777563,I777800);
DFFARX1 I_45595 (I777752,I2683,I777520,I777840,);
not I_45596 (I777848,I777840);
not I_45597 (I777865,I251701);
not I_45598 (I777882,I251704);
nor I_45599 (I777899,I777882,I251716);
nor I_45600 (I777512,I777848,I777899);
nor I_45601 (I777930,I777882,I251713);
and I_45602 (I777947,I777930,I251695);
or I_45603 (I777964,I777947,I251710);
DFFARX1 I_45604 (I777964,I2683,I777520,I777990,);
nor I_45605 (I777500,I777990,I777546);
not I_45606 (I778012,I777990);
and I_45607 (I778029,I778012,I777546);
nor I_45608 (I777494,I777571,I778029);
nand I_45609 (I778060,I778012,I777622);
nor I_45610 (I777488,I777882,I778060);
nand I_45611 (I777491,I778012,I777800);
nand I_45612 (I778105,I777622,I251704);
nor I_45613 (I777503,I777865,I778105);
not I_45614 (I778166,I2690);
DFFARX1 I_45615 (I1066179,I2683,I778166,I778192,);
DFFARX1 I_45616 (I1066203,I2683,I778166,I778209,);
not I_45617 (I778217,I778209);
not I_45618 (I778234,I1066185);
nor I_45619 (I778251,I778234,I1066194);
not I_45620 (I778268,I1066179);
nor I_45621 (I778285,I778251,I1066200);
nor I_45622 (I778302,I778209,I778285);
DFFARX1 I_45623 (I778302,I2683,I778166,I778152,);
nor I_45624 (I778333,I1066200,I1066194);
nand I_45625 (I778350,I778333,I1066185);
DFFARX1 I_45626 (I778350,I2683,I778166,I778155,);
nor I_45627 (I778381,I778268,I1066200);
nand I_45628 (I778398,I778381,I1066197);
nor I_45629 (I778415,I778192,I778398);
DFFARX1 I_45630 (I778415,I2683,I778166,I778131,);
not I_45631 (I778446,I778398);
nand I_45632 (I778143,I778209,I778446);
DFFARX1 I_45633 (I778398,I2683,I778166,I778486,);
not I_45634 (I778494,I778486);
not I_45635 (I778511,I1066200);
not I_45636 (I778528,I1066191);
nor I_45637 (I778545,I778528,I1066179);
nor I_45638 (I778158,I778494,I778545);
nor I_45639 (I778576,I778528,I1066182);
and I_45640 (I778593,I778576,I1066206);
or I_45641 (I778610,I778593,I1066188);
DFFARX1 I_45642 (I778610,I2683,I778166,I778636,);
nor I_45643 (I778146,I778636,I778192);
not I_45644 (I778658,I778636);
and I_45645 (I778675,I778658,I778192);
nor I_45646 (I778140,I778217,I778675);
nand I_45647 (I778706,I778658,I778268);
nor I_45648 (I778134,I778528,I778706);
nand I_45649 (I778137,I778658,I778446);
nand I_45650 (I778751,I778268,I1066191);
nor I_45651 (I778149,I778511,I778751);
not I_45652 (I778812,I2690);
DFFARX1 I_45653 (I947860,I2683,I778812,I778838,);
DFFARX1 I_45654 (I947842,I2683,I778812,I778855,);
not I_45655 (I778863,I778855);
not I_45656 (I778880,I947851);
nor I_45657 (I778897,I778880,I947863);
not I_45658 (I778914,I947845);
nor I_45659 (I778931,I778897,I947854);
nor I_45660 (I778948,I778855,I778931);
DFFARX1 I_45661 (I778948,I2683,I778812,I778798,);
nor I_45662 (I778979,I947854,I947863);
nand I_45663 (I778996,I778979,I947851);
DFFARX1 I_45664 (I778996,I2683,I778812,I778801,);
nor I_45665 (I779027,I778914,I947854);
nand I_45666 (I779044,I779027,I947866);
nor I_45667 (I779061,I778838,I779044);
DFFARX1 I_45668 (I779061,I2683,I778812,I778777,);
not I_45669 (I779092,I779044);
nand I_45670 (I778789,I778855,I779092);
DFFARX1 I_45671 (I779044,I2683,I778812,I779132,);
not I_45672 (I779140,I779132);
not I_45673 (I779157,I947854);
not I_45674 (I779174,I947842);
nor I_45675 (I779191,I779174,I947845);
nor I_45676 (I778804,I779140,I779191);
nor I_45677 (I779222,I779174,I947848);
and I_45678 (I779239,I779222,I947857);
or I_45679 (I779256,I779239,I947845);
DFFARX1 I_45680 (I779256,I2683,I778812,I779282,);
nor I_45681 (I778792,I779282,I778838);
not I_45682 (I779304,I779282);
and I_45683 (I779321,I779304,I778838);
nor I_45684 (I778786,I778863,I779321);
nand I_45685 (I779352,I779304,I778914);
nor I_45686 (I778780,I779174,I779352);
nand I_45687 (I778783,I779304,I779092);
nand I_45688 (I779397,I778914,I947842);
nor I_45689 (I778795,I779157,I779397);
not I_45690 (I779458,I2690);
DFFARX1 I_45691 (I886592,I2683,I779458,I779484,);
DFFARX1 I_45692 (I886574,I2683,I779458,I779501,);
not I_45693 (I779509,I779501);
not I_45694 (I779526,I886583);
nor I_45695 (I779543,I779526,I886595);
not I_45696 (I779560,I886577);
nor I_45697 (I779577,I779543,I886586);
nor I_45698 (I779594,I779501,I779577);
DFFARX1 I_45699 (I779594,I2683,I779458,I779444,);
nor I_45700 (I779625,I886586,I886595);
nand I_45701 (I779642,I779625,I886583);
DFFARX1 I_45702 (I779642,I2683,I779458,I779447,);
nor I_45703 (I779673,I779560,I886586);
nand I_45704 (I779690,I779673,I886598);
nor I_45705 (I779707,I779484,I779690);
DFFARX1 I_45706 (I779707,I2683,I779458,I779423,);
not I_45707 (I779738,I779690);
nand I_45708 (I779435,I779501,I779738);
DFFARX1 I_45709 (I779690,I2683,I779458,I779778,);
not I_45710 (I779786,I779778);
not I_45711 (I779803,I886586);
not I_45712 (I779820,I886574);
nor I_45713 (I779837,I779820,I886577);
nor I_45714 (I779450,I779786,I779837);
nor I_45715 (I779868,I779820,I886580);
and I_45716 (I779885,I779868,I886589);
or I_45717 (I779902,I779885,I886577);
DFFARX1 I_45718 (I779902,I2683,I779458,I779928,);
nor I_45719 (I779438,I779928,I779484);
not I_45720 (I779950,I779928);
and I_45721 (I779967,I779950,I779484);
nor I_45722 (I779432,I779509,I779967);
nand I_45723 (I779998,I779950,I779560);
nor I_45724 (I779426,I779820,I779998);
nand I_45725 (I779429,I779950,I779738);
nand I_45726 (I780043,I779560,I886574);
nor I_45727 (I779441,I779803,I780043);
not I_45728 (I780104,I2690);
DFFARX1 I_45729 (I350808,I2683,I780104,I780130,);
DFFARX1 I_45730 (I350805,I2683,I780104,I780147,);
not I_45731 (I780155,I780147);
not I_45732 (I780172,I350820);
nor I_45733 (I780189,I780172,I350823);
not I_45734 (I780206,I350811);
nor I_45735 (I780223,I780189,I350817);
nor I_45736 (I780240,I780147,I780223);
DFFARX1 I_45737 (I780240,I2683,I780104,I780090,);
nor I_45738 (I780271,I350817,I350823);
nand I_45739 (I780288,I780271,I350820);
DFFARX1 I_45740 (I780288,I2683,I780104,I780093,);
nor I_45741 (I780319,I780206,I350817);
nand I_45742 (I780336,I780319,I350829);
nor I_45743 (I780353,I780130,I780336);
DFFARX1 I_45744 (I780353,I2683,I780104,I780069,);
not I_45745 (I780384,I780336);
nand I_45746 (I780081,I780147,I780384);
DFFARX1 I_45747 (I780336,I2683,I780104,I780424,);
not I_45748 (I780432,I780424);
not I_45749 (I780449,I350817);
not I_45750 (I780466,I350802);
nor I_45751 (I780483,I780466,I350811);
nor I_45752 (I780096,I780432,I780483);
nor I_45753 (I780514,I780466,I350814);
and I_45754 (I780531,I780514,I350802);
or I_45755 (I780548,I780531,I350826);
DFFARX1 I_45756 (I780548,I2683,I780104,I780574,);
nor I_45757 (I780084,I780574,I780130);
not I_45758 (I780596,I780574);
and I_45759 (I780613,I780596,I780130);
nor I_45760 (I780078,I780155,I780613);
nand I_45761 (I780644,I780596,I780206);
nor I_45762 (I780072,I780466,I780644);
nand I_45763 (I780075,I780596,I780384);
nand I_45764 (I780689,I780206,I350802);
nor I_45765 (I780087,I780449,I780689);
not I_45766 (I780750,I2690);
DFFARX1 I_45767 (I891216,I2683,I780750,I780776,);
DFFARX1 I_45768 (I891198,I2683,I780750,I780793,);
not I_45769 (I780801,I780793);
not I_45770 (I780818,I891207);
nor I_45771 (I780835,I780818,I891219);
not I_45772 (I780852,I891201);
nor I_45773 (I780869,I780835,I891210);
nor I_45774 (I780886,I780793,I780869);
DFFARX1 I_45775 (I780886,I2683,I780750,I780736,);
nor I_45776 (I780917,I891210,I891219);
nand I_45777 (I780934,I780917,I891207);
DFFARX1 I_45778 (I780934,I2683,I780750,I780739,);
nor I_45779 (I780965,I780852,I891210);
nand I_45780 (I780982,I780965,I891222);
nor I_45781 (I780999,I780776,I780982);
DFFARX1 I_45782 (I780999,I2683,I780750,I780715,);
not I_45783 (I781030,I780982);
nand I_45784 (I780727,I780793,I781030);
DFFARX1 I_45785 (I780982,I2683,I780750,I781070,);
not I_45786 (I781078,I781070);
not I_45787 (I781095,I891210);
not I_45788 (I781112,I891198);
nor I_45789 (I781129,I781112,I891201);
nor I_45790 (I780742,I781078,I781129);
nor I_45791 (I781160,I781112,I891204);
and I_45792 (I781177,I781160,I891213);
or I_45793 (I781194,I781177,I891201);
DFFARX1 I_45794 (I781194,I2683,I780750,I781220,);
nor I_45795 (I780730,I781220,I780776);
not I_45796 (I781242,I781220);
and I_45797 (I781259,I781242,I780776);
nor I_45798 (I780724,I780801,I781259);
nand I_45799 (I781290,I781242,I780852);
nor I_45800 (I780718,I781112,I781290);
nand I_45801 (I780721,I781242,I781030);
nand I_45802 (I781335,I780852,I891198);
nor I_45803 (I780733,I781095,I781335);
not I_45804 (I781396,I2690);
DFFARX1 I_45805 (I359512,I2683,I781396,I781422,);
DFFARX1 I_45806 (I359509,I2683,I781396,I781439,);
not I_45807 (I781447,I781439);
not I_45808 (I781464,I359524);
nor I_45809 (I781481,I781464,I359527);
not I_45810 (I781498,I359515);
nor I_45811 (I781515,I781481,I359521);
nor I_45812 (I781532,I781439,I781515);
DFFARX1 I_45813 (I781532,I2683,I781396,I781382,);
nor I_45814 (I781563,I359521,I359527);
nand I_45815 (I781580,I781563,I359524);
DFFARX1 I_45816 (I781580,I2683,I781396,I781385,);
nor I_45817 (I781611,I781498,I359521);
nand I_45818 (I781628,I781611,I359533);
nor I_45819 (I781645,I781422,I781628);
DFFARX1 I_45820 (I781645,I2683,I781396,I781361,);
not I_45821 (I781676,I781628);
nand I_45822 (I781373,I781439,I781676);
DFFARX1 I_45823 (I781628,I2683,I781396,I781716,);
not I_45824 (I781724,I781716);
not I_45825 (I781741,I359521);
not I_45826 (I781758,I359506);
nor I_45827 (I781775,I781758,I359515);
nor I_45828 (I781388,I781724,I781775);
nor I_45829 (I781806,I781758,I359518);
and I_45830 (I781823,I781806,I359506);
or I_45831 (I781840,I781823,I359530);
DFFARX1 I_45832 (I781840,I2683,I781396,I781866,);
nor I_45833 (I781376,I781866,I781422);
not I_45834 (I781888,I781866);
and I_45835 (I781905,I781888,I781422);
nor I_45836 (I781370,I781447,I781905);
nand I_45837 (I781936,I781888,I781498);
nor I_45838 (I781364,I781758,I781936);
nand I_45839 (I781367,I781888,I781676);
nand I_45840 (I781981,I781498,I359506);
nor I_45841 (I781379,I781741,I781981);
not I_45842 (I782042,I2690);
DFFARX1 I_45843 (I853068,I2683,I782042,I782068,);
DFFARX1 I_45844 (I853050,I2683,I782042,I782085,);
not I_45845 (I782093,I782085);
not I_45846 (I782110,I853059);
nor I_45847 (I782127,I782110,I853071);
not I_45848 (I782144,I853053);
nor I_45849 (I782161,I782127,I853062);
nor I_45850 (I782178,I782085,I782161);
DFFARX1 I_45851 (I782178,I2683,I782042,I782028,);
nor I_45852 (I782209,I853062,I853071);
nand I_45853 (I782226,I782209,I853059);
DFFARX1 I_45854 (I782226,I2683,I782042,I782031,);
nor I_45855 (I782257,I782144,I853062);
nand I_45856 (I782274,I782257,I853074);
nor I_45857 (I782291,I782068,I782274);
DFFARX1 I_45858 (I782291,I2683,I782042,I782007,);
not I_45859 (I782322,I782274);
nand I_45860 (I782019,I782085,I782322);
DFFARX1 I_45861 (I782274,I2683,I782042,I782362,);
not I_45862 (I782370,I782362);
not I_45863 (I782387,I853062);
not I_45864 (I782404,I853050);
nor I_45865 (I782421,I782404,I853053);
nor I_45866 (I782034,I782370,I782421);
nor I_45867 (I782452,I782404,I853056);
and I_45868 (I782469,I782452,I853065);
or I_45869 (I782486,I782469,I853053);
DFFARX1 I_45870 (I782486,I2683,I782042,I782512,);
nor I_45871 (I782022,I782512,I782068);
not I_45872 (I782534,I782512);
and I_45873 (I782551,I782534,I782068);
nor I_45874 (I782016,I782093,I782551);
nand I_45875 (I782582,I782534,I782144);
nor I_45876 (I782010,I782404,I782582);
nand I_45877 (I782013,I782534,I782322);
nand I_45878 (I782627,I782144,I853050);
nor I_45879 (I782025,I782387,I782627);
not I_45880 (I782688,I2690);
DFFARX1 I_45881 (I873876,I2683,I782688,I782714,);
DFFARX1 I_45882 (I873858,I2683,I782688,I782731,);
not I_45883 (I782739,I782731);
not I_45884 (I782756,I873867);
nor I_45885 (I782773,I782756,I873879);
not I_45886 (I782790,I873861);
nor I_45887 (I782807,I782773,I873870);
nor I_45888 (I782824,I782731,I782807);
DFFARX1 I_45889 (I782824,I2683,I782688,I782674,);
nor I_45890 (I782855,I873870,I873879);
nand I_45891 (I782872,I782855,I873867);
DFFARX1 I_45892 (I782872,I2683,I782688,I782677,);
nor I_45893 (I782903,I782790,I873870);
nand I_45894 (I782920,I782903,I873882);
nor I_45895 (I782937,I782714,I782920);
DFFARX1 I_45896 (I782937,I2683,I782688,I782653,);
not I_45897 (I782968,I782920);
nand I_45898 (I782665,I782731,I782968);
DFFARX1 I_45899 (I782920,I2683,I782688,I783008,);
not I_45900 (I783016,I783008);
not I_45901 (I783033,I873870);
not I_45902 (I783050,I873858);
nor I_45903 (I783067,I783050,I873861);
nor I_45904 (I782680,I783016,I783067);
nor I_45905 (I783098,I783050,I873864);
and I_45906 (I783115,I783098,I873873);
or I_45907 (I783132,I783115,I873861);
DFFARX1 I_45908 (I783132,I2683,I782688,I783158,);
nor I_45909 (I782668,I783158,I782714);
not I_45910 (I783180,I783158);
and I_45911 (I783197,I783180,I782714);
nor I_45912 (I782662,I782739,I783197);
nand I_45913 (I783228,I783180,I782790);
nor I_45914 (I782656,I783050,I783228);
nand I_45915 (I782659,I783180,I782968);
nand I_45916 (I783273,I782790,I873858);
nor I_45917 (I782671,I783033,I783273);
not I_45918 (I783334,I2690);
DFFARX1 I_45919 (I482113,I2683,I783334,I783360,);
DFFARX1 I_45920 (I482125,I2683,I783334,I783377,);
not I_45921 (I783385,I783377);
not I_45922 (I783402,I482134);
nor I_45923 (I783419,I783402,I482110);
not I_45924 (I783436,I482128);
nor I_45925 (I783453,I783419,I482122);
nor I_45926 (I783470,I783377,I783453);
DFFARX1 I_45927 (I783470,I2683,I783334,I783320,);
nor I_45928 (I783501,I482122,I482110);
nand I_45929 (I783518,I783501,I482134);
DFFARX1 I_45930 (I783518,I2683,I783334,I783323,);
nor I_45931 (I783549,I783436,I482122);
nand I_45932 (I783566,I783549,I482116);
nor I_45933 (I783583,I783360,I783566);
DFFARX1 I_45934 (I783583,I2683,I783334,I783299,);
not I_45935 (I783614,I783566);
nand I_45936 (I783311,I783377,I783614);
DFFARX1 I_45937 (I783566,I2683,I783334,I783654,);
not I_45938 (I783662,I783654);
not I_45939 (I783679,I482122);
not I_45940 (I783696,I482131);
nor I_45941 (I783713,I783696,I482128);
nor I_45942 (I783326,I783662,I783713);
nor I_45943 (I783744,I783696,I482113);
and I_45944 (I783761,I783744,I482110);
or I_45945 (I783778,I783761,I482119);
DFFARX1 I_45946 (I783778,I2683,I783334,I783804,);
nor I_45947 (I783314,I783804,I783360);
not I_45948 (I783826,I783804);
and I_45949 (I783843,I783826,I783360);
nor I_45950 (I783308,I783385,I783843);
nand I_45951 (I783874,I783826,I783436);
nor I_45952 (I783302,I783696,I783874);
nand I_45953 (I783305,I783826,I783614);
nand I_45954 (I783919,I783436,I482131);
nor I_45955 (I783317,I783679,I783919);
not I_45956 (I783980,I2690);
DFFARX1 I_45957 (I294379,I2683,I783980,I784006,);
DFFARX1 I_45958 (I294385,I2683,I783980,I784023,);
not I_45959 (I784031,I784023);
not I_45960 (I784048,I294406);
nor I_45961 (I784065,I784048,I294394);
not I_45962 (I784082,I294403);
nor I_45963 (I784099,I784065,I294388);
nor I_45964 (I784116,I784023,I784099);
DFFARX1 I_45965 (I784116,I2683,I783980,I783966,);
nor I_45966 (I784147,I294388,I294394);
nand I_45967 (I784164,I784147,I294406);
DFFARX1 I_45968 (I784164,I2683,I783980,I783969,);
nor I_45969 (I784195,I784082,I294388);
nand I_45970 (I784212,I784195,I294379);
nor I_45971 (I784229,I784006,I784212);
DFFARX1 I_45972 (I784229,I2683,I783980,I783945,);
not I_45973 (I784260,I784212);
nand I_45974 (I783957,I784023,I784260);
DFFARX1 I_45975 (I784212,I2683,I783980,I784300,);
not I_45976 (I784308,I784300);
not I_45977 (I784325,I294388);
not I_45978 (I784342,I294391);
nor I_45979 (I784359,I784342,I294403);
nor I_45980 (I783972,I784308,I784359);
nor I_45981 (I784390,I784342,I294400);
and I_45982 (I784407,I784390,I294382);
or I_45983 (I784424,I784407,I294397);
DFFARX1 I_45984 (I784424,I2683,I783980,I784450,);
nor I_45985 (I783960,I784450,I784006);
not I_45986 (I784472,I784450);
and I_45987 (I784489,I784472,I784006);
nor I_45988 (I783954,I784031,I784489);
nand I_45989 (I784520,I784472,I784082);
nor I_45990 (I783948,I784342,I784520);
nand I_45991 (I783951,I784472,I784260);
nand I_45992 (I784565,I784082,I294391);
nor I_45993 (I783963,I784325,I784565);
not I_45994 (I784626,I2690);
DFFARX1 I_45995 (I940346,I2683,I784626,I784652,);
DFFARX1 I_45996 (I940328,I2683,I784626,I784669,);
not I_45997 (I784677,I784669);
not I_45998 (I784694,I940337);
nor I_45999 (I784711,I784694,I940349);
not I_46000 (I784728,I940331);
nor I_46001 (I784745,I784711,I940340);
nor I_46002 (I784762,I784669,I784745);
DFFARX1 I_46003 (I784762,I2683,I784626,I784612,);
nor I_46004 (I784793,I940340,I940349);
nand I_46005 (I784810,I784793,I940337);
DFFARX1 I_46006 (I784810,I2683,I784626,I784615,);
nor I_46007 (I784841,I784728,I940340);
nand I_46008 (I784858,I784841,I940352);
nor I_46009 (I784875,I784652,I784858);
DFFARX1 I_46010 (I784875,I2683,I784626,I784591,);
not I_46011 (I784906,I784858);
nand I_46012 (I784603,I784669,I784906);
DFFARX1 I_46013 (I784858,I2683,I784626,I784946,);
not I_46014 (I784954,I784946);
not I_46015 (I784971,I940340);
not I_46016 (I784988,I940328);
nor I_46017 (I785005,I784988,I940331);
nor I_46018 (I784618,I784954,I785005);
nor I_46019 (I785036,I784988,I940334);
and I_46020 (I785053,I785036,I940343);
or I_46021 (I785070,I785053,I940331);
DFFARX1 I_46022 (I785070,I2683,I784626,I785096,);
nor I_46023 (I784606,I785096,I784652);
not I_46024 (I785118,I785096);
and I_46025 (I785135,I785118,I784652);
nor I_46026 (I784600,I784677,I785135);
nand I_46027 (I785166,I785118,I784728);
nor I_46028 (I784594,I784988,I785166);
nand I_46029 (I784597,I785118,I784906);
nand I_46030 (I785211,I784728,I940328);
nor I_46031 (I784609,I784971,I785211);
not I_46032 (I785272,I2690);
DFFARX1 I_46033 (I43765,I2683,I785272,I785298,);
DFFARX1 I_46034 (I43771,I2683,I785272,I785315,);
not I_46035 (I785323,I785315);
not I_46036 (I785340,I43765);
nor I_46037 (I785357,I785340,I43777);
not I_46038 (I785374,I43789);
nor I_46039 (I785391,I785357,I43783);
nor I_46040 (I785408,I785315,I785391);
DFFARX1 I_46041 (I785408,I2683,I785272,I785258,);
nor I_46042 (I785439,I43783,I43777);
nand I_46043 (I785456,I785439,I43765);
DFFARX1 I_46044 (I785456,I2683,I785272,I785261,);
nor I_46045 (I785487,I785374,I43783);
nand I_46046 (I785504,I785487,I43768);
nor I_46047 (I785521,I785298,I785504);
DFFARX1 I_46048 (I785521,I2683,I785272,I785237,);
not I_46049 (I785552,I785504);
nand I_46050 (I785249,I785315,I785552);
DFFARX1 I_46051 (I785504,I2683,I785272,I785592,);
not I_46052 (I785600,I785592);
not I_46053 (I785617,I43783);
not I_46054 (I785634,I43768);
nor I_46055 (I785651,I785634,I43789);
nor I_46056 (I785264,I785600,I785651);
nor I_46057 (I785682,I785634,I43786);
and I_46058 (I785699,I785682,I43780);
or I_46059 (I785716,I785699,I43774);
DFFARX1 I_46060 (I785716,I2683,I785272,I785742,);
nor I_46061 (I785252,I785742,I785298);
not I_46062 (I785764,I785742);
and I_46063 (I785781,I785764,I785298);
nor I_46064 (I785246,I785323,I785781);
nand I_46065 (I785812,I785764,I785374);
nor I_46066 (I785240,I785634,I785812);
nand I_46067 (I785243,I785764,I785552);
nand I_46068 (I785857,I785374,I43768);
nor I_46069 (I785255,I785617,I785857);
not I_46070 (I785918,I2690);
DFFARX1 I_46071 (I111748,I2683,I785918,I785944,);
DFFARX1 I_46072 (I111754,I2683,I785918,I785961,);
not I_46073 (I785969,I785961);
not I_46074 (I785986,I111772);
nor I_46075 (I786003,I785986,I111751);
not I_46076 (I786020,I111757);
nor I_46077 (I786037,I786003,I111763);
nor I_46078 (I786054,I785961,I786037);
DFFARX1 I_46079 (I786054,I2683,I785918,I785904,);
nor I_46080 (I786085,I111763,I111751);
nand I_46081 (I786102,I786085,I111772);
DFFARX1 I_46082 (I786102,I2683,I785918,I785907,);
nor I_46083 (I786133,I786020,I111763);
nand I_46084 (I786150,I786133,I111769);
nor I_46085 (I786167,I785944,I786150);
DFFARX1 I_46086 (I786167,I2683,I785918,I785883,);
not I_46087 (I786198,I786150);
nand I_46088 (I785895,I785961,I786198);
DFFARX1 I_46089 (I786150,I2683,I785918,I786238,);
not I_46090 (I786246,I786238);
not I_46091 (I786263,I111763);
not I_46092 (I786280,I111751);
nor I_46093 (I786297,I786280,I111757);
nor I_46094 (I785910,I786246,I786297);
nor I_46095 (I786328,I786280,I111760);
and I_46096 (I786345,I786328,I111748);
or I_46097 (I786362,I786345,I111766);
DFFARX1 I_46098 (I786362,I2683,I785918,I786388,);
nor I_46099 (I785898,I786388,I785944);
not I_46100 (I786410,I786388);
and I_46101 (I786427,I786410,I785944);
nor I_46102 (I785892,I785969,I786427);
nand I_46103 (I786458,I786410,I786020);
nor I_46104 (I785886,I786280,I786458);
nand I_46105 (I785889,I786410,I786198);
nand I_46106 (I786503,I786020,I111751);
nor I_46107 (I785901,I786263,I786503);
not I_46108 (I786564,I2690);
DFFARX1 I_46109 (I619102,I2683,I786564,I786590,);
DFFARX1 I_46110 (I619099,I2683,I786564,I786607,);
not I_46111 (I786615,I786607);
not I_46112 (I786632,I619099);
nor I_46113 (I786649,I786632,I619102);
not I_46114 (I786666,I619114);
nor I_46115 (I786683,I786649,I619108);
nor I_46116 (I786700,I786607,I786683);
DFFARX1 I_46117 (I786700,I2683,I786564,I786550,);
nor I_46118 (I786731,I619108,I619102);
nand I_46119 (I786748,I786731,I619099);
DFFARX1 I_46120 (I786748,I2683,I786564,I786553,);
nor I_46121 (I786779,I786666,I619108);
nand I_46122 (I786796,I786779,I619096);
nor I_46123 (I786813,I786590,I786796);
DFFARX1 I_46124 (I786813,I2683,I786564,I786529,);
not I_46125 (I786844,I786796);
nand I_46126 (I786541,I786607,I786844);
DFFARX1 I_46127 (I786796,I2683,I786564,I786884,);
not I_46128 (I786892,I786884);
not I_46129 (I786909,I619108);
not I_46130 (I786926,I619105);
nor I_46131 (I786943,I786926,I619114);
nor I_46132 (I786556,I786892,I786943);
nor I_46133 (I786974,I786926,I619111);
and I_46134 (I786991,I786974,I619117);
or I_46135 (I787008,I786991,I619096);
DFFARX1 I_46136 (I787008,I2683,I786564,I787034,);
nor I_46137 (I786544,I787034,I786590);
not I_46138 (I787056,I787034);
and I_46139 (I787073,I787056,I786590);
nor I_46140 (I786538,I786615,I787073);
nand I_46141 (I787104,I787056,I786666);
nor I_46142 (I786532,I786926,I787104);
nand I_46143 (I786535,I787056,I786844);
nand I_46144 (I787149,I786666,I619105);
nor I_46145 (I786547,I786909,I787149);
not I_46146 (I787210,I2690);
DFFARX1 I_46147 (I210456,I2683,I787210,I787236,);
DFFARX1 I_46148 (I210468,I2683,I787210,I787253,);
not I_46149 (I787261,I787253);
not I_46150 (I787278,I210474);
nor I_46151 (I787295,I787278,I210459);
not I_46152 (I787312,I210450);
nor I_46153 (I787329,I787295,I210471);
nor I_46154 (I787346,I787253,I787329);
DFFARX1 I_46155 (I787346,I2683,I787210,I787196,);
nor I_46156 (I787377,I210471,I210459);
nand I_46157 (I787394,I787377,I210474);
DFFARX1 I_46158 (I787394,I2683,I787210,I787199,);
nor I_46159 (I787425,I787312,I210471);
nand I_46160 (I787442,I787425,I210453);
nor I_46161 (I787459,I787236,I787442);
DFFARX1 I_46162 (I787459,I2683,I787210,I787175,);
not I_46163 (I787490,I787442);
nand I_46164 (I787187,I787253,I787490);
DFFARX1 I_46165 (I787442,I2683,I787210,I787530,);
not I_46166 (I787538,I787530);
not I_46167 (I787555,I210471);
not I_46168 (I787572,I210462);
nor I_46169 (I787589,I787572,I210450);
nor I_46170 (I787202,I787538,I787589);
nor I_46171 (I787620,I787572,I210465);
and I_46172 (I787637,I787620,I210453);
or I_46173 (I787654,I787637,I210450);
DFFARX1 I_46174 (I787654,I2683,I787210,I787680,);
nor I_46175 (I787190,I787680,I787236);
not I_46176 (I787702,I787680);
and I_46177 (I787719,I787702,I787236);
nor I_46178 (I787184,I787261,I787719);
nand I_46179 (I787750,I787702,I787312);
nor I_46180 (I787178,I787572,I787750);
nand I_46181 (I787181,I787702,I787490);
nand I_46182 (I787795,I787312,I210462);
nor I_46183 (I787193,I787555,I787795);
not I_46184 (I787856,I2690);
DFFARX1 I_46185 (I170591,I2683,I787856,I787882,);
DFFARX1 I_46186 (I170603,I2683,I787856,I787899,);
not I_46187 (I787907,I787899);
not I_46188 (I787924,I170609);
nor I_46189 (I787941,I787924,I170594);
not I_46190 (I787958,I170585);
nor I_46191 (I787975,I787941,I170606);
nor I_46192 (I787992,I787899,I787975);
DFFARX1 I_46193 (I787992,I2683,I787856,I787842,);
nor I_46194 (I788023,I170606,I170594);
nand I_46195 (I788040,I788023,I170609);
DFFARX1 I_46196 (I788040,I2683,I787856,I787845,);
nor I_46197 (I788071,I787958,I170606);
nand I_46198 (I788088,I788071,I170588);
nor I_46199 (I788105,I787882,I788088);
DFFARX1 I_46200 (I788105,I2683,I787856,I787821,);
not I_46201 (I788136,I788088);
nand I_46202 (I787833,I787899,I788136);
DFFARX1 I_46203 (I788088,I2683,I787856,I788176,);
not I_46204 (I788184,I788176);
not I_46205 (I788201,I170606);
not I_46206 (I788218,I170597);
nor I_46207 (I788235,I788218,I170585);
nor I_46208 (I787848,I788184,I788235);
nor I_46209 (I788266,I788218,I170600);
and I_46210 (I788283,I788266,I170588);
or I_46211 (I788300,I788283,I170585);
DFFARX1 I_46212 (I788300,I2683,I787856,I788326,);
nor I_46213 (I787836,I788326,I787882);
not I_46214 (I788348,I788326);
and I_46215 (I788365,I788348,I787882);
nor I_46216 (I787830,I787907,I788365);
nand I_46217 (I788396,I788348,I787958);
nor I_46218 (I787824,I788218,I788396);
nand I_46219 (I787827,I788348,I788136);
nand I_46220 (I788441,I787958,I170597);
nor I_46221 (I787839,I788201,I788441);
not I_46222 (I788502,I2690);
DFFARX1 I_46223 (I927052,I2683,I788502,I788528,);
DFFARX1 I_46224 (I927034,I2683,I788502,I788545,);
not I_46225 (I788553,I788545);
not I_46226 (I788570,I927043);
nor I_46227 (I788587,I788570,I927055);
not I_46228 (I788604,I927037);
nor I_46229 (I788621,I788587,I927046);
nor I_46230 (I788638,I788545,I788621);
DFFARX1 I_46231 (I788638,I2683,I788502,I788488,);
nor I_46232 (I788669,I927046,I927055);
nand I_46233 (I788686,I788669,I927043);
DFFARX1 I_46234 (I788686,I2683,I788502,I788491,);
nor I_46235 (I788717,I788604,I927046);
nand I_46236 (I788734,I788717,I927058);
nor I_46237 (I788751,I788528,I788734);
DFFARX1 I_46238 (I788751,I2683,I788502,I788467,);
not I_46239 (I788782,I788734);
nand I_46240 (I788479,I788545,I788782);
DFFARX1 I_46241 (I788734,I2683,I788502,I788822,);
not I_46242 (I788830,I788822);
not I_46243 (I788847,I927046);
not I_46244 (I788864,I927034);
nor I_46245 (I788881,I788864,I927037);
nor I_46246 (I788494,I788830,I788881);
nor I_46247 (I788912,I788864,I927040);
and I_46248 (I788929,I788912,I927049);
or I_46249 (I788946,I788929,I927037);
DFFARX1 I_46250 (I788946,I2683,I788502,I788972,);
nor I_46251 (I788482,I788972,I788528);
not I_46252 (I788994,I788972);
and I_46253 (I789011,I788994,I788528);
nor I_46254 (I788476,I788553,I789011);
nand I_46255 (I789042,I788994,I788604);
nor I_46256 (I788470,I788864,I789042);
nand I_46257 (I788473,I788994,I788782);
nand I_46258 (I789087,I788604,I927034);
nor I_46259 (I788485,I788847,I789087);
not I_46260 (I789148,I2690);
DFFARX1 I_46261 (I1018061,I2683,I789148,I789174,);
DFFARX1 I_46262 (I1018055,I2683,I789148,I789191,);
not I_46263 (I789199,I789191);
not I_46264 (I789216,I1018064);
nor I_46265 (I789233,I789216,I1018076);
not I_46266 (I789250,I1018058);
nor I_46267 (I789267,I789233,I1018055);
nor I_46268 (I789284,I789191,I789267);
DFFARX1 I_46269 (I789284,I2683,I789148,I789134,);
nor I_46270 (I789315,I1018055,I1018076);
nand I_46271 (I789332,I789315,I1018064);
DFFARX1 I_46272 (I789332,I2683,I789148,I789137,);
nor I_46273 (I789363,I789250,I1018055);
nand I_46274 (I789380,I789363,I1018052);
nor I_46275 (I789397,I789174,I789380);
DFFARX1 I_46276 (I789397,I2683,I789148,I789113,);
not I_46277 (I789428,I789380);
nand I_46278 (I789125,I789191,I789428);
DFFARX1 I_46279 (I789380,I2683,I789148,I789468,);
not I_46280 (I789476,I789468);
not I_46281 (I789493,I1018055);
not I_46282 (I789510,I1018073);
nor I_46283 (I789527,I789510,I1018058);
nor I_46284 (I789140,I789476,I789527);
nor I_46285 (I789558,I789510,I1018067);
and I_46286 (I789575,I789558,I1018052);
or I_46287 (I789592,I789575,I1018070);
DFFARX1 I_46288 (I789592,I2683,I789148,I789618,);
nor I_46289 (I789128,I789618,I789174);
not I_46290 (I789640,I789618);
and I_46291 (I789657,I789640,I789174);
nor I_46292 (I789122,I789199,I789657);
nand I_46293 (I789688,I789640,I789250);
nor I_46294 (I789116,I789510,I789688);
nand I_46295 (I789119,I789640,I789428);
nand I_46296 (I789733,I789250,I1018073);
nor I_46297 (I789131,I789493,I789733);
not I_46298 (I789794,I2690);
DFFARX1 I_46299 (I562458,I2683,I789794,I789820,);
DFFARX1 I_46300 (I562452,I2683,I789794,I789837,);
not I_46301 (I789845,I789837);
not I_46302 (I789862,I562467);
nor I_46303 (I789879,I789862,I562452);
not I_46304 (I789896,I562461);
nor I_46305 (I789913,I789879,I562470);
nor I_46306 (I789930,I789837,I789913);
DFFARX1 I_46307 (I789930,I2683,I789794,I789780,);
nor I_46308 (I789961,I562470,I562452);
nand I_46309 (I789978,I789961,I562467);
DFFARX1 I_46310 (I789978,I2683,I789794,I789783,);
nor I_46311 (I790009,I789896,I562470);
nand I_46312 (I790026,I790009,I562455);
nor I_46313 (I790043,I789820,I790026);
DFFARX1 I_46314 (I790043,I2683,I789794,I789759,);
not I_46315 (I790074,I790026);
nand I_46316 (I789771,I789837,I790074);
DFFARX1 I_46317 (I790026,I2683,I789794,I790114,);
not I_46318 (I790122,I790114);
not I_46319 (I790139,I562470);
not I_46320 (I790156,I562464);
nor I_46321 (I790173,I790156,I562461);
nor I_46322 (I789786,I790122,I790173);
nor I_46323 (I790204,I790156,I562473);
and I_46324 (I790221,I790204,I562476);
or I_46325 (I790238,I790221,I562455);
DFFARX1 I_46326 (I790238,I2683,I789794,I790264,);
nor I_46327 (I789774,I790264,I789820);
not I_46328 (I790286,I790264);
and I_46329 (I790303,I790286,I789820);
nor I_46330 (I789768,I789845,I790303);
nand I_46331 (I790334,I790286,I789896);
nor I_46332 (I789762,I790156,I790334);
nand I_46333 (I789765,I790286,I790074);
nand I_46334 (I790379,I789896,I562464);
nor I_46335 (I789777,I790139,I790379);
not I_46336 (I790440,I2690);
DFFARX1 I_46337 (I567082,I2683,I790440,I790466,);
DFFARX1 I_46338 (I567076,I2683,I790440,I790483,);
not I_46339 (I790491,I790483);
not I_46340 (I790508,I567091);
nor I_46341 (I790525,I790508,I567076);
not I_46342 (I790542,I567085);
nor I_46343 (I790559,I790525,I567094);
nor I_46344 (I790576,I790483,I790559);
DFFARX1 I_46345 (I790576,I2683,I790440,I790426,);
nor I_46346 (I790607,I567094,I567076);
nand I_46347 (I790624,I790607,I567091);
DFFARX1 I_46348 (I790624,I2683,I790440,I790429,);
nor I_46349 (I790655,I790542,I567094);
nand I_46350 (I790672,I790655,I567079);
nor I_46351 (I790689,I790466,I790672);
DFFARX1 I_46352 (I790689,I2683,I790440,I790405,);
not I_46353 (I790720,I790672);
nand I_46354 (I790417,I790483,I790720);
DFFARX1 I_46355 (I790672,I2683,I790440,I790760,);
not I_46356 (I790768,I790760);
not I_46357 (I790785,I567094);
not I_46358 (I790802,I567088);
nor I_46359 (I790819,I790802,I567085);
nor I_46360 (I790432,I790768,I790819);
nor I_46361 (I790850,I790802,I567097);
and I_46362 (I790867,I790850,I567100);
or I_46363 (I790884,I790867,I567079);
DFFARX1 I_46364 (I790884,I2683,I790440,I790910,);
nor I_46365 (I790420,I790910,I790466);
not I_46366 (I790932,I790910);
and I_46367 (I790949,I790932,I790466);
nor I_46368 (I790414,I790491,I790949);
nand I_46369 (I790980,I790932,I790542);
nor I_46370 (I790408,I790802,I790980);
nand I_46371 (I790411,I790932,I790720);
nand I_46372 (I791025,I790542,I567088);
nor I_46373 (I790423,I790785,I791025);
not I_46374 (I791086,I2690);
DFFARX1 I_46375 (I248530,I2683,I791086,I791112,);
DFFARX1 I_46376 (I248536,I2683,I791086,I791129,);
not I_46377 (I791137,I791129);
not I_46378 (I791154,I248557);
nor I_46379 (I791171,I791154,I248545);
not I_46380 (I791188,I248554);
nor I_46381 (I791205,I791171,I248539);
nor I_46382 (I791222,I791129,I791205);
DFFARX1 I_46383 (I791222,I2683,I791086,I791072,);
nor I_46384 (I791253,I248539,I248545);
nand I_46385 (I791270,I791253,I248557);
DFFARX1 I_46386 (I791270,I2683,I791086,I791075,);
nor I_46387 (I791301,I791188,I248539);
nand I_46388 (I791318,I791301,I248530);
nor I_46389 (I791335,I791112,I791318);
DFFARX1 I_46390 (I791335,I2683,I791086,I791051,);
not I_46391 (I791366,I791318);
nand I_46392 (I791063,I791129,I791366);
DFFARX1 I_46393 (I791318,I2683,I791086,I791406,);
not I_46394 (I791414,I791406);
not I_46395 (I791431,I248539);
not I_46396 (I791448,I248542);
nor I_46397 (I791465,I791448,I248554);
nor I_46398 (I791078,I791414,I791465);
nor I_46399 (I791496,I791448,I248551);
and I_46400 (I791513,I791496,I248533);
or I_46401 (I791530,I791513,I248548);
DFFARX1 I_46402 (I791530,I2683,I791086,I791556,);
nor I_46403 (I791066,I791556,I791112);
not I_46404 (I791578,I791556);
and I_46405 (I791595,I791578,I791112);
nor I_46406 (I791060,I791137,I791595);
nand I_46407 (I791626,I791578,I791188);
nor I_46408 (I791054,I791448,I791626);
nand I_46409 (I791057,I791578,I791366);
nand I_46410 (I791671,I791188,I248542);
nor I_46411 (I791069,I791431,I791671);
not I_46412 (I791732,I2690);
DFFARX1 I_46413 (I915492,I2683,I791732,I791758,);
DFFARX1 I_46414 (I915474,I2683,I791732,I791775,);
not I_46415 (I791783,I791775);
not I_46416 (I791800,I915483);
nor I_46417 (I791817,I791800,I915495);
not I_46418 (I791834,I915477);
nor I_46419 (I791851,I791817,I915486);
nor I_46420 (I791868,I791775,I791851);
DFFARX1 I_46421 (I791868,I2683,I791732,I791718,);
nor I_46422 (I791899,I915486,I915495);
nand I_46423 (I791916,I791899,I915483);
DFFARX1 I_46424 (I791916,I2683,I791732,I791721,);
nor I_46425 (I791947,I791834,I915486);
nand I_46426 (I791964,I791947,I915498);
nor I_46427 (I791981,I791758,I791964);
DFFARX1 I_46428 (I791981,I2683,I791732,I791697,);
not I_46429 (I792012,I791964);
nand I_46430 (I791709,I791775,I792012);
DFFARX1 I_46431 (I791964,I2683,I791732,I792052,);
not I_46432 (I792060,I792052);
not I_46433 (I792077,I915486);
not I_46434 (I792094,I915474);
nor I_46435 (I792111,I792094,I915477);
nor I_46436 (I791724,I792060,I792111);
nor I_46437 (I792142,I792094,I915480);
and I_46438 (I792159,I792142,I915489);
or I_46439 (I792176,I792159,I915477);
DFFARX1 I_46440 (I792176,I2683,I791732,I792202,);
nor I_46441 (I791712,I792202,I791758);
not I_46442 (I792224,I792202);
and I_46443 (I792241,I792224,I791758);
nor I_46444 (I791706,I791783,I792241);
nand I_46445 (I792272,I792224,I791834);
nor I_46446 (I791700,I792094,I792272);
nand I_46447 (I791703,I792224,I792012);
nand I_46448 (I792317,I791834,I915474);
nor I_46449 (I791715,I792077,I792317);
not I_46450 (I792378,I2690);
DFFARX1 I_46451 (I520264,I2683,I792378,I792404,);
DFFARX1 I_46452 (I520258,I2683,I792378,I792421,);
not I_46453 (I792429,I792421);
not I_46454 (I792446,I520273);
nor I_46455 (I792463,I792446,I520258);
not I_46456 (I792480,I520267);
nor I_46457 (I792497,I792463,I520276);
nor I_46458 (I792514,I792421,I792497);
DFFARX1 I_46459 (I792514,I2683,I792378,I792364,);
nor I_46460 (I792545,I520276,I520258);
nand I_46461 (I792562,I792545,I520273);
DFFARX1 I_46462 (I792562,I2683,I792378,I792367,);
nor I_46463 (I792593,I792480,I520276);
nand I_46464 (I792610,I792593,I520261);
nor I_46465 (I792627,I792404,I792610);
DFFARX1 I_46466 (I792627,I2683,I792378,I792343,);
not I_46467 (I792658,I792610);
nand I_46468 (I792355,I792421,I792658);
DFFARX1 I_46469 (I792610,I2683,I792378,I792698,);
not I_46470 (I792706,I792698);
not I_46471 (I792723,I520276);
not I_46472 (I792740,I520270);
nor I_46473 (I792757,I792740,I520267);
nor I_46474 (I792370,I792706,I792757);
nor I_46475 (I792788,I792740,I520279);
and I_46476 (I792805,I792788,I520282);
or I_46477 (I792822,I792805,I520261);
DFFARX1 I_46478 (I792822,I2683,I792378,I792848,);
nor I_46479 (I792358,I792848,I792404);
not I_46480 (I792870,I792848);
and I_46481 (I792887,I792870,I792404);
nor I_46482 (I792352,I792429,I792887);
nand I_46483 (I792918,I792870,I792480);
nor I_46484 (I792346,I792740,I792918);
nand I_46485 (I792349,I792870,I792658);
nand I_46486 (I792963,I792480,I520270);
nor I_46487 (I792361,I792723,I792963);
not I_46488 (I793024,I2690);
DFFARX1 I_46489 (I449167,I2683,I793024,I793050,);
DFFARX1 I_46490 (I449179,I2683,I793024,I793067,);
not I_46491 (I793075,I793067);
not I_46492 (I793092,I449188);
nor I_46493 (I793109,I793092,I449164);
not I_46494 (I793126,I449182);
nor I_46495 (I793143,I793109,I449176);
nor I_46496 (I793160,I793067,I793143);
DFFARX1 I_46497 (I793160,I2683,I793024,I793010,);
nor I_46498 (I793191,I449176,I449164);
nand I_46499 (I793208,I793191,I449188);
DFFARX1 I_46500 (I793208,I2683,I793024,I793013,);
nor I_46501 (I793239,I793126,I449176);
nand I_46502 (I793256,I793239,I449170);
nor I_46503 (I793273,I793050,I793256);
DFFARX1 I_46504 (I793273,I2683,I793024,I792989,);
not I_46505 (I793304,I793256);
nand I_46506 (I793001,I793067,I793304);
DFFARX1 I_46507 (I793256,I2683,I793024,I793344,);
not I_46508 (I793352,I793344);
not I_46509 (I793369,I449176);
not I_46510 (I793386,I449185);
nor I_46511 (I793403,I793386,I449182);
nor I_46512 (I793016,I793352,I793403);
nor I_46513 (I793434,I793386,I449167);
and I_46514 (I793451,I793434,I449164);
or I_46515 (I793468,I793451,I449173);
DFFARX1 I_46516 (I793468,I2683,I793024,I793494,);
nor I_46517 (I793004,I793494,I793050);
not I_46518 (I793516,I793494);
and I_46519 (I793533,I793516,I793050);
nor I_46520 (I792998,I793075,I793533);
nand I_46521 (I793564,I793516,I793126);
nor I_46522 (I792992,I793386,I793564);
nand I_46523 (I792995,I793516,I793304);
nand I_46524 (I793609,I793126,I449185);
nor I_46525 (I793007,I793369,I793609);
not I_46526 (I793670,I2690);
DFFARX1 I_46527 (I639128,I2683,I793670,I793696,);
DFFARX1 I_46528 (I639125,I2683,I793670,I793713,);
not I_46529 (I793721,I793713);
not I_46530 (I793738,I639125);
nor I_46531 (I793755,I793738,I639128);
not I_46532 (I793772,I639140);
nor I_46533 (I793789,I793755,I639134);
nor I_46534 (I793806,I793713,I793789);
DFFARX1 I_46535 (I793806,I2683,I793670,I793656,);
nor I_46536 (I793837,I639134,I639128);
nand I_46537 (I793854,I793837,I639125);
DFFARX1 I_46538 (I793854,I2683,I793670,I793659,);
nor I_46539 (I793885,I793772,I639134);
nand I_46540 (I793902,I793885,I639122);
nor I_46541 (I793919,I793696,I793902);
DFFARX1 I_46542 (I793919,I2683,I793670,I793635,);
not I_46543 (I793950,I793902);
nand I_46544 (I793647,I793713,I793950);
DFFARX1 I_46545 (I793902,I2683,I793670,I793990,);
not I_46546 (I793998,I793990);
not I_46547 (I794015,I639134);
not I_46548 (I794032,I639131);
nor I_46549 (I794049,I794032,I639140);
nor I_46550 (I793662,I793998,I794049);
nor I_46551 (I794080,I794032,I639137);
and I_46552 (I794097,I794080,I639143);
or I_46553 (I794114,I794097,I639122);
DFFARX1 I_46554 (I794114,I2683,I793670,I794140,);
nor I_46555 (I793650,I794140,I793696);
not I_46556 (I794162,I794140);
and I_46557 (I794179,I794162,I793696);
nor I_46558 (I793644,I793721,I794179);
nand I_46559 (I794210,I794162,I793772);
nor I_46560 (I793638,I794032,I794210);
nand I_46561 (I793641,I794162,I793950);
nand I_46562 (I794255,I793772,I639131);
nor I_46563 (I793653,I794015,I794255);
not I_46564 (I794316,I2690);
DFFARX1 I_46565 (I377464,I2683,I794316,I794342,);
DFFARX1 I_46566 (I377461,I2683,I794316,I794359,);
not I_46567 (I794367,I794359);
not I_46568 (I794384,I377476);
nor I_46569 (I794401,I794384,I377479);
not I_46570 (I794418,I377467);
nor I_46571 (I794435,I794401,I377473);
nor I_46572 (I794452,I794359,I794435);
DFFARX1 I_46573 (I794452,I2683,I794316,I794302,);
nor I_46574 (I794483,I377473,I377479);
nand I_46575 (I794500,I794483,I377476);
DFFARX1 I_46576 (I794500,I2683,I794316,I794305,);
nor I_46577 (I794531,I794418,I377473);
nand I_46578 (I794548,I794531,I377485);
nor I_46579 (I794565,I794342,I794548);
DFFARX1 I_46580 (I794565,I2683,I794316,I794281,);
not I_46581 (I794596,I794548);
nand I_46582 (I794293,I794359,I794596);
DFFARX1 I_46583 (I794548,I2683,I794316,I794636,);
not I_46584 (I794644,I794636);
not I_46585 (I794661,I377473);
not I_46586 (I794678,I377458);
nor I_46587 (I794695,I794678,I377467);
nor I_46588 (I794308,I794644,I794695);
nor I_46589 (I794726,I794678,I377470);
and I_46590 (I794743,I794726,I377458);
or I_46591 (I794760,I794743,I377482);
DFFARX1 I_46592 (I794760,I2683,I794316,I794786,);
nor I_46593 (I794296,I794786,I794342);
not I_46594 (I794808,I794786);
and I_46595 (I794825,I794808,I794342);
nor I_46596 (I794290,I794367,I794825);
nand I_46597 (I794856,I794808,I794418);
nor I_46598 (I794284,I794678,I794856);
nand I_46599 (I794287,I794808,I794596);
nand I_46600 (I794901,I794418,I377458);
nor I_46601 (I794299,I794661,I794901);
not I_46602 (I794962,I2690);
DFFARX1 I_46603 (I608698,I2683,I794962,I794988,);
DFFARX1 I_46604 (I608692,I2683,I794962,I795005,);
not I_46605 (I795013,I795005);
not I_46606 (I795030,I608707);
nor I_46607 (I795047,I795030,I608692);
not I_46608 (I795064,I608701);
nor I_46609 (I795081,I795047,I608710);
nor I_46610 (I795098,I795005,I795081);
DFFARX1 I_46611 (I795098,I2683,I794962,I794948,);
nor I_46612 (I795129,I608710,I608692);
nand I_46613 (I795146,I795129,I608707);
DFFARX1 I_46614 (I795146,I2683,I794962,I794951,);
nor I_46615 (I795177,I795064,I608710);
nand I_46616 (I795194,I795177,I608695);
nor I_46617 (I795211,I794988,I795194);
DFFARX1 I_46618 (I795211,I2683,I794962,I794927,);
not I_46619 (I795242,I795194);
nand I_46620 (I794939,I795005,I795242);
DFFARX1 I_46621 (I795194,I2683,I794962,I795282,);
not I_46622 (I795290,I795282);
not I_46623 (I795307,I608710);
not I_46624 (I795324,I608704);
nor I_46625 (I795341,I795324,I608701);
nor I_46626 (I794954,I795290,I795341);
nor I_46627 (I795372,I795324,I608713);
and I_46628 (I795389,I795372,I608716);
or I_46629 (I795406,I795389,I608695);
DFFARX1 I_46630 (I795406,I2683,I794962,I795432,);
nor I_46631 (I794942,I795432,I794988);
not I_46632 (I795454,I795432);
and I_46633 (I795471,I795454,I794988);
nor I_46634 (I794936,I795013,I795471);
nand I_46635 (I795502,I795454,I795064);
nor I_46636 (I794930,I795324,I795502);
nand I_46637 (I794933,I795454,I795242);
nand I_46638 (I795547,I795064,I608704);
nor I_46639 (I794945,I795307,I795547);
not I_46640 (I795608,I2690);
DFFARX1 I_46641 (I1091764,I2683,I795608,I795634,);
DFFARX1 I_46642 (I1091788,I2683,I795608,I795651,);
not I_46643 (I795659,I795651);
not I_46644 (I795676,I1091770);
nor I_46645 (I795693,I795676,I1091779);
not I_46646 (I795710,I1091764);
nor I_46647 (I795727,I795693,I1091785);
nor I_46648 (I795744,I795651,I795727);
DFFARX1 I_46649 (I795744,I2683,I795608,I795594,);
nor I_46650 (I795775,I1091785,I1091779);
nand I_46651 (I795792,I795775,I1091770);
DFFARX1 I_46652 (I795792,I2683,I795608,I795597,);
nor I_46653 (I795823,I795710,I1091785);
nand I_46654 (I795840,I795823,I1091782);
nor I_46655 (I795857,I795634,I795840);
DFFARX1 I_46656 (I795857,I2683,I795608,I795573,);
not I_46657 (I795888,I795840);
nand I_46658 (I795585,I795651,I795888);
DFFARX1 I_46659 (I795840,I2683,I795608,I795928,);
not I_46660 (I795936,I795928);
not I_46661 (I795953,I1091785);
not I_46662 (I795970,I1091776);
nor I_46663 (I795987,I795970,I1091764);
nor I_46664 (I795600,I795936,I795987);
nor I_46665 (I796018,I795970,I1091767);
and I_46666 (I796035,I796018,I1091791);
or I_46667 (I796052,I796035,I1091773);
DFFARX1 I_46668 (I796052,I2683,I795608,I796078,);
nor I_46669 (I795588,I796078,I795634);
not I_46670 (I796100,I796078);
and I_46671 (I796117,I796100,I795634);
nor I_46672 (I795582,I795659,I796117);
nand I_46673 (I796148,I796100,I795710);
nor I_46674 (I795576,I795970,I796148);
nand I_46675 (I795579,I796100,I795888);
nand I_46676 (I796193,I795710,I1091776);
nor I_46677 (I795591,I795953,I796193);
not I_46678 (I796248,I2690);
DFFARX1 I_46679 (I327978,I2683,I796248,I796274,);
DFFARX1 I_46680 (I796274,I2683,I796248,I796291,);
not I_46681 (I796240,I796291);
not I_46682 (I796313,I796274);
DFFARX1 I_46683 (I327966,I2683,I796248,I796339,);
nand I_46684 (I796347,I796339,I327972);
not I_46685 (I796364,I327972);
not I_46686 (I796381,I327969);
nand I_46687 (I796398,I327957,I327954);
and I_46688 (I796415,I327957,I327954);
not I_46689 (I796432,I327981);
nand I_46690 (I796449,I796432,I796381);
nor I_46691 (I796222,I796449,I796347);
nor I_46692 (I796480,I796364,I796449);
nand I_46693 (I796225,I796415,I796480);
not I_46694 (I796511,I327954);
nor I_46695 (I796528,I796511,I327957);
nor I_46696 (I796545,I796528,I327981);
nor I_46697 (I796562,I796313,I796545);
DFFARX1 I_46698 (I796562,I2683,I796248,I796234,);
not I_46699 (I796593,I796528);
DFFARX1 I_46700 (I796593,I2683,I796248,I796237,);
and I_46701 (I796231,I796339,I796528);
nor I_46702 (I796638,I796511,I327963);
and I_46703 (I796655,I796638,I327960);
or I_46704 (I796672,I796655,I327975);
DFFARX1 I_46705 (I796672,I2683,I796248,I796698,);
nor I_46706 (I796706,I796698,I796432);
DFFARX1 I_46707 (I796706,I2683,I796248,I796219,);
nand I_46708 (I796737,I796698,I796339);
nand I_46709 (I796754,I796432,I796737);
nor I_46710 (I796228,I796754,I796398);
not I_46711 (I796809,I2690);
DFFARX1 I_46712 (I1008807,I2683,I796809,I796835,);
DFFARX1 I_46713 (I796835,I2683,I796809,I796852,);
not I_46714 (I796801,I796852);
not I_46715 (I796874,I796835);
DFFARX1 I_46716 (I1008804,I2683,I796809,I796900,);
nand I_46717 (I796908,I796900,I1008810);
not I_46718 (I796925,I1008810);
not I_46719 (I796942,I1008819);
nand I_46720 (I796959,I1008813,I1008807);
and I_46721 (I796976,I1008813,I1008807);
not I_46722 (I796993,I1008825);
nand I_46723 (I797010,I796993,I796942);
nor I_46724 (I796783,I797010,I796908);
nor I_46725 (I797041,I796925,I797010);
nand I_46726 (I796786,I796976,I797041);
not I_46727 (I797072,I1008822);
nor I_46728 (I797089,I797072,I1008813);
nor I_46729 (I797106,I797089,I1008825);
nor I_46730 (I797123,I796874,I797106);
DFFARX1 I_46731 (I797123,I2683,I796809,I796795,);
not I_46732 (I797154,I797089);
DFFARX1 I_46733 (I797154,I2683,I796809,I796798,);
and I_46734 (I796792,I796900,I797089);
nor I_46735 (I797199,I797072,I1008816);
and I_46736 (I797216,I797199,I1008828);
or I_46737 (I797233,I797216,I1008804);
DFFARX1 I_46738 (I797233,I2683,I796809,I797259,);
nor I_46739 (I797267,I797259,I796993);
DFFARX1 I_46740 (I797267,I2683,I796809,I796780,);
nand I_46741 (I797298,I797259,I796900);
nand I_46742 (I797315,I796993,I797298);
nor I_46743 (I796789,I797315,I796959);
not I_46744 (I797370,I2690);
DFFARX1 I_46745 (I839193,I2683,I797370,I797396,);
DFFARX1 I_46746 (I797396,I2683,I797370,I797413,);
not I_46747 (I797362,I797413);
not I_46748 (I797435,I797396);
DFFARX1 I_46749 (I839184,I2683,I797370,I797461,);
nand I_46750 (I797469,I797461,I839181);
not I_46751 (I797486,I839181);
not I_46752 (I797503,I839190);
nand I_46753 (I797520,I839199,I839181);
and I_46754 (I797537,I839199,I839181);
not I_46755 (I797554,I839178);
nand I_46756 (I797571,I797554,I797503);
nor I_46757 (I797344,I797571,I797469);
nor I_46758 (I797602,I797486,I797571);
nand I_46759 (I797347,I797537,I797602);
not I_46760 (I797633,I839187);
nor I_46761 (I797650,I797633,I839199);
nor I_46762 (I797667,I797650,I839178);
nor I_46763 (I797684,I797435,I797667);
DFFARX1 I_46764 (I797684,I2683,I797370,I797356,);
not I_46765 (I797715,I797650);
DFFARX1 I_46766 (I797715,I2683,I797370,I797359,);
and I_46767 (I797353,I797461,I797650);
nor I_46768 (I797760,I797633,I839202);
and I_46769 (I797777,I797760,I839178);
or I_46770 (I797794,I797777,I839196);
DFFARX1 I_46771 (I797794,I2683,I797370,I797820,);
nor I_46772 (I797828,I797820,I797554);
DFFARX1 I_46773 (I797828,I2683,I797370,I797341,);
nand I_46774 (I797859,I797820,I797461);
nand I_46775 (I797876,I797554,I797859);
nor I_46776 (I797350,I797876,I797520);
not I_46777 (I797931,I2690);
DFFARX1 I_46778 (I96477,I2683,I797931,I797957,);
DFFARX1 I_46779 (I797957,I2683,I797931,I797974,);
not I_46780 (I797923,I797974);
not I_46781 (I797996,I797957);
DFFARX1 I_46782 (I96465,I2683,I797931,I798022,);
nand I_46783 (I798030,I798022,I96480);
not I_46784 (I798047,I96480);
not I_46785 (I798064,I96468);
nand I_46786 (I798081,I96489,I96483);
and I_46787 (I798098,I96489,I96483);
not I_46788 (I798115,I96471);
nand I_46789 (I798132,I798115,I798064);
nor I_46790 (I797905,I798132,I798030);
nor I_46791 (I798163,I798047,I798132);
nand I_46792 (I797908,I798098,I798163);
not I_46793 (I798194,I96474);
nor I_46794 (I798211,I798194,I96489);
nor I_46795 (I798228,I798211,I96471);
nor I_46796 (I798245,I797996,I798228);
DFFARX1 I_46797 (I798245,I2683,I797931,I797917,);
not I_46798 (I798276,I798211);
DFFARX1 I_46799 (I798276,I2683,I797931,I797920,);
and I_46800 (I797914,I798022,I798211);
nor I_46801 (I798321,I798194,I96468);
and I_46802 (I798338,I798321,I96465);
or I_46803 (I798355,I798338,I96486);
DFFARX1 I_46804 (I798355,I2683,I797931,I798381,);
nor I_46805 (I798389,I798381,I798115);
DFFARX1 I_46806 (I798389,I2683,I797931,I797902,);
nand I_46807 (I798420,I798381,I798022);
nand I_46808 (I798437,I798115,I798420);
nor I_46809 (I797911,I798437,I798081);
not I_46810 (I798492,I2690);
DFFARX1 I_46811 (I697628,I2683,I798492,I798518,);
DFFARX1 I_46812 (I798518,I2683,I798492,I798535,);
not I_46813 (I798484,I798535);
not I_46814 (I798557,I798518);
DFFARX1 I_46815 (I697625,I2683,I798492,I798583,);
nand I_46816 (I798591,I798583,I697640);
not I_46817 (I798608,I697640);
not I_46818 (I798625,I697637);
nand I_46819 (I798642,I697634,I697622);
and I_46820 (I798659,I697634,I697622);
not I_46821 (I798676,I697619);
nand I_46822 (I798693,I798676,I798625);
nor I_46823 (I798466,I798693,I798591);
nor I_46824 (I798724,I798608,I798693);
nand I_46825 (I798469,I798659,I798724);
not I_46826 (I798755,I697625);
nor I_46827 (I798772,I798755,I697634);
nor I_46828 (I798789,I798772,I697619);
nor I_46829 (I798806,I798557,I798789);
DFFARX1 I_46830 (I798806,I2683,I798492,I798478,);
not I_46831 (I798837,I798772);
DFFARX1 I_46832 (I798837,I2683,I798492,I798481,);
and I_46833 (I798475,I798583,I798772);
nor I_46834 (I798882,I798755,I697631);
and I_46835 (I798899,I798882,I697619);
or I_46836 (I798916,I798899,I697622);
DFFARX1 I_46837 (I798916,I2683,I798492,I798942,);
nor I_46838 (I798950,I798942,I798676);
DFFARX1 I_46839 (I798950,I2683,I798492,I798463,);
nand I_46840 (I798981,I798942,I798583);
nand I_46841 (I798998,I798676,I798981);
nor I_46842 (I798472,I798998,I798642);
not I_46843 (I799053,I2690);
DFFARX1 I_46844 (I94896,I2683,I799053,I799079,);
DFFARX1 I_46845 (I799079,I2683,I799053,I799096,);
not I_46846 (I799045,I799096);
not I_46847 (I799118,I799079);
DFFARX1 I_46848 (I94884,I2683,I799053,I799144,);
nand I_46849 (I799152,I799144,I94899);
not I_46850 (I799169,I94899);
not I_46851 (I799186,I94887);
nand I_46852 (I799203,I94908,I94902);
and I_46853 (I799220,I94908,I94902);
not I_46854 (I799237,I94890);
nand I_46855 (I799254,I799237,I799186);
nor I_46856 (I799027,I799254,I799152);
nor I_46857 (I799285,I799169,I799254);
nand I_46858 (I799030,I799220,I799285);
not I_46859 (I799316,I94893);
nor I_46860 (I799333,I799316,I94908);
nor I_46861 (I799350,I799333,I94890);
nor I_46862 (I799367,I799118,I799350);
DFFARX1 I_46863 (I799367,I2683,I799053,I799039,);
not I_46864 (I799398,I799333);
DFFARX1 I_46865 (I799398,I2683,I799053,I799042,);
and I_46866 (I799036,I799144,I799333);
nor I_46867 (I799443,I799316,I94887);
and I_46868 (I799460,I799443,I94884);
or I_46869 (I799477,I799460,I94905);
DFFARX1 I_46870 (I799477,I2683,I799053,I799503,);
nor I_46871 (I799511,I799503,I799237);
DFFARX1 I_46872 (I799511,I2683,I799053,I799024,);
nand I_46873 (I799542,I799503,I799144);
nand I_46874 (I799559,I799237,I799542);
nor I_46875 (I799033,I799559,I799203);
not I_46876 (I799614,I2690);
DFFARX1 I_46877 (I979876,I2683,I799614,I799640,);
DFFARX1 I_46878 (I799640,I2683,I799614,I799657,);
not I_46879 (I799606,I799657);
not I_46880 (I799679,I799640);
DFFARX1 I_46881 (I979882,I2683,I799614,I799705,);
nand I_46882 (I799713,I799705,I979891);
not I_46883 (I799730,I979891);
not I_46884 (I799747,I979870);
nand I_46885 (I799764,I979873,I979873);
and I_46886 (I799781,I979873,I979873);
not I_46887 (I799798,I979885);
nand I_46888 (I799815,I799798,I799747);
nor I_46889 (I799588,I799815,I799713);
nor I_46890 (I799846,I799730,I799815);
nand I_46891 (I799591,I799781,I799846);
not I_46892 (I799877,I979879);
nor I_46893 (I799894,I799877,I979873);
nor I_46894 (I799911,I799894,I979885);
nor I_46895 (I799928,I799679,I799911);
DFFARX1 I_46896 (I799928,I2683,I799614,I799600,);
not I_46897 (I799959,I799894);
DFFARX1 I_46898 (I799959,I2683,I799614,I799603,);
and I_46899 (I799597,I799705,I799894);
nor I_46900 (I800004,I799877,I979894);
and I_46901 (I800021,I800004,I979870);
or I_46902 (I800038,I800021,I979888);
DFFARX1 I_46903 (I800038,I2683,I799614,I800064,);
nor I_46904 (I800072,I800064,I799798);
DFFARX1 I_46905 (I800072,I2683,I799614,I799585,);
nand I_46906 (I800103,I800064,I799705);
nand I_46907 (I800120,I799798,I800103);
nor I_46908 (I799594,I800120,I799764);
not I_46909 (I800175,I2690);
DFFARX1 I_46910 (I503499,I2683,I800175,I800201,);
DFFARX1 I_46911 (I800201,I2683,I800175,I800218,);
not I_46912 (I800167,I800218);
not I_46913 (I800240,I800201);
DFFARX1 I_46914 (I503511,I2683,I800175,I800266,);
nand I_46915 (I800274,I800266,I503520);
not I_46916 (I800291,I503520);
not I_46917 (I800308,I503502);
nand I_46918 (I800325,I503505,I503496);
and I_46919 (I800342,I503505,I503496);
not I_46920 (I800359,I503514);
nand I_46921 (I800376,I800359,I800308);
nor I_46922 (I800149,I800376,I800274);
nor I_46923 (I800407,I800291,I800376);
nand I_46924 (I800152,I800342,I800407);
not I_46925 (I800438,I503517);
nor I_46926 (I800455,I800438,I503505);
nor I_46927 (I800472,I800455,I503514);
nor I_46928 (I800489,I800240,I800472);
DFFARX1 I_46929 (I800489,I2683,I800175,I800161,);
not I_46930 (I800520,I800455);
DFFARX1 I_46931 (I800520,I2683,I800175,I800164,);
and I_46932 (I800158,I800266,I800455);
nor I_46933 (I800565,I800438,I503496);
and I_46934 (I800582,I800565,I503508);
or I_46935 (I800599,I800582,I503499);
DFFARX1 I_46936 (I800599,I2683,I800175,I800625,);
nor I_46937 (I800633,I800625,I800359);
DFFARX1 I_46938 (I800633,I2683,I800175,I800146,);
nand I_46939 (I800664,I800625,I800266);
nand I_46940 (I800681,I800359,I800664);
nor I_46941 (I800155,I800681,I800325);
not I_46942 (I800736,I2690);
DFFARX1 I_46943 (I786529,I2683,I800736,I800762,);
DFFARX1 I_46944 (I800762,I2683,I800736,I800779,);
not I_46945 (I800728,I800779);
not I_46946 (I800801,I800762);
DFFARX1 I_46947 (I786556,I2683,I800736,I800827,);
nand I_46948 (I800835,I800827,I786547);
not I_46949 (I800852,I786547);
not I_46950 (I800869,I786529);
nand I_46951 (I800886,I786541,I786544);
and I_46952 (I800903,I786541,I786544);
not I_46953 (I800920,I786553);
nand I_46954 (I800937,I800920,I800869);
nor I_46955 (I800710,I800937,I800835);
nor I_46956 (I800968,I800852,I800937);
nand I_46957 (I800713,I800903,I800968);
not I_46958 (I800999,I786538);
nor I_46959 (I801016,I800999,I786541);
nor I_46960 (I801033,I801016,I786553);
nor I_46961 (I801050,I800801,I801033);
DFFARX1 I_46962 (I801050,I2683,I800736,I800722,);
not I_46963 (I801081,I801016);
DFFARX1 I_46964 (I801081,I2683,I800736,I800725,);
and I_46965 (I800719,I800827,I801016);
nor I_46966 (I801126,I800999,I786532);
and I_46967 (I801143,I801126,I786535);
or I_46968 (I801160,I801143,I786550);
DFFARX1 I_46969 (I801160,I2683,I800736,I801186,);
nor I_46970 (I801194,I801186,I800920);
DFFARX1 I_46971 (I801194,I2683,I800736,I800707,);
nand I_46972 (I801225,I801186,I800827);
nand I_46973 (I801242,I800920,I801225);
nor I_46974 (I800716,I801242,I800886);
not I_46975 (I801297,I2690);
DFFARX1 I_46976 (I1028817,I2683,I801297,I801323,);
DFFARX1 I_46977 (I801323,I2683,I801297,I801340,);
not I_46978 (I801289,I801340);
not I_46979 (I801362,I801323);
DFFARX1 I_46980 (I1028802,I2683,I801297,I801388,);
nand I_46981 (I801396,I801388,I1028811);
not I_46982 (I801413,I1028811);
not I_46983 (I801430,I1028805);
nand I_46984 (I801447,I1028823,I1028820);
and I_46985 (I801464,I1028823,I1028820);
not I_46986 (I801481,I1028796);
nand I_46987 (I801498,I801481,I801430);
nor I_46988 (I801271,I801498,I801396);
nor I_46989 (I801529,I801413,I801498);
nand I_46990 (I801274,I801464,I801529);
not I_46991 (I801560,I1028799);
nor I_46992 (I801577,I801560,I1028823);
nor I_46993 (I801594,I801577,I1028796);
nor I_46994 (I801611,I801362,I801594);
DFFARX1 I_46995 (I801611,I2683,I801297,I801283,);
not I_46996 (I801642,I801577);
DFFARX1 I_46997 (I801642,I2683,I801297,I801286,);
and I_46998 (I801280,I801388,I801577);
nor I_46999 (I801687,I801560,I1028796);
and I_47000 (I801704,I801687,I1028814);
or I_47001 (I801721,I801704,I1028808);
DFFARX1 I_47002 (I801721,I2683,I801297,I801747,);
nor I_47003 (I801755,I801747,I801481);
DFFARX1 I_47004 (I801755,I2683,I801297,I801268,);
nand I_47005 (I801786,I801747,I801388);
nand I_47006 (I801803,I801481,I801786);
nor I_47007 (I801277,I801803,I801447);
not I_47008 (I801858,I2690);
DFFARX1 I_47009 (I361706,I2683,I801858,I801884,);
DFFARX1 I_47010 (I801884,I2683,I801858,I801901,);
not I_47011 (I801850,I801901);
not I_47012 (I801923,I801884);
DFFARX1 I_47013 (I361694,I2683,I801858,I801949,);
nand I_47014 (I801957,I801949,I361700);
not I_47015 (I801974,I361700);
not I_47016 (I801991,I361697);
nand I_47017 (I802008,I361685,I361682);
and I_47018 (I802025,I361685,I361682);
not I_47019 (I802042,I361709);
nand I_47020 (I802059,I802042,I801991);
nor I_47021 (I801832,I802059,I801957);
nor I_47022 (I802090,I801974,I802059);
nand I_47023 (I801835,I802025,I802090);
not I_47024 (I802121,I361682);
nor I_47025 (I802138,I802121,I361685);
nor I_47026 (I802155,I802138,I361709);
nor I_47027 (I802172,I801923,I802155);
DFFARX1 I_47028 (I802172,I2683,I801858,I801844,);
not I_47029 (I802203,I802138);
DFFARX1 I_47030 (I802203,I2683,I801858,I801847,);
and I_47031 (I801841,I801949,I802138);
nor I_47032 (I802248,I802121,I361691);
and I_47033 (I802265,I802248,I361688);
or I_47034 (I802282,I802265,I361703);
DFFARX1 I_47035 (I802282,I2683,I801858,I802308,);
nor I_47036 (I802316,I802308,I802042);
DFFARX1 I_47037 (I802316,I2683,I801858,I801829,);
nand I_47038 (I802347,I802308,I801949);
nand I_47039 (I802364,I802042,I802347);
nor I_47040 (I801838,I802364,I802008);
not I_47041 (I802419,I2690);
DFFARX1 I_47042 (I183083,I2683,I802419,I802445,);
DFFARX1 I_47043 (I802445,I2683,I802419,I802462,);
not I_47044 (I802411,I802462);
not I_47045 (I802484,I802445);
DFFARX1 I_47046 (I183098,I2683,I802419,I802510,);
nand I_47047 (I802518,I802510,I183080);
not I_47048 (I802535,I183080);
not I_47049 (I802552,I183089);
nand I_47050 (I802569,I183095,I183086);
and I_47051 (I802586,I183095,I183086);
not I_47052 (I802603,I183083);
nand I_47053 (I802620,I802603,I802552);
nor I_47054 (I802393,I802620,I802518);
nor I_47055 (I802651,I802535,I802620);
nand I_47056 (I802396,I802586,I802651);
not I_47057 (I802682,I183080);
nor I_47058 (I802699,I802682,I183095);
nor I_47059 (I802716,I802699,I183083);
nor I_47060 (I802733,I802484,I802716);
DFFARX1 I_47061 (I802733,I2683,I802419,I802405,);
not I_47062 (I802764,I802699);
DFFARX1 I_47063 (I802764,I2683,I802419,I802408,);
and I_47064 (I802402,I802510,I802699);
nor I_47065 (I802809,I802682,I183104);
and I_47066 (I802826,I802809,I183101);
or I_47067 (I802843,I802826,I183092);
DFFARX1 I_47068 (I802843,I2683,I802419,I802869,);
nor I_47069 (I802877,I802869,I802603);
DFFARX1 I_47070 (I802877,I2683,I802419,I802390,);
nand I_47071 (I802908,I802869,I802510);
nand I_47072 (I802925,I802603,I802908);
nor I_47073 (I802399,I802925,I802569);
not I_47074 (I802980,I2690);
DFFARX1 I_47075 (I203313,I2683,I802980,I803006,);
DFFARX1 I_47076 (I803006,I2683,I802980,I803023,);
not I_47077 (I802972,I803023);
not I_47078 (I803045,I803006);
DFFARX1 I_47079 (I203328,I2683,I802980,I803071,);
nand I_47080 (I803079,I803071,I203310);
not I_47081 (I803096,I203310);
not I_47082 (I803113,I203319);
nand I_47083 (I803130,I203325,I203316);
and I_47084 (I803147,I203325,I203316);
not I_47085 (I803164,I203313);
nand I_47086 (I803181,I803164,I803113);
nor I_47087 (I802954,I803181,I803079);
nor I_47088 (I803212,I803096,I803181);
nand I_47089 (I802957,I803147,I803212);
not I_47090 (I803243,I203310);
nor I_47091 (I803260,I803243,I203325);
nor I_47092 (I803277,I803260,I203313);
nor I_47093 (I803294,I803045,I803277);
DFFARX1 I_47094 (I803294,I2683,I802980,I802966,);
not I_47095 (I803325,I803260);
DFFARX1 I_47096 (I803325,I2683,I802980,I802969,);
and I_47097 (I802963,I803071,I803260);
nor I_47098 (I803370,I803243,I203334);
and I_47099 (I803387,I803370,I203331);
or I_47100 (I803404,I803387,I203322);
DFFARX1 I_47101 (I803404,I2683,I802980,I803430,);
nor I_47102 (I803438,I803430,I803164);
DFFARX1 I_47103 (I803438,I2683,I802980,I802951,);
nand I_47104 (I803469,I803430,I803071);
nand I_47105 (I803486,I803164,I803469);
nor I_47106 (I802960,I803486,I803130);
not I_47107 (I803541,I2690);
DFFARX1 I_47108 (I1058459,I2683,I803541,I803567,);
DFFARX1 I_47109 (I803567,I2683,I803541,I803584,);
not I_47110 (I803533,I803584);
not I_47111 (I803606,I803567);
DFFARX1 I_47112 (I1058453,I2683,I803541,I803632,);
nand I_47113 (I803640,I803632,I1058444);
not I_47114 (I803657,I1058444);
not I_47115 (I803674,I1058471);
nand I_47116 (I803691,I1058456,I1058465);
and I_47117 (I803708,I1058456,I1058465);
not I_47118 (I803725,I1058450);
nand I_47119 (I803742,I803725,I803674);
nor I_47120 (I803515,I803742,I803640);
nor I_47121 (I803773,I803657,I803742);
nand I_47122 (I803518,I803708,I803773);
not I_47123 (I803804,I1058468);
nor I_47124 (I803821,I803804,I1058456);
nor I_47125 (I803838,I803821,I1058450);
nor I_47126 (I803855,I803606,I803838);
DFFARX1 I_47127 (I803855,I2683,I803541,I803527,);
not I_47128 (I803886,I803821);
DFFARX1 I_47129 (I803886,I2683,I803541,I803530,);
and I_47130 (I803524,I803632,I803821);
nor I_47131 (I803931,I803804,I1058462);
and I_47132 (I803948,I803931,I1058444);
or I_47133 (I803965,I803948,I1058447);
DFFARX1 I_47134 (I803965,I2683,I803541,I803991,);
nor I_47135 (I803999,I803991,I803725);
DFFARX1 I_47136 (I803999,I2683,I803541,I803512,);
nand I_47137 (I804030,I803991,I803632);
nand I_47138 (I804047,I803725,I804030);
nor I_47139 (I803521,I804047,I803691);
not I_47140 (I804102,I2690);
DFFARX1 I_47141 (I996669,I2683,I804102,I804128,);
DFFARX1 I_47142 (I804128,I2683,I804102,I804145,);
not I_47143 (I804094,I804145);
not I_47144 (I804167,I804128);
DFFARX1 I_47145 (I996666,I2683,I804102,I804193,);
nand I_47146 (I804201,I804193,I996672);
not I_47147 (I804218,I996672);
not I_47148 (I804235,I996681);
nand I_47149 (I804252,I996675,I996669);
and I_47150 (I804269,I996675,I996669);
not I_47151 (I804286,I996687);
nand I_47152 (I804303,I804286,I804235);
nor I_47153 (I804076,I804303,I804201);
nor I_47154 (I804334,I804218,I804303);
nand I_47155 (I804079,I804269,I804334);
not I_47156 (I804365,I996684);
nor I_47157 (I804382,I804365,I996675);
nor I_47158 (I804399,I804382,I996687);
nor I_47159 (I804416,I804167,I804399);
DFFARX1 I_47160 (I804416,I2683,I804102,I804088,);
not I_47161 (I804447,I804382);
DFFARX1 I_47162 (I804447,I2683,I804102,I804091,);
and I_47163 (I804085,I804193,I804382);
nor I_47164 (I804492,I804365,I996678);
and I_47165 (I804509,I804492,I996690);
or I_47166 (I804526,I804509,I996666);
DFFARX1 I_47167 (I804526,I2683,I804102,I804552,);
nor I_47168 (I804560,I804552,I804286);
DFFARX1 I_47169 (I804560,I2683,I804102,I804073,);
nand I_47170 (I804591,I804552,I804193);
nand I_47171 (I804608,I804286,I804591);
nor I_47172 (I804082,I804608,I804252);
not I_47173 (I804663,I2690);
DFFARX1 I_47174 (I654414,I2683,I804663,I804689,);
DFFARX1 I_47175 (I804689,I2683,I804663,I804706,);
not I_47176 (I804655,I804706);
not I_47177 (I804728,I804689);
DFFARX1 I_47178 (I654411,I2683,I804663,I804754,);
nand I_47179 (I804762,I804754,I654426);
not I_47180 (I804779,I654426);
not I_47181 (I804796,I654423);
nand I_47182 (I804813,I654420,I654408);
and I_47183 (I804830,I654420,I654408);
not I_47184 (I804847,I654405);
nand I_47185 (I804864,I804847,I804796);
nor I_47186 (I804637,I804864,I804762);
nor I_47187 (I804895,I804779,I804864);
nand I_47188 (I804640,I804830,I804895);
not I_47189 (I804926,I654411);
nor I_47190 (I804943,I804926,I654420);
nor I_47191 (I804960,I804943,I654405);
nor I_47192 (I804977,I804728,I804960);
DFFARX1 I_47193 (I804977,I2683,I804663,I804649,);
not I_47194 (I805008,I804943);
DFFARX1 I_47195 (I805008,I2683,I804663,I804652,);
and I_47196 (I804646,I804754,I804943);
nor I_47197 (I805053,I804926,I654417);
and I_47198 (I805070,I805053,I654405);
or I_47199 (I805087,I805070,I654408);
DFFARX1 I_47200 (I805087,I2683,I804663,I805113,);
nor I_47201 (I805121,I805113,I804847);
DFFARX1 I_47202 (I805121,I2683,I804663,I804634,);
nand I_47203 (I805152,I805113,I804754);
nand I_47204 (I805169,I804847,I805152);
nor I_47205 (I804643,I805169,I804813);
not I_47206 (I805224,I2690);
DFFARX1 I_47207 (I360074,I2683,I805224,I805250,);
DFFARX1 I_47208 (I805250,I2683,I805224,I805267,);
not I_47209 (I805216,I805267);
not I_47210 (I805289,I805250);
DFFARX1 I_47211 (I360062,I2683,I805224,I805315,);
nand I_47212 (I805323,I805315,I360068);
not I_47213 (I805340,I360068);
not I_47214 (I805357,I360065);
nand I_47215 (I805374,I360053,I360050);
and I_47216 (I805391,I360053,I360050);
not I_47217 (I805408,I360077);
nand I_47218 (I805425,I805408,I805357);
nor I_47219 (I805198,I805425,I805323);
nor I_47220 (I805456,I805340,I805425);
nand I_47221 (I805201,I805391,I805456);
not I_47222 (I805487,I360050);
nor I_47223 (I805504,I805487,I360053);
nor I_47224 (I805521,I805504,I360077);
nor I_47225 (I805538,I805289,I805521);
DFFARX1 I_47226 (I805538,I2683,I805224,I805210,);
not I_47227 (I805569,I805504);
DFFARX1 I_47228 (I805569,I2683,I805224,I805213,);
and I_47229 (I805207,I805315,I805504);
nor I_47230 (I805614,I805487,I360059);
and I_47231 (I805631,I805614,I360056);
or I_47232 (I805648,I805631,I360071);
DFFARX1 I_47233 (I805648,I2683,I805224,I805674,);
nor I_47234 (I805682,I805674,I805408);
DFFARX1 I_47235 (I805682,I2683,I805224,I805195,);
nand I_47236 (I805713,I805674,I805315);
nand I_47237 (I805730,I805408,I805713);
nor I_47238 (I805204,I805730,I805374);
not I_47239 (I805785,I2690);
DFFARX1 I_47240 (I720637,I2683,I805785,I805811,);
DFFARX1 I_47241 (I805811,I2683,I805785,I805828,);
not I_47242 (I805777,I805828);
not I_47243 (I805850,I805811);
DFFARX1 I_47244 (I720664,I2683,I805785,I805876,);
nand I_47245 (I805884,I805876,I720655);
not I_47246 (I805901,I720655);
not I_47247 (I805918,I720637);
nand I_47248 (I805935,I720649,I720652);
and I_47249 (I805952,I720649,I720652);
not I_47250 (I805969,I720661);
nand I_47251 (I805986,I805969,I805918);
nor I_47252 (I805759,I805986,I805884);
nor I_47253 (I806017,I805901,I805986);
nand I_47254 (I805762,I805952,I806017);
not I_47255 (I806048,I720646);
nor I_47256 (I806065,I806048,I720649);
nor I_47257 (I806082,I806065,I720661);
nor I_47258 (I806099,I805850,I806082);
DFFARX1 I_47259 (I806099,I2683,I805785,I805771,);
not I_47260 (I806130,I806065);
DFFARX1 I_47261 (I806130,I2683,I805785,I805774,);
and I_47262 (I805768,I805876,I806065);
nor I_47263 (I806175,I806048,I720640);
and I_47264 (I806192,I806175,I720643);
or I_47265 (I806209,I806192,I720658);
DFFARX1 I_47266 (I806209,I2683,I805785,I806235,);
nor I_47267 (I806243,I806235,I805969);
DFFARX1 I_47268 (I806243,I2683,I805785,I805756,);
nand I_47269 (I806274,I806235,I805876);
nand I_47270 (I806291,I805969,I806274);
nor I_47271 (I805765,I806291,I805935);
not I_47272 (I806346,I2690);
DFFARX1 I_47273 (I134888,I2683,I806346,I806372,);
DFFARX1 I_47274 (I806372,I2683,I806346,I806389,);
not I_47275 (I806338,I806389);
not I_47276 (I806411,I806372);
DFFARX1 I_47277 (I134903,I2683,I806346,I806437,);
nand I_47278 (I806445,I806437,I134885);
not I_47279 (I806462,I134885);
not I_47280 (I806479,I134894);
nand I_47281 (I806496,I134900,I134891);
and I_47282 (I806513,I134900,I134891);
not I_47283 (I806530,I134888);
nand I_47284 (I806547,I806530,I806479);
nor I_47285 (I806320,I806547,I806445);
nor I_47286 (I806578,I806462,I806547);
nand I_47287 (I806323,I806513,I806578);
not I_47288 (I806609,I134885);
nor I_47289 (I806626,I806609,I134900);
nor I_47290 (I806643,I806626,I134888);
nor I_47291 (I806660,I806411,I806643);
DFFARX1 I_47292 (I806660,I2683,I806346,I806332,);
not I_47293 (I806691,I806626);
DFFARX1 I_47294 (I806691,I2683,I806346,I806335,);
and I_47295 (I806329,I806437,I806626);
nor I_47296 (I806736,I806609,I134909);
and I_47297 (I806753,I806736,I134906);
or I_47298 (I806770,I806753,I134897);
DFFARX1 I_47299 (I806770,I2683,I806346,I806796,);
nor I_47300 (I806804,I806796,I806530);
DFFARX1 I_47301 (I806804,I2683,I806346,I806317,);
nand I_47302 (I806835,I806796,I806437);
nand I_47303 (I806852,I806530,I806835);
nor I_47304 (I806326,I806852,I806496);
not I_47305 (I806907,I2690);
DFFARX1 I_47306 (I728389,I2683,I806907,I806933,);
DFFARX1 I_47307 (I806933,I2683,I806907,I806950,);
not I_47308 (I806899,I806950);
not I_47309 (I806972,I806933);
DFFARX1 I_47310 (I728416,I2683,I806907,I806998,);
nand I_47311 (I807006,I806998,I728407);
not I_47312 (I807023,I728407);
not I_47313 (I807040,I728389);
nand I_47314 (I807057,I728401,I728404);
and I_47315 (I807074,I728401,I728404);
not I_47316 (I807091,I728413);
nand I_47317 (I807108,I807091,I807040);
nor I_47318 (I806881,I807108,I807006);
nor I_47319 (I807139,I807023,I807108);
nand I_47320 (I806884,I807074,I807139);
not I_47321 (I807170,I728398);
nor I_47322 (I807187,I807170,I728401);
nor I_47323 (I807204,I807187,I728413);
nor I_47324 (I807221,I806972,I807204);
DFFARX1 I_47325 (I807221,I2683,I806907,I806893,);
not I_47326 (I807252,I807187);
DFFARX1 I_47327 (I807252,I2683,I806907,I806896,);
and I_47328 (I806890,I806998,I807187);
nor I_47329 (I807297,I807170,I728392);
and I_47330 (I807314,I807297,I728395);
or I_47331 (I807331,I807314,I728410);
DFFARX1 I_47332 (I807331,I2683,I806907,I807357,);
nor I_47333 (I807365,I807357,I807091);
DFFARX1 I_47334 (I807365,I2683,I806907,I806878,);
nand I_47335 (I807396,I807357,I806998);
nand I_47336 (I807413,I807091,I807396);
nor I_47337 (I806887,I807413,I807057);
not I_47338 (I807468,I2690);
DFFARX1 I_47339 (I918379,I2683,I807468,I807494,);
DFFARX1 I_47340 (I807494,I2683,I807468,I807511,);
not I_47341 (I807460,I807511);
not I_47342 (I807533,I807494);
DFFARX1 I_47343 (I918370,I2683,I807468,I807559,);
nand I_47344 (I807567,I807559,I918367);
not I_47345 (I807584,I918367);
not I_47346 (I807601,I918376);
nand I_47347 (I807618,I918385,I918367);
and I_47348 (I807635,I918385,I918367);
not I_47349 (I807652,I918364);
nand I_47350 (I807669,I807652,I807601);
nor I_47351 (I807442,I807669,I807567);
nor I_47352 (I807700,I807584,I807669);
nand I_47353 (I807445,I807635,I807700);
not I_47354 (I807731,I918373);
nor I_47355 (I807748,I807731,I918385);
nor I_47356 (I807765,I807748,I918364);
nor I_47357 (I807782,I807533,I807765);
DFFARX1 I_47358 (I807782,I2683,I807468,I807454,);
not I_47359 (I807813,I807748);
DFFARX1 I_47360 (I807813,I2683,I807468,I807457,);
and I_47361 (I807451,I807559,I807748);
nor I_47362 (I807858,I807731,I918388);
and I_47363 (I807875,I807858,I918364);
or I_47364 (I807892,I807875,I918382);
DFFARX1 I_47365 (I807892,I2683,I807468,I807918,);
nor I_47366 (I807926,I807918,I807652);
DFFARX1 I_47367 (I807926,I2683,I807468,I807439,);
nand I_47368 (I807957,I807918,I807559);
nand I_47369 (I807974,I807652,I807957);
nor I_47370 (I807448,I807974,I807618);
not I_47371 (I808029,I2690);
DFFARX1 I_47372 (I187843,I2683,I808029,I808055,);
DFFARX1 I_47373 (I808055,I2683,I808029,I808072,);
not I_47374 (I808021,I808072);
not I_47375 (I808094,I808055);
DFFARX1 I_47376 (I187858,I2683,I808029,I808120,);
nand I_47377 (I808128,I808120,I187840);
not I_47378 (I808145,I187840);
not I_47379 (I808162,I187849);
nand I_47380 (I808179,I187855,I187846);
and I_47381 (I808196,I187855,I187846);
not I_47382 (I808213,I187843);
nand I_47383 (I808230,I808213,I808162);
nor I_47384 (I808003,I808230,I808128);
nor I_47385 (I808261,I808145,I808230);
nand I_47386 (I808006,I808196,I808261);
not I_47387 (I808292,I187840);
nor I_47388 (I808309,I808292,I187855);
nor I_47389 (I808326,I808309,I187843);
nor I_47390 (I808343,I808094,I808326);
DFFARX1 I_47391 (I808343,I2683,I808029,I808015,);
not I_47392 (I808374,I808309);
DFFARX1 I_47393 (I808374,I2683,I808029,I808018,);
and I_47394 (I808012,I808120,I808309);
nor I_47395 (I808419,I808292,I187864);
and I_47396 (I808436,I808419,I187861);
or I_47397 (I808453,I808436,I187852);
DFFARX1 I_47398 (I808453,I2683,I808029,I808479,);
nor I_47399 (I808487,I808479,I808213);
DFFARX1 I_47400 (I808487,I2683,I808029,I808000,);
nand I_47401 (I808518,I808479,I808120);
nand I_47402 (I808535,I808213,I808518);
nor I_47403 (I808009,I808535,I808179);
not I_47404 (I808590,I2690);
DFFARX1 I_47405 (I1075119,I2683,I808590,I808616,);
DFFARX1 I_47406 (I808616,I2683,I808590,I808633,);
not I_47407 (I808582,I808633);
not I_47408 (I808655,I808616);
DFFARX1 I_47409 (I1075113,I2683,I808590,I808681,);
nand I_47410 (I808689,I808681,I1075104);
not I_47411 (I808706,I1075104);
not I_47412 (I808723,I1075131);
nand I_47413 (I808740,I1075116,I1075125);
and I_47414 (I808757,I1075116,I1075125);
not I_47415 (I808774,I1075110);
nand I_47416 (I808791,I808774,I808723);
nor I_47417 (I808564,I808791,I808689);
nor I_47418 (I808822,I808706,I808791);
nand I_47419 (I808567,I808757,I808822);
not I_47420 (I808853,I1075128);
nor I_47421 (I808870,I808853,I1075116);
nor I_47422 (I808887,I808870,I1075110);
nor I_47423 (I808904,I808655,I808887);
DFFARX1 I_47424 (I808904,I2683,I808590,I808576,);
not I_47425 (I808935,I808870);
DFFARX1 I_47426 (I808935,I2683,I808590,I808579,);
and I_47427 (I808573,I808681,I808870);
nor I_47428 (I808980,I808853,I1075122);
and I_47429 (I808997,I808980,I1075104);
or I_47430 (I809014,I808997,I1075107);
DFFARX1 I_47431 (I809014,I2683,I808590,I809040,);
nor I_47432 (I809048,I809040,I808774);
DFFARX1 I_47433 (I809048,I2683,I808590,I808561,);
nand I_47434 (I809079,I809040,I808681);
nand I_47435 (I809096,I808774,I809079);
nor I_47436 (I808570,I809096,I808740);
not I_47437 (I809151,I2690);
DFFARX1 I_47438 (I921847,I2683,I809151,I809177,);
DFFARX1 I_47439 (I809177,I2683,I809151,I809194,);
not I_47440 (I809143,I809194);
not I_47441 (I809216,I809177);
DFFARX1 I_47442 (I921838,I2683,I809151,I809242,);
nand I_47443 (I809250,I809242,I921835);
not I_47444 (I809267,I921835);
not I_47445 (I809284,I921844);
nand I_47446 (I809301,I921853,I921835);
and I_47447 (I809318,I921853,I921835);
not I_47448 (I809335,I921832);
nand I_47449 (I809352,I809335,I809284);
nor I_47450 (I809125,I809352,I809250);
nor I_47451 (I809383,I809267,I809352);
nand I_47452 (I809128,I809318,I809383);
not I_47453 (I809414,I921841);
nor I_47454 (I809431,I809414,I921853);
nor I_47455 (I809448,I809431,I921832);
nor I_47456 (I809465,I809216,I809448);
DFFARX1 I_47457 (I809465,I2683,I809151,I809137,);
not I_47458 (I809496,I809431);
DFFARX1 I_47459 (I809496,I2683,I809151,I809140,);
and I_47460 (I809134,I809242,I809431);
nor I_47461 (I809541,I809414,I921856);
and I_47462 (I809558,I809541,I921832);
or I_47463 (I809575,I809558,I921850);
DFFARX1 I_47464 (I809575,I2683,I809151,I809601,);
nor I_47465 (I809609,I809601,I809335);
DFFARX1 I_47466 (I809609,I2683,I809151,I809122,);
nand I_47467 (I809640,I809601,I809242);
nand I_47468 (I809657,I809335,I809640);
nor I_47469 (I809131,I809657,I809301);
not I_47470 (I809712,I2690);
DFFARX1 I_47471 (I337226,I2683,I809712,I809738,);
DFFARX1 I_47472 (I809738,I2683,I809712,I809755,);
not I_47473 (I809704,I809755);
not I_47474 (I809777,I809738);
DFFARX1 I_47475 (I337214,I2683,I809712,I809803,);
nand I_47476 (I809811,I809803,I337220);
not I_47477 (I809828,I337220);
not I_47478 (I809845,I337217);
nand I_47479 (I809862,I337205,I337202);
and I_47480 (I809879,I337205,I337202);
not I_47481 (I809896,I337229);
nand I_47482 (I809913,I809896,I809845);
nor I_47483 (I809686,I809913,I809811);
nor I_47484 (I809944,I809828,I809913);
nand I_47485 (I809689,I809879,I809944);
not I_47486 (I809975,I337202);
nor I_47487 (I809992,I809975,I337205);
nor I_47488 (I810009,I809992,I337229);
nor I_47489 (I810026,I809777,I810009);
DFFARX1 I_47490 (I810026,I2683,I809712,I809698,);
not I_47491 (I810057,I809992);
DFFARX1 I_47492 (I810057,I2683,I809712,I809701,);
and I_47493 (I809695,I809803,I809992);
nor I_47494 (I810102,I809975,I337211);
and I_47495 (I810119,I810102,I337208);
or I_47496 (I810136,I810119,I337223);
DFFARX1 I_47497 (I810136,I2683,I809712,I810162,);
nor I_47498 (I810170,I810162,I809896);
DFFARX1 I_47499 (I810170,I2683,I809712,I809683,);
nand I_47500 (I810201,I810162,I809803);
nand I_47501 (I810218,I809896,I810201);
nor I_47502 (I809692,I810218,I809862);
not I_47503 (I810273,I2690);
DFFARX1 I_47504 (I1468,I2683,I810273,I810299,);
DFFARX1 I_47505 (I810299,I2683,I810273,I810316,);
not I_47506 (I810265,I810316);
not I_47507 (I810338,I810299);
DFFARX1 I_47508 (I1596,I2683,I810273,I810364,);
nand I_47509 (I810372,I810364,I1828);
not I_47510 (I810389,I1828);
not I_47511 (I810406,I2580);
nand I_47512 (I810423,I1628,I2436);
and I_47513 (I810440,I1628,I2436);
not I_47514 (I810457,I1476);
nand I_47515 (I810474,I810457,I810406);
nor I_47516 (I810247,I810474,I810372);
nor I_47517 (I810505,I810389,I810474);
nand I_47518 (I810250,I810440,I810505);
not I_47519 (I810536,I1484);
nor I_47520 (I810553,I810536,I1628);
nor I_47521 (I810570,I810553,I1476);
nor I_47522 (I810587,I810338,I810570);
DFFARX1 I_47523 (I810587,I2683,I810273,I810259,);
not I_47524 (I810618,I810553);
DFFARX1 I_47525 (I810618,I2683,I810273,I810262,);
and I_47526 (I810256,I810364,I810553);
nor I_47527 (I810663,I810536,I1388);
and I_47528 (I810680,I810663,I1380);
or I_47529 (I810697,I810680,I1764);
DFFARX1 I_47530 (I810697,I2683,I810273,I810723,);
nor I_47531 (I810731,I810723,I810457);
DFFARX1 I_47532 (I810731,I2683,I810273,I810244,);
nand I_47533 (I810762,I810723,I810364);
nand I_47534 (I810779,I810457,I810762);
nor I_47535 (I810253,I810779,I810423);
not I_47536 (I810834,I2690);
DFFARX1 I_47537 (I324714,I2683,I810834,I810860,);
DFFARX1 I_47538 (I810860,I2683,I810834,I810877,);
not I_47539 (I810826,I810877);
not I_47540 (I810899,I810860);
DFFARX1 I_47541 (I324702,I2683,I810834,I810925,);
nand I_47542 (I810933,I810925,I324708);
not I_47543 (I810950,I324708);
not I_47544 (I810967,I324705);
nand I_47545 (I810984,I324693,I324690);
and I_47546 (I811001,I324693,I324690);
not I_47547 (I811018,I324717);
nand I_47548 (I811035,I811018,I810967);
nor I_47549 (I810808,I811035,I810933);
nor I_47550 (I811066,I810950,I811035);
nand I_47551 (I810811,I811001,I811066);
not I_47552 (I811097,I324690);
nor I_47553 (I811114,I811097,I324693);
nor I_47554 (I811131,I811114,I324717);
nor I_47555 (I811148,I810899,I811131);
DFFARX1 I_47556 (I811148,I2683,I810834,I810820,);
not I_47557 (I811179,I811114);
DFFARX1 I_47558 (I811179,I2683,I810834,I810823,);
and I_47559 (I810817,I810925,I811114);
nor I_47560 (I811224,I811097,I324699);
and I_47561 (I811241,I811224,I324696);
or I_47562 (I811258,I811241,I324711);
DFFARX1 I_47563 (I811258,I2683,I810834,I811284,);
nor I_47564 (I811292,I811284,I811018);
DFFARX1 I_47565 (I811292,I2683,I810834,I810805,);
nand I_47566 (I811323,I811284,I810925);
nand I_47567 (I811340,I811018,I811323);
nor I_47568 (I810814,I811340,I810984);
not I_47569 (I811395,I2690);
DFFARX1 I_47570 (I442806,I2683,I811395,I811421,);
DFFARX1 I_47571 (I811421,I2683,I811395,I811438,);
not I_47572 (I811387,I811438);
not I_47573 (I811460,I811421);
DFFARX1 I_47574 (I442821,I2683,I811395,I811486,);
nand I_47575 (I811494,I811486,I442812);
not I_47576 (I811511,I442812);
not I_47577 (I811528,I442818);
nand I_47578 (I811545,I442815,I442824);
and I_47579 (I811562,I442815,I442824);
not I_47580 (I811579,I442809);
nand I_47581 (I811596,I811579,I811528);
nor I_47582 (I811369,I811596,I811494);
nor I_47583 (I811627,I811511,I811596);
nand I_47584 (I811372,I811562,I811627);
not I_47585 (I811658,I442806);
nor I_47586 (I811675,I811658,I442815);
nor I_47587 (I811692,I811675,I442809);
nor I_47588 (I811709,I811460,I811692);
DFFARX1 I_47589 (I811709,I2683,I811395,I811381,);
not I_47590 (I811740,I811675);
DFFARX1 I_47591 (I811740,I2683,I811395,I811384,);
and I_47592 (I811378,I811486,I811675);
nor I_47593 (I811785,I811658,I442830);
and I_47594 (I811802,I811785,I442809);
or I_47595 (I811819,I811802,I442827);
DFFARX1 I_47596 (I811819,I2683,I811395,I811845,);
nor I_47597 (I811853,I811845,I811579);
DFFARX1 I_47598 (I811853,I2683,I811395,I811366,);
nand I_47599 (I811884,I811845,I811486);
nand I_47600 (I811901,I811579,I811884);
nor I_47601 (I811375,I811901,I811545);
not I_47602 (I811956,I2690);
DFFARX1 I_47603 (I527775,I2683,I811956,I811982,);
DFFARX1 I_47604 (I811982,I2683,I811956,I811999,);
not I_47605 (I811948,I811999);
not I_47606 (I812021,I811982);
DFFARX1 I_47607 (I527787,I2683,I811956,I812047,);
nand I_47608 (I812055,I812047,I527796);
not I_47609 (I812072,I527796);
not I_47610 (I812089,I527778);
nand I_47611 (I812106,I527781,I527772);
and I_47612 (I812123,I527781,I527772);
not I_47613 (I812140,I527790);
nand I_47614 (I812157,I812140,I812089);
nor I_47615 (I811930,I812157,I812055);
nor I_47616 (I812188,I812072,I812157);
nand I_47617 (I811933,I812123,I812188);
not I_47618 (I812219,I527793);
nor I_47619 (I812236,I812219,I527781);
nor I_47620 (I812253,I812236,I527790);
nor I_47621 (I812270,I812021,I812253);
DFFARX1 I_47622 (I812270,I2683,I811956,I811942,);
not I_47623 (I812301,I812236);
DFFARX1 I_47624 (I812301,I2683,I811956,I811945,);
and I_47625 (I811939,I812047,I812236);
nor I_47626 (I812346,I812219,I527772);
and I_47627 (I812363,I812346,I527784);
or I_47628 (I812380,I812363,I527775);
DFFARX1 I_47629 (I812380,I2683,I811956,I812406,);
nor I_47630 (I812414,I812406,I812140);
DFFARX1 I_47631 (I812414,I2683,I811956,I811927,);
nand I_47632 (I812445,I812406,I812047);
nand I_47633 (I812462,I812140,I812445);
nor I_47634 (I811936,I812462,I812106);
not I_47635 (I812517,I2690);
DFFARX1 I_47636 (I963012,I2683,I812517,I812543,);
DFFARX1 I_47637 (I812543,I2683,I812517,I812560,);
not I_47638 (I812509,I812560);
not I_47639 (I812582,I812543);
DFFARX1 I_47640 (I963018,I2683,I812517,I812608,);
nand I_47641 (I812616,I812608,I963027);
not I_47642 (I812633,I963027);
not I_47643 (I812650,I963006);
nand I_47644 (I812667,I963009,I963009);
and I_47645 (I812684,I963009,I963009);
not I_47646 (I812701,I963021);
nand I_47647 (I812718,I812701,I812650);
nor I_47648 (I812491,I812718,I812616);
nor I_47649 (I812749,I812633,I812718);
nand I_47650 (I812494,I812684,I812749);
not I_47651 (I812780,I963015);
nor I_47652 (I812797,I812780,I963009);
nor I_47653 (I812814,I812797,I963021);
nor I_47654 (I812831,I812582,I812814);
DFFARX1 I_47655 (I812831,I2683,I812517,I812503,);
not I_47656 (I812862,I812797);
DFFARX1 I_47657 (I812862,I2683,I812517,I812506,);
and I_47658 (I812500,I812608,I812797);
nor I_47659 (I812907,I812780,I963030);
and I_47660 (I812924,I812907,I963006);
or I_47661 (I812941,I812924,I963024);
DFFARX1 I_47662 (I812941,I2683,I812517,I812967,);
nor I_47663 (I812975,I812967,I812701);
DFFARX1 I_47664 (I812975,I2683,I812517,I812488,);
nand I_47665 (I813006,I812967,I812608);
nand I_47666 (I813023,I812701,I813006);
nor I_47667 (I812497,I813023,I812667);
not I_47668 (I813078,I2690);
DFFARX1 I_47669 (I631226,I2683,I813078,I813104,);
DFFARX1 I_47670 (I813104,I2683,I813078,I813121,);
not I_47671 (I813070,I813121);
not I_47672 (I813143,I813104);
DFFARX1 I_47673 (I631223,I2683,I813078,I813169,);
nand I_47674 (I813177,I813169,I631238);
not I_47675 (I813194,I631238);
not I_47676 (I813211,I631235);
nand I_47677 (I813228,I631232,I631220);
and I_47678 (I813245,I631232,I631220);
not I_47679 (I813262,I631217);
nand I_47680 (I813279,I813262,I813211);
nor I_47681 (I813052,I813279,I813177);
nor I_47682 (I813310,I813194,I813279);
nand I_47683 (I813055,I813245,I813310);
not I_47684 (I813341,I631223);
nor I_47685 (I813358,I813341,I631232);
nor I_47686 (I813375,I813358,I631217);
nor I_47687 (I813392,I813143,I813375);
DFFARX1 I_47688 (I813392,I2683,I813078,I813064,);
not I_47689 (I813423,I813358);
DFFARX1 I_47690 (I813423,I2683,I813078,I813067,);
and I_47691 (I813061,I813169,I813358);
nor I_47692 (I813468,I813341,I631229);
and I_47693 (I813485,I813468,I631217);
or I_47694 (I813502,I813485,I631220);
DFFARX1 I_47695 (I813502,I2683,I813078,I813528,);
nor I_47696 (I813536,I813528,I813262);
DFFARX1 I_47697 (I813536,I2683,I813078,I813049,);
nand I_47698 (I813567,I813528,I813169);
nand I_47699 (I813584,I813262,I813567);
nor I_47700 (I813058,I813584,I813228);
not I_47701 (I813639,I2690);
DFFARX1 I_47702 (I1065004,I2683,I813639,I813665,);
DFFARX1 I_47703 (I813665,I2683,I813639,I813682,);
not I_47704 (I813631,I813682);
not I_47705 (I813704,I813665);
DFFARX1 I_47706 (I1064998,I2683,I813639,I813730,);
nand I_47707 (I813738,I813730,I1064989);
not I_47708 (I813755,I1064989);
not I_47709 (I813772,I1065016);
nand I_47710 (I813789,I1065001,I1065010);
and I_47711 (I813806,I1065001,I1065010);
not I_47712 (I813823,I1064995);
nand I_47713 (I813840,I813823,I813772);
nor I_47714 (I813613,I813840,I813738);
nor I_47715 (I813871,I813755,I813840);
nand I_47716 (I813616,I813806,I813871);
not I_47717 (I813902,I1065013);
nor I_47718 (I813919,I813902,I1065001);
nor I_47719 (I813936,I813919,I1064995);
nor I_47720 (I813953,I813704,I813936);
DFFARX1 I_47721 (I813953,I2683,I813639,I813625,);
not I_47722 (I813984,I813919);
DFFARX1 I_47723 (I813984,I2683,I813639,I813628,);
and I_47724 (I813622,I813730,I813919);
nor I_47725 (I814029,I813902,I1065007);
and I_47726 (I814046,I814029,I1064989);
or I_47727 (I814063,I814046,I1064992);
DFFARX1 I_47728 (I814063,I2683,I813639,I814089,);
nor I_47729 (I814097,I814089,I813823);
DFFARX1 I_47730 (I814097,I2683,I813639,I813610,);
nand I_47731 (I814128,I814089,I813730);
nand I_47732 (I814145,I813823,I814128);
nor I_47733 (I813619,I814145,I813789);
not I_47734 (I814200,I2690);
DFFARX1 I_47735 (I186058,I2683,I814200,I814226,);
DFFARX1 I_47736 (I814226,I2683,I814200,I814243,);
not I_47737 (I814192,I814243);
not I_47738 (I814265,I814226);
DFFARX1 I_47739 (I186073,I2683,I814200,I814291,);
nand I_47740 (I814299,I814291,I186055);
not I_47741 (I814316,I186055);
not I_47742 (I814333,I186064);
nand I_47743 (I814350,I186070,I186061);
and I_47744 (I814367,I186070,I186061);
not I_47745 (I814384,I186058);
nand I_47746 (I814401,I814384,I814333);
nor I_47747 (I814174,I814401,I814299);
nor I_47748 (I814432,I814316,I814401);
nand I_47749 (I814177,I814367,I814432);
not I_47750 (I814463,I186055);
nor I_47751 (I814480,I814463,I186070);
nor I_47752 (I814497,I814480,I186058);
nor I_47753 (I814514,I814265,I814497);
DFFARX1 I_47754 (I814514,I2683,I814200,I814186,);
not I_47755 (I814545,I814480);
DFFARX1 I_47756 (I814545,I2683,I814200,I814189,);
and I_47757 (I814183,I814291,I814480);
nor I_47758 (I814590,I814463,I186079);
and I_47759 (I814607,I814590,I186076);
or I_47760 (I814624,I814607,I186067);
DFFARX1 I_47761 (I814624,I2683,I814200,I814650,);
nor I_47762 (I814658,I814650,I814384);
DFFARX1 I_47763 (I814658,I2683,I814200,I814171,);
nand I_47764 (I814689,I814650,I814291);
nand I_47765 (I814706,I814384,I814689);
nor I_47766 (I814180,I814706,I814350);
not I_47767 (I814761,I2690);
DFFARX1 I_47768 (I490780,I2683,I814761,I814787,);
DFFARX1 I_47769 (I814787,I2683,I814761,I814804,);
not I_47770 (I814753,I814804);
not I_47771 (I814826,I814787);
DFFARX1 I_47772 (I490795,I2683,I814761,I814852,);
nand I_47773 (I814860,I814852,I490786);
not I_47774 (I814877,I490786);
not I_47775 (I814894,I490792);
nand I_47776 (I814911,I490789,I490798);
and I_47777 (I814928,I490789,I490798);
not I_47778 (I814945,I490783);
nand I_47779 (I814962,I814945,I814894);
nor I_47780 (I814735,I814962,I814860);
nor I_47781 (I814993,I814877,I814962);
nand I_47782 (I814738,I814928,I814993);
not I_47783 (I815024,I490780);
nor I_47784 (I815041,I815024,I490789);
nor I_47785 (I815058,I815041,I490783);
nor I_47786 (I815075,I814826,I815058);
DFFARX1 I_47787 (I815075,I2683,I814761,I814747,);
not I_47788 (I815106,I815041);
DFFARX1 I_47789 (I815106,I2683,I814761,I814750,);
and I_47790 (I814744,I814852,I815041);
nor I_47791 (I815151,I815024,I490804);
and I_47792 (I815168,I815151,I490783);
or I_47793 (I815185,I815168,I490801);
DFFARX1 I_47794 (I815185,I2683,I814761,I815211,);
nor I_47795 (I815219,I815211,I814945);
DFFARX1 I_47796 (I815219,I2683,I814761,I814732,);
nand I_47797 (I815250,I815211,I814852);
nand I_47798 (I815267,I814945,I815250);
nor I_47799 (I814741,I815267,I814911);
not I_47800 (I815322,I2690);
DFFARX1 I_47801 (I27446,I2683,I815322,I815348,);
DFFARX1 I_47802 (I815348,I2683,I815322,I815365,);
not I_47803 (I815314,I815365);
not I_47804 (I815387,I815348);
DFFARX1 I_47805 (I27431,I2683,I815322,I815413,);
nand I_47806 (I815421,I815413,I27443);
not I_47807 (I815438,I27443);
not I_47808 (I815455,I27449);
nand I_47809 (I815472,I27437,I27428);
and I_47810 (I815489,I27437,I27428);
not I_47811 (I815506,I27434);
nand I_47812 (I815523,I815506,I815455);
nor I_47813 (I815296,I815523,I815421);
nor I_47814 (I815554,I815438,I815523);
nand I_47815 (I815299,I815489,I815554);
not I_47816 (I815585,I27440);
nor I_47817 (I815602,I815585,I27437);
nor I_47818 (I815619,I815602,I27434);
nor I_47819 (I815636,I815387,I815619);
DFFARX1 I_47820 (I815636,I2683,I815322,I815308,);
not I_47821 (I815667,I815602);
DFFARX1 I_47822 (I815667,I2683,I815322,I815311,);
and I_47823 (I815305,I815413,I815602);
nor I_47824 (I815712,I815585,I27428);
and I_47825 (I815729,I815712,I27452);
or I_47826 (I815746,I815729,I27431);
DFFARX1 I_47827 (I815746,I2683,I815322,I815772,);
nor I_47828 (I815780,I815772,I815506);
DFFARX1 I_47829 (I815780,I2683,I815322,I815293,);
nand I_47830 (I815811,I815772,I815413);
nand I_47831 (I815828,I815506,I815811);
nor I_47832 (I815302,I815828,I815472);
not I_47833 (I815883,I2690);
DFFARX1 I_47834 (I1046559,I2683,I815883,I815909,);
DFFARX1 I_47835 (I815909,I2683,I815883,I815926,);
not I_47836 (I815875,I815926);
not I_47837 (I815948,I815909);
DFFARX1 I_47838 (I1046553,I2683,I815883,I815974,);
nand I_47839 (I815982,I815974,I1046544);
not I_47840 (I815999,I1046544);
not I_47841 (I816016,I1046571);
nand I_47842 (I816033,I1046556,I1046565);
and I_47843 (I816050,I1046556,I1046565);
not I_47844 (I816067,I1046550);
nand I_47845 (I816084,I816067,I816016);
nor I_47846 (I815857,I816084,I815982);
nor I_47847 (I816115,I815999,I816084);
nand I_47848 (I815860,I816050,I816115);
not I_47849 (I816146,I1046568);
nor I_47850 (I816163,I816146,I1046556);
nor I_47851 (I816180,I816163,I1046550);
nor I_47852 (I816197,I815948,I816180);
DFFARX1 I_47853 (I816197,I2683,I815883,I815869,);
not I_47854 (I816228,I816163);
DFFARX1 I_47855 (I816228,I2683,I815883,I815872,);
and I_47856 (I815866,I815974,I816163);
nor I_47857 (I816273,I816146,I1046562);
and I_47858 (I816290,I816273,I1046544);
or I_47859 (I816307,I816290,I1046547);
DFFARX1 I_47860 (I816307,I2683,I815883,I816333,);
nor I_47861 (I816341,I816333,I816067);
DFFARX1 I_47862 (I816341,I2683,I815883,I815854,);
nand I_47863 (I816372,I816333,I815974);
nand I_47864 (I816389,I816067,I816372);
nor I_47865 (I815863,I816389,I816033);
not I_47866 (I816444,I2690);
DFFARX1 I_47867 (I578061,I2683,I816444,I816470,);
DFFARX1 I_47868 (I816470,I2683,I816444,I816487,);
not I_47869 (I816436,I816487);
not I_47870 (I816509,I816470);
DFFARX1 I_47871 (I578073,I2683,I816444,I816535,);
nand I_47872 (I816543,I816535,I578082);
not I_47873 (I816560,I578082);
not I_47874 (I816577,I578064);
nand I_47875 (I816594,I578067,I578058);
and I_47876 (I816611,I578067,I578058);
not I_47877 (I816628,I578076);
nand I_47878 (I816645,I816628,I816577);
nor I_47879 (I816418,I816645,I816543);
nor I_47880 (I816676,I816560,I816645);
nand I_47881 (I816421,I816611,I816676);
not I_47882 (I816707,I578079);
nor I_47883 (I816724,I816707,I578067);
nor I_47884 (I816741,I816724,I578076);
nor I_47885 (I816758,I816509,I816741);
DFFARX1 I_47886 (I816758,I2683,I816444,I816430,);
not I_47887 (I816789,I816724);
DFFARX1 I_47888 (I816789,I2683,I816444,I816433,);
and I_47889 (I816427,I816535,I816724);
nor I_47890 (I816834,I816707,I578058);
and I_47891 (I816851,I816834,I578070);
or I_47892 (I816868,I816851,I578061);
DFFARX1 I_47893 (I816868,I2683,I816444,I816894,);
nor I_47894 (I816902,I816894,I816628);
DFFARX1 I_47895 (I816902,I2683,I816444,I816415,);
nand I_47896 (I816933,I816894,I816535);
nand I_47897 (I816950,I816628,I816933);
nor I_47898 (I816424,I816950,I816594);
not I_47899 (I817005,I2690);
DFFARX1 I_47900 (I10434,I2683,I817005,I817031,);
DFFARX1 I_47901 (I817031,I2683,I817005,I817048,);
not I_47902 (I816997,I817048);
not I_47903 (I817070,I817031);
DFFARX1 I_47904 (I10446,I2683,I817005,I817096,);
nand I_47905 (I817104,I817096,I10443);
not I_47906 (I817121,I10443);
not I_47907 (I817138,I10434);
nand I_47908 (I817155,I10428,I10428);
and I_47909 (I817172,I10428,I10428);
not I_47910 (I817189,I10449);
nand I_47911 (I817206,I817189,I817138);
nor I_47912 (I816979,I817206,I817104);
nor I_47913 (I817237,I817121,I817206);
nand I_47914 (I816982,I817172,I817237);
not I_47915 (I817268,I10440);
nor I_47916 (I817285,I817268,I10428);
nor I_47917 (I817302,I817285,I10449);
nor I_47918 (I817319,I817070,I817302);
DFFARX1 I_47919 (I817319,I2683,I817005,I816991,);
not I_47920 (I817350,I817285);
DFFARX1 I_47921 (I817350,I2683,I817005,I816994,);
and I_47922 (I816988,I817096,I817285);
nor I_47923 (I817395,I817268,I10431);
and I_47924 (I817412,I817395,I10431);
or I_47925 (I817429,I817412,I10437);
DFFARX1 I_47926 (I817429,I2683,I817005,I817455,);
nor I_47927 (I817463,I817455,I817189);
DFFARX1 I_47928 (I817463,I2683,I817005,I816976,);
nand I_47929 (I817494,I817455,I817096);
nand I_47930 (I817511,I817189,I817494);
nor I_47931 (I816985,I817511,I817155);
not I_47932 (I817566,I2690);
DFFARX1 I_47933 (I580373,I2683,I817566,I817592,);
DFFARX1 I_47934 (I817592,I2683,I817566,I817609,);
not I_47935 (I817558,I817609);
not I_47936 (I817631,I817592);
DFFARX1 I_47937 (I580385,I2683,I817566,I817657,);
nand I_47938 (I817665,I817657,I580394);
not I_47939 (I817682,I580394);
not I_47940 (I817699,I580376);
nand I_47941 (I817716,I580379,I580370);
and I_47942 (I817733,I580379,I580370);
not I_47943 (I817750,I580388);
nand I_47944 (I817767,I817750,I817699);
nor I_47945 (I817540,I817767,I817665);
nor I_47946 (I817798,I817682,I817767);
nand I_47947 (I817543,I817733,I817798);
not I_47948 (I817829,I580391);
nor I_47949 (I817846,I817829,I580379);
nor I_47950 (I817863,I817846,I580388);
nor I_47951 (I817880,I817631,I817863);
DFFARX1 I_47952 (I817880,I2683,I817566,I817552,);
not I_47953 (I817911,I817846);
DFFARX1 I_47954 (I817911,I2683,I817566,I817555,);
and I_47955 (I817549,I817657,I817846);
nor I_47956 (I817956,I817829,I580370);
and I_47957 (I817973,I817956,I580382);
or I_47958 (I817990,I817973,I580373);
DFFARX1 I_47959 (I817990,I2683,I817566,I818016,);
nor I_47960 (I818024,I818016,I817750);
DFFARX1 I_47961 (I818024,I2683,I817566,I817537,);
nand I_47962 (I818055,I818016,I817657);
nand I_47963 (I818072,I817750,I818055);
nor I_47964 (I817546,I818072,I817716);
not I_47965 (I818127,I2690);
DFFARX1 I_47966 (I901617,I2683,I818127,I818153,);
DFFARX1 I_47967 (I818153,I2683,I818127,I818170,);
not I_47968 (I818119,I818170);
not I_47969 (I818192,I818153);
DFFARX1 I_47970 (I901608,I2683,I818127,I818218,);
nand I_47971 (I818226,I818218,I901605);
not I_47972 (I818243,I901605);
not I_47973 (I818260,I901614);
nand I_47974 (I818277,I901623,I901605);
and I_47975 (I818294,I901623,I901605);
not I_47976 (I818311,I901602);
nand I_47977 (I818328,I818311,I818260);
nor I_47978 (I818101,I818328,I818226);
nor I_47979 (I818359,I818243,I818328);
nand I_47980 (I818104,I818294,I818359);
not I_47981 (I818390,I901611);
nor I_47982 (I818407,I818390,I901623);
nor I_47983 (I818424,I818407,I901602);
nor I_47984 (I818441,I818192,I818424);
DFFARX1 I_47985 (I818441,I2683,I818127,I818113,);
not I_47986 (I818472,I818407);
DFFARX1 I_47987 (I818472,I2683,I818127,I818116,);
and I_47988 (I818110,I818218,I818407);
nor I_47989 (I818517,I818390,I901626);
and I_47990 (I818534,I818517,I901602);
or I_47991 (I818551,I818534,I901620);
DFFARX1 I_47992 (I818551,I2683,I818127,I818577,);
nor I_47993 (I818585,I818577,I818311);
DFFARX1 I_47994 (I818585,I2683,I818127,I818098,);
nand I_47995 (I818616,I818577,I818218);
nand I_47996 (I818633,I818311,I818616);
nor I_47997 (I818107,I818633,I818277);
not I_47998 (I818688,I2690);
DFFARX1 I_47999 (I109652,I2683,I818688,I818714,);
DFFARX1 I_48000 (I818714,I2683,I818688,I818731,);
not I_48001 (I818680,I818731);
not I_48002 (I818753,I818714);
DFFARX1 I_48003 (I109640,I2683,I818688,I818779,);
nand I_48004 (I818787,I818779,I109655);
not I_48005 (I818804,I109655);
not I_48006 (I818821,I109643);
nand I_48007 (I818838,I109664,I109658);
and I_48008 (I818855,I109664,I109658);
not I_48009 (I818872,I109646);
nand I_48010 (I818889,I818872,I818821);
nor I_48011 (I818662,I818889,I818787);
nor I_48012 (I818920,I818804,I818889);
nand I_48013 (I818665,I818855,I818920);
not I_48014 (I818951,I109649);
nor I_48015 (I818968,I818951,I109664);
nor I_48016 (I818985,I818968,I109646);
nor I_48017 (I819002,I818753,I818985);
DFFARX1 I_48018 (I819002,I2683,I818688,I818674,);
not I_48019 (I819033,I818968);
DFFARX1 I_48020 (I819033,I2683,I818688,I818677,);
and I_48021 (I818671,I818779,I818968);
nor I_48022 (I819078,I818951,I109643);
and I_48023 (I819095,I819078,I109640);
or I_48024 (I819112,I819095,I109661);
DFFARX1 I_48025 (I819112,I2683,I818688,I819138,);
nor I_48026 (I819146,I819138,I818872);
DFFARX1 I_48027 (I819146,I2683,I818688,I818659,);
nand I_48028 (I819177,I819138,I818779);
nand I_48029 (I819194,I818872,I819177);
nor I_48030 (I818668,I819194,I818838);
not I_48031 (I819249,I2690);
DFFARX1 I_48032 (I831679,I2683,I819249,I819275,);
DFFARX1 I_48033 (I819275,I2683,I819249,I819292,);
not I_48034 (I819241,I819292);
not I_48035 (I819314,I819275);
DFFARX1 I_48036 (I831670,I2683,I819249,I819340,);
nand I_48037 (I819348,I819340,I831667);
not I_48038 (I819365,I831667);
not I_48039 (I819382,I831676);
nand I_48040 (I819399,I831685,I831667);
and I_48041 (I819416,I831685,I831667);
not I_48042 (I819433,I831664);
nand I_48043 (I819450,I819433,I819382);
nor I_48044 (I819223,I819450,I819348);
nor I_48045 (I819481,I819365,I819450);
nand I_48046 (I819226,I819416,I819481);
not I_48047 (I819512,I831673);
nor I_48048 (I819529,I819512,I831685);
nor I_48049 (I819546,I819529,I831664);
nor I_48050 (I819563,I819314,I819546);
DFFARX1 I_48051 (I819563,I2683,I819249,I819235,);
not I_48052 (I819594,I819529);
DFFARX1 I_48053 (I819594,I2683,I819249,I819238,);
and I_48054 (I819232,I819340,I819529);
nor I_48055 (I819639,I819512,I831688);
and I_48056 (I819656,I819639,I831664);
or I_48057 (I819673,I819656,I831682);
DFFARX1 I_48058 (I819673,I2683,I819249,I819699,);
nor I_48059 (I819707,I819699,I819433);
DFFARX1 I_48060 (I819707,I2683,I819249,I819220,);
nand I_48061 (I819738,I819699,I819340);
nand I_48062 (I819755,I819433,I819738);
nor I_48063 (I819229,I819755,I819399);
not I_48064 (I819810,I2690);
DFFARX1 I_48065 (I257510,I2683,I819810,I819836,);
DFFARX1 I_48066 (I819836,I2683,I819810,I819853,);
not I_48067 (I819802,I819853);
not I_48068 (I819875,I819836);
DFFARX1 I_48069 (I257507,I2683,I819810,I819901,);
nand I_48070 (I819909,I819901,I257501);
not I_48071 (I819926,I257501);
not I_48072 (I819943,I257498);
nand I_48073 (I819960,I257492,I257489);
and I_48074 (I819977,I257492,I257489);
not I_48075 (I819994,I257504);
nand I_48076 (I820011,I819994,I819943);
nor I_48077 (I819784,I820011,I819909);
nor I_48078 (I820042,I819926,I820011);
nand I_48079 (I819787,I819977,I820042);
not I_48080 (I820073,I257516);
nor I_48081 (I820090,I820073,I257492);
nor I_48082 (I820107,I820090,I257504);
nor I_48083 (I820124,I819875,I820107);
DFFARX1 I_48084 (I820124,I2683,I819810,I819796,);
not I_48085 (I820155,I820090);
DFFARX1 I_48086 (I820155,I2683,I819810,I819799,);
and I_48087 (I819793,I819901,I820090);
nor I_48088 (I820200,I820073,I257513);
and I_48089 (I820217,I820200,I257489);
or I_48090 (I820234,I820217,I257495);
DFFARX1 I_48091 (I820234,I2683,I819810,I820260,);
nor I_48092 (I820268,I820260,I819994);
DFFARX1 I_48093 (I820268,I2683,I819810,I819781,);
nand I_48094 (I820299,I820260,I819901);
nand I_48095 (I820316,I819994,I820299);
nor I_48096 (I819790,I820316,I819960);
not I_48097 (I820371,I2690);
DFFARX1 I_48098 (I624902,I2683,I820371,I820397,);
DFFARX1 I_48099 (I820397,I2683,I820371,I820414,);
not I_48100 (I820363,I820414);
not I_48101 (I820436,I820397);
DFFARX1 I_48102 (I624899,I2683,I820371,I820462,);
nand I_48103 (I820470,I820462,I624914);
not I_48104 (I820487,I624914);
not I_48105 (I820504,I624911);
nand I_48106 (I820521,I624908,I624896);
and I_48107 (I820538,I624908,I624896);
not I_48108 (I820555,I624893);
nand I_48109 (I820572,I820555,I820504);
nor I_48110 (I820345,I820572,I820470);
nor I_48111 (I820603,I820487,I820572);
nand I_48112 (I820348,I820538,I820603);
not I_48113 (I820634,I624899);
nor I_48114 (I820651,I820634,I624908);
nor I_48115 (I820668,I820651,I624893);
nor I_48116 (I820685,I820436,I820668);
DFFARX1 I_48117 (I820685,I2683,I820371,I820357,);
not I_48118 (I820716,I820651);
DFFARX1 I_48119 (I820716,I2683,I820371,I820360,);
and I_48120 (I820354,I820462,I820651);
nor I_48121 (I820761,I820634,I624905);
and I_48122 (I820778,I820761,I624893);
or I_48123 (I820795,I820778,I624896);
DFFARX1 I_48124 (I820795,I2683,I820371,I820821,);
nor I_48125 (I820829,I820821,I820555);
DFFARX1 I_48126 (I820829,I2683,I820371,I820342,);
nand I_48127 (I820860,I820821,I820462);
nand I_48128 (I820877,I820555,I820860);
nor I_48129 (I820351,I820877,I820521);
not I_48130 (I820932,I2690);
DFFARX1 I_48131 (I273320,I2683,I820932,I820958,);
DFFARX1 I_48132 (I820958,I2683,I820932,I820975,);
not I_48133 (I820924,I820975);
not I_48134 (I820997,I820958);
DFFARX1 I_48135 (I273317,I2683,I820932,I821023,);
nand I_48136 (I821031,I821023,I273311);
not I_48137 (I821048,I273311);
not I_48138 (I821065,I273308);
nand I_48139 (I821082,I273302,I273299);
and I_48140 (I821099,I273302,I273299);
not I_48141 (I821116,I273314);
nand I_48142 (I821133,I821116,I821065);
nor I_48143 (I820906,I821133,I821031);
nor I_48144 (I821164,I821048,I821133);
nand I_48145 (I820909,I821099,I821164);
not I_48146 (I821195,I273326);
nor I_48147 (I821212,I821195,I273302);
nor I_48148 (I821229,I821212,I273314);
nor I_48149 (I821246,I820997,I821229);
DFFARX1 I_48150 (I821246,I2683,I820932,I820918,);
not I_48151 (I821277,I821212);
DFFARX1 I_48152 (I821277,I2683,I820932,I820921,);
and I_48153 (I820915,I821023,I821212);
nor I_48154 (I821322,I821195,I273323);
and I_48155 (I821339,I821322,I273299);
or I_48156 (I821356,I821339,I273305);
DFFARX1 I_48157 (I821356,I2683,I820932,I821382,);
nor I_48158 (I821390,I821382,I821116);
DFFARX1 I_48159 (I821390,I2683,I820932,I820903,);
nand I_48160 (I821421,I821382,I821023);
nand I_48161 (I821438,I821116,I821421);
nor I_48162 (I820912,I821438,I821082);
not I_48163 (I821493,I2690);
DFFARX1 I_48164 (I943811,I2683,I821493,I821519,);
DFFARX1 I_48165 (I821519,I2683,I821493,I821536,);
not I_48166 (I821485,I821536);
not I_48167 (I821558,I821519);
DFFARX1 I_48168 (I943802,I2683,I821493,I821584,);
nand I_48169 (I821592,I821584,I943799);
not I_48170 (I821609,I943799);
not I_48171 (I821626,I943808);
nand I_48172 (I821643,I943817,I943799);
and I_48173 (I821660,I943817,I943799);
not I_48174 (I821677,I943796);
nand I_48175 (I821694,I821677,I821626);
nor I_48176 (I821467,I821694,I821592);
nor I_48177 (I821725,I821609,I821694);
nand I_48178 (I821470,I821660,I821725);
not I_48179 (I821756,I943805);
nor I_48180 (I821773,I821756,I943817);
nor I_48181 (I821790,I821773,I943796);
nor I_48182 (I821807,I821558,I821790);
DFFARX1 I_48183 (I821807,I2683,I821493,I821479,);
not I_48184 (I821838,I821773);
DFFARX1 I_48185 (I821838,I2683,I821493,I821482,);
and I_48186 (I821476,I821584,I821773);
nor I_48187 (I821883,I821756,I943820);
and I_48188 (I821900,I821883,I943796);
or I_48189 (I821917,I821900,I943814);
DFFARX1 I_48190 (I821917,I2683,I821493,I821943,);
nor I_48191 (I821951,I821943,I821677);
DFFARX1 I_48192 (I821951,I2683,I821493,I821464,);
nand I_48193 (I821982,I821943,I821584);
nand I_48194 (I821999,I821677,I821982);
nor I_48195 (I821473,I821999,I821643);
not I_48196 (I822054,I2690);
DFFARX1 I_48197 (I284387,I2683,I822054,I822080,);
DFFARX1 I_48198 (I822080,I2683,I822054,I822097,);
not I_48199 (I822046,I822097);
not I_48200 (I822119,I822080);
DFFARX1 I_48201 (I284384,I2683,I822054,I822145,);
nand I_48202 (I822153,I822145,I284378);
not I_48203 (I822170,I284378);
not I_48204 (I822187,I284375);
nand I_48205 (I822204,I284369,I284366);
and I_48206 (I822221,I284369,I284366);
not I_48207 (I822238,I284381);
nand I_48208 (I822255,I822238,I822187);
nor I_48209 (I822028,I822255,I822153);
nor I_48210 (I822286,I822170,I822255);
nand I_48211 (I822031,I822221,I822286);
not I_48212 (I822317,I284393);
nor I_48213 (I822334,I822317,I284369);
nor I_48214 (I822351,I822334,I284381);
nor I_48215 (I822368,I822119,I822351);
DFFARX1 I_48216 (I822368,I2683,I822054,I822040,);
not I_48217 (I822399,I822334);
DFFARX1 I_48218 (I822399,I2683,I822054,I822043,);
and I_48219 (I822037,I822145,I822334);
nor I_48220 (I822444,I822317,I284390);
and I_48221 (I822461,I822444,I284366);
or I_48222 (I822478,I822461,I284372);
DFFARX1 I_48223 (I822478,I2683,I822054,I822504,);
nor I_48224 (I822512,I822504,I822238);
DFFARX1 I_48225 (I822512,I2683,I822054,I822025,);
nand I_48226 (I822543,I822504,I822145);
nand I_48227 (I822560,I822238,I822543);
nor I_48228 (I822034,I822560,I822204);
not I_48229 (I822615,I2690);
DFFARX1 I_48230 (I346474,I2683,I822615,I822641,);
DFFARX1 I_48231 (I822641,I2683,I822615,I822658,);
not I_48232 (I822607,I822658);
not I_48233 (I822680,I822641);
DFFARX1 I_48234 (I346462,I2683,I822615,I822706,);
nand I_48235 (I822714,I822706,I346468);
not I_48236 (I822731,I346468);
not I_48237 (I822748,I346465);
nand I_48238 (I822765,I346453,I346450);
and I_48239 (I822782,I346453,I346450);
not I_48240 (I822799,I346477);
nand I_48241 (I822816,I822799,I822748);
nor I_48242 (I822589,I822816,I822714);
nor I_48243 (I822847,I822731,I822816);
nand I_48244 (I822592,I822782,I822847);
not I_48245 (I822878,I346450);
nor I_48246 (I822895,I822878,I346453);
nor I_48247 (I822912,I822895,I346477);
nor I_48248 (I822929,I822680,I822912);
DFFARX1 I_48249 (I822929,I2683,I822615,I822601,);
not I_48250 (I822960,I822895);
DFFARX1 I_48251 (I822960,I2683,I822615,I822604,);
and I_48252 (I822598,I822706,I822895);
nor I_48253 (I823005,I822878,I346459);
and I_48254 (I823022,I823005,I346456);
or I_48255 (I823039,I823022,I346471);
DFFARX1 I_48256 (I823039,I2683,I822615,I823065,);
nor I_48257 (I823073,I823065,I822799);
DFFARX1 I_48258 (I823073,I2683,I822615,I822586,);
nand I_48259 (I823104,I823065,I822706);
nand I_48260 (I823121,I822799,I823104);
nor I_48261 (I822595,I823121,I822765);
not I_48262 (I823176,I2690);
DFFARX1 I_48263 (I719345,I2683,I823176,I823202,);
DFFARX1 I_48264 (I823202,I2683,I823176,I823219,);
not I_48265 (I823168,I823219);
not I_48266 (I823241,I823202);
DFFARX1 I_48267 (I719372,I2683,I823176,I823267,);
nand I_48268 (I823275,I823267,I719363);
not I_48269 (I823292,I719363);
not I_48270 (I823309,I719345);
nand I_48271 (I823326,I719357,I719360);
and I_48272 (I823343,I719357,I719360);
not I_48273 (I823360,I719369);
nand I_48274 (I823377,I823360,I823309);
nor I_48275 (I823150,I823377,I823275);
nor I_48276 (I823408,I823292,I823377);
nand I_48277 (I823153,I823343,I823408);
not I_48278 (I823439,I719354);
nor I_48279 (I823456,I823439,I719357);
nor I_48280 (I823473,I823456,I719369);
nor I_48281 (I823490,I823241,I823473);
DFFARX1 I_48282 (I823490,I2683,I823176,I823162,);
not I_48283 (I823521,I823456);
DFFARX1 I_48284 (I823521,I2683,I823176,I823165,);
and I_48285 (I823159,I823267,I823456);
nor I_48286 (I823566,I823439,I719348);
and I_48287 (I823583,I823566,I719351);
or I_48288 (I823600,I823583,I719366);
DFFARX1 I_48289 (I823600,I2683,I823176,I823626,);
nor I_48290 (I823634,I823626,I823360);
DFFARX1 I_48291 (I823634,I2683,I823176,I823147,);
nand I_48292 (I823665,I823626,I823267);
nand I_48293 (I823682,I823360,I823665);
nor I_48294 (I823156,I823682,I823326);
not I_48295 (I823737,I2690);
DFFARX1 I_48296 (I168803,I2683,I823737,I823763,);
DFFARX1 I_48297 (I823763,I2683,I823737,I823780,);
not I_48298 (I823729,I823780);
not I_48299 (I823802,I823763);
DFFARX1 I_48300 (I168818,I2683,I823737,I823828,);
nand I_48301 (I823836,I823828,I168800);
not I_48302 (I823853,I168800);
not I_48303 (I823870,I168809);
nand I_48304 (I823887,I168815,I168806);
and I_48305 (I823904,I168815,I168806);
not I_48306 (I823921,I168803);
nand I_48307 (I823938,I823921,I823870);
nor I_48308 (I823711,I823938,I823836);
nor I_48309 (I823969,I823853,I823938);
nand I_48310 (I823714,I823904,I823969);
not I_48311 (I824000,I168800);
nor I_48312 (I824017,I824000,I168815);
nor I_48313 (I824034,I824017,I168803);
nor I_48314 (I824051,I823802,I824034);
DFFARX1 I_48315 (I824051,I2683,I823737,I823723,);
not I_48316 (I824082,I824017);
DFFARX1 I_48317 (I824082,I2683,I823737,I823726,);
and I_48318 (I823720,I823828,I824017);
nor I_48319 (I824127,I824000,I168824);
and I_48320 (I824144,I824127,I168821);
or I_48321 (I824161,I824144,I168812);
DFFARX1 I_48322 (I824161,I2683,I823737,I824187,);
nor I_48323 (I824195,I824187,I823921);
DFFARX1 I_48324 (I824195,I2683,I823737,I823708,);
nand I_48325 (I824226,I824187,I823828);
nand I_48326 (I824243,I823921,I824226);
nor I_48327 (I823717,I824243,I823887);
not I_48328 (I824298,I2690);
DFFARX1 I_48329 (I128343,I2683,I824298,I824324,);
DFFARX1 I_48330 (I824324,I2683,I824298,I824341,);
not I_48331 (I824290,I824341);
not I_48332 (I824363,I824324);
DFFARX1 I_48333 (I128358,I2683,I824298,I824389,);
nand I_48334 (I824397,I824389,I128340);
not I_48335 (I824414,I128340);
not I_48336 (I824431,I128349);
nand I_48337 (I824448,I128355,I128346);
and I_48338 (I824465,I128355,I128346);
not I_48339 (I824482,I128343);
nand I_48340 (I824499,I824482,I824431);
nor I_48341 (I824272,I824499,I824397);
nor I_48342 (I824530,I824414,I824499);
nand I_48343 (I824275,I824465,I824530);
not I_48344 (I824561,I128340);
nor I_48345 (I824578,I824561,I128355);
nor I_48346 (I824595,I824578,I128343);
nor I_48347 (I824612,I824363,I824595);
DFFARX1 I_48348 (I824612,I2683,I824298,I824284,);
not I_48349 (I824643,I824578);
DFFARX1 I_48350 (I824643,I2683,I824298,I824287,);
and I_48351 (I824281,I824389,I824578);
nor I_48352 (I824688,I824561,I128364);
and I_48353 (I824705,I824688,I128361);
or I_48354 (I824722,I824705,I128352);
DFFARX1 I_48355 (I824722,I2683,I824298,I824748,);
nor I_48356 (I824756,I824748,I824482);
DFFARX1 I_48357 (I824756,I2683,I824298,I824269,);
nand I_48358 (I824787,I824748,I824389);
nand I_48359 (I824804,I824482,I824787);
nor I_48360 (I824278,I824804,I824448);
not I_48361 (I824859,I2690);
DFFARX1 I_48362 (I767149,I2683,I824859,I824885,);
DFFARX1 I_48363 (I824885,I2683,I824859,I824902,);
not I_48364 (I824851,I824902);
not I_48365 (I824924,I824885);
DFFARX1 I_48366 (I767176,I2683,I824859,I824950,);
nand I_48367 (I824958,I824950,I767167);
not I_48368 (I824975,I767167);
not I_48369 (I824992,I767149);
nand I_48370 (I825009,I767161,I767164);
and I_48371 (I825026,I767161,I767164);
not I_48372 (I825043,I767173);
nand I_48373 (I825060,I825043,I824992);
nor I_48374 (I824833,I825060,I824958);
nor I_48375 (I825091,I824975,I825060);
nand I_48376 (I824836,I825026,I825091);
not I_48377 (I825122,I767158);
nor I_48378 (I825139,I825122,I767161);
nor I_48379 (I825156,I825139,I767173);
nor I_48380 (I825173,I824924,I825156);
DFFARX1 I_48381 (I825173,I2683,I824859,I824845,);
not I_48382 (I825204,I825139);
DFFARX1 I_48383 (I825204,I2683,I824859,I824848,);
and I_48384 (I824842,I824950,I825139);
nor I_48385 (I825249,I825122,I767152);
and I_48386 (I825266,I825249,I767155);
or I_48387 (I825283,I825266,I767170);
DFFARX1 I_48388 (I825283,I2683,I824859,I825309,);
nor I_48389 (I825317,I825309,I825043);
DFFARX1 I_48390 (I825317,I2683,I824859,I824830,);
nand I_48391 (I825348,I825309,I824950);
nand I_48392 (I825365,I825043,I825348);
nor I_48393 (I824839,I825365,I825009);
not I_48394 (I825420,I2690);
DFFARX1 I_48395 (I1070954,I2683,I825420,I825446,);
DFFARX1 I_48396 (I825446,I2683,I825420,I825463,);
not I_48397 (I825412,I825463);
not I_48398 (I825485,I825446);
DFFARX1 I_48399 (I1070948,I2683,I825420,I825511,);
nand I_48400 (I825519,I825511,I1070939);
not I_48401 (I825536,I1070939);
not I_48402 (I825553,I1070966);
nand I_48403 (I825570,I1070951,I1070960);
and I_48404 (I825587,I1070951,I1070960);
not I_48405 (I825604,I1070945);
nand I_48406 (I825621,I825604,I825553);
nor I_48407 (I825394,I825621,I825519);
nor I_48408 (I825652,I825536,I825621);
nand I_48409 (I825397,I825587,I825652);
not I_48410 (I825683,I1070963);
nor I_48411 (I825700,I825683,I1070951);
nor I_48412 (I825717,I825700,I1070945);
nor I_48413 (I825734,I825485,I825717);
DFFARX1 I_48414 (I825734,I2683,I825420,I825406,);
not I_48415 (I825765,I825700);
DFFARX1 I_48416 (I825765,I2683,I825420,I825409,);
and I_48417 (I825403,I825511,I825700);
nor I_48418 (I825810,I825683,I1070957);
and I_48419 (I825827,I825810,I1070939);
or I_48420 (I825844,I825827,I1070942);
DFFARX1 I_48421 (I825844,I2683,I825420,I825870,);
nor I_48422 (I825878,I825870,I825604);
DFFARX1 I_48423 (I825878,I2683,I825420,I825391,);
nand I_48424 (I825909,I825870,I825511);
nand I_48425 (I825926,I825604,I825909);
nor I_48426 (I825400,I825926,I825570);
not I_48427 (I825981,I2690);
DFFARX1 I_48428 (I1024890,I2683,I825981,I826007,);
DFFARX1 I_48429 (I826007,I2683,I825981,I826024,);
not I_48430 (I825973,I826024);
not I_48431 (I826046,I826007);
DFFARX1 I_48432 (I1024875,I2683,I825981,I826072,);
nand I_48433 (I826080,I826072,I1024884);
not I_48434 (I826097,I1024884);
not I_48435 (I826114,I1024878);
nand I_48436 (I826131,I1024896,I1024893);
and I_48437 (I826148,I1024896,I1024893);
not I_48438 (I826165,I1024869);
nand I_48439 (I826182,I826165,I826114);
nor I_48440 (I825955,I826182,I826080);
nor I_48441 (I826213,I826097,I826182);
nand I_48442 (I825958,I826148,I826213);
not I_48443 (I826244,I1024872);
nor I_48444 (I826261,I826244,I1024896);
nor I_48445 (I826278,I826261,I1024869);
nor I_48446 (I826295,I826046,I826278);
DFFARX1 I_48447 (I826295,I2683,I825981,I825967,);
not I_48448 (I826326,I826261);
DFFARX1 I_48449 (I826326,I2683,I825981,I825970,);
and I_48450 (I825964,I826072,I826261);
nor I_48451 (I826371,I826244,I1024869);
and I_48452 (I826388,I826371,I1024887);
or I_48453 (I826405,I826388,I1024881);
DFFARX1 I_48454 (I826405,I2683,I825981,I826431,);
nor I_48455 (I826439,I826431,I826165);
DFFARX1 I_48456 (I826439,I2683,I825981,I825952,);
nand I_48457 (I826470,I826431,I826072);
nand I_48458 (I826487,I826165,I826470);
nor I_48459 (I825961,I826487,I826131);
not I_48460 (I826542,I2690);
DFFARX1 I_48461 (I1005917,I2683,I826542,I826568,);
DFFARX1 I_48462 (I826568,I2683,I826542,I826585,);
not I_48463 (I826534,I826585);
not I_48464 (I826607,I826568);
DFFARX1 I_48465 (I1005914,I2683,I826542,I826633,);
nand I_48466 (I826641,I826633,I1005920);
not I_48467 (I826658,I1005920);
not I_48468 (I826675,I1005929);
nand I_48469 (I826692,I1005923,I1005917);
and I_48470 (I826709,I1005923,I1005917);
not I_48471 (I826726,I1005935);
nand I_48472 (I826743,I826726,I826675);
nor I_48473 (I826516,I826743,I826641);
nor I_48474 (I826774,I826658,I826743);
nand I_48475 (I826519,I826709,I826774);
not I_48476 (I826805,I1005932);
nor I_48477 (I826822,I826805,I1005923);
nor I_48478 (I826839,I826822,I1005935);
nor I_48479 (I826856,I826607,I826839);
DFFARX1 I_48480 (I826856,I2683,I826542,I826528,);
not I_48481 (I826887,I826822);
DFFARX1 I_48482 (I826887,I2683,I826542,I826531,);
and I_48483 (I826525,I826633,I826822);
nor I_48484 (I826932,I826805,I1005926);
and I_48485 (I826949,I826932,I1005938);
or I_48486 (I826966,I826949,I1005914);
DFFARX1 I_48487 (I826966,I2683,I826542,I826992,);
nor I_48488 (I827000,I826992,I826726);
DFFARX1 I_48489 (I827000,I2683,I826542,I826513,);
nand I_48490 (I827031,I826992,I826633);
nand I_48491 (I827048,I826726,I827031);
nor I_48492 (I826522,I827048,I826692);
not I_48493 (I827103,I2690);
DFFARX1 I_48494 (I250132,I2683,I827103,I827129,);
DFFARX1 I_48495 (I827129,I2683,I827103,I827146,);
not I_48496 (I827095,I827146);
not I_48497 (I827168,I827129);
DFFARX1 I_48498 (I250129,I2683,I827103,I827194,);
nand I_48499 (I827202,I827194,I250123);
not I_48500 (I827219,I250123);
not I_48501 (I827236,I250120);
nand I_48502 (I827253,I250114,I250111);
and I_48503 (I827270,I250114,I250111);
not I_48504 (I827287,I250126);
nand I_48505 (I827304,I827287,I827236);
nor I_48506 (I827077,I827304,I827202);
nor I_48507 (I827335,I827219,I827304);
nand I_48508 (I827080,I827270,I827335);
not I_48509 (I827366,I250138);
nor I_48510 (I827383,I827366,I250114);
nor I_48511 (I827400,I827383,I250126);
nor I_48512 (I827417,I827168,I827400);
DFFARX1 I_48513 (I827417,I2683,I827103,I827089,);
not I_48514 (I827448,I827383);
DFFARX1 I_48515 (I827448,I2683,I827103,I827092,);
and I_48516 (I827086,I827194,I827383);
nor I_48517 (I827493,I827366,I250135);
and I_48518 (I827510,I827493,I250111);
or I_48519 (I827527,I827510,I250117);
DFFARX1 I_48520 (I827527,I2683,I827103,I827553,);
nor I_48521 (I827561,I827553,I827287);
DFFARX1 I_48522 (I827561,I2683,I827103,I827074,);
nand I_48523 (I827592,I827553,I827194);
nand I_48524 (I827609,I827287,I827592);
nor I_48525 (I827083,I827609,I827253);
not I_48526 (I827664,I2690);
DFFARX1 I_48527 (I833413,I2683,I827664,I827690,);
DFFARX1 I_48528 (I827690,I2683,I827664,I827707,);
not I_48529 (I827656,I827707);
not I_48530 (I827729,I827690);
DFFARX1 I_48531 (I833404,I2683,I827664,I827755,);
nand I_48532 (I827763,I827755,I833401);
not I_48533 (I827780,I833401);
not I_48534 (I827797,I833410);
nand I_48535 (I827814,I833419,I833401);
and I_48536 (I827831,I833419,I833401);
not I_48537 (I827848,I833398);
nand I_48538 (I827865,I827848,I827797);
nor I_48539 (I827638,I827865,I827763);
nor I_48540 (I827896,I827780,I827865);
nand I_48541 (I827641,I827831,I827896);
not I_48542 (I827927,I833407);
nor I_48543 (I827944,I827927,I833419);
nor I_48544 (I827961,I827944,I833398);
nor I_48545 (I827978,I827729,I827961);
DFFARX1 I_48546 (I827978,I2683,I827664,I827650,);
not I_48547 (I828009,I827944);
DFFARX1 I_48548 (I828009,I2683,I827664,I827653,);
and I_48549 (I827647,I827755,I827944);
nor I_48550 (I828054,I827927,I833422);
and I_48551 (I828071,I828054,I833398);
or I_48552 (I828088,I828071,I833416);
DFFARX1 I_48553 (I828088,I2683,I827664,I828114,);
nor I_48554 (I828122,I828114,I827848);
DFFARX1 I_48555 (I828122,I2683,I827664,I827635,);
nand I_48556 (I828153,I828114,I827755);
nand I_48557 (I828170,I827848,I828153);
nor I_48558 (I827644,I828170,I827814);
not I_48559 (I828228,I2690);
DFFARX1 I_48560 (I107556,I2683,I828228,I828254,);
and I_48561 (I828262,I828254,I107532);
DFFARX1 I_48562 (I828262,I2683,I828228,I828211,);
DFFARX1 I_48563 (I107550,I2683,I828228,I828302,);
not I_48564 (I828310,I107538);
not I_48565 (I828327,I107535);
nand I_48566 (I828344,I828327,I828310);
nor I_48567 (I828199,I828302,I828344);
DFFARX1 I_48568 (I828344,I2683,I828228,I828384,);
not I_48569 (I828220,I828384);
not I_48570 (I828406,I107544);
nand I_48571 (I828423,I828327,I828406);
DFFARX1 I_48572 (I828423,I2683,I828228,I828449,);
not I_48573 (I828457,I828449);
not I_48574 (I828474,I107535);
nand I_48575 (I828491,I828474,I107553);
and I_48576 (I828508,I828310,I828491);
nor I_48577 (I828525,I828423,I828508);
DFFARX1 I_48578 (I828525,I2683,I828228,I828196,);
DFFARX1 I_48579 (I828508,I2683,I828228,I828217,);
nor I_48580 (I828570,I107535,I107547);
nor I_48581 (I828208,I828423,I828570);
or I_48582 (I828601,I107535,I107547);
nor I_48583 (I828618,I107541,I107532);
DFFARX1 I_48584 (I828618,I2683,I828228,I828644,);
not I_48585 (I828652,I828644);
nor I_48586 (I828214,I828652,I828457);
nand I_48587 (I828683,I828652,I828302);
not I_48588 (I828700,I107541);
nand I_48589 (I828717,I828700,I828406);
nand I_48590 (I828734,I828652,I828717);
nand I_48591 (I828205,I828734,I828683);
nand I_48592 (I828202,I828717,I828601);
not I_48593 (I828806,I2690);
DFFARX1 I_48594 (I118820,I2683,I828806,I828832,);
and I_48595 (I828840,I828832,I118844);
DFFARX1 I_48596 (I828840,I2683,I828806,I828789,);
DFFARX1 I_48597 (I118820,I2683,I828806,I828880,);
not I_48598 (I828888,I118838);
not I_48599 (I828905,I118823);
nand I_48600 (I828922,I828905,I828888);
nor I_48601 (I828777,I828880,I828922);
DFFARX1 I_48602 (I828922,I2683,I828806,I828962,);
not I_48603 (I828798,I828962);
not I_48604 (I828984,I118832);
nand I_48605 (I829001,I828905,I828984);
DFFARX1 I_48606 (I829001,I2683,I828806,I829027,);
not I_48607 (I829035,I829027);
not I_48608 (I829052,I118829);
nand I_48609 (I829069,I829052,I118826);
and I_48610 (I829086,I828888,I829069);
nor I_48611 (I829103,I829001,I829086);
DFFARX1 I_48612 (I829103,I2683,I828806,I828774,);
DFFARX1 I_48613 (I829086,I2683,I828806,I828795,);
nor I_48614 (I829148,I118829,I118835);
nor I_48615 (I828786,I829001,I829148);
or I_48616 (I829179,I118829,I118835);
nor I_48617 (I829196,I118841,I118847);
DFFARX1 I_48618 (I829196,I2683,I828806,I829222,);
not I_48619 (I829230,I829222);
nor I_48620 (I828792,I829230,I829035);
nand I_48621 (I829261,I829230,I828880);
not I_48622 (I829278,I118841);
nand I_48623 (I829295,I829278,I828984);
nand I_48624 (I829312,I829230,I829295);
nand I_48625 (I828783,I829312,I829261);
nand I_48626 (I828780,I829295,I829179);
not I_48627 (I829384,I2690);
DFFARX1 I_48628 (I512759,I2683,I829384,I829410,);
and I_48629 (I829418,I829410,I512747);
DFFARX1 I_48630 (I829418,I2683,I829384,I829367,);
DFFARX1 I_48631 (I512750,I2683,I829384,I829458,);
not I_48632 (I829466,I512744);
not I_48633 (I829483,I512768);
nand I_48634 (I829500,I829483,I829466);
nor I_48635 (I829355,I829458,I829500);
DFFARX1 I_48636 (I829500,I2683,I829384,I829540,);
not I_48637 (I829376,I829540);
not I_48638 (I829562,I512756);
nand I_48639 (I829579,I829483,I829562);
DFFARX1 I_48640 (I829579,I2683,I829384,I829605,);
not I_48641 (I829613,I829605);
not I_48642 (I829630,I512765);
nand I_48643 (I829647,I829630,I512762);
and I_48644 (I829664,I829466,I829647);
nor I_48645 (I829681,I829579,I829664);
DFFARX1 I_48646 (I829681,I2683,I829384,I829352,);
DFFARX1 I_48647 (I829664,I2683,I829384,I829373,);
nor I_48648 (I829726,I512765,I512753);
nor I_48649 (I829364,I829579,I829726);
or I_48650 (I829757,I512765,I512753);
nor I_48651 (I829774,I512744,I512747);
DFFARX1 I_48652 (I829774,I2683,I829384,I829800,);
not I_48653 (I829808,I829800);
nor I_48654 (I829370,I829808,I829613);
nand I_48655 (I829839,I829808,I829458);
not I_48656 (I829856,I512744);
nand I_48657 (I829873,I829856,I829562);
nand I_48658 (I829890,I829808,I829873);
nand I_48659 (I829361,I829890,I829839);
nand I_48660 (I829358,I829873,I829757);
not I_48661 (I829962,I2690);
DFFARX1 I_48662 (I553219,I2683,I829962,I829988,);
and I_48663 (I829996,I829988,I553207);
DFFARX1 I_48664 (I829996,I2683,I829962,I829945,);
DFFARX1 I_48665 (I553210,I2683,I829962,I830036,);
not I_48666 (I830044,I553204);
not I_48667 (I830061,I553228);
nand I_48668 (I830078,I830061,I830044);
nor I_48669 (I829933,I830036,I830078);
DFFARX1 I_48670 (I830078,I2683,I829962,I830118,);
not I_48671 (I829954,I830118);
not I_48672 (I830140,I553216);
nand I_48673 (I830157,I830061,I830140);
DFFARX1 I_48674 (I830157,I2683,I829962,I830183,);
not I_48675 (I830191,I830183);
not I_48676 (I830208,I553225);
nand I_48677 (I830225,I830208,I553222);
and I_48678 (I830242,I830044,I830225);
nor I_48679 (I830259,I830157,I830242);
DFFARX1 I_48680 (I830259,I2683,I829962,I829930,);
DFFARX1 I_48681 (I830242,I2683,I829962,I829951,);
nor I_48682 (I830304,I553225,I553213);
nor I_48683 (I829942,I830157,I830304);
or I_48684 (I830335,I553225,I553213);
nor I_48685 (I830352,I553204,I553207);
DFFARX1 I_48686 (I830352,I2683,I829962,I830378,);
not I_48687 (I830386,I830378);
nor I_48688 (I829948,I830386,I830191);
nand I_48689 (I830417,I830386,I830036);
not I_48690 (I830434,I553204);
nand I_48691 (I830451,I830434,I830140);
nand I_48692 (I830468,I830386,I830451);
nand I_48693 (I829939,I830468,I830417);
nand I_48694 (I829936,I830451,I830335);
not I_48695 (I830540,I2690);
DFFARX1 I_48696 (I965203,I2683,I830540,I830566,);
and I_48697 (I830574,I830566,I965197);
DFFARX1 I_48698 (I830574,I2683,I830540,I830523,);
DFFARX1 I_48699 (I965182,I2683,I830540,I830614,);
not I_48700 (I830622,I965188);
not I_48701 (I830639,I965200);
nand I_48702 (I830656,I830639,I830622);
nor I_48703 (I830511,I830614,I830656);
DFFARX1 I_48704 (I830656,I2683,I830540,I830696,);
not I_48705 (I830532,I830696);
not I_48706 (I830718,I965182);
nand I_48707 (I830735,I830639,I830718);
DFFARX1 I_48708 (I830735,I2683,I830540,I830761,);
not I_48709 (I830769,I830761);
not I_48710 (I830786,I965206);
nand I_48711 (I830803,I830786,I965194);
and I_48712 (I830820,I830622,I830803);
nor I_48713 (I830837,I830735,I830820);
DFFARX1 I_48714 (I830837,I2683,I830540,I830508,);
DFFARX1 I_48715 (I830820,I2683,I830540,I830529,);
nor I_48716 (I830882,I965206,I965185);
nor I_48717 (I830520,I830735,I830882);
or I_48718 (I830913,I965206,I965185);
nor I_48719 (I830930,I965191,I965185);
DFFARX1 I_48720 (I830930,I2683,I830540,I830956,);
not I_48721 (I830964,I830956);
nor I_48722 (I830526,I830964,I830769);
nand I_48723 (I830995,I830964,I830614);
not I_48724 (I831012,I965191);
nand I_48725 (I831029,I831012,I830718);
nand I_48726 (I831046,I830964,I831029);
nand I_48727 (I830517,I831046,I830995);
nand I_48728 (I830514,I831029,I830913);
not I_48729 (I831118,I2690);
DFFARX1 I_48730 (I383986,I2683,I831118,I831144,);
and I_48731 (I831152,I831144,I384001);
DFFARX1 I_48732 (I831152,I2683,I831118,I831101,);
DFFARX1 I_48733 (I384004,I2683,I831118,I831192,);
not I_48734 (I831200,I383998);
not I_48735 (I831217,I384013);
nand I_48736 (I831234,I831217,I831200);
nor I_48737 (I831089,I831192,I831234);
DFFARX1 I_48738 (I831234,I2683,I831118,I831274,);
not I_48739 (I831110,I831274);
not I_48740 (I831296,I383989);
nand I_48741 (I831313,I831217,I831296);
DFFARX1 I_48742 (I831313,I2683,I831118,I831339,);
not I_48743 (I831347,I831339);
not I_48744 (I831364,I383992);
nand I_48745 (I831381,I831364,I383986);
and I_48746 (I831398,I831200,I831381);
nor I_48747 (I831415,I831313,I831398);
DFFARX1 I_48748 (I831415,I2683,I831118,I831086,);
DFFARX1 I_48749 (I831398,I2683,I831118,I831107,);
nor I_48750 (I831460,I383992,I383995);
nor I_48751 (I831098,I831313,I831460);
or I_48752 (I831491,I383992,I383995);
nor I_48753 (I831508,I384010,I384007);
DFFARX1 I_48754 (I831508,I2683,I831118,I831534,);
not I_48755 (I831542,I831534);
nor I_48756 (I831104,I831542,I831347);
nand I_48757 (I831573,I831542,I831192);
not I_48758 (I831590,I384010);
nand I_48759 (I831607,I831590,I831296);
nand I_48760 (I831624,I831542,I831607);
nand I_48761 (I831095,I831624,I831573);
nand I_48762 (I831092,I831607,I831491);
not I_48763 (I831696,I2690);
DFFARX1 I_48764 (I706431,I2683,I831696,I831722,);
and I_48765 (I831730,I831722,I706425);
DFFARX1 I_48766 (I831730,I2683,I831696,I831679,);
DFFARX1 I_48767 (I706443,I2683,I831696,I831770,);
not I_48768 (I831778,I706434);
not I_48769 (I831795,I706446);
nand I_48770 (I831812,I831795,I831778);
nor I_48771 (I831667,I831770,I831812);
DFFARX1 I_48772 (I831812,I2683,I831696,I831852,);
not I_48773 (I831688,I831852);
not I_48774 (I831874,I706452);
nand I_48775 (I831891,I831795,I831874);
DFFARX1 I_48776 (I831891,I2683,I831696,I831917,);
not I_48777 (I831925,I831917);
not I_48778 (I831942,I706428);
nand I_48779 (I831959,I831942,I706449);
and I_48780 (I831976,I831778,I831959);
nor I_48781 (I831993,I831891,I831976);
DFFARX1 I_48782 (I831993,I2683,I831696,I831664,);
DFFARX1 I_48783 (I831976,I2683,I831696,I831685,);
nor I_48784 (I832038,I706428,I706440);
nor I_48785 (I831676,I831891,I832038);
or I_48786 (I832069,I706428,I706440);
nor I_48787 (I832086,I706425,I706437);
DFFARX1 I_48788 (I832086,I2683,I831696,I832112,);
not I_48789 (I832120,I832112);
nor I_48790 (I831682,I832120,I831925);
nand I_48791 (I832151,I832120,I831770);
not I_48792 (I832168,I706425);
nand I_48793 (I832185,I832168,I831874);
nand I_48794 (I832202,I832120,I832185);
nand I_48795 (I831673,I832202,I832151);
nand I_48796 (I831670,I832185,I832069);
not I_48797 (I832274,I2690);
DFFARX1 I_48798 (I443399,I2683,I832274,I832300,);
and I_48799 (I832308,I832300,I443387);
DFFARX1 I_48800 (I832308,I2683,I832274,I832257,);
DFFARX1 I_48801 (I443402,I2683,I832274,I832348,);
not I_48802 (I832356,I443393);
not I_48803 (I832373,I443384);
nand I_48804 (I832390,I832373,I832356);
nor I_48805 (I832245,I832348,I832390);
DFFARX1 I_48806 (I832390,I2683,I832274,I832430,);
not I_48807 (I832266,I832430);
not I_48808 (I832452,I443390);
nand I_48809 (I832469,I832373,I832452);
DFFARX1 I_48810 (I832469,I2683,I832274,I832495,);
not I_48811 (I832503,I832495);
not I_48812 (I832520,I443405);
nand I_48813 (I832537,I832520,I443408);
and I_48814 (I832554,I832356,I832537);
nor I_48815 (I832571,I832469,I832554);
DFFARX1 I_48816 (I832571,I2683,I832274,I832242,);
DFFARX1 I_48817 (I832554,I2683,I832274,I832263,);
nor I_48818 (I832616,I443405,I443384);
nor I_48819 (I832254,I832469,I832616);
or I_48820 (I832647,I443405,I443384);
nor I_48821 (I832664,I443396,I443387);
DFFARX1 I_48822 (I832664,I2683,I832274,I832690,);
not I_48823 (I832698,I832690);
nor I_48824 (I832260,I832698,I832503);
nand I_48825 (I832729,I832698,I832348);
not I_48826 (I832746,I443396);
nand I_48827 (I832763,I832746,I832452);
nand I_48828 (I832780,I832698,I832763);
nand I_48829 (I832251,I832780,I832729);
nand I_48830 (I832248,I832763,I832647);
not I_48831 (I832852,I2690);
DFFARX1 I_48832 (I800149,I2683,I832852,I832878,);
and I_48833 (I832886,I832878,I800146);
DFFARX1 I_48834 (I832886,I2683,I832852,I832835,);
DFFARX1 I_48835 (I800152,I2683,I832852,I832926,);
not I_48836 (I832934,I800155);
not I_48837 (I832951,I800149);
nand I_48838 (I832968,I832951,I832934);
nor I_48839 (I832823,I832926,I832968);
DFFARX1 I_48840 (I832968,I2683,I832852,I833008,);
not I_48841 (I832844,I833008);
not I_48842 (I833030,I800164);
nand I_48843 (I833047,I832951,I833030);
DFFARX1 I_48844 (I833047,I2683,I832852,I833073,);
not I_48845 (I833081,I833073);
not I_48846 (I833098,I800161);
nand I_48847 (I833115,I833098,I800167);
and I_48848 (I833132,I832934,I833115);
nor I_48849 (I833149,I833047,I833132);
DFFARX1 I_48850 (I833149,I2683,I832852,I832820,);
DFFARX1 I_48851 (I833132,I2683,I832852,I832841,);
nor I_48852 (I833194,I800161,I800146);
nor I_48853 (I832832,I833047,I833194);
or I_48854 (I833225,I800161,I800146);
nor I_48855 (I833242,I800158,I800152);
DFFARX1 I_48856 (I833242,I2683,I832852,I833268,);
not I_48857 (I833276,I833268);
nor I_48858 (I832838,I833276,I833081);
nand I_48859 (I833307,I833276,I832926);
not I_48860 (I833324,I800158);
nand I_48861 (I833341,I833324,I833030);
nand I_48862 (I833358,I833276,I833341);
nand I_48863 (I832829,I833358,I833307);
nand I_48864 (I832826,I833341,I833225);
not I_48865 (I833430,I2690);
DFFARX1 I_48866 (I72247,I2683,I833430,I833456,);
and I_48867 (I833464,I833456,I72223);
DFFARX1 I_48868 (I833464,I2683,I833430,I833413,);
DFFARX1 I_48869 (I72241,I2683,I833430,I833504,);
not I_48870 (I833512,I72229);
not I_48871 (I833529,I72226);
nand I_48872 (I833546,I833529,I833512);
nor I_48873 (I833401,I833504,I833546);
DFFARX1 I_48874 (I833546,I2683,I833430,I833586,);
not I_48875 (I833422,I833586);
not I_48876 (I833608,I72235);
nand I_48877 (I833625,I833529,I833608);
DFFARX1 I_48878 (I833625,I2683,I833430,I833651,);
not I_48879 (I833659,I833651);
not I_48880 (I833676,I72226);
nand I_48881 (I833693,I833676,I72244);
and I_48882 (I833710,I833512,I833693);
nor I_48883 (I833727,I833625,I833710);
DFFARX1 I_48884 (I833727,I2683,I833430,I833398,);
DFFARX1 I_48885 (I833710,I2683,I833430,I833419,);
nor I_48886 (I833772,I72226,I72238);
nor I_48887 (I833410,I833625,I833772);
or I_48888 (I833803,I72226,I72238);
nor I_48889 (I833820,I72232,I72223);
DFFARX1 I_48890 (I833820,I2683,I833430,I833846,);
not I_48891 (I833854,I833846);
nor I_48892 (I833416,I833854,I833659);
nand I_48893 (I833885,I833854,I833504);
not I_48894 (I833902,I72232);
nand I_48895 (I833919,I833902,I833608);
nand I_48896 (I833936,I833854,I833919);
nand I_48897 (I833407,I833936,I833885);
nand I_48898 (I833404,I833919,I833803);
not I_48899 (I834008,I2690);
DFFARX1 I_48900 (I653354,I2683,I834008,I834034,);
and I_48901 (I834042,I834034,I653360);
DFFARX1 I_48902 (I834042,I2683,I834008,I833991,);
DFFARX1 I_48903 (I653366,I2683,I834008,I834082,);
not I_48904 (I834090,I653351);
not I_48905 (I834107,I653351);
nand I_48906 (I834124,I834107,I834090);
nor I_48907 (I833979,I834082,I834124);
DFFARX1 I_48908 (I834124,I2683,I834008,I834164,);
not I_48909 (I834000,I834164);
not I_48910 (I834186,I653369);
nand I_48911 (I834203,I834107,I834186);
DFFARX1 I_48912 (I834203,I2683,I834008,I834229,);
not I_48913 (I834237,I834229);
not I_48914 (I834254,I653363);
nand I_48915 (I834271,I834254,I653354);
and I_48916 (I834288,I834090,I834271);
nor I_48917 (I834305,I834203,I834288);
DFFARX1 I_48918 (I834305,I2683,I834008,I833976,);
DFFARX1 I_48919 (I834288,I2683,I834008,I833997,);
nor I_48920 (I834350,I653363,I653372);
nor I_48921 (I833988,I834203,I834350);
or I_48922 (I834381,I653363,I653372);
nor I_48923 (I834398,I653357,I653357);
DFFARX1 I_48924 (I834398,I2683,I834008,I834424,);
not I_48925 (I834432,I834424);
nor I_48926 (I833994,I834432,I834237);
nand I_48927 (I834463,I834432,I834082);
not I_48928 (I834480,I653357);
nand I_48929 (I834497,I834480,I834186);
nand I_48930 (I834514,I834432,I834497);
nand I_48931 (I833985,I834514,I834463);
nand I_48932 (I833982,I834497,I834381);
not I_48933 (I834586,I2690);
DFFARX1 I_48934 (I543971,I2683,I834586,I834612,);
and I_48935 (I834620,I834612,I543959);
DFFARX1 I_48936 (I834620,I2683,I834586,I834569,);
DFFARX1 I_48937 (I543962,I2683,I834586,I834660,);
not I_48938 (I834668,I543956);
not I_48939 (I834685,I543980);
nand I_48940 (I834702,I834685,I834668);
nor I_48941 (I834557,I834660,I834702);
DFFARX1 I_48942 (I834702,I2683,I834586,I834742,);
not I_48943 (I834578,I834742);
not I_48944 (I834764,I543968);
nand I_48945 (I834781,I834685,I834764);
DFFARX1 I_48946 (I834781,I2683,I834586,I834807,);
not I_48947 (I834815,I834807);
not I_48948 (I834832,I543977);
nand I_48949 (I834849,I834832,I543974);
and I_48950 (I834866,I834668,I834849);
nor I_48951 (I834883,I834781,I834866);
DFFARX1 I_48952 (I834883,I2683,I834586,I834554,);
DFFARX1 I_48953 (I834866,I2683,I834586,I834575,);
nor I_48954 (I834928,I543977,I543965);
nor I_48955 (I834566,I834781,I834928);
or I_48956 (I834959,I543977,I543965);
nor I_48957 (I834976,I543956,I543959);
DFFARX1 I_48958 (I834976,I2683,I834586,I835002,);
not I_48959 (I835010,I835002);
nor I_48960 (I834572,I835010,I834815);
nand I_48961 (I835041,I835010,I834660);
not I_48962 (I835058,I543956);
nand I_48963 (I835075,I835058,I834764);
nand I_48964 (I835092,I835010,I835075);
nand I_48965 (I834563,I835092,I835041);
nand I_48966 (I834560,I835075,I834959);
not I_48967 (I835164,I2690);
DFFARX1 I_48968 (I255408,I2683,I835164,I835190,);
and I_48969 (I835198,I835190,I255393);
DFFARX1 I_48970 (I835198,I2683,I835164,I835147,);
DFFARX1 I_48971 (I255399,I2683,I835164,I835238,);
not I_48972 (I835246,I255381);
not I_48973 (I835263,I255402);
nand I_48974 (I835280,I835263,I835246);
nor I_48975 (I835135,I835238,I835280);
DFFARX1 I_48976 (I835280,I2683,I835164,I835320,);
not I_48977 (I835156,I835320);
not I_48978 (I835342,I255405);
nand I_48979 (I835359,I835263,I835342);
DFFARX1 I_48980 (I835359,I2683,I835164,I835385,);
not I_48981 (I835393,I835385);
not I_48982 (I835410,I255396);
nand I_48983 (I835427,I835410,I255384);
and I_48984 (I835444,I835246,I835427);
nor I_48985 (I835461,I835359,I835444);
DFFARX1 I_48986 (I835461,I2683,I835164,I835132,);
DFFARX1 I_48987 (I835444,I2683,I835164,I835153,);
nor I_48988 (I835506,I255396,I255390);
nor I_48989 (I835144,I835359,I835506);
or I_48990 (I835537,I255396,I255390);
nor I_48991 (I835554,I255387,I255381);
DFFARX1 I_48992 (I835554,I2683,I835164,I835580,);
not I_48993 (I835588,I835580);
nor I_48994 (I835150,I835588,I835393);
nand I_48995 (I835619,I835588,I835238);
not I_48996 (I835636,I255387);
nand I_48997 (I835653,I835636,I835342);
nand I_48998 (I835670,I835588,I835653);
nand I_48999 (I835141,I835670,I835619);
nand I_49000 (I835138,I835653,I835537);
not I_49001 (I835742,I2690);
DFFARX1 I_49002 (I985875,I2683,I835742,I835768,);
and I_49003 (I835776,I835768,I985869);
DFFARX1 I_49004 (I835776,I2683,I835742,I835725,);
DFFARX1 I_49005 (I985854,I2683,I835742,I835816,);
not I_49006 (I835824,I985860);
not I_49007 (I835841,I985872);
nand I_49008 (I835858,I835841,I835824);
nor I_49009 (I835713,I835816,I835858);
DFFARX1 I_49010 (I835858,I2683,I835742,I835898,);
not I_49011 (I835734,I835898);
not I_49012 (I835920,I985854);
nand I_49013 (I835937,I835841,I835920);
DFFARX1 I_49014 (I835937,I2683,I835742,I835963,);
not I_49015 (I835971,I835963);
not I_49016 (I835988,I985878);
nand I_49017 (I836005,I835988,I985866);
and I_49018 (I836022,I835824,I836005);
nor I_49019 (I836039,I835937,I836022);
DFFARX1 I_49020 (I836039,I2683,I835742,I835710,);
DFFARX1 I_49021 (I836022,I2683,I835742,I835731,);
nor I_49022 (I836084,I985878,I985857);
nor I_49023 (I835722,I835937,I836084);
or I_49024 (I836115,I985878,I985857);
nor I_49025 (I836132,I985863,I985857);
DFFARX1 I_49026 (I836132,I2683,I835742,I836158,);
not I_49027 (I836166,I836158);
nor I_49028 (I835728,I836166,I835971);
nand I_49029 (I836197,I836166,I835816);
not I_49030 (I836214,I985863);
nand I_49031 (I836231,I836214,I835920);
nand I_49032 (I836248,I836166,I836231);
nand I_49033 (I835719,I836248,I836197);
nand I_49034 (I835716,I836231,I836115);
not I_49035 (I836320,I2690);
DFFARX1 I_49036 (I332850,I2683,I836320,I836346,);
and I_49037 (I836354,I836346,I332865);
DFFARX1 I_49038 (I836354,I2683,I836320,I836303,);
DFFARX1 I_49039 (I332868,I2683,I836320,I836394,);
not I_49040 (I836402,I332862);
not I_49041 (I836419,I332877);
nand I_49042 (I836436,I836419,I836402);
nor I_49043 (I836291,I836394,I836436);
DFFARX1 I_49044 (I836436,I2683,I836320,I836476,);
not I_49045 (I836312,I836476);
not I_49046 (I836498,I332853);
nand I_49047 (I836515,I836419,I836498);
DFFARX1 I_49048 (I836515,I2683,I836320,I836541,);
not I_49049 (I836549,I836541);
not I_49050 (I836566,I332856);
nand I_49051 (I836583,I836566,I332850);
and I_49052 (I836600,I836402,I836583);
nor I_49053 (I836617,I836515,I836600);
DFFARX1 I_49054 (I836617,I2683,I836320,I836288,);
DFFARX1 I_49055 (I836600,I2683,I836320,I836309,);
nor I_49056 (I836662,I332856,I332859);
nor I_49057 (I836300,I836515,I836662);
or I_49058 (I836693,I332856,I332859);
nor I_49059 (I836710,I332874,I332871);
DFFARX1 I_49060 (I836710,I2683,I836320,I836736,);
not I_49061 (I836744,I836736);
nor I_49062 (I836306,I836744,I836549);
nand I_49063 (I836775,I836744,I836394);
not I_49064 (I836792,I332874);
nand I_49065 (I836809,I836792,I836498);
nand I_49066 (I836826,I836744,I836809);
nand I_49067 (I836297,I836826,I836775);
nand I_49068 (I836294,I836809,I836693);
not I_49069 (I836898,I2690);
DFFARX1 I_49070 (I233274,I2683,I836898,I836924,);
and I_49071 (I836932,I836924,I233259);
DFFARX1 I_49072 (I836932,I2683,I836898,I836881,);
DFFARX1 I_49073 (I233265,I2683,I836898,I836972,);
not I_49074 (I836980,I233247);
not I_49075 (I836997,I233268);
nand I_49076 (I837014,I836997,I836980);
nor I_49077 (I836869,I836972,I837014);
DFFARX1 I_49078 (I837014,I2683,I836898,I837054,);
not I_49079 (I836890,I837054);
not I_49080 (I837076,I233271);
nand I_49081 (I837093,I836997,I837076);
DFFARX1 I_49082 (I837093,I2683,I836898,I837119,);
not I_49083 (I837127,I837119);
not I_49084 (I837144,I233262);
nand I_49085 (I837161,I837144,I233250);
and I_49086 (I837178,I836980,I837161);
nor I_49087 (I837195,I837093,I837178);
DFFARX1 I_49088 (I837195,I2683,I836898,I836866,);
DFFARX1 I_49089 (I837178,I2683,I836898,I836887,);
nor I_49090 (I837240,I233262,I233256);
nor I_49091 (I836878,I837093,I837240);
or I_49092 (I837271,I233262,I233256);
nor I_49093 (I837288,I233253,I233247);
DFFARX1 I_49094 (I837288,I2683,I836898,I837314,);
not I_49095 (I837322,I837314);
nor I_49096 (I836884,I837322,I837127);
nand I_49097 (I837353,I837322,I836972);
not I_49098 (I837370,I233253);
nand I_49099 (I837387,I837370,I837076);
nand I_49100 (I837404,I837322,I837387);
nand I_49101 (I836875,I837404,I837353);
nand I_49102 (I836872,I837387,I837271);
not I_49103 (I837476,I2690);
DFFARX1 I_49104 (I517961,I2683,I837476,I837502,);
and I_49105 (I837510,I837502,I517949);
DFFARX1 I_49106 (I837510,I2683,I837476,I837459,);
DFFARX1 I_49107 (I517952,I2683,I837476,I837550,);
not I_49108 (I837558,I517946);
not I_49109 (I837575,I517970);
nand I_49110 (I837592,I837575,I837558);
nor I_49111 (I837447,I837550,I837592);
DFFARX1 I_49112 (I837592,I2683,I837476,I837632,);
not I_49113 (I837468,I837632);
not I_49114 (I837654,I517958);
nand I_49115 (I837671,I837575,I837654);
DFFARX1 I_49116 (I837671,I2683,I837476,I837697,);
not I_49117 (I837705,I837697);
not I_49118 (I837722,I517967);
nand I_49119 (I837739,I837722,I517964);
and I_49120 (I837756,I837558,I837739);
nor I_49121 (I837773,I837671,I837756);
DFFARX1 I_49122 (I837773,I2683,I837476,I837444,);
DFFARX1 I_49123 (I837756,I2683,I837476,I837465,);
nor I_49124 (I837818,I517967,I517955);
nor I_49125 (I837456,I837671,I837818);
or I_49126 (I837849,I517967,I517955);
nor I_49127 (I837866,I517946,I517949);
DFFARX1 I_49128 (I837866,I2683,I837476,I837892,);
not I_49129 (I837900,I837892);
nor I_49130 (I837462,I837900,I837705);
nand I_49131 (I837931,I837900,I837550);
not I_49132 (I837948,I517946);
nand I_49133 (I837965,I837948,I837654);
nand I_49134 (I837982,I837900,I837965);
nand I_49135 (I837453,I837982,I837931);
nand I_49136 (I837450,I837965,I837849);
not I_49137 (I838054,I2690);
DFFARX1 I_49138 (I569981,I2683,I838054,I838080,);
and I_49139 (I838088,I838080,I569969);
DFFARX1 I_49140 (I838088,I2683,I838054,I838037,);
DFFARX1 I_49141 (I569972,I2683,I838054,I838128,);
not I_49142 (I838136,I569966);
not I_49143 (I838153,I569990);
nand I_49144 (I838170,I838153,I838136);
nor I_49145 (I838025,I838128,I838170);
DFFARX1 I_49146 (I838170,I2683,I838054,I838210,);
not I_49147 (I838046,I838210);
not I_49148 (I838232,I569978);
nand I_49149 (I838249,I838153,I838232);
DFFARX1 I_49150 (I838249,I2683,I838054,I838275,);
not I_49151 (I838283,I838275);
not I_49152 (I838300,I569987);
nand I_49153 (I838317,I838300,I569984);
and I_49154 (I838334,I838136,I838317);
nor I_49155 (I838351,I838249,I838334);
DFFARX1 I_49156 (I838351,I2683,I838054,I838022,);
DFFARX1 I_49157 (I838334,I2683,I838054,I838043,);
nor I_49158 (I838396,I569987,I569975);
nor I_49159 (I838034,I838249,I838396);
or I_49160 (I838427,I569987,I569975);
nor I_49161 (I838444,I569966,I569969);
DFFARX1 I_49162 (I838444,I2683,I838054,I838470,);
not I_49163 (I838478,I838470);
nor I_49164 (I838040,I838478,I838283);
nand I_49165 (I838509,I838478,I838128);
not I_49166 (I838526,I569966);
nand I_49167 (I838543,I838526,I838232);
nand I_49168 (I838560,I838478,I838543);
nand I_49169 (I838031,I838560,I838509);
nand I_49170 (I838028,I838543,I838427);
not I_49171 (I838632,I2690);
DFFARX1 I_49172 (I651773,I2683,I838632,I838658,);
and I_49173 (I838666,I838658,I651779);
DFFARX1 I_49174 (I838666,I2683,I838632,I838615,);
DFFARX1 I_49175 (I651785,I2683,I838632,I838706,);
not I_49176 (I838714,I651770);
not I_49177 (I838731,I651770);
nand I_49178 (I838748,I838731,I838714);
nor I_49179 (I838603,I838706,I838748);
DFFARX1 I_49180 (I838748,I2683,I838632,I838788,);
not I_49181 (I838624,I838788);
not I_49182 (I838810,I651788);
nand I_49183 (I838827,I838731,I838810);
DFFARX1 I_49184 (I838827,I2683,I838632,I838853,);
not I_49185 (I838861,I838853);
not I_49186 (I838878,I651782);
nand I_49187 (I838895,I838878,I651773);
and I_49188 (I838912,I838714,I838895);
nor I_49189 (I838929,I838827,I838912);
DFFARX1 I_49190 (I838929,I2683,I838632,I838600,);
DFFARX1 I_49191 (I838912,I2683,I838632,I838621,);
nor I_49192 (I838974,I651782,I651791);
nor I_49193 (I838612,I838827,I838974);
or I_49194 (I839005,I651782,I651791);
nor I_49195 (I839022,I651776,I651776);
DFFARX1 I_49196 (I839022,I2683,I838632,I839048,);
not I_49197 (I839056,I839048);
nor I_49198 (I838618,I839056,I838861);
nand I_49199 (I839087,I839056,I838706);
not I_49200 (I839104,I651776);
nand I_49201 (I839121,I839104,I838810);
nand I_49202 (I839138,I839056,I839121);
nand I_49203 (I838609,I839138,I839087);
nand I_49204 (I838606,I839121,I839005);
not I_49205 (I839210,I2690);
DFFARX1 I_49206 (I709015,I2683,I839210,I839236,);
and I_49207 (I839244,I839236,I709009);
DFFARX1 I_49208 (I839244,I2683,I839210,I839193,);
DFFARX1 I_49209 (I709027,I2683,I839210,I839284,);
not I_49210 (I839292,I709018);
not I_49211 (I839309,I709030);
nand I_49212 (I839326,I839309,I839292);
nor I_49213 (I839181,I839284,I839326);
DFFARX1 I_49214 (I839326,I2683,I839210,I839366,);
not I_49215 (I839202,I839366);
not I_49216 (I839388,I709036);
nand I_49217 (I839405,I839309,I839388);
DFFARX1 I_49218 (I839405,I2683,I839210,I839431,);
not I_49219 (I839439,I839431);
not I_49220 (I839456,I709012);
nand I_49221 (I839473,I839456,I709033);
and I_49222 (I839490,I839292,I839473);
nor I_49223 (I839507,I839405,I839490);
DFFARX1 I_49224 (I839507,I2683,I839210,I839178,);
DFFARX1 I_49225 (I839490,I2683,I839210,I839199,);
nor I_49226 (I839552,I709012,I709024);
nor I_49227 (I839190,I839405,I839552);
or I_49228 (I839583,I709012,I709024);
nor I_49229 (I839600,I709009,I709021);
DFFARX1 I_49230 (I839600,I2683,I839210,I839626,);
not I_49231 (I839634,I839626);
nor I_49232 (I839196,I839634,I839439);
nand I_49233 (I839665,I839634,I839284);
not I_49234 (I839682,I709009);
nand I_49235 (I839699,I839682,I839388);
nand I_49236 (I839716,I839634,I839699);
nand I_49237 (I839187,I839716,I839665);
nand I_49238 (I839184,I839699,I839583);
not I_49239 (I839788,I2690);
DFFARX1 I_49240 (I774261,I2683,I839788,I839814,);
and I_49241 (I839822,I839814,I774255);
DFFARX1 I_49242 (I839822,I2683,I839788,I839771,);
DFFARX1 I_49243 (I774273,I2683,I839788,I839862,);
not I_49244 (I839870,I774264);
not I_49245 (I839887,I774276);
nand I_49246 (I839904,I839887,I839870);
nor I_49247 (I839759,I839862,I839904);
DFFARX1 I_49248 (I839904,I2683,I839788,I839944,);
not I_49249 (I839780,I839944);
not I_49250 (I839966,I774282);
nand I_49251 (I839983,I839887,I839966);
DFFARX1 I_49252 (I839983,I2683,I839788,I840009,);
not I_49253 (I840017,I840009);
not I_49254 (I840034,I774258);
nand I_49255 (I840051,I840034,I774279);
and I_49256 (I840068,I839870,I840051);
nor I_49257 (I840085,I839983,I840068);
DFFARX1 I_49258 (I840085,I2683,I839788,I839756,);
DFFARX1 I_49259 (I840068,I2683,I839788,I839777,);
nor I_49260 (I840130,I774258,I774270);
nor I_49261 (I839768,I839983,I840130);
or I_49262 (I840161,I774258,I774270);
nor I_49263 (I840178,I774255,I774267);
DFFARX1 I_49264 (I840178,I2683,I839788,I840204,);
not I_49265 (I840212,I840204);
nor I_49266 (I839774,I840212,I840017);
nand I_49267 (I840243,I840212,I839862);
not I_49268 (I840260,I774255);
nand I_49269 (I840277,I840260,I839966);
nand I_49270 (I840294,I840212,I840277);
nand I_49271 (I839765,I840294,I840243);
nand I_49272 (I839762,I840277,I840161);
not I_49273 (I840366,I2690);
DFFARX1 I_49274 (I805759,I2683,I840366,I840392,);
and I_49275 (I840400,I840392,I805756);
DFFARX1 I_49276 (I840400,I2683,I840366,I840349,);
DFFARX1 I_49277 (I805762,I2683,I840366,I840440,);
not I_49278 (I840448,I805765);
not I_49279 (I840465,I805759);
nand I_49280 (I840482,I840465,I840448);
nor I_49281 (I840337,I840440,I840482);
DFFARX1 I_49282 (I840482,I2683,I840366,I840522,);
not I_49283 (I840358,I840522);
not I_49284 (I840544,I805774);
nand I_49285 (I840561,I840465,I840544);
DFFARX1 I_49286 (I840561,I2683,I840366,I840587,);
not I_49287 (I840595,I840587);
not I_49288 (I840612,I805771);
nand I_49289 (I840629,I840612,I805777);
and I_49290 (I840646,I840448,I840629);
nor I_49291 (I840663,I840561,I840646);
DFFARX1 I_49292 (I840663,I2683,I840366,I840334,);
DFFARX1 I_49293 (I840646,I2683,I840366,I840355,);
nor I_49294 (I840708,I805771,I805756);
nor I_49295 (I840346,I840561,I840708);
or I_49296 (I840739,I805771,I805756);
nor I_49297 (I840756,I805768,I805762);
DFFARX1 I_49298 (I840756,I2683,I840366,I840782,);
not I_49299 (I840790,I840782);
nor I_49300 (I840352,I840790,I840595);
nand I_49301 (I840821,I840790,I840440);
not I_49302 (I840838,I805768);
nand I_49303 (I840855,I840838,I840544);
nand I_49304 (I840872,I840790,I840855);
nand I_49305 (I840343,I840872,I840821);
nand I_49306 (I840340,I840855,I840739);
not I_49307 (I840944,I2690);
DFFARX1 I_49308 (I196170,I2683,I840944,I840970,);
and I_49309 (I840978,I840970,I196173);
DFFARX1 I_49310 (I840978,I2683,I840944,I840927,);
DFFARX1 I_49311 (I196173,I2683,I840944,I841018,);
not I_49312 (I841026,I196188);
not I_49313 (I841043,I196194);
nand I_49314 (I841060,I841043,I841026);
nor I_49315 (I840915,I841018,I841060);
DFFARX1 I_49316 (I841060,I2683,I840944,I841100,);
not I_49317 (I840936,I841100);
not I_49318 (I841122,I196182);
nand I_49319 (I841139,I841043,I841122);
DFFARX1 I_49320 (I841139,I2683,I840944,I841165,);
not I_49321 (I841173,I841165);
not I_49322 (I841190,I196179);
nand I_49323 (I841207,I841190,I196176);
and I_49324 (I841224,I841026,I841207);
nor I_49325 (I841241,I841139,I841224);
DFFARX1 I_49326 (I841241,I2683,I840944,I840912,);
DFFARX1 I_49327 (I841224,I2683,I840944,I840933,);
nor I_49328 (I841286,I196179,I196170);
nor I_49329 (I840924,I841139,I841286);
or I_49330 (I841317,I196179,I196170);
nor I_49331 (I841334,I196185,I196191);
DFFARX1 I_49332 (I841334,I2683,I840944,I841360,);
not I_49333 (I841368,I841360);
nor I_49334 (I840930,I841368,I841173);
nand I_49335 (I841399,I841368,I841018);
not I_49336 (I841416,I196185);
nand I_49337 (I841433,I841416,I841122);
nand I_49338 (I841450,I841368,I841433);
nand I_49339 (I840921,I841450,I841399);
nand I_49340 (I840918,I841433,I841317);
not I_49341 (I841522,I2690);
DFFARX1 I_49342 (I275961,I2683,I841522,I841548,);
and I_49343 (I841556,I841548,I275946);
DFFARX1 I_49344 (I841556,I2683,I841522,I841505,);
DFFARX1 I_49345 (I275952,I2683,I841522,I841596,);
not I_49346 (I841604,I275934);
not I_49347 (I841621,I275955);
nand I_49348 (I841638,I841621,I841604);
nor I_49349 (I841493,I841596,I841638);
DFFARX1 I_49350 (I841638,I2683,I841522,I841678,);
not I_49351 (I841514,I841678);
not I_49352 (I841700,I275958);
nand I_49353 (I841717,I841621,I841700);
DFFARX1 I_49354 (I841717,I2683,I841522,I841743,);
not I_49355 (I841751,I841743);
not I_49356 (I841768,I275949);
nand I_49357 (I841785,I841768,I275937);
and I_49358 (I841802,I841604,I841785);
nor I_49359 (I841819,I841717,I841802);
DFFARX1 I_49360 (I841819,I2683,I841522,I841490,);
DFFARX1 I_49361 (I841802,I2683,I841522,I841511,);
nor I_49362 (I841864,I275949,I275943);
nor I_49363 (I841502,I841717,I841864);
or I_49364 (I841895,I275949,I275943);
nor I_49365 (I841912,I275940,I275934);
DFFARX1 I_49366 (I841912,I2683,I841522,I841938,);
not I_49367 (I841946,I841938);
nor I_49368 (I841508,I841946,I841751);
nand I_49369 (I841977,I841946,I841596);
not I_49370 (I841994,I275940);
nand I_49371 (I842011,I841994,I841700);
nand I_49372 (I842028,I841946,I842011);
nand I_49373 (I841499,I842028,I841977);
nand I_49374 (I841496,I842011,I841895);
not I_49375 (I842100,I2690);
DFFARX1 I_49376 (I130125,I2683,I842100,I842126,);
and I_49377 (I842134,I842126,I130128);
DFFARX1 I_49378 (I842134,I2683,I842100,I842083,);
DFFARX1 I_49379 (I130128,I2683,I842100,I842174,);
not I_49380 (I842182,I130143);
not I_49381 (I842199,I130149);
nand I_49382 (I842216,I842199,I842182);
nor I_49383 (I842071,I842174,I842216);
DFFARX1 I_49384 (I842216,I2683,I842100,I842256,);
not I_49385 (I842092,I842256);
not I_49386 (I842278,I130137);
nand I_49387 (I842295,I842199,I842278);
DFFARX1 I_49388 (I842295,I2683,I842100,I842321,);
not I_49389 (I842329,I842321);
not I_49390 (I842346,I130134);
nand I_49391 (I842363,I842346,I130131);
and I_49392 (I842380,I842182,I842363);
nor I_49393 (I842397,I842295,I842380);
DFFARX1 I_49394 (I842397,I2683,I842100,I842068,);
DFFARX1 I_49395 (I842380,I2683,I842100,I842089,);
nor I_49396 (I842442,I130134,I130125);
nor I_49397 (I842080,I842295,I842442);
or I_49398 (I842473,I130134,I130125);
nor I_49399 (I842490,I130140,I130146);
DFFARX1 I_49400 (I842490,I2683,I842100,I842516,);
not I_49401 (I842524,I842516);
nor I_49402 (I842086,I842524,I842329);
nand I_49403 (I842555,I842524,I842174);
not I_49404 (I842572,I130140);
nand I_49405 (I842589,I842572,I842278);
nand I_49406 (I842606,I842524,I842589);
nand I_49407 (I842077,I842606,I842555);
nand I_49408 (I842074,I842589,I842473);
not I_49409 (I842678,I2690);
DFFARX1 I_49410 (I790411,I2683,I842678,I842704,);
and I_49411 (I842712,I842704,I790405);
DFFARX1 I_49412 (I842712,I2683,I842678,I842661,);
DFFARX1 I_49413 (I790423,I2683,I842678,I842752,);
not I_49414 (I842760,I790414);
not I_49415 (I842777,I790426);
nand I_49416 (I842794,I842777,I842760);
nor I_49417 (I842649,I842752,I842794);
DFFARX1 I_49418 (I842794,I2683,I842678,I842834,);
not I_49419 (I842670,I842834);
not I_49420 (I842856,I790432);
nand I_49421 (I842873,I842777,I842856);
DFFARX1 I_49422 (I842873,I2683,I842678,I842899,);
not I_49423 (I842907,I842899);
not I_49424 (I842924,I790408);
nand I_49425 (I842941,I842924,I790429);
and I_49426 (I842958,I842760,I842941);
nor I_49427 (I842975,I842873,I842958);
DFFARX1 I_49428 (I842975,I2683,I842678,I842646,);
DFFARX1 I_49429 (I842958,I2683,I842678,I842667,);
nor I_49430 (I843020,I790408,I790420);
nor I_49431 (I842658,I842873,I843020);
or I_49432 (I843051,I790408,I790420);
nor I_49433 (I843068,I790405,I790417);
DFFARX1 I_49434 (I843068,I2683,I842678,I843094,);
not I_49435 (I843102,I843094);
nor I_49436 (I842664,I843102,I842907);
nand I_49437 (I843133,I843102,I842752);
not I_49438 (I843150,I790405);
nand I_49439 (I843167,I843150,I842856);
nand I_49440 (I843184,I843102,I843167);
nand I_49441 (I842655,I843184,I843133);
nand I_49442 (I842652,I843167,I843051);
not I_49443 (I843256,I2690);
DFFARX1 I_49444 (I443977,I2683,I843256,I843282,);
and I_49445 (I843290,I843282,I443965);
DFFARX1 I_49446 (I843290,I2683,I843256,I843239,);
DFFARX1 I_49447 (I443980,I2683,I843256,I843330,);
not I_49448 (I843338,I443971);
not I_49449 (I843355,I443962);
nand I_49450 (I843372,I843355,I843338);
nor I_49451 (I843227,I843330,I843372);
DFFARX1 I_49452 (I843372,I2683,I843256,I843412,);
not I_49453 (I843248,I843412);
not I_49454 (I843434,I443968);
nand I_49455 (I843451,I843355,I843434);
DFFARX1 I_49456 (I843451,I2683,I843256,I843477,);
not I_49457 (I843485,I843477);
not I_49458 (I843502,I443983);
nand I_49459 (I843519,I843502,I443986);
and I_49460 (I843536,I843338,I843519);
nor I_49461 (I843553,I843451,I843536);
DFFARX1 I_49462 (I843553,I2683,I843256,I843224,);
DFFARX1 I_49463 (I843536,I2683,I843256,I843245,);
nor I_49464 (I843598,I443983,I443962);
nor I_49465 (I843236,I843451,I843598);
or I_49466 (I843629,I443983,I443962);
nor I_49467 (I843646,I443974,I443965);
DFFARX1 I_49468 (I843646,I2683,I843256,I843672,);
not I_49469 (I843680,I843672);
nor I_49470 (I843242,I843680,I843485);
nand I_49471 (I843711,I843680,I843330);
not I_49472 (I843728,I443974);
nand I_49473 (I843745,I843728,I843434);
nand I_49474 (I843762,I843680,I843745);
nand I_49475 (I843233,I843762,I843711);
nand I_49476 (I843230,I843745,I843629);
not I_49477 (I843834,I2690);
DFFARX1 I_49478 (I274907,I2683,I843834,I843860,);
and I_49479 (I843868,I843860,I274892);
DFFARX1 I_49480 (I843868,I2683,I843834,I843817,);
DFFARX1 I_49481 (I274898,I2683,I843834,I843908,);
not I_49482 (I843916,I274880);
not I_49483 (I843933,I274901);
nand I_49484 (I843950,I843933,I843916);
nor I_49485 (I843805,I843908,I843950);
DFFARX1 I_49486 (I843950,I2683,I843834,I843990,);
not I_49487 (I843826,I843990);
not I_49488 (I844012,I274904);
nand I_49489 (I844029,I843933,I844012);
DFFARX1 I_49490 (I844029,I2683,I843834,I844055,);
not I_49491 (I844063,I844055);
not I_49492 (I844080,I274895);
nand I_49493 (I844097,I844080,I274883);
and I_49494 (I844114,I843916,I844097);
nor I_49495 (I844131,I844029,I844114);
DFFARX1 I_49496 (I844131,I2683,I843834,I843802,);
DFFARX1 I_49497 (I844114,I2683,I843834,I843823,);
nor I_49498 (I844176,I274895,I274889);
nor I_49499 (I843814,I844029,I844176);
or I_49500 (I844207,I274895,I274889);
nor I_49501 (I844224,I274886,I274880);
DFFARX1 I_49502 (I844224,I2683,I843834,I844250,);
not I_49503 (I844258,I844250);
nor I_49504 (I843820,I844258,I844063);
nand I_49505 (I844289,I844258,I843908);
not I_49506 (I844306,I274886);
nand I_49507 (I844323,I844306,I844012);
nand I_49508 (I844340,I844258,I844323);
nand I_49509 (I843811,I844340,I844289);
nand I_49510 (I843808,I844323,I844207);
not I_49511 (I844412,I2690);
DFFARX1 I_49512 (I274380,I2683,I844412,I844438,);
and I_49513 (I844446,I844438,I274365);
DFFARX1 I_49514 (I844446,I2683,I844412,I844395,);
DFFARX1 I_49515 (I274371,I2683,I844412,I844486,);
not I_49516 (I844494,I274353);
not I_49517 (I844511,I274374);
nand I_49518 (I844528,I844511,I844494);
nor I_49519 (I844383,I844486,I844528);
DFFARX1 I_49520 (I844528,I2683,I844412,I844568,);
not I_49521 (I844404,I844568);
not I_49522 (I844590,I274377);
nand I_49523 (I844607,I844511,I844590);
DFFARX1 I_49524 (I844607,I2683,I844412,I844633,);
not I_49525 (I844641,I844633);
not I_49526 (I844658,I274368);
nand I_49527 (I844675,I844658,I274356);
and I_49528 (I844692,I844494,I844675);
nor I_49529 (I844709,I844607,I844692);
DFFARX1 I_49530 (I844709,I2683,I844412,I844380,);
DFFARX1 I_49531 (I844692,I2683,I844412,I844401,);
nor I_49532 (I844754,I274368,I274362);
nor I_49533 (I844392,I844607,I844754);
or I_49534 (I844785,I274368,I274362);
nor I_49535 (I844802,I274359,I274353);
DFFARX1 I_49536 (I844802,I2683,I844412,I844828,);
not I_49537 (I844836,I844828);
nor I_49538 (I844398,I844836,I844641);
nand I_49539 (I844867,I844836,I844486);
not I_49540 (I844884,I274359);
nand I_49541 (I844901,I844884,I844590);
nand I_49542 (I844918,I844836,I844901);
nand I_49543 (I844389,I844918,I844867);
nand I_49544 (I844386,I844901,I844785);
not I_49545 (I844990,I2690);
DFFARX1 I_49546 (I552063,I2683,I844990,I845016,);
and I_49547 (I845024,I845016,I552051);
DFFARX1 I_49548 (I845024,I2683,I844990,I844973,);
DFFARX1 I_49549 (I552054,I2683,I844990,I845064,);
not I_49550 (I845072,I552048);
not I_49551 (I845089,I552072);
nand I_49552 (I845106,I845089,I845072);
nor I_49553 (I844961,I845064,I845106);
DFFARX1 I_49554 (I845106,I2683,I844990,I845146,);
not I_49555 (I844982,I845146);
not I_49556 (I845168,I552060);
nand I_49557 (I845185,I845089,I845168);
DFFARX1 I_49558 (I845185,I2683,I844990,I845211,);
not I_49559 (I845219,I845211);
not I_49560 (I845236,I552069);
nand I_49561 (I845253,I845236,I552066);
and I_49562 (I845270,I845072,I845253);
nor I_49563 (I845287,I845185,I845270);
DFFARX1 I_49564 (I845287,I2683,I844990,I844958,);
DFFARX1 I_49565 (I845270,I2683,I844990,I844979,);
nor I_49566 (I845332,I552069,I552057);
nor I_49567 (I844970,I845185,I845332);
or I_49568 (I845363,I552069,I552057);
nor I_49569 (I845380,I552048,I552051);
DFFARX1 I_49570 (I845380,I2683,I844990,I845406,);
not I_49571 (I845414,I845406);
nor I_49572 (I844976,I845414,I845219);
nand I_49573 (I845445,I845414,I845064);
not I_49574 (I845462,I552048);
nand I_49575 (I845479,I845462,I845168);
nand I_49576 (I845496,I845414,I845479);
nand I_49577 (I844967,I845496,I845445);
nand I_49578 (I844964,I845479,I845363);
not I_49579 (I845568,I2690);
DFFARX1 I_49580 (I685501,I2683,I845568,I845594,);
and I_49581 (I845602,I845594,I685507);
DFFARX1 I_49582 (I845602,I2683,I845568,I845551,);
DFFARX1 I_49583 (I685513,I2683,I845568,I845642,);
not I_49584 (I845650,I685498);
not I_49585 (I845667,I685498);
nand I_49586 (I845684,I845667,I845650);
nor I_49587 (I845539,I845642,I845684);
DFFARX1 I_49588 (I845684,I2683,I845568,I845724,);
not I_49589 (I845560,I845724);
not I_49590 (I845746,I685516);
nand I_49591 (I845763,I845667,I845746);
DFFARX1 I_49592 (I845763,I2683,I845568,I845789,);
not I_49593 (I845797,I845789);
not I_49594 (I845814,I685510);
nand I_49595 (I845831,I845814,I685501);
and I_49596 (I845848,I845650,I845831);
nor I_49597 (I845865,I845763,I845848);
DFFARX1 I_49598 (I845865,I2683,I845568,I845536,);
DFFARX1 I_49599 (I845848,I2683,I845568,I845557,);
nor I_49600 (I845910,I685510,I685519);
nor I_49601 (I845548,I845763,I845910);
or I_49602 (I845941,I685510,I685519);
nor I_49603 (I845958,I685504,I685504);
DFFARX1 I_49604 (I845958,I2683,I845568,I845984,);
not I_49605 (I845992,I845984);
nor I_49606 (I845554,I845992,I845797);
nand I_49607 (I846023,I845992,I845642);
not I_49608 (I846040,I685504);
nand I_49609 (I846057,I846040,I845746);
nand I_49610 (I846074,I845992,I846057);
nand I_49611 (I845545,I846074,I846023);
nand I_49612 (I845542,I846057,I845941);
not I_49613 (I846146,I2690);
DFFARX1 I_49614 (I434729,I2683,I846146,I846172,);
and I_49615 (I846180,I846172,I434717);
DFFARX1 I_49616 (I846180,I2683,I846146,I846129,);
DFFARX1 I_49617 (I434732,I2683,I846146,I846220,);
not I_49618 (I846228,I434723);
not I_49619 (I846245,I434714);
nand I_49620 (I846262,I846245,I846228);
nor I_49621 (I846117,I846220,I846262);
DFFARX1 I_49622 (I846262,I2683,I846146,I846302,);
not I_49623 (I846138,I846302);
not I_49624 (I846324,I434720);
nand I_49625 (I846341,I846245,I846324);
DFFARX1 I_49626 (I846341,I2683,I846146,I846367,);
not I_49627 (I846375,I846367);
not I_49628 (I846392,I434735);
nand I_49629 (I846409,I846392,I434738);
and I_49630 (I846426,I846228,I846409);
nor I_49631 (I846443,I846341,I846426);
DFFARX1 I_49632 (I846443,I2683,I846146,I846114,);
DFFARX1 I_49633 (I846426,I2683,I846146,I846135,);
nor I_49634 (I846488,I434735,I434714);
nor I_49635 (I846126,I846341,I846488);
or I_49636 (I846519,I434735,I434714);
nor I_49637 (I846536,I434726,I434717);
DFFARX1 I_49638 (I846536,I2683,I846146,I846562,);
not I_49639 (I846570,I846562);
nor I_49640 (I846132,I846570,I846375);
nand I_49641 (I846601,I846570,I846220);
not I_49642 (I846618,I434726);
nand I_49643 (I846635,I846618,I846324);
nand I_49644 (I846652,I846570,I846635);
nand I_49645 (I846123,I846652,I846601);
nand I_49646 (I846120,I846635,I846519);
not I_49647 (I846724,I2690);
DFFARX1 I_49648 (I386162,I2683,I846724,I846750,);
and I_49649 (I846758,I846750,I386177);
DFFARX1 I_49650 (I846758,I2683,I846724,I846707,);
DFFARX1 I_49651 (I386180,I2683,I846724,I846798,);
not I_49652 (I846806,I386174);
not I_49653 (I846823,I386189);
nand I_49654 (I846840,I846823,I846806);
nor I_49655 (I846695,I846798,I846840);
DFFARX1 I_49656 (I846840,I2683,I846724,I846880,);
not I_49657 (I846716,I846880);
not I_49658 (I846902,I386165);
nand I_49659 (I846919,I846823,I846902);
DFFARX1 I_49660 (I846919,I2683,I846724,I846945,);
not I_49661 (I846953,I846945);
not I_49662 (I846970,I386168);
nand I_49663 (I846987,I846970,I386162);
and I_49664 (I847004,I846806,I846987);
nor I_49665 (I847021,I846919,I847004);
DFFARX1 I_49666 (I847021,I2683,I846724,I846692,);
DFFARX1 I_49667 (I847004,I2683,I846724,I846713,);
nor I_49668 (I847066,I386168,I386171);
nor I_49669 (I846704,I846919,I847066);
or I_49670 (I847097,I386168,I386171);
nor I_49671 (I847114,I386186,I386183);
DFFARX1 I_49672 (I847114,I2683,I846724,I847140,);
not I_49673 (I847148,I847140);
nor I_49674 (I846710,I847148,I846953);
nand I_49675 (I847179,I847148,I846798);
not I_49676 (I847196,I386186);
nand I_49677 (I847213,I847196,I846902);
nand I_49678 (I847230,I847148,I847213);
nand I_49679 (I846701,I847230,I847179);
nand I_49680 (I846698,I847213,I847097);
not I_49681 (I847302,I2690);
DFFARX1 I_49682 (I380178,I2683,I847302,I847328,);
and I_49683 (I847336,I847328,I380193);
DFFARX1 I_49684 (I847336,I2683,I847302,I847285,);
DFFARX1 I_49685 (I380196,I2683,I847302,I847376,);
not I_49686 (I847384,I380190);
not I_49687 (I847401,I380205);
nand I_49688 (I847418,I847401,I847384);
nor I_49689 (I847273,I847376,I847418);
DFFARX1 I_49690 (I847418,I2683,I847302,I847458,);
not I_49691 (I847294,I847458);
not I_49692 (I847480,I380181);
nand I_49693 (I847497,I847401,I847480);
DFFARX1 I_49694 (I847497,I2683,I847302,I847523,);
not I_49695 (I847531,I847523);
not I_49696 (I847548,I380184);
nand I_49697 (I847565,I847548,I380178);
and I_49698 (I847582,I847384,I847565);
nor I_49699 (I847599,I847497,I847582);
DFFARX1 I_49700 (I847599,I2683,I847302,I847270,);
DFFARX1 I_49701 (I847582,I2683,I847302,I847291,);
nor I_49702 (I847644,I380184,I380187);
nor I_49703 (I847282,I847497,I847644);
or I_49704 (I847675,I380184,I380187);
nor I_49705 (I847692,I380202,I380199);
DFFARX1 I_49706 (I847692,I2683,I847302,I847718,);
not I_49707 (I847726,I847718);
nor I_49708 (I847288,I847726,I847531);
nand I_49709 (I847757,I847726,I847376);
not I_49710 (I847774,I380202);
nand I_49711 (I847791,I847774,I847480);
nand I_49712 (I847808,I847726,I847791);
nand I_49713 (I847279,I847808,I847757);
nand I_49714 (I847276,I847791,I847675);
not I_49715 (I847880,I2690);
DFFARX1 I_49716 (I308108,I2683,I847880,I847906,);
and I_49717 (I847914,I847906,I308093);
DFFARX1 I_49718 (I847914,I2683,I847880,I847863,);
DFFARX1 I_49719 (I308099,I2683,I847880,I847954,);
not I_49720 (I847962,I308081);
not I_49721 (I847979,I308102);
nand I_49722 (I847996,I847979,I847962);
nor I_49723 (I847851,I847954,I847996);
DFFARX1 I_49724 (I847996,I2683,I847880,I848036,);
not I_49725 (I847872,I848036);
not I_49726 (I848058,I308105);
nand I_49727 (I848075,I847979,I848058);
DFFARX1 I_49728 (I848075,I2683,I847880,I848101,);
not I_49729 (I848109,I848101);
not I_49730 (I848126,I308096);
nand I_49731 (I848143,I848126,I308084);
and I_49732 (I848160,I847962,I848143);
nor I_49733 (I848177,I848075,I848160);
DFFARX1 I_49734 (I848177,I2683,I847880,I847848,);
DFFARX1 I_49735 (I848160,I2683,I847880,I847869,);
nor I_49736 (I848222,I308096,I308090);
nor I_49737 (I847860,I848075,I848222);
or I_49738 (I848253,I308096,I308090);
nor I_49739 (I848270,I308087,I308081);
DFFARX1 I_49740 (I848270,I2683,I847880,I848296,);
not I_49741 (I848304,I848296);
nor I_49742 (I847866,I848304,I848109);
nand I_49743 (I848335,I848304,I847954);
not I_49744 (I848352,I308087);
nand I_49745 (I848369,I848352,I848058);
nand I_49746 (I848386,I848304,I848369);
nand I_49747 (I847857,I848386,I848335);
nand I_49748 (I847854,I848369,I848253);
not I_49749 (I848458,I2690);
DFFARX1 I_49750 (I1062041,I2683,I848458,I848484,);
and I_49751 (I848492,I848484,I1062023);
DFFARX1 I_49752 (I848492,I2683,I848458,I848441,);
DFFARX1 I_49753 (I1062014,I2683,I848458,I848532,);
not I_49754 (I848540,I1062029);
not I_49755 (I848557,I1062017);
nand I_49756 (I848574,I848557,I848540);
nor I_49757 (I848429,I848532,I848574);
DFFARX1 I_49758 (I848574,I2683,I848458,I848614,);
not I_49759 (I848450,I848614);
not I_49760 (I848636,I1062026);
nand I_49761 (I848653,I848557,I848636);
DFFARX1 I_49762 (I848653,I2683,I848458,I848679,);
not I_49763 (I848687,I848679);
not I_49764 (I848704,I1062035);
nand I_49765 (I848721,I848704,I1062014);
and I_49766 (I848738,I848540,I848721);
nor I_49767 (I848755,I848653,I848738);
DFFARX1 I_49768 (I848755,I2683,I848458,I848426,);
DFFARX1 I_49769 (I848738,I2683,I848458,I848447,);
nor I_49770 (I848800,I1062035,I1062038);
nor I_49771 (I848438,I848653,I848800);
or I_49772 (I848831,I1062035,I1062038);
nor I_49773 (I848848,I1062032,I1062020);
DFFARX1 I_49774 (I848848,I2683,I848458,I848874,);
not I_49775 (I848882,I848874);
nor I_49776 (I848444,I848882,I848687);
nand I_49777 (I848913,I848882,I848532);
not I_49778 (I848930,I1062032);
nand I_49779 (I848947,I848930,I848636);
nand I_49780 (I848964,I848882,I848947);
nand I_49781 (I848435,I848964,I848913);
nand I_49782 (I848432,I848947,I848831);
not I_49783 (I849036,I2690);
DFFARX1 I_49784 (I970643,I2683,I849036,I849062,);
and I_49785 (I849070,I849062,I970637);
DFFARX1 I_49786 (I849070,I2683,I849036,I849019,);
DFFARX1 I_49787 (I970622,I2683,I849036,I849110,);
not I_49788 (I849118,I970628);
not I_49789 (I849135,I970640);
nand I_49790 (I849152,I849135,I849118);
nor I_49791 (I849007,I849110,I849152);
DFFARX1 I_49792 (I849152,I2683,I849036,I849192,);
not I_49793 (I849028,I849192);
not I_49794 (I849214,I970622);
nand I_49795 (I849231,I849135,I849214);
DFFARX1 I_49796 (I849231,I2683,I849036,I849257,);
not I_49797 (I849265,I849257);
not I_49798 (I849282,I970646);
nand I_49799 (I849299,I849282,I970634);
and I_49800 (I849316,I849118,I849299);
nor I_49801 (I849333,I849231,I849316);
DFFARX1 I_49802 (I849333,I2683,I849036,I849004,);
DFFARX1 I_49803 (I849316,I2683,I849036,I849025,);
nor I_49804 (I849378,I970646,I970625);
nor I_49805 (I849016,I849231,I849378);
or I_49806 (I849409,I970646,I970625);
nor I_49807 (I849426,I970631,I970625);
DFFARX1 I_49808 (I849426,I2683,I849036,I849452,);
not I_49809 (I849460,I849452);
nor I_49810 (I849022,I849460,I849265);
nand I_49811 (I849491,I849460,I849110);
not I_49812 (I849508,I970631);
nand I_49813 (I849525,I849508,I849214);
nand I_49814 (I849542,I849460,I849525);
nand I_49815 (I849013,I849542,I849491);
nand I_49816 (I849010,I849525,I849409);
not I_49817 (I849614,I2690);
DFFARX1 I_49818 (I976627,I2683,I849614,I849640,);
and I_49819 (I849648,I849640,I976621);
DFFARX1 I_49820 (I849648,I2683,I849614,I849597,);
DFFARX1 I_49821 (I976606,I2683,I849614,I849688,);
not I_49822 (I849696,I976612);
not I_49823 (I849713,I976624);
nand I_49824 (I849730,I849713,I849696);
nor I_49825 (I849585,I849688,I849730);
DFFARX1 I_49826 (I849730,I2683,I849614,I849770,);
not I_49827 (I849606,I849770);
not I_49828 (I849792,I976606);
nand I_49829 (I849809,I849713,I849792);
DFFARX1 I_49830 (I849809,I2683,I849614,I849835,);
not I_49831 (I849843,I849835);
not I_49832 (I849860,I976630);
nand I_49833 (I849877,I849860,I976618);
and I_49834 (I849894,I849696,I849877);
nor I_49835 (I849911,I849809,I849894);
DFFARX1 I_49836 (I849911,I2683,I849614,I849582,);
DFFARX1 I_49837 (I849894,I2683,I849614,I849603,);
nor I_49838 (I849956,I976630,I976609);
nor I_49839 (I849594,I849809,I849956);
or I_49840 (I849987,I976630,I976609);
nor I_49841 (I850004,I976615,I976609);
DFFARX1 I_49842 (I850004,I2683,I849614,I850030,);
not I_49843 (I850038,I850030);
nor I_49844 (I849600,I850038,I849843);
nand I_49845 (I850069,I850038,I849688);
not I_49846 (I850086,I976615);
nand I_49847 (I850103,I850086,I849792);
nand I_49848 (I850120,I850038,I850103);
nand I_49849 (I849591,I850120,I850069);
nand I_49850 (I849588,I850103,I849987);
not I_49851 (I850192,I2690);
DFFARX1 I_49852 (I142025,I2683,I850192,I850218,);
and I_49853 (I850226,I850218,I142028);
DFFARX1 I_49854 (I850226,I2683,I850192,I850175,);
DFFARX1 I_49855 (I142028,I2683,I850192,I850266,);
not I_49856 (I850274,I142043);
not I_49857 (I850291,I142049);
nand I_49858 (I850308,I850291,I850274);
nor I_49859 (I850163,I850266,I850308);
DFFARX1 I_49860 (I850308,I2683,I850192,I850348,);
not I_49861 (I850184,I850348);
not I_49862 (I850370,I142037);
nand I_49863 (I850387,I850291,I850370);
DFFARX1 I_49864 (I850387,I2683,I850192,I850413,);
not I_49865 (I850421,I850413);
not I_49866 (I850438,I142034);
nand I_49867 (I850455,I850438,I142031);
and I_49868 (I850472,I850274,I850455);
nor I_49869 (I850489,I850387,I850472);
DFFARX1 I_49870 (I850489,I2683,I850192,I850160,);
DFFARX1 I_49871 (I850472,I2683,I850192,I850181,);
nor I_49872 (I850534,I142034,I142025);
nor I_49873 (I850172,I850387,I850534);
or I_49874 (I850565,I142034,I142025);
nor I_49875 (I850582,I142040,I142046);
DFFARX1 I_49876 (I850582,I2683,I850192,I850608,);
not I_49877 (I850616,I850608);
nor I_49878 (I850178,I850616,I850421);
nand I_49879 (I850647,I850616,I850266);
not I_49880 (I850664,I142040);
nand I_49881 (I850681,I850664,I850370);
nand I_49882 (I850698,I850616,I850681);
nand I_49883 (I850169,I850698,I850647);
nand I_49884 (I850166,I850681,I850565);
not I_49885 (I850770,I2690);
DFFARX1 I_49886 (I271745,I2683,I850770,I850796,);
and I_49887 (I850804,I850796,I271730);
DFFARX1 I_49888 (I850804,I2683,I850770,I850753,);
DFFARX1 I_49889 (I271736,I2683,I850770,I850844,);
not I_49890 (I850852,I271718);
not I_49891 (I850869,I271739);
nand I_49892 (I850886,I850869,I850852);
nor I_49893 (I850741,I850844,I850886);
DFFARX1 I_49894 (I850886,I2683,I850770,I850926,);
not I_49895 (I850762,I850926);
not I_49896 (I850948,I271742);
nand I_49897 (I850965,I850869,I850948);
DFFARX1 I_49898 (I850965,I2683,I850770,I850991,);
not I_49899 (I850999,I850991);
not I_49900 (I851016,I271733);
nand I_49901 (I851033,I851016,I271721);
and I_49902 (I851050,I850852,I851033);
nor I_49903 (I851067,I850965,I851050);
DFFARX1 I_49904 (I851067,I2683,I850770,I850738,);
DFFARX1 I_49905 (I851050,I2683,I850770,I850759,);
nor I_49906 (I851112,I271733,I271727);
nor I_49907 (I850750,I850965,I851112);
or I_49908 (I851143,I271733,I271727);
nor I_49909 (I851160,I271724,I271718);
DFFARX1 I_49910 (I851160,I2683,I850770,I851186,);
not I_49911 (I851194,I851186);
nor I_49912 (I850756,I851194,I850999);
nand I_49913 (I851225,I851194,I850844);
not I_49914 (I851242,I271724);
nand I_49915 (I851259,I851242,I850948);
nand I_49916 (I851276,I851194,I851259);
nand I_49917 (I850747,I851276,I851225);
nand I_49918 (I850744,I851259,I851143);
not I_49919 (I851348,I2690);
DFFARX1 I_49920 (I290190,I2683,I851348,I851374,);
and I_49921 (I851382,I851374,I290175);
DFFARX1 I_49922 (I851382,I2683,I851348,I851331,);
DFFARX1 I_49923 (I290181,I2683,I851348,I851422,);
not I_49924 (I851430,I290163);
not I_49925 (I851447,I290184);
nand I_49926 (I851464,I851447,I851430);
nor I_49927 (I851319,I851422,I851464);
DFFARX1 I_49928 (I851464,I2683,I851348,I851504,);
not I_49929 (I851340,I851504);
not I_49930 (I851526,I290187);
nand I_49931 (I851543,I851447,I851526);
DFFARX1 I_49932 (I851543,I2683,I851348,I851569,);
not I_49933 (I851577,I851569);
not I_49934 (I851594,I290178);
nand I_49935 (I851611,I851594,I290166);
and I_49936 (I851628,I851430,I851611);
nor I_49937 (I851645,I851543,I851628);
DFFARX1 I_49938 (I851645,I2683,I851348,I851316,);
DFFARX1 I_49939 (I851628,I2683,I851348,I851337,);
nor I_49940 (I851690,I290178,I290172);
nor I_49941 (I851328,I851543,I851690);
or I_49942 (I851721,I290178,I290172);
nor I_49943 (I851738,I290169,I290163);
DFFARX1 I_49944 (I851738,I2683,I851348,I851764,);
not I_49945 (I851772,I851764);
nor I_49946 (I851334,I851772,I851577);
nand I_49947 (I851803,I851772,I851422);
not I_49948 (I851820,I290169);
nand I_49949 (I851837,I851820,I851526);
nand I_49950 (I851854,I851772,I851837);
nand I_49951 (I851325,I851854,I851803);
nand I_49952 (I851322,I851837,I851721);
not I_49953 (I851926,I2690);
DFFARX1 I_49954 (I597147,I2683,I851926,I851952,);
and I_49955 (I851960,I851952,I597135);
DFFARX1 I_49956 (I851960,I2683,I851926,I851909,);
DFFARX1 I_49957 (I597138,I2683,I851926,I852000,);
not I_49958 (I852008,I597132);
not I_49959 (I852025,I597156);
nand I_49960 (I852042,I852025,I852008);
nor I_49961 (I851897,I852000,I852042);
DFFARX1 I_49962 (I852042,I2683,I851926,I852082,);
not I_49963 (I851918,I852082);
not I_49964 (I852104,I597144);
nand I_49965 (I852121,I852025,I852104);
DFFARX1 I_49966 (I852121,I2683,I851926,I852147,);
not I_49967 (I852155,I852147);
not I_49968 (I852172,I597153);
nand I_49969 (I852189,I852172,I597150);
and I_49970 (I852206,I852008,I852189);
nor I_49971 (I852223,I852121,I852206);
DFFARX1 I_49972 (I852223,I2683,I851926,I851894,);
DFFARX1 I_49973 (I852206,I2683,I851926,I851915,);
nor I_49974 (I852268,I597153,I597141);
nor I_49975 (I851906,I852121,I852268);
or I_49976 (I852299,I597153,I597141);
nor I_49977 (I852316,I597132,I597135);
DFFARX1 I_49978 (I852316,I2683,I851926,I852342,);
not I_49979 (I852350,I852342);
nor I_49980 (I851912,I852350,I852155);
nand I_49981 (I852381,I852350,I852000);
not I_49982 (I852398,I597132);
nand I_49983 (I852415,I852398,I852104);
nand I_49984 (I852432,I852350,I852415);
nand I_49985 (I851903,I852432,I852381);
nand I_49986 (I851900,I852415,I852299);
not I_49987 (I852504,I2690);
DFFARX1 I_49988 (I217991,I2683,I852504,I852530,);
and I_49989 (I852538,I852530,I217976);
DFFARX1 I_49990 (I852538,I2683,I852504,I852487,);
DFFARX1 I_49991 (I217982,I2683,I852504,I852578,);
not I_49992 (I852586,I217964);
not I_49993 (I852603,I217985);
nand I_49994 (I852620,I852603,I852586);
nor I_49995 (I852475,I852578,I852620);
DFFARX1 I_49996 (I852620,I2683,I852504,I852660,);
not I_49997 (I852496,I852660);
not I_49998 (I852682,I217988);
nand I_49999 (I852699,I852603,I852682);
DFFARX1 I_50000 (I852699,I2683,I852504,I852725,);
not I_50001 (I852733,I852725);
not I_50002 (I852750,I217979);
nand I_50003 (I852767,I852750,I217967);
and I_50004 (I852784,I852586,I852767);
nor I_50005 (I852801,I852699,I852784);
DFFARX1 I_50006 (I852801,I2683,I852504,I852472,);
DFFARX1 I_50007 (I852784,I2683,I852504,I852493,);
nor I_50008 (I852846,I217979,I217973);
nor I_50009 (I852484,I852699,I852846);
or I_50010 (I852877,I217979,I217973);
nor I_50011 (I852894,I217970,I217964);
DFFARX1 I_50012 (I852894,I2683,I852504,I852920,);
not I_50013 (I852928,I852920);
nor I_50014 (I852490,I852928,I852733);
nand I_50015 (I852959,I852928,I852578);
not I_50016 (I852976,I217970);
nand I_50017 (I852993,I852976,I852682);
nand I_50018 (I853010,I852928,I852993);
nand I_50019 (I852481,I853010,I852959);
nand I_50020 (I852478,I852993,I852877);
not I_50021 (I853082,I2690);
DFFARX1 I_50022 (I662313,I2683,I853082,I853108,);
and I_50023 (I853116,I853108,I662319);
DFFARX1 I_50024 (I853116,I2683,I853082,I853065,);
DFFARX1 I_50025 (I662325,I2683,I853082,I853156,);
not I_50026 (I853164,I662310);
not I_50027 (I853181,I662310);
nand I_50028 (I853198,I853181,I853164);
nor I_50029 (I853053,I853156,I853198);
DFFARX1 I_50030 (I853198,I2683,I853082,I853238,);
not I_50031 (I853074,I853238);
not I_50032 (I853260,I662328);
nand I_50033 (I853277,I853181,I853260);
DFFARX1 I_50034 (I853277,I2683,I853082,I853303,);
not I_50035 (I853311,I853303);
not I_50036 (I853328,I662322);
nand I_50037 (I853345,I853328,I662313);
and I_50038 (I853362,I853164,I853345);
nor I_50039 (I853379,I853277,I853362);
DFFARX1 I_50040 (I853379,I2683,I853082,I853050,);
DFFARX1 I_50041 (I853362,I2683,I853082,I853071,);
nor I_50042 (I853424,I662322,I662331);
nor I_50043 (I853062,I853277,I853424);
or I_50044 (I853455,I662322,I662331);
nor I_50045 (I853472,I662316,I662316);
DFFARX1 I_50046 (I853472,I2683,I853082,I853498,);
not I_50047 (I853506,I853498);
nor I_50048 (I853068,I853506,I853311);
nand I_50049 (I853537,I853506,I853156);
not I_50050 (I853554,I662316);
nand I_50051 (I853571,I853554,I853260);
nand I_50052 (I853588,I853506,I853571);
nand I_50053 (I853059,I853588,I853537);
nand I_50054 (I853056,I853571,I853455);
not I_50055 (I853660,I2690);
DFFARX1 I_50056 (I452647,I2683,I853660,I853686,);
and I_50057 (I853694,I853686,I452635);
DFFARX1 I_50058 (I853694,I2683,I853660,I853643,);
DFFARX1 I_50059 (I452650,I2683,I853660,I853734,);
not I_50060 (I853742,I452641);
not I_50061 (I853759,I452632);
nand I_50062 (I853776,I853759,I853742);
nor I_50063 (I853631,I853734,I853776);
DFFARX1 I_50064 (I853776,I2683,I853660,I853816,);
not I_50065 (I853652,I853816);
not I_50066 (I853838,I452638);
nand I_50067 (I853855,I853759,I853838);
DFFARX1 I_50068 (I853855,I2683,I853660,I853881,);
not I_50069 (I853889,I853881);
not I_50070 (I853906,I452653);
nand I_50071 (I853923,I853906,I452656);
and I_50072 (I853940,I853742,I853923);
nor I_50073 (I853957,I853855,I853940);
DFFARX1 I_50074 (I853957,I2683,I853660,I853628,);
DFFARX1 I_50075 (I853940,I2683,I853660,I853649,);
nor I_50076 (I854002,I452653,I452632);
nor I_50077 (I853640,I853855,I854002);
or I_50078 (I854033,I452653,I452632);
nor I_50079 (I854050,I452644,I452635);
DFFARX1 I_50080 (I854050,I2683,I853660,I854076,);
not I_50081 (I854084,I854076);
nor I_50082 (I853646,I854084,I853889);
nand I_50083 (I854115,I854084,I853734);
not I_50084 (I854132,I452644);
nand I_50085 (I854149,I854132,I853838);
nand I_50086 (I854166,I854084,I854149);
nand I_50087 (I853637,I854166,I854115);
nand I_50088 (I853634,I854149,I854033);
not I_50089 (I854238,I2690);
DFFARX1 I_50090 (I11038,I2683,I854238,I854264,);
and I_50091 (I854272,I854264,I11044);
DFFARX1 I_50092 (I854272,I2683,I854238,I854221,);
DFFARX1 I_50093 (I11023,I2683,I854238,I854312,);
not I_50094 (I854320,I11029);
not I_50095 (I854337,I11035);
nand I_50096 (I854354,I854337,I854320);
nor I_50097 (I854209,I854312,I854354);
DFFARX1 I_50098 (I854354,I2683,I854238,I854394,);
not I_50099 (I854230,I854394);
not I_50100 (I854416,I11026);
nand I_50101 (I854433,I854337,I854416);
DFFARX1 I_50102 (I854433,I2683,I854238,I854459,);
not I_50103 (I854467,I854459);
not I_50104 (I854484,I11041);
nand I_50105 (I854501,I854484,I11026);
and I_50106 (I854518,I854320,I854501);
nor I_50107 (I854535,I854433,I854518);
DFFARX1 I_50108 (I854535,I2683,I854238,I854206,);
DFFARX1 I_50109 (I854518,I2683,I854238,I854227,);
nor I_50110 (I854580,I11041,I11029);
nor I_50111 (I854218,I854433,I854580);
or I_50112 (I854611,I11041,I11029);
nor I_50113 (I854628,I11032,I11023);
DFFARX1 I_50114 (I854628,I2683,I854238,I854654,);
not I_50115 (I854662,I854654);
nor I_50116 (I854224,I854662,I854467);
nand I_50117 (I854693,I854662,I854312);
not I_50118 (I854710,I11032);
nand I_50119 (I854727,I854710,I854416);
nand I_50120 (I854744,I854662,I854727);
nand I_50121 (I854215,I854744,I854693);
nand I_50122 (I854212,I854727,I854611);
not I_50123 (I854816,I2690);
DFFARX1 I_50124 (I674434,I2683,I854816,I854842,);
and I_50125 (I854850,I854842,I674440);
DFFARX1 I_50126 (I854850,I2683,I854816,I854799,);
DFFARX1 I_50127 (I674446,I2683,I854816,I854890,);
not I_50128 (I854898,I674431);
not I_50129 (I854915,I674431);
nand I_50130 (I854932,I854915,I854898);
nor I_50131 (I854787,I854890,I854932);
DFFARX1 I_50132 (I854932,I2683,I854816,I854972,);
not I_50133 (I854808,I854972);
not I_50134 (I854994,I674449);
nand I_50135 (I855011,I854915,I854994);
DFFARX1 I_50136 (I855011,I2683,I854816,I855037,);
not I_50137 (I855045,I855037);
not I_50138 (I855062,I674443);
nand I_50139 (I855079,I855062,I674434);
and I_50140 (I855096,I854898,I855079);
nor I_50141 (I855113,I855011,I855096);
DFFARX1 I_50142 (I855113,I2683,I854816,I854784,);
DFFARX1 I_50143 (I855096,I2683,I854816,I854805,);
nor I_50144 (I855158,I674443,I674452);
nor I_50145 (I854796,I855011,I855158);
or I_50146 (I855189,I674443,I674452);
nor I_50147 (I855206,I674437,I674437);
DFFARX1 I_50148 (I855206,I2683,I854816,I855232,);
not I_50149 (I855240,I855232);
nor I_50150 (I854802,I855240,I855045);
nand I_50151 (I855271,I855240,I854890);
not I_50152 (I855288,I674437);
nand I_50153 (I855305,I855288,I854994);
nand I_50154 (I855322,I855240,I855305);
nand I_50155 (I854793,I855322,I855271);
nand I_50156 (I854790,I855305,I855189);
not I_50157 (I855394,I2690);
DFFARX1 I_50158 (I109137,I2683,I855394,I855420,);
and I_50159 (I855428,I855420,I109113);
DFFARX1 I_50160 (I855428,I2683,I855394,I855377,);
DFFARX1 I_50161 (I109131,I2683,I855394,I855468,);
not I_50162 (I855476,I109119);
not I_50163 (I855493,I109116);
nand I_50164 (I855510,I855493,I855476);
nor I_50165 (I855365,I855468,I855510);
DFFARX1 I_50166 (I855510,I2683,I855394,I855550,);
not I_50167 (I855386,I855550);
not I_50168 (I855572,I109125);
nand I_50169 (I855589,I855493,I855572);
DFFARX1 I_50170 (I855589,I2683,I855394,I855615,);
not I_50171 (I855623,I855615);
not I_50172 (I855640,I109116);
nand I_50173 (I855657,I855640,I109134);
and I_50174 (I855674,I855476,I855657);
nor I_50175 (I855691,I855589,I855674);
DFFARX1 I_50176 (I855691,I2683,I855394,I855362,);
DFFARX1 I_50177 (I855674,I2683,I855394,I855383,);
nor I_50178 (I855736,I109116,I109128);
nor I_50179 (I855374,I855589,I855736);
or I_50180 (I855767,I109116,I109128);
nor I_50181 (I855784,I109122,I109113);
DFFARX1 I_50182 (I855784,I2683,I855394,I855810,);
not I_50183 (I855818,I855810);
nor I_50184 (I855380,I855818,I855623);
nand I_50185 (I855849,I855818,I855468);
not I_50186 (I855866,I109122);
nand I_50187 (I855883,I855866,I855572);
nand I_50188 (I855900,I855818,I855883);
nand I_50189 (I855371,I855900,I855849);
nand I_50190 (I855368,I855883,I855767);
not I_50191 (I855972,I2690);
DFFARX1 I_50192 (I83841,I2683,I855972,I855998,);
and I_50193 (I856006,I855998,I83817);
DFFARX1 I_50194 (I856006,I2683,I855972,I855955,);
DFFARX1 I_50195 (I83835,I2683,I855972,I856046,);
not I_50196 (I856054,I83823);
not I_50197 (I856071,I83820);
nand I_50198 (I856088,I856071,I856054);
nor I_50199 (I855943,I856046,I856088);
DFFARX1 I_50200 (I856088,I2683,I855972,I856128,);
not I_50201 (I855964,I856128);
not I_50202 (I856150,I83829);
nand I_50203 (I856167,I856071,I856150);
DFFARX1 I_50204 (I856167,I2683,I855972,I856193,);
not I_50205 (I856201,I856193);
not I_50206 (I856218,I83820);
nand I_50207 (I856235,I856218,I83838);
and I_50208 (I856252,I856054,I856235);
nor I_50209 (I856269,I856167,I856252);
DFFARX1 I_50210 (I856269,I2683,I855972,I855940,);
DFFARX1 I_50211 (I856252,I2683,I855972,I855961,);
nor I_50212 (I856314,I83820,I83832);
nor I_50213 (I855952,I856167,I856314);
or I_50214 (I856345,I83820,I83832);
nor I_50215 (I856362,I83826,I83817);
DFFARX1 I_50216 (I856362,I2683,I855972,I856388,);
not I_50217 (I856396,I856388);
nor I_50218 (I855958,I856396,I856201);
nand I_50219 (I856427,I856396,I856046);
not I_50220 (I856444,I83826);
nand I_50221 (I856461,I856444,I856150);
nand I_50222 (I856478,I856396,I856461);
nand I_50223 (I855949,I856478,I856427);
nand I_50224 (I855946,I856461,I856345);
not I_50225 (I856550,I2690);
DFFARX1 I_50226 (I383442,I2683,I856550,I856576,);
and I_50227 (I856584,I856576,I383457);
DFFARX1 I_50228 (I856584,I2683,I856550,I856533,);
DFFARX1 I_50229 (I383460,I2683,I856550,I856624,);
not I_50230 (I856632,I383454);
not I_50231 (I856649,I383469);
nand I_50232 (I856666,I856649,I856632);
nor I_50233 (I856521,I856624,I856666);
DFFARX1 I_50234 (I856666,I2683,I856550,I856706,);
not I_50235 (I856542,I856706);
not I_50236 (I856728,I383445);
nand I_50237 (I856745,I856649,I856728);
DFFARX1 I_50238 (I856745,I2683,I856550,I856771,);
not I_50239 (I856779,I856771);
not I_50240 (I856796,I383448);
nand I_50241 (I856813,I856796,I383442);
and I_50242 (I856830,I856632,I856813);
nor I_50243 (I856847,I856745,I856830);
DFFARX1 I_50244 (I856847,I2683,I856550,I856518,);
DFFARX1 I_50245 (I856830,I2683,I856550,I856539,);
nor I_50246 (I856892,I383448,I383451);
nor I_50247 (I856530,I856745,I856892);
or I_50248 (I856923,I383448,I383451);
nor I_50249 (I856940,I383466,I383463);
DFFARX1 I_50250 (I856940,I2683,I856550,I856966,);
not I_50251 (I856974,I856966);
nor I_50252 (I856536,I856974,I856779);
nand I_50253 (I857005,I856974,I856624);
not I_50254 (I857022,I383466);
nand I_50255 (I857039,I857022,I856728);
nand I_50256 (I857056,I856974,I857039);
nand I_50257 (I856527,I857056,I857005);
nand I_50258 (I856524,I857039,I856923);
not I_50259 (I857128,I2690);
DFFARX1 I_50260 (I532411,I2683,I857128,I857154,);
and I_50261 (I857162,I857154,I532399);
DFFARX1 I_50262 (I857162,I2683,I857128,I857111,);
DFFARX1 I_50263 (I532402,I2683,I857128,I857202,);
not I_50264 (I857210,I532396);
not I_50265 (I857227,I532420);
nand I_50266 (I857244,I857227,I857210);
nor I_50267 (I857099,I857202,I857244);
DFFARX1 I_50268 (I857244,I2683,I857128,I857284,);
not I_50269 (I857120,I857284);
not I_50270 (I857306,I532408);
nand I_50271 (I857323,I857227,I857306);
DFFARX1 I_50272 (I857323,I2683,I857128,I857349,);
not I_50273 (I857357,I857349);
not I_50274 (I857374,I532417);
nand I_50275 (I857391,I857374,I532414);
and I_50276 (I857408,I857210,I857391);
nor I_50277 (I857425,I857323,I857408);
DFFARX1 I_50278 (I857425,I2683,I857128,I857096,);
DFFARX1 I_50279 (I857408,I2683,I857128,I857117,);
nor I_50280 (I857470,I532417,I532405);
nor I_50281 (I857108,I857323,I857470);
or I_50282 (I857501,I532417,I532405);
nor I_50283 (I857518,I532396,I532399);
DFFARX1 I_50284 (I857518,I2683,I857128,I857544,);
not I_50285 (I857552,I857544);
nor I_50286 (I857114,I857552,I857357);
nand I_50287 (I857583,I857552,I857202);
not I_50288 (I857600,I532396);
nand I_50289 (I857617,I857600,I857306);
nand I_50290 (I857634,I857552,I857617);
nand I_50291 (I857105,I857634,I857583);
nand I_50292 (I857102,I857617,I857501);
not I_50293 (I857706,I2690);
DFFARX1 I_50294 (I611597,I2683,I857706,I857732,);
and I_50295 (I857740,I857732,I611585);
DFFARX1 I_50296 (I857740,I2683,I857706,I857689,);
DFFARX1 I_50297 (I611588,I2683,I857706,I857780,);
not I_50298 (I857788,I611582);
not I_50299 (I857805,I611606);
nand I_50300 (I857822,I857805,I857788);
nor I_50301 (I857677,I857780,I857822);
DFFARX1 I_50302 (I857822,I2683,I857706,I857862,);
not I_50303 (I857698,I857862);
not I_50304 (I857884,I611594);
nand I_50305 (I857901,I857805,I857884);
DFFARX1 I_50306 (I857901,I2683,I857706,I857927,);
not I_50307 (I857935,I857927);
not I_50308 (I857952,I611603);
nand I_50309 (I857969,I857952,I611600);
and I_50310 (I857986,I857788,I857969);
nor I_50311 (I858003,I857901,I857986);
DFFARX1 I_50312 (I858003,I2683,I857706,I857674,);
DFFARX1 I_50313 (I857986,I2683,I857706,I857695,);
nor I_50314 (I858048,I611603,I611591);
nor I_50315 (I857686,I857901,I858048);
or I_50316 (I858079,I611603,I611591);
nor I_50317 (I858096,I611582,I611585);
DFFARX1 I_50318 (I858096,I2683,I857706,I858122,);
not I_50319 (I858130,I858122);
nor I_50320 (I857692,I858130,I857935);
nand I_50321 (I858161,I858130,I857780);
not I_50322 (I858178,I611582);
nand I_50323 (I858195,I858178,I857884);
nand I_50324 (I858212,I858130,I858195);
nand I_50325 (I857683,I858212,I858161);
nand I_50326 (I857680,I858195,I858079);
not I_50327 (I858284,I2690);
DFFARX1 I_50328 (I561311,I2683,I858284,I858310,);
and I_50329 (I858318,I858310,I561299);
DFFARX1 I_50330 (I858318,I2683,I858284,I858267,);
DFFARX1 I_50331 (I561302,I2683,I858284,I858358,);
not I_50332 (I858366,I561296);
not I_50333 (I858383,I561320);
nand I_50334 (I858400,I858383,I858366);
nor I_50335 (I858255,I858358,I858400);
DFFARX1 I_50336 (I858400,I2683,I858284,I858440,);
not I_50337 (I858276,I858440);
not I_50338 (I858462,I561308);
nand I_50339 (I858479,I858383,I858462);
DFFARX1 I_50340 (I858479,I2683,I858284,I858505,);
not I_50341 (I858513,I858505);
not I_50342 (I858530,I561317);
nand I_50343 (I858547,I858530,I561314);
and I_50344 (I858564,I858366,I858547);
nor I_50345 (I858581,I858479,I858564);
DFFARX1 I_50346 (I858581,I2683,I858284,I858252,);
DFFARX1 I_50347 (I858564,I2683,I858284,I858273,);
nor I_50348 (I858626,I561317,I561305);
nor I_50349 (I858264,I858479,I858626);
or I_50350 (I858657,I561317,I561305);
nor I_50351 (I858674,I561296,I561299);
DFFARX1 I_50352 (I858674,I2683,I858284,I858700,);
not I_50353 (I858708,I858700);
nor I_50354 (I858270,I858708,I858513);
nand I_50355 (I858739,I858708,I858358);
not I_50356 (I858756,I561296);
nand I_50357 (I858773,I858756,I858462);
nand I_50358 (I858790,I858708,I858773);
nand I_50359 (I858261,I858790,I858739);
nand I_50360 (I858258,I858773,I858657);
not I_50361 (I858862,I2690);
DFFARX1 I_50362 (I564779,I2683,I858862,I858888,);
and I_50363 (I858896,I858888,I564767);
DFFARX1 I_50364 (I858896,I2683,I858862,I858845,);
DFFARX1 I_50365 (I564770,I2683,I858862,I858936,);
not I_50366 (I858944,I564764);
not I_50367 (I858961,I564788);
nand I_50368 (I858978,I858961,I858944);
nor I_50369 (I858833,I858936,I858978);
DFFARX1 I_50370 (I858978,I2683,I858862,I859018,);
not I_50371 (I858854,I859018);
not I_50372 (I859040,I564776);
nand I_50373 (I859057,I858961,I859040);
DFFARX1 I_50374 (I859057,I2683,I858862,I859083,);
not I_50375 (I859091,I859083);
not I_50376 (I859108,I564785);
nand I_50377 (I859125,I859108,I564782);
and I_50378 (I859142,I858944,I859125);
nor I_50379 (I859159,I859057,I859142);
DFFARX1 I_50380 (I859159,I2683,I858862,I858830,);
DFFARX1 I_50381 (I859142,I2683,I858862,I858851,);
nor I_50382 (I859204,I564785,I564773);
nor I_50383 (I858842,I859057,I859204);
or I_50384 (I859235,I564785,I564773);
nor I_50385 (I859252,I564764,I564767);
DFFARX1 I_50386 (I859252,I2683,I858862,I859278,);
not I_50387 (I859286,I859278);
nor I_50388 (I858848,I859286,I859091);
nand I_50389 (I859317,I859286,I858936);
not I_50390 (I859334,I564764);
nand I_50391 (I859351,I859334,I859040);
nand I_50392 (I859368,I859286,I859351);
nand I_50393 (I858839,I859368,I859317);
nand I_50394 (I858836,I859351,I859235);
not I_50395 (I859440,I2690);
DFFARX1 I_50396 (I133695,I2683,I859440,I859466,);
and I_50397 (I859474,I859466,I133698);
DFFARX1 I_50398 (I859474,I2683,I859440,I859423,);
DFFARX1 I_50399 (I133698,I2683,I859440,I859514,);
not I_50400 (I859522,I133713);
not I_50401 (I859539,I133719);
nand I_50402 (I859556,I859539,I859522);
nor I_50403 (I859411,I859514,I859556);
DFFARX1 I_50404 (I859556,I2683,I859440,I859596,);
not I_50405 (I859432,I859596);
not I_50406 (I859618,I133707);
nand I_50407 (I859635,I859539,I859618);
DFFARX1 I_50408 (I859635,I2683,I859440,I859661,);
not I_50409 (I859669,I859661);
not I_50410 (I859686,I133704);
nand I_50411 (I859703,I859686,I133701);
and I_50412 (I859720,I859522,I859703);
nor I_50413 (I859737,I859635,I859720);
DFFARX1 I_50414 (I859737,I2683,I859440,I859408,);
DFFARX1 I_50415 (I859720,I2683,I859440,I859429,);
nor I_50416 (I859782,I133704,I133695);
nor I_50417 (I859420,I859635,I859782);
or I_50418 (I859813,I133704,I133695);
nor I_50419 (I859830,I133710,I133716);
DFFARX1 I_50420 (I859830,I2683,I859440,I859856,);
not I_50421 (I859864,I859856);
nor I_50422 (I859426,I859864,I859669);
nand I_50423 (I859895,I859864,I859514);
not I_50424 (I859912,I133710);
nand I_50425 (I859929,I859912,I859618);
nand I_50426 (I859946,I859864,I859929);
nand I_50427 (I859417,I859946,I859895);
nand I_50428 (I859414,I859929,I859813);
not I_50429 (I860018,I2690);
DFFARX1 I_50430 (I344274,I2683,I860018,I860044,);
and I_50431 (I860052,I860044,I344289);
DFFARX1 I_50432 (I860052,I2683,I860018,I860001,);
DFFARX1 I_50433 (I344292,I2683,I860018,I860092,);
not I_50434 (I860100,I344286);
not I_50435 (I860117,I344301);
nand I_50436 (I860134,I860117,I860100);
nor I_50437 (I859989,I860092,I860134);
DFFARX1 I_50438 (I860134,I2683,I860018,I860174,);
not I_50439 (I860010,I860174);
not I_50440 (I860196,I344277);
nand I_50441 (I860213,I860117,I860196);
DFFARX1 I_50442 (I860213,I2683,I860018,I860239,);
not I_50443 (I860247,I860239);
not I_50444 (I860264,I344280);
nand I_50445 (I860281,I860264,I344274);
and I_50446 (I860298,I860100,I860281);
nor I_50447 (I860315,I860213,I860298);
DFFARX1 I_50448 (I860315,I2683,I860018,I859986,);
DFFARX1 I_50449 (I860298,I2683,I860018,I860007,);
nor I_50450 (I860360,I344280,I344283);
nor I_50451 (I859998,I860213,I860360);
or I_50452 (I860391,I344280,I344283);
nor I_50453 (I860408,I344298,I344295);
DFFARX1 I_50454 (I860408,I2683,I860018,I860434,);
not I_50455 (I860442,I860434);
nor I_50456 (I860004,I860442,I860247);
nand I_50457 (I860473,I860442,I860092);
not I_50458 (I860490,I344298);
nand I_50459 (I860507,I860490,I860196);
nand I_50460 (I860524,I860442,I860507);
nand I_50461 (I859995,I860524,I860473);
nand I_50462 (I859992,I860507,I860391);
not I_50463 (I860596,I2690);
DFFARX1 I_50464 (I347538,I2683,I860596,I860622,);
and I_50465 (I860630,I860622,I347553);
DFFARX1 I_50466 (I860630,I2683,I860596,I860579,);
DFFARX1 I_50467 (I347556,I2683,I860596,I860670,);
not I_50468 (I860678,I347550);
not I_50469 (I860695,I347565);
nand I_50470 (I860712,I860695,I860678);
nor I_50471 (I860567,I860670,I860712);
DFFARX1 I_50472 (I860712,I2683,I860596,I860752,);
not I_50473 (I860588,I860752);
not I_50474 (I860774,I347541);
nand I_50475 (I860791,I860695,I860774);
DFFARX1 I_50476 (I860791,I2683,I860596,I860817,);
not I_50477 (I860825,I860817);
not I_50478 (I860842,I347544);
nand I_50479 (I860859,I860842,I347538);
and I_50480 (I860876,I860678,I860859);
nor I_50481 (I860893,I860791,I860876);
DFFARX1 I_50482 (I860893,I2683,I860596,I860564,);
DFFARX1 I_50483 (I860876,I2683,I860596,I860585,);
nor I_50484 (I860938,I347544,I347547);
nor I_50485 (I860576,I860791,I860938);
or I_50486 (I860969,I347544,I347547);
nor I_50487 (I860986,I347562,I347559);
DFFARX1 I_50488 (I860986,I2683,I860596,I861012,);
not I_50489 (I861020,I861012);
nor I_50490 (I860582,I861020,I860825);
nand I_50491 (I861051,I861020,I860670);
not I_50492 (I861068,I347562);
nand I_50493 (I861085,I861068,I860774);
nand I_50494 (I861102,I861020,I861085);
nand I_50495 (I860573,I861102,I861051);
nand I_50496 (I860570,I861085,I860969);
not I_50497 (I861174,I2690);
DFFARX1 I_50498 (I763279,I2683,I861174,I861200,);
and I_50499 (I861208,I861200,I763273);
DFFARX1 I_50500 (I861208,I2683,I861174,I861157,);
DFFARX1 I_50501 (I763291,I2683,I861174,I861248,);
not I_50502 (I861256,I763282);
not I_50503 (I861273,I763294);
nand I_50504 (I861290,I861273,I861256);
nor I_50505 (I861145,I861248,I861290);
DFFARX1 I_50506 (I861290,I2683,I861174,I861330,);
not I_50507 (I861166,I861330);
not I_50508 (I861352,I763300);
nand I_50509 (I861369,I861273,I861352);
DFFARX1 I_50510 (I861369,I2683,I861174,I861395,);
not I_50511 (I861403,I861395);
not I_50512 (I861420,I763276);
nand I_50513 (I861437,I861420,I763297);
and I_50514 (I861454,I861256,I861437);
nor I_50515 (I861471,I861369,I861454);
DFFARX1 I_50516 (I861471,I2683,I861174,I861142,);
DFFARX1 I_50517 (I861454,I2683,I861174,I861163,);
nor I_50518 (I861516,I763276,I763288);
nor I_50519 (I861154,I861369,I861516);
or I_50520 (I861547,I763276,I763288);
nor I_50521 (I861564,I763273,I763285);
DFFARX1 I_50522 (I861564,I2683,I861174,I861590,);
not I_50523 (I861598,I861590);
nor I_50524 (I861160,I861598,I861403);
nand I_50525 (I861629,I861598,I861248);
not I_50526 (I861646,I763273);
nand I_50527 (I861663,I861646,I861352);
nand I_50528 (I861680,I861598,I861663);
nand I_50529 (I861151,I861680,I861629);
nand I_50530 (I861148,I861663,I861547);
not I_50531 (I861752,I2690);
DFFARX1 I_50532 (I497153,I2683,I861752,I861778,);
and I_50533 (I861786,I861778,I497141);
DFFARX1 I_50534 (I861786,I2683,I861752,I861735,);
DFFARX1 I_50535 (I497144,I2683,I861752,I861826,);
not I_50536 (I861834,I497138);
not I_50537 (I861851,I497162);
nand I_50538 (I861868,I861851,I861834);
nor I_50539 (I861723,I861826,I861868);
DFFARX1 I_50540 (I861868,I2683,I861752,I861908,);
not I_50541 (I861744,I861908);
not I_50542 (I861930,I497150);
nand I_50543 (I861947,I861851,I861930);
DFFARX1 I_50544 (I861947,I2683,I861752,I861973,);
not I_50545 (I861981,I861973);
not I_50546 (I861998,I497159);
nand I_50547 (I862015,I861998,I497156);
and I_50548 (I862032,I861834,I862015);
nor I_50549 (I862049,I861947,I862032);
DFFARX1 I_50550 (I862049,I2683,I861752,I861720,);
DFFARX1 I_50551 (I862032,I2683,I861752,I861741,);
nor I_50552 (I862094,I497159,I497147);
nor I_50553 (I861732,I861947,I862094);
or I_50554 (I862125,I497159,I497147);
nor I_50555 (I862142,I497138,I497141);
DFFARX1 I_50556 (I862142,I2683,I861752,I862168,);
not I_50557 (I862176,I862168);
nor I_50558 (I861738,I862176,I861981);
nand I_50559 (I862207,I862176,I861826);
not I_50560 (I862224,I497138);
nand I_50561 (I862241,I862224,I861930);
nand I_50562 (I862258,I862176,I862241);
nand I_50563 (I861729,I862258,I862207);
nand I_50564 (I861726,I862241,I862125);
not I_50565 (I862330,I2690);
DFFARX1 I_50566 (I372562,I2683,I862330,I862356,);
and I_50567 (I862364,I862356,I372577);
DFFARX1 I_50568 (I862364,I2683,I862330,I862313,);
DFFARX1 I_50569 (I372580,I2683,I862330,I862404,);
not I_50570 (I862412,I372574);
not I_50571 (I862429,I372589);
nand I_50572 (I862446,I862429,I862412);
nor I_50573 (I862301,I862404,I862446);
DFFARX1 I_50574 (I862446,I2683,I862330,I862486,);
not I_50575 (I862322,I862486);
not I_50576 (I862508,I372565);
nand I_50577 (I862525,I862429,I862508);
DFFARX1 I_50578 (I862525,I2683,I862330,I862551,);
not I_50579 (I862559,I862551);
not I_50580 (I862576,I372568);
nand I_50581 (I862593,I862576,I372562);
and I_50582 (I862610,I862412,I862593);
nor I_50583 (I862627,I862525,I862610);
DFFARX1 I_50584 (I862627,I2683,I862330,I862298,);
DFFARX1 I_50585 (I862610,I2683,I862330,I862319,);
nor I_50586 (I862672,I372568,I372571);
nor I_50587 (I862310,I862525,I862672);
or I_50588 (I862703,I372568,I372571);
nor I_50589 (I862720,I372586,I372583);
DFFARX1 I_50590 (I862720,I2683,I862330,I862746,);
not I_50591 (I862754,I862746);
nor I_50592 (I862316,I862754,I862559);
nand I_50593 (I862785,I862754,I862404);
not I_50594 (I862802,I372586);
nand I_50595 (I862819,I862802,I862508);
nand I_50596 (I862836,I862754,I862819);
nand I_50597 (I862307,I862836,I862785);
nand I_50598 (I862304,I862819,I862703);
not I_50599 (I862908,I2690);
DFFARX1 I_50600 (I647030,I2683,I862908,I862934,);
and I_50601 (I862942,I862934,I647036);
DFFARX1 I_50602 (I862942,I2683,I862908,I862891,);
DFFARX1 I_50603 (I647042,I2683,I862908,I862982,);
not I_50604 (I862990,I647027);
not I_50605 (I863007,I647027);
nand I_50606 (I863024,I863007,I862990);
nor I_50607 (I862879,I862982,I863024);
DFFARX1 I_50608 (I863024,I2683,I862908,I863064,);
not I_50609 (I862900,I863064);
not I_50610 (I863086,I647045);
nand I_50611 (I863103,I863007,I863086);
DFFARX1 I_50612 (I863103,I2683,I862908,I863129,);
not I_50613 (I863137,I863129);
not I_50614 (I863154,I647039);
nand I_50615 (I863171,I863154,I647030);
and I_50616 (I863188,I862990,I863171);
nor I_50617 (I863205,I863103,I863188);
DFFARX1 I_50618 (I863205,I2683,I862908,I862876,);
DFFARX1 I_50619 (I863188,I2683,I862908,I862897,);
nor I_50620 (I863250,I647039,I647048);
nor I_50621 (I862888,I863103,I863250);
or I_50622 (I863281,I647039,I647048);
nor I_50623 (I863298,I647033,I647033);
DFFARX1 I_50624 (I863298,I2683,I862908,I863324,);
not I_50625 (I863332,I863324);
nor I_50626 (I862894,I863332,I863137);
nand I_50627 (I863363,I863332,I862982);
not I_50628 (I863380,I647033);
nand I_50629 (I863397,I863380,I863086);
nand I_50630 (I863414,I863332,I863397);
nand I_50631 (I862885,I863414,I863363);
nand I_50632 (I862882,I863397,I863281);
not I_50633 (I863486,I2690);
DFFARX1 I_50634 (I59599,I2683,I863486,I863512,);
and I_50635 (I863520,I863512,I59575);
DFFARX1 I_50636 (I863520,I2683,I863486,I863469,);
DFFARX1 I_50637 (I59593,I2683,I863486,I863560,);
not I_50638 (I863568,I59581);
not I_50639 (I863585,I59578);
nand I_50640 (I863602,I863585,I863568);
nor I_50641 (I863457,I863560,I863602);
DFFARX1 I_50642 (I863602,I2683,I863486,I863642,);
not I_50643 (I863478,I863642);
not I_50644 (I863664,I59587);
nand I_50645 (I863681,I863585,I863664);
DFFARX1 I_50646 (I863681,I2683,I863486,I863707,);
not I_50647 (I863715,I863707);
not I_50648 (I863732,I59578);
nand I_50649 (I863749,I863732,I59596);
and I_50650 (I863766,I863568,I863749);
nor I_50651 (I863783,I863681,I863766);
DFFARX1 I_50652 (I863783,I2683,I863486,I863454,);
DFFARX1 I_50653 (I863766,I2683,I863486,I863475,);
nor I_50654 (I863828,I59578,I59590);
nor I_50655 (I863466,I863681,I863828);
or I_50656 (I863859,I59578,I59590);
nor I_50657 (I863876,I59584,I59575);
DFFARX1 I_50658 (I863876,I2683,I863486,I863902,);
not I_50659 (I863910,I863902);
nor I_50660 (I863472,I863910,I863715);
nand I_50661 (I863941,I863910,I863560);
not I_50662 (I863958,I59584);
nand I_50663 (I863975,I863958,I863664);
nand I_50664 (I863992,I863910,I863975);
nand I_50665 (I863463,I863992,I863941);
nand I_50666 (I863460,I863975,I863859);
not I_50667 (I864064,I2690);
DFFARX1 I_50668 (I477501,I2683,I864064,I864090,);
and I_50669 (I864098,I864090,I477489);
DFFARX1 I_50670 (I864098,I2683,I864064,I864047,);
DFFARX1 I_50671 (I477504,I2683,I864064,I864138,);
not I_50672 (I864146,I477495);
not I_50673 (I864163,I477486);
nand I_50674 (I864180,I864163,I864146);
nor I_50675 (I864035,I864138,I864180);
DFFARX1 I_50676 (I864180,I2683,I864064,I864220,);
not I_50677 (I864056,I864220);
not I_50678 (I864242,I477492);
nand I_50679 (I864259,I864163,I864242);
DFFARX1 I_50680 (I864259,I2683,I864064,I864285,);
not I_50681 (I864293,I864285);
not I_50682 (I864310,I477507);
nand I_50683 (I864327,I864310,I477510);
and I_50684 (I864344,I864146,I864327);
nor I_50685 (I864361,I864259,I864344);
DFFARX1 I_50686 (I864361,I2683,I864064,I864032,);
DFFARX1 I_50687 (I864344,I2683,I864064,I864053,);
nor I_50688 (I864406,I477507,I477486);
nor I_50689 (I864044,I864259,I864406);
or I_50690 (I864437,I477507,I477486);
nor I_50691 (I864454,I477498,I477489);
DFFARX1 I_50692 (I864454,I2683,I864064,I864480,);
not I_50693 (I864488,I864480);
nor I_50694 (I864050,I864488,I864293);
nand I_50695 (I864519,I864488,I864138);
not I_50696 (I864536,I477498);
nand I_50697 (I864553,I864536,I864242);
nand I_50698 (I864570,I864488,I864553);
nand I_50699 (I864041,I864570,I864519);
nand I_50700 (I864038,I864553,I864437);
not I_50701 (I864642,I2690);
DFFARX1 I_50702 (I349170,I2683,I864642,I864668,);
and I_50703 (I864676,I864668,I349185);
DFFARX1 I_50704 (I864676,I2683,I864642,I864625,);
DFFARX1 I_50705 (I349188,I2683,I864642,I864716,);
not I_50706 (I864724,I349182);
not I_50707 (I864741,I349197);
nand I_50708 (I864758,I864741,I864724);
nor I_50709 (I864613,I864716,I864758);
DFFARX1 I_50710 (I864758,I2683,I864642,I864798,);
not I_50711 (I864634,I864798);
not I_50712 (I864820,I349173);
nand I_50713 (I864837,I864741,I864820);
DFFARX1 I_50714 (I864837,I2683,I864642,I864863,);
not I_50715 (I864871,I864863);
not I_50716 (I864888,I349176);
nand I_50717 (I864905,I864888,I349170);
and I_50718 (I864922,I864724,I864905);
nor I_50719 (I864939,I864837,I864922);
DFFARX1 I_50720 (I864939,I2683,I864642,I864610,);
DFFARX1 I_50721 (I864922,I2683,I864642,I864631,);
nor I_50722 (I864984,I349176,I349179);
nor I_50723 (I864622,I864837,I864984);
or I_50724 (I865015,I349176,I349179);
nor I_50725 (I865032,I349194,I349191);
DFFARX1 I_50726 (I865032,I2683,I864642,I865058,);
not I_50727 (I865066,I865058);
nor I_50728 (I864628,I865066,I864871);
nand I_50729 (I865097,I865066,I864716);
not I_50730 (I865114,I349194);
nand I_50731 (I865131,I865114,I864820);
nand I_50732 (I865148,I865066,I865131);
nand I_50733 (I864619,I865148,I865097);
nand I_50734 (I864616,I865131,I865015);
not I_50735 (I865220,I2690);
DFFARX1 I_50736 (I761341,I2683,I865220,I865246,);
and I_50737 (I865254,I865246,I761335);
DFFARX1 I_50738 (I865254,I2683,I865220,I865203,);
DFFARX1 I_50739 (I761353,I2683,I865220,I865294,);
not I_50740 (I865302,I761344);
not I_50741 (I865319,I761356);
nand I_50742 (I865336,I865319,I865302);
nor I_50743 (I865191,I865294,I865336);
DFFARX1 I_50744 (I865336,I2683,I865220,I865376,);
not I_50745 (I865212,I865376);
not I_50746 (I865398,I761362);
nand I_50747 (I865415,I865319,I865398);
DFFARX1 I_50748 (I865415,I2683,I865220,I865441,);
not I_50749 (I865449,I865441);
not I_50750 (I865466,I761338);
nand I_50751 (I865483,I865466,I761359);
and I_50752 (I865500,I865302,I865483);
nor I_50753 (I865517,I865415,I865500);
DFFARX1 I_50754 (I865517,I2683,I865220,I865188,);
DFFARX1 I_50755 (I865500,I2683,I865220,I865209,);
nor I_50756 (I865562,I761338,I761350);
nor I_50757 (I865200,I865415,I865562);
or I_50758 (I865593,I761338,I761350);
nor I_50759 (I865610,I761335,I761347);
DFFARX1 I_50760 (I865610,I2683,I865220,I865636,);
not I_50761 (I865644,I865636);
nor I_50762 (I865206,I865644,I865449);
nand I_50763 (I865675,I865644,I865294);
not I_50764 (I865692,I761335);
nand I_50765 (I865709,I865692,I865398);
nand I_50766 (I865726,I865644,I865709);
nand I_50767 (I865197,I865726,I865675);
nand I_50768 (I865194,I865709,I865593);
not I_50769 (I865798,I2690);
DFFARX1 I_50770 (I517383,I2683,I865798,I865824,);
and I_50771 (I865832,I865824,I517371);
DFFARX1 I_50772 (I865832,I2683,I865798,I865781,);
DFFARX1 I_50773 (I517374,I2683,I865798,I865872,);
not I_50774 (I865880,I517368);
not I_50775 (I865897,I517392);
nand I_50776 (I865914,I865897,I865880);
nor I_50777 (I865769,I865872,I865914);
DFFARX1 I_50778 (I865914,I2683,I865798,I865954,);
not I_50779 (I865790,I865954);
not I_50780 (I865976,I517380);
nand I_50781 (I865993,I865897,I865976);
DFFARX1 I_50782 (I865993,I2683,I865798,I866019,);
not I_50783 (I866027,I866019);
not I_50784 (I866044,I517389);
nand I_50785 (I866061,I866044,I517386);
and I_50786 (I866078,I865880,I866061);
nor I_50787 (I866095,I865993,I866078);
DFFARX1 I_50788 (I866095,I2683,I865798,I865766,);
DFFARX1 I_50789 (I866078,I2683,I865798,I865787,);
nor I_50790 (I866140,I517389,I517377);
nor I_50791 (I865778,I865993,I866140);
or I_50792 (I866171,I517389,I517377);
nor I_50793 (I866188,I517368,I517371);
DFFARX1 I_50794 (I866188,I2683,I865798,I866214,);
not I_50795 (I866222,I866214);
nor I_50796 (I865784,I866222,I866027);
nand I_50797 (I866253,I866222,I865872);
not I_50798 (I866270,I517368);
nand I_50799 (I866287,I866270,I865976);
nand I_50800 (I866304,I866222,I866287);
nand I_50801 (I865775,I866304,I866253);
nand I_50802 (I865772,I866287,I866171);
not I_50803 (I866376,I2690);
DFFARX1 I_50804 (I84368,I2683,I866376,I866402,);
and I_50805 (I866410,I866402,I84344);
DFFARX1 I_50806 (I866410,I2683,I866376,I866359,);
DFFARX1 I_50807 (I84362,I2683,I866376,I866450,);
not I_50808 (I866458,I84350);
not I_50809 (I866475,I84347);
nand I_50810 (I866492,I866475,I866458);
nor I_50811 (I866347,I866450,I866492);
DFFARX1 I_50812 (I866492,I2683,I866376,I866532,);
not I_50813 (I866368,I866532);
not I_50814 (I866554,I84356);
nand I_50815 (I866571,I866475,I866554);
DFFARX1 I_50816 (I866571,I2683,I866376,I866597,);
not I_50817 (I866605,I866597);
not I_50818 (I866622,I84347);
nand I_50819 (I866639,I866622,I84365);
and I_50820 (I866656,I866458,I866639);
nor I_50821 (I866673,I866571,I866656);
DFFARX1 I_50822 (I866673,I2683,I866376,I866344,);
DFFARX1 I_50823 (I866656,I2683,I866376,I866365,);
nor I_50824 (I866718,I84347,I84359);
nor I_50825 (I866356,I866571,I866718);
or I_50826 (I866749,I84347,I84359);
nor I_50827 (I866766,I84353,I84344);
DFFARX1 I_50828 (I866766,I2683,I866376,I866792,);
not I_50829 (I866800,I866792);
nor I_50830 (I866362,I866800,I866605);
nand I_50831 (I866831,I866800,I866450);
not I_50832 (I866848,I84353);
nand I_50833 (I866865,I866848,I866554);
nand I_50834 (I866882,I866800,I866865);
nand I_50835 (I866353,I866882,I866831);
nand I_50836 (I866350,I866865,I866749);
not I_50837 (I866954,I2690);
DFFARX1 I_50838 (I238017,I2683,I866954,I866980,);
and I_50839 (I866988,I866980,I238002);
DFFARX1 I_50840 (I866988,I2683,I866954,I866937,);
DFFARX1 I_50841 (I238008,I2683,I866954,I867028,);
not I_50842 (I867036,I237990);
not I_50843 (I867053,I238011);
nand I_50844 (I867070,I867053,I867036);
nor I_50845 (I866925,I867028,I867070);
DFFARX1 I_50846 (I867070,I2683,I866954,I867110,);
not I_50847 (I866946,I867110);
not I_50848 (I867132,I238014);
nand I_50849 (I867149,I867053,I867132);
DFFARX1 I_50850 (I867149,I2683,I866954,I867175,);
not I_50851 (I867183,I867175);
not I_50852 (I867200,I238005);
nand I_50853 (I867217,I867200,I237993);
and I_50854 (I867234,I867036,I867217);
nor I_50855 (I867251,I867149,I867234);
DFFARX1 I_50856 (I867251,I2683,I866954,I866922,);
DFFARX1 I_50857 (I867234,I2683,I866954,I866943,);
nor I_50858 (I867296,I238005,I237999);
nor I_50859 (I866934,I867149,I867296);
or I_50860 (I867327,I238005,I237999);
nor I_50861 (I867344,I237996,I237990);
DFFARX1 I_50862 (I867344,I2683,I866954,I867370,);
not I_50863 (I867378,I867370);
nor I_50864 (I866940,I867378,I867183);
nand I_50865 (I867409,I867378,I867028);
not I_50866 (I867426,I237996);
nand I_50867 (I867443,I867426,I867132);
nand I_50868 (I867460,I867378,I867443);
nand I_50869 (I866931,I867460,I867409);
nand I_50870 (I866928,I867443,I867327);
not I_50871 (I867532,I2690);
DFFARX1 I_50872 (I1067396,I2683,I867532,I867558,);
and I_50873 (I867566,I867558,I1067378);
DFFARX1 I_50874 (I867566,I2683,I867532,I867515,);
DFFARX1 I_50875 (I1067369,I2683,I867532,I867606,);
not I_50876 (I867614,I1067384);
not I_50877 (I867631,I1067372);
nand I_50878 (I867648,I867631,I867614);
nor I_50879 (I867503,I867606,I867648);
DFFARX1 I_50880 (I867648,I2683,I867532,I867688,);
not I_50881 (I867524,I867688);
not I_50882 (I867710,I1067381);
nand I_50883 (I867727,I867631,I867710);
DFFARX1 I_50884 (I867727,I2683,I867532,I867753,);
not I_50885 (I867761,I867753);
not I_50886 (I867778,I1067390);
nand I_50887 (I867795,I867778,I1067369);
and I_50888 (I867812,I867614,I867795);
nor I_50889 (I867829,I867727,I867812);
DFFARX1 I_50890 (I867829,I2683,I867532,I867500,);
DFFARX1 I_50891 (I867812,I2683,I867532,I867521,);
nor I_50892 (I867874,I1067390,I1067393);
nor I_50893 (I867512,I867727,I867874);
or I_50894 (I867905,I1067390,I1067393);
nor I_50895 (I867922,I1067387,I1067375);
DFFARX1 I_50896 (I867922,I2683,I867532,I867948,);
not I_50897 (I867956,I867948);
nor I_50898 (I867518,I867956,I867761);
nand I_50899 (I867987,I867956,I867606);
not I_50900 (I868004,I1067387);
nand I_50901 (I868021,I868004,I867710);
nand I_50902 (I868038,I867956,I868021);
nand I_50903 (I867509,I868038,I867987);
nand I_50904 (I867506,I868021,I867905);
not I_50905 (I868110,I2690);
DFFARX1 I_50906 (I478657,I2683,I868110,I868136,);
and I_50907 (I868144,I868136,I478645);
DFFARX1 I_50908 (I868144,I2683,I868110,I868093,);
DFFARX1 I_50909 (I478660,I2683,I868110,I868184,);
not I_50910 (I868192,I478651);
not I_50911 (I868209,I478642);
nand I_50912 (I868226,I868209,I868192);
nor I_50913 (I868081,I868184,I868226);
DFFARX1 I_50914 (I868226,I2683,I868110,I868266,);
not I_50915 (I868102,I868266);
not I_50916 (I868288,I478648);
nand I_50917 (I868305,I868209,I868288);
DFFARX1 I_50918 (I868305,I2683,I868110,I868331,);
not I_50919 (I868339,I868331);
not I_50920 (I868356,I478663);
nand I_50921 (I868373,I868356,I478666);
and I_50922 (I868390,I868192,I868373);
nor I_50923 (I868407,I868305,I868390);
DFFARX1 I_50924 (I868407,I2683,I868110,I868078,);
DFFARX1 I_50925 (I868390,I2683,I868110,I868099,);
nor I_50926 (I868452,I478663,I478642);
nor I_50927 (I868090,I868305,I868452);
or I_50928 (I868483,I478663,I478642);
nor I_50929 (I868500,I478654,I478645);
DFFARX1 I_50930 (I868500,I2683,I868110,I868526,);
not I_50931 (I868534,I868526);
nor I_50932 (I868096,I868534,I868339);
nand I_50933 (I868565,I868534,I868184);
not I_50934 (I868582,I478654);
nand I_50935 (I868599,I868582,I868288);
nand I_50936 (I868616,I868534,I868599);
nand I_50937 (I868087,I868616,I868565);
nand I_50938 (I868084,I868599,I868483);
not I_50939 (I868688,I2690);
DFFARX1 I_50940 (I310216,I2683,I868688,I868714,);
and I_50941 (I868722,I868714,I310201);
DFFARX1 I_50942 (I868722,I2683,I868688,I868671,);
DFFARX1 I_50943 (I310207,I2683,I868688,I868762,);
not I_50944 (I868770,I310189);
not I_50945 (I868787,I310210);
nand I_50946 (I868804,I868787,I868770);
nor I_50947 (I868659,I868762,I868804);
DFFARX1 I_50948 (I868804,I2683,I868688,I868844,);
not I_50949 (I868680,I868844);
not I_50950 (I868866,I310213);
nand I_50951 (I868883,I868787,I868866);
DFFARX1 I_50952 (I868883,I2683,I868688,I868909,);
not I_50953 (I868917,I868909);
not I_50954 (I868934,I310204);
nand I_50955 (I868951,I868934,I310192);
and I_50956 (I868968,I868770,I868951);
nor I_50957 (I868985,I868883,I868968);
DFFARX1 I_50958 (I868985,I2683,I868688,I868656,);
DFFARX1 I_50959 (I868968,I2683,I868688,I868677,);
nor I_50960 (I869030,I310204,I310198);
nor I_50961 (I868668,I868883,I869030);
or I_50962 (I869061,I310204,I310198);
nor I_50963 (I869078,I310195,I310189);
DFFARX1 I_50964 (I869078,I2683,I868688,I869104,);
not I_50965 (I869112,I869104);
nor I_50966 (I868674,I869112,I868917);
nand I_50967 (I869143,I869112,I868762);
not I_50968 (I869160,I310195);
nand I_50969 (I869177,I869160,I868866);
nand I_50970 (I869194,I869112,I869177);
nand I_50971 (I868665,I869194,I869143);
nand I_50972 (I868662,I869177,I869061);
not I_50973 (I869266,I2690);
DFFARX1 I_50974 (I414555,I2683,I869266,I869292,);
and I_50975 (I869300,I869292,I414570);
DFFARX1 I_50976 (I869300,I2683,I869266,I869249,);
DFFARX1 I_50977 (I414561,I2683,I869266,I869340,);
not I_50978 (I869348,I414555);
not I_50979 (I869365,I414573);
nand I_50980 (I869382,I869365,I869348);
nor I_50981 (I869237,I869340,I869382);
DFFARX1 I_50982 (I869382,I2683,I869266,I869422,);
not I_50983 (I869258,I869422);
not I_50984 (I869444,I414564);
nand I_50985 (I869461,I869365,I869444);
DFFARX1 I_50986 (I869461,I2683,I869266,I869487,);
not I_50987 (I869495,I869487);
not I_50988 (I869512,I414576);
nand I_50989 (I869529,I869512,I414552);
and I_50990 (I869546,I869348,I869529);
nor I_50991 (I869563,I869461,I869546);
DFFARX1 I_50992 (I869563,I2683,I869266,I869234,);
DFFARX1 I_50993 (I869546,I2683,I869266,I869255,);
nor I_50994 (I869608,I414576,I414552);
nor I_50995 (I869246,I869461,I869608);
or I_50996 (I869639,I414576,I414552);
nor I_50997 (I869656,I414558,I414567);
DFFARX1 I_50998 (I869656,I2683,I869266,I869682,);
not I_50999 (I869690,I869682);
nor I_51000 (I869252,I869690,I869495);
nand I_51001 (I869721,I869690,I869340);
not I_51002 (I869738,I414558);
nand I_51003 (I869755,I869738,I869444);
nand I_51004 (I869772,I869690,I869755);
nand I_51005 (I869243,I869772,I869721);
nand I_51006 (I869240,I869755,I869639);
not I_51007 (I869844,I2690);
DFFARX1 I_51008 (I768447,I2683,I869844,I869870,);
and I_51009 (I869878,I869870,I768441);
DFFARX1 I_51010 (I869878,I2683,I869844,I869827,);
DFFARX1 I_51011 (I768459,I2683,I869844,I869918,);
not I_51012 (I869926,I768450);
not I_51013 (I869943,I768462);
nand I_51014 (I869960,I869943,I869926);
nor I_51015 (I869815,I869918,I869960);
DFFARX1 I_51016 (I869960,I2683,I869844,I870000,);
not I_51017 (I869836,I870000);
not I_51018 (I870022,I768468);
nand I_51019 (I870039,I869943,I870022);
DFFARX1 I_51020 (I870039,I2683,I869844,I870065,);
not I_51021 (I870073,I870065);
not I_51022 (I870090,I768444);
nand I_51023 (I870107,I870090,I768465);
and I_51024 (I870124,I869926,I870107);
nor I_51025 (I870141,I870039,I870124);
DFFARX1 I_51026 (I870141,I2683,I869844,I869812,);
DFFARX1 I_51027 (I870124,I2683,I869844,I869833,);
nor I_51028 (I870186,I768444,I768456);
nor I_51029 (I869824,I870039,I870186);
or I_51030 (I870217,I768444,I768456);
nor I_51031 (I870234,I768441,I768453);
DFFARX1 I_51032 (I870234,I2683,I869844,I870260,);
not I_51033 (I870268,I870260);
nor I_51034 (I869830,I870268,I870073);
nand I_51035 (I870299,I870268,I869918);
not I_51036 (I870316,I768441);
nand I_51037 (I870333,I870316,I870022);
nand I_51038 (I870350,I870268,I870333);
nand I_51039 (I869821,I870350,I870299);
nand I_51040 (I869818,I870333,I870217);
not I_51041 (I870422,I2690);
DFFARX1 I_51042 (I769739,I2683,I870422,I870448,);
and I_51043 (I870456,I870448,I769733);
DFFARX1 I_51044 (I870456,I2683,I870422,I870405,);
DFFARX1 I_51045 (I769751,I2683,I870422,I870496,);
not I_51046 (I870504,I769742);
not I_51047 (I870521,I769754);
nand I_51048 (I870538,I870521,I870504);
nor I_51049 (I870393,I870496,I870538);
DFFARX1 I_51050 (I870538,I2683,I870422,I870578,);
not I_51051 (I870414,I870578);
not I_51052 (I870600,I769760);
nand I_51053 (I870617,I870521,I870600);
DFFARX1 I_51054 (I870617,I2683,I870422,I870643,);
not I_51055 (I870651,I870643);
not I_51056 (I870668,I769736);
nand I_51057 (I870685,I870668,I769757);
and I_51058 (I870702,I870504,I870685);
nor I_51059 (I870719,I870617,I870702);
DFFARX1 I_51060 (I870719,I2683,I870422,I870390,);
DFFARX1 I_51061 (I870702,I2683,I870422,I870411,);
nor I_51062 (I870764,I769736,I769748);
nor I_51063 (I870402,I870617,I870764);
or I_51064 (I870795,I769736,I769748);
nor I_51065 (I870812,I769733,I769745);
DFFARX1 I_51066 (I870812,I2683,I870422,I870838,);
not I_51067 (I870846,I870838);
nor I_51068 (I870408,I870846,I870651);
nand I_51069 (I870877,I870846,I870496);
not I_51070 (I870894,I769733);
nand I_51071 (I870911,I870894,I870600);
nand I_51072 (I870928,I870846,I870911);
nand I_51073 (I870399,I870928,I870877);
nand I_51074 (I870396,I870911,I870795);
not I_51075 (I871000,I2690);
DFFARX1 I_51076 (I469409,I2683,I871000,I871026,);
and I_51077 (I871034,I871026,I469397);
DFFARX1 I_51078 (I871034,I2683,I871000,I870983,);
DFFARX1 I_51079 (I469412,I2683,I871000,I871074,);
not I_51080 (I871082,I469403);
not I_51081 (I871099,I469394);
nand I_51082 (I871116,I871099,I871082);
nor I_51083 (I870971,I871074,I871116);
DFFARX1 I_51084 (I871116,I2683,I871000,I871156,);
not I_51085 (I870992,I871156);
not I_51086 (I871178,I469400);
nand I_51087 (I871195,I871099,I871178);
DFFARX1 I_51088 (I871195,I2683,I871000,I871221,);
not I_51089 (I871229,I871221);
not I_51090 (I871246,I469415);
nand I_51091 (I871263,I871246,I469418);
and I_51092 (I871280,I871082,I871263);
nor I_51093 (I871297,I871195,I871280);
DFFARX1 I_51094 (I871297,I2683,I871000,I870968,);
DFFARX1 I_51095 (I871280,I2683,I871000,I870989,);
nor I_51096 (I871342,I469415,I469394);
nor I_51097 (I870980,I871195,I871342);
or I_51098 (I871373,I469415,I469394);
nor I_51099 (I871390,I469406,I469397);
DFFARX1 I_51100 (I871390,I2683,I871000,I871416,);
not I_51101 (I871424,I871416);
nor I_51102 (I870986,I871424,I871229);
nand I_51103 (I871455,I871424,I871074);
not I_51104 (I871472,I469406);
nand I_51105 (I871489,I871472,I871178);
nand I_51106 (I871506,I871424,I871489);
nand I_51107 (I870977,I871506,I871455);
nand I_51108 (I870974,I871489,I871373);
not I_51109 (I871578,I2690);
DFFARX1 I_51110 (I254354,I2683,I871578,I871604,);
and I_51111 (I871612,I871604,I254339);
DFFARX1 I_51112 (I871612,I2683,I871578,I871561,);
DFFARX1 I_51113 (I254345,I2683,I871578,I871652,);
not I_51114 (I871660,I254327);
not I_51115 (I871677,I254348);
nand I_51116 (I871694,I871677,I871660);
nor I_51117 (I871549,I871652,I871694);
DFFARX1 I_51118 (I871694,I2683,I871578,I871734,);
not I_51119 (I871570,I871734);
not I_51120 (I871756,I254351);
nand I_51121 (I871773,I871677,I871756);
DFFARX1 I_51122 (I871773,I2683,I871578,I871799,);
not I_51123 (I871807,I871799);
not I_51124 (I871824,I254342);
nand I_51125 (I871841,I871824,I254330);
and I_51126 (I871858,I871660,I871841);
nor I_51127 (I871875,I871773,I871858);
DFFARX1 I_51128 (I871875,I2683,I871578,I871546,);
DFFARX1 I_51129 (I871858,I2683,I871578,I871567,);
nor I_51130 (I871920,I254342,I254336);
nor I_51131 (I871558,I871773,I871920);
or I_51132 (I871951,I254342,I254336);
nor I_51133 (I871968,I254333,I254327);
DFFARX1 I_51134 (I871968,I2683,I871578,I871994,);
not I_51135 (I872002,I871994);
nor I_51136 (I871564,I872002,I871807);
nand I_51137 (I872033,I872002,I871652);
not I_51138 (I872050,I254333);
nand I_51139 (I872067,I872050,I871756);
nand I_51140 (I872084,I872002,I872067);
nand I_51141 (I871555,I872084,I872033);
nand I_51142 (I871552,I872067,I871951);
not I_51143 (I872156,I2690);
DFFARX1 I_51144 (I224842,I2683,I872156,I872182,);
and I_51145 (I872190,I872182,I224827);
DFFARX1 I_51146 (I872190,I2683,I872156,I872139,);
DFFARX1 I_51147 (I224833,I2683,I872156,I872230,);
not I_51148 (I872238,I224815);
not I_51149 (I872255,I224836);
nand I_51150 (I872272,I872255,I872238);
nor I_51151 (I872127,I872230,I872272);
DFFARX1 I_51152 (I872272,I2683,I872156,I872312,);
not I_51153 (I872148,I872312);
not I_51154 (I872334,I224839);
nand I_51155 (I872351,I872255,I872334);
DFFARX1 I_51156 (I872351,I2683,I872156,I872377,);
not I_51157 (I872385,I872377);
not I_51158 (I872402,I224830);
nand I_51159 (I872419,I872402,I224818);
and I_51160 (I872436,I872238,I872419);
nor I_51161 (I872453,I872351,I872436);
DFFARX1 I_51162 (I872453,I2683,I872156,I872124,);
DFFARX1 I_51163 (I872436,I2683,I872156,I872145,);
nor I_51164 (I872498,I224830,I224824);
nor I_51165 (I872136,I872351,I872498);
or I_51166 (I872529,I224830,I224824);
nor I_51167 (I872546,I224821,I224815);
DFFARX1 I_51168 (I872546,I2683,I872156,I872572,);
not I_51169 (I872580,I872572);
nor I_51170 (I872142,I872580,I872385);
nand I_51171 (I872611,I872580,I872230);
not I_51172 (I872628,I224821);
nand I_51173 (I872645,I872628,I872334);
nand I_51174 (I872662,I872580,I872645);
nand I_51175 (I872133,I872662,I872611);
nand I_51176 (I872130,I872645,I872529);
not I_51177 (I872734,I2690);
DFFARX1 I_51178 (I78044,I2683,I872734,I872760,);
and I_51179 (I872768,I872760,I78020);
DFFARX1 I_51180 (I872768,I2683,I872734,I872717,);
DFFARX1 I_51181 (I78038,I2683,I872734,I872808,);
not I_51182 (I872816,I78026);
not I_51183 (I872833,I78023);
nand I_51184 (I872850,I872833,I872816);
nor I_51185 (I872705,I872808,I872850);
DFFARX1 I_51186 (I872850,I2683,I872734,I872890,);
not I_51187 (I872726,I872890);
not I_51188 (I872912,I78032);
nand I_51189 (I872929,I872833,I872912);
DFFARX1 I_51190 (I872929,I2683,I872734,I872955,);
not I_51191 (I872963,I872955);
not I_51192 (I872980,I78023);
nand I_51193 (I872997,I872980,I78041);
and I_51194 (I873014,I872816,I872997);
nor I_51195 (I873031,I872929,I873014);
DFFARX1 I_51196 (I873031,I2683,I872734,I872702,);
DFFARX1 I_51197 (I873014,I2683,I872734,I872723,);
nor I_51198 (I873076,I78023,I78035);
nor I_51199 (I872714,I872929,I873076);
or I_51200 (I873107,I78023,I78035);
nor I_51201 (I873124,I78029,I78020);
DFFARX1 I_51202 (I873124,I2683,I872734,I873150,);
not I_51203 (I873158,I873150);
nor I_51204 (I872720,I873158,I872963);
nand I_51205 (I873189,I873158,I872808);
not I_51206 (I873206,I78029);
nand I_51207 (I873223,I873206,I872912);
nand I_51208 (I873240,I873158,I873223);
nand I_51209 (I872711,I873240,I873189);
nand I_51210 (I872708,I873223,I873107);
not I_51211 (I873312,I2690);
DFFARX1 I_51212 (I628058,I2683,I873312,I873338,);
and I_51213 (I873346,I873338,I628064);
DFFARX1 I_51214 (I873346,I2683,I873312,I873295,);
DFFARX1 I_51215 (I628070,I2683,I873312,I873386,);
not I_51216 (I873394,I628055);
not I_51217 (I873411,I628055);
nand I_51218 (I873428,I873411,I873394);
nor I_51219 (I873283,I873386,I873428);
DFFARX1 I_51220 (I873428,I2683,I873312,I873468,);
not I_51221 (I873304,I873468);
not I_51222 (I873490,I628073);
nand I_51223 (I873507,I873411,I873490);
DFFARX1 I_51224 (I873507,I2683,I873312,I873533,);
not I_51225 (I873541,I873533);
not I_51226 (I873558,I628067);
nand I_51227 (I873575,I873558,I628058);
and I_51228 (I873592,I873394,I873575);
nor I_51229 (I873609,I873507,I873592);
DFFARX1 I_51230 (I873609,I2683,I873312,I873280,);
DFFARX1 I_51231 (I873592,I2683,I873312,I873301,);
nor I_51232 (I873654,I628067,I628076);
nor I_51233 (I873292,I873507,I873654);
or I_51234 (I873685,I628067,I628076);
nor I_51235 (I873702,I628061,I628061);
DFFARX1 I_51236 (I873702,I2683,I873312,I873728,);
not I_51237 (I873736,I873728);
nor I_51238 (I873298,I873736,I873541);
nand I_51239 (I873767,I873736,I873386);
not I_51240 (I873784,I628061);
nand I_51241 (I873801,I873784,I873490);
nand I_51242 (I873818,I873736,I873801);
nand I_51243 (I873289,I873818,I873767);
nand I_51244 (I873286,I873801,I873685);
not I_51245 (I873890,I2690);
DFFARX1 I_51246 (I277015,I2683,I873890,I873916,);
and I_51247 (I873924,I873916,I277000);
DFFARX1 I_51248 (I873924,I2683,I873890,I873873,);
DFFARX1 I_51249 (I277006,I2683,I873890,I873964,);
not I_51250 (I873972,I276988);
not I_51251 (I873989,I277009);
nand I_51252 (I874006,I873989,I873972);
nor I_51253 (I873861,I873964,I874006);
DFFARX1 I_51254 (I874006,I2683,I873890,I874046,);
not I_51255 (I873882,I874046);
not I_51256 (I874068,I277012);
nand I_51257 (I874085,I873989,I874068);
DFFARX1 I_51258 (I874085,I2683,I873890,I874111,);
not I_51259 (I874119,I874111);
not I_51260 (I874136,I277003);
nand I_51261 (I874153,I874136,I276991);
and I_51262 (I874170,I873972,I874153);
nor I_51263 (I874187,I874085,I874170);
DFFARX1 I_51264 (I874187,I2683,I873890,I873858,);
DFFARX1 I_51265 (I874170,I2683,I873890,I873879,);
nor I_51266 (I874232,I277003,I276997);
nor I_51267 (I873870,I874085,I874232);
or I_51268 (I874263,I277003,I276997);
nor I_51269 (I874280,I276994,I276988);
DFFARX1 I_51270 (I874280,I2683,I873890,I874306,);
not I_51271 (I874314,I874306);
nor I_51272 (I873876,I874314,I874119);
nand I_51273 (I874345,I874314,I873964);
not I_51274 (I874362,I276994);
nand I_51275 (I874379,I874362,I874068);
nand I_51276 (I874396,I874314,I874379);
nand I_51277 (I873867,I874396,I874345);
nand I_51278 (I873864,I874379,I874263);
not I_51279 (I874468,I2690);
DFFARX1 I_51280 (I287555,I2683,I874468,I874494,);
and I_51281 (I874502,I874494,I287540);
DFFARX1 I_51282 (I874502,I2683,I874468,I874451,);
DFFARX1 I_51283 (I287546,I2683,I874468,I874542,);
not I_51284 (I874550,I287528);
not I_51285 (I874567,I287549);
nand I_51286 (I874584,I874567,I874550);
nor I_51287 (I874439,I874542,I874584);
DFFARX1 I_51288 (I874584,I2683,I874468,I874624,);
not I_51289 (I874460,I874624);
not I_51290 (I874646,I287552);
nand I_51291 (I874663,I874567,I874646);
DFFARX1 I_51292 (I874663,I2683,I874468,I874689,);
not I_51293 (I874697,I874689);
not I_51294 (I874714,I287543);
nand I_51295 (I874731,I874714,I287531);
and I_51296 (I874748,I874550,I874731);
nor I_51297 (I874765,I874663,I874748);
DFFARX1 I_51298 (I874765,I2683,I874468,I874436,);
DFFARX1 I_51299 (I874748,I2683,I874468,I874457,);
nor I_51300 (I874810,I287543,I287537);
nor I_51301 (I874448,I874663,I874810);
or I_51302 (I874841,I287543,I287537);
nor I_51303 (I874858,I287534,I287528);
DFFARX1 I_51304 (I874858,I2683,I874468,I874884,);
not I_51305 (I874892,I874884);
nor I_51306 (I874454,I874892,I874697);
nand I_51307 (I874923,I874892,I874542);
not I_51308 (I874940,I287534);
nand I_51309 (I874957,I874940,I874646);
nand I_51310 (I874974,I874892,I874957);
nand I_51311 (I874445,I874974,I874923);
nand I_51312 (I874442,I874957,I874841);
not I_51313 (I875046,I2690);
DFFARX1 I_51314 (I999580,I2683,I875046,I875072,);
and I_51315 (I875080,I875072,I999562);
DFFARX1 I_51316 (I875080,I2683,I875046,I875029,);
DFFARX1 I_51317 (I999571,I2683,I875046,I875120,);
not I_51318 (I875128,I999556);
not I_51319 (I875145,I999568);
nand I_51320 (I875162,I875145,I875128);
nor I_51321 (I875017,I875120,I875162);
DFFARX1 I_51322 (I875162,I2683,I875046,I875202,);
not I_51323 (I875038,I875202);
not I_51324 (I875224,I999559);
nand I_51325 (I875241,I875145,I875224);
DFFARX1 I_51326 (I875241,I2683,I875046,I875267,);
not I_51327 (I875275,I875267);
not I_51328 (I875292,I999556);
nand I_51329 (I875309,I875292,I999559);
and I_51330 (I875326,I875128,I875309);
nor I_51331 (I875343,I875241,I875326);
DFFARX1 I_51332 (I875343,I2683,I875046,I875014,);
DFFARX1 I_51333 (I875326,I2683,I875046,I875035,);
nor I_51334 (I875388,I999556,I999577);
nor I_51335 (I875026,I875241,I875388);
or I_51336 (I875419,I999556,I999577);
nor I_51337 (I875436,I999565,I999574);
DFFARX1 I_51338 (I875436,I2683,I875046,I875462,);
not I_51339 (I875470,I875462);
nor I_51340 (I875032,I875470,I875275);
nand I_51341 (I875501,I875470,I875120);
not I_51342 (I875518,I999565);
nand I_51343 (I875535,I875518,I875224);
nand I_51344 (I875552,I875470,I875535);
nand I_51345 (I875023,I875552,I875501);
nand I_51346 (I875020,I875535,I875419);
not I_51347 (I875624,I2690);
DFFARX1 I_51348 (I124770,I2683,I875624,I875650,);
and I_51349 (I875658,I875650,I124773);
DFFARX1 I_51350 (I875658,I2683,I875624,I875607,);
DFFARX1 I_51351 (I124773,I2683,I875624,I875698,);
not I_51352 (I875706,I124788);
not I_51353 (I875723,I124794);
nand I_51354 (I875740,I875723,I875706);
nor I_51355 (I875595,I875698,I875740);
DFFARX1 I_51356 (I875740,I2683,I875624,I875780,);
not I_51357 (I875616,I875780);
not I_51358 (I875802,I124782);
nand I_51359 (I875819,I875723,I875802);
DFFARX1 I_51360 (I875819,I2683,I875624,I875845,);
not I_51361 (I875853,I875845);
not I_51362 (I875870,I124779);
nand I_51363 (I875887,I875870,I124776);
and I_51364 (I875904,I875706,I875887);
nor I_51365 (I875921,I875819,I875904);
DFFARX1 I_51366 (I875921,I2683,I875624,I875592,);
DFFARX1 I_51367 (I875904,I2683,I875624,I875613,);
nor I_51368 (I875966,I124779,I124770);
nor I_51369 (I875604,I875819,I875966);
or I_51370 (I875997,I124779,I124770);
nor I_51371 (I876014,I124785,I124791);
DFFARX1 I_51372 (I876014,I2683,I875624,I876040,);
not I_51373 (I876048,I876040);
nor I_51374 (I875610,I876048,I875853);
nand I_51375 (I876079,I876048,I875698);
not I_51376 (I876096,I124785);
nand I_51377 (I876113,I876096,I875802);
nand I_51378 (I876130,I876048,I876113);
nand I_51379 (I875601,I876130,I876079);
nand I_51380 (I875598,I876113,I875997);
not I_51381 (I876202,I2690);
DFFARX1 I_51382 (I271218,I2683,I876202,I876228,);
and I_51383 (I876236,I876228,I271203);
DFFARX1 I_51384 (I876236,I2683,I876202,I876185,);
DFFARX1 I_51385 (I271209,I2683,I876202,I876276,);
not I_51386 (I876284,I271191);
not I_51387 (I876301,I271212);
nand I_51388 (I876318,I876301,I876284);
nor I_51389 (I876173,I876276,I876318);
DFFARX1 I_51390 (I876318,I2683,I876202,I876358,);
not I_51391 (I876194,I876358);
not I_51392 (I876380,I271215);
nand I_51393 (I876397,I876301,I876380);
DFFARX1 I_51394 (I876397,I2683,I876202,I876423,);
not I_51395 (I876431,I876423);
not I_51396 (I876448,I271206);
nand I_51397 (I876465,I876448,I271194);
and I_51398 (I876482,I876284,I876465);
nor I_51399 (I876499,I876397,I876482);
DFFARX1 I_51400 (I876499,I2683,I876202,I876170,);
DFFARX1 I_51401 (I876482,I2683,I876202,I876191,);
nor I_51402 (I876544,I271206,I271200);
nor I_51403 (I876182,I876397,I876544);
or I_51404 (I876575,I271206,I271200);
nor I_51405 (I876592,I271197,I271191);
DFFARX1 I_51406 (I876592,I2683,I876202,I876618,);
not I_51407 (I876626,I876618);
nor I_51408 (I876188,I876626,I876431);
nand I_51409 (I876657,I876626,I876276);
not I_51410 (I876674,I271197);
nand I_51411 (I876691,I876674,I876380);
nand I_51412 (I876708,I876626,I876691);
nand I_51413 (I876179,I876708,I876657);
nand I_51414 (I876176,I876691,I876575);
not I_51415 (I876780,I2690);
DFFARX1 I_51416 (I304419,I2683,I876780,I876806,);
and I_51417 (I876814,I876806,I304404);
DFFARX1 I_51418 (I876814,I2683,I876780,I876763,);
DFFARX1 I_51419 (I304410,I2683,I876780,I876854,);
not I_51420 (I876862,I304392);
not I_51421 (I876879,I304413);
nand I_51422 (I876896,I876879,I876862);
nor I_51423 (I876751,I876854,I876896);
DFFARX1 I_51424 (I876896,I2683,I876780,I876936,);
not I_51425 (I876772,I876936);
not I_51426 (I876958,I304416);
nand I_51427 (I876975,I876879,I876958);
DFFARX1 I_51428 (I876975,I2683,I876780,I877001,);
not I_51429 (I877009,I877001);
not I_51430 (I877026,I304407);
nand I_51431 (I877043,I877026,I304395);
and I_51432 (I877060,I876862,I877043);
nor I_51433 (I877077,I876975,I877060);
DFFARX1 I_51434 (I877077,I2683,I876780,I876748,);
DFFARX1 I_51435 (I877060,I2683,I876780,I876769,);
nor I_51436 (I877122,I304407,I304401);
nor I_51437 (I876760,I876975,I877122);
or I_51438 (I877153,I304407,I304401);
nor I_51439 (I877170,I304398,I304392);
DFFARX1 I_51440 (I877170,I2683,I876780,I877196,);
not I_51441 (I877204,I877196);
nor I_51442 (I876766,I877204,I877009);
nand I_51443 (I877235,I877204,I876854);
not I_51444 (I877252,I304398);
nand I_51445 (I877269,I877252,I876958);
nand I_51446 (I877286,I877204,I877269);
nand I_51447 (I876757,I877286,I877235);
nand I_51448 (I876754,I877269,I877153);
not I_51449 (I877358,I2690);
DFFARX1 I_51450 (I329586,I2683,I877358,I877384,);
and I_51451 (I877392,I877384,I329601);
DFFARX1 I_51452 (I877392,I2683,I877358,I877341,);
DFFARX1 I_51453 (I329604,I2683,I877358,I877432,);
not I_51454 (I877440,I329598);
not I_51455 (I877457,I329613);
nand I_51456 (I877474,I877457,I877440);
nor I_51457 (I877329,I877432,I877474);
DFFARX1 I_51458 (I877474,I2683,I877358,I877514,);
not I_51459 (I877350,I877514);
not I_51460 (I877536,I329589);
nand I_51461 (I877553,I877457,I877536);
DFFARX1 I_51462 (I877553,I2683,I877358,I877579,);
not I_51463 (I877587,I877579);
not I_51464 (I877604,I329592);
nand I_51465 (I877621,I877604,I329586);
and I_51466 (I877638,I877440,I877621);
nor I_51467 (I877655,I877553,I877638);
DFFARX1 I_51468 (I877655,I2683,I877358,I877326,);
DFFARX1 I_51469 (I877638,I2683,I877358,I877347,);
nor I_51470 (I877700,I329592,I329595);
nor I_51471 (I877338,I877553,I877700);
or I_51472 (I877731,I329592,I329595);
nor I_51473 (I877748,I329610,I329607);
DFFARX1 I_51474 (I877748,I2683,I877358,I877774,);
not I_51475 (I877782,I877774);
nor I_51476 (I877344,I877782,I877587);
nand I_51477 (I877813,I877782,I877432);
not I_51478 (I877830,I329610);
nand I_51479 (I877847,I877830,I877536);
nand I_51480 (I877864,I877782,I877847);
nand I_51481 (I877335,I877864,I877813);
nand I_51482 (I877332,I877847,I877731);
not I_51483 (I877936,I2690);
DFFARX1 I_51484 (I1016342,I2683,I877936,I877962,);
and I_51485 (I877970,I877962,I1016324);
DFFARX1 I_51486 (I877970,I2683,I877936,I877919,);
DFFARX1 I_51487 (I1016333,I2683,I877936,I878010,);
not I_51488 (I878018,I1016318);
not I_51489 (I878035,I1016330);
nand I_51490 (I878052,I878035,I878018);
nor I_51491 (I877907,I878010,I878052);
DFFARX1 I_51492 (I878052,I2683,I877936,I878092,);
not I_51493 (I877928,I878092);
not I_51494 (I878114,I1016321);
nand I_51495 (I878131,I878035,I878114);
DFFARX1 I_51496 (I878131,I2683,I877936,I878157,);
not I_51497 (I878165,I878157);
not I_51498 (I878182,I1016318);
nand I_51499 (I878199,I878182,I1016321);
and I_51500 (I878216,I878018,I878199);
nor I_51501 (I878233,I878131,I878216);
DFFARX1 I_51502 (I878233,I2683,I877936,I877904,);
DFFARX1 I_51503 (I878216,I2683,I877936,I877925,);
nor I_51504 (I878278,I1016318,I1016339);
nor I_51505 (I877916,I878131,I878278);
or I_51506 (I878309,I1016318,I1016339);
nor I_51507 (I878326,I1016327,I1016336);
DFFARX1 I_51508 (I878326,I2683,I877936,I878352,);
not I_51509 (I878360,I878352);
nor I_51510 (I877922,I878360,I878165);
nand I_51511 (I878391,I878360,I878010);
not I_51512 (I878408,I1016327);
nand I_51513 (I878425,I878408,I878114);
nand I_51514 (I878442,I878360,I878425);
nand I_51515 (I877913,I878442,I878391);
nand I_51516 (I877910,I878425,I878309);
not I_51517 (I878514,I2690);
DFFARX1 I_51518 (I168205,I2683,I878514,I878540,);
and I_51519 (I878548,I878540,I168208);
DFFARX1 I_51520 (I878548,I2683,I878514,I878497,);
DFFARX1 I_51521 (I168208,I2683,I878514,I878588,);
not I_51522 (I878596,I168223);
not I_51523 (I878613,I168229);
nand I_51524 (I878630,I878613,I878596);
nor I_51525 (I878485,I878588,I878630);
DFFARX1 I_51526 (I878630,I2683,I878514,I878670,);
not I_51527 (I878506,I878670);
not I_51528 (I878692,I168217);
nand I_51529 (I878709,I878613,I878692);
DFFARX1 I_51530 (I878709,I2683,I878514,I878735,);
not I_51531 (I878743,I878735);
not I_51532 (I878760,I168214);
nand I_51533 (I878777,I878760,I168211);
and I_51534 (I878794,I878596,I878777);
nor I_51535 (I878811,I878709,I878794);
DFFARX1 I_51536 (I878811,I2683,I878514,I878482,);
DFFARX1 I_51537 (I878794,I2683,I878514,I878503,);
nor I_51538 (I878856,I168214,I168205);
nor I_51539 (I878494,I878709,I878856);
or I_51540 (I878887,I168214,I168205);
nor I_51541 (I878904,I168220,I168226);
DFFARX1 I_51542 (I878904,I2683,I878514,I878930,);
not I_51543 (I878938,I878930);
nor I_51544 (I878500,I878938,I878743);
nand I_51545 (I878969,I878938,I878588);
not I_51546 (I878986,I168220);
nand I_51547 (I879003,I878986,I878692);
nand I_51548 (I879020,I878938,I879003);
nand I_51549 (I878491,I879020,I878969);
nand I_51550 (I878488,I879003,I878887);
not I_51551 (I879092,I2690);
DFFARX1 I_51552 (I638071,I2683,I879092,I879118,);
and I_51553 (I879126,I879118,I638077);
DFFARX1 I_51554 (I879126,I2683,I879092,I879075,);
DFFARX1 I_51555 (I638083,I2683,I879092,I879166,);
not I_51556 (I879174,I638068);
not I_51557 (I879191,I638068);
nand I_51558 (I879208,I879191,I879174);
nor I_51559 (I879063,I879166,I879208);
DFFARX1 I_51560 (I879208,I2683,I879092,I879248,);
not I_51561 (I879084,I879248);
not I_51562 (I879270,I638086);
nand I_51563 (I879287,I879191,I879270);
DFFARX1 I_51564 (I879287,I2683,I879092,I879313,);
not I_51565 (I879321,I879313);
not I_51566 (I879338,I638080);
nand I_51567 (I879355,I879338,I638071);
and I_51568 (I879372,I879174,I879355);
nor I_51569 (I879389,I879287,I879372);
DFFARX1 I_51570 (I879389,I2683,I879092,I879060,);
DFFARX1 I_51571 (I879372,I2683,I879092,I879081,);
nor I_51572 (I879434,I638080,I638089);
nor I_51573 (I879072,I879287,I879434);
or I_51574 (I879465,I638080,I638089);
nor I_51575 (I879482,I638074,I638074);
DFFARX1 I_51576 (I879482,I2683,I879092,I879508,);
not I_51577 (I879516,I879508);
nor I_51578 (I879078,I879516,I879321);
nand I_51579 (I879547,I879516,I879166);
not I_51580 (I879564,I638074);
nand I_51581 (I879581,I879564,I879270);
nand I_51582 (I879598,I879516,I879581);
nand I_51583 (I879069,I879598,I879547);
nand I_51584 (I879066,I879581,I879465);
not I_51585 (I879670,I2690);
DFFARX1 I_51586 (I68031,I2683,I879670,I879696,);
and I_51587 (I879704,I879696,I68007);
DFFARX1 I_51588 (I879704,I2683,I879670,I879653,);
DFFARX1 I_51589 (I68025,I2683,I879670,I879744,);
not I_51590 (I879752,I68013);
not I_51591 (I879769,I68010);
nand I_51592 (I879786,I879769,I879752);
nor I_51593 (I879641,I879744,I879786);
DFFARX1 I_51594 (I879786,I2683,I879670,I879826,);
not I_51595 (I879662,I879826);
not I_51596 (I879848,I68019);
nand I_51597 (I879865,I879769,I879848);
DFFARX1 I_51598 (I879865,I2683,I879670,I879891,);
not I_51599 (I879899,I879891);
not I_51600 (I879916,I68010);
nand I_51601 (I879933,I879916,I68028);
and I_51602 (I879950,I879752,I879933);
nor I_51603 (I879967,I879865,I879950);
DFFARX1 I_51604 (I879967,I2683,I879670,I879638,);
DFFARX1 I_51605 (I879950,I2683,I879670,I879659,);
nor I_51606 (I880012,I68010,I68022);
nor I_51607 (I879650,I879865,I880012);
or I_51608 (I880043,I68010,I68022);
nor I_51609 (I880060,I68016,I68007);
DFFARX1 I_51610 (I880060,I2683,I879670,I880086,);
not I_51611 (I880094,I880086);
nor I_51612 (I879656,I880094,I879899);
nand I_51613 (I880125,I880094,I879744);
not I_51614 (I880142,I68016);
nand I_51615 (I880159,I880142,I879848);
nand I_51616 (I880176,I880094,I880159);
nand I_51617 (I879647,I880176,I880125);
nand I_51618 (I879644,I880159,I880043);
not I_51619 (I880248,I2690);
DFFARX1 I_51620 (I591945,I2683,I880248,I880274,);
and I_51621 (I880282,I880274,I591933);
DFFARX1 I_51622 (I880282,I2683,I880248,I880231,);
DFFARX1 I_51623 (I591936,I2683,I880248,I880322,);
not I_51624 (I880330,I591930);
not I_51625 (I880347,I591954);
nand I_51626 (I880364,I880347,I880330);
nor I_51627 (I880219,I880322,I880364);
DFFARX1 I_51628 (I880364,I2683,I880248,I880404,);
not I_51629 (I880240,I880404);
not I_51630 (I880426,I591942);
nand I_51631 (I880443,I880347,I880426);
DFFARX1 I_51632 (I880443,I2683,I880248,I880469,);
not I_51633 (I880477,I880469);
not I_51634 (I880494,I591951);
nand I_51635 (I880511,I880494,I591948);
and I_51636 (I880528,I880330,I880511);
nor I_51637 (I880545,I880443,I880528);
DFFARX1 I_51638 (I880545,I2683,I880248,I880216,);
DFFARX1 I_51639 (I880528,I2683,I880248,I880237,);
nor I_51640 (I880590,I591951,I591939);
nor I_51641 (I880228,I880443,I880590);
or I_51642 (I880621,I591951,I591939);
nor I_51643 (I880638,I591930,I591933);
DFFARX1 I_51644 (I880638,I2683,I880248,I880664,);
not I_51645 (I880672,I880664);
nor I_51646 (I880234,I880672,I880477);
nand I_51647 (I880703,I880672,I880322);
not I_51648 (I880720,I591930);
nand I_51649 (I880737,I880720,I880426);
nand I_51650 (I880754,I880672,I880737);
nand I_51651 (I880225,I880754,I880703);
nand I_51652 (I880222,I880737,I880621);
not I_51653 (I880826,I2690);
DFFARX1 I_51654 (I478079,I2683,I880826,I880852,);
and I_51655 (I880860,I880852,I478067);
DFFARX1 I_51656 (I880860,I2683,I880826,I880809,);
DFFARX1 I_51657 (I478082,I2683,I880826,I880900,);
not I_51658 (I880908,I478073);
not I_51659 (I880925,I478064);
nand I_51660 (I880942,I880925,I880908);
nor I_51661 (I880797,I880900,I880942);
DFFARX1 I_51662 (I880942,I2683,I880826,I880982,);
not I_51663 (I880818,I880982);
not I_51664 (I881004,I478070);
nand I_51665 (I881021,I880925,I881004);
DFFARX1 I_51666 (I881021,I2683,I880826,I881047,);
not I_51667 (I881055,I881047);
not I_51668 (I881072,I478085);
nand I_51669 (I881089,I881072,I478088);
and I_51670 (I881106,I880908,I881089);
nor I_51671 (I881123,I881021,I881106);
DFFARX1 I_51672 (I881123,I2683,I880826,I880794,);
DFFARX1 I_51673 (I881106,I2683,I880826,I880815,);
nor I_51674 (I881168,I478085,I478064);
nor I_51675 (I880806,I881021,I881168);
or I_51676 (I881199,I478085,I478064);
nor I_51677 (I881216,I478076,I478067);
DFFARX1 I_51678 (I881216,I2683,I880826,I881242,);
not I_51679 (I881250,I881242);
nor I_51680 (I880812,I881250,I881055);
nand I_51681 (I881281,I881250,I880900);
not I_51682 (I881298,I478076);
nand I_51683 (I881315,I881298,I881004);
nand I_51684 (I881332,I881250,I881315);
nand I_51685 (I880803,I881332,I881281);
nand I_51686 (I880800,I881315,I881199);
not I_51687 (I881404,I2690);
DFFARX1 I_51688 (I756819,I2683,I881404,I881430,);
and I_51689 (I881438,I881430,I756813);
DFFARX1 I_51690 (I881438,I2683,I881404,I881387,);
DFFARX1 I_51691 (I756831,I2683,I881404,I881478,);
not I_51692 (I881486,I756822);
not I_51693 (I881503,I756834);
nand I_51694 (I881520,I881503,I881486);
nor I_51695 (I881375,I881478,I881520);
DFFARX1 I_51696 (I881520,I2683,I881404,I881560,);
not I_51697 (I881396,I881560);
not I_51698 (I881582,I756840);
nand I_51699 (I881599,I881503,I881582);
DFFARX1 I_51700 (I881599,I2683,I881404,I881625,);
not I_51701 (I881633,I881625);
not I_51702 (I881650,I756816);
nand I_51703 (I881667,I881650,I756837);
and I_51704 (I881684,I881486,I881667);
nor I_51705 (I881701,I881599,I881684);
DFFARX1 I_51706 (I881701,I2683,I881404,I881372,);
DFFARX1 I_51707 (I881684,I2683,I881404,I881393,);
nor I_51708 (I881746,I756816,I756828);
nor I_51709 (I881384,I881599,I881746);
or I_51710 (I881777,I756816,I756828);
nor I_51711 (I881794,I756813,I756825);
DFFARX1 I_51712 (I881794,I2683,I881404,I881820,);
not I_51713 (I881828,I881820);
nor I_51714 (I881390,I881828,I881633);
nand I_51715 (I881859,I881828,I881478);
not I_51716 (I881876,I756813);
nand I_51717 (I881893,I881876,I881582);
nand I_51718 (I881910,I881828,I881893);
nand I_51719 (I881381,I881910,I881859);
nand I_51720 (I881378,I881893,I881777);
not I_51721 (I881982,I2690);
DFFARX1 I_51722 (I469987,I2683,I881982,I882008,);
and I_51723 (I882016,I882008,I469975);
DFFARX1 I_51724 (I882016,I2683,I881982,I881965,);
DFFARX1 I_51725 (I469990,I2683,I881982,I882056,);
not I_51726 (I882064,I469981);
not I_51727 (I882081,I469972);
nand I_51728 (I882098,I882081,I882064);
nor I_51729 (I881953,I882056,I882098);
DFFARX1 I_51730 (I882098,I2683,I881982,I882138,);
not I_51731 (I881974,I882138);
not I_51732 (I882160,I469978);
nand I_51733 (I882177,I882081,I882160);
DFFARX1 I_51734 (I882177,I2683,I881982,I882203,);
not I_51735 (I882211,I882203);
not I_51736 (I882228,I469993);
nand I_51737 (I882245,I882228,I469996);
and I_51738 (I882262,I882064,I882245);
nor I_51739 (I882279,I882177,I882262);
DFFARX1 I_51740 (I882279,I2683,I881982,I881950,);
DFFARX1 I_51741 (I882262,I2683,I881982,I881971,);
nor I_51742 (I882324,I469993,I469972);
nor I_51743 (I881962,I882177,I882324);
or I_51744 (I882355,I469993,I469972);
nor I_51745 (I882372,I469984,I469975);
DFFARX1 I_51746 (I882372,I2683,I881982,I882398,);
not I_51747 (I882406,I882398);
nor I_51748 (I881968,I882406,I882211);
nand I_51749 (I882437,I882406,I882056);
not I_51750 (I882454,I469984);
nand I_51751 (I882471,I882454,I882160);
nand I_51752 (I882488,I882406,I882471);
nand I_51753 (I881959,I882488,I882437);
nand I_51754 (I881956,I882471,I882355);
not I_51755 (I882560,I2690);
DFFARX1 I_51756 (I546283,I2683,I882560,I882586,);
and I_51757 (I882594,I882586,I546271);
DFFARX1 I_51758 (I882594,I2683,I882560,I882543,);
DFFARX1 I_51759 (I546274,I2683,I882560,I882634,);
not I_51760 (I882642,I546268);
not I_51761 (I882659,I546292);
nand I_51762 (I882676,I882659,I882642);
nor I_51763 (I882531,I882634,I882676);
DFFARX1 I_51764 (I882676,I2683,I882560,I882716,);
not I_51765 (I882552,I882716);
not I_51766 (I882738,I546280);
nand I_51767 (I882755,I882659,I882738);
DFFARX1 I_51768 (I882755,I2683,I882560,I882781,);
not I_51769 (I882789,I882781);
not I_51770 (I882806,I546289);
nand I_51771 (I882823,I882806,I546286);
and I_51772 (I882840,I882642,I882823);
nor I_51773 (I882857,I882755,I882840);
DFFARX1 I_51774 (I882857,I2683,I882560,I882528,);
DFFARX1 I_51775 (I882840,I2683,I882560,I882549,);
nor I_51776 (I882902,I546289,I546277);
nor I_51777 (I882540,I882755,I882902);
or I_51778 (I882933,I546289,I546277);
nor I_51779 (I882950,I546268,I546271);
DFFARX1 I_51780 (I882950,I2683,I882560,I882976,);
not I_51781 (I882984,I882976);
nor I_51782 (I882546,I882984,I882789);
nand I_51783 (I883015,I882984,I882634);
not I_51784 (I883032,I546268);
nand I_51785 (I883049,I883032,I882738);
nand I_51786 (I883066,I882984,I883049);
nand I_51787 (I882537,I883066,I883015);
nand I_51788 (I882534,I883049,I882933);
not I_51789 (I883138,I2690);
DFFARX1 I_51790 (I826516,I2683,I883138,I883164,);
and I_51791 (I883172,I883164,I826513);
DFFARX1 I_51792 (I883172,I2683,I883138,I883121,);
DFFARX1 I_51793 (I826519,I2683,I883138,I883212,);
not I_51794 (I883220,I826522);
not I_51795 (I883237,I826516);
nand I_51796 (I883254,I883237,I883220);
nor I_51797 (I883109,I883212,I883254);
DFFARX1 I_51798 (I883254,I2683,I883138,I883294,);
not I_51799 (I883130,I883294);
not I_51800 (I883316,I826531);
nand I_51801 (I883333,I883237,I883316);
DFFARX1 I_51802 (I883333,I2683,I883138,I883359,);
not I_51803 (I883367,I883359);
not I_51804 (I883384,I826528);
nand I_51805 (I883401,I883384,I826534);
and I_51806 (I883418,I883220,I883401);
nor I_51807 (I883435,I883333,I883418);
DFFARX1 I_51808 (I883435,I2683,I883138,I883106,);
DFFARX1 I_51809 (I883418,I2683,I883138,I883127,);
nor I_51810 (I883480,I826528,I826513);
nor I_51811 (I883118,I883333,I883480);
or I_51812 (I883511,I826528,I826513);
nor I_51813 (I883528,I826525,I826519);
DFFARX1 I_51814 (I883528,I2683,I883138,I883554,);
not I_51815 (I883562,I883554);
nor I_51816 (I883124,I883562,I883367);
nand I_51817 (I883593,I883562,I883212);
not I_51818 (I883610,I826525);
nand I_51819 (I883627,I883610,I883316);
nand I_51820 (I883644,I883562,I883627);
nand I_51821 (I883115,I883644,I883593);
nand I_51822 (I883112,I883627,I883511);
not I_51823 (I883716,I2690);
DFFARX1 I_51824 (I289136,I2683,I883716,I883742,);
and I_51825 (I883750,I883742,I289121);
DFFARX1 I_51826 (I883750,I2683,I883716,I883699,);
DFFARX1 I_51827 (I289127,I2683,I883716,I883790,);
not I_51828 (I883798,I289109);
not I_51829 (I883815,I289130);
nand I_51830 (I883832,I883815,I883798);
nor I_51831 (I883687,I883790,I883832);
DFFARX1 I_51832 (I883832,I2683,I883716,I883872,);
not I_51833 (I883708,I883872);
not I_51834 (I883894,I289133);
nand I_51835 (I883911,I883815,I883894);
DFFARX1 I_51836 (I883911,I2683,I883716,I883937,);
not I_51837 (I883945,I883937);
not I_51838 (I883962,I289124);
nand I_51839 (I883979,I883962,I289112);
and I_51840 (I883996,I883798,I883979);
nor I_51841 (I884013,I883911,I883996);
DFFARX1 I_51842 (I884013,I2683,I883716,I883684,);
DFFARX1 I_51843 (I883996,I2683,I883716,I883705,);
nor I_51844 (I884058,I289124,I289118);
nor I_51845 (I883696,I883911,I884058);
or I_51846 (I884089,I289124,I289118);
nor I_51847 (I884106,I289115,I289109);
DFFARX1 I_51848 (I884106,I2683,I883716,I884132,);
not I_51849 (I884140,I884132);
nor I_51850 (I883702,I884140,I883945);
nand I_51851 (I884171,I884140,I883790);
not I_51852 (I884188,I289115);
nand I_51853 (I884205,I884188,I883894);
nand I_51854 (I884222,I884140,I884205);
nand I_51855 (I883693,I884222,I884171);
nand I_51856 (I883690,I884205,I884089);
not I_51857 (I884294,I2690);
DFFARX1 I_51858 (I58545,I2683,I884294,I884320,);
and I_51859 (I884328,I884320,I58521);
DFFARX1 I_51860 (I884328,I2683,I884294,I884277,);
DFFARX1 I_51861 (I58539,I2683,I884294,I884368,);
not I_51862 (I884376,I58527);
not I_51863 (I884393,I58524);
nand I_51864 (I884410,I884393,I884376);
nor I_51865 (I884265,I884368,I884410);
DFFARX1 I_51866 (I884410,I2683,I884294,I884450,);
not I_51867 (I884286,I884450);
not I_51868 (I884472,I58533);
nand I_51869 (I884489,I884393,I884472);
DFFARX1 I_51870 (I884489,I2683,I884294,I884515,);
not I_51871 (I884523,I884515);
not I_51872 (I884540,I58524);
nand I_51873 (I884557,I884540,I58542);
and I_51874 (I884574,I884376,I884557);
nor I_51875 (I884591,I884489,I884574);
DFFARX1 I_51876 (I884591,I2683,I884294,I884262,);
DFFARX1 I_51877 (I884574,I2683,I884294,I884283,);
nor I_51878 (I884636,I58524,I58536);
nor I_51879 (I884274,I884489,I884636);
or I_51880 (I884667,I58524,I58536);
nor I_51881 (I884684,I58530,I58521);
DFFARX1 I_51882 (I884684,I2683,I884294,I884710,);
not I_51883 (I884718,I884710);
nor I_51884 (I884280,I884718,I884523);
nand I_51885 (I884749,I884718,I884368);
not I_51886 (I884766,I58530);
nand I_51887 (I884783,I884766,I884472);
nand I_51888 (I884800,I884718,I884783);
nand I_51889 (I884271,I884800,I884749);
nand I_51890 (I884268,I884783,I884667);
not I_51891 (I884872,I2690);
DFFARX1 I_51892 (I23212,I2683,I884872,I884898,);
and I_51893 (I884906,I884898,I23215);
DFFARX1 I_51894 (I884906,I2683,I884872,I884855,);
DFFARX1 I_51895 (I23215,I2683,I884872,I884946,);
not I_51896 (I884954,I23218);
not I_51897 (I884971,I23233);
nand I_51898 (I884988,I884971,I884954);
nor I_51899 (I884843,I884946,I884988);
DFFARX1 I_51900 (I884988,I2683,I884872,I885028,);
not I_51901 (I884864,I885028);
not I_51902 (I885050,I23227);
nand I_51903 (I885067,I884971,I885050);
DFFARX1 I_51904 (I885067,I2683,I884872,I885093,);
not I_51905 (I885101,I885093);
not I_51906 (I885118,I23230);
nand I_51907 (I885135,I885118,I23212);
and I_51908 (I885152,I884954,I885135);
nor I_51909 (I885169,I885067,I885152);
DFFARX1 I_51910 (I885169,I2683,I884872,I884840,);
DFFARX1 I_51911 (I885152,I2683,I884872,I884861,);
nor I_51912 (I885214,I23230,I23224);
nor I_51913 (I884852,I885067,I885214);
or I_51914 (I885245,I23230,I23224);
nor I_51915 (I885262,I23221,I23236);
DFFARX1 I_51916 (I885262,I2683,I884872,I885288,);
not I_51917 (I885296,I885288);
nor I_51918 (I884858,I885296,I885101);
nand I_51919 (I885327,I885296,I884946);
not I_51920 (I885344,I23221);
nand I_51921 (I885361,I885344,I885050);
nand I_51922 (I885378,I885296,I885361);
nand I_51923 (I884849,I885378,I885327);
nand I_51924 (I884846,I885361,I885245);
not I_51925 (I885450,I2690);
DFFARX1 I_51926 (I540503,I2683,I885450,I885476,);
and I_51927 (I885484,I885476,I540491);
DFFARX1 I_51928 (I885484,I2683,I885450,I885433,);
DFFARX1 I_51929 (I540494,I2683,I885450,I885524,);
not I_51930 (I885532,I540488);
not I_51931 (I885549,I540512);
nand I_51932 (I885566,I885549,I885532);
nor I_51933 (I885421,I885524,I885566);
DFFARX1 I_51934 (I885566,I2683,I885450,I885606,);
not I_51935 (I885442,I885606);
not I_51936 (I885628,I540500);
nand I_51937 (I885645,I885549,I885628);
DFFARX1 I_51938 (I885645,I2683,I885450,I885671,);
not I_51939 (I885679,I885671);
not I_51940 (I885696,I540509);
nand I_51941 (I885713,I885696,I540506);
and I_51942 (I885730,I885532,I885713);
nor I_51943 (I885747,I885645,I885730);
DFFARX1 I_51944 (I885747,I2683,I885450,I885418,);
DFFARX1 I_51945 (I885730,I2683,I885450,I885439,);
nor I_51946 (I885792,I540509,I540497);
nor I_51947 (I885430,I885645,I885792);
or I_51948 (I885823,I540509,I540497);
nor I_51949 (I885840,I540488,I540491);
DFFARX1 I_51950 (I885840,I2683,I885450,I885866,);
not I_51951 (I885874,I885866);
nor I_51952 (I885436,I885874,I885679);
nand I_51953 (I885905,I885874,I885524);
not I_51954 (I885922,I540488);
nand I_51955 (I885939,I885922,I885628);
nand I_51956 (I885956,I885874,I885939);
nand I_51957 (I885427,I885956,I885905);
nand I_51958 (I885424,I885939,I885823);
not I_51959 (I886028,I2690);
DFFARX1 I_51960 (I196765,I2683,I886028,I886054,);
and I_51961 (I886062,I886054,I196768);
DFFARX1 I_51962 (I886062,I2683,I886028,I886011,);
DFFARX1 I_51963 (I196768,I2683,I886028,I886102,);
not I_51964 (I886110,I196783);
not I_51965 (I886127,I196789);
nand I_51966 (I886144,I886127,I886110);
nor I_51967 (I885999,I886102,I886144);
DFFARX1 I_51968 (I886144,I2683,I886028,I886184,);
not I_51969 (I886020,I886184);
not I_51970 (I886206,I196777);
nand I_51971 (I886223,I886127,I886206);
DFFARX1 I_51972 (I886223,I2683,I886028,I886249,);
not I_51973 (I886257,I886249);
not I_51974 (I886274,I196774);
nand I_51975 (I886291,I886274,I196771);
and I_51976 (I886308,I886110,I886291);
nor I_51977 (I886325,I886223,I886308);
DFFARX1 I_51978 (I886325,I2683,I886028,I885996,);
DFFARX1 I_51979 (I886308,I2683,I886028,I886017,);
nor I_51980 (I886370,I196774,I196765);
nor I_51981 (I886008,I886223,I886370);
or I_51982 (I886401,I196774,I196765);
nor I_51983 (I886418,I196780,I196786);
DFFARX1 I_51984 (I886418,I2683,I886028,I886444,);
not I_51985 (I886452,I886444);
nor I_51986 (I886014,I886452,I886257);
nand I_51987 (I886483,I886452,I886102);
not I_51988 (I886500,I196780);
nand I_51989 (I886517,I886500,I886206);
nand I_51990 (I886534,I886452,I886517);
nand I_51991 (I886005,I886534,I886483);
nand I_51992 (I886002,I886517,I886401);
not I_51993 (I886606,I2690);
DFFARX1 I_51994 (I15307,I2683,I886606,I886632,);
and I_51995 (I886640,I886632,I15310);
DFFARX1 I_51996 (I886640,I2683,I886606,I886589,);
DFFARX1 I_51997 (I15310,I2683,I886606,I886680,);
not I_51998 (I886688,I15313);
not I_51999 (I886705,I15328);
nand I_52000 (I886722,I886705,I886688);
nor I_52001 (I886577,I886680,I886722);
DFFARX1 I_52002 (I886722,I2683,I886606,I886762,);
not I_52003 (I886598,I886762);
not I_52004 (I886784,I15322);
nand I_52005 (I886801,I886705,I886784);
DFFARX1 I_52006 (I886801,I2683,I886606,I886827,);
not I_52007 (I886835,I886827);
not I_52008 (I886852,I15325);
nand I_52009 (I886869,I886852,I15307);
and I_52010 (I886886,I886688,I886869);
nor I_52011 (I886903,I886801,I886886);
DFFARX1 I_52012 (I886903,I2683,I886606,I886574,);
DFFARX1 I_52013 (I886886,I2683,I886606,I886595,);
nor I_52014 (I886948,I15325,I15319);
nor I_52015 (I886586,I886801,I886948);
or I_52016 (I886979,I15325,I15319);
nor I_52017 (I886996,I15316,I15331);
DFFARX1 I_52018 (I886996,I2683,I886606,I887022,);
not I_52019 (I887030,I887022);
nor I_52020 (I886592,I887030,I886835);
nand I_52021 (I887061,I887030,I886680);
not I_52022 (I887078,I15316);
nand I_52023 (I887095,I887078,I886784);
nand I_52024 (I887112,I887030,I887095);
nand I_52025 (I886583,I887112,I887061);
nand I_52026 (I886580,I887095,I886979);
not I_52027 (I887184,I2690);
DFFARX1 I_52028 (I379634,I2683,I887184,I887210,);
and I_52029 (I887218,I887210,I379649);
DFFARX1 I_52030 (I887218,I2683,I887184,I887167,);
DFFARX1 I_52031 (I379652,I2683,I887184,I887258,);
not I_52032 (I887266,I379646);
not I_52033 (I887283,I379661);
nand I_52034 (I887300,I887283,I887266);
nor I_52035 (I887155,I887258,I887300);
DFFARX1 I_52036 (I887300,I2683,I887184,I887340,);
not I_52037 (I887176,I887340);
not I_52038 (I887362,I379637);
nand I_52039 (I887379,I887283,I887362);
DFFARX1 I_52040 (I887379,I2683,I887184,I887405,);
not I_52041 (I887413,I887405);
not I_52042 (I887430,I379640);
nand I_52043 (I887447,I887430,I379634);
and I_52044 (I887464,I887266,I887447);
nor I_52045 (I887481,I887379,I887464);
DFFARX1 I_52046 (I887481,I2683,I887184,I887152,);
DFFARX1 I_52047 (I887464,I2683,I887184,I887173,);
nor I_52048 (I887526,I379640,I379643);
nor I_52049 (I887164,I887379,I887526);
or I_52050 (I887557,I379640,I379643);
nor I_52051 (I887574,I379658,I379655);
DFFARX1 I_52052 (I887574,I2683,I887184,I887600,);
not I_52053 (I887608,I887600);
nor I_52054 (I887170,I887608,I887413);
nand I_52055 (I887639,I887608,I887258);
not I_52056 (I887656,I379658);
nand I_52057 (I887673,I887656,I887362);
nand I_52058 (I887690,I887608,I887673);
nand I_52059 (I887161,I887690,I887639);
nand I_52060 (I887158,I887673,I887557);
not I_52061 (I887762,I2690);
DFFARX1 I_52062 (I161660,I2683,I887762,I887788,);
and I_52063 (I887796,I887788,I161663);
DFFARX1 I_52064 (I887796,I2683,I887762,I887745,);
DFFARX1 I_52065 (I161663,I2683,I887762,I887836,);
not I_52066 (I887844,I161678);
not I_52067 (I887861,I161684);
nand I_52068 (I887878,I887861,I887844);
nor I_52069 (I887733,I887836,I887878);
DFFARX1 I_52070 (I887878,I2683,I887762,I887918,);
not I_52071 (I887754,I887918);
not I_52072 (I887940,I161672);
nand I_52073 (I887957,I887861,I887940);
DFFARX1 I_52074 (I887957,I2683,I887762,I887983,);
not I_52075 (I887991,I887983);
not I_52076 (I888008,I161669);
nand I_52077 (I888025,I888008,I161666);
and I_52078 (I888042,I887844,I888025);
nor I_52079 (I888059,I887957,I888042);
DFFARX1 I_52080 (I888059,I2683,I887762,I887730,);
DFFARX1 I_52081 (I888042,I2683,I887762,I887751,);
nor I_52082 (I888104,I161669,I161660);
nor I_52083 (I887742,I887957,I888104);
or I_52084 (I888135,I161669,I161660);
nor I_52085 (I888152,I161675,I161681);
DFFARX1 I_52086 (I888152,I2683,I887762,I888178,);
not I_52087 (I888186,I888178);
nor I_52088 (I887748,I888186,I887991);
nand I_52089 (I888217,I888186,I887836);
not I_52090 (I888234,I161675);
nand I_52091 (I888251,I888234,I887940);
nand I_52092 (I888268,I888186,I888251);
nand I_52093 (I887739,I888268,I888217);
nand I_52094 (I887736,I888251,I888135);
not I_52095 (I888340,I2690);
DFFARX1 I_52096 (I288609,I2683,I888340,I888366,);
and I_52097 (I888374,I888366,I288594);
DFFARX1 I_52098 (I888374,I2683,I888340,I888323,);
DFFARX1 I_52099 (I288600,I2683,I888340,I888414,);
not I_52100 (I888422,I288582);
not I_52101 (I888439,I288603);
nand I_52102 (I888456,I888439,I888422);
nor I_52103 (I888311,I888414,I888456);
DFFARX1 I_52104 (I888456,I2683,I888340,I888496,);
not I_52105 (I888332,I888496);
not I_52106 (I888518,I288606);
nand I_52107 (I888535,I888439,I888518);
DFFARX1 I_52108 (I888535,I2683,I888340,I888561,);
not I_52109 (I888569,I888561);
not I_52110 (I888586,I288597);
nand I_52111 (I888603,I888586,I288585);
and I_52112 (I888620,I888422,I888603);
nor I_52113 (I888637,I888535,I888620);
DFFARX1 I_52114 (I888637,I2683,I888340,I888308,);
DFFARX1 I_52115 (I888620,I2683,I888340,I888329,);
nor I_52116 (I888682,I288597,I288591);
nor I_52117 (I888320,I888535,I888682);
or I_52118 (I888713,I288597,I288591);
nor I_52119 (I888730,I288588,I288582);
DFFARX1 I_52120 (I888730,I2683,I888340,I888756,);
not I_52121 (I888764,I888756);
nor I_52122 (I888326,I888764,I888569);
nand I_52123 (I888795,I888764,I888414);
not I_52124 (I888812,I288588);
nand I_52125 (I888829,I888812,I888518);
nand I_52126 (I888846,I888764,I888829);
nand I_52127 (I888317,I888846,I888795);
nand I_52128 (I888314,I888829,I888713);
not I_52129 (I888918,I2690);
DFFARX1 I_52130 (I1078106,I2683,I888918,I888944,);
and I_52131 (I888952,I888944,I1078088);
DFFARX1 I_52132 (I888952,I2683,I888918,I888901,);
DFFARX1 I_52133 (I1078079,I2683,I888918,I888992,);
not I_52134 (I889000,I1078094);
not I_52135 (I889017,I1078082);
nand I_52136 (I889034,I889017,I889000);
nor I_52137 (I888889,I888992,I889034);
DFFARX1 I_52138 (I889034,I2683,I888918,I889074,);
not I_52139 (I888910,I889074);
not I_52140 (I889096,I1078091);
nand I_52141 (I889113,I889017,I889096);
DFFARX1 I_52142 (I889113,I2683,I888918,I889139,);
not I_52143 (I889147,I889139);
not I_52144 (I889164,I1078100);
nand I_52145 (I889181,I889164,I1078079);
and I_52146 (I889198,I889000,I889181);
nor I_52147 (I889215,I889113,I889198);
DFFARX1 I_52148 (I889215,I2683,I888918,I888886,);
DFFARX1 I_52149 (I889198,I2683,I888918,I888907,);
nor I_52150 (I889260,I1078100,I1078103);
nor I_52151 (I888898,I889113,I889260);
or I_52152 (I889291,I1078100,I1078103);
nor I_52153 (I889308,I1078097,I1078085);
DFFARX1 I_52154 (I889308,I2683,I888918,I889334,);
not I_52155 (I889342,I889334);
nor I_52156 (I888904,I889342,I889147);
nand I_52157 (I889373,I889342,I888992);
not I_52158 (I889390,I1078097);
nand I_52159 (I889407,I889390,I889096);
nand I_52160 (I889424,I889342,I889407);
nand I_52161 (I888895,I889424,I889373);
nand I_52162 (I888892,I889407,I889291);
not I_52163 (I889496,I2690);
DFFARX1 I_52164 (I58018,I2683,I889496,I889522,);
and I_52165 (I889530,I889522,I57994);
DFFARX1 I_52166 (I889530,I2683,I889496,I889479,);
DFFARX1 I_52167 (I58012,I2683,I889496,I889570,);
not I_52168 (I889578,I58000);
not I_52169 (I889595,I57997);
nand I_52170 (I889612,I889595,I889578);
nor I_52171 (I889467,I889570,I889612);
DFFARX1 I_52172 (I889612,I2683,I889496,I889652,);
not I_52173 (I889488,I889652);
not I_52174 (I889674,I58006);
nand I_52175 (I889691,I889595,I889674);
DFFARX1 I_52176 (I889691,I2683,I889496,I889717,);
not I_52177 (I889725,I889717);
not I_52178 (I889742,I57997);
nand I_52179 (I889759,I889742,I58015);
and I_52180 (I889776,I889578,I889759);
nor I_52181 (I889793,I889691,I889776);
DFFARX1 I_52182 (I889793,I2683,I889496,I889464,);
DFFARX1 I_52183 (I889776,I2683,I889496,I889485,);
nor I_52184 (I889838,I57997,I58009);
nor I_52185 (I889476,I889691,I889838);
or I_52186 (I889869,I57997,I58009);
nor I_52187 (I889886,I58003,I57994);
DFFARX1 I_52188 (I889886,I2683,I889496,I889912,);
not I_52189 (I889920,I889912);
nor I_52190 (I889482,I889920,I889725);
nand I_52191 (I889951,I889920,I889570);
not I_52192 (I889968,I58003);
nand I_52193 (I889985,I889968,I889674);
nand I_52194 (I890002,I889920,I889985);
nand I_52195 (I889473,I890002,I889951);
nand I_52196 (I889470,I889985,I889869);
not I_52197 (I890074,I2690);
DFFARX1 I_52198 (I405035,I2683,I890074,I890100,);
and I_52199 (I890108,I890100,I405050);
DFFARX1 I_52200 (I890108,I2683,I890074,I890057,);
DFFARX1 I_52201 (I405041,I2683,I890074,I890148,);
not I_52202 (I890156,I405035);
not I_52203 (I890173,I405053);
nand I_52204 (I890190,I890173,I890156);
nor I_52205 (I890045,I890148,I890190);
DFFARX1 I_52206 (I890190,I2683,I890074,I890230,);
not I_52207 (I890066,I890230);
not I_52208 (I890252,I405044);
nand I_52209 (I890269,I890173,I890252);
DFFARX1 I_52210 (I890269,I2683,I890074,I890295,);
not I_52211 (I890303,I890295);
not I_52212 (I890320,I405056);
nand I_52213 (I890337,I890320,I405032);
and I_52214 (I890354,I890156,I890337);
nor I_52215 (I890371,I890269,I890354);
DFFARX1 I_52216 (I890371,I2683,I890074,I890042,);
DFFARX1 I_52217 (I890354,I2683,I890074,I890063,);
nor I_52218 (I890416,I405056,I405032);
nor I_52219 (I890054,I890269,I890416);
or I_52220 (I890447,I405056,I405032);
nor I_52221 (I890464,I405038,I405047);
DFFARX1 I_52222 (I890464,I2683,I890074,I890490,);
not I_52223 (I890498,I890490);
nor I_52224 (I890060,I890498,I890303);
nand I_52225 (I890529,I890498,I890148);
not I_52226 (I890546,I405038);
nand I_52227 (I890563,I890546,I890252);
nand I_52228 (I890580,I890498,I890563);
nand I_52229 (I890051,I890580,I890529);
nand I_52230 (I890048,I890563,I890447);
not I_52231 (I890652,I2690);
DFFARX1 I_52232 (I1025991,I2683,I890652,I890678,);
and I_52233 (I890686,I890678,I1026018);
DFFARX1 I_52234 (I890686,I2683,I890652,I890635,);
DFFARX1 I_52235 (I1026000,I2683,I890652,I890726,);
not I_52236 (I890734,I1026009);
not I_52237 (I890751,I1026012);
nand I_52238 (I890768,I890751,I890734);
nor I_52239 (I890623,I890726,I890768);
DFFARX1 I_52240 (I890768,I2683,I890652,I890808,);
not I_52241 (I890644,I890808);
not I_52242 (I890830,I1026006);
nand I_52243 (I890847,I890751,I890830);
DFFARX1 I_52244 (I890847,I2683,I890652,I890873,);
not I_52245 (I890881,I890873);
not I_52246 (I890898,I1025994);
nand I_52247 (I890915,I890898,I1025997);
and I_52248 (I890932,I890734,I890915);
nor I_52249 (I890949,I890847,I890932);
DFFARX1 I_52250 (I890949,I2683,I890652,I890620,);
DFFARX1 I_52251 (I890932,I2683,I890652,I890641,);
nor I_52252 (I890994,I1025994,I1026015);
nor I_52253 (I890632,I890847,I890994);
or I_52254 (I891025,I1025994,I1026015);
nor I_52255 (I891042,I1026003,I1025991);
DFFARX1 I_52256 (I891042,I2683,I890652,I891068,);
not I_52257 (I891076,I891068);
nor I_52258 (I890638,I891076,I890881);
nand I_52259 (I891107,I891076,I890726);
not I_52260 (I891124,I1026003);
nand I_52261 (I891141,I891124,I890830);
nand I_52262 (I891158,I891076,I891141);
nand I_52263 (I890629,I891158,I891107);
nand I_52264 (I890626,I891141,I891025);
not I_52265 (I891230,I2690);
DFFARX1 I_52266 (I352434,I2683,I891230,I891256,);
and I_52267 (I891264,I891256,I352449);
DFFARX1 I_52268 (I891264,I2683,I891230,I891213,);
DFFARX1 I_52269 (I352452,I2683,I891230,I891304,);
not I_52270 (I891312,I352446);
not I_52271 (I891329,I352461);
nand I_52272 (I891346,I891329,I891312);
nor I_52273 (I891201,I891304,I891346);
DFFARX1 I_52274 (I891346,I2683,I891230,I891386,);
not I_52275 (I891222,I891386);
not I_52276 (I891408,I352437);
nand I_52277 (I891425,I891329,I891408);
DFFARX1 I_52278 (I891425,I2683,I891230,I891451,);
not I_52279 (I891459,I891451);
not I_52280 (I891476,I352440);
nand I_52281 (I891493,I891476,I352434);
and I_52282 (I891510,I891312,I891493);
nor I_52283 (I891527,I891425,I891510);
DFFARX1 I_52284 (I891527,I2683,I891230,I891198,);
DFFARX1 I_52285 (I891510,I2683,I891230,I891219,);
nor I_52286 (I891572,I352440,I352443);
nor I_52287 (I891210,I891425,I891572);
or I_52288 (I891603,I352440,I352443);
nor I_52289 (I891620,I352458,I352455);
DFFARX1 I_52290 (I891620,I2683,I891230,I891646,);
not I_52291 (I891654,I891646);
nor I_52292 (I891216,I891654,I891459);
nand I_52293 (I891685,I891654,I891304);
not I_52294 (I891702,I352458);
nand I_52295 (I891719,I891702,I891408);
nand I_52296 (I891736,I891654,I891719);
nand I_52297 (I891207,I891736,I891685);
nand I_52298 (I891204,I891719,I891603);
not I_52299 (I891808,I2690);
DFFARX1 I_52300 (I574605,I2683,I891808,I891834,);
and I_52301 (I891842,I891834,I574593);
DFFARX1 I_52302 (I891842,I2683,I891808,I891791,);
DFFARX1 I_52303 (I574596,I2683,I891808,I891882,);
not I_52304 (I891890,I574590);
not I_52305 (I891907,I574614);
nand I_52306 (I891924,I891907,I891890);
nor I_52307 (I891779,I891882,I891924);
DFFARX1 I_52308 (I891924,I2683,I891808,I891964,);
not I_52309 (I891800,I891964);
not I_52310 (I891986,I574602);
nand I_52311 (I892003,I891907,I891986);
DFFARX1 I_52312 (I892003,I2683,I891808,I892029,);
not I_52313 (I892037,I892029);
not I_52314 (I892054,I574611);
nand I_52315 (I892071,I892054,I574608);
and I_52316 (I892088,I891890,I892071);
nor I_52317 (I892105,I892003,I892088);
DFFARX1 I_52318 (I892105,I2683,I891808,I891776,);
DFFARX1 I_52319 (I892088,I2683,I891808,I891797,);
nor I_52320 (I892150,I574611,I574599);
nor I_52321 (I891788,I892003,I892150);
or I_52322 (I892181,I574611,I574599);
nor I_52323 (I892198,I574590,I574593);
DFFARX1 I_52324 (I892198,I2683,I891808,I892224,);
not I_52325 (I892232,I892224);
nor I_52326 (I891794,I892232,I892037);
nand I_52327 (I892263,I892232,I891882);
not I_52328 (I892280,I574590);
nand I_52329 (I892297,I892280,I891986);
nand I_52330 (I892314,I892232,I892297);
nand I_52331 (I891785,I892314,I892263);
nand I_52332 (I891782,I892297,I892181);
not I_52333 (I892386,I2690);
DFFARX1 I_52334 (I1087031,I2683,I892386,I892412,);
and I_52335 (I892420,I892412,I1087013);
DFFARX1 I_52336 (I892420,I2683,I892386,I892369,);
DFFARX1 I_52337 (I1087004,I2683,I892386,I892460,);
not I_52338 (I892468,I1087019);
not I_52339 (I892485,I1087007);
nand I_52340 (I892502,I892485,I892468);
nor I_52341 (I892357,I892460,I892502);
DFFARX1 I_52342 (I892502,I2683,I892386,I892542,);
not I_52343 (I892378,I892542);
not I_52344 (I892564,I1087016);
nand I_52345 (I892581,I892485,I892564);
DFFARX1 I_52346 (I892581,I2683,I892386,I892607,);
not I_52347 (I892615,I892607);
not I_52348 (I892632,I1087025);
nand I_52349 (I892649,I892632,I1087004);
and I_52350 (I892666,I892468,I892649);
nor I_52351 (I892683,I892581,I892666);
DFFARX1 I_52352 (I892683,I2683,I892386,I892354,);
DFFARX1 I_52353 (I892666,I2683,I892386,I892375,);
nor I_52354 (I892728,I1087025,I1087028);
nor I_52355 (I892366,I892581,I892728);
or I_52356 (I892759,I1087025,I1087028);
nor I_52357 (I892776,I1087022,I1087010);
DFFARX1 I_52358 (I892776,I2683,I892386,I892802,);
not I_52359 (I892810,I892802);
nor I_52360 (I892372,I892810,I892615);
nand I_52361 (I892841,I892810,I892460);
not I_52362 (I892858,I1087022);
nand I_52363 (I892875,I892858,I892564);
nand I_52364 (I892892,I892810,I892875);
nand I_52365 (I892363,I892892,I892841);
nand I_52366 (I892360,I892875,I892759);
not I_52367 (I892964,I2690);
DFFARX1 I_52368 (I5088,I2683,I892964,I892990,);
and I_52369 (I892998,I892990,I5094);
DFFARX1 I_52370 (I892998,I2683,I892964,I892947,);
DFFARX1 I_52371 (I5073,I2683,I892964,I893038,);
not I_52372 (I893046,I5079);
not I_52373 (I893063,I5085);
nand I_52374 (I893080,I893063,I893046);
nor I_52375 (I892935,I893038,I893080);
DFFARX1 I_52376 (I893080,I2683,I892964,I893120,);
not I_52377 (I892956,I893120);
not I_52378 (I893142,I5076);
nand I_52379 (I893159,I893063,I893142);
DFFARX1 I_52380 (I893159,I2683,I892964,I893185,);
not I_52381 (I893193,I893185);
not I_52382 (I893210,I5091);
nand I_52383 (I893227,I893210,I5076);
and I_52384 (I893244,I893046,I893227);
nor I_52385 (I893261,I893159,I893244);
DFFARX1 I_52386 (I893261,I2683,I892964,I892932,);
DFFARX1 I_52387 (I893244,I2683,I892964,I892953,);
nor I_52388 (I893306,I5091,I5079);
nor I_52389 (I892944,I893159,I893306);
or I_52390 (I893337,I5091,I5079);
nor I_52391 (I893354,I5082,I5073);
DFFARX1 I_52392 (I893354,I2683,I892964,I893380,);
not I_52393 (I893388,I893380);
nor I_52394 (I892950,I893388,I893193);
nand I_52395 (I893419,I893388,I893038);
not I_52396 (I893436,I5082);
nand I_52397 (I893453,I893436,I893142);
nand I_52398 (I893470,I893388,I893453);
nand I_52399 (I892941,I893470,I893419);
nand I_52400 (I892938,I893453,I893337);
not I_52401 (I893542,I2690);
DFFARX1 I_52402 (I661259,I2683,I893542,I893568,);
and I_52403 (I893576,I893568,I661265);
DFFARX1 I_52404 (I893576,I2683,I893542,I893525,);
DFFARX1 I_52405 (I661271,I2683,I893542,I893616,);
not I_52406 (I893624,I661256);
not I_52407 (I893641,I661256);
nand I_52408 (I893658,I893641,I893624);
nor I_52409 (I893513,I893616,I893658);
DFFARX1 I_52410 (I893658,I2683,I893542,I893698,);
not I_52411 (I893534,I893698);
not I_52412 (I893720,I661274);
nand I_52413 (I893737,I893641,I893720);
DFFARX1 I_52414 (I893737,I2683,I893542,I893763,);
not I_52415 (I893771,I893763);
not I_52416 (I893788,I661268);
nand I_52417 (I893805,I893788,I661259);
and I_52418 (I893822,I893624,I893805);
nor I_52419 (I893839,I893737,I893822);
DFFARX1 I_52420 (I893839,I2683,I893542,I893510,);
DFFARX1 I_52421 (I893822,I2683,I893542,I893531,);
nor I_52422 (I893884,I661268,I661277);
nor I_52423 (I893522,I893737,I893884);
or I_52424 (I893915,I661268,I661277);
nor I_52425 (I893932,I661262,I661262);
DFFARX1 I_52426 (I893932,I2683,I893542,I893958,);
not I_52427 (I893966,I893958);
nor I_52428 (I893528,I893966,I893771);
nand I_52429 (I893997,I893966,I893616);
not I_52430 (I894014,I661262);
nand I_52431 (I894031,I894014,I893720);
nand I_52432 (I894048,I893966,I894031);
nand I_52433 (I893519,I894048,I893997);
nand I_52434 (I893516,I894031,I893915);
not I_52435 (I894120,I2690);
DFFARX1 I_52436 (I689190,I2683,I894120,I894146,);
and I_52437 (I894154,I894146,I689196);
DFFARX1 I_52438 (I894154,I2683,I894120,I894103,);
DFFARX1 I_52439 (I689202,I2683,I894120,I894194,);
not I_52440 (I894202,I689187);
not I_52441 (I894219,I689187);
nand I_52442 (I894236,I894219,I894202);
nor I_52443 (I894091,I894194,I894236);
DFFARX1 I_52444 (I894236,I2683,I894120,I894276,);
not I_52445 (I894112,I894276);
not I_52446 (I894298,I689205);
nand I_52447 (I894315,I894219,I894298);
DFFARX1 I_52448 (I894315,I2683,I894120,I894341,);
not I_52449 (I894349,I894341);
not I_52450 (I894366,I689199);
nand I_52451 (I894383,I894366,I689190);
and I_52452 (I894400,I894202,I894383);
nor I_52453 (I894417,I894315,I894400);
DFFARX1 I_52454 (I894417,I2683,I894120,I894088,);
DFFARX1 I_52455 (I894400,I2683,I894120,I894109,);
nor I_52456 (I894462,I689199,I689208);
nor I_52457 (I894100,I894315,I894462);
or I_52458 (I894493,I689199,I689208);
nor I_52459 (I894510,I689193,I689193);
DFFARX1 I_52460 (I894510,I2683,I894120,I894536,);
not I_52461 (I894544,I894536);
nor I_52462 (I894106,I894544,I894349);
nand I_52463 (I894575,I894544,I894194);
not I_52464 (I894592,I689193);
nand I_52465 (I894609,I894592,I894298);
nand I_52466 (I894626,I894544,I894609);
nand I_52467 (I894097,I894626,I894575);
nand I_52468 (I894094,I894609,I894493);
not I_52469 (I894698,I2690);
DFFARX1 I_52470 (I565357,I2683,I894698,I894724,);
and I_52471 (I894732,I894724,I565345);
DFFARX1 I_52472 (I894732,I2683,I894698,I894681,);
DFFARX1 I_52473 (I565348,I2683,I894698,I894772,);
not I_52474 (I894780,I565342);
not I_52475 (I894797,I565366);
nand I_52476 (I894814,I894797,I894780);
nor I_52477 (I894669,I894772,I894814);
DFFARX1 I_52478 (I894814,I2683,I894698,I894854,);
not I_52479 (I894690,I894854);
not I_52480 (I894876,I565354);
nand I_52481 (I894893,I894797,I894876);
DFFARX1 I_52482 (I894893,I2683,I894698,I894919,);
not I_52483 (I894927,I894919);
not I_52484 (I894944,I565363);
nand I_52485 (I894961,I894944,I565360);
and I_52486 (I894978,I894780,I894961);
nor I_52487 (I894995,I894893,I894978);
DFFARX1 I_52488 (I894995,I2683,I894698,I894666,);
DFFARX1 I_52489 (I894978,I2683,I894698,I894687,);
nor I_52490 (I895040,I565363,I565351);
nor I_52491 (I894678,I894893,I895040);
or I_52492 (I895071,I565363,I565351);
nor I_52493 (I895088,I565342,I565345);
DFFARX1 I_52494 (I895088,I2683,I894698,I895114,);
not I_52495 (I895122,I895114);
nor I_52496 (I894684,I895122,I894927);
nand I_52497 (I895153,I895122,I894772);
not I_52498 (I895170,I565342);
nand I_52499 (I895187,I895170,I894876);
nand I_52500 (I895204,I895122,I895187);
nand I_52501 (I894675,I895204,I895153);
nand I_52502 (I894672,I895187,I895071);
not I_52503 (I895276,I2690);
DFFARX1 I_52504 (I660205,I2683,I895276,I895302,);
and I_52505 (I895310,I895302,I660211);
DFFARX1 I_52506 (I895310,I2683,I895276,I895259,);
DFFARX1 I_52507 (I660217,I2683,I895276,I895350,);
not I_52508 (I895358,I660202);
not I_52509 (I895375,I660202);
nand I_52510 (I895392,I895375,I895358);
nor I_52511 (I895247,I895350,I895392);
DFFARX1 I_52512 (I895392,I2683,I895276,I895432,);
not I_52513 (I895268,I895432);
not I_52514 (I895454,I660220);
nand I_52515 (I895471,I895375,I895454);
DFFARX1 I_52516 (I895471,I2683,I895276,I895497,);
not I_52517 (I895505,I895497);
not I_52518 (I895522,I660214);
nand I_52519 (I895539,I895522,I660205);
and I_52520 (I895556,I895358,I895539);
nor I_52521 (I895573,I895471,I895556);
DFFARX1 I_52522 (I895573,I2683,I895276,I895244,);
DFFARX1 I_52523 (I895556,I2683,I895276,I895265,);
nor I_52524 (I895618,I660214,I660223);
nor I_52525 (I895256,I895471,I895618);
or I_52526 (I895649,I660214,I660223);
nor I_52527 (I895666,I660208,I660208);
DFFARX1 I_52528 (I895666,I2683,I895276,I895692,);
not I_52529 (I895700,I895692);
nor I_52530 (I895262,I895700,I895505);
nand I_52531 (I895731,I895700,I895350);
not I_52532 (I895748,I660208);
nand I_52533 (I895765,I895748,I895454);
nand I_52534 (I895782,I895700,I895765);
nand I_52535 (I895253,I895782,I895731);
nand I_52536 (I895250,I895765,I895649);
not I_52537 (I895854,I2690);
DFFARX1 I_52538 (I186650,I2683,I895854,I895880,);
and I_52539 (I895888,I895880,I186653);
DFFARX1 I_52540 (I895888,I2683,I895854,I895837,);
DFFARX1 I_52541 (I186653,I2683,I895854,I895928,);
not I_52542 (I895936,I186668);
not I_52543 (I895953,I186674);
nand I_52544 (I895970,I895953,I895936);
nor I_52545 (I895825,I895928,I895970);
DFFARX1 I_52546 (I895970,I2683,I895854,I896010,);
not I_52547 (I895846,I896010);
not I_52548 (I896032,I186662);
nand I_52549 (I896049,I895953,I896032);
DFFARX1 I_52550 (I896049,I2683,I895854,I896075,);
not I_52551 (I896083,I896075);
not I_52552 (I896100,I186659);
nand I_52553 (I896117,I896100,I186656);
and I_52554 (I896134,I895936,I896117);
nor I_52555 (I896151,I896049,I896134);
DFFARX1 I_52556 (I896151,I2683,I895854,I895822,);
DFFARX1 I_52557 (I896134,I2683,I895854,I895843,);
nor I_52558 (I896196,I186659,I186650);
nor I_52559 (I895834,I896049,I896196);
or I_52560 (I896227,I186659,I186650);
nor I_52561 (I896244,I186665,I186671);
DFFARX1 I_52562 (I896244,I2683,I895854,I896270,);
not I_52563 (I896278,I896270);
nor I_52564 (I895840,I896278,I896083);
nand I_52565 (I896309,I896278,I895928);
not I_52566 (I896326,I186665);
nand I_52567 (I896343,I896326,I896032);
nand I_52568 (I896360,I896278,I896343);
nand I_52569 (I895831,I896360,I896309);
nand I_52570 (I895828,I896343,I896227);
not I_52571 (I896432,I2690);
DFFARX1 I_52572 (I1040621,I2683,I896432,I896458,);
and I_52573 (I896466,I896458,I1040603);
DFFARX1 I_52574 (I896466,I2683,I896432,I896415,);
DFFARX1 I_52575 (I1040594,I2683,I896432,I896506,);
not I_52576 (I896514,I1040609);
not I_52577 (I896531,I1040597);
nand I_52578 (I896548,I896531,I896514);
nor I_52579 (I896403,I896506,I896548);
DFFARX1 I_52580 (I896548,I2683,I896432,I896588,);
not I_52581 (I896424,I896588);
not I_52582 (I896610,I1040606);
nand I_52583 (I896627,I896531,I896610);
DFFARX1 I_52584 (I896627,I2683,I896432,I896653,);
not I_52585 (I896661,I896653);
not I_52586 (I896678,I1040615);
nand I_52587 (I896695,I896678,I1040594);
and I_52588 (I896712,I896514,I896695);
nor I_52589 (I896729,I896627,I896712);
DFFARX1 I_52590 (I896729,I2683,I896432,I896400,);
DFFARX1 I_52591 (I896712,I2683,I896432,I896421,);
nor I_52592 (I896774,I1040615,I1040618);
nor I_52593 (I896412,I896627,I896774);
or I_52594 (I896805,I1040615,I1040618);
nor I_52595 (I896822,I1040612,I1040600);
DFFARX1 I_52596 (I896822,I2683,I896432,I896848,);
not I_52597 (I896856,I896848);
nor I_52598 (I896418,I896856,I896661);
nand I_52599 (I896887,I896856,I896506);
not I_52600 (I896904,I1040612);
nand I_52601 (I896921,I896904,I896610);
nand I_52602 (I896938,I896856,I896921);
nand I_52603 (I896409,I896938,I896887);
nand I_52604 (I896406,I896921,I896805);
not I_52605 (I897010,I2690);
DFFARX1 I_52606 (I1091196,I2683,I897010,I897036,);
and I_52607 (I897044,I897036,I1091178);
DFFARX1 I_52608 (I897044,I2683,I897010,I896993,);
DFFARX1 I_52609 (I1091169,I2683,I897010,I897084,);
not I_52610 (I897092,I1091184);
not I_52611 (I897109,I1091172);
nand I_52612 (I897126,I897109,I897092);
nor I_52613 (I896981,I897084,I897126);
DFFARX1 I_52614 (I897126,I2683,I897010,I897166,);
not I_52615 (I897002,I897166);
not I_52616 (I897188,I1091181);
nand I_52617 (I897205,I897109,I897188);
DFFARX1 I_52618 (I897205,I2683,I897010,I897231,);
not I_52619 (I897239,I897231);
not I_52620 (I897256,I1091190);
nand I_52621 (I897273,I897256,I1091169);
and I_52622 (I897290,I897092,I897273);
nor I_52623 (I897307,I897205,I897290);
DFFARX1 I_52624 (I897307,I2683,I897010,I896978,);
DFFARX1 I_52625 (I897290,I2683,I897010,I896999,);
nor I_52626 (I897352,I1091190,I1091193);
nor I_52627 (I896990,I897205,I897352);
or I_52628 (I897383,I1091190,I1091193);
nor I_52629 (I897400,I1091187,I1091175);
DFFARX1 I_52630 (I897400,I2683,I897010,I897426,);
not I_52631 (I897434,I897426);
nor I_52632 (I896996,I897434,I897239);
nand I_52633 (I897465,I897434,I897084);
not I_52634 (I897482,I1091187);
nand I_52635 (I897499,I897482,I897188);
nand I_52636 (I897516,I897434,I897499);
nand I_52637 (I896987,I897516,I897465);
nand I_52638 (I896984,I897499,I897383);
not I_52639 (I897588,I2690);
DFFARX1 I_52640 (I616799,I2683,I897588,I897614,);
and I_52641 (I897622,I897614,I616787);
DFFARX1 I_52642 (I897622,I2683,I897588,I897571,);
DFFARX1 I_52643 (I616790,I2683,I897588,I897662,);
not I_52644 (I897670,I616784);
not I_52645 (I897687,I616808);
nand I_52646 (I897704,I897687,I897670);
nor I_52647 (I897559,I897662,I897704);
DFFARX1 I_52648 (I897704,I2683,I897588,I897744,);
not I_52649 (I897580,I897744);
not I_52650 (I897766,I616796);
nand I_52651 (I897783,I897687,I897766);
DFFARX1 I_52652 (I897783,I2683,I897588,I897809,);
not I_52653 (I897817,I897809);
not I_52654 (I897834,I616805);
nand I_52655 (I897851,I897834,I616802);
and I_52656 (I897868,I897670,I897851);
nor I_52657 (I897885,I897783,I897868);
DFFARX1 I_52658 (I897885,I2683,I897588,I897556,);
DFFARX1 I_52659 (I897868,I2683,I897588,I897577,);
nor I_52660 (I897930,I616805,I616793);
nor I_52661 (I897568,I897783,I897930);
or I_52662 (I897961,I616805,I616793);
nor I_52663 (I897978,I616784,I616787);
DFFARX1 I_52664 (I897978,I2683,I897588,I898004,);
not I_52665 (I898012,I898004);
nor I_52666 (I897574,I898012,I897817);
nand I_52667 (I898043,I898012,I897662);
not I_52668 (I898060,I616784);
nand I_52669 (I898077,I898060,I897766);
nand I_52670 (I898094,I898012,I898077);
nand I_52671 (I897565,I898094,I898043);
nand I_52672 (I897562,I898077,I897961);
not I_52673 (I898166,I2690);
DFFARX1 I_52674 (I959219,I2683,I898166,I898192,);
and I_52675 (I898200,I898192,I959213);
DFFARX1 I_52676 (I898200,I2683,I898166,I898149,);
DFFARX1 I_52677 (I959198,I2683,I898166,I898240,);
not I_52678 (I898248,I959204);
not I_52679 (I898265,I959216);
nand I_52680 (I898282,I898265,I898248);
nor I_52681 (I898137,I898240,I898282);
DFFARX1 I_52682 (I898282,I2683,I898166,I898322,);
not I_52683 (I898158,I898322);
not I_52684 (I898344,I959198);
nand I_52685 (I898361,I898265,I898344);
DFFARX1 I_52686 (I898361,I2683,I898166,I898387,);
not I_52687 (I898395,I898387);
not I_52688 (I898412,I959222);
nand I_52689 (I898429,I898412,I959210);
and I_52690 (I898446,I898248,I898429);
nor I_52691 (I898463,I898361,I898446);
DFFARX1 I_52692 (I898463,I2683,I898166,I898134,);
DFFARX1 I_52693 (I898446,I2683,I898166,I898155,);
nor I_52694 (I898508,I959222,I959201);
nor I_52695 (I898146,I898361,I898508);
or I_52696 (I898539,I959222,I959201);
nor I_52697 (I898556,I959207,I959201);
DFFARX1 I_52698 (I898556,I2683,I898166,I898582,);
not I_52699 (I898590,I898582);
nor I_52700 (I898152,I898590,I898395);
nand I_52701 (I898621,I898590,I898240);
not I_52702 (I898638,I959207);
nand I_52703 (I898655,I898638,I898344);
nand I_52704 (I898672,I898590,I898655);
nand I_52705 (I898143,I898672,I898621);
nand I_52706 (I898140,I898655,I898539);
not I_52707 (I898744,I2690);
DFFARX1 I_52708 (I693406,I2683,I898744,I898770,);
and I_52709 (I898778,I898770,I693412);
DFFARX1 I_52710 (I898778,I2683,I898744,I898727,);
DFFARX1 I_52711 (I693418,I2683,I898744,I898818,);
not I_52712 (I898826,I693403);
not I_52713 (I898843,I693403);
nand I_52714 (I898860,I898843,I898826);
nor I_52715 (I898715,I898818,I898860);
DFFARX1 I_52716 (I898860,I2683,I898744,I898900,);
not I_52717 (I898736,I898900);
not I_52718 (I898922,I693421);
nand I_52719 (I898939,I898843,I898922);
DFFARX1 I_52720 (I898939,I2683,I898744,I898965,);
not I_52721 (I898973,I898965);
not I_52722 (I898990,I693415);
nand I_52723 (I899007,I898990,I693406);
and I_52724 (I899024,I898826,I899007);
nor I_52725 (I899041,I898939,I899024);
DFFARX1 I_52726 (I899041,I2683,I898744,I898712,);
DFFARX1 I_52727 (I899024,I2683,I898744,I898733,);
nor I_52728 (I899086,I693415,I693424);
nor I_52729 (I898724,I898939,I899086);
or I_52730 (I899117,I693415,I693424);
nor I_52731 (I899134,I693409,I693409);
DFFARX1 I_52732 (I899134,I2683,I898744,I899160,);
not I_52733 (I899168,I899160);
nor I_52734 (I898730,I899168,I898973);
nand I_52735 (I899199,I899168,I898818);
not I_52736 (I899216,I693409);
nand I_52737 (I899233,I899216,I898922);
nand I_52738 (I899250,I899168,I899233);
nand I_52739 (I898721,I899250,I899199);
nand I_52740 (I898718,I899233,I899117);
not I_52741 (I899322,I2690);
DFFARX1 I_52742 (I449757,I2683,I899322,I899348,);
and I_52743 (I899356,I899348,I449745);
DFFARX1 I_52744 (I899356,I2683,I899322,I899305,);
DFFARX1 I_52745 (I449760,I2683,I899322,I899396,);
not I_52746 (I899404,I449751);
not I_52747 (I899421,I449742);
nand I_52748 (I899438,I899421,I899404);
nor I_52749 (I899293,I899396,I899438);
DFFARX1 I_52750 (I899438,I2683,I899322,I899478,);
not I_52751 (I899314,I899478);
not I_52752 (I899500,I449748);
nand I_52753 (I899517,I899421,I899500);
DFFARX1 I_52754 (I899517,I2683,I899322,I899543,);
not I_52755 (I899551,I899543);
not I_52756 (I899568,I449763);
nand I_52757 (I899585,I899568,I449766);
and I_52758 (I899602,I899404,I899585);
nor I_52759 (I899619,I899517,I899602);
DFFARX1 I_52760 (I899619,I2683,I899322,I899290,);
DFFARX1 I_52761 (I899602,I2683,I899322,I899311,);
nor I_52762 (I899664,I449763,I449742);
nor I_52763 (I899302,I899517,I899664);
or I_52764 (I899695,I449763,I449742);
nor I_52765 (I899712,I449754,I449745);
DFFARX1 I_52766 (I899712,I2683,I899322,I899738,);
not I_52767 (I899746,I899738);
nor I_52768 (I899308,I899746,I899551);
nand I_52769 (I899777,I899746,I899396);
not I_52770 (I899794,I449754);
nand I_52771 (I899811,I899794,I899500);
nand I_52772 (I899828,I899746,I899811);
nand I_52773 (I899299,I899828,I899777);
nand I_52774 (I899296,I899811,I899695);
not I_52775 (I899900,I2690);
DFFARX1 I_52776 (I82260,I2683,I899900,I899926,);
and I_52777 (I899934,I899926,I82236);
DFFARX1 I_52778 (I899934,I2683,I899900,I899883,);
DFFARX1 I_52779 (I82254,I2683,I899900,I899974,);
not I_52780 (I899982,I82242);
not I_52781 (I899999,I82239);
nand I_52782 (I900016,I899999,I899982);
nor I_52783 (I899871,I899974,I900016);
DFFARX1 I_52784 (I900016,I2683,I899900,I900056,);
not I_52785 (I899892,I900056);
not I_52786 (I900078,I82248);
nand I_52787 (I900095,I899999,I900078);
DFFARX1 I_52788 (I900095,I2683,I899900,I900121,);
not I_52789 (I900129,I900121);
not I_52790 (I900146,I82239);
nand I_52791 (I900163,I900146,I82257);
and I_52792 (I900180,I899982,I900163);
nor I_52793 (I900197,I900095,I900180);
DFFARX1 I_52794 (I900197,I2683,I899900,I899868,);
DFFARX1 I_52795 (I900180,I2683,I899900,I899889,);
nor I_52796 (I900242,I82239,I82251);
nor I_52797 (I899880,I900095,I900242);
or I_52798 (I900273,I82239,I82251);
nor I_52799 (I900290,I82245,I82236);
DFFARX1 I_52800 (I900290,I2683,I899900,I900316,);
not I_52801 (I900324,I900316);
nor I_52802 (I899886,I900324,I900129);
nand I_52803 (I900355,I900324,I899974);
not I_52804 (I900372,I82245);
nand I_52805 (I900389,I900372,I900078);
nand I_52806 (I900406,I900324,I900389);
nand I_52807 (I899877,I900406,I900355);
nand I_52808 (I899874,I900389,I900273);
not I_52809 (I900478,I2690);
DFFARX1 I_52810 (I60126,I2683,I900478,I900504,);
and I_52811 (I900512,I900504,I60102);
DFFARX1 I_52812 (I900512,I2683,I900478,I900461,);
DFFARX1 I_52813 (I60120,I2683,I900478,I900552,);
not I_52814 (I900560,I60108);
not I_52815 (I900577,I60105);
nand I_52816 (I900594,I900577,I900560);
nor I_52817 (I900449,I900552,I900594);
DFFARX1 I_52818 (I900594,I2683,I900478,I900634,);
not I_52819 (I900470,I900634);
not I_52820 (I900656,I60114);
nand I_52821 (I900673,I900577,I900656);
DFFARX1 I_52822 (I900673,I2683,I900478,I900699,);
not I_52823 (I900707,I900699);
not I_52824 (I900724,I60105);
nand I_52825 (I900741,I900724,I60123);
and I_52826 (I900758,I900560,I900741);
nor I_52827 (I900775,I900673,I900758);
DFFARX1 I_52828 (I900775,I2683,I900478,I900446,);
DFFARX1 I_52829 (I900758,I2683,I900478,I900467,);
nor I_52830 (I900820,I60105,I60117);
nor I_52831 (I900458,I900673,I900820);
or I_52832 (I900851,I60105,I60117);
nor I_52833 (I900868,I60111,I60102);
DFFARX1 I_52834 (I900868,I2683,I900478,I900894,);
not I_52835 (I900902,I900894);
nor I_52836 (I900464,I900902,I900707);
nand I_52837 (I900933,I900902,I900552);
not I_52838 (I900950,I60111);
nand I_52839 (I900967,I900950,I900656);
nand I_52840 (I900984,I900902,I900967);
nand I_52841 (I900455,I900984,I900933);
nand I_52842 (I900452,I900967,I900851);
not I_52843 (I901056,I2690);
DFFARX1 I_52844 (I824833,I2683,I901056,I901082,);
and I_52845 (I901090,I901082,I824830);
DFFARX1 I_52846 (I901090,I2683,I901056,I901039,);
DFFARX1 I_52847 (I824836,I2683,I901056,I901130,);
not I_52848 (I901138,I824839);
not I_52849 (I901155,I824833);
nand I_52850 (I901172,I901155,I901138);
nor I_52851 (I901027,I901130,I901172);
DFFARX1 I_52852 (I901172,I2683,I901056,I901212,);
not I_52853 (I901048,I901212);
not I_52854 (I901234,I824848);
nand I_52855 (I901251,I901155,I901234);
DFFARX1 I_52856 (I901251,I2683,I901056,I901277,);
not I_52857 (I901285,I901277);
not I_52858 (I901302,I824845);
nand I_52859 (I901319,I901302,I824851);
and I_52860 (I901336,I901138,I901319);
nor I_52861 (I901353,I901251,I901336);
DFFARX1 I_52862 (I901353,I2683,I901056,I901024,);
DFFARX1 I_52863 (I901336,I2683,I901056,I901045,);
nor I_52864 (I901398,I824845,I824830);
nor I_52865 (I901036,I901251,I901398);
or I_52866 (I901429,I824845,I824830);
nor I_52867 (I901446,I824842,I824836);
DFFARX1 I_52868 (I901446,I2683,I901056,I901472,);
not I_52869 (I901480,I901472);
nor I_52870 (I901042,I901480,I901285);
nand I_52871 (I901511,I901480,I901130);
not I_52872 (I901528,I824842);
nand I_52873 (I901545,I901528,I901234);
nand I_52874 (I901562,I901480,I901545);
nand I_52875 (I901033,I901562,I901511);
nand I_52876 (I901030,I901545,I901429);
not I_52877 (I901634,I2690);
DFFARX1 I_52878 (I495997,I2683,I901634,I901660,);
and I_52879 (I901668,I901660,I495985);
DFFARX1 I_52880 (I901668,I2683,I901634,I901617,);
DFFARX1 I_52881 (I496000,I2683,I901634,I901708,);
not I_52882 (I901716,I495991);
not I_52883 (I901733,I495982);
nand I_52884 (I901750,I901733,I901716);
nor I_52885 (I901605,I901708,I901750);
DFFARX1 I_52886 (I901750,I2683,I901634,I901790,);
not I_52887 (I901626,I901790);
not I_52888 (I901812,I495988);
nand I_52889 (I901829,I901733,I901812);
DFFARX1 I_52890 (I901829,I2683,I901634,I901855,);
not I_52891 (I901863,I901855);
not I_52892 (I901880,I496003);
nand I_52893 (I901897,I901880,I496006);
and I_52894 (I901914,I901716,I901897);
nor I_52895 (I901931,I901829,I901914);
DFFARX1 I_52896 (I901931,I2683,I901634,I901602,);
DFFARX1 I_52897 (I901914,I2683,I901634,I901623,);
nor I_52898 (I901976,I496003,I495982);
nor I_52899 (I901614,I901829,I901976);
or I_52900 (I902007,I496003,I495982);
nor I_52901 (I902024,I495994,I495985);
DFFARX1 I_52902 (I902024,I2683,I901634,I902050,);
not I_52903 (I902058,I902050);
nor I_52904 (I901620,I902058,I901863);
nand I_52905 (I902089,I902058,I901708);
not I_52906 (I902106,I495994);
nand I_52907 (I902123,I902106,I901812);
nand I_52908 (I902140,I902058,I902123);
nand I_52909 (I901611,I902140,I902089);
nand I_52910 (I901608,I902123,I902007);
not I_52911 (I902212,I2690);
DFFARX1 I_52912 (I815857,I2683,I902212,I902238,);
and I_52913 (I902246,I902238,I815854);
DFFARX1 I_52914 (I902246,I2683,I902212,I902195,);
DFFARX1 I_52915 (I815860,I2683,I902212,I902286,);
not I_52916 (I902294,I815863);
not I_52917 (I902311,I815857);
nand I_52918 (I902328,I902311,I902294);
nor I_52919 (I902183,I902286,I902328);
DFFARX1 I_52920 (I902328,I2683,I902212,I902368,);
not I_52921 (I902204,I902368);
not I_52922 (I902390,I815872);
nand I_52923 (I902407,I902311,I902390);
DFFARX1 I_52924 (I902407,I2683,I902212,I902433,);
not I_52925 (I902441,I902433);
not I_52926 (I902458,I815869);
nand I_52927 (I902475,I902458,I815875);
and I_52928 (I902492,I902294,I902475);
nor I_52929 (I902509,I902407,I902492);
DFFARX1 I_52930 (I902509,I2683,I902212,I902180,);
DFFARX1 I_52931 (I902492,I2683,I902212,I902201,);
nor I_52932 (I902554,I815869,I815854);
nor I_52933 (I902192,I902407,I902554);
or I_52934 (I902585,I815869,I815854);
nor I_52935 (I902602,I815866,I815860);
DFFARX1 I_52936 (I902602,I2683,I902212,I902628,);
not I_52937 (I902636,I902628);
nor I_52938 (I902198,I902636,I902441);
nand I_52939 (I902667,I902636,I902286);
not I_52940 (I902684,I815866);
nand I_52941 (I902701,I902684,I902390);
nand I_52942 (I902718,I902636,I902701);
nand I_52943 (I902189,I902718,I902667);
nand I_52944 (I902186,I902701,I902585);
not I_52945 (I902790,I2690);
DFFARX1 I_52946 (I788473,I2683,I902790,I902816,);
and I_52947 (I902824,I902816,I788467);
DFFARX1 I_52948 (I902824,I2683,I902790,I902773,);
DFFARX1 I_52949 (I788485,I2683,I902790,I902864,);
not I_52950 (I902872,I788476);
not I_52951 (I902889,I788488);
nand I_52952 (I902906,I902889,I902872);
nor I_52953 (I902761,I902864,I902906);
DFFARX1 I_52954 (I902906,I2683,I902790,I902946,);
not I_52955 (I902782,I902946);
not I_52956 (I902968,I788494);
nand I_52957 (I902985,I902889,I902968);
DFFARX1 I_52958 (I902985,I2683,I902790,I903011,);
not I_52959 (I903019,I903011);
not I_52960 (I903036,I788470);
nand I_52961 (I903053,I903036,I788491);
and I_52962 (I903070,I902872,I903053);
nor I_52963 (I903087,I902985,I903070);
DFFARX1 I_52964 (I903087,I2683,I902790,I902758,);
DFFARX1 I_52965 (I903070,I2683,I902790,I902779,);
nor I_52966 (I903132,I788470,I788482);
nor I_52967 (I902770,I902985,I903132);
or I_52968 (I903163,I788470,I788482);
nor I_52969 (I903180,I788467,I788479);
DFFARX1 I_52970 (I903180,I2683,I902790,I903206,);
not I_52971 (I903214,I903206);
nor I_52972 (I902776,I903214,I903019);
nand I_52973 (I903245,I903214,I902864);
not I_52974 (I903262,I788467);
nand I_52975 (I903279,I903262,I902968);
nand I_52976 (I903296,I903214,I903279);
nand I_52977 (I902767,I903296,I903245);
nand I_52978 (I902764,I903279,I903163);
not I_52979 (I903368,I2690);
DFFARX1 I_52980 (I335026,I2683,I903368,I903394,);
and I_52981 (I903402,I903394,I335041);
DFFARX1 I_52982 (I903402,I2683,I903368,I903351,);
DFFARX1 I_52983 (I335044,I2683,I903368,I903442,);
not I_52984 (I903450,I335038);
not I_52985 (I903467,I335053);
nand I_52986 (I903484,I903467,I903450);
nor I_52987 (I903339,I903442,I903484);
DFFARX1 I_52988 (I903484,I2683,I903368,I903524,);
not I_52989 (I903360,I903524);
not I_52990 (I903546,I335029);
nand I_52991 (I903563,I903467,I903546);
DFFARX1 I_52992 (I903563,I2683,I903368,I903589,);
not I_52993 (I903597,I903589);
not I_52994 (I903614,I335032);
nand I_52995 (I903631,I903614,I335026);
and I_52996 (I903648,I903450,I903631);
nor I_52997 (I903665,I903563,I903648);
DFFARX1 I_52998 (I903665,I2683,I903368,I903336,);
DFFARX1 I_52999 (I903648,I2683,I903368,I903357,);
nor I_53000 (I903710,I335032,I335035);
nor I_53001 (I903348,I903563,I903710);
or I_53002 (I903741,I335032,I335035);
nor I_53003 (I903758,I335050,I335047);
DFFARX1 I_53004 (I903758,I2683,I903368,I903784,);
not I_53005 (I903792,I903784);
nor I_53006 (I903354,I903792,I903597);
nand I_53007 (I903823,I903792,I903442);
not I_53008 (I903840,I335050);
nand I_53009 (I903857,I903840,I903546);
nand I_53010 (I903874,I903792,I903857);
nand I_53011 (I903345,I903874,I903823);
nand I_53012 (I903342,I903857,I903741);
not I_53013 (I903946,I2690);
DFFARX1 I_53014 (I967923,I2683,I903946,I903972,);
and I_53015 (I903980,I903972,I967917);
DFFARX1 I_53016 (I903980,I2683,I903946,I903929,);
DFFARX1 I_53017 (I967902,I2683,I903946,I904020,);
not I_53018 (I904028,I967908);
not I_53019 (I904045,I967920);
nand I_53020 (I904062,I904045,I904028);
nor I_53021 (I903917,I904020,I904062);
DFFARX1 I_53022 (I904062,I2683,I903946,I904102,);
not I_53023 (I903938,I904102);
not I_53024 (I904124,I967902);
nand I_53025 (I904141,I904045,I904124);
DFFARX1 I_53026 (I904141,I2683,I903946,I904167,);
not I_53027 (I904175,I904167);
not I_53028 (I904192,I967926);
nand I_53029 (I904209,I904192,I967914);
and I_53030 (I904226,I904028,I904209);
nor I_53031 (I904243,I904141,I904226);
DFFARX1 I_53032 (I904243,I2683,I903946,I903914,);
DFFARX1 I_53033 (I904226,I2683,I903946,I903935,);
nor I_53034 (I904288,I967926,I967905);
nor I_53035 (I903926,I904141,I904288);
or I_53036 (I904319,I967926,I967905);
nor I_53037 (I904336,I967911,I967905);
DFFARX1 I_53038 (I904336,I2683,I903946,I904362,);
not I_53039 (I904370,I904362);
nor I_53040 (I903932,I904370,I904175);
nand I_53041 (I904401,I904370,I904020);
not I_53042 (I904418,I967911);
nand I_53043 (I904435,I904418,I904124);
nand I_53044 (I904452,I904370,I904435);
nand I_53045 (I903923,I904452,I904401);
nand I_53046 (I903920,I904435,I904319);
not I_53047 (I904524,I2690);
DFFARX1 I_53048 (I671799,I2683,I904524,I904550,);
and I_53049 (I904558,I904550,I671805);
DFFARX1 I_53050 (I904558,I2683,I904524,I904507,);
DFFARX1 I_53051 (I671811,I2683,I904524,I904598,);
not I_53052 (I904606,I671796);
not I_53053 (I904623,I671796);
nand I_53054 (I904640,I904623,I904606);
nor I_53055 (I904495,I904598,I904640);
DFFARX1 I_53056 (I904640,I2683,I904524,I904680,);
not I_53057 (I904516,I904680);
not I_53058 (I904702,I671814);
nand I_53059 (I904719,I904623,I904702);
DFFARX1 I_53060 (I904719,I2683,I904524,I904745,);
not I_53061 (I904753,I904745);
not I_53062 (I904770,I671808);
nand I_53063 (I904787,I904770,I671799);
and I_53064 (I904804,I904606,I904787);
nor I_53065 (I904821,I904719,I904804);
DFFARX1 I_53066 (I904821,I2683,I904524,I904492,);
DFFARX1 I_53067 (I904804,I2683,I904524,I904513,);
nor I_53068 (I904866,I671808,I671817);
nor I_53069 (I904504,I904719,I904866);
or I_53070 (I904897,I671808,I671817);
nor I_53071 (I904914,I671802,I671802);
DFFARX1 I_53072 (I904914,I2683,I904524,I904940,);
not I_53073 (I904948,I904940);
nor I_53074 (I904510,I904948,I904753);
nand I_53075 (I904979,I904948,I904598);
not I_53076 (I904996,I671802);
nand I_53077 (I905013,I904996,I904702);
nand I_53078 (I905030,I904948,I905013);
nand I_53079 (I904501,I905030,I904979);
nand I_53080 (I904498,I905013,I904897);
not I_53081 (I905102,I2690);
DFFARX1 I_53082 (I128935,I2683,I905102,I905128,);
and I_53083 (I905136,I905128,I128938);
DFFARX1 I_53084 (I905136,I2683,I905102,I905085,);
DFFARX1 I_53085 (I128938,I2683,I905102,I905176,);
not I_53086 (I905184,I128953);
not I_53087 (I905201,I128959);
nand I_53088 (I905218,I905201,I905184);
nor I_53089 (I905073,I905176,I905218);
DFFARX1 I_53090 (I905218,I2683,I905102,I905258,);
not I_53091 (I905094,I905258);
not I_53092 (I905280,I128947);
nand I_53093 (I905297,I905201,I905280);
DFFARX1 I_53094 (I905297,I2683,I905102,I905323,);
not I_53095 (I905331,I905323);
not I_53096 (I905348,I128944);
nand I_53097 (I905365,I905348,I128941);
and I_53098 (I905382,I905184,I905365);
nor I_53099 (I905399,I905297,I905382);
DFFARX1 I_53100 (I905399,I2683,I905102,I905070,);
DFFARX1 I_53101 (I905382,I2683,I905102,I905091,);
nor I_53102 (I905444,I128944,I128935);
nor I_53103 (I905082,I905297,I905444);
or I_53104 (I905475,I128944,I128935);
nor I_53105 (I905492,I128950,I128956);
DFFARX1 I_53106 (I905492,I2683,I905102,I905518,);
not I_53107 (I905526,I905518);
nor I_53108 (I905088,I905526,I905331);
nand I_53109 (I905557,I905526,I905176);
not I_53110 (I905574,I128950);
nand I_53111 (I905591,I905574,I905280);
nand I_53112 (I905608,I905526,I905591);
nand I_53113 (I905079,I905608,I905557);
nand I_53114 (I905076,I905591,I905475);
not I_53115 (I905680,I2690);
DFFARX1 I_53116 (I547439,I2683,I905680,I905706,);
and I_53117 (I905714,I905706,I547427);
DFFARX1 I_53118 (I905714,I2683,I905680,I905663,);
DFFARX1 I_53119 (I547430,I2683,I905680,I905754,);
not I_53120 (I905762,I547424);
not I_53121 (I905779,I547448);
nand I_53122 (I905796,I905779,I905762);
nor I_53123 (I905651,I905754,I905796);
DFFARX1 I_53124 (I905796,I2683,I905680,I905836,);
not I_53125 (I905672,I905836);
not I_53126 (I905858,I547436);
nand I_53127 (I905875,I905779,I905858);
DFFARX1 I_53128 (I905875,I2683,I905680,I905901,);
not I_53129 (I905909,I905901);
not I_53130 (I905926,I547445);
nand I_53131 (I905943,I905926,I547442);
and I_53132 (I905960,I905762,I905943);
nor I_53133 (I905977,I905875,I905960);
DFFARX1 I_53134 (I905977,I2683,I905680,I905648,);
DFFARX1 I_53135 (I905960,I2683,I905680,I905669,);
nor I_53136 (I906022,I547445,I547433);
nor I_53137 (I905660,I905875,I906022);
or I_53138 (I906053,I547445,I547433);
nor I_53139 (I906070,I547424,I547427);
DFFARX1 I_53140 (I906070,I2683,I905680,I906096,);
not I_53141 (I906104,I906096);
nor I_53142 (I905666,I906104,I905909);
nand I_53143 (I906135,I906104,I905754);
not I_53144 (I906152,I547424);
nand I_53145 (I906169,I906152,I905858);
nand I_53146 (I906186,I906104,I906169);
nand I_53147 (I905657,I906186,I906135);
nand I_53148 (I905654,I906169,I906053);
not I_53149 (I906258,I2690);
DFFARX1 I_53150 (I688136,I2683,I906258,I906284,);
and I_53151 (I906292,I906284,I688142);
DFFARX1 I_53152 (I906292,I2683,I906258,I906241,);
DFFARX1 I_53153 (I688148,I2683,I906258,I906332,);
not I_53154 (I906340,I688133);
not I_53155 (I906357,I688133);
nand I_53156 (I906374,I906357,I906340);
nor I_53157 (I906229,I906332,I906374);
DFFARX1 I_53158 (I906374,I2683,I906258,I906414,);
not I_53159 (I906250,I906414);
not I_53160 (I906436,I688151);
nand I_53161 (I906453,I906357,I906436);
DFFARX1 I_53162 (I906453,I2683,I906258,I906479,);
not I_53163 (I906487,I906479);
not I_53164 (I906504,I688145);
nand I_53165 (I906521,I906504,I688136);
and I_53166 (I906538,I906340,I906521);
nor I_53167 (I906555,I906453,I906538);
DFFARX1 I_53168 (I906555,I2683,I906258,I906226,);
DFFARX1 I_53169 (I906538,I2683,I906258,I906247,);
nor I_53170 (I906600,I688145,I688154);
nor I_53171 (I906238,I906453,I906600);
or I_53172 (I906631,I688145,I688154);
nor I_53173 (I906648,I688139,I688139);
DFFARX1 I_53174 (I906648,I2683,I906258,I906674,);
not I_53175 (I906682,I906674);
nor I_53176 (I906244,I906682,I906487);
nand I_53177 (I906713,I906682,I906332);
not I_53178 (I906730,I688139);
nand I_53179 (I906747,I906730,I906436);
nand I_53180 (I906764,I906682,I906747);
nand I_53181 (I906235,I906764,I906713);
nand I_53182 (I906232,I906747,I906631);
not I_53183 (I906836,I2690);
DFFARX1 I_53184 (I664421,I2683,I906836,I906862,);
and I_53185 (I906870,I906862,I664427);
DFFARX1 I_53186 (I906870,I2683,I906836,I906819,);
DFFARX1 I_53187 (I664433,I2683,I906836,I906910,);
not I_53188 (I906918,I664418);
not I_53189 (I906935,I664418);
nand I_53190 (I906952,I906935,I906918);
nor I_53191 (I906807,I906910,I906952);
DFFARX1 I_53192 (I906952,I2683,I906836,I906992,);
not I_53193 (I906828,I906992);
not I_53194 (I907014,I664436);
nand I_53195 (I907031,I906935,I907014);
DFFARX1 I_53196 (I907031,I2683,I906836,I907057,);
not I_53197 (I907065,I907057);
not I_53198 (I907082,I664430);
nand I_53199 (I907099,I907082,I664421);
and I_53200 (I907116,I906918,I907099);
nor I_53201 (I907133,I907031,I907116);
DFFARX1 I_53202 (I907133,I2683,I906836,I906804,);
DFFARX1 I_53203 (I907116,I2683,I906836,I906825,);
nor I_53204 (I907178,I664430,I664439);
nor I_53205 (I906816,I907031,I907178);
or I_53206 (I907209,I664430,I664439);
nor I_53207 (I907226,I664424,I664424);
DFFARX1 I_53208 (I907226,I2683,I906836,I907252,);
not I_53209 (I907260,I907252);
nor I_53210 (I906822,I907260,I907065);
nand I_53211 (I907291,I907260,I906910);
not I_53212 (I907308,I664424);
nand I_53213 (I907325,I907308,I907014);
nand I_53214 (I907342,I907260,I907325);
nand I_53215 (I906813,I907342,I907291);
nand I_53216 (I906810,I907325,I907209);
not I_53217 (I907414,I2690);
DFFARX1 I_53218 (I621734,I2683,I907414,I907440,);
and I_53219 (I907448,I907440,I621740);
DFFARX1 I_53220 (I907448,I2683,I907414,I907397,);
DFFARX1 I_53221 (I621746,I2683,I907414,I907488,);
not I_53222 (I907496,I621731);
not I_53223 (I907513,I621731);
nand I_53224 (I907530,I907513,I907496);
nor I_53225 (I907385,I907488,I907530);
DFFARX1 I_53226 (I907530,I2683,I907414,I907570,);
not I_53227 (I907406,I907570);
not I_53228 (I907592,I621749);
nand I_53229 (I907609,I907513,I907592);
DFFARX1 I_53230 (I907609,I2683,I907414,I907635,);
not I_53231 (I907643,I907635);
not I_53232 (I907660,I621743);
nand I_53233 (I907677,I907660,I621734);
and I_53234 (I907694,I907496,I907677);
nor I_53235 (I907711,I907609,I907694);
DFFARX1 I_53236 (I907711,I2683,I907414,I907382,);
DFFARX1 I_53237 (I907694,I2683,I907414,I907403,);
nor I_53238 (I907756,I621743,I621752);
nor I_53239 (I907394,I907609,I907756);
or I_53240 (I907787,I621743,I621752);
nor I_53241 (I907804,I621737,I621737);
DFFARX1 I_53242 (I907804,I2683,I907414,I907830,);
not I_53243 (I907838,I907830);
nor I_53244 (I907400,I907838,I907643);
nand I_53245 (I907869,I907838,I907488);
not I_53246 (I907886,I621737);
nand I_53247 (I907903,I907886,I907592);
nand I_53248 (I907920,I907838,I907903);
nand I_53249 (I907391,I907920,I907869);
nand I_53250 (I907388,I907903,I907787);
not I_53251 (I907992,I2690);
DFFARX1 I_53252 (I400870,I2683,I907992,I908018,);
and I_53253 (I908026,I908018,I400885);
DFFARX1 I_53254 (I908026,I2683,I907992,I907975,);
DFFARX1 I_53255 (I400876,I2683,I907992,I908066,);
not I_53256 (I908074,I400870);
not I_53257 (I908091,I400888);
nand I_53258 (I908108,I908091,I908074);
nor I_53259 (I907963,I908066,I908108);
DFFARX1 I_53260 (I908108,I2683,I907992,I908148,);
not I_53261 (I907984,I908148);
not I_53262 (I908170,I400879);
nand I_53263 (I908187,I908091,I908170);
DFFARX1 I_53264 (I908187,I2683,I907992,I908213,);
not I_53265 (I908221,I908213);
not I_53266 (I908238,I400891);
nand I_53267 (I908255,I908238,I400867);
and I_53268 (I908272,I908074,I908255);
nor I_53269 (I908289,I908187,I908272);
DFFARX1 I_53270 (I908289,I2683,I907992,I907960,);
DFFARX1 I_53271 (I908272,I2683,I907992,I907981,);
nor I_53272 (I908334,I400891,I400867);
nor I_53273 (I907972,I908187,I908334);
or I_53274 (I908365,I400891,I400867);
nor I_53275 (I908382,I400873,I400882);
DFFARX1 I_53276 (I908382,I2683,I907992,I908408,);
not I_53277 (I908416,I908408);
nor I_53278 (I907978,I908416,I908221);
nand I_53279 (I908447,I908416,I908066);
not I_53280 (I908464,I400873);
nand I_53281 (I908481,I908464,I908170);
nand I_53282 (I908498,I908416,I908481);
nand I_53283 (I907969,I908498,I908447);
nand I_53284 (I907966,I908481,I908365);
not I_53285 (I908570,I2690);
DFFARX1 I_53286 (I8063,I2683,I908570,I908596,);
and I_53287 (I908604,I908596,I8069);
DFFARX1 I_53288 (I908604,I2683,I908570,I908553,);
DFFARX1 I_53289 (I8048,I2683,I908570,I908644,);
not I_53290 (I908652,I8054);
not I_53291 (I908669,I8060);
nand I_53292 (I908686,I908669,I908652);
nor I_53293 (I908541,I908644,I908686);
DFFARX1 I_53294 (I908686,I2683,I908570,I908726,);
not I_53295 (I908562,I908726);
not I_53296 (I908748,I8051);
nand I_53297 (I908765,I908669,I908748);
DFFARX1 I_53298 (I908765,I2683,I908570,I908791,);
not I_53299 (I908799,I908791);
not I_53300 (I908816,I8066);
nand I_53301 (I908833,I908816,I8051);
and I_53302 (I908850,I908652,I908833);
nor I_53303 (I908867,I908765,I908850);
DFFARX1 I_53304 (I908867,I2683,I908570,I908538,);
DFFARX1 I_53305 (I908850,I2683,I908570,I908559,);
nor I_53306 (I908912,I8066,I8054);
nor I_53307 (I908550,I908765,I908912);
or I_53308 (I908943,I8066,I8054);
nor I_53309 (I908960,I8057,I8048);
DFFARX1 I_53310 (I908960,I2683,I908570,I908986,);
not I_53311 (I908994,I908986);
nor I_53312 (I908556,I908994,I908799);
nand I_53313 (I909025,I908994,I908644);
not I_53314 (I909042,I8057);
nand I_53315 (I909059,I909042,I908748);
nand I_53316 (I909076,I908994,I909059);
nand I_53317 (I908547,I909076,I909025);
nand I_53318 (I908544,I909059,I908943);
not I_53319 (I909148,I2690);
DFFARX1 I_53320 (I53275,I2683,I909148,I909174,);
and I_53321 (I909182,I909174,I53251);
DFFARX1 I_53322 (I909182,I2683,I909148,I909131,);
DFFARX1 I_53323 (I53269,I2683,I909148,I909222,);
not I_53324 (I909230,I53257);
not I_53325 (I909247,I53254);
nand I_53326 (I909264,I909247,I909230);
nor I_53327 (I909119,I909222,I909264);
DFFARX1 I_53328 (I909264,I2683,I909148,I909304,);
not I_53329 (I909140,I909304);
not I_53330 (I909326,I53263);
nand I_53331 (I909343,I909247,I909326);
DFFARX1 I_53332 (I909343,I2683,I909148,I909369,);
not I_53333 (I909377,I909369);
not I_53334 (I909394,I53254);
nand I_53335 (I909411,I909394,I53272);
and I_53336 (I909428,I909230,I909411);
nor I_53337 (I909445,I909343,I909428);
DFFARX1 I_53338 (I909445,I2683,I909148,I909116,);
DFFARX1 I_53339 (I909428,I2683,I909148,I909137,);
nor I_53340 (I909490,I53254,I53266);
nor I_53341 (I909128,I909343,I909490);
or I_53342 (I909521,I53254,I53266);
nor I_53343 (I909538,I53260,I53251);
DFFARX1 I_53344 (I909538,I2683,I909148,I909564,);
not I_53345 (I909572,I909564);
nor I_53346 (I909134,I909572,I909377);
nand I_53347 (I909603,I909572,I909222);
not I_53348 (I909620,I53260);
nand I_53349 (I909637,I909620,I909326);
nand I_53350 (I909654,I909572,I909637);
nand I_53351 (I909125,I909654,I909603);
nand I_53352 (I909122,I909637,I909521);
not I_53353 (I909726,I2690);
DFFARX1 I_53354 (I798466,I2683,I909726,I909752,);
and I_53355 (I909760,I909752,I798463);
DFFARX1 I_53356 (I909760,I2683,I909726,I909709,);
DFFARX1 I_53357 (I798469,I2683,I909726,I909800,);
not I_53358 (I909808,I798472);
not I_53359 (I909825,I798466);
nand I_53360 (I909842,I909825,I909808);
nor I_53361 (I909697,I909800,I909842);
DFFARX1 I_53362 (I909842,I2683,I909726,I909882,);
not I_53363 (I909718,I909882);
not I_53364 (I909904,I798481);
nand I_53365 (I909921,I909825,I909904);
DFFARX1 I_53366 (I909921,I2683,I909726,I909947,);
not I_53367 (I909955,I909947);
not I_53368 (I909972,I798478);
nand I_53369 (I909989,I909972,I798484);
and I_53370 (I910006,I909808,I909989);
nor I_53371 (I910023,I909921,I910006);
DFFARX1 I_53372 (I910023,I2683,I909726,I909694,);
DFFARX1 I_53373 (I910006,I2683,I909726,I909715,);
nor I_53374 (I910068,I798478,I798463);
nor I_53375 (I909706,I909921,I910068);
or I_53376 (I910099,I798478,I798463);
nor I_53377 (I910116,I798475,I798469);
DFFARX1 I_53378 (I910116,I2683,I909726,I910142,);
not I_53379 (I910150,I910142);
nor I_53380 (I909712,I910150,I909955);
nand I_53381 (I910181,I910150,I909800);
not I_53382 (I910198,I798475);
nand I_53383 (I910215,I910198,I909904);
nand I_53384 (I910232,I910150,I910215);
nand I_53385 (I909703,I910232,I910181);
nand I_53386 (I909700,I910215,I910099);
not I_53387 (I910304,I2690);
DFFARX1 I_53388 (I969011,I2683,I910304,I910330,);
and I_53389 (I910338,I910330,I969005);
DFFARX1 I_53390 (I910338,I2683,I910304,I910287,);
DFFARX1 I_53391 (I968990,I2683,I910304,I910378,);
not I_53392 (I910386,I968996);
not I_53393 (I910403,I969008);
nand I_53394 (I910420,I910403,I910386);
nor I_53395 (I910275,I910378,I910420);
DFFARX1 I_53396 (I910420,I2683,I910304,I910460,);
not I_53397 (I910296,I910460);
not I_53398 (I910482,I968990);
nand I_53399 (I910499,I910403,I910482);
DFFARX1 I_53400 (I910499,I2683,I910304,I910525,);
not I_53401 (I910533,I910525);
not I_53402 (I910550,I969014);
nand I_53403 (I910567,I910550,I969002);
and I_53404 (I910584,I910386,I910567);
nor I_53405 (I910601,I910499,I910584);
DFFARX1 I_53406 (I910601,I2683,I910304,I910272,);
DFFARX1 I_53407 (I910584,I2683,I910304,I910293,);
nor I_53408 (I910646,I969014,I968993);
nor I_53409 (I910284,I910499,I910646);
or I_53410 (I910677,I969014,I968993);
nor I_53411 (I910694,I968999,I968993);
DFFARX1 I_53412 (I910694,I2683,I910304,I910720,);
not I_53413 (I910728,I910720);
nor I_53414 (I910290,I910728,I910533);
nand I_53415 (I910759,I910728,I910378);
not I_53416 (I910776,I968999);
nand I_53417 (I910793,I910776,I910482);
nand I_53418 (I910810,I910728,I910793);
nand I_53419 (I910281,I910810,I910759);
nand I_53420 (I910278,I910793,I910677);
not I_53421 (I910882,I2690);
DFFARX1 I_53422 (I403250,I2683,I910882,I910908,);
and I_53423 (I910916,I910908,I403265);
DFFARX1 I_53424 (I910916,I2683,I910882,I910865,);
DFFARX1 I_53425 (I403256,I2683,I910882,I910956,);
not I_53426 (I910964,I403250);
not I_53427 (I910981,I403268);
nand I_53428 (I910998,I910981,I910964);
nor I_53429 (I910853,I910956,I910998);
DFFARX1 I_53430 (I910998,I2683,I910882,I911038,);
not I_53431 (I910874,I911038);
not I_53432 (I911060,I403259);
nand I_53433 (I911077,I910981,I911060);
DFFARX1 I_53434 (I911077,I2683,I910882,I911103,);
not I_53435 (I911111,I911103);
not I_53436 (I911128,I403271);
nand I_53437 (I911145,I911128,I403247);
and I_53438 (I911162,I910964,I911145);
nor I_53439 (I911179,I911077,I911162);
DFFARX1 I_53440 (I911179,I2683,I910882,I910850,);
DFFARX1 I_53441 (I911162,I2683,I910882,I910871,);
nor I_53442 (I911224,I403271,I403247);
nor I_53443 (I910862,I911077,I911224);
or I_53444 (I911255,I403271,I403247);
nor I_53445 (I911272,I403253,I403262);
DFFARX1 I_53446 (I911272,I2683,I910882,I911298,);
not I_53447 (I911306,I911298);
nor I_53448 (I910868,I911306,I911111);
nand I_53449 (I911337,I911306,I910956);
not I_53450 (I911354,I403253);
nand I_53451 (I911371,I911354,I911060);
nand I_53452 (I911388,I911306,I911371);
nand I_53453 (I910859,I911388,I911337);
nand I_53454 (I910856,I911371,I911255);
not I_53455 (I911460,I2690);
DFFARX1 I_53456 (I401465,I2683,I911460,I911486,);
and I_53457 (I911494,I911486,I401480);
DFFARX1 I_53458 (I911494,I2683,I911460,I911443,);
DFFARX1 I_53459 (I401471,I2683,I911460,I911534,);
not I_53460 (I911542,I401465);
not I_53461 (I911559,I401483);
nand I_53462 (I911576,I911559,I911542);
nor I_53463 (I911431,I911534,I911576);
DFFARX1 I_53464 (I911576,I2683,I911460,I911616,);
not I_53465 (I911452,I911616);
not I_53466 (I911638,I401474);
nand I_53467 (I911655,I911559,I911638);
DFFARX1 I_53468 (I911655,I2683,I911460,I911681,);
not I_53469 (I911689,I911681);
not I_53470 (I911706,I401486);
nand I_53471 (I911723,I911706,I401462);
and I_53472 (I911740,I911542,I911723);
nor I_53473 (I911757,I911655,I911740);
DFFARX1 I_53474 (I911757,I2683,I911460,I911428,);
DFFARX1 I_53475 (I911740,I2683,I911460,I911449,);
nor I_53476 (I911802,I401486,I401462);
nor I_53477 (I911440,I911655,I911802);
or I_53478 (I911833,I401486,I401462);
nor I_53479 (I911850,I401468,I401477);
DFFARX1 I_53480 (I911850,I2683,I911460,I911876,);
not I_53481 (I911884,I911876);
nor I_53482 (I911446,I911884,I911689);
nand I_53483 (I911915,I911884,I911534);
not I_53484 (I911932,I401468);
nand I_53485 (I911949,I911932,I911638);
nand I_53486 (I911966,I911884,I911949);
nand I_53487 (I911437,I911966,I911915);
nand I_53488 (I911434,I911949,I911833);
not I_53489 (I912038,I2690);
DFFARX1 I_53490 (I44292,I2683,I912038,I912064,);
and I_53491 (I912072,I912064,I44295);
DFFARX1 I_53492 (I912072,I2683,I912038,I912021,);
DFFARX1 I_53493 (I44295,I2683,I912038,I912112,);
not I_53494 (I912120,I44298);
not I_53495 (I912137,I44313);
nand I_53496 (I912154,I912137,I912120);
nor I_53497 (I912009,I912112,I912154);
DFFARX1 I_53498 (I912154,I2683,I912038,I912194,);
not I_53499 (I912030,I912194);
not I_53500 (I912216,I44307);
nand I_53501 (I912233,I912137,I912216);
DFFARX1 I_53502 (I912233,I2683,I912038,I912259,);
not I_53503 (I912267,I912259);
not I_53504 (I912284,I44310);
nand I_53505 (I912301,I912284,I44292);
and I_53506 (I912318,I912120,I912301);
nor I_53507 (I912335,I912233,I912318);
DFFARX1 I_53508 (I912335,I2683,I912038,I912006,);
DFFARX1 I_53509 (I912318,I2683,I912038,I912027,);
nor I_53510 (I912380,I44310,I44304);
nor I_53511 (I912018,I912233,I912380);
or I_53512 (I912411,I44310,I44304);
nor I_53513 (I912428,I44301,I44316);
DFFARX1 I_53514 (I912428,I2683,I912038,I912454,);
not I_53515 (I912462,I912454);
nor I_53516 (I912024,I912462,I912267);
nand I_53517 (I912493,I912462,I912112);
not I_53518 (I912510,I44301);
nand I_53519 (I912527,I912510,I912216);
nand I_53520 (I912544,I912462,I912527);
nand I_53521 (I912015,I912544,I912493);
nand I_53522 (I912012,I912527,I912411);
not I_53523 (I912616,I2690);
DFFARX1 I_53524 (I381810,I2683,I912616,I912642,);
and I_53525 (I912650,I912642,I381825);
DFFARX1 I_53526 (I912650,I2683,I912616,I912599,);
DFFARX1 I_53527 (I381828,I2683,I912616,I912690,);
not I_53528 (I912698,I381822);
not I_53529 (I912715,I381837);
nand I_53530 (I912732,I912715,I912698);
nor I_53531 (I912587,I912690,I912732);
DFFARX1 I_53532 (I912732,I2683,I912616,I912772,);
not I_53533 (I912608,I912772);
not I_53534 (I912794,I381813);
nand I_53535 (I912811,I912715,I912794);
DFFARX1 I_53536 (I912811,I2683,I912616,I912837,);
not I_53537 (I912845,I912837);
not I_53538 (I912862,I381816);
nand I_53539 (I912879,I912862,I381810);
and I_53540 (I912896,I912698,I912879);
nor I_53541 (I912913,I912811,I912896);
DFFARX1 I_53542 (I912913,I2683,I912616,I912584,);
DFFARX1 I_53543 (I912896,I2683,I912616,I912605,);
nor I_53544 (I912958,I381816,I381819);
nor I_53545 (I912596,I912811,I912958);
or I_53546 (I912989,I381816,I381819);
nor I_53547 (I913006,I381834,I381831);
DFFARX1 I_53548 (I913006,I2683,I912616,I913032,);
not I_53549 (I913040,I913032);
nor I_53550 (I912602,I913040,I912845);
nand I_53551 (I913071,I913040,I912690);
not I_53552 (I913088,I381834);
nand I_53553 (I913105,I913088,I912794);
nand I_53554 (I913122,I913040,I913105);
nand I_53555 (I912593,I913122,I913071);
nand I_53556 (I912590,I913105,I912989);
not I_53557 (I913194,I2690);
DFFARX1 I_53558 (I993800,I2683,I913194,I913220,);
and I_53559 (I913228,I913220,I993782);
DFFARX1 I_53560 (I913228,I2683,I913194,I913177,);
DFFARX1 I_53561 (I993791,I2683,I913194,I913268,);
not I_53562 (I913276,I993776);
not I_53563 (I913293,I993788);
nand I_53564 (I913310,I913293,I913276);
nor I_53565 (I913165,I913268,I913310);
DFFARX1 I_53566 (I913310,I2683,I913194,I913350,);
not I_53567 (I913186,I913350);
not I_53568 (I913372,I993779);
nand I_53569 (I913389,I913293,I913372);
DFFARX1 I_53570 (I913389,I2683,I913194,I913415,);
not I_53571 (I913423,I913415);
not I_53572 (I913440,I993776);
nand I_53573 (I913457,I913440,I993779);
and I_53574 (I913474,I913276,I913457);
nor I_53575 (I913491,I913389,I913474);
DFFARX1 I_53576 (I913491,I2683,I913194,I913162,);
DFFARX1 I_53577 (I913474,I2683,I913194,I913183,);
nor I_53578 (I913536,I993776,I993797);
nor I_53579 (I913174,I913389,I913536);
or I_53580 (I913567,I993776,I993797);
nor I_53581 (I913584,I993785,I993794);
DFFARX1 I_53582 (I913584,I2683,I913194,I913610,);
not I_53583 (I913618,I913610);
nor I_53584 (I913180,I913618,I913423);
nand I_53585 (I913649,I913618,I913268);
not I_53586 (I913666,I993785);
nand I_53587 (I913683,I913666,I913372);
nand I_53588 (I913700,I913618,I913683);
nand I_53589 (I913171,I913700,I913649);
nand I_53590 (I913168,I913683,I913567);
not I_53591 (I913772,I2690);
DFFARX1 I_53592 (I300203,I2683,I913772,I913798,);
and I_53593 (I913806,I913798,I300188);
DFFARX1 I_53594 (I913806,I2683,I913772,I913755,);
DFFARX1 I_53595 (I300194,I2683,I913772,I913846,);
not I_53596 (I913854,I300176);
not I_53597 (I913871,I300197);
nand I_53598 (I913888,I913871,I913854);
nor I_53599 (I913743,I913846,I913888);
DFFARX1 I_53600 (I913888,I2683,I913772,I913928,);
not I_53601 (I913764,I913928);
not I_53602 (I913950,I300200);
nand I_53603 (I913967,I913871,I913950);
DFFARX1 I_53604 (I913967,I2683,I913772,I913993,);
not I_53605 (I914001,I913993);
not I_53606 (I914018,I300191);
nand I_53607 (I914035,I914018,I300179);
and I_53608 (I914052,I913854,I914035);
nor I_53609 (I914069,I913967,I914052);
DFFARX1 I_53610 (I914069,I2683,I913772,I913740,);
DFFARX1 I_53611 (I914052,I2683,I913772,I913761,);
nor I_53612 (I914114,I300191,I300185);
nor I_53613 (I913752,I913967,I914114);
or I_53614 (I914145,I300191,I300185);
nor I_53615 (I914162,I300182,I300176);
DFFARX1 I_53616 (I914162,I2683,I913772,I914188,);
not I_53617 (I914196,I914188);
nor I_53618 (I913758,I914196,I914001);
nand I_53619 (I914227,I914196,I913846);
not I_53620 (I914244,I300182);
nand I_53621 (I914261,I914244,I913950);
nand I_53622 (I914278,I914196,I914261);
nand I_53623 (I913749,I914278,I914227);
nand I_53624 (I913746,I914261,I914145);
not I_53625 (I914350,I2690);
DFFARX1 I_53626 (I253827,I2683,I914350,I914376,);
and I_53627 (I914384,I914376,I253812);
DFFARX1 I_53628 (I914384,I2683,I914350,I914333,);
DFFARX1 I_53629 (I253818,I2683,I914350,I914424,);
not I_53630 (I914432,I253800);
not I_53631 (I914449,I253821);
nand I_53632 (I914466,I914449,I914432);
nor I_53633 (I914321,I914424,I914466);
DFFARX1 I_53634 (I914466,I2683,I914350,I914506,);
not I_53635 (I914342,I914506);
not I_53636 (I914528,I253824);
nand I_53637 (I914545,I914449,I914528);
DFFARX1 I_53638 (I914545,I2683,I914350,I914571,);
not I_53639 (I914579,I914571);
not I_53640 (I914596,I253815);
nand I_53641 (I914613,I914596,I253803);
and I_53642 (I914630,I914432,I914613);
nor I_53643 (I914647,I914545,I914630);
DFFARX1 I_53644 (I914647,I2683,I914350,I914318,);
DFFARX1 I_53645 (I914630,I2683,I914350,I914339,);
nor I_53646 (I914692,I253815,I253809);
nor I_53647 (I914330,I914545,I914692);
or I_53648 (I914723,I253815,I253809);
nor I_53649 (I914740,I253806,I253800);
DFFARX1 I_53650 (I914740,I2683,I914350,I914766,);
not I_53651 (I914774,I914766);
nor I_53652 (I914336,I914774,I914579);
nand I_53653 (I914805,I914774,I914424);
not I_53654 (I914822,I253806);
nand I_53655 (I914839,I914822,I914528);
nand I_53656 (I914856,I914774,I914839);
nand I_53657 (I914327,I914856,I914805);
nand I_53658 (I914324,I914839,I914723);
not I_53659 (I914928,I2690);
DFFARX1 I_53660 (I259624,I2683,I914928,I914954,);
and I_53661 (I914962,I914954,I259609);
DFFARX1 I_53662 (I914962,I2683,I914928,I914911,);
DFFARX1 I_53663 (I259615,I2683,I914928,I915002,);
not I_53664 (I915010,I259597);
not I_53665 (I915027,I259618);
nand I_53666 (I915044,I915027,I915010);
nor I_53667 (I914899,I915002,I915044);
DFFARX1 I_53668 (I915044,I2683,I914928,I915084,);
not I_53669 (I914920,I915084);
not I_53670 (I915106,I259621);
nand I_53671 (I915123,I915027,I915106);
DFFARX1 I_53672 (I915123,I2683,I914928,I915149,);
not I_53673 (I915157,I915149);
not I_53674 (I915174,I259612);
nand I_53675 (I915191,I915174,I259600);
and I_53676 (I915208,I915010,I915191);
nor I_53677 (I915225,I915123,I915208);
DFFARX1 I_53678 (I915225,I2683,I914928,I914896,);
DFFARX1 I_53679 (I915208,I2683,I914928,I914917,);
nor I_53680 (I915270,I259612,I259606);
nor I_53681 (I914908,I915123,I915270);
or I_53682 (I915301,I259612,I259606);
nor I_53683 (I915318,I259603,I259597);
DFFARX1 I_53684 (I915318,I2683,I914928,I915344,);
not I_53685 (I915352,I915344);
nor I_53686 (I914914,I915352,I915157);
nand I_53687 (I915383,I915352,I915002);
not I_53688 (I915400,I259603);
nand I_53689 (I915417,I915400,I915106);
nand I_53690 (I915434,I915352,I915417);
nand I_53691 (I914905,I915434,I915383);
nand I_53692 (I914902,I915417,I915301);
not I_53693 (I915506,I2690);
DFFARX1 I_53694 (I326322,I2683,I915506,I915532,);
and I_53695 (I915540,I915532,I326337);
DFFARX1 I_53696 (I915540,I2683,I915506,I915489,);
DFFARX1 I_53697 (I326340,I2683,I915506,I915580,);
not I_53698 (I915588,I326334);
not I_53699 (I915605,I326349);
nand I_53700 (I915622,I915605,I915588);
nor I_53701 (I915477,I915580,I915622);
DFFARX1 I_53702 (I915622,I2683,I915506,I915662,);
not I_53703 (I915498,I915662);
not I_53704 (I915684,I326325);
nand I_53705 (I915701,I915605,I915684);
DFFARX1 I_53706 (I915701,I2683,I915506,I915727,);
not I_53707 (I915735,I915727);
not I_53708 (I915752,I326328);
nand I_53709 (I915769,I915752,I326322);
and I_53710 (I915786,I915588,I915769);
nor I_53711 (I915803,I915701,I915786);
DFFARX1 I_53712 (I915803,I2683,I915506,I915474,);
DFFARX1 I_53713 (I915786,I2683,I915506,I915495,);
nor I_53714 (I915848,I326328,I326331);
nor I_53715 (I915486,I915701,I915848);
or I_53716 (I915879,I326328,I326331);
nor I_53717 (I915896,I326346,I326343);
DFFARX1 I_53718 (I915896,I2683,I915506,I915922,);
not I_53719 (I915930,I915922);
nor I_53720 (I915492,I915930,I915735);
nand I_53721 (I915961,I915930,I915580);
not I_53722 (I915978,I326346);
nand I_53723 (I915995,I915978,I915684);
nand I_53724 (I916012,I915930,I915995);
nand I_53725 (I915483,I916012,I915961);
nand I_53726 (I915480,I915995,I915879);
not I_53727 (I916084,I2690);
DFFARX1 I_53728 (I432417,I2683,I916084,I916110,);
and I_53729 (I916118,I916110,I432405);
DFFARX1 I_53730 (I916118,I2683,I916084,I916067,);
DFFARX1 I_53731 (I432420,I2683,I916084,I916158,);
not I_53732 (I916166,I432411);
not I_53733 (I916183,I432402);
nand I_53734 (I916200,I916183,I916166);
nor I_53735 (I916055,I916158,I916200);
DFFARX1 I_53736 (I916200,I2683,I916084,I916240,);
not I_53737 (I916076,I916240);
not I_53738 (I916262,I432408);
nand I_53739 (I916279,I916183,I916262);
DFFARX1 I_53740 (I916279,I2683,I916084,I916305,);
not I_53741 (I916313,I916305);
not I_53742 (I916330,I432423);
nand I_53743 (I916347,I916330,I432426);
and I_53744 (I916364,I916166,I916347);
nor I_53745 (I916381,I916279,I916364);
DFFARX1 I_53746 (I916381,I2683,I916084,I916052,);
DFFARX1 I_53747 (I916364,I2683,I916084,I916073,);
nor I_53748 (I916426,I432423,I432402);
nor I_53749 (I916064,I916279,I916426);
or I_53750 (I916457,I432423,I432402);
nor I_53751 (I916474,I432414,I432405);
DFFARX1 I_53752 (I916474,I2683,I916084,I916500,);
not I_53753 (I916508,I916500);
nor I_53754 (I916070,I916508,I916313);
nand I_53755 (I916539,I916508,I916158);
not I_53756 (I916556,I432414);
nand I_53757 (I916573,I916556,I916262);
nand I_53758 (I916590,I916508,I916573);
nand I_53759 (I916061,I916590,I916539);
nand I_53760 (I916058,I916573,I916457);
not I_53761 (I916662,I2690);
DFFARX1 I_53762 (I568825,I2683,I916662,I916688,);
and I_53763 (I916696,I916688,I568813);
DFFARX1 I_53764 (I916696,I2683,I916662,I916645,);
DFFARX1 I_53765 (I568816,I2683,I916662,I916736,);
not I_53766 (I916744,I568810);
not I_53767 (I916761,I568834);
nand I_53768 (I916778,I916761,I916744);
nor I_53769 (I916633,I916736,I916778);
DFFARX1 I_53770 (I916778,I2683,I916662,I916818,);
not I_53771 (I916654,I916818);
not I_53772 (I916840,I568822);
nand I_53773 (I916857,I916761,I916840);
DFFARX1 I_53774 (I916857,I2683,I916662,I916883,);
not I_53775 (I916891,I916883);
not I_53776 (I916908,I568831);
nand I_53777 (I916925,I916908,I568828);
and I_53778 (I916942,I916744,I916925);
nor I_53779 (I916959,I916857,I916942);
DFFARX1 I_53780 (I916959,I2683,I916662,I916630,);
DFFARX1 I_53781 (I916942,I2683,I916662,I916651,);
nor I_53782 (I917004,I568831,I568819);
nor I_53783 (I916642,I916857,I917004);
or I_53784 (I917035,I568831,I568819);
nor I_53785 (I917052,I568810,I568813);
DFFARX1 I_53786 (I917052,I2683,I916662,I917078,);
not I_53787 (I917086,I917078);
nor I_53788 (I916648,I917086,I916891);
nand I_53789 (I917117,I917086,I916736);
not I_53790 (I917134,I568810);
nand I_53791 (I917151,I917134,I916840);
nand I_53792 (I917168,I917086,I917151);
nand I_53793 (I916639,I917168,I917117);
nand I_53794 (I916636,I917151,I917035);
not I_53795 (I917240,I2690);
DFFARX1 I_53796 (I175940,I2683,I917240,I917266,);
and I_53797 (I917274,I917266,I175943);
DFFARX1 I_53798 (I917274,I2683,I917240,I917223,);
DFFARX1 I_53799 (I175943,I2683,I917240,I917314,);
not I_53800 (I917322,I175958);
not I_53801 (I917339,I175964);
nand I_53802 (I917356,I917339,I917322);
nor I_53803 (I917211,I917314,I917356);
DFFARX1 I_53804 (I917356,I2683,I917240,I917396,);
not I_53805 (I917232,I917396);
not I_53806 (I917418,I175952);
nand I_53807 (I917435,I917339,I917418);
DFFARX1 I_53808 (I917435,I2683,I917240,I917461,);
not I_53809 (I917469,I917461);
not I_53810 (I917486,I175949);
nand I_53811 (I917503,I917486,I175946);
and I_53812 (I917520,I917322,I917503);
nor I_53813 (I917537,I917435,I917520);
DFFARX1 I_53814 (I917537,I2683,I917240,I917208,);
DFFARX1 I_53815 (I917520,I2683,I917240,I917229,);
nor I_53816 (I917582,I175949,I175940);
nor I_53817 (I917220,I917435,I917582);
or I_53818 (I917613,I175949,I175940);
nor I_53819 (I917630,I175955,I175961);
DFFARX1 I_53820 (I917630,I2683,I917240,I917656,);
not I_53821 (I917664,I917656);
nor I_53822 (I917226,I917664,I917469);
nand I_53823 (I917695,I917664,I917314);
not I_53824 (I917712,I175955);
nand I_53825 (I917729,I917712,I917418);
nand I_53826 (I917746,I917664,I917729);
nand I_53827 (I917217,I917746,I917695);
nand I_53828 (I917214,I917729,I917613);
not I_53829 (I917818,I2690);
DFFARX1 I_53830 (I977171,I2683,I917818,I917844,);
and I_53831 (I917852,I917844,I977165);
DFFARX1 I_53832 (I917852,I2683,I917818,I917801,);
DFFARX1 I_53833 (I977150,I2683,I917818,I917892,);
not I_53834 (I917900,I977156);
not I_53835 (I917917,I977168);
nand I_53836 (I917934,I917917,I917900);
nor I_53837 (I917789,I917892,I917934);
DFFARX1 I_53838 (I917934,I2683,I917818,I917974,);
not I_53839 (I917810,I917974);
not I_53840 (I917996,I977150);
nand I_53841 (I918013,I917917,I917996);
DFFARX1 I_53842 (I918013,I2683,I917818,I918039,);
not I_53843 (I918047,I918039);
not I_53844 (I918064,I977174);
nand I_53845 (I918081,I918064,I977162);
and I_53846 (I918098,I917900,I918081);
nor I_53847 (I918115,I918013,I918098);
DFFARX1 I_53848 (I918115,I2683,I917818,I917786,);
DFFARX1 I_53849 (I918098,I2683,I917818,I917807,);
nor I_53850 (I918160,I977174,I977153);
nor I_53851 (I917798,I918013,I918160);
or I_53852 (I918191,I977174,I977153);
nor I_53853 (I918208,I977159,I977153);
DFFARX1 I_53854 (I918208,I2683,I917818,I918234,);
not I_53855 (I918242,I918234);
nor I_53856 (I917804,I918242,I918047);
nand I_53857 (I918273,I918242,I917892);
not I_53858 (I918290,I977159);
nand I_53859 (I918307,I918290,I917996);
nand I_53860 (I918324,I918242,I918307);
nand I_53861 (I917795,I918324,I918273);
nand I_53862 (I917792,I918307,I918191);
not I_53863 (I918396,I2690);
DFFARX1 I_53864 (I40076,I2683,I918396,I918422,);
and I_53865 (I918430,I918422,I40079);
DFFARX1 I_53866 (I918430,I2683,I918396,I918379,);
DFFARX1 I_53867 (I40079,I2683,I918396,I918470,);
not I_53868 (I918478,I40082);
not I_53869 (I918495,I40097);
nand I_53870 (I918512,I918495,I918478);
nor I_53871 (I918367,I918470,I918512);
DFFARX1 I_53872 (I918512,I2683,I918396,I918552,);
not I_53873 (I918388,I918552);
not I_53874 (I918574,I40091);
nand I_53875 (I918591,I918495,I918574);
DFFARX1 I_53876 (I918591,I2683,I918396,I918617,);
not I_53877 (I918625,I918617);
not I_53878 (I918642,I40094);
nand I_53879 (I918659,I918642,I40076);
and I_53880 (I918676,I918478,I918659);
nor I_53881 (I918693,I918591,I918676);
DFFARX1 I_53882 (I918693,I2683,I918396,I918364,);
DFFARX1 I_53883 (I918676,I2683,I918396,I918385,);
nor I_53884 (I918738,I40094,I40088);
nor I_53885 (I918376,I918591,I918738);
or I_53886 (I918769,I40094,I40088);
nor I_53887 (I918786,I40085,I40100);
DFFARX1 I_53888 (I918786,I2683,I918396,I918812,);
not I_53889 (I918820,I918812);
nor I_53890 (I918382,I918820,I918625);
nand I_53891 (I918851,I918820,I918470);
not I_53892 (I918868,I40085);
nand I_53893 (I918885,I918868,I918574);
nand I_53894 (I918902,I918820,I918885);
nand I_53895 (I918373,I918902,I918851);
nand I_53896 (I918370,I918885,I918769);
not I_53897 (I918974,I2690);
DFFARX1 I_53898 (I16888,I2683,I918974,I919000,);
and I_53899 (I919008,I919000,I16891);
DFFARX1 I_53900 (I919008,I2683,I918974,I918957,);
DFFARX1 I_53901 (I16891,I2683,I918974,I919048,);
not I_53902 (I919056,I16894);
not I_53903 (I919073,I16909);
nand I_53904 (I919090,I919073,I919056);
nor I_53905 (I918945,I919048,I919090);
DFFARX1 I_53906 (I919090,I2683,I918974,I919130,);
not I_53907 (I918966,I919130);
not I_53908 (I919152,I16903);
nand I_53909 (I919169,I919073,I919152);
DFFARX1 I_53910 (I919169,I2683,I918974,I919195,);
not I_53911 (I919203,I919195);
not I_53912 (I919220,I16906);
nand I_53913 (I919237,I919220,I16888);
and I_53914 (I919254,I919056,I919237);
nor I_53915 (I919271,I919169,I919254);
DFFARX1 I_53916 (I919271,I2683,I918974,I918942,);
DFFARX1 I_53917 (I919254,I2683,I918974,I918963,);
nor I_53918 (I919316,I16906,I16900);
nor I_53919 (I918954,I919169,I919316);
or I_53920 (I919347,I16906,I16900);
nor I_53921 (I919364,I16897,I16912);
DFFARX1 I_53922 (I919364,I2683,I918974,I919390,);
not I_53923 (I919398,I919390);
nor I_53924 (I918960,I919398,I919203);
nand I_53925 (I919429,I919398,I919048);
not I_53926 (I919446,I16897);
nand I_53927 (I919463,I919446,I919152);
nand I_53928 (I919480,I919398,I919463);
nand I_53929 (I918951,I919480,I919429);
nand I_53930 (I918948,I919463,I919347);
not I_53931 (I919552,I2690);
DFFARX1 I_53932 (I211667,I2683,I919552,I919578,);
and I_53933 (I919586,I919578,I211652);
DFFARX1 I_53934 (I919586,I2683,I919552,I919535,);
DFFARX1 I_53935 (I211658,I2683,I919552,I919626,);
not I_53936 (I919634,I211640);
not I_53937 (I919651,I211661);
nand I_53938 (I919668,I919651,I919634);
nor I_53939 (I919523,I919626,I919668);
DFFARX1 I_53940 (I919668,I2683,I919552,I919708,);
not I_53941 (I919544,I919708);
not I_53942 (I919730,I211664);
nand I_53943 (I919747,I919651,I919730);
DFFARX1 I_53944 (I919747,I2683,I919552,I919773,);
not I_53945 (I919781,I919773);
not I_53946 (I919798,I211655);
nand I_53947 (I919815,I919798,I211643);
and I_53948 (I919832,I919634,I919815);
nor I_53949 (I919849,I919747,I919832);
DFFARX1 I_53950 (I919849,I2683,I919552,I919520,);
DFFARX1 I_53951 (I919832,I2683,I919552,I919541,);
nor I_53952 (I919894,I211655,I211649);
nor I_53953 (I919532,I919747,I919894);
or I_53954 (I919925,I211655,I211649);
nor I_53955 (I919942,I211646,I211640);
DFFARX1 I_53956 (I919942,I2683,I919552,I919968,);
not I_53957 (I919976,I919968);
nor I_53958 (I919538,I919976,I919781);
nand I_53959 (I920007,I919976,I919626);
not I_53960 (I920024,I211646);
nand I_53961 (I920041,I920024,I919730);
nand I_53962 (I920058,I919976,I920041);
nand I_53963 (I919529,I920058,I920007);
nand I_53964 (I919526,I920041,I919925);
not I_53965 (I920130,I2690);
DFFARX1 I_53966 (I1009984,I2683,I920130,I920156,);
and I_53967 (I920164,I920156,I1009966);
DFFARX1 I_53968 (I920164,I2683,I920130,I920113,);
DFFARX1 I_53969 (I1009975,I2683,I920130,I920204,);
not I_53970 (I920212,I1009960);
not I_53971 (I920229,I1009972);
nand I_53972 (I920246,I920229,I920212);
nor I_53973 (I920101,I920204,I920246);
DFFARX1 I_53974 (I920246,I2683,I920130,I920286,);
not I_53975 (I920122,I920286);
not I_53976 (I920308,I1009963);
nand I_53977 (I920325,I920229,I920308);
DFFARX1 I_53978 (I920325,I2683,I920130,I920351,);
not I_53979 (I920359,I920351);
not I_53980 (I920376,I1009960);
nand I_53981 (I920393,I920376,I1009963);
and I_53982 (I920410,I920212,I920393);
nor I_53983 (I920427,I920325,I920410);
DFFARX1 I_53984 (I920427,I2683,I920130,I920098,);
DFFARX1 I_53985 (I920410,I2683,I920130,I920119,);
nor I_53986 (I920472,I1009960,I1009981);
nor I_53987 (I920110,I920325,I920472);
or I_53988 (I920503,I1009960,I1009981);
nor I_53989 (I920520,I1009969,I1009978);
DFFARX1 I_53990 (I920520,I2683,I920130,I920546,);
not I_53991 (I920554,I920546);
nor I_53992 (I920116,I920554,I920359);
nand I_53993 (I920585,I920554,I920204);
not I_53994 (I920602,I1009969);
nand I_53995 (I920619,I920602,I920308);
nand I_53996 (I920636,I920554,I920619);
nand I_53997 (I920107,I920636,I920585);
nand I_53998 (I920104,I920619,I920503);
not I_53999 (I920708,I2690);
DFFARX1 I_54000 (I580963,I2683,I920708,I920734,);
and I_54001 (I920742,I920734,I580951);
DFFARX1 I_54002 (I920742,I2683,I920708,I920691,);
DFFARX1 I_54003 (I580954,I2683,I920708,I920782,);
not I_54004 (I920790,I580948);
not I_54005 (I920807,I580972);
nand I_54006 (I920824,I920807,I920790);
nor I_54007 (I920679,I920782,I920824);
DFFARX1 I_54008 (I920824,I2683,I920708,I920864,);
not I_54009 (I920700,I920864);
not I_54010 (I920886,I580960);
nand I_54011 (I920903,I920807,I920886);
DFFARX1 I_54012 (I920903,I2683,I920708,I920929,);
not I_54013 (I920937,I920929);
not I_54014 (I920954,I580969);
nand I_54015 (I920971,I920954,I580966);
and I_54016 (I920988,I920790,I920971);
nor I_54017 (I921005,I920903,I920988);
DFFARX1 I_54018 (I921005,I2683,I920708,I920676,);
DFFARX1 I_54019 (I920988,I2683,I920708,I920697,);
nor I_54020 (I921050,I580969,I580957);
nor I_54021 (I920688,I920903,I921050);
or I_54022 (I921081,I580969,I580957);
nor I_54023 (I921098,I580948,I580951);
DFFARX1 I_54024 (I921098,I2683,I920708,I921124,);
not I_54025 (I921132,I921124);
nor I_54026 (I920694,I921132,I920937);
nand I_54027 (I921163,I921132,I920782);
not I_54028 (I921180,I580948);
nand I_54029 (I921197,I921180,I920886);
nand I_54030 (I921214,I921132,I921197);
nand I_54031 (I920685,I921214,I921163);
nand I_54032 (I920682,I921197,I921081);
not I_54033 (I921286,I2690);
DFFARX1 I_54034 (I230639,I2683,I921286,I921312,);
and I_54035 (I921320,I921312,I230624);
DFFARX1 I_54036 (I921320,I2683,I921286,I921269,);
DFFARX1 I_54037 (I230630,I2683,I921286,I921360,);
not I_54038 (I921368,I230612);
not I_54039 (I921385,I230633);
nand I_54040 (I921402,I921385,I921368);
nor I_54041 (I921257,I921360,I921402);
DFFARX1 I_54042 (I921402,I2683,I921286,I921442,);
not I_54043 (I921278,I921442);
not I_54044 (I921464,I230636);
nand I_54045 (I921481,I921385,I921464);
DFFARX1 I_54046 (I921481,I2683,I921286,I921507,);
not I_54047 (I921515,I921507);
not I_54048 (I921532,I230627);
nand I_54049 (I921549,I921532,I230615);
and I_54050 (I921566,I921368,I921549);
nor I_54051 (I921583,I921481,I921566);
DFFARX1 I_54052 (I921583,I2683,I921286,I921254,);
DFFARX1 I_54053 (I921566,I2683,I921286,I921275,);
nor I_54054 (I921628,I230627,I230621);
nor I_54055 (I921266,I921481,I921628);
or I_54056 (I921659,I230627,I230621);
nor I_54057 (I921676,I230618,I230612);
DFFARX1 I_54058 (I921676,I2683,I921286,I921702,);
not I_54059 (I921710,I921702);
nor I_54060 (I921272,I921710,I921515);
nand I_54061 (I921741,I921710,I921360);
not I_54062 (I921758,I230618);
nand I_54063 (I921775,I921758,I921464);
nand I_54064 (I921792,I921710,I921775);
nand I_54065 (I921263,I921792,I921741);
nand I_54066 (I921260,I921775,I921659);
not I_54067 (I921864,I2690);
DFFARX1 I_54068 (I558421,I2683,I921864,I921890,);
and I_54069 (I921898,I921890,I558409);
DFFARX1 I_54070 (I921898,I2683,I921864,I921847,);
DFFARX1 I_54071 (I558412,I2683,I921864,I921938,);
not I_54072 (I921946,I558406);
not I_54073 (I921963,I558430);
nand I_54074 (I921980,I921963,I921946);
nor I_54075 (I921835,I921938,I921980);
DFFARX1 I_54076 (I921980,I2683,I921864,I922020,);
not I_54077 (I921856,I922020);
not I_54078 (I922042,I558418);
nand I_54079 (I922059,I921963,I922042);
DFFARX1 I_54080 (I922059,I2683,I921864,I922085,);
not I_54081 (I922093,I922085);
not I_54082 (I922110,I558427);
nand I_54083 (I922127,I922110,I558424);
and I_54084 (I922144,I921946,I922127);
nor I_54085 (I922161,I922059,I922144);
DFFARX1 I_54086 (I922161,I2683,I921864,I921832,);
DFFARX1 I_54087 (I922144,I2683,I921864,I921853,);
nor I_54088 (I922206,I558427,I558415);
nor I_54089 (I921844,I922059,I922206);
or I_54090 (I922237,I558427,I558415);
nor I_54091 (I922254,I558406,I558409);
DFFARX1 I_54092 (I922254,I2683,I921864,I922280,);
not I_54093 (I922288,I922280);
nor I_54094 (I921850,I922288,I922093);
nand I_54095 (I922319,I922288,I921938);
not I_54096 (I922336,I558406);
nand I_54097 (I922353,I922336,I922042);
nand I_54098 (I922370,I922288,I922353);
nand I_54099 (I921841,I922370,I922319);
nand I_54100 (I921838,I922353,I922237);
not I_54101 (I922442,I2690);
DFFARX1 I_54102 (I305473,I2683,I922442,I922468,);
and I_54103 (I922476,I922468,I305458);
DFFARX1 I_54104 (I922476,I2683,I922442,I922425,);
DFFARX1 I_54105 (I305464,I2683,I922442,I922516,);
not I_54106 (I922524,I305446);
not I_54107 (I922541,I305467);
nand I_54108 (I922558,I922541,I922524);
nor I_54109 (I922413,I922516,I922558);
DFFARX1 I_54110 (I922558,I2683,I922442,I922598,);
not I_54111 (I922434,I922598);
not I_54112 (I922620,I305470);
nand I_54113 (I922637,I922541,I922620);
DFFARX1 I_54114 (I922637,I2683,I922442,I922663,);
not I_54115 (I922671,I922663);
not I_54116 (I922688,I305461);
nand I_54117 (I922705,I922688,I305449);
and I_54118 (I922722,I922524,I922705);
nor I_54119 (I922739,I922637,I922722);
DFFARX1 I_54120 (I922739,I2683,I922442,I922410,);
DFFARX1 I_54121 (I922722,I2683,I922442,I922431,);
nor I_54122 (I922784,I305461,I305455);
nor I_54123 (I922422,I922637,I922784);
or I_54124 (I922815,I305461,I305455);
nor I_54125 (I922832,I305452,I305446);
DFFARX1 I_54126 (I922832,I2683,I922442,I922858,);
not I_54127 (I922866,I922858);
nor I_54128 (I922428,I922866,I922671);
nand I_54129 (I922897,I922866,I922516);
not I_54130 (I922914,I305452);
nand I_54131 (I922931,I922914,I922620);
nand I_54132 (I922948,I922866,I922931);
nand I_54133 (I922419,I922948,I922897);
nand I_54134 (I922416,I922931,I922815);
not I_54135 (I923020,I2690);
DFFARX1 I_54136 (I572871,I2683,I923020,I923046,);
and I_54137 (I923054,I923046,I572859);
DFFARX1 I_54138 (I923054,I2683,I923020,I923003,);
DFFARX1 I_54139 (I572862,I2683,I923020,I923094,);
not I_54140 (I923102,I572856);
not I_54141 (I923119,I572880);
nand I_54142 (I923136,I923119,I923102);
nor I_54143 (I922991,I923094,I923136);
DFFARX1 I_54144 (I923136,I2683,I923020,I923176,);
not I_54145 (I923012,I923176);
not I_54146 (I923198,I572868);
nand I_54147 (I923215,I923119,I923198);
DFFARX1 I_54148 (I923215,I2683,I923020,I923241,);
not I_54149 (I923249,I923241);
not I_54150 (I923266,I572877);
nand I_54151 (I923283,I923266,I572874);
and I_54152 (I923300,I923102,I923283);
nor I_54153 (I923317,I923215,I923300);
DFFARX1 I_54154 (I923317,I2683,I923020,I922988,);
DFFARX1 I_54155 (I923300,I2683,I923020,I923009,);
nor I_54156 (I923362,I572877,I572865);
nor I_54157 (I923000,I923215,I923362);
or I_54158 (I923393,I572877,I572865);
nor I_54159 (I923410,I572856,I572859);
DFFARX1 I_54160 (I923410,I2683,I923020,I923436,);
not I_54161 (I923444,I923436);
nor I_54162 (I923006,I923444,I923249);
nand I_54163 (I923475,I923444,I923094);
not I_54164 (I923492,I572856);
nand I_54165 (I923509,I923492,I923198);
nand I_54166 (I923526,I923444,I923509);
nand I_54167 (I922997,I923526,I923475);
nand I_54168 (I922994,I923509,I923393);
not I_54169 (I923598,I2690);
DFFARX1 I_54170 (I1100716,I2683,I923598,I923624,);
and I_54171 (I923632,I923624,I1100698);
DFFARX1 I_54172 (I923632,I2683,I923598,I923581,);
DFFARX1 I_54173 (I1100689,I2683,I923598,I923672,);
not I_54174 (I923680,I1100704);
not I_54175 (I923697,I1100692);
nand I_54176 (I923714,I923697,I923680);
nor I_54177 (I923569,I923672,I923714);
DFFARX1 I_54178 (I923714,I2683,I923598,I923754,);
not I_54179 (I923590,I923754);
not I_54180 (I923776,I1100701);
nand I_54181 (I923793,I923697,I923776);
DFFARX1 I_54182 (I923793,I2683,I923598,I923819,);
not I_54183 (I923827,I923819);
not I_54184 (I923844,I1100710);
nand I_54185 (I923861,I923844,I1100689);
and I_54186 (I923878,I923680,I923861);
nor I_54187 (I923895,I923793,I923878);
DFFARX1 I_54188 (I923895,I2683,I923598,I923566,);
DFFARX1 I_54189 (I923878,I2683,I923598,I923587,);
nor I_54190 (I923940,I1100710,I1100713);
nor I_54191 (I923578,I923793,I923940);
or I_54192 (I923971,I1100710,I1100713);
nor I_54193 (I923988,I1100707,I1100695);
DFFARX1 I_54194 (I923988,I2683,I923598,I924014,);
not I_54195 (I924022,I924014);
nor I_54196 (I923584,I924022,I923827);
nand I_54197 (I924053,I924022,I923672);
not I_54198 (I924070,I1100707);
nand I_54199 (I924087,I924070,I923776);
nand I_54200 (I924104,I924022,I924087);
nand I_54201 (I923575,I924104,I924053);
nand I_54202 (I923572,I924087,I923971);
not I_54203 (I924176,I2690);
DFFARX1 I_54204 (I771677,I2683,I924176,I924202,);
and I_54205 (I924210,I924202,I771671);
DFFARX1 I_54206 (I924210,I2683,I924176,I924159,);
DFFARX1 I_54207 (I771689,I2683,I924176,I924250,);
not I_54208 (I924258,I771680);
not I_54209 (I924275,I771692);
nand I_54210 (I924292,I924275,I924258);
nor I_54211 (I924147,I924250,I924292);
DFFARX1 I_54212 (I924292,I2683,I924176,I924332,);
not I_54213 (I924168,I924332);
not I_54214 (I924354,I771698);
nand I_54215 (I924371,I924275,I924354);
DFFARX1 I_54216 (I924371,I2683,I924176,I924397,);
not I_54217 (I924405,I924397);
not I_54218 (I924422,I771674);
nand I_54219 (I924439,I924422,I771695);
and I_54220 (I924456,I924258,I924439);
nor I_54221 (I924473,I924371,I924456);
DFFARX1 I_54222 (I924473,I2683,I924176,I924144,);
DFFARX1 I_54223 (I924456,I2683,I924176,I924165,);
nor I_54224 (I924518,I771674,I771686);
nor I_54225 (I924156,I924371,I924518);
or I_54226 (I924549,I771674,I771686);
nor I_54227 (I924566,I771671,I771683);
DFFARX1 I_54228 (I924566,I2683,I924176,I924592,);
not I_54229 (I924600,I924592);
nor I_54230 (I924162,I924600,I924405);
nand I_54231 (I924631,I924600,I924250);
not I_54232 (I924648,I771671);
nand I_54233 (I924665,I924648,I924354);
nand I_54234 (I924682,I924600,I924665);
nand I_54235 (I924153,I924682,I924631);
nand I_54236 (I924150,I924665,I924549);
not I_54237 (I924754,I2690);
DFFARX1 I_54238 (I1008250,I2683,I924754,I924780,);
and I_54239 (I924788,I924780,I1008232);
DFFARX1 I_54240 (I924788,I2683,I924754,I924737,);
DFFARX1 I_54241 (I1008241,I2683,I924754,I924828,);
not I_54242 (I924836,I1008226);
not I_54243 (I924853,I1008238);
nand I_54244 (I924870,I924853,I924836);
nor I_54245 (I924725,I924828,I924870);
DFFARX1 I_54246 (I924870,I2683,I924754,I924910,);
not I_54247 (I924746,I924910);
not I_54248 (I924932,I1008229);
nand I_54249 (I924949,I924853,I924932);
DFFARX1 I_54250 (I924949,I2683,I924754,I924975,);
not I_54251 (I924983,I924975);
not I_54252 (I925000,I1008226);
nand I_54253 (I925017,I925000,I1008229);
and I_54254 (I925034,I924836,I925017);
nor I_54255 (I925051,I924949,I925034);
DFFARX1 I_54256 (I925051,I2683,I924754,I924722,);
DFFARX1 I_54257 (I925034,I2683,I924754,I924743,);
nor I_54258 (I925096,I1008226,I1008247);
nor I_54259 (I924734,I924949,I925096);
or I_54260 (I925127,I1008226,I1008247);
nor I_54261 (I925144,I1008235,I1008244);
DFFARX1 I_54262 (I925144,I2683,I924754,I925170,);
not I_54263 (I925178,I925170);
nor I_54264 (I924740,I925178,I924983);
nand I_54265 (I925209,I925178,I924828);
not I_54266 (I925226,I1008235);
nand I_54267 (I925243,I925226,I924932);
nand I_54268 (I925260,I925178,I925243);
nand I_54269 (I924731,I925260,I925209);
nand I_54270 (I924728,I925243,I925127);
not I_54271 (I925332,I2690);
DFFARX1 I_54272 (I417530,I2683,I925332,I925358,);
and I_54273 (I925366,I925358,I417545);
DFFARX1 I_54274 (I925366,I2683,I925332,I925315,);
DFFARX1 I_54275 (I417536,I2683,I925332,I925406,);
not I_54276 (I925414,I417530);
not I_54277 (I925431,I417548);
nand I_54278 (I925448,I925431,I925414);
nor I_54279 (I925303,I925406,I925448);
DFFARX1 I_54280 (I925448,I2683,I925332,I925488,);
not I_54281 (I925324,I925488);
not I_54282 (I925510,I417539);
nand I_54283 (I925527,I925431,I925510);
DFFARX1 I_54284 (I925527,I2683,I925332,I925553,);
not I_54285 (I925561,I925553);
not I_54286 (I925578,I417551);
nand I_54287 (I925595,I925578,I417527);
and I_54288 (I925612,I925414,I925595);
nor I_54289 (I925629,I925527,I925612);
DFFARX1 I_54290 (I925629,I2683,I925332,I925300,);
DFFARX1 I_54291 (I925612,I2683,I925332,I925321,);
nor I_54292 (I925674,I417551,I417527);
nor I_54293 (I925312,I925527,I925674);
or I_54294 (I925705,I417551,I417527);
nor I_54295 (I925722,I417533,I417542);
DFFARX1 I_54296 (I925722,I2683,I925332,I925748,);
not I_54297 (I925756,I925748);
nor I_54298 (I925318,I925756,I925561);
nand I_54299 (I925787,I925756,I925406);
not I_54300 (I925804,I417533);
nand I_54301 (I925821,I925804,I925510);
nand I_54302 (I925838,I925756,I925821);
nand I_54303 (I925309,I925838,I925787);
nand I_54304 (I925306,I925821,I925705);
not I_54305 (I925910,I2690);
DFFARX1 I_54306 (I542815,I2683,I925910,I925936,);
and I_54307 (I925944,I925936,I542803);
DFFARX1 I_54308 (I925944,I2683,I925910,I925893,);
DFFARX1 I_54309 (I542806,I2683,I925910,I925984,);
not I_54310 (I925992,I542800);
not I_54311 (I926009,I542824);
nand I_54312 (I926026,I926009,I925992);
nor I_54313 (I925881,I925984,I926026);
DFFARX1 I_54314 (I926026,I2683,I925910,I926066,);
not I_54315 (I925902,I926066);
not I_54316 (I926088,I542812);
nand I_54317 (I926105,I926009,I926088);
DFFARX1 I_54318 (I926105,I2683,I925910,I926131,);
not I_54319 (I926139,I926131);
not I_54320 (I926156,I542821);
nand I_54321 (I926173,I926156,I542818);
and I_54322 (I926190,I925992,I926173);
nor I_54323 (I926207,I926105,I926190);
DFFARX1 I_54324 (I926207,I2683,I925910,I925878,);
DFFARX1 I_54325 (I926190,I2683,I925910,I925899,);
nor I_54326 (I926252,I542821,I542809);
nor I_54327 (I925890,I926105,I926252);
or I_54328 (I926283,I542821,I542809);
nor I_54329 (I926300,I542800,I542803);
DFFARX1 I_54330 (I926300,I2683,I925910,I926326,);
not I_54331 (I926334,I926326);
nor I_54332 (I925896,I926334,I926139);
nand I_54333 (I926365,I926334,I925984);
not I_54334 (I926382,I542800);
nand I_54335 (I926399,I926382,I926088);
nand I_54336 (I926416,I926334,I926399);
nand I_54337 (I925887,I926416,I926365);
nand I_54338 (I925884,I926399,I926283);
not I_54339 (I926488,I2690);
DFFARX1 I_54340 (I331218,I2683,I926488,I926514,);
and I_54341 (I926522,I926514,I331233);
DFFARX1 I_54342 (I926522,I2683,I926488,I926471,);
DFFARX1 I_54343 (I331236,I2683,I926488,I926562,);
not I_54344 (I926570,I331230);
not I_54345 (I926587,I331245);
nand I_54346 (I926604,I926587,I926570);
nor I_54347 (I926459,I926562,I926604);
DFFARX1 I_54348 (I926604,I2683,I926488,I926644,);
not I_54349 (I926480,I926644);
not I_54350 (I926666,I331221);
nand I_54351 (I926683,I926587,I926666);
DFFARX1 I_54352 (I926683,I2683,I926488,I926709,);
not I_54353 (I926717,I926709);
not I_54354 (I926734,I331224);
nand I_54355 (I926751,I926734,I331218);
and I_54356 (I926768,I926570,I926751);
nor I_54357 (I926785,I926683,I926768);
DFFARX1 I_54358 (I926785,I2683,I926488,I926456,);
DFFARX1 I_54359 (I926768,I2683,I926488,I926477,);
nor I_54360 (I926830,I331224,I331227);
nor I_54361 (I926468,I926683,I926830);
or I_54362 (I926861,I331224,I331227);
nor I_54363 (I926878,I331242,I331239);
DFFARX1 I_54364 (I926878,I2683,I926488,I926904,);
not I_54365 (I926912,I926904);
nor I_54366 (I926474,I926912,I926717);
nand I_54367 (I926943,I926912,I926562);
not I_54368 (I926960,I331242);
nand I_54369 (I926977,I926960,I926666);
nand I_54370 (I926994,I926912,I926977);
nand I_54371 (I926465,I926994,I926943);
nand I_54372 (I926462,I926977,I926861);
not I_54373 (I927066,I2690);
DFFARX1 I_54374 (I727749,I2683,I927066,I927092,);
and I_54375 (I927100,I927092,I727743);
DFFARX1 I_54376 (I927100,I2683,I927066,I927049,);
DFFARX1 I_54377 (I727761,I2683,I927066,I927140,);
not I_54378 (I927148,I727752);
not I_54379 (I927165,I727764);
nand I_54380 (I927182,I927165,I927148);
nor I_54381 (I927037,I927140,I927182);
DFFARX1 I_54382 (I927182,I2683,I927066,I927222,);
not I_54383 (I927058,I927222);
not I_54384 (I927244,I727770);
nand I_54385 (I927261,I927165,I927244);
DFFARX1 I_54386 (I927261,I2683,I927066,I927287,);
not I_54387 (I927295,I927287);
not I_54388 (I927312,I727746);
nand I_54389 (I927329,I927312,I727767);
and I_54390 (I927346,I927148,I927329);
nor I_54391 (I927363,I927261,I927346);
DFFARX1 I_54392 (I927363,I2683,I927066,I927034,);
DFFARX1 I_54393 (I927346,I2683,I927066,I927055,);
nor I_54394 (I927408,I727746,I727758);
nor I_54395 (I927046,I927261,I927408);
or I_54396 (I927439,I727746,I727758);
nor I_54397 (I927456,I727743,I727755);
DFFARX1 I_54398 (I927456,I2683,I927066,I927482,);
not I_54399 (I927490,I927482);
nor I_54400 (I927052,I927490,I927295);
nand I_54401 (I927521,I927490,I927140);
not I_54402 (I927538,I727743);
nand I_54403 (I927555,I927538,I927244);
nand I_54404 (I927572,I927490,I927555);
nand I_54405 (I927043,I927572,I927521);
nand I_54406 (I927040,I927555,I927439);
not I_54407 (I927644,I2690);
DFFARX1 I_54408 (I510447,I2683,I927644,I927670,);
and I_54409 (I927678,I927670,I510435);
DFFARX1 I_54410 (I927678,I2683,I927644,I927627,);
DFFARX1 I_54411 (I510438,I2683,I927644,I927718,);
not I_54412 (I927726,I510432);
not I_54413 (I927743,I510456);
nand I_54414 (I927760,I927743,I927726);
nor I_54415 (I927615,I927718,I927760);
DFFARX1 I_54416 (I927760,I2683,I927644,I927800,);
not I_54417 (I927636,I927800);
not I_54418 (I927822,I510444);
nand I_54419 (I927839,I927743,I927822);
DFFARX1 I_54420 (I927839,I2683,I927644,I927865,);
not I_54421 (I927873,I927865);
not I_54422 (I927890,I510453);
nand I_54423 (I927907,I927890,I510450);
and I_54424 (I927924,I927726,I927907);
nor I_54425 (I927941,I927839,I927924);
DFFARX1 I_54426 (I927941,I2683,I927644,I927612,);
DFFARX1 I_54427 (I927924,I2683,I927644,I927633,);
nor I_54428 (I927986,I510453,I510441);
nor I_54429 (I927624,I927839,I927986);
or I_54430 (I928017,I510453,I510441);
nor I_54431 (I928034,I510432,I510435);
DFFARX1 I_54432 (I928034,I2683,I927644,I928060,);
not I_54433 (I928068,I928060);
nor I_54434 (I927630,I928068,I927873);
nand I_54435 (I928099,I928068,I927718);
not I_54436 (I928116,I510432);
nand I_54437 (I928133,I928116,I927822);
nand I_54438 (I928150,I928068,I928133);
nand I_54439 (I927621,I928150,I928099);
nand I_54440 (I927618,I928133,I928017);
not I_54441 (I928222,I2690);
DFFARX1 I_54442 (I648084,I2683,I928222,I928248,);
and I_54443 (I928256,I928248,I648090);
DFFARX1 I_54444 (I928256,I2683,I928222,I928205,);
DFFARX1 I_54445 (I648096,I2683,I928222,I928296,);
not I_54446 (I928304,I648081);
not I_54447 (I928321,I648081);
nand I_54448 (I928338,I928321,I928304);
nor I_54449 (I928193,I928296,I928338);
DFFARX1 I_54450 (I928338,I2683,I928222,I928378,);
not I_54451 (I928214,I928378);
not I_54452 (I928400,I648099);
nand I_54453 (I928417,I928321,I928400);
DFFARX1 I_54454 (I928417,I2683,I928222,I928443,);
not I_54455 (I928451,I928443);
not I_54456 (I928468,I648093);
nand I_54457 (I928485,I928468,I648084);
and I_54458 (I928502,I928304,I928485);
nor I_54459 (I928519,I928417,I928502);
DFFARX1 I_54460 (I928519,I2683,I928222,I928190,);
DFFARX1 I_54461 (I928502,I2683,I928222,I928211,);
nor I_54462 (I928564,I648093,I648102);
nor I_54463 (I928202,I928417,I928564);
or I_54464 (I928595,I648093,I648102);
nor I_54465 (I928612,I648087,I648087);
DFFARX1 I_54466 (I928612,I2683,I928222,I928638,);
not I_54467 (I928646,I928638);
nor I_54468 (I928208,I928646,I928451);
nand I_54469 (I928677,I928646,I928296);
not I_54470 (I928694,I648087);
nand I_54471 (I928711,I928694,I928400);
nand I_54472 (I928728,I928646,I928711);
nand I_54473 (I928199,I928728,I928677);
nand I_54474 (I928196,I928711,I928595);
not I_54475 (I928800,I2690);
DFFARX1 I_54476 (I765863,I2683,I928800,I928826,);
and I_54477 (I928834,I928826,I765857);
DFFARX1 I_54478 (I928834,I2683,I928800,I928783,);
DFFARX1 I_54479 (I765875,I2683,I928800,I928874,);
not I_54480 (I928882,I765866);
not I_54481 (I928899,I765878);
nand I_54482 (I928916,I928899,I928882);
nor I_54483 (I928771,I928874,I928916);
DFFARX1 I_54484 (I928916,I2683,I928800,I928956,);
not I_54485 (I928792,I928956);
not I_54486 (I928978,I765884);
nand I_54487 (I928995,I928899,I928978);
DFFARX1 I_54488 (I928995,I2683,I928800,I929021,);
not I_54489 (I929029,I929021);
not I_54490 (I929046,I765860);
nand I_54491 (I929063,I929046,I765881);
and I_54492 (I929080,I928882,I929063);
nor I_54493 (I929097,I928995,I929080);
DFFARX1 I_54494 (I929097,I2683,I928800,I928768,);
DFFARX1 I_54495 (I929080,I2683,I928800,I928789,);
nor I_54496 (I929142,I765860,I765872);
nor I_54497 (I928780,I928995,I929142);
or I_54498 (I929173,I765860,I765872);
nor I_54499 (I929190,I765857,I765869);
DFFARX1 I_54500 (I929190,I2683,I928800,I929216,);
not I_54501 (I929224,I929216);
nor I_54502 (I928786,I929224,I929029);
nand I_54503 (I929255,I929224,I928874);
not I_54504 (I929272,I765857);
nand I_54505 (I929289,I929272,I928978);
nand I_54506 (I929306,I929224,I929289);
nand I_54507 (I928777,I929306,I929255);
nand I_54508 (I928774,I929289,I929173);
not I_54509 (I929378,I2690);
DFFARX1 I_54510 (I45346,I2683,I929378,I929404,);
and I_54511 (I929412,I929404,I45349);
DFFARX1 I_54512 (I929412,I2683,I929378,I929361,);
DFFARX1 I_54513 (I45349,I2683,I929378,I929452,);
not I_54514 (I929460,I45352);
not I_54515 (I929477,I45367);
nand I_54516 (I929494,I929477,I929460);
nor I_54517 (I929349,I929452,I929494);
DFFARX1 I_54518 (I929494,I2683,I929378,I929534,);
not I_54519 (I929370,I929534);
not I_54520 (I929556,I45361);
nand I_54521 (I929573,I929477,I929556);
DFFARX1 I_54522 (I929573,I2683,I929378,I929599,);
not I_54523 (I929607,I929599);
not I_54524 (I929624,I45364);
nand I_54525 (I929641,I929624,I45346);
and I_54526 (I929658,I929460,I929641);
nor I_54527 (I929675,I929573,I929658);
DFFARX1 I_54528 (I929675,I2683,I929378,I929346,);
DFFARX1 I_54529 (I929658,I2683,I929378,I929367,);
nor I_54530 (I929720,I45364,I45358);
nor I_54531 (I929358,I929573,I929720);
or I_54532 (I929751,I45364,I45358);
nor I_54533 (I929768,I45355,I45370);
DFFARX1 I_54534 (I929768,I2683,I929378,I929794,);
not I_54535 (I929802,I929794);
nor I_54536 (I929364,I929802,I929607);
nand I_54537 (I929833,I929802,I929452);
not I_54538 (I929850,I45355);
nand I_54539 (I929867,I929850,I929556);
nand I_54540 (I929884,I929802,I929867);
nand I_54541 (I929355,I929884,I929833);
nand I_54542 (I929352,I929867,I929751);
not I_54543 (I929956,I2690);
DFFARX1 I_54544 (I272799,I2683,I929956,I929982,);
and I_54545 (I929990,I929982,I272784);
DFFARX1 I_54546 (I929990,I2683,I929956,I929939,);
DFFARX1 I_54547 (I272790,I2683,I929956,I930030,);
not I_54548 (I930038,I272772);
not I_54549 (I930055,I272793);
nand I_54550 (I930072,I930055,I930038);
nor I_54551 (I929927,I930030,I930072);
DFFARX1 I_54552 (I930072,I2683,I929956,I930112,);
not I_54553 (I929948,I930112);
not I_54554 (I930134,I272796);
nand I_54555 (I930151,I930055,I930134);
DFFARX1 I_54556 (I930151,I2683,I929956,I930177,);
not I_54557 (I930185,I930177);
not I_54558 (I930202,I272787);
nand I_54559 (I930219,I930202,I272775);
and I_54560 (I930236,I930038,I930219);
nor I_54561 (I930253,I930151,I930236);
DFFARX1 I_54562 (I930253,I2683,I929956,I929924,);
DFFARX1 I_54563 (I930236,I2683,I929956,I929945,);
nor I_54564 (I930298,I272787,I272781);
nor I_54565 (I929936,I930151,I930298);
or I_54566 (I930329,I272787,I272781);
nor I_54567 (I930346,I272778,I272772);
DFFARX1 I_54568 (I930346,I2683,I929956,I930372,);
not I_54569 (I930380,I930372);
nor I_54570 (I929942,I930380,I930185);
nand I_54571 (I930411,I930380,I930030);
not I_54572 (I930428,I272778);
nand I_54573 (I930445,I930428,I930134);
nand I_54574 (I930462,I930380,I930445);
nand I_54575 (I929933,I930462,I930411);
nand I_54576 (I929930,I930445,I930329);
not I_54577 (I930534,I2690);
DFFARX1 I_54578 (I501777,I2683,I930534,I930560,);
and I_54579 (I930568,I930560,I501765);
DFFARX1 I_54580 (I930568,I2683,I930534,I930517,);
DFFARX1 I_54581 (I501768,I2683,I930534,I930608,);
not I_54582 (I930616,I501762);
not I_54583 (I930633,I501786);
nand I_54584 (I930650,I930633,I930616);
nor I_54585 (I930505,I930608,I930650);
DFFARX1 I_54586 (I930650,I2683,I930534,I930690,);
not I_54587 (I930526,I930690);
not I_54588 (I930712,I501774);
nand I_54589 (I930729,I930633,I930712);
DFFARX1 I_54590 (I930729,I2683,I930534,I930755,);
not I_54591 (I930763,I930755);
not I_54592 (I930780,I501783);
nand I_54593 (I930797,I930780,I501780);
and I_54594 (I930814,I930616,I930797);
nor I_54595 (I930831,I930729,I930814);
DFFARX1 I_54596 (I930831,I2683,I930534,I930502,);
DFFARX1 I_54597 (I930814,I2683,I930534,I930523,);
nor I_54598 (I930876,I501783,I501771);
nor I_54599 (I930514,I930729,I930876);
or I_54600 (I930907,I501783,I501771);
nor I_54601 (I930924,I501762,I501765);
DFFARX1 I_54602 (I930924,I2683,I930534,I930950,);
not I_54603 (I930958,I930950);
nor I_54604 (I930520,I930958,I930763);
nand I_54605 (I930989,I930958,I930608);
not I_54606 (I931006,I501762);
nand I_54607 (I931023,I931006,I930712);
nand I_54608 (I931040,I930958,I931023);
nand I_54609 (I930511,I931040,I930989);
nand I_54610 (I930508,I931023,I930907);
not I_54611 (I931112,I2690);
DFFARX1 I_54612 (I1007672,I2683,I931112,I931138,);
and I_54613 (I931146,I931138,I1007654);
DFFARX1 I_54614 (I931146,I2683,I931112,I931095,);
DFFARX1 I_54615 (I1007663,I2683,I931112,I931186,);
not I_54616 (I931194,I1007648);
not I_54617 (I931211,I1007660);
nand I_54618 (I931228,I931211,I931194);
nor I_54619 (I931083,I931186,I931228);
DFFARX1 I_54620 (I931228,I2683,I931112,I931268,);
not I_54621 (I931104,I931268);
not I_54622 (I931290,I1007651);
nand I_54623 (I931307,I931211,I931290);
DFFARX1 I_54624 (I931307,I2683,I931112,I931333,);
not I_54625 (I931341,I931333);
not I_54626 (I931358,I1007648);
nand I_54627 (I931375,I931358,I1007651);
and I_54628 (I931392,I931194,I931375);
nor I_54629 (I931409,I931307,I931392);
DFFARX1 I_54630 (I931409,I2683,I931112,I931080,);
DFFARX1 I_54631 (I931392,I2683,I931112,I931101,);
nor I_54632 (I931454,I1007648,I1007669);
nor I_54633 (I931092,I931307,I931454);
or I_54634 (I931485,I1007648,I1007669);
nor I_54635 (I931502,I1007657,I1007666);
DFFARX1 I_54636 (I931502,I2683,I931112,I931528,);
not I_54637 (I931536,I931528);
nor I_54638 (I931098,I931536,I931341);
nand I_54639 (I931567,I931536,I931186);
not I_54640 (I931584,I1007657);
nand I_54641 (I931601,I931584,I931290);
nand I_54642 (I931618,I931536,I931601);
nand I_54643 (I931089,I931618,I931567);
nand I_54644 (I931086,I931601,I931485);
not I_54645 (I931690,I2690);
DFFARX1 I_54646 (I390514,I2683,I931690,I931716,);
and I_54647 (I931724,I931716,I390529);
DFFARX1 I_54648 (I931724,I2683,I931690,I931673,);
DFFARX1 I_54649 (I390532,I2683,I931690,I931764,);
not I_54650 (I931772,I390526);
not I_54651 (I931789,I390541);
nand I_54652 (I931806,I931789,I931772);
nor I_54653 (I931661,I931764,I931806);
DFFARX1 I_54654 (I931806,I2683,I931690,I931846,);
not I_54655 (I931682,I931846);
not I_54656 (I931868,I390517);
nand I_54657 (I931885,I931789,I931868);
DFFARX1 I_54658 (I931885,I2683,I931690,I931911,);
not I_54659 (I931919,I931911);
not I_54660 (I931936,I390520);
nand I_54661 (I931953,I931936,I390514);
and I_54662 (I931970,I931772,I931953);
nor I_54663 (I931987,I931885,I931970);
DFFARX1 I_54664 (I931987,I2683,I931690,I931658,);
DFFARX1 I_54665 (I931970,I2683,I931690,I931679,);
nor I_54666 (I932032,I390520,I390523);
nor I_54667 (I931670,I931885,I932032);
or I_54668 (I932063,I390520,I390523);
nor I_54669 (I932080,I390538,I390535);
DFFARX1 I_54670 (I932080,I2683,I931690,I932106,);
not I_54671 (I932114,I932106);
nor I_54672 (I931676,I932114,I931919);
nand I_54673 (I932145,I932114,I931764);
not I_54674 (I932162,I390538);
nand I_54675 (I932179,I932162,I931868);
nand I_54676 (I932196,I932114,I932179);
nand I_54677 (I931667,I932196,I932145);
nand I_54678 (I931664,I932179,I932063);
not I_54679 (I932268,I2690);
DFFARX1 I_54680 (I158090,I2683,I932268,I932294,);
and I_54681 (I932302,I932294,I158093);
DFFARX1 I_54682 (I932302,I2683,I932268,I932251,);
DFFARX1 I_54683 (I158093,I2683,I932268,I932342,);
not I_54684 (I932350,I158108);
not I_54685 (I932367,I158114);
nand I_54686 (I932384,I932367,I932350);
nor I_54687 (I932239,I932342,I932384);
DFFARX1 I_54688 (I932384,I2683,I932268,I932424,);
not I_54689 (I932260,I932424);
not I_54690 (I932446,I158102);
nand I_54691 (I932463,I932367,I932446);
DFFARX1 I_54692 (I932463,I2683,I932268,I932489,);
not I_54693 (I932497,I932489);
not I_54694 (I932514,I158099);
nand I_54695 (I932531,I932514,I158096);
and I_54696 (I932548,I932350,I932531);
nor I_54697 (I932565,I932463,I932548);
DFFARX1 I_54698 (I932565,I2683,I932268,I932236,);
DFFARX1 I_54699 (I932548,I2683,I932268,I932257,);
nor I_54700 (I932610,I158099,I158090);
nor I_54701 (I932248,I932463,I932610);
or I_54702 (I932641,I158099,I158090);
nor I_54703 (I932658,I158105,I158111);
DFFARX1 I_54704 (I932658,I2683,I932268,I932684,);
not I_54705 (I932692,I932684);
nor I_54706 (I932254,I932692,I932497);
nand I_54707 (I932723,I932692,I932342);
not I_54708 (I932740,I158105);
nand I_54709 (I932757,I932740,I932446);
nand I_54710 (I932774,I932692,I932757);
nand I_54711 (I932245,I932774,I932723);
nand I_54712 (I932242,I932757,I932641);
not I_54713 (I932846,I2690);
DFFARX1 I_54714 (I83314,I2683,I932846,I932872,);
and I_54715 (I932880,I932872,I83290);
DFFARX1 I_54716 (I932880,I2683,I932846,I932829,);
DFFARX1 I_54717 (I83308,I2683,I932846,I932920,);
not I_54718 (I932928,I83296);
not I_54719 (I932945,I83293);
nand I_54720 (I932962,I932945,I932928);
nor I_54721 (I932817,I932920,I932962);
DFFARX1 I_54722 (I932962,I2683,I932846,I933002,);
not I_54723 (I932838,I933002);
not I_54724 (I933024,I83302);
nand I_54725 (I933041,I932945,I933024);
DFFARX1 I_54726 (I933041,I2683,I932846,I933067,);
not I_54727 (I933075,I933067);
not I_54728 (I933092,I83293);
nand I_54729 (I933109,I933092,I83311);
and I_54730 (I933126,I932928,I933109);
nor I_54731 (I933143,I933041,I933126);
DFFARX1 I_54732 (I933143,I2683,I932846,I932814,);
DFFARX1 I_54733 (I933126,I2683,I932846,I932835,);
nor I_54734 (I933188,I83293,I83305);
nor I_54735 (I932826,I933041,I933188);
or I_54736 (I933219,I83293,I83305);
nor I_54737 (I933236,I83299,I83290);
DFFARX1 I_54738 (I933236,I2683,I932846,I933262,);
not I_54739 (I933270,I933262);
nor I_54740 (I932832,I933270,I933075);
nand I_54741 (I933301,I933270,I932920);
not I_54742 (I933318,I83299);
nand I_54743 (I933335,I933318,I933024);
nand I_54744 (I933352,I933270,I933335);
nand I_54745 (I932823,I933352,I933301);
nand I_54746 (I932820,I933335,I933219);
not I_54747 (I933424,I2690);
DFFARX1 I_54748 (I341010,I2683,I933424,I933450,);
and I_54749 (I933458,I933450,I341025);
DFFARX1 I_54750 (I933458,I2683,I933424,I933407,);
DFFARX1 I_54751 (I341028,I2683,I933424,I933498,);
not I_54752 (I933506,I341022);
not I_54753 (I933523,I341037);
nand I_54754 (I933540,I933523,I933506);
nor I_54755 (I933395,I933498,I933540);
DFFARX1 I_54756 (I933540,I2683,I933424,I933580,);
not I_54757 (I933416,I933580);
not I_54758 (I933602,I341013);
nand I_54759 (I933619,I933523,I933602);
DFFARX1 I_54760 (I933619,I2683,I933424,I933645,);
not I_54761 (I933653,I933645);
not I_54762 (I933670,I341016);
nand I_54763 (I933687,I933670,I341010);
and I_54764 (I933704,I933506,I933687);
nor I_54765 (I933721,I933619,I933704);
DFFARX1 I_54766 (I933721,I2683,I933424,I933392,);
DFFARX1 I_54767 (I933704,I2683,I933424,I933413,);
nor I_54768 (I933766,I341016,I341019);
nor I_54769 (I933404,I933619,I933766);
or I_54770 (I933797,I341016,I341019);
nor I_54771 (I933814,I341034,I341031);
DFFARX1 I_54772 (I933814,I2683,I933424,I933840,);
not I_54773 (I933848,I933840);
nor I_54774 (I933410,I933848,I933653);
nand I_54775 (I933879,I933848,I933498);
not I_54776 (I933896,I341034);
nand I_54777 (I933913,I933896,I933602);
nand I_54778 (I933930,I933848,I933913);
nand I_54779 (I933401,I933930,I933879);
nand I_54780 (I933398,I933913,I933797);
not I_54781 (I934002,I2690);
DFFARX1 I_54782 (I103867,I2683,I934002,I934028,);
and I_54783 (I934036,I934028,I103843);
DFFARX1 I_54784 (I934036,I2683,I934002,I933985,);
DFFARX1 I_54785 (I103861,I2683,I934002,I934076,);
not I_54786 (I934084,I103849);
not I_54787 (I934101,I103846);
nand I_54788 (I934118,I934101,I934084);
nor I_54789 (I933973,I934076,I934118);
DFFARX1 I_54790 (I934118,I2683,I934002,I934158,);
not I_54791 (I933994,I934158);
not I_54792 (I934180,I103855);
nand I_54793 (I934197,I934101,I934180);
DFFARX1 I_54794 (I934197,I2683,I934002,I934223,);
not I_54795 (I934231,I934223);
not I_54796 (I934248,I103846);
nand I_54797 (I934265,I934248,I103864);
and I_54798 (I934282,I934084,I934265);
nor I_54799 (I934299,I934197,I934282);
DFFARX1 I_54800 (I934299,I2683,I934002,I933970,);
DFFARX1 I_54801 (I934282,I2683,I934002,I933991,);
nor I_54802 (I934344,I103846,I103858);
nor I_54803 (I933982,I934197,I934344);
or I_54804 (I934375,I103846,I103858);
nor I_54805 (I934392,I103852,I103843);
DFFARX1 I_54806 (I934392,I2683,I934002,I934418,);
not I_54807 (I934426,I934418);
nor I_54808 (I933988,I934426,I934231);
nand I_54809 (I934457,I934426,I934076);
not I_54810 (I934474,I103852);
nand I_54811 (I934491,I934474,I934180);
nand I_54812 (I934508,I934426,I934491);
nand I_54813 (I933979,I934508,I934457);
nand I_54814 (I933976,I934491,I934375);
not I_54815 (I934580,I2690);
DFFARX1 I_54816 (I1044786,I2683,I934580,I934606,);
and I_54817 (I934614,I934606,I1044768);
DFFARX1 I_54818 (I934614,I2683,I934580,I934563,);
DFFARX1 I_54819 (I1044759,I2683,I934580,I934654,);
not I_54820 (I934662,I1044774);
not I_54821 (I934679,I1044762);
nand I_54822 (I934696,I934679,I934662);
nor I_54823 (I934551,I934654,I934696);
DFFARX1 I_54824 (I934696,I2683,I934580,I934736,);
not I_54825 (I934572,I934736);
not I_54826 (I934758,I1044771);
nand I_54827 (I934775,I934679,I934758);
DFFARX1 I_54828 (I934775,I2683,I934580,I934801,);
not I_54829 (I934809,I934801);
not I_54830 (I934826,I1044780);
nand I_54831 (I934843,I934826,I1044759);
and I_54832 (I934860,I934662,I934843);
nor I_54833 (I934877,I934775,I934860);
DFFARX1 I_54834 (I934877,I2683,I934580,I934548,);
DFFARX1 I_54835 (I934860,I2683,I934580,I934569,);
nor I_54836 (I934922,I1044780,I1044783);
nor I_54837 (I934560,I934775,I934922);
or I_54838 (I934953,I1044780,I1044783);
nor I_54839 (I934970,I1044777,I1044765);
DFFARX1 I_54840 (I934970,I2683,I934580,I934996,);
not I_54841 (I935004,I934996);
nor I_54842 (I934566,I935004,I934809);
nand I_54843 (I935035,I935004,I934654);
not I_54844 (I935052,I1044777);
nand I_54845 (I935069,I935052,I934758);
nand I_54846 (I935086,I935004,I935069);
nand I_54847 (I934557,I935086,I935035);
nand I_54848 (I934554,I935069,I934953);
not I_54849 (I935158,I2690);
DFFARX1 I_54850 (I977715,I2683,I935158,I935184,);
and I_54851 (I935192,I935184,I977709);
DFFARX1 I_54852 (I935192,I2683,I935158,I935141,);
DFFARX1 I_54853 (I977694,I2683,I935158,I935232,);
not I_54854 (I935240,I977700);
not I_54855 (I935257,I977712);
nand I_54856 (I935274,I935257,I935240);
nor I_54857 (I935129,I935232,I935274);
DFFARX1 I_54858 (I935274,I2683,I935158,I935314,);
not I_54859 (I935150,I935314);
not I_54860 (I935336,I977694);
nand I_54861 (I935353,I935257,I935336);
DFFARX1 I_54862 (I935353,I2683,I935158,I935379,);
not I_54863 (I935387,I935379);
not I_54864 (I935404,I977718);
nand I_54865 (I935421,I935404,I977706);
and I_54866 (I935438,I935240,I935421);
nor I_54867 (I935455,I935353,I935438);
DFFARX1 I_54868 (I935455,I2683,I935158,I935126,);
DFFARX1 I_54869 (I935438,I2683,I935158,I935147,);
nor I_54870 (I935500,I977718,I977697);
nor I_54871 (I935138,I935353,I935500);
or I_54872 (I935531,I977718,I977697);
nor I_54873 (I935548,I977703,I977697);
DFFARX1 I_54874 (I935548,I2683,I935158,I935574,);
not I_54875 (I935582,I935574);
nor I_54876 (I935144,I935582,I935387);
nand I_54877 (I935613,I935582,I935232);
not I_54878 (I935630,I977703);
nand I_54879 (I935647,I935630,I935336);
nand I_54880 (I935664,I935582,I935647);
nand I_54881 (I935135,I935664,I935613);
nand I_54882 (I935132,I935647,I935531);
not I_54883 (I935736,I2690);
DFFARX1 I_54884 (I955955,I2683,I935736,I935762,);
and I_54885 (I935770,I935762,I955949);
DFFARX1 I_54886 (I935770,I2683,I935736,I935719,);
DFFARX1 I_54887 (I955934,I2683,I935736,I935810,);
not I_54888 (I935818,I955940);
not I_54889 (I935835,I955952);
nand I_54890 (I935852,I935835,I935818);
nor I_54891 (I935707,I935810,I935852);
DFFARX1 I_54892 (I935852,I2683,I935736,I935892,);
not I_54893 (I935728,I935892);
not I_54894 (I935914,I955934);
nand I_54895 (I935931,I935835,I935914);
DFFARX1 I_54896 (I935931,I2683,I935736,I935957,);
not I_54897 (I935965,I935957);
not I_54898 (I935982,I955958);
nand I_54899 (I935999,I935982,I955946);
and I_54900 (I936016,I935818,I935999);
nor I_54901 (I936033,I935931,I936016);
DFFARX1 I_54902 (I936033,I2683,I935736,I935704,);
DFFARX1 I_54903 (I936016,I2683,I935736,I935725,);
nor I_54904 (I936078,I955958,I955937);
nor I_54905 (I935716,I935931,I936078);
or I_54906 (I936109,I955958,I955937);
nor I_54907 (I936126,I955943,I955937);
DFFARX1 I_54908 (I936126,I2683,I935736,I936152,);
not I_54909 (I936160,I936152);
nor I_54910 (I935722,I936160,I935965);
nand I_54911 (I936191,I936160,I935810);
not I_54912 (I936208,I955943);
nand I_54913 (I936225,I936208,I935914);
nand I_54914 (I936242,I936160,I936225);
nand I_54915 (I935713,I936242,I936191);
nand I_54916 (I935710,I936225,I936109);
not I_54917 (I936314,I2690);
DFFARX1 I_54918 (I550329,I2683,I936314,I936340,);
and I_54919 (I936348,I936340,I550317);
DFFARX1 I_54920 (I936348,I2683,I936314,I936297,);
DFFARX1 I_54921 (I550320,I2683,I936314,I936388,);
not I_54922 (I936396,I550314);
not I_54923 (I936413,I550338);
nand I_54924 (I936430,I936413,I936396);
nor I_54925 (I936285,I936388,I936430);
DFFARX1 I_54926 (I936430,I2683,I936314,I936470,);
not I_54927 (I936306,I936470);
not I_54928 (I936492,I550326);
nand I_54929 (I936509,I936413,I936492);
DFFARX1 I_54930 (I936509,I2683,I936314,I936535,);
not I_54931 (I936543,I936535);
not I_54932 (I936560,I550335);
nand I_54933 (I936577,I936560,I550332);
and I_54934 (I936594,I936396,I936577);
nor I_54935 (I936611,I936509,I936594);
DFFARX1 I_54936 (I936611,I2683,I936314,I936282,);
DFFARX1 I_54937 (I936594,I2683,I936314,I936303,);
nor I_54938 (I936656,I550335,I550323);
nor I_54939 (I936294,I936509,I936656);
or I_54940 (I936687,I550335,I550323);
nor I_54941 (I936704,I550314,I550317);
DFFARX1 I_54942 (I936704,I2683,I936314,I936730,);
not I_54943 (I936738,I936730);
nor I_54944 (I936300,I936738,I936543);
nand I_54945 (I936769,I936738,I936388);
not I_54946 (I936786,I550314);
nand I_54947 (I936803,I936786,I936492);
nand I_54948 (I936820,I936738,I936803);
nand I_54949 (I936291,I936820,I936769);
nand I_54950 (I936288,I936803,I936687);
not I_54951 (I936892,I2690);
DFFARX1 I_54952 (I311270,I2683,I936892,I936918,);
and I_54953 (I936926,I936918,I311255);
DFFARX1 I_54954 (I936926,I2683,I936892,I936875,);
DFFARX1 I_54955 (I311261,I2683,I936892,I936966,);
not I_54956 (I936974,I311243);
not I_54957 (I936991,I311264);
nand I_54958 (I937008,I936991,I936974);
nor I_54959 (I936863,I936966,I937008);
DFFARX1 I_54960 (I937008,I2683,I936892,I937048,);
not I_54961 (I936884,I937048);
not I_54962 (I937070,I311267);
nand I_54963 (I937087,I936991,I937070);
DFFARX1 I_54964 (I937087,I2683,I936892,I937113,);
not I_54965 (I937121,I937113);
not I_54966 (I937138,I311258);
nand I_54967 (I937155,I937138,I311246);
and I_54968 (I937172,I936974,I937155);
nor I_54969 (I937189,I937087,I937172);
DFFARX1 I_54970 (I937189,I2683,I936892,I936860,);
DFFARX1 I_54971 (I937172,I2683,I936892,I936881,);
nor I_54972 (I937234,I311258,I311252);
nor I_54973 (I936872,I937087,I937234);
or I_54974 (I937265,I311258,I311252);
nor I_54975 (I937282,I311249,I311243);
DFFARX1 I_54976 (I937282,I2683,I936892,I937308,);
not I_54977 (I937316,I937308);
nor I_54978 (I936878,I937316,I937121);
nand I_54979 (I937347,I937316,I936966);
not I_54980 (I937364,I311249);
nand I_54981 (I937381,I937364,I937070);
nand I_54982 (I937398,I937316,I937381);
nand I_54983 (I936869,I937398,I937347);
nand I_54984 (I936866,I937381,I937265);
not I_54985 (I937470,I2690);
DFFARX1 I_54986 (I794933,I2683,I937470,I937496,);
and I_54987 (I937504,I937496,I794927);
DFFARX1 I_54988 (I937504,I2683,I937470,I937453,);
DFFARX1 I_54989 (I794945,I2683,I937470,I937544,);
not I_54990 (I937552,I794936);
not I_54991 (I937569,I794948);
nand I_54992 (I937586,I937569,I937552);
nor I_54993 (I937441,I937544,I937586);
DFFARX1 I_54994 (I937586,I2683,I937470,I937626,);
not I_54995 (I937462,I937626);
not I_54996 (I937648,I794954);
nand I_54997 (I937665,I937569,I937648);
DFFARX1 I_54998 (I937665,I2683,I937470,I937691,);
not I_54999 (I937699,I937691);
not I_55000 (I937716,I794930);
nand I_55001 (I937733,I937716,I794951);
and I_55002 (I937750,I937552,I937733);
nor I_55003 (I937767,I937665,I937750);
DFFARX1 I_55004 (I937767,I2683,I937470,I937438,);
DFFARX1 I_55005 (I937750,I2683,I937470,I937459,);
nor I_55006 (I937812,I794930,I794942);
nor I_55007 (I937450,I937665,I937812);
or I_55008 (I937843,I794930,I794942);
nor I_55009 (I937860,I794927,I794939);
DFFARX1 I_55010 (I937860,I2683,I937470,I937886,);
not I_55011 (I937894,I937886);
nor I_55012 (I937456,I937894,I937699);
nand I_55013 (I937925,I937894,I937544);
not I_55014 (I937942,I794927);
nand I_55015 (I937959,I937942,I937648);
nand I_55016 (I937976,I937894,I937959);
nand I_55017 (I937447,I937976,I937925);
nand I_55018 (I937444,I937959,I937843);
not I_55019 (I938048,I2690);
DFFARX1 I_55020 (I995534,I2683,I938048,I938074,);
and I_55021 (I938082,I938074,I995516);
DFFARX1 I_55022 (I938082,I2683,I938048,I938031,);
DFFARX1 I_55023 (I995525,I2683,I938048,I938122,);
not I_55024 (I938130,I995510);
not I_55025 (I938147,I995522);
nand I_55026 (I938164,I938147,I938130);
nor I_55027 (I938019,I938122,I938164);
DFFARX1 I_55028 (I938164,I2683,I938048,I938204,);
not I_55029 (I938040,I938204);
not I_55030 (I938226,I995513);
nand I_55031 (I938243,I938147,I938226);
DFFARX1 I_55032 (I938243,I2683,I938048,I938269,);
not I_55033 (I938277,I938269);
not I_55034 (I938294,I995510);
nand I_55035 (I938311,I938294,I995513);
and I_55036 (I938328,I938130,I938311);
nor I_55037 (I938345,I938243,I938328);
DFFARX1 I_55038 (I938345,I2683,I938048,I938016,);
DFFARX1 I_55039 (I938328,I2683,I938048,I938037,);
nor I_55040 (I938390,I995510,I995531);
nor I_55041 (I938028,I938243,I938390);
or I_55042 (I938421,I995510,I995531);
nor I_55043 (I938438,I995519,I995528);
DFFARX1 I_55044 (I938438,I2683,I938048,I938464,);
not I_55045 (I938472,I938464);
nor I_55046 (I938034,I938472,I938277);
nand I_55047 (I938503,I938472,I938122);
not I_55048 (I938520,I995519);
nand I_55049 (I938537,I938520,I938226);
nand I_55050 (I938554,I938472,I938537);
nand I_55051 (I938025,I938554,I938503);
nand I_55052 (I938022,I938537,I938421);
not I_55053 (I938626,I2690);
DFFARX1 I_55054 (I506979,I2683,I938626,I938652,);
and I_55055 (I938660,I938652,I506967);
DFFARX1 I_55056 (I938660,I2683,I938626,I938609,);
DFFARX1 I_55057 (I506970,I2683,I938626,I938700,);
not I_55058 (I938708,I506964);
not I_55059 (I938725,I506988);
nand I_55060 (I938742,I938725,I938708);
nor I_55061 (I938597,I938700,I938742);
DFFARX1 I_55062 (I938742,I2683,I938626,I938782,);
not I_55063 (I938618,I938782);
not I_55064 (I938804,I506976);
nand I_55065 (I938821,I938725,I938804);
DFFARX1 I_55066 (I938821,I2683,I938626,I938847,);
not I_55067 (I938855,I938847);
not I_55068 (I938872,I506985);
nand I_55069 (I938889,I938872,I506982);
and I_55070 (I938906,I938708,I938889);
nor I_55071 (I938923,I938821,I938906);
DFFARX1 I_55072 (I938923,I2683,I938626,I938594,);
DFFARX1 I_55073 (I938906,I2683,I938626,I938615,);
nor I_55074 (I938968,I506985,I506973);
nor I_55075 (I938606,I938821,I938968);
or I_55076 (I938999,I506985,I506973);
nor I_55077 (I939016,I506964,I506967);
DFFARX1 I_55078 (I939016,I2683,I938626,I939042,);
not I_55079 (I939050,I939042);
nor I_55080 (I938612,I939050,I938855);
nand I_55081 (I939081,I939050,I938700);
not I_55082 (I939098,I506964);
nand I_55083 (I939115,I939098,I938804);
nand I_55084 (I939132,I939050,I939115);
nand I_55085 (I938603,I939132,I939081);
nand I_55086 (I938600,I939115,I938999);
not I_55087 (I939204,I2690);
DFFARX1 I_55088 (I393778,I2683,I939204,I939230,);
and I_55089 (I939238,I939230,I393793);
DFFARX1 I_55090 (I939238,I2683,I939204,I939187,);
DFFARX1 I_55091 (I393796,I2683,I939204,I939278,);
not I_55092 (I939286,I393790);
not I_55093 (I939303,I393805);
nand I_55094 (I939320,I939303,I939286);
nor I_55095 (I939175,I939278,I939320);
DFFARX1 I_55096 (I939320,I2683,I939204,I939360,);
not I_55097 (I939196,I939360);
not I_55098 (I939382,I393781);
nand I_55099 (I939399,I939303,I939382);
DFFARX1 I_55100 (I939399,I2683,I939204,I939425,);
not I_55101 (I939433,I939425);
not I_55102 (I939450,I393784);
nand I_55103 (I939467,I939450,I393778);
and I_55104 (I939484,I939286,I939467);
nor I_55105 (I939501,I939399,I939484);
DFFARX1 I_55106 (I939501,I2683,I939204,I939172,);
DFFARX1 I_55107 (I939484,I2683,I939204,I939193,);
nor I_55108 (I939546,I393784,I393787);
nor I_55109 (I939184,I939399,I939546);
or I_55110 (I939577,I393784,I393787);
nor I_55111 (I939594,I393802,I393799);
DFFARX1 I_55112 (I939594,I2683,I939204,I939620,);
not I_55113 (I939628,I939620);
nor I_55114 (I939190,I939628,I939433);
nand I_55115 (I939659,I939628,I939278);
not I_55116 (I939676,I393802);
nand I_55117 (I939693,I939676,I939382);
nand I_55118 (I939710,I939628,I939693);
nand I_55119 (I939181,I939710,I939659);
nand I_55120 (I939178,I939693,I939577);
not I_55121 (I939782,I2690);
DFFARX1 I_55122 (I35333,I2683,I939782,I939808,);
and I_55123 (I939816,I939808,I35336);
DFFARX1 I_55124 (I939816,I2683,I939782,I939765,);
DFFARX1 I_55125 (I35336,I2683,I939782,I939856,);
not I_55126 (I939864,I35339);
not I_55127 (I939881,I35354);
nand I_55128 (I939898,I939881,I939864);
nor I_55129 (I939753,I939856,I939898);
DFFARX1 I_55130 (I939898,I2683,I939782,I939938,);
not I_55131 (I939774,I939938);
not I_55132 (I939960,I35348);
nand I_55133 (I939977,I939881,I939960);
DFFARX1 I_55134 (I939977,I2683,I939782,I940003,);
not I_55135 (I940011,I940003);
not I_55136 (I940028,I35351);
nand I_55137 (I940045,I940028,I35333);
and I_55138 (I940062,I939864,I940045);
nor I_55139 (I940079,I939977,I940062);
DFFARX1 I_55140 (I940079,I2683,I939782,I939750,);
DFFARX1 I_55141 (I940062,I2683,I939782,I939771,);
nor I_55142 (I940124,I35351,I35345);
nor I_55143 (I939762,I939977,I940124);
or I_55144 (I940155,I35351,I35345);
nor I_55145 (I940172,I35342,I35357);
DFFARX1 I_55146 (I940172,I2683,I939782,I940198,);
not I_55147 (I940206,I940198);
nor I_55148 (I939768,I940206,I940011);
nand I_55149 (I940237,I940206,I939856);
not I_55150 (I940254,I35342);
nand I_55151 (I940271,I940254,I939960);
nand I_55152 (I940288,I940206,I940271);
nand I_55153 (I939759,I940288,I940237);
nand I_55154 (I939756,I940271,I940155);
not I_55155 (I940360,I2690);
DFFARX1 I_55156 (I225369,I2683,I940360,I940386,);
and I_55157 (I940394,I940386,I225354);
DFFARX1 I_55158 (I940394,I2683,I940360,I940343,);
DFFARX1 I_55159 (I225360,I2683,I940360,I940434,);
not I_55160 (I940442,I225342);
not I_55161 (I940459,I225363);
nand I_55162 (I940476,I940459,I940442);
nor I_55163 (I940331,I940434,I940476);
DFFARX1 I_55164 (I940476,I2683,I940360,I940516,);
not I_55165 (I940352,I940516);
not I_55166 (I940538,I225366);
nand I_55167 (I940555,I940459,I940538);
DFFARX1 I_55168 (I940555,I2683,I940360,I940581,);
not I_55169 (I940589,I940581);
not I_55170 (I940606,I225357);
nand I_55171 (I940623,I940606,I225345);
and I_55172 (I940640,I940442,I940623);
nor I_55173 (I940657,I940555,I940640);
DFFARX1 I_55174 (I940657,I2683,I940360,I940328,);
DFFARX1 I_55175 (I940640,I2683,I940360,I940349,);
nor I_55176 (I940702,I225357,I225351);
nor I_55177 (I940340,I940555,I940702);
or I_55178 (I940733,I225357,I225351);
nor I_55179 (I940750,I225348,I225342);
DFFARX1 I_55180 (I940750,I2683,I940360,I940776,);
not I_55181 (I940784,I940776);
nor I_55182 (I940346,I940784,I940589);
nand I_55183 (I940815,I940784,I940434);
not I_55184 (I940832,I225348);
nand I_55185 (I940849,I940832,I940538);
nand I_55186 (I940866,I940784,I940849);
nand I_55187 (I940337,I940866,I940815);
nand I_55188 (I940334,I940849,I940733);
not I_55189 (I940938,I2690);
DFFARX1 I_55190 (I133100,I2683,I940938,I940964,);
and I_55191 (I940972,I940964,I133103);
DFFARX1 I_55192 (I940972,I2683,I940938,I940921,);
DFFARX1 I_55193 (I133103,I2683,I940938,I941012,);
not I_55194 (I941020,I133118);
not I_55195 (I941037,I133124);
nand I_55196 (I941054,I941037,I941020);
nor I_55197 (I940909,I941012,I941054);
DFFARX1 I_55198 (I941054,I2683,I940938,I941094,);
not I_55199 (I940930,I941094);
not I_55200 (I941116,I133112);
nand I_55201 (I941133,I941037,I941116);
DFFARX1 I_55202 (I941133,I2683,I940938,I941159,);
not I_55203 (I941167,I941159);
not I_55204 (I941184,I133109);
nand I_55205 (I941201,I941184,I133106);
and I_55206 (I941218,I941020,I941201);
nor I_55207 (I941235,I941133,I941218);
DFFARX1 I_55208 (I941235,I2683,I940938,I940906,);
DFFARX1 I_55209 (I941218,I2683,I940938,I940927,);
nor I_55210 (I941280,I133109,I133100);
nor I_55211 (I940918,I941133,I941280);
or I_55212 (I941311,I133109,I133100);
nor I_55213 (I941328,I133115,I133121);
DFFARX1 I_55214 (I941328,I2683,I940938,I941354,);
not I_55215 (I941362,I941354);
nor I_55216 (I940924,I941362,I941167);
nand I_55217 (I941393,I941362,I941012);
not I_55218 (I941410,I133115);
nand I_55219 (I941427,I941410,I941116);
nand I_55220 (I941444,I941362,I941427);
nand I_55221 (I940915,I941444,I941393);
nand I_55222 (I940912,I941427,I941311);
not I_55223 (I941516,I2690);
DFFARX1 I_55224 (I24266,I2683,I941516,I941542,);
and I_55225 (I941550,I941542,I24269);
DFFARX1 I_55226 (I941550,I2683,I941516,I941499,);
DFFARX1 I_55227 (I24269,I2683,I941516,I941590,);
not I_55228 (I941598,I24272);
not I_55229 (I941615,I24287);
nand I_55230 (I941632,I941615,I941598);
nor I_55231 (I941487,I941590,I941632);
DFFARX1 I_55232 (I941632,I2683,I941516,I941672,);
not I_55233 (I941508,I941672);
not I_55234 (I941694,I24281);
nand I_55235 (I941711,I941615,I941694);
DFFARX1 I_55236 (I941711,I2683,I941516,I941737,);
not I_55237 (I941745,I941737);
not I_55238 (I941762,I24284);
nand I_55239 (I941779,I941762,I24266);
and I_55240 (I941796,I941598,I941779);
nor I_55241 (I941813,I941711,I941796);
DFFARX1 I_55242 (I941813,I2683,I941516,I941484,);
DFFARX1 I_55243 (I941796,I2683,I941516,I941505,);
nor I_55244 (I941858,I24284,I24278);
nor I_55245 (I941496,I941711,I941858);
or I_55246 (I941889,I24284,I24278);
nor I_55247 (I941906,I24275,I24290);
DFFARX1 I_55248 (I941906,I2683,I941516,I941932,);
not I_55249 (I941940,I941932);
nor I_55250 (I941502,I941940,I941745);
nand I_55251 (I941971,I941940,I941590);
not I_55252 (I941988,I24275);
nand I_55253 (I942005,I941988,I941694);
nand I_55254 (I942022,I941940,I942005);
nand I_55255 (I941493,I942022,I941971);
nand I_55256 (I941490,I942005,I941889);
not I_55257 (I942094,I2690);
DFFARX1 I_55258 (I1060256,I2683,I942094,I942120,);
and I_55259 (I942128,I942120,I1060238);
DFFARX1 I_55260 (I942128,I2683,I942094,I942077,);
DFFARX1 I_55261 (I1060229,I2683,I942094,I942168,);
not I_55262 (I942176,I1060244);
not I_55263 (I942193,I1060232);
nand I_55264 (I942210,I942193,I942176);
nor I_55265 (I942065,I942168,I942210);
DFFARX1 I_55266 (I942210,I2683,I942094,I942250,);
not I_55267 (I942086,I942250);
not I_55268 (I942272,I1060241);
nand I_55269 (I942289,I942193,I942272);
DFFARX1 I_55270 (I942289,I2683,I942094,I942315,);
not I_55271 (I942323,I942315);
not I_55272 (I942340,I1060250);
nand I_55273 (I942357,I942340,I1060229);
and I_55274 (I942374,I942176,I942357);
nor I_55275 (I942391,I942289,I942374);
DFFARX1 I_55276 (I942391,I2683,I942094,I942062,);
DFFARX1 I_55277 (I942374,I2683,I942094,I942083,);
nor I_55278 (I942436,I1060250,I1060253);
nor I_55279 (I942074,I942289,I942436);
or I_55280 (I942467,I1060250,I1060253);
nor I_55281 (I942484,I1060247,I1060235);
DFFARX1 I_55282 (I942484,I2683,I942094,I942510,);
not I_55283 (I942518,I942510);
nor I_55284 (I942080,I942518,I942323);
nand I_55285 (I942549,I942518,I942168);
not I_55286 (I942566,I1060247);
nand I_55287 (I942583,I942566,I942272);
nand I_55288 (I942600,I942518,I942583);
nand I_55289 (I942071,I942600,I942549);
nand I_55290 (I942068,I942583,I942467);
not I_55291 (I942672,I2690);
DFFARX1 I_55292 (I343186,I2683,I942672,I942698,);
and I_55293 (I942706,I942698,I343201);
DFFARX1 I_55294 (I942706,I2683,I942672,I942655,);
DFFARX1 I_55295 (I343204,I2683,I942672,I942746,);
not I_55296 (I942754,I343198);
not I_55297 (I942771,I343213);
nand I_55298 (I942788,I942771,I942754);
nor I_55299 (I942643,I942746,I942788);
DFFARX1 I_55300 (I942788,I2683,I942672,I942828,);
not I_55301 (I942664,I942828);
not I_55302 (I942850,I343189);
nand I_55303 (I942867,I942771,I942850);
DFFARX1 I_55304 (I942867,I2683,I942672,I942893,);
not I_55305 (I942901,I942893);
not I_55306 (I942918,I343192);
nand I_55307 (I942935,I942918,I343186);
and I_55308 (I942952,I942754,I942935);
nor I_55309 (I942969,I942867,I942952);
DFFARX1 I_55310 (I942969,I2683,I942672,I942640,);
DFFARX1 I_55311 (I942952,I2683,I942672,I942661,);
nor I_55312 (I943014,I343192,I343195);
nor I_55313 (I942652,I942867,I943014);
or I_55314 (I943045,I343192,I343195);
nor I_55315 (I943062,I343210,I343207);
DFFARX1 I_55316 (I943062,I2683,I942672,I943088,);
not I_55317 (I943096,I943088);
nor I_55318 (I942658,I943096,I942901);
nand I_55319 (I943127,I943096,I942746);
not I_55320 (I943144,I343210);
nand I_55321 (I943161,I943144,I942850);
nand I_55322 (I943178,I943096,I943161);
nand I_55323 (I942649,I943178,I943127);
nand I_55324 (I942646,I943161,I943045);
not I_55325 (I943250,I2690);
DFFARX1 I_55326 (I1069181,I2683,I943250,I943276,);
and I_55327 (I943284,I943276,I1069163);
DFFARX1 I_55328 (I943284,I2683,I943250,I943233,);
DFFARX1 I_55329 (I1069154,I2683,I943250,I943324,);
not I_55330 (I943332,I1069169);
not I_55331 (I943349,I1069157);
nand I_55332 (I943366,I943349,I943332);
nor I_55333 (I943221,I943324,I943366);
DFFARX1 I_55334 (I943366,I2683,I943250,I943406,);
not I_55335 (I943242,I943406);
not I_55336 (I943428,I1069166);
nand I_55337 (I943445,I943349,I943428);
DFFARX1 I_55338 (I943445,I2683,I943250,I943471,);
not I_55339 (I943479,I943471);
not I_55340 (I943496,I1069175);
nand I_55341 (I943513,I943496,I1069154);
and I_55342 (I943530,I943332,I943513);
nor I_55343 (I943547,I943445,I943530);
DFFARX1 I_55344 (I943547,I2683,I943250,I943218,);
DFFARX1 I_55345 (I943530,I2683,I943250,I943239,);
nor I_55346 (I943592,I1069175,I1069178);
nor I_55347 (I943230,I943445,I943592);
or I_55348 (I943623,I1069175,I1069178);
nor I_55349 (I943640,I1069172,I1069160);
DFFARX1 I_55350 (I943640,I2683,I943250,I943666,);
not I_55351 (I943674,I943666);
nor I_55352 (I943236,I943674,I943479);
nand I_55353 (I943705,I943674,I943324);
not I_55354 (I943722,I1069172);
nand I_55355 (I943739,I943722,I943428);
nand I_55356 (I943756,I943674,I943739);
nand I_55357 (I943227,I943756,I943705);
nand I_55358 (I943224,I943739,I943623);
not I_55359 (I943828,I2690);
DFFARX1 I_55360 (I623315,I2683,I943828,I943854,);
and I_55361 (I943862,I943854,I623321);
DFFARX1 I_55362 (I943862,I2683,I943828,I943811,);
DFFARX1 I_55363 (I623327,I2683,I943828,I943902,);
not I_55364 (I943910,I623312);
not I_55365 (I943927,I623312);
nand I_55366 (I943944,I943927,I943910);
nor I_55367 (I943799,I943902,I943944);
DFFARX1 I_55368 (I943944,I2683,I943828,I943984,);
not I_55369 (I943820,I943984);
not I_55370 (I944006,I623330);
nand I_55371 (I944023,I943927,I944006);
DFFARX1 I_55372 (I944023,I2683,I943828,I944049,);
not I_55373 (I944057,I944049);
not I_55374 (I944074,I623324);
nand I_55375 (I944091,I944074,I623315);
and I_55376 (I944108,I943910,I944091);
nor I_55377 (I944125,I944023,I944108);
DFFARX1 I_55378 (I944125,I2683,I943828,I943796,);
DFFARX1 I_55379 (I944108,I2683,I943828,I943817,);
nor I_55380 (I944170,I623324,I623333);
nor I_55381 (I943808,I944023,I944170);
or I_55382 (I944201,I623324,I623333);
nor I_55383 (I944218,I623318,I623318);
DFFARX1 I_55384 (I944218,I2683,I943828,I944244,);
not I_55385 (I944252,I944244);
nor I_55386 (I943814,I944252,I944057);
nand I_55387 (I944283,I944252,I943902);
not I_55388 (I944300,I623318);
nand I_55389 (I944317,I944300,I944006);
nand I_55390 (I944334,I944252,I944317);
nand I_55391 (I943805,I944334,I944283);
nand I_55392 (I943802,I944317,I944201);
not I_55393 (I944406,I2690);
DFFARX1 I_55394 (I349714,I2683,I944406,I944432,);
and I_55395 (I944440,I944432,I349729);
DFFARX1 I_55396 (I944440,I2683,I944406,I944389,);
DFFARX1 I_55397 (I349732,I2683,I944406,I944480,);
not I_55398 (I944488,I349726);
not I_55399 (I944505,I349741);
nand I_55400 (I944522,I944505,I944488);
nor I_55401 (I944377,I944480,I944522);
DFFARX1 I_55402 (I944522,I2683,I944406,I944562,);
not I_55403 (I944398,I944562);
not I_55404 (I944584,I349717);
nand I_55405 (I944601,I944505,I944584);
DFFARX1 I_55406 (I944601,I2683,I944406,I944627,);
not I_55407 (I944635,I944627);
not I_55408 (I944652,I349720);
nand I_55409 (I944669,I944652,I349714);
and I_55410 (I944686,I944488,I944669);
nor I_55411 (I944703,I944601,I944686);
DFFARX1 I_55412 (I944703,I2683,I944406,I944374,);
DFFARX1 I_55413 (I944686,I2683,I944406,I944395,);
nor I_55414 (I944748,I349720,I349723);
nor I_55415 (I944386,I944601,I944748);
or I_55416 (I944779,I349720,I349723);
nor I_55417 (I944796,I349738,I349735);
DFFARX1 I_55418 (I944796,I2683,I944406,I944822,);
not I_55419 (I944830,I944822);
nor I_55420 (I944392,I944830,I944635);
nand I_55421 (I944861,I944830,I944480);
not I_55422 (I944878,I349738);
nand I_55423 (I944895,I944878,I944584);
nand I_55424 (I944912,I944830,I944895);
nand I_55425 (I944383,I944912,I944861);
nand I_55426 (I944380,I944895,I944779);
not I_55427 (I944984,I2690);
DFFARX1 I_55428 (I253300,I2683,I944984,I945010,);
and I_55429 (I945018,I945010,I253285);
DFFARX1 I_55430 (I945018,I2683,I944984,I944967,);
DFFARX1 I_55431 (I253291,I2683,I944984,I945058,);
not I_55432 (I945066,I253273);
not I_55433 (I945083,I253294);
nand I_55434 (I945100,I945083,I945066);
nor I_55435 (I944955,I945058,I945100);
DFFARX1 I_55436 (I945100,I2683,I944984,I945140,);
not I_55437 (I944976,I945140);
not I_55438 (I945162,I253297);
nand I_55439 (I945179,I945083,I945162);
DFFARX1 I_55440 (I945179,I2683,I944984,I945205,);
not I_55441 (I945213,I945205);
not I_55442 (I945230,I253288);
nand I_55443 (I945247,I945230,I253276);
and I_55444 (I945264,I945066,I945247);
nor I_55445 (I945281,I945179,I945264);
DFFARX1 I_55446 (I945281,I2683,I944984,I944952,);
DFFARX1 I_55447 (I945264,I2683,I944984,I944973,);
nor I_55448 (I945326,I253288,I253282);
nor I_55449 (I944964,I945179,I945326);
or I_55450 (I945357,I253288,I253282);
nor I_55451 (I945374,I253279,I253273);
DFFARX1 I_55452 (I945374,I2683,I944984,I945400,);
not I_55453 (I945408,I945400);
nor I_55454 (I944970,I945408,I945213);
nand I_55455 (I945439,I945408,I945058);
not I_55456 (I945456,I253279);
nand I_55457 (I945473,I945456,I945162);
nand I_55458 (I945490,I945408,I945473);
nand I_55459 (I944961,I945490,I945439);
nand I_55460 (I944958,I945473,I945357);
not I_55461 (I945562,I2690);
DFFARX1 I_55462 (I111245,I2683,I945562,I945588,);
and I_55463 (I945596,I945588,I111221);
DFFARX1 I_55464 (I945596,I2683,I945562,I945545,);
DFFARX1 I_55465 (I111239,I2683,I945562,I945636,);
not I_55466 (I945644,I111227);
not I_55467 (I945661,I111224);
nand I_55468 (I945678,I945661,I945644);
nor I_55469 (I945533,I945636,I945678);
DFFARX1 I_55470 (I945678,I2683,I945562,I945718,);
not I_55471 (I945554,I945718);
not I_55472 (I945740,I111233);
nand I_55473 (I945757,I945661,I945740);
DFFARX1 I_55474 (I945757,I2683,I945562,I945783,);
not I_55475 (I945791,I945783);
not I_55476 (I945808,I111224);
nand I_55477 (I945825,I945808,I111242);
and I_55478 (I945842,I945644,I945825);
nor I_55479 (I945859,I945757,I945842);
DFFARX1 I_55480 (I945859,I2683,I945562,I945530,);
DFFARX1 I_55481 (I945842,I2683,I945562,I945551,);
nor I_55482 (I945904,I111224,I111236);
nor I_55483 (I945542,I945757,I945904);
or I_55484 (I945935,I111224,I111236);
nor I_55485 (I945952,I111230,I111221);
DFFARX1 I_55486 (I945952,I2683,I945562,I945978,);
not I_55487 (I945986,I945978);
nor I_55488 (I945548,I945986,I945791);
nand I_55489 (I946017,I945986,I945636);
not I_55490 (I946034,I111230);
nand I_55491 (I946051,I946034,I945740);
nand I_55492 (I946068,I945986,I946051);
nand I_55493 (I945539,I946068,I946017);
nand I_55494 (I945536,I946051,I945935);
not I_55495 (I946140,I2690);
DFFARX1 I_55496 (I340466,I2683,I946140,I946166,);
and I_55497 (I946174,I946166,I340481);
DFFARX1 I_55498 (I946174,I2683,I946140,I946123,);
DFFARX1 I_55499 (I340484,I2683,I946140,I946214,);
not I_55500 (I946222,I340478);
not I_55501 (I946239,I340493);
nand I_55502 (I946256,I946239,I946222);
nor I_55503 (I946111,I946214,I946256);
DFFARX1 I_55504 (I946256,I2683,I946140,I946296,);
not I_55505 (I946132,I946296);
not I_55506 (I946318,I340469);
nand I_55507 (I946335,I946239,I946318);
DFFARX1 I_55508 (I946335,I2683,I946140,I946361,);
not I_55509 (I946369,I946361);
not I_55510 (I946386,I340472);
nand I_55511 (I946403,I946386,I340466);
and I_55512 (I946420,I946222,I946403);
nor I_55513 (I946437,I946335,I946420);
DFFARX1 I_55514 (I946437,I2683,I946140,I946108,);
DFFARX1 I_55515 (I946420,I2683,I946140,I946129,);
nor I_55516 (I946482,I340472,I340475);
nor I_55517 (I946120,I946335,I946482);
or I_55518 (I946513,I340472,I340475);
nor I_55519 (I946530,I340490,I340487);
DFFARX1 I_55520 (I946530,I2683,I946140,I946556,);
not I_55521 (I946564,I946556);
nor I_55522 (I946126,I946564,I946369);
nand I_55523 (I946595,I946564,I946214);
not I_55524 (I946612,I340490);
nand I_55525 (I946629,I946612,I946318);
nand I_55526 (I946646,I946564,I946629);
nand I_55527 (I946117,I946646,I946595);
nand I_55528 (I946114,I946629,I946513);
not I_55529 (I946718,I2690);
DFFARX1 I_55530 (I770385,I2683,I946718,I946744,);
and I_55531 (I946752,I946744,I770379);
DFFARX1 I_55532 (I946752,I2683,I946718,I946701,);
DFFARX1 I_55533 (I770397,I2683,I946718,I946792,);
not I_55534 (I946800,I770388);
not I_55535 (I946817,I770400);
nand I_55536 (I946834,I946817,I946800);
nor I_55537 (I946689,I946792,I946834);
DFFARX1 I_55538 (I946834,I2683,I946718,I946874,);
not I_55539 (I946710,I946874);
not I_55540 (I946896,I770406);
nand I_55541 (I946913,I946817,I946896);
DFFARX1 I_55542 (I946913,I2683,I946718,I946939,);
not I_55543 (I946947,I946939);
not I_55544 (I946964,I770382);
nand I_55545 (I946981,I946964,I770403);
and I_55546 (I946998,I946800,I946981);
nor I_55547 (I947015,I946913,I946998);
DFFARX1 I_55548 (I947015,I2683,I946718,I946686,);
DFFARX1 I_55549 (I946998,I2683,I946718,I946707,);
nor I_55550 (I947060,I770382,I770394);
nor I_55551 (I946698,I946913,I947060);
or I_55552 (I947091,I770382,I770394);
nor I_55553 (I947108,I770379,I770391);
DFFARX1 I_55554 (I947108,I2683,I946718,I947134,);
not I_55555 (I947142,I947134);
nor I_55556 (I946704,I947142,I946947);
nand I_55557 (I947173,I947142,I946792);
not I_55558 (I947190,I770379);
nand I_55559 (I947207,I947190,I946896);
nand I_55560 (I947224,I947142,I947207);
nand I_55561 (I946695,I947224,I947173);
nand I_55562 (I946692,I947207,I947091);
not I_55563 (I947296,I2690);
DFFARX1 I_55564 (I787181,I2683,I947296,I947322,);
and I_55565 (I947330,I947322,I787175);
DFFARX1 I_55566 (I947330,I2683,I947296,I947279,);
DFFARX1 I_55567 (I787193,I2683,I947296,I947370,);
not I_55568 (I947378,I787184);
not I_55569 (I947395,I787196);
nand I_55570 (I947412,I947395,I947378);
nor I_55571 (I947267,I947370,I947412);
DFFARX1 I_55572 (I947412,I2683,I947296,I947452,);
not I_55573 (I947288,I947452);
not I_55574 (I947474,I787202);
nand I_55575 (I947491,I947395,I947474);
DFFARX1 I_55576 (I947491,I2683,I947296,I947517,);
not I_55577 (I947525,I947517);
not I_55578 (I947542,I787178);
nand I_55579 (I947559,I947542,I787199);
and I_55580 (I947576,I947378,I947559);
nor I_55581 (I947593,I947491,I947576);
DFFARX1 I_55582 (I947593,I2683,I947296,I947264,);
DFFARX1 I_55583 (I947576,I2683,I947296,I947285,);
nor I_55584 (I947638,I787178,I787190);
nor I_55585 (I947276,I947491,I947638);
or I_55586 (I947669,I787178,I787190);
nor I_55587 (I947686,I787175,I787187);
DFFARX1 I_55588 (I947686,I2683,I947296,I947712,);
not I_55589 (I947720,I947712);
nor I_55590 (I947282,I947720,I947525);
nand I_55591 (I947751,I947720,I947370);
not I_55592 (I947768,I787175);
nand I_55593 (I947785,I947768,I947474);
nand I_55594 (I947802,I947720,I947785);
nand I_55595 (I947273,I947802,I947751);
nand I_55596 (I947270,I947785,I947669);
not I_55597 (I947874,I2690);
DFFARX1 I_55598 (I445133,I2683,I947874,I947900,);
and I_55599 (I947908,I947900,I445121);
DFFARX1 I_55600 (I947908,I2683,I947874,I947857,);
DFFARX1 I_55601 (I445136,I2683,I947874,I947948,);
not I_55602 (I947956,I445127);
not I_55603 (I947973,I445118);
nand I_55604 (I947990,I947973,I947956);
nor I_55605 (I947845,I947948,I947990);
DFFARX1 I_55606 (I947990,I2683,I947874,I948030,);
not I_55607 (I947866,I948030);
not I_55608 (I948052,I445124);
nand I_55609 (I948069,I947973,I948052);
DFFARX1 I_55610 (I948069,I2683,I947874,I948095,);
not I_55611 (I948103,I948095);
not I_55612 (I948120,I445139);
nand I_55613 (I948137,I948120,I445142);
and I_55614 (I948154,I947956,I948137);
nor I_55615 (I948171,I948069,I948154);
DFFARX1 I_55616 (I948171,I2683,I947874,I947842,);
DFFARX1 I_55617 (I948154,I2683,I947874,I947863,);
nor I_55618 (I948216,I445139,I445118);
nor I_55619 (I947854,I948069,I948216);
or I_55620 (I948247,I445139,I445118);
nor I_55621 (I948264,I445130,I445121);
DFFARX1 I_55622 (I948264,I2683,I947874,I948290,);
not I_55623 (I948298,I948290);
nor I_55624 (I947860,I948298,I948103);
nand I_55625 (I948329,I948298,I947948);
not I_55626 (I948346,I445130);
nand I_55627 (I948363,I948346,I948052);
nand I_55628 (I948380,I948298,I948363);
nand I_55629 (I947851,I948380,I948329);
nand I_55630 (I947848,I948363,I948247);
not I_55631 (I948452,I2690);
DFFARX1 I_55632 (I812491,I2683,I948452,I948478,);
and I_55633 (I948486,I948478,I812488);
DFFARX1 I_55634 (I948486,I2683,I948452,I948435,);
DFFARX1 I_55635 (I812494,I2683,I948452,I948526,);
not I_55636 (I948534,I812497);
not I_55637 (I948551,I812491);
nand I_55638 (I948568,I948551,I948534);
nor I_55639 (I948423,I948526,I948568);
DFFARX1 I_55640 (I948568,I2683,I948452,I948608,);
not I_55641 (I948444,I948608);
not I_55642 (I948630,I812506);
nand I_55643 (I948647,I948551,I948630);
DFFARX1 I_55644 (I948647,I2683,I948452,I948673,);
not I_55645 (I948681,I948673);
not I_55646 (I948698,I812503);
nand I_55647 (I948715,I948698,I812509);
and I_55648 (I948732,I948534,I948715);
nor I_55649 (I948749,I948647,I948732);
DFFARX1 I_55650 (I948749,I2683,I948452,I948420,);
DFFARX1 I_55651 (I948732,I2683,I948452,I948441,);
nor I_55652 (I948794,I812503,I812488);
nor I_55653 (I948432,I948647,I948794);
or I_55654 (I948825,I812503,I812488);
nor I_55655 (I948842,I812500,I812494);
DFFARX1 I_55656 (I948842,I2683,I948452,I948868,);
not I_55657 (I948876,I948868);
nor I_55658 (I948438,I948876,I948681);
nand I_55659 (I948907,I948876,I948526);
not I_55660 (I948924,I812500);
nand I_55661 (I948941,I948924,I948630);
nand I_55662 (I948958,I948876,I948941);
nand I_55663 (I948429,I948958,I948907);
nand I_55664 (I948426,I948941,I948825);
not I_55665 (I949030,I2690);
DFFARX1 I_55666 (I815296,I2683,I949030,I949056,);
and I_55667 (I949064,I949056,I815293);
DFFARX1 I_55668 (I949064,I2683,I949030,I949013,);
DFFARX1 I_55669 (I815299,I2683,I949030,I949104,);
not I_55670 (I949112,I815302);
not I_55671 (I949129,I815296);
nand I_55672 (I949146,I949129,I949112);
nor I_55673 (I949001,I949104,I949146);
DFFARX1 I_55674 (I949146,I2683,I949030,I949186,);
not I_55675 (I949022,I949186);
not I_55676 (I949208,I815311);
nand I_55677 (I949225,I949129,I949208);
DFFARX1 I_55678 (I949225,I2683,I949030,I949251,);
not I_55679 (I949259,I949251);
not I_55680 (I949276,I815308);
nand I_55681 (I949293,I949276,I815314);
and I_55682 (I949310,I949112,I949293);
nor I_55683 (I949327,I949225,I949310);
DFFARX1 I_55684 (I949327,I2683,I949030,I948998,);
DFFARX1 I_55685 (I949310,I2683,I949030,I949019,);
nor I_55686 (I949372,I815308,I815293);
nor I_55687 (I949010,I949225,I949372);
or I_55688 (I949403,I815308,I815293);
nor I_55689 (I949420,I815305,I815299);
DFFARX1 I_55690 (I949420,I2683,I949030,I949446,);
not I_55691 (I949454,I949446);
nor I_55692 (I949016,I949454,I949259);
nand I_55693 (I949485,I949454,I949104);
not I_55694 (I949502,I815305);
nand I_55695 (I949519,I949502,I949208);
nand I_55696 (I949536,I949454,I949519);
nand I_55697 (I949007,I949536,I949485);
nand I_55698 (I949004,I949519,I949403);
not I_55699 (I949608,I2690);
DFFARX1 I_55700 (I155115,I2683,I949608,I949634,);
and I_55701 (I949642,I949634,I155118);
DFFARX1 I_55702 (I949642,I2683,I949608,I949591,);
DFFARX1 I_55703 (I155118,I2683,I949608,I949682,);
not I_55704 (I949690,I155133);
not I_55705 (I949707,I155139);
nand I_55706 (I949724,I949707,I949690);
nor I_55707 (I949579,I949682,I949724);
DFFARX1 I_55708 (I949724,I2683,I949608,I949764,);
not I_55709 (I949600,I949764);
not I_55710 (I949786,I155127);
nand I_55711 (I949803,I949707,I949786);
DFFARX1 I_55712 (I949803,I2683,I949608,I949829,);
not I_55713 (I949837,I949829);
not I_55714 (I949854,I155124);
nand I_55715 (I949871,I949854,I155121);
and I_55716 (I949888,I949690,I949871);
nor I_55717 (I949905,I949803,I949888);
DFFARX1 I_55718 (I949905,I2683,I949608,I949576,);
DFFARX1 I_55719 (I949888,I2683,I949608,I949597,);
nor I_55720 (I949950,I155124,I155115);
nor I_55721 (I949588,I949803,I949950);
or I_55722 (I949981,I155124,I155115);
nor I_55723 (I949998,I155130,I155136);
DFFARX1 I_55724 (I949998,I2683,I949608,I950024,);
not I_55725 (I950032,I950024);
nor I_55726 (I949594,I950032,I949837);
nand I_55727 (I950063,I950032,I949682);
not I_55728 (I950080,I155130);
nand I_55729 (I950097,I950080,I949786);
nand I_55730 (I950114,I950032,I950097);
nand I_55731 (I949585,I950114,I950063);
nand I_55732 (I949582,I950097,I949981);
not I_55733 (I950186,I2690);
DFFARX1 I_55734 (I74882,I2683,I950186,I950212,);
and I_55735 (I950220,I950212,I74858);
DFFARX1 I_55736 (I950220,I2683,I950186,I950169,);
DFFARX1 I_55737 (I74876,I2683,I950186,I950260,);
not I_55738 (I950268,I74864);
not I_55739 (I950285,I74861);
nand I_55740 (I950302,I950285,I950268);
nor I_55741 (I950157,I950260,I950302);
DFFARX1 I_55742 (I950302,I2683,I950186,I950342,);
not I_55743 (I950178,I950342);
not I_55744 (I950364,I74870);
nand I_55745 (I950381,I950285,I950364);
DFFARX1 I_55746 (I950381,I2683,I950186,I950407,);
not I_55747 (I950415,I950407);
not I_55748 (I950432,I74861);
nand I_55749 (I950449,I950432,I74879);
and I_55750 (I950466,I950268,I950449);
nor I_55751 (I950483,I950381,I950466);
DFFARX1 I_55752 (I950483,I2683,I950186,I950154,);
DFFARX1 I_55753 (I950466,I2683,I950186,I950175,);
nor I_55754 (I950528,I74861,I74873);
nor I_55755 (I950166,I950381,I950528);
or I_55756 (I950559,I74861,I74873);
nor I_55757 (I950576,I74867,I74858);
DFFARX1 I_55758 (I950576,I2683,I950186,I950602,);
not I_55759 (I950610,I950602);
nor I_55760 (I950172,I950610,I950415);
nand I_55761 (I950641,I950610,I950260);
not I_55762 (I950658,I74867);
nand I_55763 (I950675,I950658,I950364);
nand I_55764 (I950692,I950610,I950675);
nand I_55765 (I950163,I950692,I950641);
nand I_55766 (I950160,I950675,I950559);
not I_55767 (I950764,I2690);
DFFARX1 I_55768 (I545705,I2683,I950764,I950790,);
and I_55769 (I950798,I950790,I545693);
DFFARX1 I_55770 (I950798,I2683,I950764,I950747,);
DFFARX1 I_55771 (I545696,I2683,I950764,I950838,);
not I_55772 (I950846,I545690);
not I_55773 (I950863,I545714);
nand I_55774 (I950880,I950863,I950846);
nor I_55775 (I950735,I950838,I950880);
DFFARX1 I_55776 (I950880,I2683,I950764,I950920,);
not I_55777 (I950756,I950920);
not I_55778 (I950942,I545702);
nand I_55779 (I950959,I950863,I950942);
DFFARX1 I_55780 (I950959,I2683,I950764,I950985,);
not I_55781 (I950993,I950985);
not I_55782 (I951010,I545711);
nand I_55783 (I951027,I951010,I545708);
and I_55784 (I951044,I950846,I951027);
nor I_55785 (I951061,I950959,I951044);
DFFARX1 I_55786 (I951061,I2683,I950764,I950732,);
DFFARX1 I_55787 (I951044,I2683,I950764,I950753,);
nor I_55788 (I951106,I545711,I545699);
nor I_55789 (I950744,I950959,I951106);
or I_55790 (I951137,I545711,I545699);
nor I_55791 (I951154,I545690,I545693);
DFFARX1 I_55792 (I951154,I2683,I950764,I951180,);
not I_55793 (I951188,I951180);
nor I_55794 (I950750,I951188,I950993);
nand I_55795 (I951219,I951188,I950838);
not I_55796 (I951236,I545690);
nand I_55797 (I951253,I951236,I950942);
nand I_55798 (I951270,I951188,I951253);
nand I_55799 (I950741,I951270,I951219);
nand I_55800 (I950738,I951253,I951137);
not I_55801 (I951342,I2690);
DFFARX1 I_55802 (I108083,I2683,I951342,I951368,);
and I_55803 (I951376,I951368,I108059);
DFFARX1 I_55804 (I951376,I2683,I951342,I951325,);
DFFARX1 I_55805 (I108077,I2683,I951342,I951416,);
not I_55806 (I951424,I108065);
not I_55807 (I951441,I108062);
nand I_55808 (I951458,I951441,I951424);
nor I_55809 (I951313,I951416,I951458);
DFFARX1 I_55810 (I951458,I2683,I951342,I951498,);
not I_55811 (I951334,I951498);
not I_55812 (I951520,I108071);
nand I_55813 (I951537,I951441,I951520);
DFFARX1 I_55814 (I951537,I2683,I951342,I951563,);
not I_55815 (I951571,I951563);
not I_55816 (I951588,I108062);
nand I_55817 (I951605,I951588,I108080);
and I_55818 (I951622,I951424,I951605);
nor I_55819 (I951639,I951537,I951622);
DFFARX1 I_55820 (I951639,I2683,I951342,I951310,);
DFFARX1 I_55821 (I951622,I2683,I951342,I951331,);
nor I_55822 (I951684,I108062,I108074);
nor I_55823 (I951322,I951537,I951684);
or I_55824 (I951715,I108062,I108074);
nor I_55825 (I951732,I108068,I108059);
DFFARX1 I_55826 (I951732,I2683,I951342,I951758,);
not I_55827 (I951766,I951758);
nor I_55828 (I951328,I951766,I951571);
nand I_55829 (I951797,I951766,I951416);
not I_55830 (I951814,I108068);
nand I_55831 (I951831,I951814,I951520);
nand I_55832 (I951848,I951766,I951831);
nand I_55833 (I951319,I951848,I951797);
nand I_55834 (I951316,I951831,I951715);
not I_55835 (I951920,I2690);
DFFARX1 I_55836 (I588477,I2683,I951920,I951946,);
and I_55837 (I951954,I951946,I588465);
DFFARX1 I_55838 (I951954,I2683,I951920,I951903,);
DFFARX1 I_55839 (I588468,I2683,I951920,I951994,);
not I_55840 (I952002,I588462);
not I_55841 (I952019,I588486);
nand I_55842 (I952036,I952019,I952002);
nor I_55843 (I951891,I951994,I952036);
DFFARX1 I_55844 (I952036,I2683,I951920,I952076,);
not I_55845 (I951912,I952076);
not I_55846 (I952098,I588474);
nand I_55847 (I952115,I952019,I952098);
DFFARX1 I_55848 (I952115,I2683,I951920,I952141,);
not I_55849 (I952149,I952141);
not I_55850 (I952166,I588483);
nand I_55851 (I952183,I952166,I588480);
and I_55852 (I952200,I952002,I952183);
nor I_55853 (I952217,I952115,I952200);
DFFARX1 I_55854 (I952217,I2683,I951920,I951888,);
DFFARX1 I_55855 (I952200,I2683,I951920,I951909,);
nor I_55856 (I952262,I588483,I588471);
nor I_55857 (I951900,I952115,I952262);
or I_55858 (I952293,I588483,I588471);
nor I_55859 (I952310,I588462,I588465);
DFFARX1 I_55860 (I952310,I2683,I951920,I952336,);
not I_55861 (I952344,I952336);
nor I_55862 (I951906,I952344,I952149);
nand I_55863 (I952375,I952344,I951994);
not I_55864 (I952392,I588462);
nand I_55865 (I952409,I952392,I952098);
nand I_55866 (I952426,I952344,I952409);
nand I_55867 (I951897,I952426,I952375);
nand I_55868 (I951894,I952409,I952293);
not I_55869 (I952498,I2690);
DFFARX1 I_55870 (I152735,I2683,I952498,I952524,);
and I_55871 (I952532,I952524,I152738);
DFFARX1 I_55872 (I952532,I2683,I952498,I952481,);
DFFARX1 I_55873 (I152738,I2683,I952498,I952572,);
not I_55874 (I952580,I152753);
not I_55875 (I952597,I152759);
nand I_55876 (I952614,I952597,I952580);
nor I_55877 (I952469,I952572,I952614);
DFFARX1 I_55878 (I952614,I2683,I952498,I952654,);
not I_55879 (I952490,I952654);
not I_55880 (I952676,I152747);
nand I_55881 (I952693,I952597,I952676);
DFFARX1 I_55882 (I952693,I2683,I952498,I952719,);
not I_55883 (I952727,I952719);
not I_55884 (I952744,I152744);
nand I_55885 (I952761,I952744,I152741);
and I_55886 (I952778,I952580,I952761);
nor I_55887 (I952795,I952693,I952778);
DFFARX1 I_55888 (I952795,I2683,I952498,I952466,);
DFFARX1 I_55889 (I952778,I2683,I952498,I952487,);
nor I_55890 (I952840,I152744,I152735);
nor I_55891 (I952478,I952693,I952840);
or I_55892 (I952871,I152744,I152735);
nor I_55893 (I952888,I152750,I152756);
DFFARX1 I_55894 (I952888,I2683,I952498,I952914,);
not I_55895 (I952922,I952914);
nor I_55896 (I952484,I952922,I952727);
nand I_55897 (I952953,I952922,I952572);
not I_55898 (I952970,I152750);
nand I_55899 (I952987,I952970,I952676);
nand I_55900 (I953004,I952922,I952987);
nand I_55901 (I952475,I953004,I952953);
nand I_55902 (I952472,I952987,I952871);
not I_55903 (I953076,I2690);
DFFARX1 I_55904 (I455537,I2683,I953076,I953102,);
and I_55905 (I953110,I953102,I455525);
DFFARX1 I_55906 (I953110,I2683,I953076,I953059,);
DFFARX1 I_55907 (I455540,I2683,I953076,I953150,);
not I_55908 (I953158,I455531);
not I_55909 (I953175,I455522);
nand I_55910 (I953192,I953175,I953158);
nor I_55911 (I953047,I953150,I953192);
DFFARX1 I_55912 (I953192,I2683,I953076,I953232,);
not I_55913 (I953068,I953232);
not I_55914 (I953254,I455528);
nand I_55915 (I953271,I953175,I953254);
DFFARX1 I_55916 (I953271,I2683,I953076,I953297,);
not I_55917 (I953305,I953297);
not I_55918 (I953322,I455543);
nand I_55919 (I953339,I953322,I455546);
and I_55920 (I953356,I953158,I953339);
nor I_55921 (I953373,I953271,I953356);
DFFARX1 I_55922 (I953373,I2683,I953076,I953044,);
DFFARX1 I_55923 (I953356,I2683,I953076,I953065,);
nor I_55924 (I953418,I455543,I455522);
nor I_55925 (I953056,I953271,I953418);
or I_55926 (I953449,I455543,I455522);
nor I_55927 (I953466,I455534,I455525);
DFFARX1 I_55928 (I953466,I2683,I953076,I953492,);
not I_55929 (I953500,I953492);
nor I_55930 (I953062,I953500,I953305);
nand I_55931 (I953531,I953500,I953150);
not I_55932 (I953548,I455534);
nand I_55933 (I953565,I953548,I953254);
nand I_55934 (I953582,I953500,I953565);
nand I_55935 (I953053,I953582,I953531);
nand I_55936 (I953050,I953565,I953449);
not I_55937 (I953654,I2690);
DFFARX1 I_55938 (I80152,I2683,I953654,I953680,);
and I_55939 (I953688,I953680,I80128);
DFFARX1 I_55940 (I953688,I2683,I953654,I953637,);
DFFARX1 I_55941 (I80146,I2683,I953654,I953728,);
not I_55942 (I953736,I80134);
not I_55943 (I953753,I80131);
nand I_55944 (I953770,I953753,I953736);
nor I_55945 (I953625,I953728,I953770);
DFFARX1 I_55946 (I953770,I2683,I953654,I953810,);
not I_55947 (I953646,I953810);
not I_55948 (I953832,I80140);
nand I_55949 (I953849,I953753,I953832);
DFFARX1 I_55950 (I953849,I2683,I953654,I953875,);
not I_55951 (I953883,I953875);
not I_55952 (I953900,I80131);
nand I_55953 (I953917,I953900,I80149);
and I_55954 (I953934,I953736,I953917);
nor I_55955 (I953951,I953849,I953934);
DFFARX1 I_55956 (I953951,I2683,I953654,I953622,);
DFFARX1 I_55957 (I953934,I2683,I953654,I953643,);
nor I_55958 (I953996,I80131,I80143);
nor I_55959 (I953634,I953849,I953996);
or I_55960 (I954027,I80131,I80143);
nor I_55961 (I954044,I80137,I80128);
DFFARX1 I_55962 (I954044,I2683,I953654,I954070,);
not I_55963 (I954078,I954070);
nor I_55964 (I953640,I954078,I953883);
nand I_55965 (I954109,I954078,I953728);
not I_55966 (I954126,I80137);
nand I_55967 (I954143,I954126,I953832);
nand I_55968 (I954160,I954078,I954143);
nand I_55969 (I953631,I954160,I954109);
nand I_55970 (I953628,I954143,I954027);
not I_55971 (I954232,I2690);
DFFARX1 I_55972 (I299149,I2683,I954232,I954258,);
and I_55973 (I954266,I954258,I299134);
DFFARX1 I_55974 (I954266,I2683,I954232,I954215,);
DFFARX1 I_55975 (I299140,I2683,I954232,I954306,);
not I_55976 (I954314,I299122);
not I_55977 (I954331,I299143);
nand I_55978 (I954348,I954331,I954314);
nor I_55979 (I954203,I954306,I954348);
DFFARX1 I_55980 (I954348,I2683,I954232,I954388,);
not I_55981 (I954224,I954388);
not I_55982 (I954410,I299146);
nand I_55983 (I954427,I954331,I954410);
DFFARX1 I_55984 (I954427,I2683,I954232,I954453,);
not I_55985 (I954461,I954453);
not I_55986 (I954478,I299137);
nand I_55987 (I954495,I954478,I299125);
and I_55988 (I954512,I954314,I954495);
nor I_55989 (I954529,I954427,I954512);
DFFARX1 I_55990 (I954529,I2683,I954232,I954200,);
DFFARX1 I_55991 (I954512,I2683,I954232,I954221,);
nor I_55992 (I954574,I299137,I299131);
nor I_55993 (I954212,I954427,I954574);
or I_55994 (I954605,I299137,I299131);
nor I_55995 (I954622,I299128,I299122);
DFFARX1 I_55996 (I954622,I2683,I954232,I954648,);
not I_55997 (I954656,I954648);
nor I_55998 (I954218,I954656,I954461);
nand I_55999 (I954687,I954656,I954306);
not I_56000 (I954704,I299128);
nand I_56001 (I954721,I954704,I954410);
nand I_56002 (I954738,I954656,I954721);
nand I_56003 (I954209,I954738,I954687);
nand I_56004 (I954206,I954721,I954605);
not I_56005 (I954810,I2690);
DFFARX1 I_56006 (I122985,I2683,I954810,I954836,);
and I_56007 (I954844,I954836,I122988);
DFFARX1 I_56008 (I954844,I2683,I954810,I954793,);
DFFARX1 I_56009 (I122988,I2683,I954810,I954884,);
not I_56010 (I954892,I123003);
not I_56011 (I954909,I123009);
nand I_56012 (I954926,I954909,I954892);
nor I_56013 (I954781,I954884,I954926);
DFFARX1 I_56014 (I954926,I2683,I954810,I954966,);
not I_56015 (I954802,I954966);
not I_56016 (I954988,I122997);
nand I_56017 (I955005,I954909,I954988);
DFFARX1 I_56018 (I955005,I2683,I954810,I955031,);
not I_56019 (I955039,I955031);
not I_56020 (I955056,I122994);
nand I_56021 (I955073,I955056,I122991);
and I_56022 (I955090,I954892,I955073);
nor I_56023 (I955107,I955005,I955090);
DFFARX1 I_56024 (I955107,I2683,I954810,I954778,);
DFFARX1 I_56025 (I955090,I2683,I954810,I954799,);
nor I_56026 (I955152,I122994,I122985);
nor I_56027 (I954790,I955005,I955152);
or I_56028 (I955183,I122994,I122985);
nor I_56029 (I955200,I123000,I123006);
DFFARX1 I_56030 (I955200,I2683,I954810,I955226,);
not I_56031 (I955234,I955226);
nor I_56032 (I954796,I955234,I955039);
nand I_56033 (I955265,I955234,I954884);
not I_56034 (I955282,I123000);
nand I_56035 (I955299,I955282,I954988);
nand I_56036 (I955316,I955234,I955299);
nand I_56037 (I954787,I955316,I955265);
nand I_56038 (I954784,I955299,I955183);
not I_56039 (I955388,I2690);
DFFARX1 I_56040 (I804076,I2683,I955388,I955414,);
and I_56041 (I955422,I955414,I804073);
DFFARX1 I_56042 (I955422,I2683,I955388,I955371,);
DFFARX1 I_56043 (I804079,I2683,I955388,I955462,);
not I_56044 (I955470,I804082);
not I_56045 (I955487,I804076);
nand I_56046 (I955504,I955487,I955470);
nor I_56047 (I955359,I955462,I955504);
DFFARX1 I_56048 (I955504,I2683,I955388,I955544,);
not I_56049 (I955380,I955544);
not I_56050 (I955566,I804091);
nand I_56051 (I955583,I955487,I955566);
DFFARX1 I_56052 (I955583,I2683,I955388,I955609,);
not I_56053 (I955617,I955609);
not I_56054 (I955634,I804088);
nand I_56055 (I955651,I955634,I804094);
and I_56056 (I955668,I955470,I955651);
nor I_56057 (I955685,I955583,I955668);
DFFARX1 I_56058 (I955685,I2683,I955388,I955356,);
DFFARX1 I_56059 (I955668,I2683,I955388,I955377,);
nor I_56060 (I955730,I804088,I804073);
nor I_56061 (I955368,I955583,I955730);
or I_56062 (I955761,I804088,I804073);
nor I_56063 (I955778,I804085,I804079);
DFFARX1 I_56064 (I955778,I2683,I955388,I955804,);
not I_56065 (I955812,I955804);
nor I_56066 (I955374,I955812,I955617);
nand I_56067 (I955843,I955812,I955462);
not I_56068 (I955860,I804085);
nand I_56069 (I955877,I955860,I955566);
nand I_56070 (I955894,I955812,I955877);
nand I_56071 (I955365,I955894,I955843);
nand I_56072 (I955362,I955877,I955761);
not I_56073 (I955966,I2690);
DFFARX1 I_56074 (I381290,I2683,I955966,I955992,);
nand I_56075 (I956000,I955992,I381287);
DFFARX1 I_56076 (I381266,I2683,I955966,I956026,);
DFFARX1 I_56077 (I956026,I2683,I955966,I956043,);
not I_56078 (I955958,I956043);
not I_56079 (I956065,I381281);
nor I_56080 (I956082,I381281,I381284);
not I_56081 (I956099,I381275);
nand I_56082 (I956116,I956065,I956099);
nor I_56083 (I956133,I381275,I381281);
and I_56084 (I955937,I956133,I956000);
not I_56085 (I956164,I381272);
nand I_56086 (I956181,I956164,I381293);
nor I_56087 (I956198,I381272,I381269);
not I_56088 (I956215,I956198);
nand I_56089 (I955940,I956082,I956215);
DFFARX1 I_56090 (I956198,I2683,I955966,I955955,);
nor I_56091 (I956260,I381278,I381275);
nor I_56092 (I956277,I956260,I381284);
and I_56093 (I956294,I956277,I956181);
DFFARX1 I_56094 (I956294,I2683,I955966,I955952,);
nor I_56095 (I955949,I956260,I956116);
or I_56096 (I955946,I956198,I956260);
nor I_56097 (I956353,I381278,I381266);
DFFARX1 I_56098 (I956353,I2683,I955966,I956379,);
not I_56099 (I956387,I956379);
nand I_56100 (I956404,I956387,I956065);
nor I_56101 (I956421,I956404,I381284);
DFFARX1 I_56102 (I956421,I2683,I955966,I955934,);
nor I_56103 (I956452,I956387,I956116);
nor I_56104 (I955943,I956260,I956452);
not I_56105 (I956510,I2690);
DFFARX1 I_56106 (I697098,I2683,I956510,I956536,);
nand I_56107 (I956544,I956536,I697092);
DFFARX1 I_56108 (I697095,I2683,I956510,I956570,);
DFFARX1 I_56109 (I956570,I2683,I956510,I956587,);
not I_56110 (I956502,I956587);
not I_56111 (I956609,I697101);
nor I_56112 (I956626,I697101,I697095);
not I_56113 (I956643,I697104);
nand I_56114 (I956660,I956609,I956643);
nor I_56115 (I956677,I697104,I697101);
and I_56116 (I956481,I956677,I956544);
not I_56117 (I956708,I697113);
nand I_56118 (I956725,I956708,I697107);
nor I_56119 (I956742,I697113,I697110);
not I_56120 (I956759,I956742);
nand I_56121 (I956484,I956626,I956759);
DFFARX1 I_56122 (I956742,I2683,I956510,I956499,);
nor I_56123 (I956804,I697092,I697104);
nor I_56124 (I956821,I956804,I697095);
and I_56125 (I956838,I956821,I956725);
DFFARX1 I_56126 (I956838,I2683,I956510,I956496,);
nor I_56127 (I956493,I956804,I956660);
or I_56128 (I956490,I956742,I956804);
nor I_56129 (I956897,I697092,I697098);
DFFARX1 I_56130 (I956897,I2683,I956510,I956923,);
not I_56131 (I956931,I956923);
nand I_56132 (I956948,I956931,I956609);
nor I_56133 (I956965,I956948,I697095);
DFFARX1 I_56134 (I956965,I2683,I956510,I956478,);
nor I_56135 (I956996,I956931,I956660);
nor I_56136 (I956487,I956804,I956996);
not I_56137 (I957054,I2690);
DFFARX1 I_56138 (I1092981,I2683,I957054,I957080,);
nand I_56139 (I957088,I957080,I1092966);
DFFARX1 I_56140 (I1092960,I2683,I957054,I957114,);
DFFARX1 I_56141 (I957114,I2683,I957054,I957131,);
not I_56142 (I957046,I957131);
not I_56143 (I957153,I1092954);
nor I_56144 (I957170,I1092954,I1092975);
not I_56145 (I957187,I1092963);
nand I_56146 (I957204,I957153,I957187);
nor I_56147 (I957221,I1092963,I1092954);
and I_56148 (I957025,I957221,I957088);
not I_56149 (I957252,I1092972);
nand I_56150 (I957269,I957252,I1092978);
nor I_56151 (I957286,I1092972,I1092969);
not I_56152 (I957303,I957286);
nand I_56153 (I957028,I957170,I957303);
DFFARX1 I_56154 (I957286,I2683,I957054,I957043,);
nor I_56155 (I957348,I1092957,I1092963);
nor I_56156 (I957365,I957348,I1092975);
and I_56157 (I957382,I957365,I957269);
DFFARX1 I_56158 (I957382,I2683,I957054,I957040,);
nor I_56159 (I957037,I957348,I957204);
or I_56160 (I957034,I957286,I957348);
nor I_56161 (I957441,I1092957,I1092954);
DFFARX1 I_56162 (I957441,I2683,I957054,I957467,);
not I_56163 (I957475,I957467);
nand I_56164 (I957492,I957475,I957153);
nor I_56165 (I957509,I957492,I1092975);
DFFARX1 I_56166 (I957509,I2683,I957054,I957022,);
nor I_56167 (I957540,I957475,I957204);
nor I_56168 (I957031,I957348,I957540);
not I_56169 (I957598,I2690);
DFFARX1 I_56170 (I1024335,I2683,I957598,I957624,);
nand I_56171 (I957632,I957624,I1024320);
DFFARX1 I_56172 (I1024332,I2683,I957598,I957658,);
DFFARX1 I_56173 (I957658,I2683,I957598,I957675,);
not I_56174 (I957590,I957675);
not I_56175 (I957697,I1024326);
nor I_56176 (I957714,I1024326,I1024317);
not I_56177 (I957731,I1024311);
nand I_56178 (I957748,I957697,I957731);
nor I_56179 (I957765,I1024311,I1024326);
and I_56180 (I957569,I957765,I957632);
not I_56181 (I957796,I1024323);
nand I_56182 (I957813,I957796,I1024308);
nor I_56183 (I957830,I1024323,I1024329);
not I_56184 (I957847,I957830);
nand I_56185 (I957572,I957714,I957847);
DFFARX1 I_56186 (I957830,I2683,I957598,I957587,);
nor I_56187 (I957892,I1024314,I1024311);
nor I_56188 (I957909,I957892,I1024317);
and I_56189 (I957926,I957909,I957813);
DFFARX1 I_56190 (I957926,I2683,I957598,I957584,);
nor I_56191 (I957581,I957892,I957748);
or I_56192 (I957578,I957830,I957892);
nor I_56193 (I957985,I1024314,I1024308);
DFFARX1 I_56194 (I957985,I2683,I957598,I958011,);
not I_56195 (I958019,I958011);
nand I_56196 (I958036,I958019,I957697);
nor I_56197 (I958053,I958036,I1024317);
DFFARX1 I_56198 (I958053,I2683,I957598,I957566,);
nor I_56199 (I958084,I958019,I957748);
nor I_56200 (I957575,I957892,I958084);
not I_56201 (I958142,I2690);
DFFARX1 I_56202 (I124184,I2683,I958142,I958168,);
nand I_56203 (I958176,I958168,I124199);
DFFARX1 I_56204 (I124196,I2683,I958142,I958202,);
DFFARX1 I_56205 (I958202,I2683,I958142,I958219,);
not I_56206 (I958134,I958219);
not I_56207 (I958241,I124175);
nor I_56208 (I958258,I124175,I124181);
not I_56209 (I958275,I124187);
nand I_56210 (I958292,I958241,I958275);
nor I_56211 (I958309,I124187,I124175);
and I_56212 (I958113,I958309,I958176);
not I_56213 (I958340,I124193);
nand I_56214 (I958357,I958340,I124175);
nor I_56215 (I958374,I124193,I124178);
not I_56216 (I958391,I958374);
nand I_56217 (I958116,I958258,I958391);
DFFARX1 I_56218 (I958374,I2683,I958142,I958131,);
nor I_56219 (I958436,I124178,I124187);
nor I_56220 (I958453,I958436,I124181);
and I_56221 (I958470,I958453,I958357);
DFFARX1 I_56222 (I958470,I2683,I958142,I958128,);
nor I_56223 (I958125,I958436,I958292);
or I_56224 (I958122,I958374,I958436);
nor I_56225 (I958529,I124178,I124190);
DFFARX1 I_56226 (I958529,I2683,I958142,I958555,);
not I_56227 (I958563,I958555);
nand I_56228 (I958580,I958563,I958241);
nor I_56229 (I958597,I958580,I124181);
DFFARX1 I_56230 (I958597,I2683,I958142,I958110,);
nor I_56231 (I958628,I958563,I958292);
nor I_56232 (I958119,I958436,I958628);
not I_56233 (I958686,I2690);
DFFARX1 I_56234 (I563033,I2683,I958686,I958712,);
nand I_56235 (I958720,I958712,I563048);
DFFARX1 I_56236 (I563042,I2683,I958686,I958746,);
DFFARX1 I_56237 (I958746,I2683,I958686,I958763,);
not I_56238 (I958678,I958763);
not I_56239 (I958785,I563045);
nor I_56240 (I958802,I563045,I563051);
not I_56241 (I958819,I563033);
nand I_56242 (I958836,I958785,I958819);
nor I_56243 (I958853,I563033,I563045);
and I_56244 (I958657,I958853,I958720);
not I_56245 (I958884,I563030);
nand I_56246 (I958901,I958884,I563036);
nor I_56247 (I958918,I563030,I563030);
not I_56248 (I958935,I958918);
nand I_56249 (I958660,I958802,I958935);
DFFARX1 I_56250 (I958918,I2683,I958686,I958675,);
nor I_56251 (I958980,I563039,I563033);
nor I_56252 (I958997,I958980,I563051);
and I_56253 (I959014,I958997,I958901);
DFFARX1 I_56254 (I959014,I2683,I958686,I958672,);
nor I_56255 (I958669,I958980,I958836);
or I_56256 (I958666,I958918,I958980);
nor I_56257 (I959073,I563039,I563054);
DFFARX1 I_56258 (I959073,I2683,I958686,I959099,);
not I_56259 (I959107,I959099);
nand I_56260 (I959124,I959107,I958785);
nor I_56261 (I959141,I959124,I563051);
DFFARX1 I_56262 (I959141,I2683,I958686,I958654,);
nor I_56263 (I959172,I959107,I958836);
nor I_56264 (I958663,I958980,I959172);
not I_56265 (I959230,I2690);
DFFARX1 I_56266 (I743247,I2683,I959230,I959256,);
nand I_56267 (I959264,I959256,I743247);
DFFARX1 I_56268 (I743259,I2683,I959230,I959290,);
DFFARX1 I_56269 (I959290,I2683,I959230,I959307,);
not I_56270 (I959222,I959307);
not I_56271 (I959329,I743253);
nor I_56272 (I959346,I743253,I743274);
not I_56273 (I959363,I743262);
nand I_56274 (I959380,I959329,I959363);
nor I_56275 (I959397,I743262,I743253);
and I_56276 (I959201,I959397,I959264);
not I_56277 (I959428,I743256);
nand I_56278 (I959445,I959428,I743271);
nor I_56279 (I959462,I743256,I743265);
not I_56280 (I959479,I959462);
nand I_56281 (I959204,I959346,I959479);
DFFARX1 I_56282 (I959462,I2683,I959230,I959219,);
nor I_56283 (I959524,I743268,I743262);
nor I_56284 (I959541,I959524,I743274);
and I_56285 (I959558,I959541,I959445);
DFFARX1 I_56286 (I959558,I2683,I959230,I959216,);
nor I_56287 (I959213,I959524,I959380);
or I_56288 (I959210,I959462,I959524);
nor I_56289 (I959617,I743268,I743250);
DFFARX1 I_56290 (I959617,I2683,I959230,I959643,);
not I_56291 (I959651,I959643);
nand I_56292 (I959668,I959651,I959329);
nor I_56293 (I959685,I959668,I743274);
DFFARX1 I_56294 (I959685,I2683,I959230,I959198,);
nor I_56295 (I959716,I959651,I959380);
nor I_56296 (I959207,I959524,I959716);
not I_56297 (I959774,I2690);
DFFARX1 I_56298 (I781361,I2683,I959774,I959800,);
nand I_56299 (I959808,I959800,I781361);
DFFARX1 I_56300 (I781373,I2683,I959774,I959834,);
DFFARX1 I_56301 (I959834,I2683,I959774,I959851,);
not I_56302 (I959766,I959851);
not I_56303 (I959873,I781367);
nor I_56304 (I959890,I781367,I781388);
not I_56305 (I959907,I781376);
nand I_56306 (I959924,I959873,I959907);
nor I_56307 (I959941,I781376,I781367);
and I_56308 (I959745,I959941,I959808);
not I_56309 (I959972,I781370);
nand I_56310 (I959989,I959972,I781385);
nor I_56311 (I960006,I781370,I781379);
not I_56312 (I960023,I960006);
nand I_56313 (I959748,I959890,I960023);
DFFARX1 I_56314 (I960006,I2683,I959774,I959763,);
nor I_56315 (I960068,I781382,I781376);
nor I_56316 (I960085,I960068,I781388);
and I_56317 (I960102,I960085,I959989);
DFFARX1 I_56318 (I960102,I2683,I959774,I959760,);
nor I_56319 (I959757,I960068,I959924);
or I_56320 (I959754,I960006,I960068);
nor I_56321 (I960161,I781382,I781364);
DFFARX1 I_56322 (I960161,I2683,I959774,I960187,);
not I_56323 (I960195,I960187);
nand I_56324 (I960212,I960195,I959873);
nor I_56325 (I960229,I960212,I781388);
DFFARX1 I_56326 (I960229,I2683,I959774,I959742,);
nor I_56327 (I960260,I960195,I959924);
nor I_56328 (I959751,I960068,I960260);
not I_56329 (I960318,I2690);
DFFARX1 I_56330 (I291229,I2683,I960318,I960344,);
nand I_56331 (I960352,I960344,I291232);
DFFARX1 I_56332 (I291226,I2683,I960318,I960378,);
DFFARX1 I_56333 (I960378,I2683,I960318,I960395,);
not I_56334 (I960310,I960395);
not I_56335 (I960417,I291235);
nor I_56336 (I960434,I291235,I291220);
not I_56337 (I960451,I291244);
nand I_56338 (I960468,I960417,I960451);
nor I_56339 (I960485,I291244,I291235);
and I_56340 (I960289,I960485,I960352);
not I_56341 (I960516,I291223);
nand I_56342 (I960533,I960516,I291241);
nor I_56343 (I960550,I291223,I291217);
not I_56344 (I960567,I960550);
nand I_56345 (I960292,I960434,I960567);
DFFARX1 I_56346 (I960550,I2683,I960318,I960307,);
nor I_56347 (I960612,I291238,I291244);
nor I_56348 (I960629,I960612,I291220);
and I_56349 (I960646,I960629,I960533);
DFFARX1 I_56350 (I960646,I2683,I960318,I960304,);
nor I_56351 (I960301,I960612,I960468);
or I_56352 (I960298,I960550,I960612);
nor I_56353 (I960705,I291238,I291217);
DFFARX1 I_56354 (I960705,I2683,I960318,I960731,);
not I_56355 (I960739,I960731);
nand I_56356 (I960756,I960739,I960417);
nor I_56357 (I960773,I960756,I291220);
DFFARX1 I_56358 (I960773,I2683,I960318,I960286,);
nor I_56359 (I960804,I960739,I960468);
nor I_56360 (I960295,I960612,I960804);
not I_56361 (I960862,I2690);
DFFARX1 I_56362 (I1059661,I2683,I960862,I960888,);
nand I_56363 (I960896,I960888,I1059646);
DFFARX1 I_56364 (I1059640,I2683,I960862,I960922,);
DFFARX1 I_56365 (I960922,I2683,I960862,I960939,);
not I_56366 (I960854,I960939);
not I_56367 (I960961,I1059634);
nor I_56368 (I960978,I1059634,I1059655);
not I_56369 (I960995,I1059643);
nand I_56370 (I961012,I960961,I960995);
nor I_56371 (I961029,I1059643,I1059634);
and I_56372 (I960833,I961029,I960896);
not I_56373 (I961060,I1059652);
nand I_56374 (I961077,I961060,I1059658);
nor I_56375 (I961094,I1059652,I1059649);
not I_56376 (I961111,I961094);
nand I_56377 (I960836,I960978,I961111);
DFFARX1 I_56378 (I961094,I2683,I960862,I960851,);
nor I_56379 (I961156,I1059637,I1059643);
nor I_56380 (I961173,I961156,I1059655);
and I_56381 (I961190,I961173,I961077);
DFFARX1 I_56382 (I961190,I2683,I960862,I960848,);
nor I_56383 (I960845,I961156,I961012);
or I_56384 (I960842,I961094,I961156);
nor I_56385 (I961249,I1059637,I1059634);
DFFARX1 I_56386 (I961249,I2683,I960862,I961275,);
not I_56387 (I961283,I961275);
nand I_56388 (I961300,I961283,I960961);
nor I_56389 (I961317,I961300,I1059655);
DFFARX1 I_56390 (I961317,I2683,I960862,I960830,);
nor I_56391 (I961348,I961283,I961012);
nor I_56392 (I960839,I961156,I961348);
not I_56393 (I961406,I2690);
DFFARX1 I_56394 (I801286,I2683,I961406,I961432,);
nand I_56395 (I961440,I961432,I801274);
DFFARX1 I_56396 (I801268,I2683,I961406,I961466,);
DFFARX1 I_56397 (I961466,I2683,I961406,I961483,);
not I_56398 (I961398,I961483);
not I_56399 (I961505,I801268);
nor I_56400 (I961522,I801268,I801280);
not I_56401 (I961539,I801277);
nand I_56402 (I961556,I961505,I961539);
nor I_56403 (I961573,I801277,I801268);
and I_56404 (I961377,I961573,I961440);
not I_56405 (I961604,I801271);
nand I_56406 (I961621,I961604,I801283);
nor I_56407 (I961638,I801271,I801289);
not I_56408 (I961655,I961638);
nand I_56409 (I961380,I961522,I961655);
DFFARX1 I_56410 (I961638,I2683,I961406,I961395,);
nor I_56411 (I961700,I801274,I801277);
nor I_56412 (I961717,I961700,I801280);
and I_56413 (I961734,I961717,I961621);
DFFARX1 I_56414 (I961734,I2683,I961406,I961392,);
nor I_56415 (I961389,I961700,I961556);
or I_56416 (I961386,I961638,I961700);
nor I_56417 (I961793,I801274,I801271);
DFFARX1 I_56418 (I961793,I2683,I961406,I961819,);
not I_56419 (I961827,I961819);
nand I_56420 (I961844,I961827,I961505);
nor I_56421 (I961861,I961844,I801280);
DFFARX1 I_56422 (I961861,I2683,I961406,I961374,);
nor I_56423 (I961892,I961827,I961556);
nor I_56424 (I961383,I961700,I961892);
not I_56425 (I961950,I2690);
DFFARX1 I_56426 (I721929,I2683,I961950,I961976,);
nand I_56427 (I961984,I961976,I721929);
DFFARX1 I_56428 (I721941,I2683,I961950,I962010,);
DFFARX1 I_56429 (I962010,I2683,I961950,I962027,);
not I_56430 (I961942,I962027);
not I_56431 (I962049,I721935);
nor I_56432 (I962066,I721935,I721956);
not I_56433 (I962083,I721944);
nand I_56434 (I962100,I962049,I962083);
nor I_56435 (I962117,I721944,I721935);
and I_56436 (I961921,I962117,I961984);
not I_56437 (I962148,I721938);
nand I_56438 (I962165,I962148,I721953);
nor I_56439 (I962182,I721938,I721947);
not I_56440 (I962199,I962182);
nand I_56441 (I961924,I962066,I962199);
DFFARX1 I_56442 (I962182,I2683,I961950,I961939,);
nor I_56443 (I962244,I721950,I721944);
nor I_56444 (I962261,I962244,I721956);
and I_56445 (I962278,I962261,I962165);
DFFARX1 I_56446 (I962278,I2683,I961950,I961936,);
nor I_56447 (I961933,I962244,I962100);
or I_56448 (I961930,I962182,I962244);
nor I_56449 (I962337,I721950,I721932);
DFFARX1 I_56450 (I962337,I2683,I961950,I962363,);
not I_56451 (I962371,I962363);
nand I_56452 (I962388,I962371,I962049);
nor I_56453 (I962405,I962388,I721956);
DFFARX1 I_56454 (I962405,I2683,I961950,I961918,);
nor I_56455 (I962436,I962371,I962100);
nor I_56456 (I961927,I962244,I962436);
not I_56457 (I962494,I2690);
DFFARX1 I_56458 (I22694,I2683,I962494,I962520,);
nand I_56459 (I962528,I962520,I22688);
DFFARX1 I_56460 (I22709,I2683,I962494,I962554,);
DFFARX1 I_56461 (I962554,I2683,I962494,I962571,);
not I_56462 (I962486,I962571);
not I_56463 (I962593,I22697);
nor I_56464 (I962610,I22697,I22706);
not I_56465 (I962627,I22685);
nand I_56466 (I962644,I962593,I962627);
nor I_56467 (I962661,I22685,I22697);
and I_56468 (I962465,I962661,I962528);
not I_56469 (I962692,I22703);
nand I_56470 (I962709,I962692,I22691);
nor I_56471 (I962726,I22703,I22685);
not I_56472 (I962743,I962726);
nand I_56473 (I962468,I962610,I962743);
DFFARX1 I_56474 (I962726,I2683,I962494,I962483,);
nor I_56475 (I962788,I22688,I22685);
nor I_56476 (I962805,I962788,I22706);
and I_56477 (I962822,I962805,I962709);
DFFARX1 I_56478 (I962822,I2683,I962494,I962480,);
nor I_56479 (I962477,I962788,I962644);
or I_56480 (I962474,I962726,I962788);
nor I_56481 (I962881,I22688,I22700);
DFFARX1 I_56482 (I962881,I2683,I962494,I962907,);
not I_56483 (I962915,I962907);
nand I_56484 (I962932,I962915,I962593);
nor I_56485 (I962949,I962932,I22706);
DFFARX1 I_56486 (I962949,I2683,I962494,I962462,);
nor I_56487 (I962980,I962915,I962644);
nor I_56488 (I962471,I962788,I962980);
not I_56489 (I963038,I2690);
DFFARX1 I_56490 (I1053116,I2683,I963038,I963064,);
nand I_56491 (I963072,I963064,I1053101);
DFFARX1 I_56492 (I1053095,I2683,I963038,I963098,);
DFFARX1 I_56493 (I963098,I2683,I963038,I963115,);
not I_56494 (I963030,I963115);
not I_56495 (I963137,I1053089);
nor I_56496 (I963154,I1053089,I1053110);
not I_56497 (I963171,I1053098);
nand I_56498 (I963188,I963137,I963171);
nor I_56499 (I963205,I1053098,I1053089);
and I_56500 (I963009,I963205,I963072);
not I_56501 (I963236,I1053107);
nand I_56502 (I963253,I963236,I1053113);
nor I_56503 (I963270,I1053107,I1053104);
not I_56504 (I963287,I963270);
nand I_56505 (I963012,I963154,I963287);
DFFARX1 I_56506 (I963270,I2683,I963038,I963027,);
nor I_56507 (I963332,I1053092,I1053098);
nor I_56508 (I963349,I963332,I1053110);
and I_56509 (I963366,I963349,I963253);
DFFARX1 I_56510 (I963366,I2683,I963038,I963024,);
nor I_56511 (I963021,I963332,I963188);
or I_56512 (I963018,I963270,I963332);
nor I_56513 (I963425,I1053092,I1053089);
DFFARX1 I_56514 (I963425,I2683,I963038,I963451,);
not I_56515 (I963459,I963451);
nand I_56516 (I963476,I963459,I963137);
nor I_56517 (I963493,I963476,I1053110);
DFFARX1 I_56518 (I963493,I2683,I963038,I963006,);
nor I_56519 (I963524,I963459,I963188);
nor I_56520 (I963015,I963332,I963524);
not I_56521 (I963582,I2690);
DFFARX1 I_56522 (I902204,I2683,I963582,I963608,);
nand I_56523 (I963616,I963608,I902183);
DFFARX1 I_56524 (I902180,I2683,I963582,I963642,);
DFFARX1 I_56525 (I963642,I2683,I963582,I963659,);
not I_56526 (I963574,I963659);
not I_56527 (I963681,I902192);
nor I_56528 (I963698,I902192,I902201);
not I_56529 (I963715,I902189);
nand I_56530 (I963732,I963681,I963715);
nor I_56531 (I963749,I902189,I902192);
and I_56532 (I963553,I963749,I963616);
not I_56533 (I963780,I902198);
nand I_56534 (I963797,I963780,I902195);
nor I_56535 (I963814,I902198,I902180);
not I_56536 (I963831,I963814);
nand I_56537 (I963556,I963698,I963831);
DFFARX1 I_56538 (I963814,I2683,I963582,I963571,);
nor I_56539 (I963876,I902183,I902189);
nor I_56540 (I963893,I963876,I902201);
and I_56541 (I963910,I963893,I963797);
DFFARX1 I_56542 (I963910,I2683,I963582,I963568,);
nor I_56543 (I963565,I963876,I963732);
or I_56544 (I963562,I963814,I963876);
nor I_56545 (I963969,I902183,I902186);
DFFARX1 I_56546 (I963969,I2683,I963582,I963995,);
not I_56547 (I964003,I963995);
nand I_56548 (I964020,I964003,I963681);
nor I_56549 (I964037,I964020,I902201);
DFFARX1 I_56550 (I964037,I2683,I963582,I963550,);
nor I_56551 (I964068,I964003,I963732);
nor I_56552 (I963559,I963876,I964068);
not I_56553 (I964126,I2690);
DFFARX1 I_56554 (I424667,I2683,I964126,I964152,);
nand I_56555 (I964160,I964152,I424691);
DFFARX1 I_56556 (I424670,I2683,I964126,I964186,);
DFFARX1 I_56557 (I964186,I2683,I964126,I964203,);
not I_56558 (I964118,I964203);
not I_56559 (I964225,I424673);
nor I_56560 (I964242,I424673,I424688);
not I_56561 (I964259,I424679);
nand I_56562 (I964276,I964225,I964259);
nor I_56563 (I964293,I424679,I424673);
and I_56564 (I964097,I964293,I964160);
not I_56565 (I964324,I424676);
nand I_56566 (I964341,I964324,I424670);
nor I_56567 (I964358,I424676,I424685);
not I_56568 (I964375,I964358);
nand I_56569 (I964100,I964242,I964375);
DFFARX1 I_56570 (I964358,I2683,I964126,I964115,);
nor I_56571 (I964420,I424682,I424679);
nor I_56572 (I964437,I964420,I424688);
and I_56573 (I964454,I964437,I964341);
DFFARX1 I_56574 (I964454,I2683,I964126,I964112,);
nor I_56575 (I964109,I964420,I964276);
or I_56576 (I964106,I964358,I964420);
nor I_56577 (I964513,I424682,I424667);
DFFARX1 I_56578 (I964513,I2683,I964126,I964539,);
not I_56579 (I964547,I964539);
nand I_56580 (I964564,I964547,I964225);
nor I_56581 (I964581,I964564,I424688);
DFFARX1 I_56582 (I964581,I2683,I964126,I964094,);
nor I_56583 (I964612,I964547,I964276);
nor I_56584 (I964103,I964420,I964612);
not I_56585 (I964670,I2690);
DFFARX1 I_56586 (I569391,I2683,I964670,I964696,);
nand I_56587 (I964704,I964696,I569406);
DFFARX1 I_56588 (I569400,I2683,I964670,I964730,);
DFFARX1 I_56589 (I964730,I2683,I964670,I964747,);
not I_56590 (I964662,I964747);
not I_56591 (I964769,I569403);
nor I_56592 (I964786,I569403,I569409);
not I_56593 (I964803,I569391);
nand I_56594 (I964820,I964769,I964803);
nor I_56595 (I964837,I569391,I569403);
and I_56596 (I964641,I964837,I964704);
not I_56597 (I964868,I569388);
nand I_56598 (I964885,I964868,I569394);
nor I_56599 (I964902,I569388,I569388);
not I_56600 (I964919,I964902);
nand I_56601 (I964644,I964786,I964919);
DFFARX1 I_56602 (I964902,I2683,I964670,I964659,);
nor I_56603 (I964964,I569397,I569391);
nor I_56604 (I964981,I964964,I569409);
and I_56605 (I964998,I964981,I964885);
DFFARX1 I_56606 (I964998,I2683,I964670,I964656,);
nor I_56607 (I964653,I964964,I964820);
or I_56608 (I964650,I964902,I964964);
nor I_56609 (I965057,I569397,I569412);
DFFARX1 I_56610 (I965057,I2683,I964670,I965083,);
not I_56611 (I965091,I965083);
nand I_56612 (I965108,I965091,I964769);
nor I_56613 (I965125,I965108,I569409);
DFFARX1 I_56614 (I965125,I2683,I964670,I964638,);
nor I_56615 (I965156,I965091,I964820);
nor I_56616 (I964647,I964964,I965156);
not I_56617 (I965214,I2690);
DFFARX1 I_56618 (I318186,I2683,I965214,I965240,);
nand I_56619 (I965248,I965240,I318183);
DFFARX1 I_56620 (I318162,I2683,I965214,I965274,);
DFFARX1 I_56621 (I965274,I2683,I965214,I965291,);
not I_56622 (I965206,I965291);
not I_56623 (I965313,I318177);
nor I_56624 (I965330,I318177,I318180);
not I_56625 (I965347,I318171);
nand I_56626 (I965364,I965313,I965347);
nor I_56627 (I965381,I318171,I318177);
and I_56628 (I965185,I965381,I965248);
not I_56629 (I965412,I318168);
nand I_56630 (I965429,I965412,I318189);
nor I_56631 (I965446,I318168,I318165);
not I_56632 (I965463,I965446);
nand I_56633 (I965188,I965330,I965463);
DFFARX1 I_56634 (I965446,I2683,I965214,I965203,);
nor I_56635 (I965508,I318174,I318171);
nor I_56636 (I965525,I965508,I318180);
and I_56637 (I965542,I965525,I965429);
DFFARX1 I_56638 (I965542,I2683,I965214,I965200,);
nor I_56639 (I965197,I965508,I965364);
or I_56640 (I965194,I965446,I965508);
nor I_56641 (I965601,I318174,I318162);
DFFARX1 I_56642 (I965601,I2683,I965214,I965627,);
not I_56643 (I965635,I965627);
nand I_56644 (I965652,I965635,I965313);
nor I_56645 (I965669,I965652,I318180);
DFFARX1 I_56646 (I965669,I2683,I965214,I965182,);
nor I_56647 (I965700,I965635,I965364);
nor I_56648 (I965191,I965508,I965700);
not I_56649 (I965758,I2690);
DFFARX1 I_56650 (I609273,I2683,I965758,I965784,);
nand I_56651 (I965792,I965784,I609288);
DFFARX1 I_56652 (I609282,I2683,I965758,I965818,);
DFFARX1 I_56653 (I965818,I2683,I965758,I965835,);
not I_56654 (I965750,I965835);
not I_56655 (I965857,I609285);
nor I_56656 (I965874,I609285,I609291);
not I_56657 (I965891,I609273);
nand I_56658 (I965908,I965857,I965891);
nor I_56659 (I965925,I609273,I609285);
and I_56660 (I965729,I965925,I965792);
not I_56661 (I965956,I609270);
nand I_56662 (I965973,I965956,I609276);
nor I_56663 (I965990,I609270,I609270);
not I_56664 (I966007,I965990);
nand I_56665 (I965732,I965874,I966007);
DFFARX1 I_56666 (I965990,I2683,I965758,I965747,);
nor I_56667 (I966052,I609279,I609273);
nor I_56668 (I966069,I966052,I609291);
and I_56669 (I966086,I966069,I965973);
DFFARX1 I_56670 (I966086,I2683,I965758,I965744,);
nor I_56671 (I965741,I966052,I965908);
or I_56672 (I965738,I965990,I966052);
nor I_56673 (I966145,I609279,I609294);
DFFARX1 I_56674 (I966145,I2683,I965758,I966171,);
not I_56675 (I966179,I966171);
nand I_56676 (I966196,I966179,I965857);
nor I_56677 (I966213,I966196,I609291);
DFFARX1 I_56678 (I966213,I2683,I965758,I965726,);
nor I_56679 (I966244,I966179,I965908);
nor I_56680 (I965735,I966052,I966244);
not I_56681 (I966302,I2690);
DFFARX1 I_56682 (I82784,I2683,I966302,I966328,);
nand I_56683 (I966336,I966328,I82766);
DFFARX1 I_56684 (I82763,I2683,I966302,I966362,);
DFFARX1 I_56685 (I966362,I2683,I966302,I966379,);
not I_56686 (I966294,I966379);
not I_56687 (I966401,I82781);
nor I_56688 (I966418,I82781,I82775);
not I_56689 (I966435,I82763);
nand I_56690 (I966452,I966401,I966435);
nor I_56691 (I966469,I82763,I82781);
and I_56692 (I966273,I966469,I966336);
not I_56693 (I966500,I82772);
nand I_56694 (I966517,I966500,I82778);
nor I_56695 (I966534,I82772,I82766);
not I_56696 (I966551,I966534);
nand I_56697 (I966276,I966418,I966551);
DFFARX1 I_56698 (I966534,I2683,I966302,I966291,);
nor I_56699 (I966596,I82769,I82763);
nor I_56700 (I966613,I966596,I82775);
and I_56701 (I966630,I966613,I966517);
DFFARX1 I_56702 (I966630,I2683,I966302,I966288,);
nor I_56703 (I966285,I966596,I966452);
or I_56704 (I966282,I966534,I966596);
nor I_56705 (I966689,I82769,I82787);
DFFARX1 I_56706 (I966689,I2683,I966302,I966715,);
not I_56707 (I966723,I966715);
nand I_56708 (I966740,I966723,I966401);
nor I_56709 (I966757,I966740,I82775);
DFFARX1 I_56710 (I966757,I2683,I966302,I966270,);
nor I_56711 (I966788,I966723,I966452);
nor I_56712 (I966279,I966596,I966788);
not I_56713 (I966846,I2690);
DFFARX1 I_56714 (I740017,I2683,I966846,I966872,);
nand I_56715 (I966880,I966872,I740017);
DFFARX1 I_56716 (I740029,I2683,I966846,I966906,);
DFFARX1 I_56717 (I966906,I2683,I966846,I966923,);
not I_56718 (I966838,I966923);
not I_56719 (I966945,I740023);
nor I_56720 (I966962,I740023,I740044);
not I_56721 (I966979,I740032);
nand I_56722 (I966996,I966945,I966979);
nor I_56723 (I967013,I740032,I740023);
and I_56724 (I966817,I967013,I966880);
not I_56725 (I967044,I740026);
nand I_56726 (I967061,I967044,I740041);
nor I_56727 (I967078,I740026,I740035);
not I_56728 (I967095,I967078);
nand I_56729 (I966820,I966962,I967095);
DFFARX1 I_56730 (I967078,I2683,I966846,I966835,);
nor I_56731 (I967140,I740038,I740032);
nor I_56732 (I967157,I967140,I740044);
and I_56733 (I967174,I967157,I967061);
DFFARX1 I_56734 (I967174,I2683,I966846,I966832,);
nor I_56735 (I966829,I967140,I966996);
or I_56736 (I966826,I967078,I967140);
nor I_56737 (I967233,I740038,I740020);
DFFARX1 I_56738 (I967233,I2683,I966846,I967259,);
not I_56739 (I967267,I967259);
nand I_56740 (I967284,I967267,I966945);
nor I_56741 (I967301,I967284,I740044);
DFFARX1 I_56742 (I967301,I2683,I966846,I966814,);
nor I_56743 (I967332,I967267,I966996);
nor I_56744 (I966823,I967140,I967332);
not I_56745 (I967390,I2690);
DFFARX1 I_56746 (I935150,I2683,I967390,I967416,);
nand I_56747 (I967424,I967416,I935129);
DFFARX1 I_56748 (I935126,I2683,I967390,I967450,);
DFFARX1 I_56749 (I967450,I2683,I967390,I967467,);
not I_56750 (I967382,I967467);
not I_56751 (I967489,I935138);
nor I_56752 (I967506,I935138,I935147);
not I_56753 (I967523,I935135);
nand I_56754 (I967540,I967489,I967523);
nor I_56755 (I967557,I935135,I935138);
and I_56756 (I967361,I967557,I967424);
not I_56757 (I967588,I935144);
nand I_56758 (I967605,I967588,I935141);
nor I_56759 (I967622,I935144,I935126);
not I_56760 (I967639,I967622);
nand I_56761 (I967364,I967506,I967639);
DFFARX1 I_56762 (I967622,I2683,I967390,I967379,);
nor I_56763 (I967684,I935129,I935135);
nor I_56764 (I967701,I967684,I935147);
and I_56765 (I967718,I967701,I967605);
DFFARX1 I_56766 (I967718,I2683,I967390,I967376,);
nor I_56767 (I967373,I967684,I967540);
or I_56768 (I967370,I967622,I967684);
nor I_56769 (I967777,I935129,I935132);
DFFARX1 I_56770 (I967777,I2683,I967390,I967803,);
not I_56771 (I967811,I967803);
nand I_56772 (I967828,I967811,I967489);
nor I_56773 (I967845,I967828,I935147);
DFFARX1 I_56774 (I967845,I2683,I967390,I967358,);
nor I_56775 (I967876,I967811,I967540);
nor I_56776 (I967367,I967684,I967876);
not I_56777 (I967934,I2690);
DFFARX1 I_56778 (I227462,I2683,I967934,I967960,);
nand I_56779 (I967968,I967960,I227465);
DFFARX1 I_56780 (I227459,I2683,I967934,I967994,);
DFFARX1 I_56781 (I967994,I2683,I967934,I968011,);
not I_56782 (I967926,I968011);
not I_56783 (I968033,I227468);
nor I_56784 (I968050,I227468,I227453);
not I_56785 (I968067,I227477);
nand I_56786 (I968084,I968033,I968067);
nor I_56787 (I968101,I227477,I227468);
and I_56788 (I967905,I968101,I967968);
not I_56789 (I968132,I227456);
nand I_56790 (I968149,I968132,I227474);
nor I_56791 (I968166,I227456,I227450);
not I_56792 (I968183,I968166);
nand I_56793 (I967908,I968050,I968183);
DFFARX1 I_56794 (I968166,I2683,I967934,I967923,);
nor I_56795 (I968228,I227471,I227477);
nor I_56796 (I968245,I968228,I227453);
and I_56797 (I968262,I968245,I968149);
DFFARX1 I_56798 (I968262,I2683,I967934,I967920,);
nor I_56799 (I967917,I968228,I968084);
or I_56800 (I967914,I968166,I968228);
nor I_56801 (I968321,I227471,I227450);
DFFARX1 I_56802 (I968321,I2683,I967934,I968347,);
not I_56803 (I968355,I968347);
nand I_56804 (I968372,I968355,I968033);
nor I_56805 (I968389,I968372,I227453);
DFFARX1 I_56806 (I968389,I2683,I967934,I967902,);
nor I_56807 (I968420,I968355,I968084);
nor I_56808 (I967911,I968228,I968420);
not I_56809 (I968478,I2690);
DFFARX1 I_56810 (I234840,I2683,I968478,I968504,);
nand I_56811 (I968512,I968504,I234843);
DFFARX1 I_56812 (I234837,I2683,I968478,I968538,);
DFFARX1 I_56813 (I968538,I2683,I968478,I968555,);
not I_56814 (I968470,I968555);
not I_56815 (I968577,I234846);
nor I_56816 (I968594,I234846,I234831);
not I_56817 (I968611,I234855);
nand I_56818 (I968628,I968577,I968611);
nor I_56819 (I968645,I234855,I234846);
and I_56820 (I968449,I968645,I968512);
not I_56821 (I968676,I234834);
nand I_56822 (I968693,I968676,I234852);
nor I_56823 (I968710,I234834,I234828);
not I_56824 (I968727,I968710);
nand I_56825 (I968452,I968594,I968727);
DFFARX1 I_56826 (I968710,I2683,I968478,I968467,);
nor I_56827 (I968772,I234849,I234855);
nor I_56828 (I968789,I968772,I234831);
and I_56829 (I968806,I968789,I968693);
DFFARX1 I_56830 (I968806,I2683,I968478,I968464,);
nor I_56831 (I968461,I968772,I968628);
or I_56832 (I968458,I968710,I968772);
nor I_56833 (I968865,I234849,I234828);
DFFARX1 I_56834 (I968865,I2683,I968478,I968891,);
not I_56835 (I968899,I968891);
nand I_56836 (I968916,I968899,I968577);
nor I_56837 (I968933,I968916,I234831);
DFFARX1 I_56838 (I968933,I2683,I968478,I968446,);
nor I_56839 (I968964,I968899,I968628);
nor I_56840 (I968455,I968772,I968964);
not I_56841 (I969022,I2690);
DFFARX1 I_56842 (I684977,I2683,I969022,I969048,);
nand I_56843 (I969056,I969048,I684971);
DFFARX1 I_56844 (I684974,I2683,I969022,I969082,);
DFFARX1 I_56845 (I969082,I2683,I969022,I969099,);
not I_56846 (I969014,I969099);
not I_56847 (I969121,I684980);
nor I_56848 (I969138,I684980,I684974);
not I_56849 (I969155,I684983);
nand I_56850 (I969172,I969121,I969155);
nor I_56851 (I969189,I684983,I684980);
and I_56852 (I968993,I969189,I969056);
not I_56853 (I969220,I684992);
nand I_56854 (I969237,I969220,I684986);
nor I_56855 (I969254,I684992,I684989);
not I_56856 (I969271,I969254);
nand I_56857 (I968996,I969138,I969271);
DFFARX1 I_56858 (I969254,I2683,I969022,I969011,);
nor I_56859 (I969316,I684971,I684983);
nor I_56860 (I969333,I969316,I684974);
and I_56861 (I969350,I969333,I969237);
DFFARX1 I_56862 (I969350,I2683,I969022,I969008,);
nor I_56863 (I969005,I969316,I969172);
or I_56864 (I969002,I969254,I969316);
nor I_56865 (I969409,I684971,I684977);
DFFARX1 I_56866 (I969409,I2683,I969022,I969435,);
not I_56867 (I969443,I969435);
nand I_56868 (I969460,I969443,I969121);
nor I_56869 (I969477,I969460,I684974);
DFFARX1 I_56870 (I969477,I2683,I969022,I968990,);
nor I_56871 (I969508,I969443,I969172);
nor I_56872 (I968999,I969316,I969508);
not I_56873 (I969566,I2690);
DFFARX1 I_56874 (I519683,I2683,I969566,I969592,);
nand I_56875 (I969600,I969592,I519698);
DFFARX1 I_56876 (I519692,I2683,I969566,I969626,);
DFFARX1 I_56877 (I969626,I2683,I969566,I969643,);
not I_56878 (I969558,I969643);
not I_56879 (I969665,I519695);
nor I_56880 (I969682,I519695,I519701);
not I_56881 (I969699,I519683);
nand I_56882 (I969716,I969665,I969699);
nor I_56883 (I969733,I519683,I519695);
and I_56884 (I969537,I969733,I969600);
not I_56885 (I969764,I519680);
nand I_56886 (I969781,I969764,I519686);
nor I_56887 (I969798,I519680,I519680);
not I_56888 (I969815,I969798);
nand I_56889 (I969540,I969682,I969815);
DFFARX1 I_56890 (I969798,I2683,I969566,I969555,);
nor I_56891 (I969860,I519689,I519683);
nor I_56892 (I969877,I969860,I519701);
and I_56893 (I969894,I969877,I969781);
DFFARX1 I_56894 (I969894,I2683,I969566,I969552,);
nor I_56895 (I969549,I969860,I969716);
or I_56896 (I969546,I969798,I969860);
nor I_56897 (I969953,I519689,I519704);
DFFARX1 I_56898 (I969953,I2683,I969566,I969979,);
not I_56899 (I969987,I969979);
nand I_56900 (I970004,I969987,I969665);
nor I_56901 (I970021,I970004,I519701);
DFFARX1 I_56902 (I970021,I2683,I969566,I969534,);
nor I_56903 (I970052,I969987,I969716);
nor I_56904 (I969543,I969860,I970052);
not I_56905 (I970110,I2690);
DFFARX1 I_56906 (I534711,I2683,I970110,I970136,);
nand I_56907 (I970144,I970136,I534726);
DFFARX1 I_56908 (I534720,I2683,I970110,I970170,);
DFFARX1 I_56909 (I970170,I2683,I970110,I970187,);
not I_56910 (I970102,I970187);
not I_56911 (I970209,I534723);
nor I_56912 (I970226,I534723,I534729);
not I_56913 (I970243,I534711);
nand I_56914 (I970260,I970209,I970243);
nor I_56915 (I970277,I534711,I534723);
and I_56916 (I970081,I970277,I970144);
not I_56917 (I970308,I534708);
nand I_56918 (I970325,I970308,I534714);
nor I_56919 (I970342,I534708,I534708);
not I_56920 (I970359,I970342);
nand I_56921 (I970084,I970226,I970359);
DFFARX1 I_56922 (I970342,I2683,I970110,I970099,);
nor I_56923 (I970404,I534717,I534711);
nor I_56924 (I970421,I970404,I534729);
and I_56925 (I970438,I970421,I970325);
DFFARX1 I_56926 (I970438,I2683,I970110,I970096,);
nor I_56927 (I970093,I970404,I970260);
or I_56928 (I970090,I970342,I970404);
nor I_56929 (I970497,I534717,I534732);
DFFARX1 I_56930 (I970497,I2683,I970110,I970523,);
not I_56931 (I970531,I970523);
nand I_56932 (I970548,I970531,I970209);
nor I_56933 (I970565,I970548,I534729);
DFFARX1 I_56934 (I970565,I2683,I970110,I970078,);
nor I_56935 (I970596,I970531,I970260);
nor I_56936 (I970087,I970404,I970596);
not I_56937 (I970654,I2690);
DFFARX1 I_56938 (I362794,I2683,I970654,I970680,);
nand I_56939 (I970688,I970680,I362791);
DFFARX1 I_56940 (I362770,I2683,I970654,I970714,);
DFFARX1 I_56941 (I970714,I2683,I970654,I970731,);
not I_56942 (I970646,I970731);
not I_56943 (I970753,I362785);
nor I_56944 (I970770,I362785,I362788);
not I_56945 (I970787,I362779);
nand I_56946 (I970804,I970753,I970787);
nor I_56947 (I970821,I362779,I362785);
and I_56948 (I970625,I970821,I970688);
not I_56949 (I970852,I362776);
nand I_56950 (I970869,I970852,I362797);
nor I_56951 (I970886,I362776,I362773);
not I_56952 (I970903,I970886);
nand I_56953 (I970628,I970770,I970903);
DFFARX1 I_56954 (I970886,I2683,I970654,I970643,);
nor I_56955 (I970948,I362782,I362779);
nor I_56956 (I970965,I970948,I362788);
and I_56957 (I970982,I970965,I970869);
DFFARX1 I_56958 (I970982,I2683,I970654,I970640,);
nor I_56959 (I970637,I970948,I970804);
or I_56960 (I970634,I970886,I970948);
nor I_56961 (I971041,I362782,I362770);
DFFARX1 I_56962 (I971041,I2683,I970654,I971067,);
not I_56963 (I971075,I971067);
nand I_56964 (I971092,I971075,I970753);
nor I_56965 (I971109,I971092,I362788);
DFFARX1 I_56966 (I971109,I2683,I970654,I970622,);
nor I_56967 (I971140,I971075,I970804);
nor I_56968 (I970631,I970948,I971140);
not I_56969 (I971198,I2690);
DFFARX1 I_56970 (I521995,I2683,I971198,I971224,);
nand I_56971 (I971232,I971224,I522010);
DFFARX1 I_56972 (I522004,I2683,I971198,I971258,);
DFFARX1 I_56973 (I971258,I2683,I971198,I971275,);
not I_56974 (I971190,I971275);
not I_56975 (I971297,I522007);
nor I_56976 (I971314,I522007,I522013);
not I_56977 (I971331,I521995);
nand I_56978 (I971348,I971297,I971331);
nor I_56979 (I971365,I521995,I522007);
and I_56980 (I971169,I971365,I971232);
not I_56981 (I971396,I521992);
nand I_56982 (I971413,I971396,I521998);
nor I_56983 (I971430,I521992,I521992);
not I_56984 (I971447,I971430);
nand I_56985 (I971172,I971314,I971447);
DFFARX1 I_56986 (I971430,I2683,I971198,I971187,);
nor I_56987 (I971492,I522001,I521995);
nor I_56988 (I971509,I971492,I522013);
and I_56989 (I971526,I971509,I971413);
DFFARX1 I_56990 (I971526,I2683,I971198,I971184,);
nor I_56991 (I971181,I971492,I971348);
or I_56992 (I971178,I971430,I971492);
nor I_56993 (I971585,I522001,I522016);
DFFARX1 I_56994 (I971585,I2683,I971198,I971611,);
not I_56995 (I971619,I971611);
nand I_56996 (I971636,I971619,I971297);
nor I_56997 (I971653,I971636,I522013);
DFFARX1 I_56998 (I971653,I2683,I971198,I971166,);
nor I_56999 (I971684,I971619,I971348);
nor I_57000 (I971175,I971492,I971684);
not I_57001 (I971742,I2690);
DFFARX1 I_57002 (I192609,I2683,I971742,I971768,);
nand I_57003 (I971776,I971768,I192624);
DFFARX1 I_57004 (I192621,I2683,I971742,I971802,);
DFFARX1 I_57005 (I971802,I2683,I971742,I971819,);
not I_57006 (I971734,I971819);
not I_57007 (I971841,I192600);
nor I_57008 (I971858,I192600,I192606);
not I_57009 (I971875,I192612);
nand I_57010 (I971892,I971841,I971875);
nor I_57011 (I971909,I192612,I192600);
and I_57012 (I971713,I971909,I971776);
not I_57013 (I971940,I192618);
nand I_57014 (I971957,I971940,I192600);
nor I_57015 (I971974,I192618,I192603);
not I_57016 (I971991,I971974);
nand I_57017 (I971716,I971858,I971991);
DFFARX1 I_57018 (I971974,I2683,I971742,I971731,);
nor I_57019 (I972036,I192603,I192612);
nor I_57020 (I972053,I972036,I192606);
and I_57021 (I972070,I972053,I971957);
DFFARX1 I_57022 (I972070,I2683,I971742,I971728,);
nor I_57023 (I971725,I972036,I971892);
or I_57024 (I971722,I971974,I972036);
nor I_57025 (I972129,I192603,I192615);
DFFARX1 I_57026 (I972129,I2683,I971742,I972155,);
not I_57027 (I972163,I972155);
nand I_57028 (I972180,I972163,I971841);
nor I_57029 (I972197,I972180,I192606);
DFFARX1 I_57030 (I972197,I2683,I971742,I971710,);
nor I_57031 (I972228,I972163,I971892);
nor I_57032 (I971719,I972036,I972228);
not I_57033 (I972286,I2690);
DFFARX1 I_57034 (I278581,I2683,I972286,I972312,);
nand I_57035 (I972320,I972312,I278584);
DFFARX1 I_57036 (I278578,I2683,I972286,I972346,);
DFFARX1 I_57037 (I972346,I2683,I972286,I972363,);
not I_57038 (I972278,I972363);
not I_57039 (I972385,I278587);
nor I_57040 (I972402,I278587,I278572);
not I_57041 (I972419,I278596);
nand I_57042 (I972436,I972385,I972419);
nor I_57043 (I972453,I278596,I278587);
and I_57044 (I972257,I972453,I972320);
not I_57045 (I972484,I278575);
nand I_57046 (I972501,I972484,I278593);
nor I_57047 (I972518,I278575,I278569);
not I_57048 (I972535,I972518);
nand I_57049 (I972260,I972402,I972535);
DFFARX1 I_57050 (I972518,I2683,I972286,I972275,);
nor I_57051 (I972580,I278590,I278596);
nor I_57052 (I972597,I972580,I278572);
and I_57053 (I972614,I972597,I972501);
DFFARX1 I_57054 (I972614,I2683,I972286,I972272,);
nor I_57055 (I972269,I972580,I972436);
or I_57056 (I972266,I972518,I972580);
nor I_57057 (I972673,I278590,I278569);
DFFARX1 I_57058 (I972673,I2683,I972286,I972699,);
not I_57059 (I972707,I972699);
nand I_57060 (I972724,I972707,I972385);
nor I_57061 (I972741,I972724,I278572);
DFFARX1 I_57062 (I972741,I2683,I972286,I972254,);
nor I_57063 (I972772,I972707,I972436);
nor I_57064 (I972263,I972580,I972772);
not I_57065 (I972830,I2690);
DFFARX1 I_57066 (I231678,I2683,I972830,I972856,);
nand I_57067 (I972864,I972856,I231681);
DFFARX1 I_57068 (I231675,I2683,I972830,I972890,);
DFFARX1 I_57069 (I972890,I2683,I972830,I972907,);
not I_57070 (I972822,I972907);
not I_57071 (I972929,I231684);
nor I_57072 (I972946,I231684,I231669);
not I_57073 (I972963,I231693);
nand I_57074 (I972980,I972929,I972963);
nor I_57075 (I972997,I231693,I231684);
and I_57076 (I972801,I972997,I972864);
not I_57077 (I973028,I231672);
nand I_57078 (I973045,I973028,I231690);
nor I_57079 (I973062,I231672,I231666);
not I_57080 (I973079,I973062);
nand I_57081 (I972804,I972946,I973079);
DFFARX1 I_57082 (I973062,I2683,I972830,I972819,);
nor I_57083 (I973124,I231687,I231693);
nor I_57084 (I973141,I973124,I231669);
and I_57085 (I973158,I973141,I973045);
DFFARX1 I_57086 (I973158,I2683,I972830,I972816,);
nor I_57087 (I972813,I973124,I972980);
or I_57088 (I972810,I973062,I973124);
nor I_57089 (I973217,I231687,I231666);
DFFARX1 I_57090 (I973217,I2683,I972830,I973243,);
not I_57091 (I973251,I973243);
nand I_57092 (I973268,I973251,I972929);
nor I_57093 (I973285,I973268,I231669);
DFFARX1 I_57094 (I973285,I2683,I972830,I972798,);
nor I_57095 (I973316,I973251,I972980);
nor I_57096 (I972807,I973124,I973316);
not I_57097 (I973374,I2690);
DFFARX1 I_57098 (I942086,I2683,I973374,I973400,);
nand I_57099 (I973408,I973400,I942065);
DFFARX1 I_57100 (I942062,I2683,I973374,I973434,);
DFFARX1 I_57101 (I973434,I2683,I973374,I973451,);
not I_57102 (I973366,I973451);
not I_57103 (I973473,I942074);
nor I_57104 (I973490,I942074,I942083);
not I_57105 (I973507,I942071);
nand I_57106 (I973524,I973473,I973507);
nor I_57107 (I973541,I942071,I942074);
and I_57108 (I973345,I973541,I973408);
not I_57109 (I973572,I942080);
nand I_57110 (I973589,I973572,I942077);
nor I_57111 (I973606,I942080,I942062);
not I_57112 (I973623,I973606);
nand I_57113 (I973348,I973490,I973623);
DFFARX1 I_57114 (I973606,I2683,I973374,I973363,);
nor I_57115 (I973668,I942065,I942071);
nor I_57116 (I973685,I973668,I942083);
and I_57117 (I973702,I973685,I973589);
DFFARX1 I_57118 (I973702,I2683,I973374,I973360,);
nor I_57119 (I973357,I973668,I973524);
or I_57120 (I973354,I973606,I973668);
nor I_57121 (I973761,I942065,I942068);
DFFARX1 I_57122 (I973761,I2683,I973374,I973787,);
not I_57123 (I973795,I973787);
nand I_57124 (I973812,I973795,I973473);
nor I_57125 (I973829,I973812,I942083);
DFFARX1 I_57126 (I973829,I2683,I973374,I973342,);
nor I_57127 (I973860,I973795,I973524);
nor I_57128 (I973351,I973668,I973860);
not I_57129 (I973918,I2690);
DFFARX1 I_57130 (I436469,I2683,I973918,I973944,);
nand I_57131 (I973952,I973944,I436457);
DFFARX1 I_57132 (I436463,I2683,I973918,I973978,);
DFFARX1 I_57133 (I973978,I2683,I973918,I973995,);
not I_57134 (I973910,I973995);
not I_57135 (I974017,I436448);
nor I_57136 (I974034,I436448,I436460);
not I_57137 (I974051,I436451);
nand I_57138 (I974068,I974017,I974051);
nor I_57139 (I974085,I436451,I436448);
and I_57140 (I973889,I974085,I973952);
not I_57141 (I974116,I436466);
nand I_57142 (I974133,I974116,I436448);
nor I_57143 (I974150,I436466,I436472);
not I_57144 (I974167,I974150);
nand I_57145 (I973892,I974034,I974167);
DFFARX1 I_57146 (I974150,I2683,I973918,I973907,);
nor I_57147 (I974212,I436454,I436451);
nor I_57148 (I974229,I974212,I436460);
and I_57149 (I974246,I974229,I974133);
DFFARX1 I_57150 (I974246,I2683,I973918,I973904,);
nor I_57151 (I973901,I974212,I974068);
or I_57152 (I973898,I974150,I974212);
nor I_57153 (I974305,I436454,I436451);
DFFARX1 I_57154 (I974305,I2683,I973918,I974331,);
not I_57155 (I974339,I974331);
nand I_57156 (I974356,I974339,I974017);
nor I_57157 (I974373,I974356,I436460);
DFFARX1 I_57158 (I974373,I2683,I973918,I973886,);
nor I_57159 (I974404,I974339,I974068);
nor I_57160 (I973895,I974212,I974404);
not I_57161 (I974462,I2690);
DFFARX1 I_57162 (I593089,I2683,I974462,I974488,);
nand I_57163 (I974496,I974488,I593104);
DFFARX1 I_57164 (I593098,I2683,I974462,I974522,);
DFFARX1 I_57165 (I974522,I2683,I974462,I974539,);
not I_57166 (I974454,I974539);
not I_57167 (I974561,I593101);
nor I_57168 (I974578,I593101,I593107);
not I_57169 (I974595,I593089);
nand I_57170 (I974612,I974561,I974595);
nor I_57171 (I974629,I593089,I593101);
and I_57172 (I974433,I974629,I974496);
not I_57173 (I974660,I593086);
nand I_57174 (I974677,I974660,I593092);
nor I_57175 (I974694,I593086,I593086);
not I_57176 (I974711,I974694);
nand I_57177 (I974436,I974578,I974711);
DFFARX1 I_57178 (I974694,I2683,I974462,I974451,);
nor I_57179 (I974756,I593095,I593089);
nor I_57180 (I974773,I974756,I593107);
and I_57181 (I974790,I974773,I974677);
DFFARX1 I_57182 (I974790,I2683,I974462,I974448,);
nor I_57183 (I974445,I974756,I974612);
or I_57184 (I974442,I974694,I974756);
nor I_57185 (I974849,I593095,I593110);
DFFARX1 I_57186 (I974849,I2683,I974462,I974875,);
not I_57187 (I974883,I974875);
nand I_57188 (I974900,I974883,I974561);
nor I_57189 (I974917,I974900,I593107);
DFFARX1 I_57190 (I974917,I2683,I974462,I974430,);
nor I_57191 (I974948,I974883,I974612);
nor I_57192 (I974439,I974756,I974948);
not I_57193 (I975006,I2690);
DFFARX1 I_57194 (I655465,I2683,I975006,I975032,);
nand I_57195 (I975040,I975032,I655459);
DFFARX1 I_57196 (I655462,I2683,I975006,I975066,);
DFFARX1 I_57197 (I975066,I2683,I975006,I975083,);
not I_57198 (I974998,I975083);
not I_57199 (I975105,I655468);
nor I_57200 (I975122,I655468,I655462);
not I_57201 (I975139,I655471);
nand I_57202 (I975156,I975105,I975139);
nor I_57203 (I975173,I655471,I655468);
and I_57204 (I974977,I975173,I975040);
not I_57205 (I975204,I655480);
nand I_57206 (I975221,I975204,I655474);
nor I_57207 (I975238,I655480,I655477);
not I_57208 (I975255,I975238);
nand I_57209 (I974980,I975122,I975255);
DFFARX1 I_57210 (I975238,I2683,I975006,I974995,);
nor I_57211 (I975300,I655459,I655471);
nor I_57212 (I975317,I975300,I655462);
and I_57213 (I975334,I975317,I975221);
DFFARX1 I_57214 (I975334,I2683,I975006,I974992,);
nor I_57215 (I974989,I975300,I975156);
or I_57216 (I974986,I975238,I975300);
nor I_57217 (I975393,I655459,I655465);
DFFARX1 I_57218 (I975393,I2683,I975006,I975419,);
not I_57219 (I975427,I975419);
nand I_57220 (I975444,I975427,I975105);
nor I_57221 (I975461,I975444,I655462);
DFFARX1 I_57222 (I975461,I2683,I975006,I974974,);
nor I_57223 (I975492,I975427,I975156);
nor I_57224 (I974983,I975300,I975492);
not I_57225 (I975550,I2690);
DFFARX1 I_57226 (I248015,I2683,I975550,I975576,);
nand I_57227 (I975584,I975576,I248018);
DFFARX1 I_57228 (I248012,I2683,I975550,I975610,);
DFFARX1 I_57229 (I975610,I2683,I975550,I975627,);
not I_57230 (I975542,I975627);
not I_57231 (I975649,I248021);
nor I_57232 (I975666,I248021,I248006);
not I_57233 (I975683,I248030);
nand I_57234 (I975700,I975649,I975683);
nor I_57235 (I975717,I248030,I248021);
and I_57236 (I975521,I975717,I975584);
not I_57237 (I975748,I248009);
nand I_57238 (I975765,I975748,I248027);
nor I_57239 (I975782,I248009,I248003);
not I_57240 (I975799,I975782);
nand I_57241 (I975524,I975666,I975799);
DFFARX1 I_57242 (I975782,I2683,I975550,I975539,);
nor I_57243 (I975844,I248024,I248030);
nor I_57244 (I975861,I975844,I248006);
and I_57245 (I975878,I975861,I975765);
DFFARX1 I_57246 (I975878,I2683,I975550,I975536,);
nor I_57247 (I975533,I975844,I975700);
or I_57248 (I975530,I975782,I975844);
nor I_57249 (I975937,I248024,I248003);
DFFARX1 I_57250 (I975937,I2683,I975550,I975963,);
not I_57251 (I975971,I975963);
nand I_57252 (I975988,I975971,I975649);
nor I_57253 (I976005,I975988,I248006);
DFFARX1 I_57254 (I976005,I2683,I975550,I975518,);
nor I_57255 (I976036,I975971,I975700);
nor I_57256 (I975527,I975844,I976036);
not I_57257 (I976094,I2690);
DFFARX1 I_57258 (I363882,I2683,I976094,I976120,);
nand I_57259 (I976128,I976120,I363879);
DFFARX1 I_57260 (I363858,I2683,I976094,I976154,);
DFFARX1 I_57261 (I976154,I2683,I976094,I976171,);
not I_57262 (I976086,I976171);
not I_57263 (I976193,I363873);
nor I_57264 (I976210,I363873,I363876);
not I_57265 (I976227,I363867);
nand I_57266 (I976244,I976193,I976227);
nor I_57267 (I976261,I363867,I363873);
and I_57268 (I976065,I976261,I976128);
not I_57269 (I976292,I363864);
nand I_57270 (I976309,I976292,I363885);
nor I_57271 (I976326,I363864,I363861);
not I_57272 (I976343,I976326);
nand I_57273 (I976068,I976210,I976343);
DFFARX1 I_57274 (I976326,I2683,I976094,I976083,);
nor I_57275 (I976388,I363870,I363867);
nor I_57276 (I976405,I976388,I363876);
and I_57277 (I976422,I976405,I976309);
DFFARX1 I_57278 (I976422,I2683,I976094,I976080,);
nor I_57279 (I976077,I976388,I976244);
or I_57280 (I976074,I976326,I976388);
nor I_57281 (I976481,I363870,I363858);
DFFARX1 I_57282 (I976481,I2683,I976094,I976507,);
not I_57283 (I976515,I976507);
nand I_57284 (I976532,I976515,I976193);
nor I_57285 (I976549,I976532,I363876);
DFFARX1 I_57286 (I976549,I2683,I976094,I976062,);
nor I_57287 (I976580,I976515,I976244);
nor I_57288 (I976071,I976388,I976580);
not I_57289 (I976638,I2690);
DFFARX1 I_57290 (I571125,I2683,I976638,I976664,);
nand I_57291 (I976672,I976664,I571140);
DFFARX1 I_57292 (I571134,I2683,I976638,I976698,);
DFFARX1 I_57293 (I976698,I2683,I976638,I976715,);
not I_57294 (I976630,I976715);
not I_57295 (I976737,I571137);
nor I_57296 (I976754,I571137,I571143);
not I_57297 (I976771,I571125);
nand I_57298 (I976788,I976737,I976771);
nor I_57299 (I976805,I571125,I571137);
and I_57300 (I976609,I976805,I976672);
not I_57301 (I976836,I571122);
nand I_57302 (I976853,I976836,I571128);
nor I_57303 (I976870,I571122,I571122);
not I_57304 (I976887,I976870);
nand I_57305 (I976612,I976754,I976887);
DFFARX1 I_57306 (I976870,I2683,I976638,I976627,);
nor I_57307 (I976932,I571131,I571125);
nor I_57308 (I976949,I976932,I571143);
and I_57309 (I976966,I976949,I976853);
DFFARX1 I_57310 (I976966,I2683,I976638,I976624,);
nor I_57311 (I976621,I976932,I976788);
or I_57312 (I976618,I976870,I976932);
nor I_57313 (I977025,I571131,I571146);
DFFARX1 I_57314 (I977025,I2683,I976638,I977051,);
not I_57315 (I977059,I977051);
nand I_57316 (I977076,I977059,I976737);
nor I_57317 (I977093,I977076,I571143);
DFFARX1 I_57318 (I977093,I2683,I976638,I976606,);
nor I_57319 (I977124,I977059,I976788);
nor I_57320 (I976615,I976932,I977124);
not I_57321 (I977182,I2690);
DFFARX1 I_57322 (I631750,I2683,I977182,I977208,);
nand I_57323 (I977216,I977208,I631744);
DFFARX1 I_57324 (I631747,I2683,I977182,I977242,);
DFFARX1 I_57325 (I977242,I2683,I977182,I977259,);
not I_57326 (I977174,I977259);
not I_57327 (I977281,I631753);
nor I_57328 (I977298,I631753,I631747);
not I_57329 (I977315,I631756);
nand I_57330 (I977332,I977281,I977315);
nor I_57331 (I977349,I631756,I631753);
and I_57332 (I977153,I977349,I977216);
not I_57333 (I977380,I631765);
nand I_57334 (I977397,I977380,I631759);
nor I_57335 (I977414,I631765,I631762);
not I_57336 (I977431,I977414);
nand I_57337 (I977156,I977298,I977431);
DFFARX1 I_57338 (I977414,I2683,I977182,I977171,);
nor I_57339 (I977476,I631744,I631756);
nor I_57340 (I977493,I977476,I631747);
and I_57341 (I977510,I977493,I977397);
DFFARX1 I_57342 (I977510,I2683,I977182,I977168,);
nor I_57343 (I977165,I977476,I977332);
or I_57344 (I977162,I977414,I977476);
nor I_57345 (I977569,I631744,I631750);
DFFARX1 I_57346 (I977569,I2683,I977182,I977595,);
not I_57347 (I977603,I977595);
nand I_57348 (I977620,I977603,I977281);
nor I_57349 (I977637,I977620,I631747);
DFFARX1 I_57350 (I977637,I2683,I977182,I977150,);
nor I_57351 (I977668,I977603,I977332);
nor I_57352 (I977159,I977476,I977668);
not I_57353 (I977726,I2690);
DFFARX1 I_57354 (I1064421,I2683,I977726,I977752,);
nand I_57355 (I977760,I977752,I1064406);
DFFARX1 I_57356 (I1064400,I2683,I977726,I977786,);
DFFARX1 I_57357 (I977786,I2683,I977726,I977803,);
not I_57358 (I977718,I977803);
not I_57359 (I977825,I1064394);
nor I_57360 (I977842,I1064394,I1064415);
not I_57361 (I977859,I1064403);
nand I_57362 (I977876,I977825,I977859);
nor I_57363 (I977893,I1064403,I1064394);
and I_57364 (I977697,I977893,I977760);
not I_57365 (I977924,I1064412);
nand I_57366 (I977941,I977924,I1064418);
nor I_57367 (I977958,I1064412,I1064409);
not I_57368 (I977975,I977958);
nand I_57369 (I977700,I977842,I977975);
DFFARX1 I_57370 (I977958,I2683,I977726,I977715,);
nor I_57371 (I978020,I1064397,I1064403);
nor I_57372 (I978037,I978020,I1064415);
and I_57373 (I978054,I978037,I977941);
DFFARX1 I_57374 (I978054,I2683,I977726,I977712,);
nor I_57375 (I977709,I978020,I977876);
or I_57376 (I977706,I977958,I978020);
nor I_57377 (I978113,I1064397,I1064394);
DFFARX1 I_57378 (I978113,I2683,I977726,I978139,);
not I_57379 (I978147,I978139);
nand I_57380 (I978164,I978147,I977825);
nor I_57381 (I978181,I978164,I1064415);
DFFARX1 I_57382 (I978181,I2683,I977726,I977694,);
nor I_57383 (I978212,I978147,I977876);
nor I_57384 (I977703,I978020,I978212);
not I_57385 (I978270,I2690);
DFFARX1 I_57386 (I206294,I2683,I978270,I978296,);
nand I_57387 (I978304,I978296,I206309);
DFFARX1 I_57388 (I206306,I2683,I978270,I978330,);
DFFARX1 I_57389 (I978330,I2683,I978270,I978347,);
not I_57390 (I978262,I978347);
not I_57391 (I978369,I206285);
nor I_57392 (I978386,I206285,I206291);
not I_57393 (I978403,I206297);
nand I_57394 (I978420,I978369,I978403);
nor I_57395 (I978437,I206297,I206285);
and I_57396 (I978241,I978437,I978304);
not I_57397 (I978468,I206303);
nand I_57398 (I978485,I978468,I206285);
nor I_57399 (I978502,I206303,I206288);
not I_57400 (I978519,I978502);
nand I_57401 (I978244,I978386,I978519);
DFFARX1 I_57402 (I978502,I2683,I978270,I978259,);
nor I_57403 (I978564,I206288,I206297);
nor I_57404 (I978581,I978564,I206291);
and I_57405 (I978598,I978581,I978485);
DFFARX1 I_57406 (I978598,I2683,I978270,I978256,);
nor I_57407 (I978253,I978564,I978420);
or I_57408 (I978250,I978502,I978564);
nor I_57409 (I978657,I206288,I206300);
DFFARX1 I_57410 (I978657,I2683,I978270,I978683,);
not I_57411 (I978691,I978683);
nand I_57412 (I978708,I978691,I978369);
nor I_57413 (I978725,I978708,I206291);
DFFARX1 I_57414 (I978725,I2683,I978270,I978238,);
nor I_57415 (I978756,I978691,I978420);
nor I_57416 (I978247,I978564,I978756);
not I_57417 (I978814,I2690);
DFFARX1 I_57418 (I88581,I2683,I978814,I978840,);
nand I_57419 (I978848,I978840,I88563);
DFFARX1 I_57420 (I88560,I2683,I978814,I978874,);
DFFARX1 I_57421 (I978874,I2683,I978814,I978891,);
not I_57422 (I978806,I978891);
not I_57423 (I978913,I88578);
nor I_57424 (I978930,I88578,I88572);
not I_57425 (I978947,I88560);
nand I_57426 (I978964,I978913,I978947);
nor I_57427 (I978981,I88560,I88578);
and I_57428 (I978785,I978981,I978848);
not I_57429 (I979012,I88569);
nand I_57430 (I979029,I979012,I88575);
nor I_57431 (I979046,I88569,I88563);
not I_57432 (I979063,I979046);
nand I_57433 (I978788,I978930,I979063);
DFFARX1 I_57434 (I979046,I2683,I978814,I978803,);
nor I_57435 (I979108,I88566,I88560);
nor I_57436 (I979125,I979108,I88572);
and I_57437 (I979142,I979125,I979029);
DFFARX1 I_57438 (I979142,I2683,I978814,I978800,);
nor I_57439 (I978797,I979108,I978964);
or I_57440 (I978794,I979046,I979108);
nor I_57441 (I979201,I88566,I88584);
DFFARX1 I_57442 (I979201,I2683,I978814,I979227,);
not I_57443 (I979235,I979227);
nand I_57444 (I979252,I979235,I978913);
nor I_57445 (I979269,I979252,I88572);
DFFARX1 I_57446 (I979269,I2683,I978814,I978782,);
nor I_57447 (I979300,I979235,I978964);
nor I_57448 (I978791,I979108,I979300);
not I_57449 (I979358,I2690);
DFFARX1 I_57450 (I463635,I2683,I979358,I979384,);
nand I_57451 (I979392,I979384,I463623);
DFFARX1 I_57452 (I463629,I2683,I979358,I979418,);
DFFARX1 I_57453 (I979418,I2683,I979358,I979435,);
not I_57454 (I979350,I979435);
not I_57455 (I979457,I463614);
nor I_57456 (I979474,I463614,I463626);
not I_57457 (I979491,I463617);
nand I_57458 (I979508,I979457,I979491);
nor I_57459 (I979525,I463617,I463614);
and I_57460 (I979329,I979525,I979392);
not I_57461 (I979556,I463632);
nand I_57462 (I979573,I979556,I463614);
nor I_57463 (I979590,I463632,I463638);
not I_57464 (I979607,I979590);
nand I_57465 (I979332,I979474,I979607);
DFFARX1 I_57466 (I979590,I2683,I979358,I979347,);
nor I_57467 (I979652,I463620,I463617);
nor I_57468 (I979669,I979652,I463626);
and I_57469 (I979686,I979669,I979573);
DFFARX1 I_57470 (I979686,I2683,I979358,I979344,);
nor I_57471 (I979341,I979652,I979508);
or I_57472 (I979338,I979590,I979652);
nor I_57473 (I979745,I463620,I463617);
DFFARX1 I_57474 (I979745,I2683,I979358,I979771,);
not I_57475 (I979779,I979771);
nand I_57476 (I979796,I979779,I979457);
nor I_57477 (I979813,I979796,I463626);
DFFARX1 I_57478 (I979813,I2683,I979358,I979326,);
nor I_57479 (I979844,I979779,I979508);
nor I_57480 (I979335,I979652,I979844);
not I_57481 (I979902,I2690);
DFFARX1 I_57482 (I777485,I2683,I979902,I979928,);
nand I_57483 (I979936,I979928,I777485);
DFFARX1 I_57484 (I777497,I2683,I979902,I979962,);
DFFARX1 I_57485 (I979962,I2683,I979902,I979979,);
not I_57486 (I979894,I979979);
not I_57487 (I980001,I777491);
nor I_57488 (I980018,I777491,I777512);
not I_57489 (I980035,I777500);
nand I_57490 (I980052,I980001,I980035);
nor I_57491 (I980069,I777500,I777491);
and I_57492 (I979873,I980069,I979936);
not I_57493 (I980100,I777494);
nand I_57494 (I980117,I980100,I777509);
nor I_57495 (I980134,I777494,I777503);
not I_57496 (I980151,I980134);
nand I_57497 (I979876,I980018,I980151);
DFFARX1 I_57498 (I980134,I2683,I979902,I979891,);
nor I_57499 (I980196,I777506,I777500);
nor I_57500 (I980213,I980196,I777512);
and I_57501 (I980230,I980213,I980117);
DFFARX1 I_57502 (I980230,I2683,I979902,I979888,);
nor I_57503 (I979885,I980196,I980052);
or I_57504 (I979882,I980134,I980196);
nor I_57505 (I980289,I777506,I777488);
DFFARX1 I_57506 (I980289,I2683,I979902,I980315,);
not I_57507 (I980323,I980315);
nand I_57508 (I980340,I980323,I980001);
nor I_57509 (I980357,I980340,I777512);
DFFARX1 I_57510 (I980357,I2683,I979902,I979870,);
nor I_57511 (I980388,I980323,I980052);
nor I_57512 (I979879,I980196,I980388);
not I_57513 (I980446,I2690);
DFFARX1 I_57514 (I538179,I2683,I980446,I980472,);
nand I_57515 (I980480,I980472,I538194);
DFFARX1 I_57516 (I538188,I2683,I980446,I980506,);
DFFARX1 I_57517 (I980506,I2683,I980446,I980523,);
not I_57518 (I980438,I980523);
not I_57519 (I980545,I538191);
nor I_57520 (I980562,I538191,I538197);
not I_57521 (I980579,I538179);
nand I_57522 (I980596,I980545,I980579);
nor I_57523 (I980613,I538179,I538191);
and I_57524 (I980417,I980613,I980480);
not I_57525 (I980644,I538176);
nand I_57526 (I980661,I980644,I538182);
nor I_57527 (I980678,I538176,I538176);
not I_57528 (I980695,I980678);
nand I_57529 (I980420,I980562,I980695);
DFFARX1 I_57530 (I980678,I2683,I980446,I980435,);
nor I_57531 (I980740,I538185,I538179);
nor I_57532 (I980757,I980740,I538197);
and I_57533 (I980774,I980757,I980661);
DFFARX1 I_57534 (I980774,I2683,I980446,I980432,);
nor I_57535 (I980429,I980740,I980596);
or I_57536 (I980426,I980678,I980740);
nor I_57537 (I980833,I538185,I538200);
DFFARX1 I_57538 (I980833,I2683,I980446,I980859,);
not I_57539 (I980867,I980859);
nand I_57540 (I980884,I980867,I980545);
nor I_57541 (I980901,I980884,I538197);
DFFARX1 I_57542 (I980901,I2683,I980446,I980414,);
nor I_57543 (I980932,I980867,I980596);
nor I_57544 (I980423,I980740,I980932);
not I_57545 (I980990,I2690);
DFFARX1 I_57546 (I64866,I2683,I980990,I981016,);
nand I_57547 (I981024,I981016,I64848);
DFFARX1 I_57548 (I64845,I2683,I980990,I981050,);
DFFARX1 I_57549 (I981050,I2683,I980990,I981067,);
not I_57550 (I980982,I981067);
not I_57551 (I981089,I64863);
nor I_57552 (I981106,I64863,I64857);
not I_57553 (I981123,I64845);
nand I_57554 (I981140,I981089,I981123);
nor I_57555 (I981157,I64845,I64863);
and I_57556 (I980961,I981157,I981024);
not I_57557 (I981188,I64854);
nand I_57558 (I981205,I981188,I64860);
nor I_57559 (I981222,I64854,I64848);
not I_57560 (I981239,I981222);
nand I_57561 (I980964,I981106,I981239);
DFFARX1 I_57562 (I981222,I2683,I980990,I980979,);
nor I_57563 (I981284,I64851,I64845);
nor I_57564 (I981301,I981284,I64857);
and I_57565 (I981318,I981301,I981205);
DFFARX1 I_57566 (I981318,I2683,I980990,I980976,);
nor I_57567 (I980973,I981284,I981140);
or I_57568 (I980970,I981222,I981284);
nor I_57569 (I981377,I64851,I64869);
DFFARX1 I_57570 (I981377,I2683,I980990,I981403,);
not I_57571 (I981411,I981403);
nand I_57572 (I981428,I981411,I981089);
nor I_57573 (I981445,I981428,I64857);
DFFARX1 I_57574 (I981445,I2683,I980990,I980958,);
nor I_57575 (I981476,I981411,I981140);
nor I_57576 (I980967,I981284,I981476);
not I_57577 (I981534,I2690);
DFFARX1 I_57578 (I141439,I2683,I981534,I981560,);
nand I_57579 (I981568,I981560,I141454);
DFFARX1 I_57580 (I141451,I2683,I981534,I981594,);
DFFARX1 I_57581 (I981594,I2683,I981534,I981611,);
not I_57582 (I981526,I981611);
not I_57583 (I981633,I141430);
nor I_57584 (I981650,I141430,I141436);
not I_57585 (I981667,I141442);
nand I_57586 (I981684,I981633,I981667);
nor I_57587 (I981701,I141442,I141430);
and I_57588 (I981505,I981701,I981568);
not I_57589 (I981732,I141448);
nand I_57590 (I981749,I981732,I141430);
nor I_57591 (I981766,I141448,I141433);
not I_57592 (I981783,I981766);
nand I_57593 (I981508,I981650,I981783);
DFFARX1 I_57594 (I981766,I2683,I981534,I981523,);
nor I_57595 (I981828,I141433,I141442);
nor I_57596 (I981845,I981828,I141436);
and I_57597 (I981862,I981845,I981749);
DFFARX1 I_57598 (I981862,I2683,I981534,I981520,);
nor I_57599 (I981517,I981828,I981684);
or I_57600 (I981514,I981766,I981828);
nor I_57601 (I981921,I141433,I141445);
DFFARX1 I_57602 (I981921,I2683,I981534,I981947,);
not I_57603 (I981955,I981947);
nand I_57604 (I981972,I981955,I981633);
nor I_57605 (I981989,I981972,I141436);
DFFARX1 I_57606 (I981989,I2683,I981534,I981502,);
nor I_57607 (I982020,I981955,I981684);
nor I_57608 (I981511,I981828,I982020);
not I_57609 (I982078,I2690);
DFFARX1 I_57610 (I1050736,I2683,I982078,I982104,);
nand I_57611 (I982112,I982104,I1050721);
DFFARX1 I_57612 (I1050715,I2683,I982078,I982138,);
DFFARX1 I_57613 (I982138,I2683,I982078,I982155,);
not I_57614 (I982070,I982155);
not I_57615 (I982177,I1050709);
nor I_57616 (I982194,I1050709,I1050730);
not I_57617 (I982211,I1050718);
nand I_57618 (I982228,I982177,I982211);
nor I_57619 (I982245,I1050718,I1050709);
and I_57620 (I982049,I982245,I982112);
not I_57621 (I982276,I1050727);
nand I_57622 (I982293,I982276,I1050733);
nor I_57623 (I982310,I1050727,I1050724);
not I_57624 (I982327,I982310);
nand I_57625 (I982052,I982194,I982327);
DFFARX1 I_57626 (I982310,I2683,I982078,I982067,);
nor I_57627 (I982372,I1050712,I1050718);
nor I_57628 (I982389,I982372,I1050730);
and I_57629 (I982406,I982389,I982293);
DFFARX1 I_57630 (I982406,I2683,I982078,I982064,);
nor I_57631 (I982061,I982372,I982228);
or I_57632 (I982058,I982310,I982372);
nor I_57633 (I982465,I1050712,I1050709);
DFFARX1 I_57634 (I982465,I2683,I982078,I982491,);
not I_57635 (I982499,I982491);
nand I_57636 (I982516,I982499,I982177);
nor I_57637 (I982533,I982516,I1050730);
DFFARX1 I_57638 (I982533,I2683,I982078,I982046,);
nor I_57639 (I982564,I982499,I982228);
nor I_57640 (I982055,I982372,I982564);
not I_57641 (I982622,I2690);
DFFARX1 I_57642 (I51164,I2683,I982622,I982648,);
nand I_57643 (I982656,I982648,I51146);
DFFARX1 I_57644 (I51143,I2683,I982622,I982682,);
DFFARX1 I_57645 (I982682,I2683,I982622,I982699,);
not I_57646 (I982614,I982699);
not I_57647 (I982721,I51161);
nor I_57648 (I982738,I51161,I51155);
not I_57649 (I982755,I51143);
nand I_57650 (I982772,I982721,I982755);
nor I_57651 (I982789,I51143,I51161);
and I_57652 (I982593,I982789,I982656);
not I_57653 (I982820,I51152);
nand I_57654 (I982837,I982820,I51158);
nor I_57655 (I982854,I51152,I51146);
not I_57656 (I982871,I982854);
nand I_57657 (I982596,I982738,I982871);
DFFARX1 I_57658 (I982854,I2683,I982622,I982611,);
nor I_57659 (I982916,I51149,I51143);
nor I_57660 (I982933,I982916,I51155);
and I_57661 (I982950,I982933,I982837);
DFFARX1 I_57662 (I982950,I2683,I982622,I982608,);
nor I_57663 (I982605,I982916,I982772);
or I_57664 (I982602,I982854,I982916);
nor I_57665 (I983009,I51149,I51167);
DFFARX1 I_57666 (I983009,I2683,I982622,I983035,);
not I_57667 (I983043,I983035);
nand I_57668 (I983060,I983043,I982721);
nor I_57669 (I983077,I983060,I51155);
DFFARX1 I_57670 (I983077,I2683,I982622,I982590,);
nor I_57671 (I983108,I983043,I982772);
nor I_57672 (I982599,I982916,I983108);
not I_57673 (I983166,I2690);
DFFARX1 I_57674 (I640182,I2683,I983166,I983192,);
nand I_57675 (I983200,I983192,I640176);
DFFARX1 I_57676 (I640179,I2683,I983166,I983226,);
DFFARX1 I_57677 (I983226,I2683,I983166,I983243,);
not I_57678 (I983158,I983243);
not I_57679 (I983265,I640185);
nor I_57680 (I983282,I640185,I640179);
not I_57681 (I983299,I640188);
nand I_57682 (I983316,I983265,I983299);
nor I_57683 (I983333,I640188,I640185);
and I_57684 (I983137,I983333,I983200);
not I_57685 (I983364,I640197);
nand I_57686 (I983381,I983364,I640191);
nor I_57687 (I983398,I640197,I640194);
not I_57688 (I983415,I983398);
nand I_57689 (I983140,I983282,I983415);
DFFARX1 I_57690 (I983398,I2683,I983166,I983155,);
nor I_57691 (I983460,I640176,I640188);
nor I_57692 (I983477,I983460,I640179);
and I_57693 (I983494,I983477,I983381);
DFFARX1 I_57694 (I983494,I2683,I983166,I983152,);
nor I_57695 (I983149,I983460,I983316);
or I_57696 (I983146,I983398,I983460);
nor I_57697 (I983553,I640176,I640182);
DFFARX1 I_57698 (I983553,I2683,I983166,I983579,);
not I_57699 (I983587,I983579);
nand I_57700 (I983604,I983587,I983265);
nor I_57701 (I983621,I983604,I640179);
DFFARX1 I_57702 (I983621,I2683,I983166,I983134,);
nor I_57703 (I983652,I983587,I983316);
nor I_57704 (I983143,I983460,I983652);
not I_57705 (I983710,I2690);
DFFARX1 I_57706 (I387818,I2683,I983710,I983736,);
nand I_57707 (I983744,I983736,I387815);
DFFARX1 I_57708 (I387794,I2683,I983710,I983770,);
DFFARX1 I_57709 (I983770,I2683,I983710,I983787,);
not I_57710 (I983702,I983787);
not I_57711 (I983809,I387809);
nor I_57712 (I983826,I387809,I387812);
not I_57713 (I983843,I387803);
nand I_57714 (I983860,I983809,I983843);
nor I_57715 (I983877,I387803,I387809);
and I_57716 (I983681,I983877,I983744);
not I_57717 (I983908,I387800);
nand I_57718 (I983925,I983908,I387821);
nor I_57719 (I983942,I387800,I387797);
not I_57720 (I983959,I983942);
nand I_57721 (I983684,I983826,I983959);
DFFARX1 I_57722 (I983942,I2683,I983710,I983699,);
nor I_57723 (I984004,I387806,I387803);
nor I_57724 (I984021,I984004,I387812);
and I_57725 (I984038,I984021,I983925);
DFFARX1 I_57726 (I984038,I2683,I983710,I983696,);
nor I_57727 (I983693,I984004,I983860);
or I_57728 (I983690,I983942,I984004);
nor I_57729 (I984097,I387806,I387794);
DFFARX1 I_57730 (I984097,I2683,I983710,I984123,);
not I_57731 (I984131,I984123);
nand I_57732 (I984148,I984131,I983809);
nor I_57733 (I984165,I984148,I387812);
DFFARX1 I_57734 (I984165,I2683,I983710,I983678,);
nor I_57735 (I984196,I984131,I983860);
nor I_57736 (I983687,I984004,I984196);
not I_57737 (I984254,I2690);
DFFARX1 I_57738 (I617943,I2683,I984254,I984280,);
nand I_57739 (I984288,I984280,I617958);
DFFARX1 I_57740 (I617952,I2683,I984254,I984314,);
DFFARX1 I_57741 (I984314,I2683,I984254,I984331,);
not I_57742 (I984246,I984331);
not I_57743 (I984353,I617955);
nor I_57744 (I984370,I617955,I617961);
not I_57745 (I984387,I617943);
nand I_57746 (I984404,I984353,I984387);
nor I_57747 (I984421,I617943,I617955);
and I_57748 (I984225,I984421,I984288);
not I_57749 (I984452,I617940);
nand I_57750 (I984469,I984452,I617946);
nor I_57751 (I984486,I617940,I617940);
not I_57752 (I984503,I984486);
nand I_57753 (I984228,I984370,I984503);
DFFARX1 I_57754 (I984486,I2683,I984254,I984243,);
nor I_57755 (I984548,I617949,I617943);
nor I_57756 (I984565,I984548,I617961);
and I_57757 (I984582,I984565,I984469);
DFFARX1 I_57758 (I984582,I2683,I984254,I984240,);
nor I_57759 (I984237,I984548,I984404);
or I_57760 (I984234,I984486,I984548);
nor I_57761 (I984641,I617949,I617964);
DFFARX1 I_57762 (I984641,I2683,I984254,I984667,);
not I_57763 (I984675,I984667);
nand I_57764 (I984692,I984675,I984353);
nor I_57765 (I984709,I984692,I617961);
DFFARX1 I_57766 (I984709,I2683,I984254,I984222,);
nor I_57767 (I984740,I984675,I984404);
nor I_57768 (I984231,I984548,I984740);
not I_57769 (I984798,I2690);
DFFARX1 I_57770 (I846716,I2683,I984798,I984824,);
nand I_57771 (I984832,I984824,I846695);
DFFARX1 I_57772 (I846692,I2683,I984798,I984858,);
DFFARX1 I_57773 (I984858,I2683,I984798,I984875,);
not I_57774 (I984790,I984875);
not I_57775 (I984897,I846704);
nor I_57776 (I984914,I846704,I846713);
not I_57777 (I984931,I846701);
nand I_57778 (I984948,I984897,I984931);
nor I_57779 (I984965,I846701,I846704);
and I_57780 (I984769,I984965,I984832);
not I_57781 (I984996,I846710);
nand I_57782 (I985013,I984996,I846707);
nor I_57783 (I985030,I846710,I846692);
not I_57784 (I985047,I985030);
nand I_57785 (I984772,I984914,I985047);
DFFARX1 I_57786 (I985030,I2683,I984798,I984787,);
nor I_57787 (I985092,I846695,I846701);
nor I_57788 (I985109,I985092,I846713);
and I_57789 (I985126,I985109,I985013);
DFFARX1 I_57790 (I985126,I2683,I984798,I984784,);
nor I_57791 (I984781,I985092,I984948);
or I_57792 (I984778,I985030,I985092);
nor I_57793 (I985185,I846695,I846698);
DFFARX1 I_57794 (I985185,I2683,I984798,I985211,);
not I_57795 (I985219,I985211);
nand I_57796 (I985236,I985219,I984897);
nor I_57797 (I985253,I985236,I846713);
DFFARX1 I_57798 (I985253,I2683,I984798,I984766,);
nor I_57799 (I985284,I985219,I984948);
nor I_57800 (I984775,I985092,I985284);
not I_57801 (I985342,I2690);
DFFARX1 I_57802 (I1049546,I2683,I985342,I985368,);
nand I_57803 (I985376,I985368,I1049531);
DFFARX1 I_57804 (I1049525,I2683,I985342,I985402,);
DFFARX1 I_57805 (I985402,I2683,I985342,I985419,);
not I_57806 (I985334,I985419);
not I_57807 (I985441,I1049519);
nor I_57808 (I985458,I1049519,I1049540);
not I_57809 (I985475,I1049528);
nand I_57810 (I985492,I985441,I985475);
nor I_57811 (I985509,I1049528,I1049519);
and I_57812 (I985313,I985509,I985376);
not I_57813 (I985540,I1049537);
nand I_57814 (I985557,I985540,I1049543);
nor I_57815 (I985574,I1049537,I1049534);
not I_57816 (I985591,I985574);
nand I_57817 (I985316,I985458,I985591);
DFFARX1 I_57818 (I985574,I2683,I985342,I985331,);
nor I_57819 (I985636,I1049522,I1049528);
nor I_57820 (I985653,I985636,I1049540);
and I_57821 (I985670,I985653,I985557);
DFFARX1 I_57822 (I985670,I2683,I985342,I985328,);
nor I_57823 (I985325,I985636,I985492);
or I_57824 (I985322,I985574,I985636);
nor I_57825 (I985729,I1049522,I1049519);
DFFARX1 I_57826 (I985729,I2683,I985342,I985755,);
not I_57827 (I985763,I985755);
nand I_57828 (I985780,I985763,I985441);
nor I_57829 (I985797,I985780,I1049540);
DFFARX1 I_57830 (I985797,I2683,I985342,I985310,);
nor I_57831 (I985828,I985763,I985492);
nor I_57832 (I985319,I985636,I985828);
not I_57833 (I985886,I2690);
DFFARX1 I_57834 (I865212,I2683,I985886,I985912,);
nand I_57835 (I985920,I985912,I865191);
DFFARX1 I_57836 (I865188,I2683,I985886,I985946,);
DFFARX1 I_57837 (I985946,I2683,I985886,I985963,);
not I_57838 (I985878,I985963);
not I_57839 (I985985,I865200);
nor I_57840 (I986002,I865200,I865209);
not I_57841 (I986019,I865197);
nand I_57842 (I986036,I985985,I986019);
nor I_57843 (I986053,I865197,I865200);
and I_57844 (I985857,I986053,I985920);
not I_57845 (I986084,I865206);
nand I_57846 (I986101,I986084,I865203);
nor I_57847 (I986118,I865206,I865188);
not I_57848 (I986135,I986118);
nand I_57849 (I985860,I986002,I986135);
DFFARX1 I_57850 (I986118,I2683,I985886,I985875,);
nor I_57851 (I986180,I865191,I865197);
nor I_57852 (I986197,I986180,I865209);
and I_57853 (I986214,I986197,I986101);
DFFARX1 I_57854 (I986214,I2683,I985886,I985872,);
nor I_57855 (I985869,I986180,I986036);
or I_57856 (I985866,I986118,I986180);
nor I_57857 (I986273,I865191,I865194);
DFFARX1 I_57858 (I986273,I2683,I985886,I986299,);
not I_57859 (I986307,I986299);
nand I_57860 (I986324,I986307,I985985);
nor I_57861 (I986341,I986324,I865209);
DFFARX1 I_57862 (I986341,I2683,I985886,I985854,);
nor I_57863 (I986372,I986307,I986036);
nor I_57864 (I985863,I986180,I986372);
not I_57865 (I986430,I2690);
DFFARX1 I_57866 (I923012,I2683,I986430,I986456,);
nand I_57867 (I986464,I986456,I922991);
DFFARX1 I_57868 (I922988,I2683,I986430,I986490,);
DFFARX1 I_57869 (I986490,I2683,I986430,I986507,);
not I_57870 (I986422,I986507);
not I_57871 (I986529,I923000);
nor I_57872 (I986546,I923000,I923009);
not I_57873 (I986563,I922997);
nand I_57874 (I986580,I986529,I986563);
nor I_57875 (I986597,I922997,I923000);
and I_57876 (I986401,I986597,I986464);
not I_57877 (I986628,I923006);
nand I_57878 (I986645,I986628,I923003);
nor I_57879 (I986662,I923006,I922988);
not I_57880 (I986679,I986662);
nand I_57881 (I986404,I986546,I986679);
DFFARX1 I_57882 (I986662,I2683,I986430,I986419,);
nor I_57883 (I986724,I922991,I922997);
nor I_57884 (I986741,I986724,I923009);
and I_57885 (I986758,I986741,I986645);
DFFARX1 I_57886 (I986758,I2683,I986430,I986416,);
nor I_57887 (I986413,I986724,I986580);
or I_57888 (I986410,I986662,I986724);
nor I_57889 (I986817,I922991,I922994);
DFFARX1 I_57890 (I986817,I2683,I986430,I986843,);
not I_57891 (I986851,I986843);
nand I_57892 (I986868,I986851,I986529);
nor I_57893 (I986885,I986868,I923009);
DFFARX1 I_57894 (I986885,I2683,I986430,I986398,);
nor I_57895 (I986916,I986851,I986580);
nor I_57896 (I986407,I986724,I986916);
not I_57897 (I986974,I2690);
DFFARX1 I_57898 (I376394,I2683,I986974,I987000,);
nand I_57899 (I987008,I987000,I376391);
DFFARX1 I_57900 (I376370,I2683,I986974,I987034,);
DFFARX1 I_57901 (I987034,I2683,I986974,I987051,);
not I_57902 (I986966,I987051);
not I_57903 (I987073,I376385);
nor I_57904 (I987090,I376385,I376388);
not I_57905 (I987107,I376379);
nand I_57906 (I987124,I987073,I987107);
nor I_57907 (I987141,I376379,I376385);
and I_57908 (I986945,I987141,I987008);
not I_57909 (I987172,I376376);
nand I_57910 (I987189,I987172,I376397);
nor I_57911 (I987206,I376376,I376373);
not I_57912 (I987223,I987206);
nand I_57913 (I986948,I987090,I987223);
DFFARX1 I_57914 (I987206,I2683,I986974,I986963,);
nor I_57915 (I987268,I376382,I376379);
nor I_57916 (I987285,I987268,I376388);
and I_57917 (I987302,I987285,I987189);
DFFARX1 I_57918 (I987302,I2683,I986974,I986960,);
nor I_57919 (I986957,I987268,I987124);
or I_57920 (I986954,I987206,I987268);
nor I_57921 (I987361,I376382,I376370);
DFFARX1 I_57922 (I987361,I2683,I986974,I987387,);
not I_57923 (I987395,I987387);
nand I_57924 (I987412,I987395,I987073);
nor I_57925 (I987429,I987412,I376388);
DFFARX1 I_57926 (I987429,I2683,I986974,I986942,);
nor I_57927 (I987460,I987395,I987124);
nor I_57928 (I986951,I987268,I987460);
not I_57929 (I987518,I2690);
DFFARX1 I_57930 (I265406,I2683,I987518,I987544,);
nand I_57931 (I987552,I987544,I265409);
DFFARX1 I_57932 (I265403,I2683,I987518,I987578,);
DFFARX1 I_57933 (I987578,I2683,I987518,I987595,);
not I_57934 (I987510,I987595);
not I_57935 (I987617,I265412);
nor I_57936 (I987634,I265412,I265397);
not I_57937 (I987651,I265421);
nand I_57938 (I987668,I987617,I987651);
nor I_57939 (I987685,I265421,I265412);
and I_57940 (I987489,I987685,I987552);
not I_57941 (I987716,I265400);
nand I_57942 (I987733,I987716,I265418);
nor I_57943 (I987750,I265400,I265394);
not I_57944 (I987767,I987750);
nand I_57945 (I987492,I987634,I987767);
DFFARX1 I_57946 (I987750,I2683,I987518,I987507,);
nor I_57947 (I987812,I265415,I265421);
nor I_57948 (I987829,I987812,I265397);
and I_57949 (I987846,I987829,I987733);
DFFARX1 I_57950 (I987846,I2683,I987518,I987504,);
nor I_57951 (I987501,I987812,I987668);
or I_57952 (I987498,I987750,I987812);
nor I_57953 (I987905,I265415,I265394);
DFFARX1 I_57954 (I987905,I2683,I987518,I987931,);
not I_57955 (I987939,I987931);
nand I_57956 (I987956,I987939,I987617);
nor I_57957 (I987973,I987956,I265397);
DFFARX1 I_57958 (I987973,I2683,I987518,I987486,);
nor I_57959 (I988004,I987939,I987668);
nor I_57960 (I987495,I987812,I988004);
not I_57961 (I988062,I2690);
DFFARX1 I_57962 (I494269,I2683,I988062,I988088,);
nand I_57963 (I988096,I988088,I494257);
DFFARX1 I_57964 (I494263,I2683,I988062,I988122,);
DFFARX1 I_57965 (I988122,I2683,I988062,I988139,);
not I_57966 (I988054,I988139);
not I_57967 (I988161,I494248);
nor I_57968 (I988178,I494248,I494260);
not I_57969 (I988195,I494251);
nand I_57970 (I988212,I988161,I988195);
nor I_57971 (I988229,I494251,I494248);
and I_57972 (I988033,I988229,I988096);
not I_57973 (I988260,I494266);
nand I_57974 (I988277,I988260,I494248);
nor I_57975 (I988294,I494266,I494272);
not I_57976 (I988311,I988294);
nand I_57977 (I988036,I988178,I988311);
DFFARX1 I_57978 (I988294,I2683,I988062,I988051,);
nor I_57979 (I988356,I494254,I494251);
nor I_57980 (I988373,I988356,I494260);
and I_57981 (I988390,I988373,I988277);
DFFARX1 I_57982 (I988390,I2683,I988062,I988048,);
nor I_57983 (I988045,I988356,I988212);
or I_57984 (I988042,I988294,I988356);
nor I_57985 (I988449,I494254,I494251);
DFFARX1 I_57986 (I988449,I2683,I988062,I988475,);
not I_57987 (I988483,I988475);
nand I_57988 (I988500,I988483,I988161);
nor I_57989 (I988517,I988500,I494260);
DFFARX1 I_57990 (I988517,I2683,I988062,I988030,);
nor I_57991 (I988548,I988483,I988212);
nor I_57992 (I988039,I988356,I988548);
not I_57993 (I988606,I2690);
DFFARX1 I_57994 (I1048948,I2683,I988606,I988632,);
nand I_57995 (I988640,I988632,I1048939);
not I_57996 (I988657,I988640);
DFFARX1 I_57997 (I1048924,I2683,I988606,I988683,);
not I_57998 (I988691,I988683);
not I_57999 (I988708,I1048927);
or I_58000 (I988725,I1048936,I1048927);
nor I_58001 (I988742,I1048936,I1048927);
or I_58002 (I988759,I1048933,I1048936);
DFFARX1 I_58003 (I988759,I2683,I988606,I988598,);
not I_58004 (I988790,I1048945);
nand I_58005 (I988807,I988790,I1048924);
nand I_58006 (I988824,I988708,I988807);
and I_58007 (I988577,I988691,I988824);
nor I_58008 (I988855,I1048945,I1048930);
and I_58009 (I988872,I988691,I988855);
nor I_58010 (I988583,I988657,I988872);
DFFARX1 I_58011 (I988855,I2683,I988606,I988912,);
not I_58012 (I988920,I988912);
nor I_58013 (I988592,I988691,I988920);
or I_58014 (I988951,I988759,I1048951);
nor I_58015 (I988968,I1048951,I1048933);
nand I_58016 (I988985,I988824,I988968);
nand I_58017 (I989002,I988951,I988985);
DFFARX1 I_58018 (I989002,I2683,I988606,I988595,);
nor I_58019 (I989033,I988968,I988725);
DFFARX1 I_58020 (I989033,I2683,I988606,I988574,);
nor I_58021 (I989064,I1048951,I1048942);
DFFARX1 I_58022 (I989064,I2683,I988606,I989090,);
DFFARX1 I_58023 (I989090,I2683,I988606,I988589,);
not I_58024 (I989112,I989090);
nand I_58025 (I988586,I989112,I988640);
nand I_58026 (I988580,I989112,I988742);
not I_58027 (I989184,I2690);
DFFARX1 I_58028 (I742607,I2683,I989184,I989210,);
nand I_58029 (I989218,I989210,I742628);
not I_58030 (I989235,I989218);
DFFARX1 I_58031 (I742601,I2683,I989184,I989261,);
not I_58032 (I989269,I989261);
not I_58033 (I989286,I742622);
or I_58034 (I989303,I742613,I742622);
nor I_58035 (I989320,I742613,I742622);
or I_58036 (I989337,I742616,I742613);
DFFARX1 I_58037 (I989337,I2683,I989184,I989176,);
not I_58038 (I989368,I742604);
nand I_58039 (I989385,I989368,I742619);
nand I_58040 (I989402,I989286,I989385);
and I_58041 (I989155,I989269,I989402);
nor I_58042 (I989433,I742604,I742601);
and I_58043 (I989450,I989269,I989433);
nor I_58044 (I989161,I989235,I989450);
DFFARX1 I_58045 (I989433,I2683,I989184,I989490,);
not I_58046 (I989498,I989490);
nor I_58047 (I989170,I989269,I989498);
or I_58048 (I989529,I989337,I742625);
nor I_58049 (I989546,I742625,I742616);
nand I_58050 (I989563,I989402,I989546);
nand I_58051 (I989580,I989529,I989563);
DFFARX1 I_58052 (I989580,I2683,I989184,I989173,);
nor I_58053 (I989611,I989546,I989303);
DFFARX1 I_58054 (I989611,I2683,I989184,I989152,);
nor I_58055 (I989642,I742625,I742610);
DFFARX1 I_58056 (I989642,I2683,I989184,I989668,);
DFFARX1 I_58057 (I989668,I2683,I989184,I989167,);
not I_58058 (I989690,I989668);
nand I_58059 (I989164,I989690,I989218);
nand I_58060 (I989158,I989690,I989320);
not I_58061 (I989762,I2690);
DFFARX1 I_58062 (I364405,I2683,I989762,I989788,);
nand I_58063 (I989796,I989788,I364414);
not I_58064 (I989813,I989796);
DFFARX1 I_58065 (I364402,I2683,I989762,I989839,);
not I_58066 (I989847,I989839);
not I_58067 (I989864,I364408);
or I_58068 (I989881,I364402,I364408);
nor I_58069 (I989898,I364402,I364408);
or I_58070 (I989915,I364417,I364402);
DFFARX1 I_58071 (I989915,I2683,I989762,I989754,);
not I_58072 (I989946,I364411);
nand I_58073 (I989963,I989946,I364426);
nand I_58074 (I989980,I989864,I989963);
and I_58075 (I989733,I989847,I989980);
nor I_58076 (I990011,I364411,I364429);
and I_58077 (I990028,I989847,I990011);
nor I_58078 (I989739,I989813,I990028);
DFFARX1 I_58079 (I990011,I2683,I989762,I990068,);
not I_58080 (I990076,I990068);
nor I_58081 (I989748,I989847,I990076);
or I_58082 (I990107,I989915,I364420);
nor I_58083 (I990124,I364420,I364417);
nand I_58084 (I990141,I989980,I990124);
nand I_58085 (I990158,I990107,I990141);
DFFARX1 I_58086 (I990158,I2683,I989762,I989751,);
nor I_58087 (I990189,I990124,I989881);
DFFARX1 I_58088 (I990189,I2683,I989762,I989730,);
nor I_58089 (I990220,I364420,I364423);
DFFARX1 I_58090 (I990220,I2683,I989762,I990246,);
DFFARX1 I_58091 (I990246,I2683,I989762,I989745,);
not I_58092 (I990268,I990246);
nand I_58093 (I989742,I990268,I989796);
nand I_58094 (I989736,I990268,I989898);
not I_58095 (I990340,I2690);
DFFARX1 I_58096 (I927630,I2683,I990340,I990366,);
nand I_58097 (I990374,I990366,I927615);
not I_58098 (I990391,I990374);
DFFARX1 I_58099 (I927618,I2683,I990340,I990417,);
not I_58100 (I990425,I990417);
not I_58101 (I990442,I927633);
or I_58102 (I990459,I927636,I927633);
nor I_58103 (I990476,I927636,I927633);
or I_58104 (I990493,I927612,I927636);
DFFARX1 I_58105 (I990493,I2683,I990340,I990332,);
not I_58106 (I990524,I927624);
nand I_58107 (I990541,I990524,I927627);
nand I_58108 (I990558,I990442,I990541);
and I_58109 (I990311,I990425,I990558);
nor I_58110 (I990589,I927624,I927621);
and I_58111 (I990606,I990425,I990589);
nor I_58112 (I990317,I990391,I990606);
DFFARX1 I_58113 (I990589,I2683,I990340,I990646,);
not I_58114 (I990654,I990646);
nor I_58115 (I990326,I990425,I990654);
or I_58116 (I990685,I990493,I927612);
nor I_58117 (I990702,I927612,I927612);
nand I_58118 (I990719,I990558,I990702);
nand I_58119 (I990736,I990685,I990719);
DFFARX1 I_58120 (I990736,I2683,I990340,I990329,);
nor I_58121 (I990767,I990702,I990459);
DFFARX1 I_58122 (I990767,I2683,I990340,I990308,);
nor I_58123 (I990798,I927612,I927615);
DFFARX1 I_58124 (I990798,I2683,I990340,I990824,);
DFFARX1 I_58125 (I990824,I2683,I990340,I990323,);
not I_58126 (I990846,I990824);
nand I_58127 (I990320,I990846,I990374);
nand I_58128 (I990314,I990846,I990476);
not I_58129 (I990918,I2690);
DFFARX1 I_58130 (I116455,I2683,I990918,I990944,);
nand I_58131 (I990952,I990944,I116464);
not I_58132 (I990969,I990952);
DFFARX1 I_58133 (I116446,I2683,I990918,I990995,);
not I_58134 (I991003,I990995);
not I_58135 (I991020,I116452);
or I_58136 (I991037,I116461,I116452);
nor I_58137 (I991054,I116461,I116452);
or I_58138 (I991071,I116449,I116461);
DFFARX1 I_58139 (I991071,I2683,I990918,I990910,);
not I_58140 (I991102,I116467);
nand I_58141 (I991119,I991102,I116440);
nand I_58142 (I991136,I991020,I991119);
and I_58143 (I990889,I991003,I991136);
nor I_58144 (I991167,I116467,I116443);
and I_58145 (I991184,I991003,I991167);
nor I_58146 (I990895,I990969,I991184);
DFFARX1 I_58147 (I991167,I2683,I990918,I991224,);
not I_58148 (I991232,I991224);
nor I_58149 (I990904,I991003,I991232);
or I_58150 (I991263,I991071,I116458);
nor I_58151 (I991280,I116458,I116449);
nand I_58152 (I991297,I991136,I991280);
nand I_58153 (I991314,I991263,I991297);
DFFARX1 I_58154 (I991314,I2683,I990918,I990907,);
nor I_58155 (I991345,I991280,I991037);
DFFARX1 I_58156 (I991345,I2683,I990918,I990886,);
nor I_58157 (I991376,I116458,I116440);
DFFARX1 I_58158 (I991376,I2683,I990918,I991402,);
DFFARX1 I_58159 (I991402,I2683,I990918,I990901,);
not I_58160 (I991424,I991402);
nand I_58161 (I990898,I991424,I990952);
nand I_58162 (I990892,I991424,I991054);
not I_58163 (I991496,I2690);
DFFARX1 I_58164 (I512166,I2683,I991496,I991522,);
nand I_58165 (I991530,I991522,I512169);
not I_58166 (I991547,I991530);
DFFARX1 I_58167 (I512181,I2683,I991496,I991573,);
not I_58168 (I991581,I991573);
not I_58169 (I991598,I512166);
or I_58170 (I991615,I512175,I512166);
nor I_58171 (I991632,I512175,I512166);
or I_58172 (I991649,I512184,I512175);
DFFARX1 I_58173 (I991649,I2683,I991496,I991488,);
not I_58174 (I991680,I512187);
nand I_58175 (I991697,I991680,I512169);
nand I_58176 (I991714,I991598,I991697);
and I_58177 (I991467,I991581,I991714);
nor I_58178 (I991745,I512187,I512172);
and I_58179 (I991762,I991581,I991745);
nor I_58180 (I991473,I991547,I991762);
DFFARX1 I_58181 (I991745,I2683,I991496,I991802,);
not I_58182 (I991810,I991802);
nor I_58183 (I991482,I991581,I991810);
or I_58184 (I991841,I991649,I512178);
nor I_58185 (I991858,I512178,I512184);
nand I_58186 (I991875,I991714,I991858);
nand I_58187 (I991892,I991841,I991875);
DFFARX1 I_58188 (I991892,I2683,I991496,I991485,);
nor I_58189 (I991923,I991858,I991615);
DFFARX1 I_58190 (I991923,I2683,I991496,I991464,);
nor I_58191 (I991954,I512178,I512190);
DFFARX1 I_58192 (I991954,I2683,I991496,I991980,);
DFFARX1 I_58193 (I991980,I2683,I991496,I991479,);
not I_58194 (I992002,I991980);
nand I_58195 (I991476,I992002,I991530);
nand I_58196 (I991470,I992002,I991632);
not I_58197 (I992074,I2690);
DFFARX1 I_58198 (I279102,I2683,I992074,I992100,);
nand I_58199 (I992108,I992100,I279123);
not I_58200 (I992125,I992108);
DFFARX1 I_58201 (I279117,I2683,I992074,I992151,);
not I_58202 (I992159,I992151);
not I_58203 (I992176,I279105);
or I_58204 (I992193,I279120,I279105);
nor I_58205 (I992210,I279120,I279105);
or I_58206 (I992227,I279111,I279120);
DFFARX1 I_58207 (I992227,I2683,I992074,I992066,);
not I_58208 (I992258,I279099);
nand I_58209 (I992275,I992258,I279096);
nand I_58210 (I992292,I992176,I992275);
and I_58211 (I992045,I992159,I992292);
nor I_58212 (I992323,I279099,I279108);
and I_58213 (I992340,I992159,I992323);
nor I_58214 (I992051,I992125,I992340);
DFFARX1 I_58215 (I992323,I2683,I992074,I992380,);
not I_58216 (I992388,I992380);
nor I_58217 (I992060,I992159,I992388);
or I_58218 (I992419,I992227,I279114);
nor I_58219 (I992436,I279114,I279111);
nand I_58220 (I992453,I992292,I992436);
nand I_58221 (I992470,I992419,I992453);
DFFARX1 I_58222 (I992470,I2683,I992074,I992063,);
nor I_58223 (I992501,I992436,I992193);
DFFARX1 I_58224 (I992501,I2683,I992074,I992042,);
nor I_58225 (I992532,I279114,I279096);
DFFARX1 I_58226 (I992532,I2683,I992074,I992558,);
DFFARX1 I_58227 (I992558,I2683,I992074,I992057,);
not I_58228 (I992580,I992558);
nand I_58229 (I992054,I992580,I992108);
nand I_58230 (I992048,I992580,I992210);
not I_58231 (I992652,I2690);
DFFARX1 I_58232 (I604068,I2683,I992652,I992678,);
nand I_58233 (I992686,I992678,I604071);
not I_58234 (I992703,I992686);
DFFARX1 I_58235 (I604083,I2683,I992652,I992729,);
not I_58236 (I992737,I992729);
not I_58237 (I992754,I604068);
or I_58238 (I992771,I604077,I604068);
nor I_58239 (I992788,I604077,I604068);
or I_58240 (I992805,I604086,I604077);
DFFARX1 I_58241 (I992805,I2683,I992652,I992644,);
not I_58242 (I992836,I604089);
nand I_58243 (I992853,I992836,I604071);
nand I_58244 (I992870,I992754,I992853);
and I_58245 (I992623,I992737,I992870);
nor I_58246 (I992901,I604089,I604074);
and I_58247 (I992918,I992737,I992901);
nor I_58248 (I992629,I992703,I992918);
DFFARX1 I_58249 (I992901,I2683,I992652,I992958,);
not I_58250 (I992966,I992958);
nor I_58251 (I992638,I992737,I992966);
or I_58252 (I992997,I992805,I604080);
nor I_58253 (I993014,I604080,I604086);
nand I_58254 (I993031,I992870,I993014);
nand I_58255 (I993048,I992997,I993031);
DFFARX1 I_58256 (I993048,I2683,I992652,I992641,);
nor I_58257 (I993079,I993014,I992771);
DFFARX1 I_58258 (I993079,I2683,I992652,I992620,);
nor I_58259 (I993110,I604080,I604092);
DFFARX1 I_58260 (I993110,I2683,I992652,I993136,);
DFFARX1 I_58261 (I993136,I2683,I992652,I992635,);
not I_58262 (I993158,I993136);
nand I_58263 (I992632,I993158,I992686);
nand I_58264 (I992626,I993158,I992788);
not I_58265 (I993230,I2690);
DFFARX1 I_58266 (I101220,I2683,I993230,I993256,);
nand I_58267 (I993264,I993256,I101211);
not I_58268 (I993281,I993264);
DFFARX1 I_58269 (I101208,I2683,I993230,I993307,);
not I_58270 (I993315,I993307);
not I_58271 (I993332,I101217);
or I_58272 (I993349,I101208,I101217);
nor I_58273 (I993366,I101208,I101217);
or I_58274 (I993383,I101214,I101208);
DFFARX1 I_58275 (I993383,I2683,I993230,I993222,);
not I_58276 (I993414,I101223);
nand I_58277 (I993431,I993414,I101232);
nand I_58278 (I993448,I993332,I993431);
and I_58279 (I993201,I993315,I993448);
nor I_58280 (I993479,I101223,I101226);
and I_58281 (I993496,I993315,I993479);
nor I_58282 (I993207,I993281,I993496);
DFFARX1 I_58283 (I993479,I2683,I993230,I993536,);
not I_58284 (I993544,I993536);
nor I_58285 (I993216,I993315,I993544);
or I_58286 (I993575,I993383,I101211);
nor I_58287 (I993592,I101211,I101214);
nand I_58288 (I993609,I993448,I993592);
nand I_58289 (I993626,I993575,I993609);
DFFARX1 I_58290 (I993626,I2683,I993230,I993219,);
nor I_58291 (I993657,I993592,I993349);
DFFARX1 I_58292 (I993657,I2683,I993230,I993198,);
nor I_58293 (I993688,I101211,I101229);
DFFARX1 I_58294 (I993688,I2683,I993230,I993714,);
DFFARX1 I_58295 (I993714,I2683,I993230,I993213,);
not I_58296 (I993736,I993714);
nand I_58297 (I993210,I993736,I993264);
nand I_58298 (I993204,I993736,I993366);
not I_58299 (I993808,I2690);
DFFARX1 I_58300 (I392693,I2683,I993808,I993834,);
nand I_58301 (I993842,I993834,I392702);
not I_58302 (I993859,I993842);
DFFARX1 I_58303 (I392690,I2683,I993808,I993885,);
not I_58304 (I993893,I993885);
not I_58305 (I993910,I392696);
or I_58306 (I993927,I392690,I392696);
nor I_58307 (I993944,I392690,I392696);
or I_58308 (I993961,I392705,I392690);
DFFARX1 I_58309 (I993961,I2683,I993808,I993800,);
not I_58310 (I993992,I392699);
nand I_58311 (I994009,I993992,I392714);
nand I_58312 (I994026,I993910,I994009);
and I_58313 (I993779,I993893,I994026);
nor I_58314 (I994057,I392699,I392717);
and I_58315 (I994074,I993893,I994057);
nor I_58316 (I993785,I993859,I994074);
DFFARX1 I_58317 (I994057,I2683,I993808,I994114,);
not I_58318 (I994122,I994114);
nor I_58319 (I993794,I993893,I994122);
or I_58320 (I994153,I993961,I392708);
nor I_58321 (I994170,I392708,I392705);
nand I_58322 (I994187,I994026,I994170);
nand I_58323 (I994204,I994153,I994187);
DFFARX1 I_58324 (I994204,I2683,I993808,I993797,);
nor I_58325 (I994235,I994170,I993927);
DFFARX1 I_58326 (I994235,I2683,I993808,I993776,);
nor I_58327 (I994266,I392708,I392711);
DFFARX1 I_58328 (I994266,I2683,I993808,I994292,);
DFFARX1 I_58329 (I994292,I2683,I993808,I993791,);
not I_58330 (I994314,I994292);
nand I_58331 (I993788,I994314,I993842);
nand I_58332 (I993782,I994314,I993944);
not I_58333 (I994386,I2690);
DFFARX1 I_58334 (I1069773,I2683,I994386,I994412,);
nand I_58335 (I994420,I994412,I1069764);
not I_58336 (I994437,I994420);
DFFARX1 I_58337 (I1069749,I2683,I994386,I994463,);
not I_58338 (I994471,I994463);
not I_58339 (I994488,I1069752);
or I_58340 (I994505,I1069761,I1069752);
nor I_58341 (I994522,I1069761,I1069752);
or I_58342 (I994539,I1069758,I1069761);
DFFARX1 I_58343 (I994539,I2683,I994386,I994378,);
not I_58344 (I994570,I1069770);
nand I_58345 (I994587,I994570,I1069749);
nand I_58346 (I994604,I994488,I994587);
and I_58347 (I994357,I994471,I994604);
nor I_58348 (I994635,I1069770,I1069755);
and I_58349 (I994652,I994471,I994635);
nor I_58350 (I994363,I994437,I994652);
DFFARX1 I_58351 (I994635,I2683,I994386,I994692,);
not I_58352 (I994700,I994692);
nor I_58353 (I994372,I994471,I994700);
or I_58354 (I994731,I994539,I1069776);
nor I_58355 (I994748,I1069776,I1069758);
nand I_58356 (I994765,I994604,I994748);
nand I_58357 (I994782,I994731,I994765);
DFFARX1 I_58358 (I994782,I2683,I994386,I994375,);
nor I_58359 (I994813,I994748,I994505);
DFFARX1 I_58360 (I994813,I2683,I994386,I994354,);
nor I_58361 (I994844,I1069776,I1069767);
DFFARX1 I_58362 (I994844,I2683,I994386,I994870,);
DFFARX1 I_58363 (I994870,I2683,I994386,I994369,);
not I_58364 (I994892,I994870);
nand I_58365 (I994366,I994892,I994420);
nand I_58366 (I994360,I994892,I994522);
not I_58367 (I994964,I2690);
DFFARX1 I_58368 (I907400,I2683,I994964,I994990,);
nand I_58369 (I994998,I994990,I907385);
not I_58370 (I995015,I994998);
DFFARX1 I_58371 (I907388,I2683,I994964,I995041,);
not I_58372 (I995049,I995041);
not I_58373 (I995066,I907403);
or I_58374 (I995083,I907406,I907403);
nor I_58375 (I995100,I907406,I907403);
or I_58376 (I995117,I907382,I907406);
DFFARX1 I_58377 (I995117,I2683,I994964,I994956,);
not I_58378 (I995148,I907394);
nand I_58379 (I995165,I995148,I907397);
nand I_58380 (I995182,I995066,I995165);
and I_58381 (I994935,I995049,I995182);
nor I_58382 (I995213,I907394,I907391);
and I_58383 (I995230,I995049,I995213);
nor I_58384 (I994941,I995015,I995230);
DFFARX1 I_58385 (I995213,I2683,I994964,I995270,);
not I_58386 (I995278,I995270);
nor I_58387 (I994950,I995049,I995278);
or I_58388 (I995309,I995117,I907382);
nor I_58389 (I995326,I907382,I907382);
nand I_58390 (I995343,I995182,I995326);
nand I_58391 (I995360,I995309,I995343);
DFFARX1 I_58392 (I995360,I2683,I994964,I994953,);
nor I_58393 (I995391,I995326,I995083);
DFFARX1 I_58394 (I995391,I2683,I994964,I994932,);
nor I_58395 (I995422,I907382,I907385);
DFFARX1 I_58396 (I995422,I2683,I994964,I995448,);
DFFARX1 I_58397 (I995448,I2683,I994964,I994947,);
not I_58398 (I995470,I995448);
nand I_58399 (I994944,I995470,I994998);
nand I_58400 (I994938,I995470,I995100);
not I_58401 (I995542,I2690);
DFFARX1 I_58402 (I734855,I2683,I995542,I995568,);
nand I_58403 (I995576,I995568,I734876);
not I_58404 (I995593,I995576);
DFFARX1 I_58405 (I734849,I2683,I995542,I995619,);
not I_58406 (I995627,I995619);
not I_58407 (I995644,I734870);
or I_58408 (I995661,I734861,I734870);
nor I_58409 (I995678,I734861,I734870);
or I_58410 (I995695,I734864,I734861);
DFFARX1 I_58411 (I995695,I2683,I995542,I995534,);
not I_58412 (I995726,I734852);
nand I_58413 (I995743,I995726,I734867);
nand I_58414 (I995760,I995644,I995743);
and I_58415 (I995513,I995627,I995760);
nor I_58416 (I995791,I734852,I734849);
and I_58417 (I995808,I995627,I995791);
nor I_58418 (I995519,I995593,I995808);
DFFARX1 I_58419 (I995791,I2683,I995542,I995848,);
not I_58420 (I995856,I995848);
nor I_58421 (I995528,I995627,I995856);
or I_58422 (I995887,I995695,I734873);
nor I_58423 (I995904,I734873,I734864);
nand I_58424 (I995921,I995760,I995904);
nand I_58425 (I995938,I995887,I995921);
DFFARX1 I_58426 (I995938,I2683,I995542,I995531,);
nor I_58427 (I995969,I995904,I995661);
DFFARX1 I_58428 (I995969,I2683,I995542,I995510,);
nor I_58429 (I996000,I734873,I734858);
DFFARX1 I_58430 (I996000,I2683,I995542,I996026,);
DFFARX1 I_58431 (I996026,I2683,I995542,I995525,);
not I_58432 (I996048,I996026);
nand I_58433 (I995522,I996048,I995576);
nand I_58434 (I995516,I996048,I995678);
not I_58435 (I996120,I2690);
DFFARX1 I_58436 (I751005,I2683,I996120,I996146,);
nand I_58437 (I996154,I996146,I751026);
not I_58438 (I996171,I996154);
DFFARX1 I_58439 (I750999,I2683,I996120,I996197,);
not I_58440 (I996205,I996197);
not I_58441 (I996222,I751020);
or I_58442 (I996239,I751011,I751020);
nor I_58443 (I996256,I751011,I751020);
or I_58444 (I996273,I751014,I751011);
DFFARX1 I_58445 (I996273,I2683,I996120,I996112,);
not I_58446 (I996304,I751002);
nand I_58447 (I996321,I996304,I751017);
nand I_58448 (I996338,I996222,I996321);
and I_58449 (I996091,I996205,I996338);
nor I_58450 (I996369,I751002,I750999);
and I_58451 (I996386,I996205,I996369);
nor I_58452 (I996097,I996171,I996386);
DFFARX1 I_58453 (I996369,I2683,I996120,I996426,);
not I_58454 (I996434,I996426);
nor I_58455 (I996106,I996205,I996434);
or I_58456 (I996465,I996273,I751023);
nor I_58457 (I996482,I751023,I751014);
nand I_58458 (I996499,I996338,I996482);
nand I_58459 (I996516,I996465,I996499);
DFFARX1 I_58460 (I996516,I2683,I996120,I996109,);
nor I_58461 (I996547,I996482,I996239);
DFFARX1 I_58462 (I996547,I2683,I996120,I996088,);
nor I_58463 (I996578,I751023,I751008);
DFFARX1 I_58464 (I996578,I2683,I996120,I996604,);
DFFARX1 I_58465 (I996604,I2683,I996120,I996103,);
not I_58466 (I996626,I996604);
nand I_58467 (I996100,I996626,I996154);
nand I_58468 (I996094,I996626,I996256);
not I_58469 (I996698,I2690);
DFFARX1 I_58470 (I452057,I2683,I996698,I996724,);
nand I_58471 (I996732,I996724,I452072);
not I_58472 (I996749,I996732);
DFFARX1 I_58473 (I452054,I2683,I996698,I996775,);
not I_58474 (I996783,I996775);
not I_58475 (I996800,I452063);
or I_58476 (I996817,I452057,I452063);
nor I_58477 (I996834,I452057,I452063);
or I_58478 (I996851,I452054,I452057);
DFFARX1 I_58479 (I996851,I2683,I996698,I996690,);
not I_58480 (I996882,I452075);
nand I_58481 (I996899,I996882,I452078);
nand I_58482 (I996916,I996800,I996899);
and I_58483 (I996669,I996783,I996916);
nor I_58484 (I996947,I452075,I452060);
and I_58485 (I996964,I996783,I996947);
nor I_58486 (I996675,I996749,I996964);
DFFARX1 I_58487 (I996947,I2683,I996698,I997004,);
not I_58488 (I997012,I997004);
nor I_58489 (I996684,I996783,I997012);
or I_58490 (I997043,I996851,I452066);
nor I_58491 (I997060,I452066,I452054);
nand I_58492 (I997077,I996916,I997060);
nand I_58493 (I997094,I997043,I997077);
DFFARX1 I_58494 (I997094,I2683,I996698,I996687,);
nor I_58495 (I997125,I997060,I996817);
DFFARX1 I_58496 (I997125,I2683,I996698,I996666,);
nor I_58497 (I997156,I452066,I452069);
DFFARX1 I_58498 (I997156,I2683,I996698,I997182,);
DFFARX1 I_58499 (I997182,I2683,I996698,I996681,);
not I_58500 (I997204,I997182);
nand I_58501 (I996678,I997204,I996732);
nand I_58502 (I996672,I997204,I996834);
not I_58503 (I997276,I2690);
DFFARX1 I_58504 (I756173,I2683,I997276,I997302,);
nand I_58505 (I997310,I997302,I756194);
not I_58506 (I997327,I997310);
DFFARX1 I_58507 (I756167,I2683,I997276,I997353,);
not I_58508 (I997361,I997353);
not I_58509 (I997378,I756188);
or I_58510 (I997395,I756179,I756188);
nor I_58511 (I997412,I756179,I756188);
or I_58512 (I997429,I756182,I756179);
DFFARX1 I_58513 (I997429,I2683,I997276,I997268,);
not I_58514 (I997460,I756170);
nand I_58515 (I997477,I997460,I756185);
nand I_58516 (I997494,I997378,I997477);
and I_58517 (I997247,I997361,I997494);
nor I_58518 (I997525,I756170,I756167);
and I_58519 (I997542,I997361,I997525);
nor I_58520 (I997253,I997327,I997542);
DFFARX1 I_58521 (I997525,I2683,I997276,I997582,);
not I_58522 (I997590,I997582);
nor I_58523 (I997262,I997361,I997590);
or I_58524 (I997621,I997429,I756191);
nor I_58525 (I997638,I756191,I756182);
nand I_58526 (I997655,I997494,I997638);
nand I_58527 (I997672,I997621,I997655);
DFFARX1 I_58528 (I997672,I2683,I997276,I997265,);
nor I_58529 (I997703,I997638,I997395);
DFFARX1 I_58530 (I997703,I2683,I997276,I997244,);
nor I_58531 (I997734,I756191,I756176);
DFFARX1 I_58532 (I997734,I2683,I997276,I997760,);
DFFARX1 I_58533 (I997760,I2683,I997276,I997259,);
not I_58534 (I997782,I997760);
nand I_58535 (I997256,I997782,I997310);
nand I_58536 (I997250,I997782,I997412);
not I_58537 (I997854,I2690);
DFFARX1 I_58538 (I782659,I2683,I997854,I997880,);
nand I_58539 (I997888,I997880,I782680);
not I_58540 (I997905,I997888);
DFFARX1 I_58541 (I782653,I2683,I997854,I997931,);
not I_58542 (I997939,I997931);
not I_58543 (I997956,I782674);
or I_58544 (I997973,I782665,I782674);
nor I_58545 (I997990,I782665,I782674);
or I_58546 (I998007,I782668,I782665);
DFFARX1 I_58547 (I998007,I2683,I997854,I997846,);
not I_58548 (I998038,I782656);
nand I_58549 (I998055,I998038,I782671);
nand I_58550 (I998072,I997956,I998055);
and I_58551 (I997825,I997939,I998072);
nor I_58552 (I998103,I782656,I782653);
and I_58553 (I998120,I997939,I998103);
nor I_58554 (I997831,I997905,I998120);
DFFARX1 I_58555 (I998103,I2683,I997854,I998160,);
not I_58556 (I998168,I998160);
nor I_58557 (I997840,I997939,I998168);
or I_58558 (I998199,I998007,I782677);
nor I_58559 (I998216,I782677,I782668);
nand I_58560 (I998233,I998072,I998216);
nand I_58561 (I998250,I998199,I998233);
DFFARX1 I_58562 (I998250,I2683,I997854,I997843,);
nor I_58563 (I998281,I998216,I997973);
DFFARX1 I_58564 (I998281,I2683,I997854,I997822,);
nor I_58565 (I998312,I782677,I782662);
DFFARX1 I_58566 (I998312,I2683,I997854,I998338,);
DFFARX1 I_58567 (I998338,I2683,I997854,I997837,);
not I_58568 (I998360,I998338);
nand I_58569 (I997834,I998360,I997888);
nand I_58570 (I997828,I998360,I997990);
not I_58571 (I998432,I2690);
DFFARX1 I_58572 (I398487,I2683,I998432,I998458,);
nand I_58573 (I998466,I998458,I398496);
not I_58574 (I998483,I998466);
DFFARX1 I_58575 (I398508,I2683,I998432,I998509,);
not I_58576 (I998517,I998509);
not I_58577 (I998534,I398499);
or I_58578 (I998551,I398493,I398499);
nor I_58579 (I998568,I398493,I398499);
or I_58580 (I998585,I398487,I398493);
DFFARX1 I_58581 (I998585,I2683,I998432,I998424,);
not I_58582 (I998616,I398490);
nand I_58583 (I998633,I998616,I398502);
nand I_58584 (I998650,I998534,I998633);
and I_58585 (I998403,I998517,I998650);
nor I_58586 (I998681,I398490,I398511);
and I_58587 (I998698,I998517,I998681);
nor I_58588 (I998409,I998483,I998698);
DFFARX1 I_58589 (I998681,I2683,I998432,I998738,);
not I_58590 (I998746,I998738);
nor I_58591 (I998418,I998517,I998746);
or I_58592 (I998777,I998585,I398505);
nor I_58593 (I998794,I398505,I398487);
nand I_58594 (I998811,I998650,I998794);
nand I_58595 (I998828,I998777,I998811);
DFFARX1 I_58596 (I998828,I2683,I998432,I998421,);
nor I_58597 (I998859,I998794,I998551);
DFFARX1 I_58598 (I998859,I2683,I998432,I998400,);
nor I_58599 (I998890,I398505,I398490);
DFFARX1 I_58600 (I998890,I2683,I998432,I998916,);
DFFARX1 I_58601 (I998916,I2683,I998432,I998415,);
not I_58602 (I998938,I998916);
nand I_58603 (I998412,I998938,I998466);
nand I_58604 (I998406,I998938,I998568);
not I_58605 (I999010,I2690);
DFFARX1 I_58606 (I30069,I2683,I999010,I999036,);
nand I_58607 (I999044,I999036,I30063);
not I_58608 (I999061,I999044);
DFFARX1 I_58609 (I30081,I2683,I999010,I999087,);
not I_58610 (I999095,I999087);
not I_58611 (I999112,I30084);
or I_58612 (I999129,I30087,I30084);
nor I_58613 (I999146,I30087,I30084);
or I_58614 (I999163,I30072,I30087);
DFFARX1 I_58615 (I999163,I2683,I999010,I999002,);
not I_58616 (I999194,I30075);
nand I_58617 (I999211,I999194,I30078);
nand I_58618 (I999228,I999112,I999211);
and I_58619 (I998981,I999095,I999228);
nor I_58620 (I999259,I30075,I30066);
and I_58621 (I999276,I999095,I999259);
nor I_58622 (I998987,I999061,I999276);
DFFARX1 I_58623 (I999259,I2683,I999010,I999316,);
not I_58624 (I999324,I999316);
nor I_58625 (I998996,I999095,I999324);
or I_58626 (I999355,I999163,I30066);
nor I_58627 (I999372,I30066,I30072);
nand I_58628 (I999389,I999228,I999372);
nand I_58629 (I999406,I999355,I999389);
DFFARX1 I_58630 (I999406,I2683,I999010,I998999,);
nor I_58631 (I999437,I999372,I999129);
DFFARX1 I_58632 (I999437,I2683,I999010,I998978,);
nor I_58633 (I999468,I30066,I30063);
DFFARX1 I_58634 (I999468,I2683,I999010,I999494,);
DFFARX1 I_58635 (I999494,I2683,I999010,I998993,);
not I_58636 (I999516,I999494);
nand I_58637 (I998990,I999516,I999044);
nand I_58638 (I998984,I999516,I999146);
not I_58639 (I999588,I2690);
DFFARX1 I_58640 (I570544,I2683,I999588,I999614,);
nand I_58641 (I999622,I999614,I570547);
not I_58642 (I999639,I999622);
DFFARX1 I_58643 (I570559,I2683,I999588,I999665,);
not I_58644 (I999673,I999665);
not I_58645 (I999690,I570544);
or I_58646 (I999707,I570553,I570544);
nor I_58647 (I999724,I570553,I570544);
or I_58648 (I999741,I570562,I570553);
DFFARX1 I_58649 (I999741,I2683,I999588,I999580,);
not I_58650 (I999772,I570565);
nand I_58651 (I999789,I999772,I570547);
nand I_58652 (I999806,I999690,I999789);
and I_58653 (I999559,I999673,I999806);
nor I_58654 (I999837,I570565,I570550);
and I_58655 (I999854,I999673,I999837);
nor I_58656 (I999565,I999639,I999854);
DFFARX1 I_58657 (I999837,I2683,I999588,I999894,);
not I_58658 (I999902,I999894);
nor I_58659 (I999574,I999673,I999902);
or I_58660 (I999933,I999741,I570556);
nor I_58661 (I999950,I570556,I570562);
nand I_58662 (I999967,I999806,I999950);
nand I_58663 (I999984,I999933,I999967);
DFFARX1 I_58664 (I999984,I2683,I999588,I999577,);
nor I_58665 (I1000015,I999950,I999707);
DFFARX1 I_58666 (I1000015,I2683,I999588,I999556,);
nor I_58667 (I1000046,I570556,I570568);
DFFARX1 I_58668 (I1000046,I2683,I999588,I1000072,);
DFFARX1 I_58669 (I1000072,I2683,I999588,I999571,);
not I_58670 (I1000094,I1000072);
nand I_58671 (I999568,I1000094,I999622);
nand I_58672 (I999562,I1000094,I999724);
not I_58673 (I1000166,I2690);
DFFARX1 I_58674 (I703847,I2683,I1000166,I1000192,);
nand I_58675 (I1000200,I1000192,I703868);
not I_58676 (I1000217,I1000200);
DFFARX1 I_58677 (I703841,I2683,I1000166,I1000243,);
not I_58678 (I1000251,I1000243);
not I_58679 (I1000268,I703862);
or I_58680 (I1000285,I703853,I703862);
nor I_58681 (I1000302,I703853,I703862);
or I_58682 (I1000319,I703856,I703853);
DFFARX1 I_58683 (I1000319,I2683,I1000166,I1000158,);
not I_58684 (I1000350,I703844);
nand I_58685 (I1000367,I1000350,I703859);
nand I_58686 (I1000384,I1000268,I1000367);
and I_58687 (I1000137,I1000251,I1000384);
nor I_58688 (I1000415,I703844,I703841);
and I_58689 (I1000432,I1000251,I1000415);
nor I_58690 (I1000143,I1000217,I1000432);
DFFARX1 I_58691 (I1000415,I2683,I1000166,I1000472,);
not I_58692 (I1000480,I1000472);
nor I_58693 (I1000152,I1000251,I1000480);
or I_58694 (I1000511,I1000319,I703865);
nor I_58695 (I1000528,I703865,I703856);
nand I_58696 (I1000545,I1000384,I1000528);
nand I_58697 (I1000562,I1000511,I1000545);
DFFARX1 I_58698 (I1000562,I2683,I1000166,I1000155,);
nor I_58699 (I1000593,I1000528,I1000285);
DFFARX1 I_58700 (I1000593,I2683,I1000166,I1000134,);
nor I_58701 (I1000624,I703865,I703850);
DFFARX1 I_58702 (I1000624,I2683,I1000166,I1000650,);
DFFARX1 I_58703 (I1000650,I2683,I1000166,I1000149,);
not I_58704 (I1000672,I1000650);
nand I_58705 (I1000146,I1000672,I1000200);
nand I_58706 (I1000140,I1000672,I1000302);
not I_58707 (I1000744,I2690);
DFFARX1 I_58708 (I410387,I2683,I1000744,I1000770,);
nand I_58709 (I1000778,I1000770,I410396);
not I_58710 (I1000795,I1000778);
DFFARX1 I_58711 (I410408,I2683,I1000744,I1000821,);
not I_58712 (I1000829,I1000821);
not I_58713 (I1000846,I410399);
or I_58714 (I1000863,I410393,I410399);
nor I_58715 (I1000880,I410393,I410399);
or I_58716 (I1000897,I410387,I410393);
DFFARX1 I_58717 (I1000897,I2683,I1000744,I1000736,);
not I_58718 (I1000928,I410390);
nand I_58719 (I1000945,I1000928,I410402);
nand I_58720 (I1000962,I1000846,I1000945);
and I_58721 (I1000715,I1000829,I1000962);
nor I_58722 (I1000993,I410390,I410411);
and I_58723 (I1001010,I1000829,I1000993);
nor I_58724 (I1000721,I1000795,I1001010);
DFFARX1 I_58725 (I1000993,I2683,I1000744,I1001050,);
not I_58726 (I1001058,I1001050);
nor I_58727 (I1000730,I1000829,I1001058);
or I_58728 (I1001089,I1000897,I410405);
nor I_58729 (I1001106,I410405,I410387);
nand I_58730 (I1001123,I1000962,I1001106);
nand I_58731 (I1001140,I1001089,I1001123);
DFFARX1 I_58732 (I1001140,I2683,I1000744,I1000733,);
nor I_58733 (I1001171,I1001106,I1000863);
DFFARX1 I_58734 (I1001171,I2683,I1000744,I1000712,);
nor I_58735 (I1001202,I410405,I410390);
DFFARX1 I_58736 (I1001202,I2683,I1000744,I1001228,);
DFFARX1 I_58737 (I1001228,I2683,I1000744,I1000727,);
not I_58738 (I1001250,I1001228);
nand I_58739 (I1000724,I1001250,I1000778);
nand I_58740 (I1000718,I1001250,I1000880);
not I_58741 (I1001322,I2690);
DFFARX1 I_58742 (I947282,I2683,I1001322,I1001348,);
nand I_58743 (I1001356,I1001348,I947267);
not I_58744 (I1001373,I1001356);
DFFARX1 I_58745 (I947270,I2683,I1001322,I1001399,);
not I_58746 (I1001407,I1001399);
not I_58747 (I1001424,I947285);
or I_58748 (I1001441,I947288,I947285);
nor I_58749 (I1001458,I947288,I947285);
or I_58750 (I1001475,I947264,I947288);
DFFARX1 I_58751 (I1001475,I2683,I1001322,I1001314,);
not I_58752 (I1001506,I947276);
nand I_58753 (I1001523,I1001506,I947279);
nand I_58754 (I1001540,I1001424,I1001523);
and I_58755 (I1001293,I1001407,I1001540);
nor I_58756 (I1001571,I947276,I947273);
and I_58757 (I1001588,I1001407,I1001571);
nor I_58758 (I1001299,I1001373,I1001588);
DFFARX1 I_58759 (I1001571,I2683,I1001322,I1001628,);
not I_58760 (I1001636,I1001628);
nor I_58761 (I1001308,I1001407,I1001636);
or I_58762 (I1001667,I1001475,I947264);
nor I_58763 (I1001684,I947264,I947264);
nand I_58764 (I1001701,I1001540,I1001684);
nand I_58765 (I1001718,I1001667,I1001701);
DFFARX1 I_58766 (I1001718,I2683,I1001322,I1001311,);
nor I_58767 (I1001749,I1001684,I1001441);
DFFARX1 I_58768 (I1001749,I2683,I1001322,I1001290,);
nor I_58769 (I1001780,I947264,I947267);
DFFARX1 I_58770 (I1001780,I2683,I1001322,I1001806,);
DFFARX1 I_58771 (I1001806,I2683,I1001322,I1001305,);
not I_58772 (I1001828,I1001806);
nand I_58773 (I1001302,I1001828,I1001356);
nand I_58774 (I1001296,I1001828,I1001458);
not I_58775 (I1001900,I2690);
DFFARX1 I_58776 (I949016,I2683,I1001900,I1001926,);
nand I_58777 (I1001934,I1001926,I949001);
not I_58778 (I1001951,I1001934);
DFFARX1 I_58779 (I949004,I2683,I1001900,I1001977,);
not I_58780 (I1001985,I1001977);
not I_58781 (I1002002,I949019);
or I_58782 (I1002019,I949022,I949019);
nor I_58783 (I1002036,I949022,I949019);
or I_58784 (I1002053,I948998,I949022);
DFFARX1 I_58785 (I1002053,I2683,I1001900,I1001892,);
not I_58786 (I1002084,I949010);
nand I_58787 (I1002101,I1002084,I949013);
nand I_58788 (I1002118,I1002002,I1002101);
and I_58789 (I1001871,I1001985,I1002118);
nor I_58790 (I1002149,I949010,I949007);
and I_58791 (I1002166,I1001985,I1002149);
nor I_58792 (I1001877,I1001951,I1002166);
DFFARX1 I_58793 (I1002149,I2683,I1001900,I1002206,);
not I_58794 (I1002214,I1002206);
nor I_58795 (I1001886,I1001985,I1002214);
or I_58796 (I1002245,I1002053,I948998);
nor I_58797 (I1002262,I948998,I948998);
nand I_58798 (I1002279,I1002118,I1002262);
nand I_58799 (I1002296,I1002245,I1002279);
DFFARX1 I_58800 (I1002296,I2683,I1001900,I1001889,);
nor I_58801 (I1002327,I1002262,I1002019);
DFFARX1 I_58802 (I1002327,I2683,I1001900,I1001868,);
nor I_58803 (I1002358,I948998,I949001);
DFFARX1 I_58804 (I1002358,I2683,I1001900,I1002384,);
DFFARX1 I_58805 (I1002384,I2683,I1001900,I1001883,);
not I_58806 (I1002406,I1002384);
nand I_58807 (I1001880,I1002406,I1001934);
nand I_58808 (I1001874,I1002406,I1002036);
not I_58809 (I1002478,I2690);
DFFARX1 I_58810 (I885436,I2683,I1002478,I1002504,);
nand I_58811 (I1002512,I1002504,I885421);
not I_58812 (I1002529,I1002512);
DFFARX1 I_58813 (I885424,I2683,I1002478,I1002555,);
not I_58814 (I1002563,I1002555);
not I_58815 (I1002580,I885439);
or I_58816 (I1002597,I885442,I885439);
nor I_58817 (I1002614,I885442,I885439);
or I_58818 (I1002631,I885418,I885442);
DFFARX1 I_58819 (I1002631,I2683,I1002478,I1002470,);
not I_58820 (I1002662,I885430);
nand I_58821 (I1002679,I1002662,I885433);
nand I_58822 (I1002696,I1002580,I1002679);
and I_58823 (I1002449,I1002563,I1002696);
nor I_58824 (I1002727,I885430,I885427);
and I_58825 (I1002744,I1002563,I1002727);
nor I_58826 (I1002455,I1002529,I1002744);
DFFARX1 I_58827 (I1002727,I2683,I1002478,I1002784,);
not I_58828 (I1002792,I1002784);
nor I_58829 (I1002464,I1002563,I1002792);
or I_58830 (I1002823,I1002631,I885418);
nor I_58831 (I1002840,I885418,I885418);
nand I_58832 (I1002857,I1002696,I1002840);
nand I_58833 (I1002874,I1002823,I1002857);
DFFARX1 I_58834 (I1002874,I2683,I1002478,I1002467,);
nor I_58835 (I1002905,I1002840,I1002597);
DFFARX1 I_58836 (I1002905,I2683,I1002478,I1002446,);
nor I_58837 (I1002936,I885418,I885421);
DFFARX1 I_58838 (I1002936,I2683,I1002478,I1002962,);
DFFARX1 I_58839 (I1002962,I2683,I1002478,I1002461,);
not I_58840 (I1002984,I1002962);
nand I_58841 (I1002458,I1002984,I1002512);
nand I_58842 (I1002452,I1002984,I1002614);
not I_58843 (I1003056,I2690);
DFFARX1 I_58844 (I265927,I2683,I1003056,I1003082,);
nand I_58845 (I1003090,I1003082,I265948);
not I_58846 (I1003107,I1003090);
DFFARX1 I_58847 (I265942,I2683,I1003056,I1003133,);
not I_58848 (I1003141,I1003133);
not I_58849 (I1003158,I265930);
or I_58850 (I1003175,I265945,I265930);
nor I_58851 (I1003192,I265945,I265930);
or I_58852 (I1003209,I265936,I265945);
DFFARX1 I_58853 (I1003209,I2683,I1003056,I1003048,);
not I_58854 (I1003240,I265924);
nand I_58855 (I1003257,I1003240,I265921);
nand I_58856 (I1003274,I1003158,I1003257);
and I_58857 (I1003027,I1003141,I1003274);
nor I_58858 (I1003305,I265924,I265933);
and I_58859 (I1003322,I1003141,I1003305);
nor I_58860 (I1003033,I1003107,I1003322);
DFFARX1 I_58861 (I1003305,I2683,I1003056,I1003362,);
not I_58862 (I1003370,I1003362);
nor I_58863 (I1003042,I1003141,I1003370);
or I_58864 (I1003401,I1003209,I265939);
nor I_58865 (I1003418,I265939,I265936);
nand I_58866 (I1003435,I1003274,I1003418);
nand I_58867 (I1003452,I1003401,I1003435);
DFFARX1 I_58868 (I1003452,I2683,I1003056,I1003045,);
nor I_58869 (I1003483,I1003418,I1003175);
DFFARX1 I_58870 (I1003483,I2683,I1003056,I1003024,);
nor I_58871 (I1003514,I265939,I265921);
DFFARX1 I_58872 (I1003514,I2683,I1003056,I1003540,);
DFFARX1 I_58873 (I1003540,I2683,I1003056,I1003039,);
not I_58874 (I1003562,I1003540);
nand I_58875 (I1003036,I1003562,I1003090);
nand I_58876 (I1003030,I1003562,I1003192);
not I_58877 (I1003634,I2690);
DFFARX1 I_58878 (I373653,I2683,I1003634,I1003660,);
nand I_58879 (I1003668,I1003660,I373662);
not I_58880 (I1003685,I1003668);
DFFARX1 I_58881 (I373650,I2683,I1003634,I1003711,);
not I_58882 (I1003719,I1003711);
not I_58883 (I1003736,I373656);
or I_58884 (I1003753,I373650,I373656);
nor I_58885 (I1003770,I373650,I373656);
or I_58886 (I1003787,I373665,I373650);
DFFARX1 I_58887 (I1003787,I2683,I1003634,I1003626,);
not I_58888 (I1003818,I373659);
nand I_58889 (I1003835,I1003818,I373674);
nand I_58890 (I1003852,I1003736,I1003835);
and I_58891 (I1003605,I1003719,I1003852);
nor I_58892 (I1003883,I373659,I373677);
and I_58893 (I1003900,I1003719,I1003883);
nor I_58894 (I1003611,I1003685,I1003900);
DFFARX1 I_58895 (I1003883,I2683,I1003634,I1003940,);
not I_58896 (I1003948,I1003940);
nor I_58897 (I1003620,I1003719,I1003948);
or I_58898 (I1003979,I1003787,I373668);
nor I_58899 (I1003996,I373668,I373665);
nand I_58900 (I1004013,I1003852,I1003996);
nand I_58901 (I1004030,I1003979,I1004013);
DFFARX1 I_58902 (I1004030,I2683,I1003634,I1003623,);
nor I_58903 (I1004061,I1003996,I1003753);
DFFARX1 I_58904 (I1004061,I2683,I1003634,I1003602,);
nor I_58905 (I1004092,I373668,I373671);
DFFARX1 I_58906 (I1004092,I2683,I1003634,I1004118,);
DFFARX1 I_58907 (I1004118,I2683,I1003634,I1003617,);
not I_58908 (I1004140,I1004118);
nand I_58909 (I1003614,I1004140,I1003668);
nand I_58910 (I1003608,I1004140,I1003770);
not I_58911 (I1004212,I2690);
DFFARX1 I_58912 (I324149,I2683,I1004212,I1004238,);
nand I_58913 (I1004246,I1004238,I324158);
not I_58914 (I1004263,I1004246);
DFFARX1 I_58915 (I324146,I2683,I1004212,I1004289,);
not I_58916 (I1004297,I1004289);
not I_58917 (I1004314,I324152);
or I_58918 (I1004331,I324146,I324152);
nor I_58919 (I1004348,I324146,I324152);
or I_58920 (I1004365,I324161,I324146);
DFFARX1 I_58921 (I1004365,I2683,I1004212,I1004204,);
not I_58922 (I1004396,I324155);
nand I_58923 (I1004413,I1004396,I324170);
nand I_58924 (I1004430,I1004314,I1004413);
and I_58925 (I1004183,I1004297,I1004430);
nor I_58926 (I1004461,I324155,I324173);
and I_58927 (I1004478,I1004297,I1004461);
nor I_58928 (I1004189,I1004263,I1004478);
DFFARX1 I_58929 (I1004461,I2683,I1004212,I1004518,);
not I_58930 (I1004526,I1004518);
nor I_58931 (I1004198,I1004297,I1004526);
or I_58932 (I1004557,I1004365,I324164);
nor I_58933 (I1004574,I324164,I324161);
nand I_58934 (I1004591,I1004430,I1004574);
nand I_58935 (I1004608,I1004557,I1004591);
DFFARX1 I_58936 (I1004608,I2683,I1004212,I1004201,);
nor I_58937 (I1004639,I1004574,I1004331);
DFFARX1 I_58938 (I1004639,I2683,I1004212,I1004180,);
nor I_58939 (I1004670,I324164,I324167);
DFFARX1 I_58940 (I1004670,I2683,I1004212,I1004696,);
DFFARX1 I_58941 (I1004696,I2683,I1004212,I1004195,);
not I_58942 (I1004718,I1004696);
nand I_58943 (I1004192,I1004718,I1004246);
nand I_58944 (I1004186,I1004718,I1004348);
not I_58945 (I1004790,I2690);
DFFARX1 I_58946 (I576902,I2683,I1004790,I1004816,);
nand I_58947 (I1004824,I1004816,I576905);
not I_58948 (I1004841,I1004824);
DFFARX1 I_58949 (I576917,I2683,I1004790,I1004867,);
not I_58950 (I1004875,I1004867);
not I_58951 (I1004892,I576902);
or I_58952 (I1004909,I576911,I576902);
nor I_58953 (I1004926,I576911,I576902);
or I_58954 (I1004943,I576920,I576911);
DFFARX1 I_58955 (I1004943,I2683,I1004790,I1004782,);
not I_58956 (I1004974,I576923);
nand I_58957 (I1004991,I1004974,I576905);
nand I_58958 (I1005008,I1004892,I1004991);
and I_58959 (I1004761,I1004875,I1005008);
nor I_58960 (I1005039,I576923,I576908);
and I_58961 (I1005056,I1004875,I1005039);
nor I_58962 (I1004767,I1004841,I1005056);
DFFARX1 I_58963 (I1005039,I2683,I1004790,I1005096,);
not I_58964 (I1005104,I1005096);
nor I_58965 (I1004776,I1004875,I1005104);
or I_58966 (I1005135,I1004943,I576914);
nor I_58967 (I1005152,I576914,I576920);
nand I_58968 (I1005169,I1005008,I1005152);
nand I_58969 (I1005186,I1005135,I1005169);
DFFARX1 I_58970 (I1005186,I2683,I1004790,I1004779,);
nor I_58971 (I1005217,I1005152,I1004909);
DFFARX1 I_58972 (I1005217,I2683,I1004790,I1004758,);
nor I_58973 (I1005248,I576914,I576926);
DFFARX1 I_58974 (I1005248,I2683,I1004790,I1005274,);
DFFARX1 I_58975 (I1005274,I2683,I1004790,I1004773,);
not I_58976 (I1005296,I1005274);
nand I_58977 (I1004770,I1005296,I1004824);
nand I_58978 (I1004764,I1005296,I1004926);
not I_58979 (I1005368,I2690);
DFFARX1 I_58980 (I243793,I2683,I1005368,I1005394,);
nand I_58981 (I1005402,I1005394,I243814);
not I_58982 (I1005419,I1005402);
DFFARX1 I_58983 (I243808,I2683,I1005368,I1005445,);
not I_58984 (I1005453,I1005445);
not I_58985 (I1005470,I243796);
or I_58986 (I1005487,I243811,I243796);
nor I_58987 (I1005504,I243811,I243796);
or I_58988 (I1005521,I243802,I243811);
DFFARX1 I_58989 (I1005521,I2683,I1005368,I1005360,);
not I_58990 (I1005552,I243790);
nand I_58991 (I1005569,I1005552,I243787);
nand I_58992 (I1005586,I1005470,I1005569);
and I_58993 (I1005339,I1005453,I1005586);
nor I_58994 (I1005617,I243790,I243799);
and I_58995 (I1005634,I1005453,I1005617);
nor I_58996 (I1005345,I1005419,I1005634);
DFFARX1 I_58997 (I1005617,I2683,I1005368,I1005674,);
not I_58998 (I1005682,I1005674);
nor I_58999 (I1005354,I1005453,I1005682);
or I_59000 (I1005713,I1005521,I243805);
nor I_59001 (I1005730,I243805,I243802);
nand I_59002 (I1005747,I1005586,I1005730);
nand I_59003 (I1005764,I1005713,I1005747);
DFFARX1 I_59004 (I1005764,I2683,I1005368,I1005357,);
nor I_59005 (I1005795,I1005730,I1005487);
DFFARX1 I_59006 (I1005795,I2683,I1005368,I1005336,);
nor I_59007 (I1005826,I243805,I243787);
DFFARX1 I_59008 (I1005826,I2683,I1005368,I1005852,);
DFFARX1 I_59009 (I1005852,I2683,I1005368,I1005351,);
not I_59010 (I1005874,I1005852);
nand I_59011 (I1005348,I1005874,I1005402);
nand I_59012 (I1005342,I1005874,I1005504);
not I_59013 (I1005946,I2690);
DFFARX1 I_59014 (I37447,I2683,I1005946,I1005972,);
nand I_59015 (I1005980,I1005972,I37441);
not I_59016 (I1005997,I1005980);
DFFARX1 I_59017 (I37459,I2683,I1005946,I1006023,);
not I_59018 (I1006031,I1006023);
not I_59019 (I1006048,I37462);
or I_59020 (I1006065,I37465,I37462);
nor I_59021 (I1006082,I37465,I37462);
or I_59022 (I1006099,I37450,I37465);
DFFARX1 I_59023 (I1006099,I2683,I1005946,I1005938,);
not I_59024 (I1006130,I37453);
nand I_59025 (I1006147,I1006130,I37456);
nand I_59026 (I1006164,I1006048,I1006147);
and I_59027 (I1005917,I1006031,I1006164);
nor I_59028 (I1006195,I37453,I37444);
and I_59029 (I1006212,I1006031,I1006195);
nor I_59030 (I1005923,I1005997,I1006212);
DFFARX1 I_59031 (I1006195,I2683,I1005946,I1006252,);
not I_59032 (I1006260,I1006252);
nor I_59033 (I1005932,I1006031,I1006260);
or I_59034 (I1006291,I1006099,I37444);
nor I_59035 (I1006308,I37444,I37450);
nand I_59036 (I1006325,I1006164,I1006308);
nand I_59037 (I1006342,I1006291,I1006325);
DFFARX1 I_59038 (I1006342,I2683,I1005946,I1005935,);
nor I_59039 (I1006373,I1006308,I1006065);
DFFARX1 I_59040 (I1006373,I2683,I1005946,I1005914,);
nor I_59041 (I1006404,I37444,I37441);
DFFARX1 I_59042 (I1006404,I2683,I1005946,I1006430,);
DFFARX1 I_59043 (I1006430,I2683,I1005946,I1005929,);
not I_59044 (I1006452,I1006430);
nand I_59045 (I1005926,I1006452,I1005980);
nand I_59046 (I1005920,I1006452,I1006082);
not I_59047 (I1006524,I2690);
DFFARX1 I_59048 (I99639,I2683,I1006524,I1006550,);
nand I_59049 (I1006558,I1006550,I99630);
not I_59050 (I1006575,I1006558);
DFFARX1 I_59051 (I99627,I2683,I1006524,I1006601,);
not I_59052 (I1006609,I1006601);
not I_59053 (I1006626,I99636);
or I_59054 (I1006643,I99627,I99636);
nor I_59055 (I1006660,I99627,I99636);
or I_59056 (I1006677,I99633,I99627);
DFFARX1 I_59057 (I1006677,I2683,I1006524,I1006516,);
not I_59058 (I1006708,I99642);
nand I_59059 (I1006725,I1006708,I99651);
nand I_59060 (I1006742,I1006626,I1006725);
and I_59061 (I1006495,I1006609,I1006742);
nor I_59062 (I1006773,I99642,I99645);
and I_59063 (I1006790,I1006609,I1006773);
nor I_59064 (I1006501,I1006575,I1006790);
DFFARX1 I_59065 (I1006773,I2683,I1006524,I1006830,);
not I_59066 (I1006838,I1006830);
nor I_59067 (I1006510,I1006609,I1006838);
or I_59068 (I1006869,I1006677,I99630);
nor I_59069 (I1006886,I99630,I99633);
nand I_59070 (I1006903,I1006742,I1006886);
nand I_59071 (I1006920,I1006869,I1006903);
DFFARX1 I_59072 (I1006920,I2683,I1006524,I1006513,);
nor I_59073 (I1006951,I1006886,I1006643);
DFFARX1 I_59074 (I1006951,I2683,I1006524,I1006492,);
nor I_59075 (I1006982,I99630,I99648);
DFFARX1 I_59076 (I1006982,I2683,I1006524,I1007008,);
DFFARX1 I_59077 (I1007008,I2683,I1006524,I1006507,);
not I_59078 (I1007030,I1007008);
nand I_59079 (I1006504,I1007030,I1006558);
nand I_59080 (I1006498,I1007030,I1006660);
not I_59081 (I1007102,I2690);
DFFARX1 I_59082 (I427047,I2683,I1007102,I1007128,);
nand I_59083 (I1007136,I1007128,I427056);
not I_59084 (I1007153,I1007136);
DFFARX1 I_59085 (I427068,I2683,I1007102,I1007179,);
not I_59086 (I1007187,I1007179);
not I_59087 (I1007204,I427059);
or I_59088 (I1007221,I427053,I427059);
nor I_59089 (I1007238,I427053,I427059);
or I_59090 (I1007255,I427047,I427053);
DFFARX1 I_59091 (I1007255,I2683,I1007102,I1007094,);
not I_59092 (I1007286,I427050);
nand I_59093 (I1007303,I1007286,I427062);
nand I_59094 (I1007320,I1007204,I1007303);
and I_59095 (I1007073,I1007187,I1007320);
nor I_59096 (I1007351,I427050,I427071);
and I_59097 (I1007368,I1007187,I1007351);
nor I_59098 (I1007079,I1007153,I1007368);
DFFARX1 I_59099 (I1007351,I2683,I1007102,I1007408,);
not I_59100 (I1007416,I1007408);
nor I_59101 (I1007088,I1007187,I1007416);
or I_59102 (I1007447,I1007255,I427065);
nor I_59103 (I1007464,I427065,I427047);
nand I_59104 (I1007481,I1007320,I1007464);
nand I_59105 (I1007498,I1007447,I1007481);
DFFARX1 I_59106 (I1007498,I2683,I1007102,I1007091,);
nor I_59107 (I1007529,I1007464,I1007221);
DFFARX1 I_59108 (I1007529,I2683,I1007102,I1007070,);
nor I_59109 (I1007560,I427065,I427050);
DFFARX1 I_59110 (I1007560,I2683,I1007102,I1007586,);
DFFARX1 I_59111 (I1007586,I2683,I1007102,I1007085,);
not I_59112 (I1007608,I1007586);
nand I_59113 (I1007082,I1007608,I1007136);
nand I_59114 (I1007076,I1007608,I1007238);
not I_59115 (I1007680,I2690);
DFFARX1 I_59116 (I399082,I2683,I1007680,I1007706,);
nand I_59117 (I1007714,I1007706,I399091);
not I_59118 (I1007731,I1007714);
DFFARX1 I_59119 (I399103,I2683,I1007680,I1007757,);
not I_59120 (I1007765,I1007757);
not I_59121 (I1007782,I399094);
or I_59122 (I1007799,I399088,I399094);
nor I_59123 (I1007816,I399088,I399094);
or I_59124 (I1007833,I399082,I399088);
DFFARX1 I_59125 (I1007833,I2683,I1007680,I1007672,);
not I_59126 (I1007864,I399085);
nand I_59127 (I1007881,I1007864,I399097);
nand I_59128 (I1007898,I1007782,I1007881);
and I_59129 (I1007651,I1007765,I1007898);
nor I_59130 (I1007929,I399085,I399106);
and I_59131 (I1007946,I1007765,I1007929);
nor I_59132 (I1007657,I1007731,I1007946);
DFFARX1 I_59133 (I1007929,I2683,I1007680,I1007986,);
not I_59134 (I1007994,I1007986);
nor I_59135 (I1007666,I1007765,I1007994);
or I_59136 (I1008025,I1007833,I399100);
nor I_59137 (I1008042,I399100,I399082);
nand I_59138 (I1008059,I1007898,I1008042);
nand I_59139 (I1008076,I1008025,I1008059);
DFFARX1 I_59140 (I1008076,I2683,I1007680,I1007669,);
nor I_59141 (I1008107,I1008042,I1007799);
DFFARX1 I_59142 (I1008107,I2683,I1007680,I1007648,);
nor I_59143 (I1008138,I399100,I399085);
DFFARX1 I_59144 (I1008138,I2683,I1007680,I1008164,);
DFFARX1 I_59145 (I1008164,I2683,I1007680,I1007663,);
not I_59146 (I1008186,I1008164);
nand I_59147 (I1007660,I1008186,I1007714);
nand I_59148 (I1007654,I1008186,I1007816);
not I_59149 (I1008258,I2690);
DFFARX1 I_59150 (I439341,I2683,I1008258,I1008284,);
nand I_59151 (I1008292,I1008284,I439356);
not I_59152 (I1008309,I1008292);
DFFARX1 I_59153 (I439338,I2683,I1008258,I1008335,);
not I_59154 (I1008343,I1008335);
not I_59155 (I1008360,I439347);
or I_59156 (I1008377,I439341,I439347);
nor I_59157 (I1008394,I439341,I439347);
or I_59158 (I1008411,I439338,I439341);
DFFARX1 I_59159 (I1008411,I2683,I1008258,I1008250,);
not I_59160 (I1008442,I439359);
nand I_59161 (I1008459,I1008442,I439362);
nand I_59162 (I1008476,I1008360,I1008459);
and I_59163 (I1008229,I1008343,I1008476);
nor I_59164 (I1008507,I439359,I439344);
and I_59165 (I1008524,I1008343,I1008507);
nor I_59166 (I1008235,I1008309,I1008524);
DFFARX1 I_59167 (I1008507,I2683,I1008258,I1008564,);
not I_59168 (I1008572,I1008564);
nor I_59169 (I1008244,I1008343,I1008572);
or I_59170 (I1008603,I1008411,I439350);
nor I_59171 (I1008620,I439350,I439338);
nand I_59172 (I1008637,I1008476,I1008620);
nand I_59173 (I1008654,I1008603,I1008637);
DFFARX1 I_59174 (I1008654,I2683,I1008258,I1008247,);
nor I_59175 (I1008685,I1008620,I1008377);
DFFARX1 I_59176 (I1008685,I2683,I1008258,I1008226,);
nor I_59177 (I1008716,I439350,I439353);
DFFARX1 I_59178 (I1008716,I2683,I1008258,I1008742,);
DFFARX1 I_59179 (I1008742,I2683,I1008258,I1008241,);
not I_59180 (I1008764,I1008742);
nand I_59181 (I1008238,I1008764,I1008292);
nand I_59182 (I1008232,I1008764,I1008394);
not I_59183 (I1008836,I2690);
DFFARX1 I_59184 (I348085,I2683,I1008836,I1008862,);
nand I_59185 (I1008870,I1008862,I348094);
not I_59186 (I1008887,I1008870);
DFFARX1 I_59187 (I348082,I2683,I1008836,I1008913,);
not I_59188 (I1008921,I1008913);
not I_59189 (I1008938,I348088);
or I_59190 (I1008955,I348082,I348088);
nor I_59191 (I1008972,I348082,I348088);
or I_59192 (I1008989,I348097,I348082);
DFFARX1 I_59193 (I1008989,I2683,I1008836,I1008828,);
not I_59194 (I1009020,I348091);
nand I_59195 (I1009037,I1009020,I348106);
nand I_59196 (I1009054,I1008938,I1009037);
and I_59197 (I1008807,I1008921,I1009054);
nor I_59198 (I1009085,I348091,I348109);
and I_59199 (I1009102,I1008921,I1009085);
nor I_59200 (I1008813,I1008887,I1009102);
DFFARX1 I_59201 (I1009085,I2683,I1008836,I1009142,);
not I_59202 (I1009150,I1009142);
nor I_59203 (I1008822,I1008921,I1009150);
or I_59204 (I1009181,I1008989,I348100);
nor I_59205 (I1009198,I348100,I348097);
nand I_59206 (I1009215,I1009054,I1009198);
nand I_59207 (I1009232,I1009181,I1009215);
DFFARX1 I_59208 (I1009232,I2683,I1008836,I1008825,);
nor I_59209 (I1009263,I1009198,I1008955);
DFFARX1 I_59210 (I1009263,I2683,I1008836,I1008804,);
nor I_59211 (I1009294,I348100,I348103);
DFFARX1 I_59212 (I1009294,I2683,I1008836,I1009320,);
DFFARX1 I_59213 (I1009320,I2683,I1008836,I1008819,);
not I_59214 (I1009342,I1009320);
nand I_59215 (I1008816,I1009342,I1008870);
nand I_59216 (I1008810,I1009342,I1008972);
not I_59217 (I1009414,I2690);
DFFARX1 I_59218 (I704493,I2683,I1009414,I1009440,);
nand I_59219 (I1009448,I1009440,I704514);
not I_59220 (I1009465,I1009448);
DFFARX1 I_59221 (I704487,I2683,I1009414,I1009491,);
not I_59222 (I1009499,I1009491);
not I_59223 (I1009516,I704508);
or I_59224 (I1009533,I704499,I704508);
nor I_59225 (I1009550,I704499,I704508);
or I_59226 (I1009567,I704502,I704499);
DFFARX1 I_59227 (I1009567,I2683,I1009414,I1009406,);
not I_59228 (I1009598,I704490);
nand I_59229 (I1009615,I1009598,I704505);
nand I_59230 (I1009632,I1009516,I1009615);
and I_59231 (I1009385,I1009499,I1009632);
nor I_59232 (I1009663,I704490,I704487);
and I_59233 (I1009680,I1009499,I1009663);
nor I_59234 (I1009391,I1009465,I1009680);
DFFARX1 I_59235 (I1009663,I2683,I1009414,I1009720,);
not I_59236 (I1009728,I1009720);
nor I_59237 (I1009400,I1009499,I1009728);
or I_59238 (I1009759,I1009567,I704511);
nor I_59239 (I1009776,I704511,I704502);
nand I_59240 (I1009793,I1009632,I1009776);
nand I_59241 (I1009810,I1009759,I1009793);
DFFARX1 I_59242 (I1009810,I2683,I1009414,I1009403,);
nor I_59243 (I1009841,I1009776,I1009533);
DFFARX1 I_59244 (I1009841,I2683,I1009414,I1009382,);
nor I_59245 (I1009872,I704511,I704496);
DFFARX1 I_59246 (I1009872,I2683,I1009414,I1009898,);
DFFARX1 I_59247 (I1009898,I2683,I1009414,I1009397,);
not I_59248 (I1009920,I1009898);
nand I_59249 (I1009394,I1009920,I1009448);
nand I_59250 (I1009388,I1009920,I1009550);
not I_59251 (I1009992,I2690);
DFFARX1 I_59252 (I705785,I2683,I1009992,I1010018,);
nand I_59253 (I1010026,I1010018,I705806);
not I_59254 (I1010043,I1010026);
DFFARX1 I_59255 (I705779,I2683,I1009992,I1010069,);
not I_59256 (I1010077,I1010069);
not I_59257 (I1010094,I705800);
or I_59258 (I1010111,I705791,I705800);
nor I_59259 (I1010128,I705791,I705800);
or I_59260 (I1010145,I705794,I705791);
DFFARX1 I_59261 (I1010145,I2683,I1009992,I1009984,);
not I_59262 (I1010176,I705782);
nand I_59263 (I1010193,I1010176,I705797);
nand I_59264 (I1010210,I1010094,I1010193);
and I_59265 (I1009963,I1010077,I1010210);
nor I_59266 (I1010241,I705782,I705779);
and I_59267 (I1010258,I1010077,I1010241);
nor I_59268 (I1009969,I1010043,I1010258);
DFFARX1 I_59269 (I1010241,I2683,I1009992,I1010298,);
not I_59270 (I1010306,I1010298);
nor I_59271 (I1009978,I1010077,I1010306);
or I_59272 (I1010337,I1010145,I705803);
nor I_59273 (I1010354,I705803,I705794);
nand I_59274 (I1010371,I1010210,I1010354);
nand I_59275 (I1010388,I1010337,I1010371);
DFFARX1 I_59276 (I1010388,I2683,I1009992,I1009981,);
nor I_59277 (I1010419,I1010354,I1010111);
DFFARX1 I_59278 (I1010419,I2683,I1009992,I1009960,);
nor I_59279 (I1010450,I705803,I705788);
DFFARX1 I_59280 (I1010450,I2683,I1009992,I1010476,);
DFFARX1 I_59281 (I1010476,I2683,I1009992,I1009975,);
not I_59282 (I1010498,I1010476);
nand I_59283 (I1009972,I1010498,I1010026);
nand I_59284 (I1009966,I1010498,I1010128);
not I_59285 (I1010570,I2690);
DFFARX1 I_59286 (I905088,I2683,I1010570,I1010596,);
nand I_59287 (I1010604,I1010596,I905073);
not I_59288 (I1010621,I1010604);
DFFARX1 I_59289 (I905076,I2683,I1010570,I1010647,);
not I_59290 (I1010655,I1010647);
not I_59291 (I1010672,I905091);
or I_59292 (I1010689,I905094,I905091);
nor I_59293 (I1010706,I905094,I905091);
or I_59294 (I1010723,I905070,I905094);
DFFARX1 I_59295 (I1010723,I2683,I1010570,I1010562,);
not I_59296 (I1010754,I905082);
nand I_59297 (I1010771,I1010754,I905085);
nand I_59298 (I1010788,I1010672,I1010771);
and I_59299 (I1010541,I1010655,I1010788);
nor I_59300 (I1010819,I905082,I905079);
and I_59301 (I1010836,I1010655,I1010819);
nor I_59302 (I1010547,I1010621,I1010836);
DFFARX1 I_59303 (I1010819,I2683,I1010570,I1010876,);
not I_59304 (I1010884,I1010876);
nor I_59305 (I1010556,I1010655,I1010884);
or I_59306 (I1010915,I1010723,I905070);
nor I_59307 (I1010932,I905070,I905070);
nand I_59308 (I1010949,I1010788,I1010932);
nand I_59309 (I1010966,I1010915,I1010949);
DFFARX1 I_59310 (I1010966,I2683,I1010570,I1010559,);
nor I_59311 (I1010997,I1010932,I1010689);
DFFARX1 I_59312 (I1010997,I2683,I1010570,I1010538,);
nor I_59313 (I1011028,I905070,I905073);
DFFARX1 I_59314 (I1011028,I2683,I1010570,I1011054,);
DFFARX1 I_59315 (I1011054,I2683,I1010570,I1010553,);
not I_59316 (I1011076,I1011054);
nand I_59317 (I1010550,I1011076,I1010604);
nand I_59318 (I1010544,I1011076,I1010706);
not I_59319 (I1011148,I2690);
DFFARX1 I_59320 (I1047758,I2683,I1011148,I1011174,);
nand I_59321 (I1011182,I1011174,I1047749);
not I_59322 (I1011199,I1011182);
DFFARX1 I_59323 (I1047734,I2683,I1011148,I1011225,);
not I_59324 (I1011233,I1011225);
not I_59325 (I1011250,I1047737);
or I_59326 (I1011267,I1047746,I1047737);
nor I_59327 (I1011284,I1047746,I1047737);
or I_59328 (I1011301,I1047743,I1047746);
DFFARX1 I_59329 (I1011301,I2683,I1011148,I1011140,);
not I_59330 (I1011332,I1047755);
nand I_59331 (I1011349,I1011332,I1047734);
nand I_59332 (I1011366,I1011250,I1011349);
and I_59333 (I1011119,I1011233,I1011366);
nor I_59334 (I1011397,I1047755,I1047740);
and I_59335 (I1011414,I1011233,I1011397);
nor I_59336 (I1011125,I1011199,I1011414);
DFFARX1 I_59337 (I1011397,I2683,I1011148,I1011454,);
not I_59338 (I1011462,I1011454);
nor I_59339 (I1011134,I1011233,I1011462);
or I_59340 (I1011493,I1011301,I1047761);
nor I_59341 (I1011510,I1047761,I1047743);
nand I_59342 (I1011527,I1011366,I1011510);
nand I_59343 (I1011544,I1011493,I1011527);
DFFARX1 I_59344 (I1011544,I2683,I1011148,I1011137,);
nor I_59345 (I1011575,I1011510,I1011267);
DFFARX1 I_59346 (I1011575,I2683,I1011148,I1011116,);
nor I_59347 (I1011606,I1047761,I1047752);
DFFARX1 I_59348 (I1011606,I2683,I1011148,I1011632,);
DFFARX1 I_59349 (I1011632,I2683,I1011148,I1011131,);
not I_59350 (I1011654,I1011632);
nand I_59351 (I1011128,I1011654,I1011182);
nand I_59352 (I1011122,I1011654,I1011284);
not I_59353 (I1011726,I2690);
DFFARX1 I_59354 (I682866,I2683,I1011726,I1011752,);
nand I_59355 (I1011760,I1011752,I682866);
not I_59356 (I1011777,I1011760);
DFFARX1 I_59357 (I682872,I2683,I1011726,I1011803,);
not I_59358 (I1011811,I1011803);
not I_59359 (I1011828,I682884);
or I_59360 (I1011845,I682869,I682884);
nor I_59361 (I1011862,I682869,I682884);
or I_59362 (I1011879,I682863,I682869);
DFFARX1 I_59363 (I1011879,I2683,I1011726,I1011718,);
not I_59364 (I1011910,I682881);
nand I_59365 (I1011927,I1011910,I682875);
nand I_59366 (I1011944,I1011828,I1011927);
and I_59367 (I1011697,I1011811,I1011944);
nor I_59368 (I1011975,I682881,I682863);
and I_59369 (I1011992,I1011811,I1011975);
nor I_59370 (I1011703,I1011777,I1011992);
DFFARX1 I_59371 (I1011975,I2683,I1011726,I1012032,);
not I_59372 (I1012040,I1012032);
nor I_59373 (I1011712,I1011811,I1012040);
or I_59374 (I1012071,I1011879,I682878);
nor I_59375 (I1012088,I682878,I682863);
nand I_59376 (I1012105,I1011944,I1012088);
nand I_59377 (I1012122,I1012071,I1012105);
DFFARX1 I_59378 (I1012122,I2683,I1011726,I1011715,);
nor I_59379 (I1012153,I1012088,I1011845);
DFFARX1 I_59380 (I1012153,I2683,I1011726,I1011694,);
nor I_59381 (I1012184,I682878,I682869);
DFFARX1 I_59382 (I1012184,I2683,I1011726,I1012210,);
DFFARX1 I_59383 (I1012210,I2683,I1011726,I1011709,);
not I_59384 (I1012232,I1012210);
nand I_59385 (I1011706,I1012232,I1011760);
nand I_59386 (I1011700,I1012232,I1011862);
not I_59387 (I1012304,I2690);
DFFARX1 I_59388 (I890638,I2683,I1012304,I1012330,);
nand I_59389 (I1012338,I1012330,I890623);
not I_59390 (I1012355,I1012338);
DFFARX1 I_59391 (I890626,I2683,I1012304,I1012381,);
not I_59392 (I1012389,I1012381);
not I_59393 (I1012406,I890641);
or I_59394 (I1012423,I890644,I890641);
nor I_59395 (I1012440,I890644,I890641);
or I_59396 (I1012457,I890620,I890644);
DFFARX1 I_59397 (I1012457,I2683,I1012304,I1012296,);
not I_59398 (I1012488,I890632);
nand I_59399 (I1012505,I1012488,I890635);
nand I_59400 (I1012522,I1012406,I1012505);
and I_59401 (I1012275,I1012389,I1012522);
nor I_59402 (I1012553,I890632,I890629);
and I_59403 (I1012570,I1012389,I1012553);
nor I_59404 (I1012281,I1012355,I1012570);
DFFARX1 I_59405 (I1012553,I2683,I1012304,I1012610,);
not I_59406 (I1012618,I1012610);
nor I_59407 (I1012290,I1012389,I1012618);
or I_59408 (I1012649,I1012457,I890620);
nor I_59409 (I1012666,I890620,I890620);
nand I_59410 (I1012683,I1012522,I1012666);
nand I_59411 (I1012700,I1012649,I1012683);
DFFARX1 I_59412 (I1012700,I2683,I1012304,I1012293,);
nor I_59413 (I1012731,I1012666,I1012423);
DFFARX1 I_59414 (I1012731,I2683,I1012304,I1012272,);
nor I_59415 (I1012762,I890620,I890623);
DFFARX1 I_59416 (I1012762,I2683,I1012304,I1012788,);
DFFARX1 I_59417 (I1012788,I2683,I1012304,I1012287,);
not I_59418 (I1012810,I1012788);
nand I_59419 (I1012284,I1012810,I1012338);
nand I_59420 (I1012278,I1012810,I1012440);
not I_59421 (I1012882,I2690);
DFFARX1 I_59422 (I765217,I2683,I1012882,I1012908,);
nand I_59423 (I1012916,I1012908,I765238);
not I_59424 (I1012933,I1012916);
DFFARX1 I_59425 (I765211,I2683,I1012882,I1012959,);
not I_59426 (I1012967,I1012959);
not I_59427 (I1012984,I765232);
or I_59428 (I1013001,I765223,I765232);
nor I_59429 (I1013018,I765223,I765232);
or I_59430 (I1013035,I765226,I765223);
DFFARX1 I_59431 (I1013035,I2683,I1012882,I1012874,);
not I_59432 (I1013066,I765214);
nand I_59433 (I1013083,I1013066,I765229);
nand I_59434 (I1013100,I1012984,I1013083);
and I_59435 (I1012853,I1012967,I1013100);
nor I_59436 (I1013131,I765214,I765211);
and I_59437 (I1013148,I1012967,I1013131);
nor I_59438 (I1012859,I1012933,I1013148);
DFFARX1 I_59439 (I1013131,I2683,I1012882,I1013188,);
not I_59440 (I1013196,I1013188);
nor I_59441 (I1012868,I1012967,I1013196);
or I_59442 (I1013227,I1013035,I765235);
nor I_59443 (I1013244,I765235,I765226);
nand I_59444 (I1013261,I1013100,I1013244);
nand I_59445 (I1013278,I1013227,I1013261);
DFFARX1 I_59446 (I1013278,I2683,I1012882,I1012871,);
nor I_59447 (I1013309,I1013244,I1013001);
DFFARX1 I_59448 (I1013309,I2683,I1012882,I1012850,);
nor I_59449 (I1013340,I765235,I765220);
DFFARX1 I_59450 (I1013340,I2683,I1012882,I1013366,);
DFFARX1 I_59451 (I1013366,I2683,I1012882,I1012865,);
not I_59452 (I1013388,I1013366);
nand I_59453 (I1012862,I1013388,I1012916);
nand I_59454 (I1012856,I1013388,I1013018);
not I_59455 (I1013460,I2690);
DFFARX1 I_59456 (I338837,I2683,I1013460,I1013486,);
nand I_59457 (I1013494,I1013486,I338846);
not I_59458 (I1013511,I1013494);
DFFARX1 I_59459 (I338834,I2683,I1013460,I1013537,);
not I_59460 (I1013545,I1013537);
not I_59461 (I1013562,I338840);
or I_59462 (I1013579,I338834,I338840);
nor I_59463 (I1013596,I338834,I338840);
or I_59464 (I1013613,I338849,I338834);
DFFARX1 I_59465 (I1013613,I2683,I1013460,I1013452,);
not I_59466 (I1013644,I338843);
nand I_59467 (I1013661,I1013644,I338858);
nand I_59468 (I1013678,I1013562,I1013661);
and I_59469 (I1013431,I1013545,I1013678);
nor I_59470 (I1013709,I338843,I338861);
and I_59471 (I1013726,I1013545,I1013709);
nor I_59472 (I1013437,I1013511,I1013726);
DFFARX1 I_59473 (I1013709,I2683,I1013460,I1013766,);
not I_59474 (I1013774,I1013766);
nor I_59475 (I1013446,I1013545,I1013774);
or I_59476 (I1013805,I1013613,I338852);
nor I_59477 (I1013822,I338852,I338849);
nand I_59478 (I1013839,I1013678,I1013822);
nand I_59479 (I1013856,I1013805,I1013839);
DFFARX1 I_59480 (I1013856,I2683,I1013460,I1013449,);
nor I_59481 (I1013887,I1013822,I1013579);
DFFARX1 I_59482 (I1013887,I2683,I1013460,I1013428,);
nor I_59483 (I1013918,I338852,I338855);
DFFARX1 I_59484 (I1013918,I2683,I1013460,I1013944,);
DFFARX1 I_59485 (I1013944,I2683,I1013460,I1013443,);
not I_59486 (I1013966,I1013944);
nand I_59487 (I1013440,I1013966,I1013494);
nand I_59488 (I1013434,I1013966,I1013596);
not I_59489 (I1014038,I2690);
DFFARX1 I_59490 (I894684,I2683,I1014038,I1014064,);
nand I_59491 (I1014072,I1014064,I894669);
not I_59492 (I1014089,I1014072);
DFFARX1 I_59493 (I894672,I2683,I1014038,I1014115,);
not I_59494 (I1014123,I1014115);
not I_59495 (I1014140,I894687);
or I_59496 (I1014157,I894690,I894687);
nor I_59497 (I1014174,I894690,I894687);
or I_59498 (I1014191,I894666,I894690);
DFFARX1 I_59499 (I1014191,I2683,I1014038,I1014030,);
not I_59500 (I1014222,I894678);
nand I_59501 (I1014239,I1014222,I894681);
nand I_59502 (I1014256,I1014140,I1014239);
and I_59503 (I1014009,I1014123,I1014256);
nor I_59504 (I1014287,I894678,I894675);
and I_59505 (I1014304,I1014123,I1014287);
nor I_59506 (I1014015,I1014089,I1014304);
DFFARX1 I_59507 (I1014287,I2683,I1014038,I1014344,);
not I_59508 (I1014352,I1014344);
nor I_59509 (I1014024,I1014123,I1014352);
or I_59510 (I1014383,I1014191,I894666);
nor I_59511 (I1014400,I894666,I894666);
nand I_59512 (I1014417,I1014256,I1014400);
nand I_59513 (I1014434,I1014383,I1014417);
DFFARX1 I_59514 (I1014434,I2683,I1014038,I1014027,);
nor I_59515 (I1014465,I1014400,I1014157);
DFFARX1 I_59516 (I1014465,I2683,I1014038,I1014006,);
nor I_59517 (I1014496,I894666,I894669);
DFFARX1 I_59518 (I1014496,I2683,I1014038,I1014522,);
DFFARX1 I_59519 (I1014522,I2683,I1014038,I1014021,);
not I_59520 (I1014544,I1014522);
nand I_59521 (I1014018,I1014544,I1014072);
nand I_59522 (I1014012,I1014544,I1014174);
not I_59523 (I1014616,I2690);
DFFARX1 I_59524 (I87518,I2683,I1014616,I1014642,);
nand I_59525 (I1014650,I1014642,I87509);
not I_59526 (I1014667,I1014650);
DFFARX1 I_59527 (I87506,I2683,I1014616,I1014693,);
not I_59528 (I1014701,I1014693);
not I_59529 (I1014718,I87515);
or I_59530 (I1014735,I87506,I87515);
nor I_59531 (I1014752,I87506,I87515);
or I_59532 (I1014769,I87512,I87506);
DFFARX1 I_59533 (I1014769,I2683,I1014616,I1014608,);
not I_59534 (I1014800,I87521);
nand I_59535 (I1014817,I1014800,I87530);
nand I_59536 (I1014834,I1014718,I1014817);
and I_59537 (I1014587,I1014701,I1014834);
nor I_59538 (I1014865,I87521,I87524);
and I_59539 (I1014882,I1014701,I1014865);
nor I_59540 (I1014593,I1014667,I1014882);
DFFARX1 I_59541 (I1014865,I2683,I1014616,I1014922,);
not I_59542 (I1014930,I1014922);
nor I_59543 (I1014602,I1014701,I1014930);
or I_59544 (I1014961,I1014769,I87509);
nor I_59545 (I1014978,I87509,I87512);
nand I_59546 (I1014995,I1014834,I1014978);
nand I_59547 (I1015012,I1014961,I1014995);
DFFARX1 I_59548 (I1015012,I2683,I1014616,I1014605,);
nor I_59549 (I1015043,I1014978,I1014735);
DFFARX1 I_59550 (I1015043,I2683,I1014616,I1014584,);
nor I_59551 (I1015074,I87509,I87527);
DFFARX1 I_59552 (I1015074,I2683,I1014616,I1015100,);
DFFARX1 I_59553 (I1015100,I2683,I1014616,I1014599,);
not I_59554 (I1015122,I1015100);
nand I_59555 (I1014596,I1015122,I1014650);
nand I_59556 (I1014590,I1015122,I1014752);
not I_59557 (I1015194,I2690);
DFFARX1 I_59558 (I41663,I2683,I1015194,I1015220,);
nand I_59559 (I1015228,I1015220,I41657);
not I_59560 (I1015245,I1015228);
DFFARX1 I_59561 (I41675,I2683,I1015194,I1015271,);
not I_59562 (I1015279,I1015271);
not I_59563 (I1015296,I41678);
or I_59564 (I1015313,I41681,I41678);
nor I_59565 (I1015330,I41681,I41678);
or I_59566 (I1015347,I41666,I41681);
DFFARX1 I_59567 (I1015347,I2683,I1015194,I1015186,);
not I_59568 (I1015378,I41669);
nand I_59569 (I1015395,I1015378,I41672);
nand I_59570 (I1015412,I1015296,I1015395);
and I_59571 (I1015165,I1015279,I1015412);
nor I_59572 (I1015443,I41669,I41660);
and I_59573 (I1015460,I1015279,I1015443);
nor I_59574 (I1015171,I1015245,I1015460);
DFFARX1 I_59575 (I1015443,I2683,I1015194,I1015500,);
not I_59576 (I1015508,I1015500);
nor I_59577 (I1015180,I1015279,I1015508);
or I_59578 (I1015539,I1015347,I41660);
nor I_59579 (I1015556,I41660,I41666);
nand I_59580 (I1015573,I1015412,I1015556);
nand I_59581 (I1015590,I1015539,I1015573);
DFFARX1 I_59582 (I1015590,I2683,I1015194,I1015183,);
nor I_59583 (I1015621,I1015556,I1015313);
DFFARX1 I_59584 (I1015621,I2683,I1015194,I1015162,);
nor I_59585 (I1015652,I41660,I41657);
DFFARX1 I_59586 (I1015652,I2683,I1015194,I1015678,);
DFFARX1 I_59587 (I1015678,I2683,I1015194,I1015177,);
not I_59588 (I1015700,I1015678);
nand I_59589 (I1015174,I1015700,I1015228);
nand I_59590 (I1015168,I1015700,I1015330);
not I_59591 (I1015772,I2690);
DFFARX1 I_59592 (I320341,I2683,I1015772,I1015798,);
nand I_59593 (I1015806,I1015798,I320350);
not I_59594 (I1015823,I1015806);
DFFARX1 I_59595 (I320338,I2683,I1015772,I1015849,);
not I_59596 (I1015857,I1015849);
not I_59597 (I1015874,I320344);
or I_59598 (I1015891,I320338,I320344);
nor I_59599 (I1015908,I320338,I320344);
or I_59600 (I1015925,I320353,I320338);
DFFARX1 I_59601 (I1015925,I2683,I1015772,I1015764,);
not I_59602 (I1015956,I320347);
nand I_59603 (I1015973,I1015956,I320362);
nand I_59604 (I1015990,I1015874,I1015973);
and I_59605 (I1015743,I1015857,I1015990);
nor I_59606 (I1016021,I320347,I320365);
and I_59607 (I1016038,I1015857,I1016021);
nor I_59608 (I1015749,I1015823,I1016038);
DFFARX1 I_59609 (I1016021,I2683,I1015772,I1016078,);
not I_59610 (I1016086,I1016078);
nor I_59611 (I1015758,I1015857,I1016086);
or I_59612 (I1016117,I1015925,I320356);
nor I_59613 (I1016134,I320356,I320353);
nand I_59614 (I1016151,I1015990,I1016134);
nand I_59615 (I1016168,I1016117,I1016151);
DFFARX1 I_59616 (I1016168,I2683,I1015772,I1015761,);
nor I_59617 (I1016199,I1016134,I1015891);
DFFARX1 I_59618 (I1016199,I2683,I1015772,I1015740,);
nor I_59619 (I1016230,I320356,I320359);
DFFARX1 I_59620 (I1016230,I2683,I1015772,I1016256,);
DFFARX1 I_59621 (I1016256,I2683,I1015772,I1015755,);
not I_59622 (I1016278,I1016256);
nand I_59623 (I1015752,I1016278,I1015806);
nand I_59624 (I1015746,I1016278,I1015908);
not I_59625 (I1016350,I2690);
DFFARX1 I_59626 (I158685,I2683,I1016350,I1016376,);
nand I_59627 (I1016384,I1016376,I158688);
not I_59628 (I1016401,I1016384);
DFFARX1 I_59629 (I158697,I2683,I1016350,I1016427,);
not I_59630 (I1016435,I1016427);
not I_59631 (I1016452,I158700);
or I_59632 (I1016469,I158691,I158700);
nor I_59633 (I1016486,I158691,I158700);
or I_59634 (I1016503,I158703,I158691);
DFFARX1 I_59635 (I1016503,I2683,I1016350,I1016342,);
not I_59636 (I1016534,I158688);
nand I_59637 (I1016551,I1016534,I158694);
nand I_59638 (I1016568,I1016452,I1016551);
and I_59639 (I1016321,I1016435,I1016568);
nor I_59640 (I1016599,I158688,I158706);
and I_59641 (I1016616,I1016435,I1016599);
nor I_59642 (I1016327,I1016401,I1016616);
DFFARX1 I_59643 (I1016599,I2683,I1016350,I1016656,);
not I_59644 (I1016664,I1016656);
nor I_59645 (I1016336,I1016435,I1016664);
or I_59646 (I1016695,I1016503,I158685);
nor I_59647 (I1016712,I158685,I158703);
nand I_59648 (I1016729,I1016568,I1016712);
nand I_59649 (I1016746,I1016695,I1016729);
DFFARX1 I_59650 (I1016746,I2683,I1016350,I1016339,);
nor I_59651 (I1016777,I1016712,I1016469);
DFFARX1 I_59652 (I1016777,I2683,I1016350,I1016318,);
nor I_59653 (I1016808,I158685,I158709);
DFFARX1 I_59654 (I1016808,I2683,I1016350,I1016834,);
DFFARX1 I_59655 (I1016834,I2683,I1016350,I1016333,);
not I_59656 (I1016856,I1016834);
nand I_59657 (I1016330,I1016856,I1016384);
nand I_59658 (I1016324,I1016856,I1016486);
not I_59659 (I1016928,I2690);
DFFARX1 I_59660 (I559562,I2683,I1016928,I1016954,);
nand I_59661 (I1016962,I1016954,I559565);
not I_59662 (I1016979,I1016962);
DFFARX1 I_59663 (I559577,I2683,I1016928,I1017005,);
not I_59664 (I1017013,I1017005);
not I_59665 (I1017030,I559562);
or I_59666 (I1017047,I559571,I559562);
nor I_59667 (I1017064,I559571,I559562);
or I_59668 (I1017081,I559580,I559571);
DFFARX1 I_59669 (I1017081,I2683,I1016928,I1016920,);
not I_59670 (I1017112,I559583);
nand I_59671 (I1017129,I1017112,I559565);
nand I_59672 (I1017146,I1017030,I1017129);
and I_59673 (I1016899,I1017013,I1017146);
nor I_59674 (I1017177,I559583,I559568);
and I_59675 (I1017194,I1017013,I1017177);
nor I_59676 (I1016905,I1016979,I1017194);
DFFARX1 I_59677 (I1017177,I2683,I1016928,I1017234,);
not I_59678 (I1017242,I1017234);
nor I_59679 (I1016914,I1017013,I1017242);
or I_59680 (I1017273,I1017081,I559574);
nor I_59681 (I1017290,I559574,I559580);
nand I_59682 (I1017307,I1017146,I1017290);
nand I_59683 (I1017324,I1017273,I1017307);
DFFARX1 I_59684 (I1017324,I2683,I1016928,I1016917,);
nor I_59685 (I1017355,I1017290,I1017047);
DFFARX1 I_59686 (I1017355,I2683,I1016928,I1016896,);
nor I_59687 (I1017386,I559574,I559586);
DFFARX1 I_59688 (I1017386,I2683,I1016928,I1017412,);
DFFARX1 I_59689 (I1017412,I2683,I1016928,I1016911,);
not I_59690 (I1017434,I1017412);
nand I_59691 (I1016908,I1017434,I1016962);
nand I_59692 (I1016902,I1017434,I1017064);
not I_59693 (I1017506,I2690);
DFFARX1 I_59694 (I441075,I2683,I1017506,I1017532,);
nand I_59695 (I1017540,I1017532,I441090);
not I_59696 (I1017557,I1017540);
DFFARX1 I_59697 (I441072,I2683,I1017506,I1017583,);
not I_59698 (I1017591,I1017583);
not I_59699 (I1017608,I441081);
or I_59700 (I1017625,I441075,I441081);
nor I_59701 (I1017642,I441075,I441081);
or I_59702 (I1017659,I441072,I441075);
DFFARX1 I_59703 (I1017659,I2683,I1017506,I1017498,);
not I_59704 (I1017690,I441093);
nand I_59705 (I1017707,I1017690,I441096);
nand I_59706 (I1017724,I1017608,I1017707);
and I_59707 (I1017477,I1017591,I1017724);
nor I_59708 (I1017755,I441093,I441078);
and I_59709 (I1017772,I1017591,I1017755);
nor I_59710 (I1017483,I1017557,I1017772);
DFFARX1 I_59711 (I1017755,I2683,I1017506,I1017812,);
not I_59712 (I1017820,I1017812);
nor I_59713 (I1017492,I1017591,I1017820);
or I_59714 (I1017851,I1017659,I441084);
nor I_59715 (I1017868,I441084,I441072);
nand I_59716 (I1017885,I1017724,I1017868);
nand I_59717 (I1017902,I1017851,I1017885);
DFFARX1 I_59718 (I1017902,I2683,I1017506,I1017495,);
nor I_59719 (I1017933,I1017868,I1017625);
DFFARX1 I_59720 (I1017933,I2683,I1017506,I1017474,);
nor I_59721 (I1017964,I441084,I441087);
DFFARX1 I_59722 (I1017964,I2683,I1017506,I1017990,);
DFFARX1 I_59723 (I1017990,I2683,I1017506,I1017489,);
not I_59724 (I1018012,I1017990);
nand I_59725 (I1017486,I1018012,I1017540);
nand I_59726 (I1017480,I1018012,I1017642);
not I_59727 (I1018084,I2690);
DFFARX1 I_59728 (I338293,I2683,I1018084,I1018110,);
nand I_59729 (I1018118,I1018110,I338302);
not I_59730 (I1018135,I1018118);
DFFARX1 I_59731 (I338290,I2683,I1018084,I1018161,);
not I_59732 (I1018169,I1018161);
not I_59733 (I1018186,I338296);
or I_59734 (I1018203,I338290,I338296);
nor I_59735 (I1018220,I338290,I338296);
or I_59736 (I1018237,I338305,I338290);
DFFARX1 I_59737 (I1018237,I2683,I1018084,I1018076,);
not I_59738 (I1018268,I338299);
nand I_59739 (I1018285,I1018268,I338314);
nand I_59740 (I1018302,I1018186,I1018285);
and I_59741 (I1018055,I1018169,I1018302);
nor I_59742 (I1018333,I338299,I338317);
and I_59743 (I1018350,I1018169,I1018333);
nor I_59744 (I1018061,I1018135,I1018350);
DFFARX1 I_59745 (I1018333,I2683,I1018084,I1018390,);
not I_59746 (I1018398,I1018390);
nor I_59747 (I1018070,I1018169,I1018398);
or I_59748 (I1018429,I1018237,I338308);
nor I_59749 (I1018446,I338308,I338305);
nand I_59750 (I1018463,I1018302,I1018446);
nand I_59751 (I1018480,I1018429,I1018463);
DFFARX1 I_59752 (I1018480,I2683,I1018084,I1018073,);
nor I_59753 (I1018511,I1018446,I1018203);
DFFARX1 I_59754 (I1018511,I2683,I1018084,I1018052,);
nor I_59755 (I1018542,I338308,I338311);
DFFARX1 I_59756 (I1018542,I2683,I1018084,I1018568,);
DFFARX1 I_59757 (I1018568,I2683,I1018084,I1018067,);
not I_59758 (I1018590,I1018568);
nand I_59759 (I1018064,I1018590,I1018118);
nand I_59760 (I1018058,I1018590,I1018220);
not I_59761 (I1018662,I2690);
DFFARX1 I_59762 (I1090003,I2683,I1018662,I1018688,);
nand I_59763 (I1018696,I1018688,I1089994);
not I_59764 (I1018713,I1018696);
DFFARX1 I_59765 (I1089979,I2683,I1018662,I1018739,);
not I_59766 (I1018747,I1018739);
not I_59767 (I1018764,I1089982);
or I_59768 (I1018781,I1089991,I1089982);
nor I_59769 (I1018798,I1089991,I1089982);
or I_59770 (I1018815,I1089988,I1089991);
DFFARX1 I_59771 (I1018815,I2683,I1018662,I1018654,);
not I_59772 (I1018846,I1090000);
nand I_59773 (I1018863,I1018846,I1089979);
nand I_59774 (I1018880,I1018764,I1018863);
and I_59775 (I1018633,I1018747,I1018880);
nor I_59776 (I1018911,I1090000,I1089985);
and I_59777 (I1018928,I1018747,I1018911);
nor I_59778 (I1018639,I1018713,I1018928);
DFFARX1 I_59779 (I1018911,I2683,I1018662,I1018968,);
not I_59780 (I1018976,I1018968);
nor I_59781 (I1018648,I1018747,I1018976);
or I_59782 (I1019007,I1018815,I1090006);
nor I_59783 (I1019024,I1090006,I1089988);
nand I_59784 (I1019041,I1018880,I1019024);
nand I_59785 (I1019058,I1019007,I1019041);
DFFARX1 I_59786 (I1019058,I2683,I1018662,I1018651,);
nor I_59787 (I1019089,I1019024,I1018781);
DFFARX1 I_59788 (I1019089,I2683,I1018662,I1018630,);
nor I_59789 (I1019120,I1090006,I1089997);
DFFARX1 I_59790 (I1019120,I2683,I1018662,I1019146,);
DFFARX1 I_59791 (I1019146,I2683,I1018662,I1018645,);
not I_59792 (I1019168,I1019146);
nand I_59793 (I1018642,I1019168,I1018696);
nand I_59794 (I1018636,I1019168,I1018798);
not I_59795 (I1019240,I2690);
DFFARX1 I_59796 (I504652,I2683,I1019240,I1019266,);
nand I_59797 (I1019274,I1019266,I504655);
not I_59798 (I1019291,I1019274);
DFFARX1 I_59799 (I504667,I2683,I1019240,I1019317,);
not I_59800 (I1019325,I1019317);
not I_59801 (I1019342,I504652);
or I_59802 (I1019359,I504661,I504652);
nor I_59803 (I1019376,I504661,I504652);
or I_59804 (I1019393,I504670,I504661);
DFFARX1 I_59805 (I1019393,I2683,I1019240,I1019232,);
not I_59806 (I1019424,I504673);
nand I_59807 (I1019441,I1019424,I504655);
nand I_59808 (I1019458,I1019342,I1019441);
and I_59809 (I1019211,I1019325,I1019458);
nor I_59810 (I1019489,I504673,I504658);
and I_59811 (I1019506,I1019325,I1019489);
nor I_59812 (I1019217,I1019291,I1019506);
DFFARX1 I_59813 (I1019489,I2683,I1019240,I1019546,);
not I_59814 (I1019554,I1019546);
nor I_59815 (I1019226,I1019325,I1019554);
or I_59816 (I1019585,I1019393,I504664);
nor I_59817 (I1019602,I504664,I504670);
nand I_59818 (I1019619,I1019458,I1019602);
nand I_59819 (I1019636,I1019585,I1019619);
DFFARX1 I_59820 (I1019636,I2683,I1019240,I1019229,);
nor I_59821 (I1019667,I1019602,I1019359);
DFFARX1 I_59822 (I1019667,I2683,I1019240,I1019208,);
nor I_59823 (I1019698,I504664,I504676);
DFFARX1 I_59824 (I1019698,I2683,I1019240,I1019724,);
DFFARX1 I_59825 (I1019724,I2683,I1019240,I1019223,);
not I_59826 (I1019746,I1019724);
nand I_59827 (I1019220,I1019746,I1019274);
nand I_59828 (I1019214,I1019746,I1019376);
not I_59829 (I1019818,I2690);
DFFARX1 I_59830 (I532974,I2683,I1019818,I1019844,);
nand I_59831 (I1019852,I1019844,I532977);
not I_59832 (I1019869,I1019852);
DFFARX1 I_59833 (I532989,I2683,I1019818,I1019895,);
not I_59834 (I1019903,I1019895);
not I_59835 (I1019920,I532974);
or I_59836 (I1019937,I532983,I532974);
nor I_59837 (I1019954,I532983,I532974);
or I_59838 (I1019971,I532992,I532983);
DFFARX1 I_59839 (I1019971,I2683,I1019818,I1019810,);
not I_59840 (I1020002,I532995);
nand I_59841 (I1020019,I1020002,I532977);
nand I_59842 (I1020036,I1019920,I1020019);
and I_59843 (I1019789,I1019903,I1020036);
nor I_59844 (I1020067,I532995,I532980);
and I_59845 (I1020084,I1019903,I1020067);
nor I_59846 (I1019795,I1019869,I1020084);
DFFARX1 I_59847 (I1020067,I2683,I1019818,I1020124,);
not I_59848 (I1020132,I1020124);
nor I_59849 (I1019804,I1019903,I1020132);
or I_59850 (I1020163,I1019971,I532986);
nor I_59851 (I1020180,I532986,I532992);
nand I_59852 (I1020197,I1020036,I1020180);
nand I_59853 (I1020214,I1020163,I1020197);
DFFARX1 I_59854 (I1020214,I2683,I1019818,I1019807,);
nor I_59855 (I1020245,I1020180,I1019937);
DFFARX1 I_59856 (I1020245,I2683,I1019818,I1019786,);
nor I_59857 (I1020276,I532986,I532998);
DFFARX1 I_59858 (I1020276,I2683,I1019818,I1020302,);
DFFARX1 I_59859 (I1020302,I2683,I1019818,I1019801,);
not I_59860 (I1020324,I1020302);
nand I_59861 (I1019798,I1020324,I1019852);
nand I_59862 (I1019792,I1020324,I1019954);
not I_59863 (I1020396,I2690);
DFFARX1 I_59864 (I270143,I2683,I1020396,I1020422,);
nand I_59865 (I1020430,I1020422,I270164);
not I_59866 (I1020447,I1020430);
DFFARX1 I_59867 (I270158,I2683,I1020396,I1020473,);
not I_59868 (I1020481,I1020473);
not I_59869 (I1020498,I270146);
or I_59870 (I1020515,I270161,I270146);
nor I_59871 (I1020532,I270161,I270146);
or I_59872 (I1020549,I270152,I270161);
DFFARX1 I_59873 (I1020549,I2683,I1020396,I1020388,);
not I_59874 (I1020580,I270140);
nand I_59875 (I1020597,I1020580,I270137);
nand I_59876 (I1020614,I1020498,I1020597);
and I_59877 (I1020367,I1020481,I1020614);
nor I_59878 (I1020645,I270140,I270149);
and I_59879 (I1020662,I1020481,I1020645);
nor I_59880 (I1020373,I1020447,I1020662);
DFFARX1 I_59881 (I1020645,I2683,I1020396,I1020702,);
not I_59882 (I1020710,I1020702);
nor I_59883 (I1020382,I1020481,I1020710);
or I_59884 (I1020741,I1020549,I270155);
nor I_59885 (I1020758,I270155,I270152);
nand I_59886 (I1020775,I1020614,I1020758);
nand I_59887 (I1020792,I1020741,I1020775);
DFFARX1 I_59888 (I1020792,I2683,I1020396,I1020385,);
nor I_59889 (I1020823,I1020758,I1020515);
DFFARX1 I_59890 (I1020823,I2683,I1020396,I1020364,);
nor I_59891 (I1020854,I270155,I270137);
DFFARX1 I_59892 (I1020854,I2683,I1020396,I1020880,);
DFFARX1 I_59893 (I1020880,I2683,I1020396,I1020379,);
not I_59894 (I1020902,I1020880);
nand I_59895 (I1020376,I1020902,I1020430);
nand I_59896 (I1020370,I1020902,I1020532);
not I_59897 (I1020977,I2690);
DFFARX1 I_59898 (I639652,I2683,I1020977,I1021003,);
nand I_59899 (I1021011,I1021003,I639670);
not I_59900 (I1021028,I1021011);
DFFARX1 I_59901 (I639649,I2683,I1020977,I1021054,);
not I_59902 (I1021062,I1021054);
nor I_59903 (I1021079,I639664,I639658);
not I_59904 (I1021096,I1021079);
DFFARX1 I_59905 (I1021096,I2683,I1020977,I1020963,);
or I_59906 (I1021127,I639655,I639664);
DFFARX1 I_59907 (I1021127,I2683,I1020977,I1020966,);
not I_59908 (I1021158,I639655);
nor I_59909 (I1021175,I1021158,I639661);
nor I_59910 (I1021192,I1021175,I639658);
nor I_59911 (I1021209,I639661,I639649);
nor I_59912 (I1021226,I1021062,I1021209);
nor I_59913 (I1020951,I1021028,I1021226);
not I_59914 (I1021257,I1021209);
nand I_59915 (I1020954,I1021257,I1021011);
nand I_59916 (I1020948,I1021257,I1021079);
nor I_59917 (I1020945,I1021209,I1021192);
nor I_59918 (I1021316,I639652,I639655);
not I_59919 (I1021333,I1021316);
DFFARX1 I_59920 (I1021316,I2683,I1020977,I1021359,);
not I_59921 (I1020969,I1021359);
nor I_59922 (I1021381,I639652,I639667);
DFFARX1 I_59923 (I1021381,I2683,I1020977,I1021407,);
and I_59924 (I1021415,I1021407,I639664);
nor I_59925 (I1021432,I1021415,I1021333);
DFFARX1 I_59926 (I1021432,I2683,I1020977,I1020960,);
nor I_59927 (I1021463,I1021407,I1021192);
DFFARX1 I_59928 (I1021463,I2683,I1020977,I1020942,);
nor I_59929 (I1020957,I1021407,I1021096);
not I_59930 (I1021538,I2690);
DFFARX1 I_59931 (I73301,I2683,I1021538,I1021564,);
nand I_59932 (I1021572,I1021564,I73292);
not I_59933 (I1021589,I1021572);
DFFARX1 I_59934 (I73280,I2683,I1021538,I1021615,);
not I_59935 (I1021623,I1021615);
nor I_59936 (I1021640,I73283,I73280);
not I_59937 (I1021657,I1021640);
DFFARX1 I_59938 (I1021657,I2683,I1021538,I1021524,);
or I_59939 (I1021688,I73277,I73283);
DFFARX1 I_59940 (I1021688,I2683,I1021538,I1021527,);
not I_59941 (I1021719,I73286);
nor I_59942 (I1021736,I1021719,I73277);
nor I_59943 (I1021753,I1021736,I73280);
nor I_59944 (I1021770,I73277,I73289);
nor I_59945 (I1021787,I1021623,I1021770);
nor I_59946 (I1021512,I1021589,I1021787);
not I_59947 (I1021818,I1021770);
nand I_59948 (I1021515,I1021818,I1021572);
nand I_59949 (I1021509,I1021818,I1021640);
nor I_59950 (I1021506,I1021770,I1021753);
nor I_59951 (I1021877,I73295,I73277);
not I_59952 (I1021894,I1021877);
DFFARX1 I_59953 (I1021877,I2683,I1021538,I1021920,);
not I_59954 (I1021530,I1021920);
nor I_59955 (I1021942,I73295,I73298);
DFFARX1 I_59956 (I1021942,I2683,I1021538,I1021968,);
and I_59957 (I1021976,I1021968,I73283);
nor I_59958 (I1021993,I1021976,I1021894);
DFFARX1 I_59959 (I1021993,I2683,I1021538,I1021521,);
nor I_59960 (I1022024,I1021968,I1021753);
DFFARX1 I_59961 (I1022024,I2683,I1021538,I1021503,);
nor I_59962 (I1021518,I1021968,I1021657);
not I_59963 (I1022099,I2690);
DFFARX1 I_59964 (I351911,I2683,I1022099,I1022125,);
nand I_59965 (I1022133,I1022125,I351893);
not I_59966 (I1022150,I1022133);
DFFARX1 I_59967 (I351890,I2683,I1022099,I1022176,);
not I_59968 (I1022184,I1022176);
nor I_59969 (I1022201,I351896,I351890);
not I_59970 (I1022218,I1022201);
DFFARX1 I_59971 (I1022218,I2683,I1022099,I1022085,);
or I_59972 (I1022249,I351899,I351896);
DFFARX1 I_59973 (I1022249,I2683,I1022099,I1022088,);
not I_59974 (I1022280,I351905);
nor I_59975 (I1022297,I1022280,I351917);
nor I_59976 (I1022314,I1022297,I351890);
nor I_59977 (I1022331,I351917,I351902);
nor I_59978 (I1022348,I1022184,I1022331);
nor I_59979 (I1022073,I1022150,I1022348);
not I_59980 (I1022379,I1022331);
nand I_59981 (I1022076,I1022379,I1022133);
nand I_59982 (I1022070,I1022379,I1022201);
nor I_59983 (I1022067,I1022331,I1022314);
nor I_59984 (I1022438,I351908,I351899);
not I_59985 (I1022455,I1022438);
DFFARX1 I_59986 (I1022438,I2683,I1022099,I1022481,);
not I_59987 (I1022091,I1022481);
nor I_59988 (I1022503,I351908,I351914);
DFFARX1 I_59989 (I1022503,I2683,I1022099,I1022529,);
and I_59990 (I1022537,I1022529,I351896);
nor I_59991 (I1022554,I1022537,I1022455);
DFFARX1 I_59992 (I1022554,I2683,I1022099,I1022082,);
nor I_59993 (I1022585,I1022529,I1022314);
DFFARX1 I_59994 (I1022585,I2683,I1022099,I1022064,);
nor I_59995 (I1022079,I1022529,I1022218);
not I_59996 (I1022660,I2690);
DFFARX1 I_59997 (I546864,I2683,I1022660,I1022686,);
nand I_59998 (I1022694,I1022686,I546849);
not I_59999 (I1022711,I1022694);
DFFARX1 I_60000 (I546867,I2683,I1022660,I1022737,);
not I_60001 (I1022745,I1022737);
nor I_60002 (I1022762,I546846,I546861);
not I_60003 (I1022779,I1022762);
DFFARX1 I_60004 (I1022779,I2683,I1022660,I1022646,);
or I_60005 (I1022810,I546858,I546846);
DFFARX1 I_60006 (I1022810,I2683,I1022660,I1022649,);
not I_60007 (I1022841,I546846);
nor I_60008 (I1022858,I1022841,I546855);
nor I_60009 (I1022875,I1022858,I546861);
nor I_60010 (I1022892,I546855,I546849);
nor I_60011 (I1022909,I1022745,I1022892);
nor I_60012 (I1022634,I1022711,I1022909);
not I_60013 (I1022940,I1022892);
nand I_60014 (I1022637,I1022940,I1022694);
nand I_60015 (I1022631,I1022940,I1022762);
nor I_60016 (I1022628,I1022892,I1022875);
nor I_60017 (I1022999,I546852,I546858);
not I_60018 (I1023016,I1022999);
DFFARX1 I_60019 (I1022999,I2683,I1022660,I1023042,);
not I_60020 (I1022652,I1023042);
nor I_60021 (I1023064,I546852,I546870);
DFFARX1 I_60022 (I1023064,I2683,I1022660,I1023090,);
and I_60023 (I1023098,I1023090,I546846);
nor I_60024 (I1023115,I1023098,I1023016);
DFFARX1 I_60025 (I1023115,I2683,I1022660,I1022643,);
nor I_60026 (I1023146,I1023090,I1022875);
DFFARX1 I_60027 (I1023146,I2683,I1022660,I1022625,);
nor I_60028 (I1022640,I1023090,I1022779);
not I_60029 (I1023221,I2690);
DFFARX1 I_60030 (I321991,I2683,I1023221,I1023247,);
nand I_60031 (I1023255,I1023247,I321973);
not I_60032 (I1023272,I1023255);
DFFARX1 I_60033 (I321970,I2683,I1023221,I1023298,);
not I_60034 (I1023306,I1023298);
nor I_60035 (I1023323,I321976,I321970);
not I_60036 (I1023340,I1023323);
DFFARX1 I_60037 (I1023340,I2683,I1023221,I1023207,);
or I_60038 (I1023371,I321979,I321976);
DFFARX1 I_60039 (I1023371,I2683,I1023221,I1023210,);
not I_60040 (I1023402,I321985);
nor I_60041 (I1023419,I1023402,I321997);
nor I_60042 (I1023436,I1023419,I321970);
nor I_60043 (I1023453,I321997,I321982);
nor I_60044 (I1023470,I1023306,I1023453);
nor I_60045 (I1023195,I1023272,I1023470);
not I_60046 (I1023501,I1023453);
nand I_60047 (I1023198,I1023501,I1023255);
nand I_60048 (I1023192,I1023501,I1023323);
nor I_60049 (I1023189,I1023453,I1023436);
nor I_60050 (I1023560,I321988,I321979);
not I_60051 (I1023577,I1023560);
DFFARX1 I_60052 (I1023560,I2683,I1023221,I1023603,);
not I_60053 (I1023213,I1023603);
nor I_60054 (I1023625,I321988,I321994);
DFFARX1 I_60055 (I1023625,I2683,I1023221,I1023651,);
and I_60056 (I1023659,I1023651,I321976);
nor I_60057 (I1023676,I1023659,I1023577);
DFFARX1 I_60058 (I1023676,I2683,I1023221,I1023204,);
nor I_60059 (I1023707,I1023651,I1023436);
DFFARX1 I_60060 (I1023707,I2683,I1023221,I1023186,);
nor I_60061 (I1023201,I1023651,I1023340);
not I_60062 (I1023782,I2690);
DFFARX1 I_60063 (I862879,I2683,I1023782,I1023808,);
nand I_60064 (I1023816,I1023808,I862876);
not I_60065 (I1023833,I1023816);
DFFARX1 I_60066 (I862879,I2683,I1023782,I1023859,);
not I_60067 (I1023867,I1023859);
nor I_60068 (I1023884,I862897,I862891);
not I_60069 (I1023901,I1023884);
DFFARX1 I_60070 (I1023901,I2683,I1023782,I1023768,);
or I_60071 (I1023932,I862900,I862897);
DFFARX1 I_60072 (I1023932,I2683,I1023782,I1023771,);
not I_60073 (I1023963,I862888);
nor I_60074 (I1023980,I1023963,I862885);
nor I_60075 (I1023997,I1023980,I862891);
nor I_60076 (I1024014,I862885,I862876);
nor I_60077 (I1024031,I1023867,I1024014);
nor I_60078 (I1023756,I1023833,I1024031);
not I_60079 (I1024062,I1024014);
nand I_60080 (I1023759,I1024062,I1023816);
nand I_60081 (I1023753,I1024062,I1023884);
nor I_60082 (I1023750,I1024014,I1023997);
nor I_60083 (I1024121,I862882,I862900);
not I_60084 (I1024138,I1024121);
DFFARX1 I_60085 (I1024121,I2683,I1023782,I1024164,);
not I_60086 (I1023774,I1024164);
nor I_60087 (I1024186,I862882,I862894);
DFFARX1 I_60088 (I1024186,I2683,I1023782,I1024212,);
and I_60089 (I1024220,I1024212,I862897);
nor I_60090 (I1024237,I1024220,I1024138);
DFFARX1 I_60091 (I1024237,I2683,I1023782,I1023765,);
nor I_60092 (I1024268,I1024212,I1023997);
DFFARX1 I_60093 (I1024268,I2683,I1023782,I1023747,);
nor I_60094 (I1023762,I1024212,I1023901);
not I_60095 (I1024343,I2690);
DFFARX1 I_60096 (I700635,I2683,I1024343,I1024369,);
nand I_60097 (I1024377,I1024369,I700617);
not I_60098 (I1024394,I1024377);
DFFARX1 I_60099 (I700629,I2683,I1024343,I1024420,);
not I_60100 (I1024428,I1024420);
nor I_60101 (I1024445,I700611,I700611);
not I_60102 (I1024462,I1024445);
DFFARX1 I_60103 (I1024462,I2683,I1024343,I1024329,);
or I_60104 (I1024493,I700623,I700611);
DFFARX1 I_60105 (I1024493,I2683,I1024343,I1024332,);
not I_60106 (I1024524,I700638);
nor I_60107 (I1024541,I1024524,I700626);
nor I_60108 (I1024558,I1024541,I700611);
nor I_60109 (I1024575,I700626,I700614);
nor I_60110 (I1024592,I1024428,I1024575);
nor I_60111 (I1024317,I1024394,I1024592);
not I_60112 (I1024623,I1024575);
nand I_60113 (I1024320,I1024623,I1024377);
nand I_60114 (I1024314,I1024623,I1024445);
nor I_60115 (I1024311,I1024575,I1024558);
nor I_60116 (I1024682,I700620,I700623);
not I_60117 (I1024699,I1024682);
DFFARX1 I_60118 (I1024682,I2683,I1024343,I1024725,);
not I_60119 (I1024335,I1024725);
nor I_60120 (I1024747,I700620,I700632);
DFFARX1 I_60121 (I1024747,I2683,I1024343,I1024773,);
and I_60122 (I1024781,I1024773,I700611);
nor I_60123 (I1024798,I1024781,I1024699);
DFFARX1 I_60124 (I1024798,I2683,I1024343,I1024326,);
nor I_60125 (I1024829,I1024773,I1024558);
DFFARX1 I_60126 (I1024829,I2683,I1024343,I1024308,);
nor I_60127 (I1024323,I1024773,I1024462);
not I_60128 (I1024904,I2690);
DFFARX1 I_60129 (I292292,I2683,I1024904,I1024930,);
nand I_60130 (I1024938,I1024930,I292271);
not I_60131 (I1024955,I1024938);
DFFARX1 I_60132 (I292280,I2683,I1024904,I1024981,);
not I_60133 (I1024989,I1024981);
nor I_60134 (I1025006,I292274,I292286);
not I_60135 (I1025023,I1025006);
DFFARX1 I_60136 (I1025023,I2683,I1024904,I1024890,);
or I_60137 (I1025054,I292277,I292274);
DFFARX1 I_60138 (I1025054,I2683,I1024904,I1024893,);
not I_60139 (I1025085,I292298);
nor I_60140 (I1025102,I1025085,I292283);
nor I_60141 (I1025119,I1025102,I292286);
nor I_60142 (I1025136,I292283,I292271);
nor I_60143 (I1025153,I1024989,I1025136);
nor I_60144 (I1024878,I1024955,I1025153);
not I_60145 (I1025184,I1025136);
nand I_60146 (I1024881,I1025184,I1024938);
nand I_60147 (I1024875,I1025184,I1025006);
nor I_60148 (I1024872,I1025136,I1025119);
nor I_60149 (I1025243,I292289,I292277);
not I_60150 (I1025260,I1025243);
DFFARX1 I_60151 (I1025243,I2683,I1024904,I1025286,);
not I_60152 (I1024896,I1025286);
nor I_60153 (I1025308,I292289,I292295);
DFFARX1 I_60154 (I1025308,I2683,I1024904,I1025334,);
and I_60155 (I1025342,I1025334,I292274);
nor I_60156 (I1025359,I1025342,I1025260);
DFFARX1 I_60157 (I1025359,I2683,I1024904,I1024887,);
nor I_60158 (I1025390,I1025334,I1025119);
DFFARX1 I_60159 (I1025390,I2683,I1024904,I1024869,);
nor I_60160 (I1024884,I1025334,I1025023);
not I_60161 (I1025465,I2690);
DFFARX1 I_60162 (I65923,I2683,I1025465,I1025491,);
nand I_60163 (I1025499,I1025491,I65914);
not I_60164 (I1025516,I1025499);
DFFARX1 I_60165 (I65902,I2683,I1025465,I1025542,);
not I_60166 (I1025550,I1025542);
nor I_60167 (I1025567,I65905,I65902);
not I_60168 (I1025584,I1025567);
DFFARX1 I_60169 (I1025584,I2683,I1025465,I1025451,);
or I_60170 (I1025615,I65899,I65905);
DFFARX1 I_60171 (I1025615,I2683,I1025465,I1025454,);
not I_60172 (I1025646,I65908);
nor I_60173 (I1025663,I1025646,I65899);
nor I_60174 (I1025680,I1025663,I65902);
nor I_60175 (I1025697,I65899,I65911);
nor I_60176 (I1025714,I1025550,I1025697);
nor I_60177 (I1025439,I1025516,I1025714);
not I_60178 (I1025745,I1025697);
nand I_60179 (I1025442,I1025745,I1025499);
nand I_60180 (I1025436,I1025745,I1025567);
nor I_60181 (I1025433,I1025697,I1025680);
nor I_60182 (I1025804,I65917,I65899);
not I_60183 (I1025821,I1025804);
DFFARX1 I_60184 (I1025804,I2683,I1025465,I1025847,);
not I_60185 (I1025457,I1025847);
nor I_60186 (I1025869,I65917,I65920);
DFFARX1 I_60187 (I1025869,I2683,I1025465,I1025895,);
and I_60188 (I1025903,I1025895,I65905);
nor I_60189 (I1025920,I1025903,I1025821);
DFFARX1 I_60190 (I1025920,I2683,I1025465,I1025448,);
nor I_60191 (I1025951,I1025895,I1025680);
DFFARX1 I_60192 (I1025951,I2683,I1025465,I1025430,);
nor I_60193 (I1025445,I1025895,I1025584);
not I_60194 (I1026026,I2690);
DFFARX1 I_60195 (I795597,I2683,I1026026,I1026052,);
nand I_60196 (I1026060,I1026052,I795579);
not I_60197 (I1026077,I1026060);
DFFARX1 I_60198 (I795591,I2683,I1026026,I1026103,);
not I_60199 (I1026111,I1026103);
nor I_60200 (I1026128,I795573,I795573);
not I_60201 (I1026145,I1026128);
DFFARX1 I_60202 (I1026145,I2683,I1026026,I1026012,);
or I_60203 (I1026176,I795585,I795573);
DFFARX1 I_60204 (I1026176,I2683,I1026026,I1026015,);
not I_60205 (I1026207,I795600);
nor I_60206 (I1026224,I1026207,I795588);
nor I_60207 (I1026241,I1026224,I795573);
nor I_60208 (I1026258,I795588,I795576);
nor I_60209 (I1026275,I1026111,I1026258);
nor I_60210 (I1026000,I1026077,I1026275);
not I_60211 (I1026306,I1026258);
nand I_60212 (I1026003,I1026306,I1026060);
nand I_60213 (I1025997,I1026306,I1026128);
nor I_60214 (I1025994,I1026258,I1026241);
nor I_60215 (I1026365,I795582,I795585);
not I_60216 (I1026382,I1026365);
DFFARX1 I_60217 (I1026365,I2683,I1026026,I1026408,);
not I_60218 (I1026018,I1026408);
nor I_60219 (I1026430,I795582,I795594);
DFFARX1 I_60220 (I1026430,I2683,I1026026,I1026456,);
and I_60221 (I1026464,I1026456,I795573);
nor I_60222 (I1026481,I1026464,I1026382);
DFFARX1 I_60223 (I1026481,I2683,I1026026,I1026009,);
nor I_60224 (I1026512,I1026456,I1026241);
DFFARX1 I_60225 (I1026512,I2683,I1026026,I1025991,);
nor I_60226 (I1026006,I1026456,I1026145);
not I_60227 (I1026587,I2690);
DFFARX1 I_60228 (I1001299,I2683,I1026587,I1026613,);
nand I_60229 (I1026621,I1026613,I1001302);
not I_60230 (I1026638,I1026621);
DFFARX1 I_60231 (I1001308,I2683,I1026587,I1026664,);
not I_60232 (I1026672,I1026664);
nor I_60233 (I1026689,I1001305,I1001290);
not I_60234 (I1026706,I1026689);
DFFARX1 I_60235 (I1026706,I2683,I1026587,I1026573,);
or I_60236 (I1026737,I1001314,I1001305);
DFFARX1 I_60237 (I1026737,I2683,I1026587,I1026576,);
not I_60238 (I1026768,I1001293);
nor I_60239 (I1026785,I1026768,I1001296);
nor I_60240 (I1026802,I1026785,I1001290);
nor I_60241 (I1026819,I1001296,I1001290);
nor I_60242 (I1026836,I1026672,I1026819);
nor I_60243 (I1026561,I1026638,I1026836);
not I_60244 (I1026867,I1026819);
nand I_60245 (I1026564,I1026867,I1026621);
nand I_60246 (I1026558,I1026867,I1026689);
nor I_60247 (I1026555,I1026819,I1026802);
nor I_60248 (I1026926,I1001293,I1001314);
not I_60249 (I1026943,I1026926);
DFFARX1 I_60250 (I1026926,I2683,I1026587,I1026969,);
not I_60251 (I1026579,I1026969);
nor I_60252 (I1026991,I1001293,I1001311);
DFFARX1 I_60253 (I1026991,I2683,I1026587,I1027017,);
and I_60254 (I1027025,I1027017,I1001305);
nor I_60255 (I1027042,I1027025,I1026943);
DFFARX1 I_60256 (I1027042,I2683,I1026587,I1026570,);
nor I_60257 (I1027073,I1027017,I1026802);
DFFARX1 I_60258 (I1027073,I2683,I1026587,I1026552,);
nor I_60259 (I1026567,I1027017,I1026706);
not I_60260 (I1027148,I2690);
DFFARX1 I_60261 (I870971,I2683,I1027148,I1027174,);
nand I_60262 (I1027182,I1027174,I870968);
not I_60263 (I1027199,I1027182);
DFFARX1 I_60264 (I870971,I2683,I1027148,I1027225,);
not I_60265 (I1027233,I1027225);
nor I_60266 (I1027250,I870989,I870983);
not I_60267 (I1027267,I1027250);
DFFARX1 I_60268 (I1027267,I2683,I1027148,I1027134,);
or I_60269 (I1027298,I870992,I870989);
DFFARX1 I_60270 (I1027298,I2683,I1027148,I1027137,);
not I_60271 (I1027329,I870980);
nor I_60272 (I1027346,I1027329,I870977);
nor I_60273 (I1027363,I1027346,I870983);
nor I_60274 (I1027380,I870977,I870968);
nor I_60275 (I1027397,I1027233,I1027380);
nor I_60276 (I1027122,I1027199,I1027397);
not I_60277 (I1027428,I1027380);
nand I_60278 (I1027125,I1027428,I1027182);
nand I_60279 (I1027119,I1027428,I1027250);
nor I_60280 (I1027116,I1027380,I1027363);
nor I_60281 (I1027487,I870974,I870992);
not I_60282 (I1027504,I1027487);
DFFARX1 I_60283 (I1027487,I2683,I1027148,I1027530,);
not I_60284 (I1027140,I1027530);
nor I_60285 (I1027552,I870974,I870986);
DFFARX1 I_60286 (I1027552,I2683,I1027148,I1027578,);
and I_60287 (I1027586,I1027578,I870989);
nor I_60288 (I1027603,I1027586,I1027504);
DFFARX1 I_60289 (I1027603,I2683,I1027148,I1027131,);
nor I_60290 (I1027634,I1027578,I1027363);
DFFARX1 I_60291 (I1027634,I2683,I1027148,I1027113,);
nor I_60292 (I1027128,I1027578,I1027267);
not I_60293 (I1027709,I2690);
DFFARX1 I_60294 (I998987,I2683,I1027709,I1027735,);
nand I_60295 (I1027743,I1027735,I998990);
not I_60296 (I1027760,I1027743);
DFFARX1 I_60297 (I998996,I2683,I1027709,I1027786,);
not I_60298 (I1027794,I1027786);
nor I_60299 (I1027811,I998993,I998978);
not I_60300 (I1027828,I1027811);
DFFARX1 I_60301 (I1027828,I2683,I1027709,I1027695,);
or I_60302 (I1027859,I999002,I998993);
DFFARX1 I_60303 (I1027859,I2683,I1027709,I1027698,);
not I_60304 (I1027890,I998981);
nor I_60305 (I1027907,I1027890,I998984);
nor I_60306 (I1027924,I1027907,I998978);
nor I_60307 (I1027941,I998984,I998978);
nor I_60308 (I1027958,I1027794,I1027941);
nor I_60309 (I1027683,I1027760,I1027958);
not I_60310 (I1027989,I1027941);
nand I_60311 (I1027686,I1027989,I1027743);
nand I_60312 (I1027680,I1027989,I1027811);
nor I_60313 (I1027677,I1027941,I1027924);
nor I_60314 (I1028048,I998981,I999002);
not I_60315 (I1028065,I1028048);
DFFARX1 I_60316 (I1028048,I2683,I1027709,I1028091,);
not I_60317 (I1027701,I1028091);
nor I_60318 (I1028113,I998981,I998999);
DFFARX1 I_60319 (I1028113,I2683,I1027709,I1028139,);
and I_60320 (I1028147,I1028139,I998993);
nor I_60321 (I1028164,I1028147,I1028065);
DFFARX1 I_60322 (I1028164,I2683,I1027709,I1027692,);
nor I_60323 (I1028195,I1028139,I1027924);
DFFARX1 I_60324 (I1028195,I2683,I1027709,I1027674,);
nor I_60325 (I1027689,I1028139,I1027828);
not I_60326 (I1028270,I2690);
DFFARX1 I_60327 (I940909,I2683,I1028270,I1028296,);
nand I_60328 (I1028304,I1028296,I940906);
not I_60329 (I1028321,I1028304);
DFFARX1 I_60330 (I940909,I2683,I1028270,I1028347,);
not I_60331 (I1028355,I1028347);
nor I_60332 (I1028372,I940927,I940921);
not I_60333 (I1028389,I1028372);
DFFARX1 I_60334 (I1028389,I2683,I1028270,I1028256,);
or I_60335 (I1028420,I940930,I940927);
DFFARX1 I_60336 (I1028420,I2683,I1028270,I1028259,);
not I_60337 (I1028451,I940918);
nor I_60338 (I1028468,I1028451,I940915);
nor I_60339 (I1028485,I1028468,I940921);
nor I_60340 (I1028502,I940915,I940906);
nor I_60341 (I1028519,I1028355,I1028502);
nor I_60342 (I1028244,I1028321,I1028519);
not I_60343 (I1028550,I1028502);
nand I_60344 (I1028247,I1028550,I1028304);
nand I_60345 (I1028241,I1028550,I1028372);
nor I_60346 (I1028238,I1028502,I1028485);
nor I_60347 (I1028609,I940912,I940930);
not I_60348 (I1028626,I1028609);
DFFARX1 I_60349 (I1028609,I2683,I1028270,I1028652,);
not I_60350 (I1028262,I1028652);
nor I_60351 (I1028674,I940912,I940924);
DFFARX1 I_60352 (I1028674,I2683,I1028270,I1028700,);
and I_60353 (I1028708,I1028700,I940927);
nor I_60354 (I1028725,I1028708,I1028626);
DFFARX1 I_60355 (I1028725,I2683,I1028270,I1028253,);
nor I_60356 (I1028756,I1028700,I1028485);
DFFARX1 I_60357 (I1028756,I2683,I1028270,I1028235,);
nor I_60358 (I1028250,I1028700,I1028389);
not I_60359 (I1028831,I2690);
DFFARX1 I_60360 (I323623,I2683,I1028831,I1028857,);
nand I_60361 (I1028865,I1028857,I323605);
not I_60362 (I1028882,I1028865);
DFFARX1 I_60363 (I323602,I2683,I1028831,I1028908,);
not I_60364 (I1028916,I1028908);
nor I_60365 (I1028933,I323608,I323602);
not I_60366 (I1028950,I1028933);
DFFARX1 I_60367 (I1028950,I2683,I1028831,I1028817,);
or I_60368 (I1028981,I323611,I323608);
DFFARX1 I_60369 (I1028981,I2683,I1028831,I1028820,);
not I_60370 (I1029012,I323617);
nor I_60371 (I1029029,I1029012,I323629);
nor I_60372 (I1029046,I1029029,I323602);
nor I_60373 (I1029063,I323629,I323614);
nor I_60374 (I1029080,I1028916,I1029063);
nor I_60375 (I1028805,I1028882,I1029080);
not I_60376 (I1029111,I1029063);
nand I_60377 (I1028808,I1029111,I1028865);
nand I_60378 (I1028802,I1029111,I1028933);
nor I_60379 (I1028799,I1029063,I1029046);
nor I_60380 (I1029170,I323620,I323611);
not I_60381 (I1029187,I1029170);
DFFARX1 I_60382 (I1029170,I2683,I1028831,I1029213,);
not I_60383 (I1028823,I1029213);
nor I_60384 (I1029235,I323620,I323626);
DFFARX1 I_60385 (I1029235,I2683,I1028831,I1029261,);
and I_60386 (I1029269,I1029261,I323608);
nor I_60387 (I1029286,I1029269,I1029187);
DFFARX1 I_60388 (I1029286,I2683,I1028831,I1028814,);
nor I_60389 (I1029317,I1029261,I1029046);
DFFARX1 I_60390 (I1029317,I2683,I1028831,I1028796,);
nor I_60391 (I1028811,I1029261,I1028950);
not I_60392 (I1029392,I2690);
DFFARX1 I_60393 (I450344,I2683,I1029392,I1029418,);
nand I_60394 (I1029426,I1029418,I450323);
not I_60395 (I1029443,I1029426);
DFFARX1 I_60396 (I450335,I2683,I1029392,I1029469,);
not I_60397 (I1029477,I1029469);
nor I_60398 (I1029494,I450323,I450332);
not I_60399 (I1029511,I1029494);
DFFARX1 I_60400 (I1029511,I2683,I1029392,I1029378,);
or I_60401 (I1029542,I450326,I450323);
DFFARX1 I_60402 (I1029542,I2683,I1029392,I1029381,);
not I_60403 (I1029573,I450329);
nor I_60404 (I1029590,I1029573,I450320);
nor I_60405 (I1029607,I1029590,I450332);
nor I_60406 (I1029624,I450320,I450338);
nor I_60407 (I1029641,I1029477,I1029624);
nor I_60408 (I1029366,I1029443,I1029641);
not I_60409 (I1029672,I1029624);
nand I_60410 (I1029369,I1029672,I1029426);
nand I_60411 (I1029363,I1029672,I1029494);
nor I_60412 (I1029360,I1029624,I1029607);
nor I_60413 (I1029731,I450341,I450326);
not I_60414 (I1029748,I1029731);
DFFARX1 I_60415 (I1029731,I2683,I1029392,I1029774,);
not I_60416 (I1029384,I1029774);
nor I_60417 (I1029796,I450341,I450320);
DFFARX1 I_60418 (I1029796,I2683,I1029392,I1029822,);
and I_60419 (I1029830,I1029822,I450323);
nor I_60420 (I1029847,I1029830,I1029748);
DFFARX1 I_60421 (I1029847,I2683,I1029392,I1029375,);
nor I_60422 (I1029878,I1029822,I1029607);
DFFARX1 I_60423 (I1029878,I2683,I1029392,I1029357,);
nor I_60424 (I1029372,I1029822,I1029511);
not I_60425 (I1029953,I2690);
DFFARX1 I_60426 (I439940,I2683,I1029953,I1029979,);
nand I_60427 (I1029987,I1029979,I439919);
not I_60428 (I1030004,I1029987);
DFFARX1 I_60429 (I439931,I2683,I1029953,I1030030,);
not I_60430 (I1030038,I1030030);
nor I_60431 (I1030055,I439919,I439928);
not I_60432 (I1030072,I1030055);
DFFARX1 I_60433 (I1030072,I2683,I1029953,I1029939,);
or I_60434 (I1030103,I439922,I439919);
DFFARX1 I_60435 (I1030103,I2683,I1029953,I1029942,);
not I_60436 (I1030134,I439925);
nor I_60437 (I1030151,I1030134,I439916);
nor I_60438 (I1030168,I1030151,I439928);
nor I_60439 (I1030185,I439916,I439934);
nor I_60440 (I1030202,I1030038,I1030185);
nor I_60441 (I1029927,I1030004,I1030202);
not I_60442 (I1030233,I1030185);
nand I_60443 (I1029930,I1030233,I1029987);
nand I_60444 (I1029924,I1030233,I1030055);
nor I_60445 (I1029921,I1030185,I1030168);
nor I_60446 (I1030292,I439937,I439922);
not I_60447 (I1030309,I1030292);
DFFARX1 I_60448 (I1030292,I2683,I1029953,I1030335,);
not I_60449 (I1029945,I1030335);
nor I_60450 (I1030357,I439937,I439916);
DFFARX1 I_60451 (I1030357,I2683,I1029953,I1030383,);
and I_60452 (I1030391,I1030383,I439919);
nor I_60453 (I1030408,I1030391,I1030309);
DFFARX1 I_60454 (I1030408,I2683,I1029953,I1029936,);
nor I_60455 (I1030439,I1030383,I1030168);
DFFARX1 I_60456 (I1030439,I2683,I1029953,I1029918,);
nor I_60457 (I1029933,I1030383,I1030072);
not I_60458 (I1030514,I2690);
DFFARX1 I_60459 (I370386,I2683,I1030514,I1030540,);
DFFARX1 I_60460 (I370392,I2683,I1030514,I1030557,);
not I_60461 (I1030565,I1030557);
nor I_60462 (I1030482,I1030540,I1030565);
DFFARX1 I_60463 (I1030565,I2683,I1030514,I1030497,);
nor I_60464 (I1030610,I370401,I370386);
and I_60465 (I1030627,I1030610,I370413);
nor I_60466 (I1030644,I1030627,I370401);
not I_60467 (I1030661,I370401);
and I_60468 (I1030678,I1030661,I370389);
nand I_60469 (I1030695,I1030678,I370410);
nor I_60470 (I1030712,I1030661,I1030695);
DFFARX1 I_60471 (I1030712,I2683,I1030514,I1030479,);
not I_60472 (I1030743,I1030695);
nand I_60473 (I1030760,I1030565,I1030743);
nand I_60474 (I1030491,I1030627,I1030743);
DFFARX1 I_60475 (I1030661,I2683,I1030514,I1030506,);
not I_60476 (I1030805,I370398);
nor I_60477 (I1030822,I1030805,I370389);
nor I_60478 (I1030839,I1030822,I1030644);
DFFARX1 I_60479 (I1030839,I2683,I1030514,I1030503,);
not I_60480 (I1030870,I1030822);
DFFARX1 I_60481 (I1030870,I2683,I1030514,I1030896,);
not I_60482 (I1030904,I1030896);
nor I_60483 (I1030500,I1030904,I1030822);
nor I_60484 (I1030935,I1030805,I370395);
and I_60485 (I1030952,I1030935,I370407);
or I_60486 (I1030969,I1030952,I370404);
DFFARX1 I_60487 (I1030969,I2683,I1030514,I1030995,);
not I_60488 (I1031003,I1030995);
nand I_60489 (I1031020,I1031003,I1030743);
not I_60490 (I1030494,I1031020);
nand I_60491 (I1030488,I1031020,I1030760);
nand I_60492 (I1030485,I1031003,I1030627);
not I_60493 (I1031109,I2690);
DFFARX1 I_60494 (I868659,I2683,I1031109,I1031135,);
DFFARX1 I_60495 (I868671,I2683,I1031109,I1031152,);
not I_60496 (I1031160,I1031152);
nor I_60497 (I1031077,I1031135,I1031160);
DFFARX1 I_60498 (I1031160,I2683,I1031109,I1031092,);
nor I_60499 (I1031205,I868668,I868662);
and I_60500 (I1031222,I1031205,I868656);
nor I_60501 (I1031239,I1031222,I868668);
not I_60502 (I1031256,I868668);
and I_60503 (I1031273,I1031256,I868665);
nand I_60504 (I1031290,I1031273,I868656);
nor I_60505 (I1031307,I1031256,I1031290);
DFFARX1 I_60506 (I1031307,I2683,I1031109,I1031074,);
not I_60507 (I1031338,I1031290);
nand I_60508 (I1031355,I1031160,I1031338);
nand I_60509 (I1031086,I1031222,I1031338);
DFFARX1 I_60510 (I1031256,I2683,I1031109,I1031101,);
not I_60511 (I1031400,I868680);
nor I_60512 (I1031417,I1031400,I868665);
nor I_60513 (I1031434,I1031417,I1031239);
DFFARX1 I_60514 (I1031434,I2683,I1031109,I1031098,);
not I_60515 (I1031465,I1031417);
DFFARX1 I_60516 (I1031465,I2683,I1031109,I1031491,);
not I_60517 (I1031499,I1031491);
nor I_60518 (I1031095,I1031499,I1031417);
nor I_60519 (I1031530,I1031400,I868674);
and I_60520 (I1031547,I1031530,I868677);
or I_60521 (I1031564,I1031547,I868659);
DFFARX1 I_60522 (I1031564,I2683,I1031109,I1031590,);
not I_60523 (I1031598,I1031590);
nand I_60524 (I1031615,I1031598,I1031338);
not I_60525 (I1031089,I1031615);
nand I_60526 (I1031083,I1031615,I1031355);
nand I_60527 (I1031080,I1031598,I1031222);
not I_60528 (I1031704,I2690);
DFFARX1 I_60529 (I516233,I2683,I1031704,I1031730,);
DFFARX1 I_60530 (I516215,I2683,I1031704,I1031747,);
not I_60531 (I1031755,I1031747);
nor I_60532 (I1031672,I1031730,I1031755);
DFFARX1 I_60533 (I1031755,I2683,I1031704,I1031687,);
nor I_60534 (I1031800,I516221,I516224);
and I_60535 (I1031817,I1031800,I516212);
nor I_60536 (I1031834,I1031817,I516221);
not I_60537 (I1031851,I516221);
and I_60538 (I1031868,I1031851,I516230);
nand I_60539 (I1031885,I1031868,I516218);
nor I_60540 (I1031902,I1031851,I1031885);
DFFARX1 I_60541 (I1031902,I2683,I1031704,I1031669,);
not I_60542 (I1031933,I1031885);
nand I_60543 (I1031950,I1031755,I1031933);
nand I_60544 (I1031681,I1031817,I1031933);
DFFARX1 I_60545 (I1031851,I2683,I1031704,I1031696,);
not I_60546 (I1031995,I516215);
nor I_60547 (I1032012,I1031995,I516230);
nor I_60548 (I1032029,I1032012,I1031834);
DFFARX1 I_60549 (I1032029,I2683,I1031704,I1031693,);
not I_60550 (I1032060,I1032012);
DFFARX1 I_60551 (I1032060,I2683,I1031704,I1032086,);
not I_60552 (I1032094,I1032086);
nor I_60553 (I1031690,I1032094,I1032012);
nor I_60554 (I1032125,I1031995,I516227);
and I_60555 (I1032142,I1032125,I516236);
or I_60556 (I1032159,I1032142,I516212);
DFFARX1 I_60557 (I1032159,I2683,I1031704,I1032185,);
not I_60558 (I1032193,I1032185);
nand I_60559 (I1032210,I1032193,I1031933);
not I_60560 (I1031684,I1032210);
nand I_60561 (I1031678,I1032210,I1031950);
nand I_60562 (I1031675,I1032193,I1031817);
not I_60563 (I1032299,I2690);
DFFARX1 I_60564 (I233795,I2683,I1032299,I1032325,);
DFFARX1 I_60565 (I233789,I2683,I1032299,I1032342,);
not I_60566 (I1032350,I1032342);
nor I_60567 (I1032267,I1032325,I1032350);
DFFARX1 I_60568 (I1032350,I2683,I1032299,I1032282,);
nor I_60569 (I1032395,I233777,I233798);
and I_60570 (I1032412,I1032395,I233792);
nor I_60571 (I1032429,I1032412,I233777);
not I_60572 (I1032446,I233777);
and I_60573 (I1032463,I1032446,I233774);
nand I_60574 (I1032480,I1032463,I233786);
nor I_60575 (I1032497,I1032446,I1032480);
DFFARX1 I_60576 (I1032497,I2683,I1032299,I1032264,);
not I_60577 (I1032528,I1032480);
nand I_60578 (I1032545,I1032350,I1032528);
nand I_60579 (I1032276,I1032412,I1032528);
DFFARX1 I_60580 (I1032446,I2683,I1032299,I1032291,);
not I_60581 (I1032590,I233801);
nor I_60582 (I1032607,I1032590,I233774);
nor I_60583 (I1032624,I1032607,I1032429);
DFFARX1 I_60584 (I1032624,I2683,I1032299,I1032288,);
not I_60585 (I1032655,I1032607);
DFFARX1 I_60586 (I1032655,I2683,I1032299,I1032681,);
not I_60587 (I1032689,I1032681);
nor I_60588 (I1032285,I1032689,I1032607);
nor I_60589 (I1032720,I1032590,I233783);
and I_60590 (I1032737,I1032720,I233780);
or I_60591 (I1032754,I1032737,I233774);
DFFARX1 I_60592 (I1032754,I2683,I1032299,I1032780,);
not I_60593 (I1032788,I1032780);
nand I_60594 (I1032805,I1032788,I1032528);
not I_60595 (I1032279,I1032805);
nand I_60596 (I1032273,I1032805,I1032545);
nand I_60597 (I1032270,I1032788,I1032412);
not I_60598 (I1032894,I2690);
DFFARX1 I_60599 (I77514,I2683,I1032894,I1032920,);
DFFARX1 I_60600 (I77502,I2683,I1032894,I1032937,);
not I_60601 (I1032945,I1032937);
nor I_60602 (I1032862,I1032920,I1032945);
DFFARX1 I_60603 (I1032945,I2683,I1032894,I1032877,);
nor I_60604 (I1032990,I77493,I77517);
and I_60605 (I1033007,I1032990,I77496);
nor I_60606 (I1033024,I1033007,I77493);
not I_60607 (I1033041,I77493);
and I_60608 (I1033058,I1033041,I77499);
nand I_60609 (I1033075,I1033058,I77511);
nor I_60610 (I1033092,I1033041,I1033075);
DFFARX1 I_60611 (I1033092,I2683,I1032894,I1032859,);
not I_60612 (I1033123,I1033075);
nand I_60613 (I1033140,I1032945,I1033123);
nand I_60614 (I1032871,I1033007,I1033123);
DFFARX1 I_60615 (I1033041,I2683,I1032894,I1032886,);
not I_60616 (I1033185,I77493);
nor I_60617 (I1033202,I1033185,I77499);
nor I_60618 (I1033219,I1033202,I1033024);
DFFARX1 I_60619 (I1033219,I2683,I1032894,I1032883,);
not I_60620 (I1033250,I1033202);
DFFARX1 I_60621 (I1033250,I2683,I1032894,I1033276,);
not I_60622 (I1033284,I1033276);
nor I_60623 (I1032880,I1033284,I1033202);
nor I_60624 (I1033315,I1033185,I77496);
and I_60625 (I1033332,I1033315,I77505);
or I_60626 (I1033349,I1033332,I77508);
DFFARX1 I_60627 (I1033349,I2683,I1032894,I1033375,);
not I_60628 (I1033383,I1033375);
nand I_60629 (I1033400,I1033383,I1033123);
not I_60630 (I1032874,I1033400);
nand I_60631 (I1032868,I1033400,I1033140);
nand I_60632 (I1032865,I1033383,I1033007);
not I_60633 (I1033489,I2690);
DFFARX1 I_60634 (I679710,I2683,I1033489,I1033515,);
DFFARX1 I_60635 (I679707,I2683,I1033489,I1033532,);
not I_60636 (I1033540,I1033532);
nor I_60637 (I1033457,I1033515,I1033540);
DFFARX1 I_60638 (I1033540,I2683,I1033489,I1033472,);
nor I_60639 (I1033585,I679722,I679704);
and I_60640 (I1033602,I1033585,I679701);
nor I_60641 (I1033619,I1033602,I679722);
not I_60642 (I1033636,I679722);
and I_60643 (I1033653,I1033636,I679707);
nand I_60644 (I1033670,I1033653,I679719);
nor I_60645 (I1033687,I1033636,I1033670);
DFFARX1 I_60646 (I1033687,I2683,I1033489,I1033454,);
not I_60647 (I1033718,I1033670);
nand I_60648 (I1033735,I1033540,I1033718);
nand I_60649 (I1033466,I1033602,I1033718);
DFFARX1 I_60650 (I1033636,I2683,I1033489,I1033481,);
not I_60651 (I1033780,I679713);
nor I_60652 (I1033797,I1033780,I679707);
nor I_60653 (I1033814,I1033797,I1033619);
DFFARX1 I_60654 (I1033814,I2683,I1033489,I1033478,);
not I_60655 (I1033845,I1033797);
DFFARX1 I_60656 (I1033845,I2683,I1033489,I1033871,);
not I_60657 (I1033879,I1033871);
nor I_60658 (I1033475,I1033879,I1033797);
nor I_60659 (I1033910,I1033780,I679701);
and I_60660 (I1033927,I1033910,I679716);
or I_60661 (I1033944,I1033927,I679704);
DFFARX1 I_60662 (I1033944,I2683,I1033489,I1033970,);
not I_60663 (I1033978,I1033970);
nand I_60664 (I1033995,I1033978,I1033718);
not I_60665 (I1033469,I1033995);
nand I_60666 (I1033463,I1033995,I1033735);
nand I_60667 (I1033460,I1033978,I1033602);
not I_60668 (I1034084,I2690);
DFFARX1 I_60669 (I1004198,I2683,I1034084,I1034110,);
DFFARX1 I_60670 (I1004189,I2683,I1034084,I1034127,);
not I_60671 (I1034135,I1034127);
nor I_60672 (I1034052,I1034110,I1034135);
DFFARX1 I_60673 (I1034135,I2683,I1034084,I1034067,);
nor I_60674 (I1034180,I1004180,I1004195);
and I_60675 (I1034197,I1034180,I1004183);
nor I_60676 (I1034214,I1034197,I1004180);
not I_60677 (I1034231,I1004180);
and I_60678 (I1034248,I1034231,I1004186);
nand I_60679 (I1034265,I1034248,I1004204);
nor I_60680 (I1034282,I1034231,I1034265);
DFFARX1 I_60681 (I1034282,I2683,I1034084,I1034049,);
not I_60682 (I1034313,I1034265);
nand I_60683 (I1034330,I1034135,I1034313);
nand I_60684 (I1034061,I1034197,I1034313);
DFFARX1 I_60685 (I1034231,I2683,I1034084,I1034076,);
not I_60686 (I1034375,I1004180);
nor I_60687 (I1034392,I1034375,I1004186);
nor I_60688 (I1034409,I1034392,I1034214);
DFFARX1 I_60689 (I1034409,I2683,I1034084,I1034073,);
not I_60690 (I1034440,I1034392);
DFFARX1 I_60691 (I1034440,I2683,I1034084,I1034466,);
not I_60692 (I1034474,I1034466);
nor I_60693 (I1034070,I1034474,I1034392);
nor I_60694 (I1034505,I1034375,I1004183);
and I_60695 (I1034522,I1034505,I1004192);
or I_60696 (I1034539,I1034522,I1004201);
DFFARX1 I_60697 (I1034539,I2683,I1034084,I1034565,);
not I_60698 (I1034573,I1034565);
nand I_60699 (I1034590,I1034573,I1034313);
not I_60700 (I1034064,I1034590);
nand I_60701 (I1034058,I1034590,I1034330);
nand I_60702 (I1034055,I1034573,I1034197);
not I_60703 (I1034679,I2690);
DFFARX1 I_60704 (I38513,I2683,I1034679,I1034705,);
DFFARX1 I_60705 (I38495,I2683,I1034679,I1034722,);
not I_60706 (I1034730,I1034722);
nor I_60707 (I1034647,I1034705,I1034730);
DFFARX1 I_60708 (I1034730,I2683,I1034679,I1034662,);
nor I_60709 (I1034775,I38495,I38510);
and I_60710 (I1034792,I1034775,I38504);
nor I_60711 (I1034809,I1034792,I38495);
not I_60712 (I1034826,I38495);
and I_60713 (I1034843,I1034826,I38498);
nand I_60714 (I1034860,I1034843,I38501);
nor I_60715 (I1034877,I1034826,I1034860);
DFFARX1 I_60716 (I1034877,I2683,I1034679,I1034644,);
not I_60717 (I1034908,I1034860);
nand I_60718 (I1034925,I1034730,I1034908);
nand I_60719 (I1034656,I1034792,I1034908);
DFFARX1 I_60720 (I1034826,I2683,I1034679,I1034671,);
not I_60721 (I1034970,I38507);
nor I_60722 (I1034987,I1034970,I38498);
nor I_60723 (I1035004,I1034987,I1034809);
DFFARX1 I_60724 (I1035004,I2683,I1034679,I1034668,);
not I_60725 (I1035035,I1034987);
DFFARX1 I_60726 (I1035035,I2683,I1034679,I1035061,);
not I_60727 (I1035069,I1035061);
nor I_60728 (I1034665,I1035069,I1034987);
nor I_60729 (I1035100,I1034970,I38519);
and I_60730 (I1035117,I1035100,I38516);
or I_60731 (I1035134,I1035117,I38498);
DFFARX1 I_60732 (I1035134,I2683,I1034679,I1035160,);
not I_60733 (I1035168,I1035160);
nand I_60734 (I1035185,I1035168,I1034908);
not I_60735 (I1034659,I1035185);
nand I_60736 (I1034653,I1035185,I1034925);
nand I_60737 (I1034650,I1035168,I1034792);
not I_60738 (I1035274,I2690);
DFFARX1 I_60739 (I625956,I2683,I1035274,I1035300,);
DFFARX1 I_60740 (I625953,I2683,I1035274,I1035317,);
not I_60741 (I1035325,I1035317);
nor I_60742 (I1035242,I1035300,I1035325);
DFFARX1 I_60743 (I1035325,I2683,I1035274,I1035257,);
nor I_60744 (I1035370,I625968,I625950);
and I_60745 (I1035387,I1035370,I625947);
nor I_60746 (I1035404,I1035387,I625968);
not I_60747 (I1035421,I625968);
and I_60748 (I1035438,I1035421,I625953);
nand I_60749 (I1035455,I1035438,I625965);
nor I_60750 (I1035472,I1035421,I1035455);
DFFARX1 I_60751 (I1035472,I2683,I1035274,I1035239,);
not I_60752 (I1035503,I1035455);
nand I_60753 (I1035520,I1035325,I1035503);
nand I_60754 (I1035251,I1035387,I1035503);
DFFARX1 I_60755 (I1035421,I2683,I1035274,I1035266,);
not I_60756 (I1035565,I625959);
nor I_60757 (I1035582,I1035565,I625953);
nor I_60758 (I1035599,I1035582,I1035404);
DFFARX1 I_60759 (I1035599,I2683,I1035274,I1035263,);
not I_60760 (I1035630,I1035582);
DFFARX1 I_60761 (I1035630,I2683,I1035274,I1035656,);
not I_60762 (I1035664,I1035656);
nor I_60763 (I1035260,I1035664,I1035582);
nor I_60764 (I1035695,I1035565,I625947);
and I_60765 (I1035712,I1035695,I625962);
or I_60766 (I1035729,I1035712,I625950);
DFFARX1 I_60767 (I1035729,I2683,I1035274,I1035755,);
not I_60768 (I1035763,I1035755);
nand I_60769 (I1035780,I1035763,I1035503);
not I_60770 (I1035254,I1035780);
nand I_60771 (I1035248,I1035780,I1035520);
nand I_60772 (I1035245,I1035763,I1035387);
not I_60773 (I1035869,I2690);
DFFARX1 I_60774 (I25338,I2683,I1035869,I1035895,);
DFFARX1 I_60775 (I25320,I2683,I1035869,I1035912,);
not I_60776 (I1035920,I1035912);
nor I_60777 (I1035837,I1035895,I1035920);
DFFARX1 I_60778 (I1035920,I2683,I1035869,I1035852,);
nor I_60779 (I1035965,I25320,I25335);
and I_60780 (I1035982,I1035965,I25329);
nor I_60781 (I1035999,I1035982,I25320);
not I_60782 (I1036016,I25320);
and I_60783 (I1036033,I1036016,I25323);
nand I_60784 (I1036050,I1036033,I25326);
nor I_60785 (I1036067,I1036016,I1036050);
DFFARX1 I_60786 (I1036067,I2683,I1035869,I1035834,);
not I_60787 (I1036098,I1036050);
nand I_60788 (I1036115,I1035920,I1036098);
nand I_60789 (I1035846,I1035982,I1036098);
DFFARX1 I_60790 (I1036016,I2683,I1035869,I1035861,);
not I_60791 (I1036160,I25332);
nor I_60792 (I1036177,I1036160,I25323);
nor I_60793 (I1036194,I1036177,I1035999);
DFFARX1 I_60794 (I1036194,I2683,I1035869,I1035858,);
not I_60795 (I1036225,I1036177);
DFFARX1 I_60796 (I1036225,I2683,I1035869,I1036251,);
not I_60797 (I1036259,I1036251);
nor I_60798 (I1035855,I1036259,I1036177);
nor I_60799 (I1036290,I1036160,I25344);
and I_60800 (I1036307,I1036290,I25341);
or I_60801 (I1036324,I1036307,I25323);
DFFARX1 I_60802 (I1036324,I2683,I1035869,I1036350,);
not I_60803 (I1036358,I1036350);
nand I_60804 (I1036375,I1036358,I1036098);
not I_60805 (I1035849,I1036375);
nand I_60806 (I1035843,I1036375,I1036115);
nand I_60807 (I1035840,I1036358,I1035982);
not I_60808 (I1036464,I2690);
DFFARX1 I_60809 (I461901,I2683,I1036464,I1036490,);
DFFARX1 I_60810 (I461895,I2683,I1036464,I1036507,);
not I_60811 (I1036515,I1036507);
nor I_60812 (I1036432,I1036490,I1036515);
DFFARX1 I_60813 (I1036515,I2683,I1036464,I1036447,);
nor I_60814 (I1036560,I461892,I461883);
and I_60815 (I1036577,I1036560,I461880);
nor I_60816 (I1036594,I1036577,I461892);
not I_60817 (I1036611,I461892);
and I_60818 (I1036628,I1036611,I461886);
nand I_60819 (I1036645,I1036628,I461898);
nor I_60820 (I1036662,I1036611,I1036645);
DFFARX1 I_60821 (I1036662,I2683,I1036464,I1036429,);
not I_60822 (I1036693,I1036645);
nand I_60823 (I1036710,I1036515,I1036693);
nand I_60824 (I1036441,I1036577,I1036693);
DFFARX1 I_60825 (I1036611,I2683,I1036464,I1036456,);
not I_60826 (I1036755,I461904);
nor I_60827 (I1036772,I1036755,I461886);
nor I_60828 (I1036789,I1036772,I1036594);
DFFARX1 I_60829 (I1036789,I2683,I1036464,I1036453,);
not I_60830 (I1036820,I1036772);
DFFARX1 I_60831 (I1036820,I2683,I1036464,I1036846,);
not I_60832 (I1036854,I1036846);
nor I_60833 (I1036450,I1036854,I1036772);
nor I_60834 (I1036885,I1036755,I461883);
and I_60835 (I1036902,I1036885,I461889);
or I_60836 (I1036919,I1036902,I461880);
DFFARX1 I_60837 (I1036919,I2683,I1036464,I1036945,);
not I_60838 (I1036953,I1036945);
nand I_60839 (I1036970,I1036953,I1036693);
not I_60840 (I1036444,I1036970);
nand I_60841 (I1036438,I1036970,I1036710);
nand I_60842 (I1036435,I1036953,I1036577);
not I_60843 (I1037059,I2690);
DFFARX1 I_60844 (I140835,I2683,I1037059,I1037085,);
DFFARX1 I_60845 (I140838,I2683,I1037059,I1037102,);
not I_60846 (I1037110,I1037102);
nor I_60847 (I1037027,I1037085,I1037110);
DFFARX1 I_60848 (I1037110,I2683,I1037059,I1037042,);
nor I_60849 (I1037155,I140844,I140838);
and I_60850 (I1037172,I1037155,I140841);
nor I_60851 (I1037189,I1037172,I140844);
not I_60852 (I1037206,I140844);
and I_60853 (I1037223,I1037206,I140835);
nand I_60854 (I1037240,I1037223,I140853);
nor I_60855 (I1037257,I1037206,I1037240);
DFFARX1 I_60856 (I1037257,I2683,I1037059,I1037024,);
not I_60857 (I1037288,I1037240);
nand I_60858 (I1037305,I1037110,I1037288);
nand I_60859 (I1037036,I1037172,I1037288);
DFFARX1 I_60860 (I1037206,I2683,I1037059,I1037051,);
not I_60861 (I1037350,I140847);
nor I_60862 (I1037367,I1037350,I140835);
nor I_60863 (I1037384,I1037367,I1037189);
DFFARX1 I_60864 (I1037384,I2683,I1037059,I1037048,);
not I_60865 (I1037415,I1037367);
DFFARX1 I_60866 (I1037415,I2683,I1037059,I1037441,);
not I_60867 (I1037449,I1037441);
nor I_60868 (I1037045,I1037449,I1037367);
nor I_60869 (I1037480,I1037350,I140850);
and I_60870 (I1037497,I1037480,I140856);
or I_60871 (I1037514,I1037497,I140859);
DFFARX1 I_60872 (I1037514,I2683,I1037059,I1037540,);
not I_60873 (I1037548,I1037540);
nand I_60874 (I1037565,I1037548,I1037288);
not I_60875 (I1037039,I1037565);
nand I_60876 (I1037033,I1037565,I1037305);
nand I_60877 (I1037030,I1037548,I1037172);
not I_60878 (I1037654,I2690);
DFFARX1 I_60879 (I916055,I2683,I1037654,I1037680,);
DFFARX1 I_60880 (I916067,I2683,I1037654,I1037697,);
not I_60881 (I1037705,I1037697);
nor I_60882 (I1037622,I1037680,I1037705);
DFFARX1 I_60883 (I1037705,I2683,I1037654,I1037637,);
nor I_60884 (I1037750,I916064,I916058);
and I_60885 (I1037767,I1037750,I916052);
nor I_60886 (I1037784,I1037767,I916064);
not I_60887 (I1037801,I916064);
and I_60888 (I1037818,I1037801,I916061);
nand I_60889 (I1037835,I1037818,I916052);
nor I_60890 (I1037852,I1037801,I1037835);
DFFARX1 I_60891 (I1037852,I2683,I1037654,I1037619,);
not I_60892 (I1037883,I1037835);
nand I_60893 (I1037900,I1037705,I1037883);
nand I_60894 (I1037631,I1037767,I1037883);
DFFARX1 I_60895 (I1037801,I2683,I1037654,I1037646,);
not I_60896 (I1037945,I916076);
nor I_60897 (I1037962,I1037945,I916061);
nor I_60898 (I1037979,I1037962,I1037784);
DFFARX1 I_60899 (I1037979,I2683,I1037654,I1037643,);
not I_60900 (I1038010,I1037962);
DFFARX1 I_60901 (I1038010,I2683,I1037654,I1038036,);
not I_60902 (I1038044,I1038036);
nor I_60903 (I1037640,I1038044,I1037962);
nor I_60904 (I1038075,I1037945,I916070);
and I_60905 (I1038092,I1038075,I916073);
or I_60906 (I1038109,I1038092,I916055);
DFFARX1 I_60907 (I1038109,I2683,I1037654,I1038135,);
not I_60908 (I1038143,I1038135);
nand I_60909 (I1038160,I1038143,I1037883);
not I_60910 (I1037634,I1038160);
nand I_60911 (I1037628,I1038160,I1037900);
nand I_60912 (I1037625,I1038143,I1037767);
not I_60913 (I1038249,I2690);
DFFARX1 I_60914 (I620159,I2683,I1038249,I1038275,);
DFFARX1 I_60915 (I620156,I2683,I1038249,I1038292,);
not I_60916 (I1038300,I1038292);
nor I_60917 (I1038217,I1038275,I1038300);
DFFARX1 I_60918 (I1038300,I2683,I1038249,I1038232,);
nor I_60919 (I1038345,I620171,I620153);
and I_60920 (I1038362,I1038345,I620150);
nor I_60921 (I1038379,I1038362,I620171);
not I_60922 (I1038396,I620171);
and I_60923 (I1038413,I1038396,I620156);
nand I_60924 (I1038430,I1038413,I620168);
nor I_60925 (I1038447,I1038396,I1038430);
DFFARX1 I_60926 (I1038447,I2683,I1038249,I1038214,);
not I_60927 (I1038478,I1038430);
nand I_60928 (I1038495,I1038300,I1038478);
nand I_60929 (I1038226,I1038362,I1038478);
DFFARX1 I_60930 (I1038396,I2683,I1038249,I1038241,);
not I_60931 (I1038540,I620162);
nor I_60932 (I1038557,I1038540,I620156);
nor I_60933 (I1038574,I1038557,I1038379);
DFFARX1 I_60934 (I1038574,I2683,I1038249,I1038238,);
not I_60935 (I1038605,I1038557);
DFFARX1 I_60936 (I1038605,I2683,I1038249,I1038631,);
not I_60937 (I1038639,I1038631);
nor I_60938 (I1038235,I1038639,I1038557);
nor I_60939 (I1038670,I1038540,I620150);
and I_60940 (I1038687,I1038670,I620165);
or I_60941 (I1038704,I1038687,I620153);
DFFARX1 I_60942 (I1038704,I2683,I1038249,I1038730,);
not I_60943 (I1038738,I1038730);
nand I_60944 (I1038755,I1038738,I1038478);
not I_60945 (I1038229,I1038755);
nand I_60946 (I1038223,I1038755,I1038495);
nand I_60947 (I1038220,I1038738,I1038362);
not I_60948 (I1038844,I2690);
DFFARX1 I_60949 (I665481,I2683,I1038844,I1038870,);
DFFARX1 I_60950 (I665478,I2683,I1038844,I1038887,);
not I_60951 (I1038895,I1038887);
nor I_60952 (I1038812,I1038870,I1038895);
DFFARX1 I_60953 (I1038895,I2683,I1038844,I1038827,);
nor I_60954 (I1038940,I665493,I665475);
and I_60955 (I1038957,I1038940,I665472);
nor I_60956 (I1038974,I1038957,I665493);
not I_60957 (I1038991,I665493);
and I_60958 (I1039008,I1038991,I665478);
nand I_60959 (I1039025,I1039008,I665490);
nor I_60960 (I1039042,I1038991,I1039025);
DFFARX1 I_60961 (I1039042,I2683,I1038844,I1038809,);
not I_60962 (I1039073,I1039025);
nand I_60963 (I1039090,I1038895,I1039073);
nand I_60964 (I1038821,I1038957,I1039073);
DFFARX1 I_60965 (I1038991,I2683,I1038844,I1038836,);
not I_60966 (I1039135,I665484);
nor I_60967 (I1039152,I1039135,I665478);
nor I_60968 (I1039169,I1039152,I1038974);
DFFARX1 I_60969 (I1039169,I2683,I1038844,I1038833,);
not I_60970 (I1039200,I1039152);
DFFARX1 I_60971 (I1039200,I2683,I1038844,I1039226,);
not I_60972 (I1039234,I1039226);
nor I_60973 (I1038830,I1039234,I1039152);
nor I_60974 (I1039265,I1039135,I665472);
and I_60975 (I1039282,I1039265,I665487);
or I_60976 (I1039299,I1039282,I665475);
DFFARX1 I_60977 (I1039299,I2683,I1038844,I1039325,);
not I_60978 (I1039333,I1039325);
nand I_60979 (I1039350,I1039333,I1039073);
not I_60980 (I1038824,I1039350);
nand I_60981 (I1038818,I1039350,I1039090);
nand I_60982 (I1038815,I1039333,I1038957);
not I_60983 (I1039439,I2690);
DFFARX1 I_60984 (I505251,I2683,I1039439,I1039465,);
DFFARX1 I_60985 (I505233,I2683,I1039439,I1039482,);
not I_60986 (I1039490,I1039482);
nor I_60987 (I1039407,I1039465,I1039490);
DFFARX1 I_60988 (I1039490,I2683,I1039439,I1039422,);
nor I_60989 (I1039535,I505239,I505242);
and I_60990 (I1039552,I1039535,I505230);
nor I_60991 (I1039569,I1039552,I505239);
not I_60992 (I1039586,I505239);
and I_60993 (I1039603,I1039586,I505248);
nand I_60994 (I1039620,I1039603,I505236);
nor I_60995 (I1039637,I1039586,I1039620);
DFFARX1 I_60996 (I1039637,I2683,I1039439,I1039404,);
not I_60997 (I1039668,I1039620);
nand I_60998 (I1039685,I1039490,I1039668);
nand I_60999 (I1039416,I1039552,I1039668);
DFFARX1 I_61000 (I1039586,I2683,I1039439,I1039431,);
not I_61001 (I1039730,I505233);
nor I_61002 (I1039747,I1039730,I505248);
nor I_61003 (I1039764,I1039747,I1039569);
DFFARX1 I_61004 (I1039764,I2683,I1039439,I1039428,);
not I_61005 (I1039795,I1039747);
DFFARX1 I_61006 (I1039795,I2683,I1039439,I1039821,);
not I_61007 (I1039829,I1039821);
nor I_61008 (I1039425,I1039829,I1039747);
nor I_61009 (I1039860,I1039730,I505245);
and I_61010 (I1039877,I1039860,I505254);
or I_61011 (I1039894,I1039877,I505230);
DFFARX1 I_61012 (I1039894,I2683,I1039439,I1039920,);
not I_61013 (I1039928,I1039920);
nand I_61014 (I1039945,I1039928,I1039668);
not I_61015 (I1039419,I1039945);
nand I_61016 (I1039413,I1039945,I1039685);
nand I_61017 (I1039410,I1039928,I1039552);
not I_61018 (I1040034,I2690);
DFFARX1 I_61019 (I1016914,I2683,I1040034,I1040060,);
DFFARX1 I_61020 (I1016905,I2683,I1040034,I1040077,);
not I_61021 (I1040085,I1040077);
nor I_61022 (I1040002,I1040060,I1040085);
DFFARX1 I_61023 (I1040085,I2683,I1040034,I1040017,);
nor I_61024 (I1040130,I1016896,I1016911);
and I_61025 (I1040147,I1040130,I1016899);
nor I_61026 (I1040164,I1040147,I1016896);
not I_61027 (I1040181,I1016896);
and I_61028 (I1040198,I1040181,I1016902);
nand I_61029 (I1040215,I1040198,I1016920);
nor I_61030 (I1040232,I1040181,I1040215);
DFFARX1 I_61031 (I1040232,I2683,I1040034,I1039999,);
not I_61032 (I1040263,I1040215);
nand I_61033 (I1040280,I1040085,I1040263);
nand I_61034 (I1040011,I1040147,I1040263);
DFFARX1 I_61035 (I1040181,I2683,I1040034,I1040026,);
not I_61036 (I1040325,I1016896);
nor I_61037 (I1040342,I1040325,I1016902);
nor I_61038 (I1040359,I1040342,I1040164);
DFFARX1 I_61039 (I1040359,I2683,I1040034,I1040023,);
not I_61040 (I1040390,I1040342);
DFFARX1 I_61041 (I1040390,I2683,I1040034,I1040416,);
not I_61042 (I1040424,I1040416);
nor I_61043 (I1040020,I1040424,I1040342);
nor I_61044 (I1040455,I1040325,I1016899);
and I_61045 (I1040472,I1040455,I1016908);
or I_61046 (I1040489,I1040472,I1016917);
DFFARX1 I_61047 (I1040489,I2683,I1040034,I1040515,);
not I_61048 (I1040523,I1040515);
nand I_61049 (I1040540,I1040523,I1040263);
not I_61050 (I1040014,I1040540);
nand I_61051 (I1040008,I1040540,I1040280);
nand I_61052 (I1040005,I1040523,I1040147);
not I_61053 (I1040629,I2690);
DFFARX1 I_61054 (I627010,I2683,I1040629,I1040655,);
DFFARX1 I_61055 (I627007,I2683,I1040629,I1040672,);
not I_61056 (I1040680,I1040672);
nor I_61057 (I1040597,I1040655,I1040680);
DFFARX1 I_61058 (I1040680,I2683,I1040629,I1040612,);
nor I_61059 (I1040725,I627022,I627004);
and I_61060 (I1040742,I1040725,I627001);
nor I_61061 (I1040759,I1040742,I627022);
not I_61062 (I1040776,I627022);
and I_61063 (I1040793,I1040776,I627007);
nand I_61064 (I1040810,I1040793,I627019);
nor I_61065 (I1040827,I1040776,I1040810);
DFFARX1 I_61066 (I1040827,I2683,I1040629,I1040594,);
not I_61067 (I1040858,I1040810);
nand I_61068 (I1040875,I1040680,I1040858);
nand I_61069 (I1040606,I1040742,I1040858);
DFFARX1 I_61070 (I1040776,I2683,I1040629,I1040621,);
not I_61071 (I1040920,I627013);
nor I_61072 (I1040937,I1040920,I627007);
nor I_61073 (I1040954,I1040937,I1040759);
DFFARX1 I_61074 (I1040954,I2683,I1040629,I1040618,);
not I_61075 (I1040985,I1040937);
DFFARX1 I_61076 (I1040985,I2683,I1040629,I1041011,);
not I_61077 (I1041019,I1041011);
nor I_61078 (I1040615,I1041019,I1040937);
nor I_61079 (I1041050,I1040920,I627001);
and I_61080 (I1041067,I1041050,I627016);
or I_61081 (I1041084,I1041067,I627004);
DFFARX1 I_61082 (I1041084,I2683,I1040629,I1041110,);
not I_61083 (I1041118,I1041110);
nand I_61084 (I1041135,I1041118,I1040858);
not I_61085 (I1040609,I1041135);
nand I_61086 (I1040603,I1041135,I1040875);
nand I_61087 (I1040600,I1041118,I1040742);
not I_61088 (I1041224,I2690);
DFFARX1 I_61089 (I794287,I2683,I1041224,I1041250,);
DFFARX1 I_61090 (I794305,I2683,I1041224,I1041267,);
not I_61091 (I1041275,I1041267);
nor I_61092 (I1041192,I1041250,I1041275);
DFFARX1 I_61093 (I1041275,I2683,I1041224,I1041207,);
nor I_61094 (I1041320,I794284,I794296);
and I_61095 (I1041337,I1041320,I794281);
nor I_61096 (I1041354,I1041337,I794284);
not I_61097 (I1041371,I794284);
and I_61098 (I1041388,I1041371,I794290);
nand I_61099 (I1041405,I1041388,I794302);
nor I_61100 (I1041422,I1041371,I1041405);
DFFARX1 I_61101 (I1041422,I2683,I1041224,I1041189,);
not I_61102 (I1041453,I1041405);
nand I_61103 (I1041470,I1041275,I1041453);
nand I_61104 (I1041201,I1041337,I1041453);
DFFARX1 I_61105 (I1041371,I2683,I1041224,I1041216,);
not I_61106 (I1041515,I794293);
nor I_61107 (I1041532,I1041515,I794290);
nor I_61108 (I1041549,I1041532,I1041354);
DFFARX1 I_61109 (I1041549,I2683,I1041224,I1041213,);
not I_61110 (I1041580,I1041532);
DFFARX1 I_61111 (I1041580,I2683,I1041224,I1041606,);
not I_61112 (I1041614,I1041606);
nor I_61113 (I1041210,I1041614,I1041532);
nor I_61114 (I1041645,I1041515,I794281);
and I_61115 (I1041662,I1041645,I794308);
or I_61116 (I1041679,I1041662,I794299);
DFFARX1 I_61117 (I1041679,I2683,I1041224,I1041705,);
not I_61118 (I1041713,I1041705);
nand I_61119 (I1041730,I1041713,I1041453);
not I_61120 (I1041204,I1041730);
nand I_61121 (I1041198,I1041730,I1041470);
nand I_61122 (I1041195,I1041713,I1041337);
not I_61123 (I1041819,I2690);
DFFARX1 I_61124 (I99121,I2683,I1041819,I1041845,);
DFFARX1 I_61125 (I99109,I2683,I1041819,I1041862,);
not I_61126 (I1041870,I1041862);
nor I_61127 (I1041787,I1041845,I1041870);
DFFARX1 I_61128 (I1041870,I2683,I1041819,I1041802,);
nor I_61129 (I1041915,I99100,I99124);
and I_61130 (I1041932,I1041915,I99103);
nor I_61131 (I1041949,I1041932,I99100);
not I_61132 (I1041966,I99100);
and I_61133 (I1041983,I1041966,I99106);
nand I_61134 (I1042000,I1041983,I99118);
nor I_61135 (I1042017,I1041966,I1042000);
DFFARX1 I_61136 (I1042017,I2683,I1041819,I1041784,);
not I_61137 (I1042048,I1042000);
nand I_61138 (I1042065,I1041870,I1042048);
nand I_61139 (I1041796,I1041932,I1042048);
DFFARX1 I_61140 (I1041966,I2683,I1041819,I1041811,);
not I_61141 (I1042110,I99100);
nor I_61142 (I1042127,I1042110,I99106);
nor I_61143 (I1042144,I1042127,I1041949);
DFFARX1 I_61144 (I1042144,I2683,I1041819,I1041808,);
not I_61145 (I1042175,I1042127);
DFFARX1 I_61146 (I1042175,I2683,I1041819,I1042201,);
not I_61147 (I1042209,I1042201);
nor I_61148 (I1041805,I1042209,I1042127);
nor I_61149 (I1042240,I1042110,I99103);
and I_61150 (I1042257,I1042240,I99112);
or I_61151 (I1042274,I1042257,I99115);
DFFARX1 I_61152 (I1042274,I2683,I1041819,I1042300,);
not I_61153 (I1042308,I1042300);
nand I_61154 (I1042325,I1042308,I1042048);
not I_61155 (I1041799,I1042325);
nand I_61156 (I1041793,I1042325,I1042065);
nand I_61157 (I1041790,I1042308,I1041932);
not I_61158 (I1042414,I2690);
DFFARX1 I_61159 (I62231,I2683,I1042414,I1042440,);
DFFARX1 I_61160 (I62219,I2683,I1042414,I1042457,);
not I_61161 (I1042465,I1042457);
nor I_61162 (I1042382,I1042440,I1042465);
DFFARX1 I_61163 (I1042465,I2683,I1042414,I1042397,);
nor I_61164 (I1042510,I62210,I62234);
and I_61165 (I1042527,I1042510,I62213);
nor I_61166 (I1042544,I1042527,I62210);
not I_61167 (I1042561,I62210);
and I_61168 (I1042578,I1042561,I62216);
nand I_61169 (I1042595,I1042578,I62228);
nor I_61170 (I1042612,I1042561,I1042595);
DFFARX1 I_61171 (I1042612,I2683,I1042414,I1042379,);
not I_61172 (I1042643,I1042595);
nand I_61173 (I1042660,I1042465,I1042643);
nand I_61174 (I1042391,I1042527,I1042643);
DFFARX1 I_61175 (I1042561,I2683,I1042414,I1042406,);
not I_61176 (I1042705,I62210);
nor I_61177 (I1042722,I1042705,I62216);
nor I_61178 (I1042739,I1042722,I1042544);
DFFARX1 I_61179 (I1042739,I2683,I1042414,I1042403,);
not I_61180 (I1042770,I1042722);
DFFARX1 I_61181 (I1042770,I2683,I1042414,I1042796,);
not I_61182 (I1042804,I1042796);
nor I_61183 (I1042400,I1042804,I1042722);
nor I_61184 (I1042835,I1042705,I62213);
and I_61185 (I1042852,I1042835,I62222);
or I_61186 (I1042869,I1042852,I62225);
DFFARX1 I_61187 (I1042869,I2683,I1042414,I1042895,);
not I_61188 (I1042903,I1042895);
nand I_61189 (I1042920,I1042903,I1042643);
not I_61190 (I1042394,I1042920);
nand I_61191 (I1042388,I1042920,I1042660);
nand I_61192 (I1042385,I1042903,I1042527);
not I_61193 (I1043009,I2690);
DFFARX1 I_61194 (I2636,I2683,I1043009,I1043035,);
DFFARX1 I_61195 (I1556,I2683,I1043009,I1043052,);
not I_61196 (I1043060,I1043052);
nor I_61197 (I1042977,I1043035,I1043060);
DFFARX1 I_61198 (I1043060,I2683,I1043009,I1042992,);
nor I_61199 (I1043105,I2180,I2092);
and I_61200 (I1043122,I1043105,I1868);
nor I_61201 (I1043139,I1043122,I2180);
not I_61202 (I1043156,I2180);
and I_61203 (I1043173,I1043156,I2324);
nand I_61204 (I1043190,I1043173,I1972);
nor I_61205 (I1043207,I1043156,I1043190);
DFFARX1 I_61206 (I1043207,I2683,I1043009,I1042974,);
not I_61207 (I1043238,I1043190);
nand I_61208 (I1043255,I1043060,I1043238);
nand I_61209 (I1042986,I1043122,I1043238);
DFFARX1 I_61210 (I1043156,I2683,I1043009,I1043001,);
not I_61211 (I1043300,I1516);
nor I_61212 (I1043317,I1043300,I2324);
nor I_61213 (I1043334,I1043317,I1043139);
DFFARX1 I_61214 (I1043334,I2683,I1043009,I1042998,);
not I_61215 (I1043365,I1043317);
DFFARX1 I_61216 (I1043365,I2683,I1043009,I1043391,);
not I_61217 (I1043399,I1043391);
nor I_61218 (I1042995,I1043399,I1043317);
nor I_61219 (I1043430,I1043300,I2220);
and I_61220 (I1043447,I1043430,I1820);
or I_61221 (I1043464,I1043447,I2300);
DFFARX1 I_61222 (I1043464,I2683,I1043009,I1043490,);
not I_61223 (I1043498,I1043490);
nand I_61224 (I1043515,I1043498,I1043238);
not I_61225 (I1042989,I1043515);
nand I_61226 (I1042983,I1043515,I1043255);
nand I_61227 (I1042980,I1043498,I1043122);
not I_61228 (I1043604,I2690);
DFFARX1 I_61229 (I966270,I2683,I1043604,I1043630,);
DFFARX1 I_61230 (I966273,I2683,I1043604,I1043647,);
not I_61231 (I1043655,I1043647);
nor I_61232 (I1043572,I1043630,I1043655);
DFFARX1 I_61233 (I1043655,I2683,I1043604,I1043587,);
nor I_61234 (I1043700,I966273,I966288);
and I_61235 (I1043717,I1043700,I966282);
nor I_61236 (I1043734,I1043717,I966273);
not I_61237 (I1043751,I966273);
and I_61238 (I1043768,I1043751,I966291);
nand I_61239 (I1043785,I1043768,I966279);
nor I_61240 (I1043802,I1043751,I1043785);
DFFARX1 I_61241 (I1043802,I2683,I1043604,I1043569,);
not I_61242 (I1043833,I1043785);
nand I_61243 (I1043850,I1043655,I1043833);
nand I_61244 (I1043581,I1043717,I1043833);
DFFARX1 I_61245 (I1043751,I2683,I1043604,I1043596,);
not I_61246 (I1043895,I966285);
nor I_61247 (I1043912,I1043895,I966291);
nor I_61248 (I1043929,I1043912,I1043734);
DFFARX1 I_61249 (I1043929,I2683,I1043604,I1043593,);
not I_61250 (I1043960,I1043912);
DFFARX1 I_61251 (I1043960,I2683,I1043604,I1043986,);
not I_61252 (I1043994,I1043986);
nor I_61253 (I1043590,I1043994,I1043912);
nor I_61254 (I1044025,I1043895,I966270);
and I_61255 (I1044042,I1044025,I966294);
or I_61256 (I1044059,I1044042,I966276);
DFFARX1 I_61257 (I1044059,I2683,I1043604,I1044085,);
not I_61258 (I1044093,I1044085);
nand I_61259 (I1044110,I1044093,I1043833);
not I_61260 (I1043584,I1044110);
nand I_61261 (I1043578,I1044110,I1043850);
nand I_61262 (I1043575,I1044093,I1043717);
not I_61263 (I1044199,I2690);
DFFARX1 I_61264 (I997262,I2683,I1044199,I1044225,);
DFFARX1 I_61265 (I997253,I2683,I1044199,I1044242,);
not I_61266 (I1044250,I1044242);
nor I_61267 (I1044167,I1044225,I1044250);
DFFARX1 I_61268 (I1044250,I2683,I1044199,I1044182,);
nor I_61269 (I1044295,I997244,I997259);
and I_61270 (I1044312,I1044295,I997247);
nor I_61271 (I1044329,I1044312,I997244);
not I_61272 (I1044346,I997244);
and I_61273 (I1044363,I1044346,I997250);
nand I_61274 (I1044380,I1044363,I997268);
nor I_61275 (I1044397,I1044346,I1044380);
DFFARX1 I_61276 (I1044397,I2683,I1044199,I1044164,);
not I_61277 (I1044428,I1044380);
nand I_61278 (I1044445,I1044250,I1044428);
nand I_61279 (I1044176,I1044312,I1044428);
DFFARX1 I_61280 (I1044346,I2683,I1044199,I1044191,);
not I_61281 (I1044490,I997244);
nor I_61282 (I1044507,I1044490,I997250);
nor I_61283 (I1044524,I1044507,I1044329);
DFFARX1 I_61284 (I1044524,I2683,I1044199,I1044188,);
not I_61285 (I1044555,I1044507);
DFFARX1 I_61286 (I1044555,I2683,I1044199,I1044581,);
not I_61287 (I1044589,I1044581);
nor I_61288 (I1044185,I1044589,I1044507);
nor I_61289 (I1044620,I1044490,I997247);
and I_61290 (I1044637,I1044620,I997256);
or I_61291 (I1044654,I1044637,I997265);
DFFARX1 I_61292 (I1044654,I2683,I1044199,I1044680,);
not I_61293 (I1044688,I1044680);
nand I_61294 (I1044705,I1044688,I1044428);
not I_61295 (I1044179,I1044705);
nand I_61296 (I1044173,I1044705,I1044445);
nand I_61297 (I1044170,I1044688,I1044312);
not I_61298 (I1044794,I2690);
DFFARX1 I_61299 (I624375,I2683,I1044794,I1044820,);
DFFARX1 I_61300 (I624372,I2683,I1044794,I1044837,);
not I_61301 (I1044845,I1044837);
nor I_61302 (I1044762,I1044820,I1044845);
DFFARX1 I_61303 (I1044845,I2683,I1044794,I1044777,);
nor I_61304 (I1044890,I624387,I624369);
and I_61305 (I1044907,I1044890,I624366);
nor I_61306 (I1044924,I1044907,I624387);
not I_61307 (I1044941,I624387);
and I_61308 (I1044958,I1044941,I624372);
nand I_61309 (I1044975,I1044958,I624384);
nor I_61310 (I1044992,I1044941,I1044975);
DFFARX1 I_61311 (I1044992,I2683,I1044794,I1044759,);
not I_61312 (I1045023,I1044975);
nand I_61313 (I1045040,I1044845,I1045023);
nand I_61314 (I1044771,I1044907,I1045023);
DFFARX1 I_61315 (I1044941,I2683,I1044794,I1044786,);
not I_61316 (I1045085,I624378);
nor I_61317 (I1045102,I1045085,I624372);
nor I_61318 (I1045119,I1045102,I1044924);
DFFARX1 I_61319 (I1045119,I2683,I1044794,I1044783,);
not I_61320 (I1045150,I1045102);
DFFARX1 I_61321 (I1045150,I2683,I1044794,I1045176,);
not I_61322 (I1045184,I1045176);
nor I_61323 (I1044780,I1045184,I1045102);
nor I_61324 (I1045215,I1045085,I624366);
and I_61325 (I1045232,I1045215,I624381);
or I_61326 (I1045249,I1045232,I624369);
DFFARX1 I_61327 (I1045249,I2683,I1044794,I1045275,);
not I_61328 (I1045283,I1045275);
nand I_61329 (I1045300,I1045283,I1045023);
not I_61330 (I1044774,I1045300);
nand I_61331 (I1044768,I1045300,I1045040);
nand I_61332 (I1044765,I1045283,I1044907);
not I_61333 (I1045389,I2690);
DFFARX1 I_61334 (I980958,I2683,I1045389,I1045415,);
DFFARX1 I_61335 (I980961,I2683,I1045389,I1045432,);
not I_61336 (I1045440,I1045432);
nor I_61337 (I1045357,I1045415,I1045440);
DFFARX1 I_61338 (I1045440,I2683,I1045389,I1045372,);
nor I_61339 (I1045485,I980961,I980976);
and I_61340 (I1045502,I1045485,I980970);
nor I_61341 (I1045519,I1045502,I980961);
not I_61342 (I1045536,I980961);
and I_61343 (I1045553,I1045536,I980979);
nand I_61344 (I1045570,I1045553,I980967);
nor I_61345 (I1045587,I1045536,I1045570);
DFFARX1 I_61346 (I1045587,I2683,I1045389,I1045354,);
not I_61347 (I1045618,I1045570);
nand I_61348 (I1045635,I1045440,I1045618);
nand I_61349 (I1045366,I1045502,I1045618);
DFFARX1 I_61350 (I1045536,I2683,I1045389,I1045381,);
not I_61351 (I1045680,I980973);
nor I_61352 (I1045697,I1045680,I980979);
nor I_61353 (I1045714,I1045697,I1045519);
DFFARX1 I_61354 (I1045714,I2683,I1045389,I1045378,);
not I_61355 (I1045745,I1045697);
DFFARX1 I_61356 (I1045745,I2683,I1045389,I1045771,);
not I_61357 (I1045779,I1045771);
nor I_61358 (I1045375,I1045779,I1045697);
nor I_61359 (I1045810,I1045680,I980958);
and I_61360 (I1045827,I1045810,I980982);
or I_61361 (I1045844,I1045827,I980964);
DFFARX1 I_61362 (I1045844,I2683,I1045389,I1045870,);
not I_61363 (I1045878,I1045870);
nand I_61364 (I1045895,I1045878,I1045618);
not I_61365 (I1045369,I1045895);
nand I_61366 (I1045363,I1045895,I1045635);
nand I_61367 (I1045360,I1045878,I1045502);
not I_61368 (I1045984,I2690);
DFFARX1 I_61369 (I776199,I2683,I1045984,I1046010,);
DFFARX1 I_61370 (I776217,I2683,I1045984,I1046027,);
not I_61371 (I1046035,I1046027);
nor I_61372 (I1045952,I1046010,I1046035);
DFFARX1 I_61373 (I1046035,I2683,I1045984,I1045967,);
nor I_61374 (I1046080,I776196,I776208);
and I_61375 (I1046097,I1046080,I776193);
nor I_61376 (I1046114,I1046097,I776196);
not I_61377 (I1046131,I776196);
and I_61378 (I1046148,I1046131,I776202);
nand I_61379 (I1046165,I1046148,I776214);
nor I_61380 (I1046182,I1046131,I1046165);
DFFARX1 I_61381 (I1046182,I2683,I1045984,I1045949,);
not I_61382 (I1046213,I1046165);
nand I_61383 (I1046230,I1046035,I1046213);
nand I_61384 (I1045961,I1046097,I1046213);
DFFARX1 I_61385 (I1046131,I2683,I1045984,I1045976,);
not I_61386 (I1046275,I776205);
nor I_61387 (I1046292,I1046275,I776202);
nor I_61388 (I1046309,I1046292,I1046114);
DFFARX1 I_61389 (I1046309,I2683,I1045984,I1045973,);
not I_61390 (I1046340,I1046292);
DFFARX1 I_61391 (I1046340,I2683,I1045984,I1046366,);
not I_61392 (I1046374,I1046366);
nor I_61393 (I1045970,I1046374,I1046292);
nor I_61394 (I1046405,I1046275,I776193);
and I_61395 (I1046422,I1046405,I776220);
or I_61396 (I1046439,I1046422,I776211);
DFFARX1 I_61397 (I1046439,I2683,I1045984,I1046465,);
not I_61398 (I1046473,I1046465);
nand I_61399 (I1046490,I1046473,I1046213);
not I_61400 (I1045964,I1046490);
nand I_61401 (I1045958,I1046490,I1046230);
nand I_61402 (I1045955,I1046473,I1046097);
not I_61403 (I1046579,I2690);
DFFARX1 I_61404 (I505829,I2683,I1046579,I1046605,);
DFFARX1 I_61405 (I505811,I2683,I1046579,I1046622,);
not I_61406 (I1046630,I1046622);
nor I_61407 (I1046547,I1046605,I1046630);
DFFARX1 I_61408 (I1046630,I2683,I1046579,I1046562,);
nor I_61409 (I1046675,I505817,I505820);
and I_61410 (I1046692,I1046675,I505808);
nor I_61411 (I1046709,I1046692,I505817);
not I_61412 (I1046726,I505817);
and I_61413 (I1046743,I1046726,I505826);
nand I_61414 (I1046760,I1046743,I505814);
nor I_61415 (I1046777,I1046726,I1046760);
DFFARX1 I_61416 (I1046777,I2683,I1046579,I1046544,);
not I_61417 (I1046808,I1046760);
nand I_61418 (I1046825,I1046630,I1046808);
nand I_61419 (I1046556,I1046692,I1046808);
DFFARX1 I_61420 (I1046726,I2683,I1046579,I1046571,);
not I_61421 (I1046870,I505811);
nor I_61422 (I1046887,I1046870,I505826);
nor I_61423 (I1046904,I1046887,I1046709);
DFFARX1 I_61424 (I1046904,I2683,I1046579,I1046568,);
not I_61425 (I1046935,I1046887);
DFFARX1 I_61426 (I1046935,I2683,I1046579,I1046961,);
not I_61427 (I1046969,I1046961);
nor I_61428 (I1046565,I1046969,I1046887);
nor I_61429 (I1047000,I1046870,I505823);
and I_61430 (I1047017,I1047000,I505832);
or I_61431 (I1047034,I1047017,I505808);
DFFARX1 I_61432 (I1047034,I2683,I1046579,I1047060,);
not I_61433 (I1047068,I1047060);
nand I_61434 (I1047085,I1047068,I1046808);
not I_61435 (I1046559,I1047085);
nand I_61436 (I1046553,I1047085,I1046825);
nand I_61437 (I1046550,I1047068,I1046692);
not I_61438 (I1047174,I2690);
DFFARX1 I_61439 (I26919,I2683,I1047174,I1047200,);
DFFARX1 I_61440 (I26901,I2683,I1047174,I1047217,);
not I_61441 (I1047225,I1047217);
nor I_61442 (I1047142,I1047200,I1047225);
DFFARX1 I_61443 (I1047225,I2683,I1047174,I1047157,);
nor I_61444 (I1047270,I26901,I26916);
and I_61445 (I1047287,I1047270,I26910);
nor I_61446 (I1047304,I1047287,I26901);
not I_61447 (I1047321,I26901);
and I_61448 (I1047338,I1047321,I26904);
nand I_61449 (I1047355,I1047338,I26907);
nor I_61450 (I1047372,I1047321,I1047355);
DFFARX1 I_61451 (I1047372,I2683,I1047174,I1047139,);
not I_61452 (I1047403,I1047355);
nand I_61453 (I1047420,I1047225,I1047403);
nand I_61454 (I1047151,I1047287,I1047403);
DFFARX1 I_61455 (I1047321,I2683,I1047174,I1047166,);
not I_61456 (I1047465,I26913);
nor I_61457 (I1047482,I1047465,I26904);
nor I_61458 (I1047499,I1047482,I1047304);
DFFARX1 I_61459 (I1047499,I2683,I1047174,I1047163,);
not I_61460 (I1047530,I1047482);
DFFARX1 I_61461 (I1047530,I2683,I1047174,I1047556,);
not I_61462 (I1047564,I1047556);
nor I_61463 (I1047160,I1047564,I1047482);
nor I_61464 (I1047595,I1047465,I26925);
and I_61465 (I1047612,I1047595,I26922);
or I_61466 (I1047629,I1047612,I26904);
DFFARX1 I_61467 (I1047629,I2683,I1047174,I1047655,);
not I_61468 (I1047663,I1047655);
nand I_61469 (I1047680,I1047663,I1047403);
not I_61470 (I1047154,I1047680);
nand I_61471 (I1047148,I1047680,I1047420);
nand I_61472 (I1047145,I1047663,I1047287);
not I_61473 (I1047769,I2690);
DFFARX1 I_61474 (I7456,I2683,I1047769,I1047795,);
DFFARX1 I_61475 (I7453,I2683,I1047769,I1047812,);
not I_61476 (I1047820,I1047812);
nor I_61477 (I1047737,I1047795,I1047820);
DFFARX1 I_61478 (I1047820,I2683,I1047769,I1047752,);
nor I_61479 (I1047865,I7471,I7468);
and I_61480 (I1047882,I1047865,I7459);
nor I_61481 (I1047899,I1047882,I7471);
not I_61482 (I1047916,I7471);
and I_61483 (I1047933,I1047916,I7456);
nand I_61484 (I1047950,I1047933,I7465);
nor I_61485 (I1047967,I1047916,I1047950);
DFFARX1 I_61486 (I1047967,I2683,I1047769,I1047734,);
not I_61487 (I1047998,I1047950);
nand I_61488 (I1048015,I1047820,I1047998);
nand I_61489 (I1047746,I1047882,I1047998);
DFFARX1 I_61490 (I1047916,I2683,I1047769,I1047761,);
not I_61491 (I1048060,I7474);
nor I_61492 (I1048077,I1048060,I7456);
nor I_61493 (I1048094,I1048077,I1047899);
DFFARX1 I_61494 (I1048094,I2683,I1047769,I1047758,);
not I_61495 (I1048125,I1048077);
DFFARX1 I_61496 (I1048125,I2683,I1047769,I1048151,);
not I_61497 (I1048159,I1048151);
nor I_61498 (I1047755,I1048159,I1048077);
nor I_61499 (I1048190,I1048060,I7453);
and I_61500 (I1048207,I1048190,I7459);
or I_61501 (I1048224,I1048207,I7462);
DFFARX1 I_61502 (I1048224,I2683,I1047769,I1048250,);
not I_61503 (I1048258,I1048250);
nand I_61504 (I1048275,I1048258,I1047998);
not I_61505 (I1047749,I1048275);
nand I_61506 (I1047743,I1048275,I1048015);
nand I_61507 (I1047740,I1048258,I1047882);
not I_61508 (I1048364,I2690);
DFFARX1 I_61509 (I126555,I2683,I1048364,I1048390,);
DFFARX1 I_61510 (I126558,I2683,I1048364,I1048407,);
not I_61511 (I1048415,I1048407);
nor I_61512 (I1048332,I1048390,I1048415);
DFFARX1 I_61513 (I1048415,I2683,I1048364,I1048347,);
nor I_61514 (I1048460,I126564,I126558);
and I_61515 (I1048477,I1048460,I126561);
nor I_61516 (I1048494,I1048477,I126564);
not I_61517 (I1048511,I126564);
and I_61518 (I1048528,I1048511,I126555);
nand I_61519 (I1048545,I1048528,I126573);
nor I_61520 (I1048562,I1048511,I1048545);
DFFARX1 I_61521 (I1048562,I2683,I1048364,I1048329,);
not I_61522 (I1048593,I1048545);
nand I_61523 (I1048610,I1048415,I1048593);
nand I_61524 (I1048341,I1048477,I1048593);
DFFARX1 I_61525 (I1048511,I2683,I1048364,I1048356,);
not I_61526 (I1048655,I126567);
nor I_61527 (I1048672,I1048655,I126555);
nor I_61528 (I1048689,I1048672,I1048494);
DFFARX1 I_61529 (I1048689,I2683,I1048364,I1048353,);
not I_61530 (I1048720,I1048672);
DFFARX1 I_61531 (I1048720,I2683,I1048364,I1048746,);
not I_61532 (I1048754,I1048746);
nor I_61533 (I1048350,I1048754,I1048672);
nor I_61534 (I1048785,I1048655,I126570);
and I_61535 (I1048802,I1048785,I126576);
or I_61536 (I1048819,I1048802,I126579);
DFFARX1 I_61537 (I1048819,I2683,I1048364,I1048845,);
not I_61538 (I1048853,I1048845);
nand I_61539 (I1048870,I1048853,I1048593);
not I_61540 (I1048344,I1048870);
nand I_61541 (I1048338,I1048870,I1048610);
nand I_61542 (I1048335,I1048853,I1048477);
not I_61543 (I1048959,I2690);
DFFARX1 I_61544 (I614493,I2683,I1048959,I1048985,);
DFFARX1 I_61545 (I614475,I2683,I1048959,I1049002,);
not I_61546 (I1049010,I1049002);
nor I_61547 (I1048927,I1048985,I1049010);
DFFARX1 I_61548 (I1049010,I2683,I1048959,I1048942,);
nor I_61549 (I1049055,I614481,I614484);
and I_61550 (I1049072,I1049055,I614472);
nor I_61551 (I1049089,I1049072,I614481);
not I_61552 (I1049106,I614481);
and I_61553 (I1049123,I1049106,I614490);
nand I_61554 (I1049140,I1049123,I614478);
nor I_61555 (I1049157,I1049106,I1049140);
DFFARX1 I_61556 (I1049157,I2683,I1048959,I1048924,);
not I_61557 (I1049188,I1049140);
nand I_61558 (I1049205,I1049010,I1049188);
nand I_61559 (I1048936,I1049072,I1049188);
DFFARX1 I_61560 (I1049106,I2683,I1048959,I1048951,);
not I_61561 (I1049250,I614475);
nor I_61562 (I1049267,I1049250,I614490);
nor I_61563 (I1049284,I1049267,I1049089);
DFFARX1 I_61564 (I1049284,I2683,I1048959,I1048948,);
not I_61565 (I1049315,I1049267);
DFFARX1 I_61566 (I1049315,I2683,I1048959,I1049341,);
not I_61567 (I1049349,I1049341);
nor I_61568 (I1048945,I1049349,I1049267);
nor I_61569 (I1049380,I1049250,I614487);
and I_61570 (I1049397,I1049380,I614496);
or I_61571 (I1049414,I1049397,I614472);
DFFARX1 I_61572 (I1049414,I2683,I1048959,I1049440,);
not I_61573 (I1049448,I1049440);
nand I_61574 (I1049465,I1049448,I1049188);
not I_61575 (I1048939,I1049465);
nand I_61576 (I1048933,I1049465,I1049205);
nand I_61577 (I1048930,I1049448,I1049072);
not I_61578 (I1049554,I2690);
DFFARX1 I_61579 (I91743,I2683,I1049554,I1049580,);
DFFARX1 I_61580 (I91731,I2683,I1049554,I1049597,);
not I_61581 (I1049605,I1049597);
nor I_61582 (I1049522,I1049580,I1049605);
DFFARX1 I_61583 (I1049605,I2683,I1049554,I1049537,);
nor I_61584 (I1049650,I91722,I91746);
and I_61585 (I1049667,I1049650,I91725);
nor I_61586 (I1049684,I1049667,I91722);
not I_61587 (I1049701,I91722);
and I_61588 (I1049718,I1049701,I91728);
nand I_61589 (I1049735,I1049718,I91740);
nor I_61590 (I1049752,I1049701,I1049735);
DFFARX1 I_61591 (I1049752,I2683,I1049554,I1049519,);
not I_61592 (I1049783,I1049735);
nand I_61593 (I1049800,I1049605,I1049783);
nand I_61594 (I1049531,I1049667,I1049783);
DFFARX1 I_61595 (I1049701,I2683,I1049554,I1049546,);
not I_61596 (I1049845,I91722);
nor I_61597 (I1049862,I1049845,I91728);
nor I_61598 (I1049879,I1049862,I1049684);
DFFARX1 I_61599 (I1049879,I2683,I1049554,I1049543,);
not I_61600 (I1049910,I1049862);
DFFARX1 I_61601 (I1049910,I2683,I1049554,I1049936,);
not I_61602 (I1049944,I1049936);
nor I_61603 (I1049540,I1049944,I1049862);
nor I_61604 (I1049975,I1049845,I91725);
and I_61605 (I1049992,I1049975,I91734);
or I_61606 (I1050009,I1049992,I91737);
DFFARX1 I_61607 (I1050009,I2683,I1049554,I1050035,);
not I_61608 (I1050043,I1050035);
nand I_61609 (I1050060,I1050043,I1049783);
not I_61610 (I1049534,I1050060);
nand I_61611 (I1049528,I1050060,I1049800);
nand I_61612 (I1049525,I1050043,I1049667);
not I_61613 (I1050149,I2690);
DFFARX1 I_61614 (I373106,I2683,I1050149,I1050175,);
DFFARX1 I_61615 (I373112,I2683,I1050149,I1050192,);
not I_61616 (I1050200,I1050192);
nor I_61617 (I1050117,I1050175,I1050200);
DFFARX1 I_61618 (I1050200,I2683,I1050149,I1050132,);
nor I_61619 (I1050245,I373121,I373106);
and I_61620 (I1050262,I1050245,I373133);
nor I_61621 (I1050279,I1050262,I373121);
not I_61622 (I1050296,I373121);
and I_61623 (I1050313,I1050296,I373109);
nand I_61624 (I1050330,I1050313,I373130);
nor I_61625 (I1050347,I1050296,I1050330);
DFFARX1 I_61626 (I1050347,I2683,I1050149,I1050114,);
not I_61627 (I1050378,I1050330);
nand I_61628 (I1050395,I1050200,I1050378);
nand I_61629 (I1050126,I1050262,I1050378);
DFFARX1 I_61630 (I1050296,I2683,I1050149,I1050141,);
not I_61631 (I1050440,I373118);
nor I_61632 (I1050457,I1050440,I373109);
nor I_61633 (I1050474,I1050457,I1050279);
DFFARX1 I_61634 (I1050474,I2683,I1050149,I1050138,);
not I_61635 (I1050505,I1050457);
DFFARX1 I_61636 (I1050505,I2683,I1050149,I1050531,);
not I_61637 (I1050539,I1050531);
nor I_61638 (I1050135,I1050539,I1050457);
nor I_61639 (I1050570,I1050440,I373115);
and I_61640 (I1050587,I1050570,I373127);
or I_61641 (I1050604,I1050587,I373124);
DFFARX1 I_61642 (I1050604,I2683,I1050149,I1050630,);
not I_61643 (I1050638,I1050630);
nand I_61644 (I1050655,I1050638,I1050378);
not I_61645 (I1050129,I1050655);
nand I_61646 (I1050123,I1050655,I1050395);
nand I_61647 (I1050120,I1050638,I1050262);
not I_61648 (I1050744,I2690);
DFFARX1 I_61649 (I142620,I2683,I1050744,I1050770,);
DFFARX1 I_61650 (I142623,I2683,I1050744,I1050787,);
not I_61651 (I1050795,I1050787);
nor I_61652 (I1050712,I1050770,I1050795);
DFFARX1 I_61653 (I1050795,I2683,I1050744,I1050727,);
nor I_61654 (I1050840,I142629,I142623);
and I_61655 (I1050857,I1050840,I142626);
nor I_61656 (I1050874,I1050857,I142629);
not I_61657 (I1050891,I142629);
and I_61658 (I1050908,I1050891,I142620);
nand I_61659 (I1050925,I1050908,I142638);
nor I_61660 (I1050942,I1050891,I1050925);
DFFARX1 I_61661 (I1050942,I2683,I1050744,I1050709,);
not I_61662 (I1050973,I1050925);
nand I_61663 (I1050990,I1050795,I1050973);
nand I_61664 (I1050721,I1050857,I1050973);
DFFARX1 I_61665 (I1050891,I2683,I1050744,I1050736,);
not I_61666 (I1051035,I142632);
nor I_61667 (I1051052,I1051035,I142620);
nor I_61668 (I1051069,I1051052,I1050874);
DFFARX1 I_61669 (I1051069,I2683,I1050744,I1050733,);
not I_61670 (I1051100,I1051052);
DFFARX1 I_61671 (I1051100,I2683,I1050744,I1051126,);
not I_61672 (I1051134,I1051126);
nor I_61673 (I1050730,I1051134,I1051052);
nor I_61674 (I1051165,I1051035,I142635);
and I_61675 (I1051182,I1051165,I142641);
or I_61676 (I1051199,I1051182,I142644);
DFFARX1 I_61677 (I1051199,I2683,I1050744,I1051225,);
not I_61678 (I1051233,I1051225);
nand I_61679 (I1051250,I1051233,I1050973);
not I_61680 (I1050724,I1051250);
nand I_61681 (I1050718,I1051250,I1050990);
nand I_61682 (I1050715,I1051233,I1050857);
not I_61683 (I1051339,I2690);
DFFARX1 I_61684 (I649671,I2683,I1051339,I1051365,);
DFFARX1 I_61685 (I649668,I2683,I1051339,I1051382,);
not I_61686 (I1051390,I1051382);
nor I_61687 (I1051307,I1051365,I1051390);
DFFARX1 I_61688 (I1051390,I2683,I1051339,I1051322,);
nor I_61689 (I1051435,I649683,I649665);
and I_61690 (I1051452,I1051435,I649662);
nor I_61691 (I1051469,I1051452,I649683);
not I_61692 (I1051486,I649683);
and I_61693 (I1051503,I1051486,I649668);
nand I_61694 (I1051520,I1051503,I649680);
nor I_61695 (I1051537,I1051486,I1051520);
DFFARX1 I_61696 (I1051537,I2683,I1051339,I1051304,);
not I_61697 (I1051568,I1051520);
nand I_61698 (I1051585,I1051390,I1051568);
nand I_61699 (I1051316,I1051452,I1051568);
DFFARX1 I_61700 (I1051486,I2683,I1051339,I1051331,);
not I_61701 (I1051630,I649674);
nor I_61702 (I1051647,I1051630,I649668);
nor I_61703 (I1051664,I1051647,I1051469);
DFFARX1 I_61704 (I1051664,I2683,I1051339,I1051328,);
not I_61705 (I1051695,I1051647);
DFFARX1 I_61706 (I1051695,I2683,I1051339,I1051721,);
not I_61707 (I1051729,I1051721);
nor I_61708 (I1051325,I1051729,I1051647);
nor I_61709 (I1051760,I1051630,I649662);
and I_61710 (I1051777,I1051760,I649677);
or I_61711 (I1051794,I1051777,I649665);
DFFARX1 I_61712 (I1051794,I2683,I1051339,I1051820,);
not I_61713 (I1051828,I1051820);
nand I_61714 (I1051845,I1051828,I1051568);
not I_61715 (I1051319,I1051845);
nand I_61716 (I1051313,I1051845,I1051585);
nand I_61717 (I1051310,I1051828,I1051452);
not I_61718 (I1051934,I2690);
DFFARX1 I_61719 (I566519,I2683,I1051934,I1051960,);
DFFARX1 I_61720 (I566501,I2683,I1051934,I1051977,);
not I_61721 (I1051985,I1051977);
nor I_61722 (I1051902,I1051960,I1051985);
DFFARX1 I_61723 (I1051985,I2683,I1051934,I1051917,);
nor I_61724 (I1052030,I566507,I566510);
and I_61725 (I1052047,I1052030,I566498);
nor I_61726 (I1052064,I1052047,I566507);
not I_61727 (I1052081,I566507);
and I_61728 (I1052098,I1052081,I566516);
nand I_61729 (I1052115,I1052098,I566504);
nor I_61730 (I1052132,I1052081,I1052115);
DFFARX1 I_61731 (I1052132,I2683,I1051934,I1051899,);
not I_61732 (I1052163,I1052115);
nand I_61733 (I1052180,I1051985,I1052163);
nand I_61734 (I1051911,I1052047,I1052163);
DFFARX1 I_61735 (I1052081,I2683,I1051934,I1051926,);
not I_61736 (I1052225,I566501);
nor I_61737 (I1052242,I1052225,I566516);
nor I_61738 (I1052259,I1052242,I1052064);
DFFARX1 I_61739 (I1052259,I2683,I1051934,I1051923,);
not I_61740 (I1052290,I1052242);
DFFARX1 I_61741 (I1052290,I2683,I1051934,I1052316,);
not I_61742 (I1052324,I1052316);
nor I_61743 (I1051920,I1052324,I1052242);
nor I_61744 (I1052355,I1052225,I566513);
and I_61745 (I1052372,I1052355,I566522);
or I_61746 (I1052389,I1052372,I566498);
DFFARX1 I_61747 (I1052389,I2683,I1051934,I1052415,);
not I_61748 (I1052423,I1052415);
nand I_61749 (I1052440,I1052423,I1052163);
not I_61750 (I1051914,I1052440);
nand I_61751 (I1051908,I1052440,I1052180);
nand I_61752 (I1051905,I1052423,I1052047);
not I_61753 (I1052529,I2690);
DFFARX1 I_61754 (I522591,I2683,I1052529,I1052555,);
DFFARX1 I_61755 (I522573,I2683,I1052529,I1052572,);
not I_61756 (I1052580,I1052572);
nor I_61757 (I1052497,I1052555,I1052580);
DFFARX1 I_61758 (I1052580,I2683,I1052529,I1052512,);
nor I_61759 (I1052625,I522579,I522582);
and I_61760 (I1052642,I1052625,I522570);
nor I_61761 (I1052659,I1052642,I522579);
not I_61762 (I1052676,I522579);
and I_61763 (I1052693,I1052676,I522588);
nand I_61764 (I1052710,I1052693,I522576);
nor I_61765 (I1052727,I1052676,I1052710);
DFFARX1 I_61766 (I1052727,I2683,I1052529,I1052494,);
not I_61767 (I1052758,I1052710);
nand I_61768 (I1052775,I1052580,I1052758);
nand I_61769 (I1052506,I1052642,I1052758);
DFFARX1 I_61770 (I1052676,I2683,I1052529,I1052521,);
not I_61771 (I1052820,I522573);
nor I_61772 (I1052837,I1052820,I522588);
nor I_61773 (I1052854,I1052837,I1052659);
DFFARX1 I_61774 (I1052854,I2683,I1052529,I1052518,);
not I_61775 (I1052885,I1052837);
DFFARX1 I_61776 (I1052885,I2683,I1052529,I1052911,);
not I_61777 (I1052919,I1052911);
nor I_61778 (I1052515,I1052919,I1052837);
nor I_61779 (I1052950,I1052820,I522585);
and I_61780 (I1052967,I1052950,I522594);
or I_61781 (I1052984,I1052967,I522570);
DFFARX1 I_61782 (I1052984,I2683,I1052529,I1053010,);
not I_61783 (I1053018,I1053010);
nand I_61784 (I1053035,I1053018,I1052758);
not I_61785 (I1052509,I1053035);
nand I_61786 (I1052503,I1053035,I1052775);
nand I_61787 (I1052500,I1053018,I1052642);
not I_61788 (I1053124,I2690);
DFFARX1 I_61789 (I429427,I2683,I1053124,I1053150,);
DFFARX1 I_61790 (I429430,I2683,I1053124,I1053167,);
not I_61791 (I1053175,I1053167);
nor I_61792 (I1053092,I1053150,I1053175);
DFFARX1 I_61793 (I1053175,I2683,I1053124,I1053107,);
nor I_61794 (I1053220,I429433,I429451);
and I_61795 (I1053237,I1053220,I429436);
nor I_61796 (I1053254,I1053237,I429433);
not I_61797 (I1053271,I429433);
and I_61798 (I1053288,I1053271,I429445);
nand I_61799 (I1053305,I1053288,I429448);
nor I_61800 (I1053322,I1053271,I1053305);
DFFARX1 I_61801 (I1053322,I2683,I1053124,I1053089,);
not I_61802 (I1053353,I1053305);
nand I_61803 (I1053370,I1053175,I1053353);
nand I_61804 (I1053101,I1053237,I1053353);
DFFARX1 I_61805 (I1053271,I2683,I1053124,I1053116,);
not I_61806 (I1053415,I429439);
nor I_61807 (I1053432,I1053415,I429445);
nor I_61808 (I1053449,I1053432,I1053254);
DFFARX1 I_61809 (I1053449,I2683,I1053124,I1053113,);
not I_61810 (I1053480,I1053432);
DFFARX1 I_61811 (I1053480,I2683,I1053124,I1053506,);
not I_61812 (I1053514,I1053506);
nor I_61813 (I1053110,I1053514,I1053432);
nor I_61814 (I1053545,I1053415,I429427);
and I_61815 (I1053562,I1053545,I429442);
or I_61816 (I1053579,I1053562,I429430);
DFFARX1 I_61817 (I1053579,I2683,I1053124,I1053605,);
not I_61818 (I1053613,I1053605);
nand I_61819 (I1053630,I1053613,I1053353);
not I_61820 (I1053104,I1053630);
nand I_61821 (I1053098,I1053630,I1053370);
nand I_61822 (I1053095,I1053613,I1053237);
not I_61823 (I1053719,I2690);
DFFARX1 I_61824 (I921257,I2683,I1053719,I1053745,);
DFFARX1 I_61825 (I921269,I2683,I1053719,I1053762,);
not I_61826 (I1053770,I1053762);
nor I_61827 (I1053687,I1053745,I1053770);
DFFARX1 I_61828 (I1053770,I2683,I1053719,I1053702,);
nor I_61829 (I1053815,I921266,I921260);
and I_61830 (I1053832,I1053815,I921254);
nor I_61831 (I1053849,I1053832,I921266);
not I_61832 (I1053866,I921266);
and I_61833 (I1053883,I1053866,I921263);
nand I_61834 (I1053900,I1053883,I921254);
nor I_61835 (I1053917,I1053866,I1053900);
DFFARX1 I_61836 (I1053917,I2683,I1053719,I1053684,);
not I_61837 (I1053948,I1053900);
nand I_61838 (I1053965,I1053770,I1053948);
nand I_61839 (I1053696,I1053832,I1053948);
DFFARX1 I_61840 (I1053866,I2683,I1053719,I1053711,);
not I_61841 (I1054010,I921278);
nor I_61842 (I1054027,I1054010,I921263);
nor I_61843 (I1054044,I1054027,I1053849);
DFFARX1 I_61844 (I1054044,I2683,I1053719,I1053708,);
not I_61845 (I1054075,I1054027);
DFFARX1 I_61846 (I1054075,I2683,I1053719,I1054101,);
not I_61847 (I1054109,I1054101);
nor I_61848 (I1053705,I1054109,I1054027);
nor I_61849 (I1054140,I1054010,I921272);
and I_61850 (I1054157,I1054140,I921275);
or I_61851 (I1054174,I1054157,I921257);
DFFARX1 I_61852 (I1054174,I2683,I1053719,I1054200,);
not I_61853 (I1054208,I1054200);
nand I_61854 (I1054225,I1054208,I1053948);
not I_61855 (I1053699,I1054225);
nand I_61856 (I1053693,I1054225,I1053965);
nand I_61857 (I1053690,I1054208,I1053832);
not I_61858 (I1054314,I2690);
DFFARX1 I_61859 (I618539,I2683,I1054314,I1054340,);
DFFARX1 I_61860 (I618521,I2683,I1054314,I1054357,);
not I_61861 (I1054365,I1054357);
nor I_61862 (I1054282,I1054340,I1054365);
DFFARX1 I_61863 (I1054365,I2683,I1054314,I1054297,);
nor I_61864 (I1054410,I618527,I618530);
and I_61865 (I1054427,I1054410,I618518);
nor I_61866 (I1054444,I1054427,I618527);
not I_61867 (I1054461,I618527);
and I_61868 (I1054478,I1054461,I618536);
nand I_61869 (I1054495,I1054478,I618524);
nor I_61870 (I1054512,I1054461,I1054495);
DFFARX1 I_61871 (I1054512,I2683,I1054314,I1054279,);
not I_61872 (I1054543,I1054495);
nand I_61873 (I1054560,I1054365,I1054543);
nand I_61874 (I1054291,I1054427,I1054543);
DFFARX1 I_61875 (I1054461,I2683,I1054314,I1054306,);
not I_61876 (I1054605,I618521);
nor I_61877 (I1054622,I1054605,I618536);
nor I_61878 (I1054639,I1054622,I1054444);
DFFARX1 I_61879 (I1054639,I2683,I1054314,I1054303,);
not I_61880 (I1054670,I1054622);
DFFARX1 I_61881 (I1054670,I2683,I1054314,I1054696,);
not I_61882 (I1054704,I1054696);
nor I_61883 (I1054300,I1054704,I1054622);
nor I_61884 (I1054735,I1054605,I618533);
and I_61885 (I1054752,I1054735,I618542);
or I_61886 (I1054769,I1054752,I618518);
DFFARX1 I_61887 (I1054769,I2683,I1054314,I1054795,);
not I_61888 (I1054803,I1054795);
nand I_61889 (I1054820,I1054803,I1054543);
not I_61890 (I1054294,I1054820);
nand I_61891 (I1054288,I1054820,I1054560);
nand I_61892 (I1054285,I1054803,I1054427);
not I_61893 (I1054909,I2690);
DFFARX1 I_61894 (I887733,I2683,I1054909,I1054935,);
DFFARX1 I_61895 (I887745,I2683,I1054909,I1054952,);
not I_61896 (I1054960,I1054952);
nor I_61897 (I1054877,I1054935,I1054960);
DFFARX1 I_61898 (I1054960,I2683,I1054909,I1054892,);
nor I_61899 (I1055005,I887742,I887736);
and I_61900 (I1055022,I1055005,I887730);
nor I_61901 (I1055039,I1055022,I887742);
not I_61902 (I1055056,I887742);
and I_61903 (I1055073,I1055056,I887739);
nand I_61904 (I1055090,I1055073,I887730);
nor I_61905 (I1055107,I1055056,I1055090);
DFFARX1 I_61906 (I1055107,I2683,I1054909,I1054874,);
not I_61907 (I1055138,I1055090);
nand I_61908 (I1055155,I1054960,I1055138);
nand I_61909 (I1054886,I1055022,I1055138);
DFFARX1 I_61910 (I1055056,I2683,I1054909,I1054901,);
not I_61911 (I1055200,I887754);
nor I_61912 (I1055217,I1055200,I887739);
nor I_61913 (I1055234,I1055217,I1055039);
DFFARX1 I_61914 (I1055234,I2683,I1054909,I1054898,);
not I_61915 (I1055265,I1055217);
DFFARX1 I_61916 (I1055265,I2683,I1054909,I1055291,);
not I_61917 (I1055299,I1055291);
nor I_61918 (I1054895,I1055299,I1055217);
nor I_61919 (I1055330,I1055200,I887748);
and I_61920 (I1055347,I1055330,I887751);
or I_61921 (I1055364,I1055347,I887733);
DFFARX1 I_61922 (I1055364,I2683,I1054909,I1055390,);
not I_61923 (I1055398,I1055390);
nand I_61924 (I1055415,I1055398,I1055138);
not I_61925 (I1054889,I1055415);
nand I_61926 (I1054883,I1055415,I1055155);
nand I_61927 (I1054880,I1055398,I1055022);
not I_61928 (I1055504,I2690);
DFFARX1 I_61929 (I821476,I2683,I1055504,I1055530,);
DFFARX1 I_61930 (I821467,I2683,I1055504,I1055547,);
not I_61931 (I1055555,I1055547);
nor I_61932 (I1055472,I1055530,I1055555);
DFFARX1 I_61933 (I1055555,I2683,I1055504,I1055487,);
nor I_61934 (I1055600,I821473,I821482);
and I_61935 (I1055617,I1055600,I821485);
nor I_61936 (I1055634,I1055617,I821473);
not I_61937 (I1055651,I821473);
and I_61938 (I1055668,I1055651,I821464);
nand I_61939 (I1055685,I1055668,I821470);
nor I_61940 (I1055702,I1055651,I1055685);
DFFARX1 I_61941 (I1055702,I2683,I1055504,I1055469,);
not I_61942 (I1055733,I1055685);
nand I_61943 (I1055750,I1055555,I1055733);
nand I_61944 (I1055481,I1055617,I1055733);
DFFARX1 I_61945 (I1055651,I2683,I1055504,I1055496,);
not I_61946 (I1055795,I821479);
nor I_61947 (I1055812,I1055795,I821464);
nor I_61948 (I1055829,I1055812,I1055634);
DFFARX1 I_61949 (I1055829,I2683,I1055504,I1055493,);
not I_61950 (I1055860,I1055812);
DFFARX1 I_61951 (I1055860,I2683,I1055504,I1055886,);
not I_61952 (I1055894,I1055886);
nor I_61953 (I1055490,I1055894,I1055812);
nor I_61954 (I1055925,I1055795,I821464);
and I_61955 (I1055942,I1055925,I821467);
or I_61956 (I1055959,I1055942,I821470);
DFFARX1 I_61957 (I1055959,I2683,I1055504,I1055985,);
not I_61958 (I1055993,I1055985);
nand I_61959 (I1056010,I1055993,I1055733);
not I_61960 (I1055484,I1056010);
nand I_61961 (I1055478,I1056010,I1055750);
nand I_61962 (I1055475,I1055993,I1055617);
not I_61963 (I1056099,I2690);
DFFARX1 I_61964 (I950735,I2683,I1056099,I1056125,);
DFFARX1 I_61965 (I950747,I2683,I1056099,I1056142,);
not I_61966 (I1056150,I1056142);
nor I_61967 (I1056067,I1056125,I1056150);
DFFARX1 I_61968 (I1056150,I2683,I1056099,I1056082,);
nor I_61969 (I1056195,I950744,I950738);
and I_61970 (I1056212,I1056195,I950732);
nor I_61971 (I1056229,I1056212,I950744);
not I_61972 (I1056246,I950744);
and I_61973 (I1056263,I1056246,I950741);
nand I_61974 (I1056280,I1056263,I950732);
nor I_61975 (I1056297,I1056246,I1056280);
DFFARX1 I_61976 (I1056297,I2683,I1056099,I1056064,);
not I_61977 (I1056328,I1056280);
nand I_61978 (I1056345,I1056150,I1056328);
nand I_61979 (I1056076,I1056212,I1056328);
DFFARX1 I_61980 (I1056246,I2683,I1056099,I1056091,);
not I_61981 (I1056390,I950756);
nor I_61982 (I1056407,I1056390,I950741);
nor I_61983 (I1056424,I1056407,I1056229);
DFFARX1 I_61984 (I1056424,I2683,I1056099,I1056088,);
not I_61985 (I1056455,I1056407);
DFFARX1 I_61986 (I1056455,I2683,I1056099,I1056481,);
not I_61987 (I1056489,I1056481);
nor I_61988 (I1056085,I1056489,I1056407);
nor I_61989 (I1056520,I1056390,I950750);
and I_61990 (I1056537,I1056520,I950753);
or I_61991 (I1056554,I1056537,I950735);
DFFARX1 I_61992 (I1056554,I2683,I1056099,I1056580,);
not I_61993 (I1056588,I1056580);
nand I_61994 (I1056605,I1056588,I1056328);
not I_61995 (I1056079,I1056605);
nand I_61996 (I1056073,I1056605,I1056345);
nand I_61997 (I1056070,I1056588,I1056212);
not I_61998 (I1056694,I2690);
DFFARX1 I_61999 (I572299,I2683,I1056694,I1056720,);
DFFARX1 I_62000 (I572281,I2683,I1056694,I1056737,);
not I_62001 (I1056745,I1056737);
nor I_62002 (I1056662,I1056720,I1056745);
DFFARX1 I_62003 (I1056745,I2683,I1056694,I1056677,);
nor I_62004 (I1056790,I572287,I572290);
and I_62005 (I1056807,I1056790,I572278);
nor I_62006 (I1056824,I1056807,I572287);
not I_62007 (I1056841,I572287);
and I_62008 (I1056858,I1056841,I572296);
nand I_62009 (I1056875,I1056858,I572284);
nor I_62010 (I1056892,I1056841,I1056875);
DFFARX1 I_62011 (I1056892,I2683,I1056694,I1056659,);
not I_62012 (I1056923,I1056875);
nand I_62013 (I1056940,I1056745,I1056923);
nand I_62014 (I1056671,I1056807,I1056923);
DFFARX1 I_62015 (I1056841,I2683,I1056694,I1056686,);
not I_62016 (I1056985,I572281);
nor I_62017 (I1057002,I1056985,I572296);
nor I_62018 (I1057019,I1057002,I1056824);
DFFARX1 I_62019 (I1057019,I2683,I1056694,I1056683,);
not I_62020 (I1057050,I1057002);
DFFARX1 I_62021 (I1057050,I2683,I1056694,I1057076,);
not I_62022 (I1057084,I1057076);
nor I_62023 (I1056680,I1057084,I1057002);
nor I_62024 (I1057115,I1056985,I572293);
and I_62025 (I1057132,I1057115,I572302);
or I_62026 (I1057149,I1057132,I572278);
DFFARX1 I_62027 (I1057149,I2683,I1056694,I1057175,);
not I_62028 (I1057183,I1057175);
nand I_62029 (I1057200,I1057183,I1056923);
not I_62030 (I1056674,I1057200);
nand I_62031 (I1056668,I1057200,I1056940);
nand I_62032 (I1056665,I1057183,I1056807);
not I_62033 (I1057289,I2690);
DFFARX1 I_62034 (I112894,I2683,I1057289,I1057315,);
DFFARX1 I_62035 (I112870,I2683,I1057289,I1057332,);
not I_62036 (I1057340,I1057332);
nor I_62037 (I1057257,I1057315,I1057340);
DFFARX1 I_62038 (I1057340,I2683,I1057289,I1057272,);
nor I_62039 (I1057385,I112897,I112879);
and I_62040 (I1057402,I1057385,I112891);
nor I_62041 (I1057419,I1057402,I112897);
not I_62042 (I1057436,I112897);
and I_62043 (I1057453,I1057436,I112873);
nand I_62044 (I1057470,I1057453,I112888);
nor I_62045 (I1057487,I1057436,I1057470);
DFFARX1 I_62046 (I1057487,I2683,I1057289,I1057254,);
not I_62047 (I1057518,I1057470);
nand I_62048 (I1057535,I1057340,I1057518);
nand I_62049 (I1057266,I1057402,I1057518);
DFFARX1 I_62050 (I1057436,I2683,I1057289,I1057281,);
not I_62051 (I1057580,I112882);
nor I_62052 (I1057597,I1057580,I112873);
nor I_62053 (I1057614,I1057597,I1057419);
DFFARX1 I_62054 (I1057614,I2683,I1057289,I1057278,);
not I_62055 (I1057645,I1057597);
DFFARX1 I_62056 (I1057645,I2683,I1057289,I1057671,);
not I_62057 (I1057679,I1057671);
nor I_62058 (I1057275,I1057679,I1057597);
nor I_62059 (I1057710,I1057580,I112885);
and I_62060 (I1057727,I1057710,I112876);
or I_62061 (I1057744,I1057727,I112870);
DFFARX1 I_62062 (I1057744,I2683,I1057289,I1057770,);
not I_62063 (I1057778,I1057770);
nand I_62064 (I1057795,I1057778,I1057518);
not I_62065 (I1057269,I1057795);
nand I_62066 (I1057263,I1057795,I1057535);
nand I_62067 (I1057260,I1057778,I1057402);
not I_62068 (I1057884,I2690);
DFFARX1 I_62069 (I208070,I2683,I1057884,I1057910,);
DFFARX1 I_62070 (I208073,I2683,I1057884,I1057927,);
not I_62071 (I1057935,I1057927);
nor I_62072 (I1057852,I1057910,I1057935);
DFFARX1 I_62073 (I1057935,I2683,I1057884,I1057867,);
nor I_62074 (I1057980,I208079,I208073);
and I_62075 (I1057997,I1057980,I208076);
nor I_62076 (I1058014,I1057997,I208079);
not I_62077 (I1058031,I208079);
and I_62078 (I1058048,I1058031,I208070);
nand I_62079 (I1058065,I1058048,I208088);
nor I_62080 (I1058082,I1058031,I1058065);
DFFARX1 I_62081 (I1058082,I2683,I1057884,I1057849,);
not I_62082 (I1058113,I1058065);
nand I_62083 (I1058130,I1057935,I1058113);
nand I_62084 (I1057861,I1057997,I1058113);
DFFARX1 I_62085 (I1058031,I2683,I1057884,I1057876,);
not I_62086 (I1058175,I208082);
nor I_62087 (I1058192,I1058175,I208070);
nor I_62088 (I1058209,I1058192,I1058014);
DFFARX1 I_62089 (I1058209,I2683,I1057884,I1057873,);
not I_62090 (I1058240,I1058192);
DFFARX1 I_62091 (I1058240,I2683,I1057884,I1058266,);
not I_62092 (I1058274,I1058266);
nor I_62093 (I1057870,I1058274,I1058192);
nor I_62094 (I1058305,I1058175,I208085);
and I_62095 (I1058322,I1058305,I208091);
or I_62096 (I1058339,I1058322,I208094);
DFFARX1 I_62097 (I1058339,I2683,I1057884,I1058365,);
not I_62098 (I1058373,I1058365);
nand I_62099 (I1058390,I1058373,I1058113);
not I_62100 (I1057864,I1058390);
nand I_62101 (I1057858,I1058390,I1058130);
nand I_62102 (I1057855,I1058373,I1057997);
not I_62103 (I1058479,I2690);
DFFARX1 I_62104 (I2428,I2683,I1058479,I1058505,);
DFFARX1 I_62105 (I1564,I2683,I1058479,I1058522,);
not I_62106 (I1058530,I1058522);
nor I_62107 (I1058447,I1058505,I1058530);
DFFARX1 I_62108 (I1058530,I2683,I1058479,I1058462,);
nor I_62109 (I1058575,I1932,I1788);
and I_62110 (I1058592,I1058575,I2316);
nor I_62111 (I1058609,I1058592,I1932);
not I_62112 (I1058626,I1932);
and I_62113 (I1058643,I1058626,I2604);
nand I_62114 (I1058660,I1058643,I1372);
nor I_62115 (I1058677,I1058626,I1058660);
DFFARX1 I_62116 (I1058677,I2683,I1058479,I1058444,);
not I_62117 (I1058708,I1058660);
nand I_62118 (I1058725,I1058530,I1058708);
nand I_62119 (I1058456,I1058592,I1058708);
DFFARX1 I_62120 (I1058626,I2683,I1058479,I1058471,);
not I_62121 (I1058770,I1548);
nor I_62122 (I1058787,I1058770,I2604);
nor I_62123 (I1058804,I1058787,I1058609);
DFFARX1 I_62124 (I1058804,I2683,I1058479,I1058468,);
not I_62125 (I1058835,I1058787);
DFFARX1 I_62126 (I1058835,I2683,I1058479,I1058861,);
not I_62127 (I1058869,I1058861);
nor I_62128 (I1058465,I1058869,I1058787);
nor I_62129 (I1058900,I1058770,I2500);
and I_62130 (I1058917,I1058900,I1604);
or I_62131 (I1058934,I1058917,I2244);
DFFARX1 I_62132 (I1058934,I2683,I1058479,I1058960,);
not I_62133 (I1058968,I1058960);
nand I_62134 (I1058985,I1058968,I1058708);
not I_62135 (I1058459,I1058985);
nand I_62136 (I1058453,I1058985,I1058725);
nand I_62137 (I1058450,I1058968,I1058592);
not I_62138 (I1059074,I2690);
DFFARX1 I_62139 (I12690,I2683,I1059074,I1059100,);
DFFARX1 I_62140 (I12672,I2683,I1059074,I1059117,);
not I_62141 (I1059125,I1059117);
nor I_62142 (I1059042,I1059100,I1059125);
DFFARX1 I_62143 (I1059125,I2683,I1059074,I1059057,);
nor I_62144 (I1059170,I12672,I12687);
and I_62145 (I1059187,I1059170,I12681);
nor I_62146 (I1059204,I1059187,I12672);
not I_62147 (I1059221,I12672);
and I_62148 (I1059238,I1059221,I12675);
nand I_62149 (I1059255,I1059238,I12678);
nor I_62150 (I1059272,I1059221,I1059255);
DFFARX1 I_62151 (I1059272,I2683,I1059074,I1059039,);
not I_62152 (I1059303,I1059255);
nand I_62153 (I1059320,I1059125,I1059303);
nand I_62154 (I1059051,I1059187,I1059303);
DFFARX1 I_62155 (I1059221,I2683,I1059074,I1059066,);
not I_62156 (I1059365,I12684);
nor I_62157 (I1059382,I1059365,I12675);
nor I_62158 (I1059399,I1059382,I1059204);
DFFARX1 I_62159 (I1059399,I2683,I1059074,I1059063,);
not I_62160 (I1059430,I1059382);
DFFARX1 I_62161 (I1059430,I2683,I1059074,I1059456,);
not I_62162 (I1059464,I1059456);
nor I_62163 (I1059060,I1059464,I1059382);
nor I_62164 (I1059495,I1059365,I12696);
and I_62165 (I1059512,I1059495,I12693);
or I_62166 (I1059529,I1059512,I12675);
DFFARX1 I_62167 (I1059529,I2683,I1059074,I1059555,);
not I_62168 (I1059563,I1059555);
nand I_62169 (I1059580,I1059563,I1059303);
not I_62170 (I1059054,I1059580);
nand I_62171 (I1059048,I1059580,I1059320);
nand I_62172 (I1059045,I1059563,I1059187);
not I_62173 (I1059669,I2690);
DFFARX1 I_62174 (I761987,I2683,I1059669,I1059695,);
DFFARX1 I_62175 (I762005,I2683,I1059669,I1059712,);
not I_62176 (I1059720,I1059712);
nor I_62177 (I1059637,I1059695,I1059720);
DFFARX1 I_62178 (I1059720,I2683,I1059669,I1059652,);
nor I_62179 (I1059765,I761984,I761996);
and I_62180 (I1059782,I1059765,I761981);
nor I_62181 (I1059799,I1059782,I761984);
not I_62182 (I1059816,I761984);
and I_62183 (I1059833,I1059816,I761990);
nand I_62184 (I1059850,I1059833,I762002);
nor I_62185 (I1059867,I1059816,I1059850);
DFFARX1 I_62186 (I1059867,I2683,I1059669,I1059634,);
not I_62187 (I1059898,I1059850);
nand I_62188 (I1059915,I1059720,I1059898);
nand I_62189 (I1059646,I1059782,I1059898);
DFFARX1 I_62190 (I1059816,I2683,I1059669,I1059661,);
not I_62191 (I1059960,I761993);
nor I_62192 (I1059977,I1059960,I761990);
nor I_62193 (I1059994,I1059977,I1059799);
DFFARX1 I_62194 (I1059994,I2683,I1059669,I1059658,);
not I_62195 (I1060025,I1059977);
DFFARX1 I_62196 (I1060025,I2683,I1059669,I1060051,);
not I_62197 (I1060059,I1060051);
nor I_62198 (I1059655,I1060059,I1059977);
nor I_62199 (I1060090,I1059960,I761981);
and I_62200 (I1060107,I1060090,I762008);
or I_62201 (I1060124,I1060107,I761999);
DFFARX1 I_62202 (I1060124,I2683,I1059669,I1060150,);
not I_62203 (I1060158,I1060150);
nand I_62204 (I1060175,I1060158,I1059898);
not I_62205 (I1059649,I1060175);
nand I_62206 (I1059643,I1060175,I1059915);
nand I_62207 (I1059640,I1060158,I1059782);
not I_62208 (I1060264,I2690);
DFFARX1 I_62209 (I386706,I2683,I1060264,I1060290,);
DFFARX1 I_62210 (I386712,I2683,I1060264,I1060307,);
not I_62211 (I1060315,I1060307);
nor I_62212 (I1060232,I1060290,I1060315);
DFFARX1 I_62213 (I1060315,I2683,I1060264,I1060247,);
nor I_62214 (I1060360,I386721,I386706);
and I_62215 (I1060377,I1060360,I386733);
nor I_62216 (I1060394,I1060377,I386721);
not I_62217 (I1060411,I386721);
and I_62218 (I1060428,I1060411,I386709);
nand I_62219 (I1060445,I1060428,I386730);
nor I_62220 (I1060462,I1060411,I1060445);
DFFARX1 I_62221 (I1060462,I2683,I1060264,I1060229,);
not I_62222 (I1060493,I1060445);
nand I_62223 (I1060510,I1060315,I1060493);
nand I_62224 (I1060241,I1060377,I1060493);
DFFARX1 I_62225 (I1060411,I2683,I1060264,I1060256,);
not I_62226 (I1060555,I386718);
nor I_62227 (I1060572,I1060555,I386709);
nor I_62228 (I1060589,I1060572,I1060394);
DFFARX1 I_62229 (I1060589,I2683,I1060264,I1060253,);
not I_62230 (I1060620,I1060572);
DFFARX1 I_62231 (I1060620,I2683,I1060264,I1060646,);
not I_62232 (I1060654,I1060646);
nor I_62233 (I1060250,I1060654,I1060572);
nor I_62234 (I1060685,I1060555,I386715);
and I_62235 (I1060702,I1060685,I386727);
or I_62236 (I1060719,I1060702,I386724);
DFFARX1 I_62237 (I1060719,I2683,I1060264,I1060745,);
not I_62238 (I1060753,I1060745);
nand I_62239 (I1060770,I1060753,I1060493);
not I_62240 (I1060244,I1060770);
nand I_62241 (I1060238,I1060770,I1060510);
nand I_62242 (I1060235,I1060753,I1060377);
not I_62243 (I1060859,I2690);
DFFARX1 I_62244 (I229052,I2683,I1060859,I1060885,);
DFFARX1 I_62245 (I229046,I2683,I1060859,I1060902,);
not I_62246 (I1060910,I1060902);
nor I_62247 (I1060827,I1060885,I1060910);
DFFARX1 I_62248 (I1060910,I2683,I1060859,I1060842,);
nor I_62249 (I1060955,I229034,I229055);
and I_62250 (I1060972,I1060955,I229049);
nor I_62251 (I1060989,I1060972,I229034);
not I_62252 (I1061006,I229034);
and I_62253 (I1061023,I1061006,I229031);
nand I_62254 (I1061040,I1061023,I229043);
nor I_62255 (I1061057,I1061006,I1061040);
DFFARX1 I_62256 (I1061057,I2683,I1060859,I1060824,);
not I_62257 (I1061088,I1061040);
nand I_62258 (I1061105,I1060910,I1061088);
nand I_62259 (I1060836,I1060972,I1061088);
DFFARX1 I_62260 (I1061006,I2683,I1060859,I1060851,);
not I_62261 (I1061150,I229058);
nor I_62262 (I1061167,I1061150,I229031);
nor I_62263 (I1061184,I1061167,I1060989);
DFFARX1 I_62264 (I1061184,I2683,I1060859,I1060848,);
not I_62265 (I1061215,I1061167);
DFFARX1 I_62266 (I1061215,I2683,I1060859,I1061241,);
not I_62267 (I1061249,I1061241);
nor I_62268 (I1060845,I1061249,I1061167);
nor I_62269 (I1061280,I1061150,I229040);
and I_62270 (I1061297,I1061280,I229037);
or I_62271 (I1061314,I1061297,I229031);
DFFARX1 I_62272 (I1061314,I2683,I1060859,I1061340,);
not I_62273 (I1061348,I1061340);
nand I_62274 (I1061365,I1061348,I1061088);
not I_62275 (I1060839,I1061365);
nand I_62276 (I1060833,I1061365,I1061105);
nand I_62277 (I1060830,I1061348,I1060972);
not I_62278 (I1061454,I2690);
DFFARX1 I_62279 (I51691,I2683,I1061454,I1061480,);
DFFARX1 I_62280 (I51679,I2683,I1061454,I1061497,);
not I_62281 (I1061505,I1061497);
nor I_62282 (I1061422,I1061480,I1061505);
DFFARX1 I_62283 (I1061505,I2683,I1061454,I1061437,);
nor I_62284 (I1061550,I51670,I51694);
and I_62285 (I1061567,I1061550,I51673);
nor I_62286 (I1061584,I1061567,I51670);
not I_62287 (I1061601,I51670);
and I_62288 (I1061618,I1061601,I51676);
nand I_62289 (I1061635,I1061618,I51688);
nor I_62290 (I1061652,I1061601,I1061635);
DFFARX1 I_62291 (I1061652,I2683,I1061454,I1061419,);
not I_62292 (I1061683,I1061635);
nand I_62293 (I1061700,I1061505,I1061683);
nand I_62294 (I1061431,I1061567,I1061683);
DFFARX1 I_62295 (I1061601,I2683,I1061454,I1061446,);
not I_62296 (I1061745,I51670);
nor I_62297 (I1061762,I1061745,I51676);
nor I_62298 (I1061779,I1061762,I1061584);
DFFARX1 I_62299 (I1061779,I2683,I1061454,I1061443,);
not I_62300 (I1061810,I1061762);
DFFARX1 I_62301 (I1061810,I2683,I1061454,I1061836,);
not I_62302 (I1061844,I1061836);
nor I_62303 (I1061440,I1061844,I1061762);
nor I_62304 (I1061875,I1061745,I51673);
and I_62305 (I1061892,I1061875,I51682);
or I_62306 (I1061909,I1061892,I51685);
DFFARX1 I_62307 (I1061909,I2683,I1061454,I1061935,);
not I_62308 (I1061943,I1061935);
nand I_62309 (I1061960,I1061943,I1061683);
not I_62310 (I1061434,I1061960);
nand I_62311 (I1061428,I1061960,I1061700);
nand I_62312 (I1061425,I1061943,I1061567);
not I_62313 (I1062049,I2690);
DFFARX1 I_62314 (I193790,I2683,I1062049,I1062075,);
DFFARX1 I_62315 (I193793,I2683,I1062049,I1062092,);
not I_62316 (I1062100,I1062092);
nor I_62317 (I1062017,I1062075,I1062100);
DFFARX1 I_62318 (I1062100,I2683,I1062049,I1062032,);
nor I_62319 (I1062145,I193799,I193793);
and I_62320 (I1062162,I1062145,I193796);
nor I_62321 (I1062179,I1062162,I193799);
not I_62322 (I1062196,I193799);
and I_62323 (I1062213,I1062196,I193790);
nand I_62324 (I1062230,I1062213,I193808);
nor I_62325 (I1062247,I1062196,I1062230);
DFFARX1 I_62326 (I1062247,I2683,I1062049,I1062014,);
not I_62327 (I1062278,I1062230);
nand I_62328 (I1062295,I1062100,I1062278);
nand I_62329 (I1062026,I1062162,I1062278);
DFFARX1 I_62330 (I1062196,I2683,I1062049,I1062041,);
not I_62331 (I1062340,I193802);
nor I_62332 (I1062357,I1062340,I193790);
nor I_62333 (I1062374,I1062357,I1062179);
DFFARX1 I_62334 (I1062374,I2683,I1062049,I1062038,);
not I_62335 (I1062405,I1062357);
DFFARX1 I_62336 (I1062405,I2683,I1062049,I1062431,);
not I_62337 (I1062439,I1062431);
nor I_62338 (I1062035,I1062439,I1062357);
nor I_62339 (I1062470,I1062340,I193805);
and I_62340 (I1062487,I1062470,I193811);
or I_62341 (I1062504,I1062487,I193814);
DFFARX1 I_62342 (I1062504,I2683,I1062049,I1062530,);
not I_62343 (I1062538,I1062530);
nand I_62344 (I1062555,I1062538,I1062278);
not I_62345 (I1062029,I1062555);
nand I_62346 (I1062023,I1062555,I1062295);
nand I_62347 (I1062020,I1062538,I1062162);
not I_62348 (I1062644,I2690);
DFFARX1 I_62349 (I385618,I2683,I1062644,I1062670,);
DFFARX1 I_62350 (I385624,I2683,I1062644,I1062687,);
not I_62351 (I1062695,I1062687);
nor I_62352 (I1062612,I1062670,I1062695);
DFFARX1 I_62353 (I1062695,I2683,I1062644,I1062627,);
nor I_62354 (I1062740,I385633,I385618);
and I_62355 (I1062757,I1062740,I385645);
nor I_62356 (I1062774,I1062757,I385633);
not I_62357 (I1062791,I385633);
and I_62358 (I1062808,I1062791,I385621);
nand I_62359 (I1062825,I1062808,I385642);
nor I_62360 (I1062842,I1062791,I1062825);
DFFARX1 I_62361 (I1062842,I2683,I1062644,I1062609,);
not I_62362 (I1062873,I1062825);
nand I_62363 (I1062890,I1062695,I1062873);
nand I_62364 (I1062621,I1062757,I1062873);
DFFARX1 I_62365 (I1062791,I2683,I1062644,I1062636,);
not I_62366 (I1062935,I385630);
nor I_62367 (I1062952,I1062935,I385621);
nor I_62368 (I1062969,I1062952,I1062774);
DFFARX1 I_62369 (I1062969,I2683,I1062644,I1062633,);
not I_62370 (I1063000,I1062952);
DFFARX1 I_62371 (I1063000,I2683,I1062644,I1063026,);
not I_62372 (I1063034,I1063026);
nor I_62373 (I1062630,I1063034,I1062952);
nor I_62374 (I1063065,I1062935,I385627);
and I_62375 (I1063082,I1063065,I385639);
or I_62376 (I1063099,I1063082,I385636);
DFFARX1 I_62377 (I1063099,I2683,I1062644,I1063125,);
not I_62378 (I1063133,I1063125);
nand I_62379 (I1063150,I1063133,I1062873);
not I_62380 (I1062624,I1063150);
nand I_62381 (I1062618,I1063150,I1062890);
nand I_62382 (I1062615,I1063133,I1062757);
not I_62383 (I1063239,I2690);
DFFARX1 I_62384 (I336114,I2683,I1063239,I1063265,);
DFFARX1 I_62385 (I336120,I2683,I1063239,I1063282,);
not I_62386 (I1063290,I1063282);
nor I_62387 (I1063207,I1063265,I1063290);
DFFARX1 I_62388 (I1063290,I2683,I1063239,I1063222,);
nor I_62389 (I1063335,I336129,I336114);
and I_62390 (I1063352,I1063335,I336141);
nor I_62391 (I1063369,I1063352,I336129);
not I_62392 (I1063386,I336129);
and I_62393 (I1063403,I1063386,I336117);
nand I_62394 (I1063420,I1063403,I336138);
nor I_62395 (I1063437,I1063386,I1063420);
DFFARX1 I_62396 (I1063437,I2683,I1063239,I1063204,);
not I_62397 (I1063468,I1063420);
nand I_62398 (I1063485,I1063290,I1063468);
nand I_62399 (I1063216,I1063352,I1063468);
DFFARX1 I_62400 (I1063386,I2683,I1063239,I1063231,);
not I_62401 (I1063530,I336126);
nor I_62402 (I1063547,I1063530,I336117);
nor I_62403 (I1063564,I1063547,I1063369);
DFFARX1 I_62404 (I1063564,I2683,I1063239,I1063228,);
not I_62405 (I1063595,I1063547);
DFFARX1 I_62406 (I1063595,I2683,I1063239,I1063621,);
not I_62407 (I1063629,I1063621);
nor I_62408 (I1063225,I1063629,I1063547);
nor I_62409 (I1063660,I1063530,I336123);
and I_62410 (I1063677,I1063660,I336135);
or I_62411 (I1063694,I1063677,I336132);
DFFARX1 I_62412 (I1063694,I2683,I1063239,I1063720,);
not I_62413 (I1063728,I1063720);
nand I_62414 (I1063745,I1063728,I1063468);
not I_62415 (I1063219,I1063745);
nand I_62416 (I1063213,I1063745,I1063485);
nand I_62417 (I1063210,I1063728,I1063352);
not I_62418 (I1063834,I2690);
DFFARX1 I_62419 (I413957,I2683,I1063834,I1063860,);
DFFARX1 I_62420 (I413960,I2683,I1063834,I1063877,);
not I_62421 (I1063885,I1063877);
nor I_62422 (I1063802,I1063860,I1063885);
DFFARX1 I_62423 (I1063885,I2683,I1063834,I1063817,);
nor I_62424 (I1063930,I413963,I413981);
and I_62425 (I1063947,I1063930,I413966);
nor I_62426 (I1063964,I1063947,I413963);
not I_62427 (I1063981,I413963);
and I_62428 (I1063998,I1063981,I413975);
nand I_62429 (I1064015,I1063998,I413978);
nor I_62430 (I1064032,I1063981,I1064015);
DFFARX1 I_62431 (I1064032,I2683,I1063834,I1063799,);
not I_62432 (I1064063,I1064015);
nand I_62433 (I1064080,I1063885,I1064063);
nand I_62434 (I1063811,I1063947,I1064063);
DFFARX1 I_62435 (I1063981,I2683,I1063834,I1063826,);
not I_62436 (I1064125,I413969);
nor I_62437 (I1064142,I1064125,I413975);
nor I_62438 (I1064159,I1064142,I1063964);
DFFARX1 I_62439 (I1064159,I2683,I1063834,I1063823,);
not I_62440 (I1064190,I1064142);
DFFARX1 I_62441 (I1064190,I2683,I1063834,I1064216,);
not I_62442 (I1064224,I1064216);
nor I_62443 (I1063820,I1064224,I1064142);
nor I_62444 (I1064255,I1064125,I413957);
and I_62445 (I1064272,I1064255,I413972);
or I_62446 (I1064289,I1064272,I413960);
DFFARX1 I_62447 (I1064289,I2683,I1063834,I1064315,);
not I_62448 (I1064323,I1064315);
nand I_62449 (I1064340,I1064323,I1064063);
not I_62450 (I1063814,I1064340);
nand I_62451 (I1063808,I1064340,I1064080);
nand I_62452 (I1063805,I1064323,I1063947);
not I_62453 (I1064429,I2690);
DFFARX1 I_62454 (I332306,I2683,I1064429,I1064455,);
DFFARX1 I_62455 (I332312,I2683,I1064429,I1064472,);
not I_62456 (I1064480,I1064472);
nor I_62457 (I1064397,I1064455,I1064480);
DFFARX1 I_62458 (I1064480,I2683,I1064429,I1064412,);
nor I_62459 (I1064525,I332321,I332306);
and I_62460 (I1064542,I1064525,I332333);
nor I_62461 (I1064559,I1064542,I332321);
not I_62462 (I1064576,I332321);
and I_62463 (I1064593,I1064576,I332309);
nand I_62464 (I1064610,I1064593,I332330);
nor I_62465 (I1064627,I1064576,I1064610);
DFFARX1 I_62466 (I1064627,I2683,I1064429,I1064394,);
not I_62467 (I1064658,I1064610);
nand I_62468 (I1064675,I1064480,I1064658);
nand I_62469 (I1064406,I1064542,I1064658);
DFFARX1 I_62470 (I1064576,I2683,I1064429,I1064421,);
not I_62471 (I1064720,I332318);
nor I_62472 (I1064737,I1064720,I332309);
nor I_62473 (I1064754,I1064737,I1064559);
DFFARX1 I_62474 (I1064754,I2683,I1064429,I1064418,);
not I_62475 (I1064785,I1064737);
DFFARX1 I_62476 (I1064785,I2683,I1064429,I1064811,);
not I_62477 (I1064819,I1064811);
nor I_62478 (I1064415,I1064819,I1064737);
nor I_62479 (I1064850,I1064720,I332315);
and I_62480 (I1064867,I1064850,I332327);
or I_62481 (I1064884,I1064867,I332324);
DFFARX1 I_62482 (I1064884,I2683,I1064429,I1064910,);
not I_62483 (I1064918,I1064910);
nand I_62484 (I1064935,I1064918,I1064658);
not I_62485 (I1064409,I1064935);
nand I_62486 (I1064403,I1064935,I1064675);
nand I_62487 (I1064400,I1064918,I1064542);
not I_62488 (I1065024,I2690);
DFFARX1 I_62489 (I52745,I2683,I1065024,I1065050,);
DFFARX1 I_62490 (I52733,I2683,I1065024,I1065067,);
not I_62491 (I1065075,I1065067);
nor I_62492 (I1064992,I1065050,I1065075);
DFFARX1 I_62493 (I1065075,I2683,I1065024,I1065007,);
nor I_62494 (I1065120,I52724,I52748);
and I_62495 (I1065137,I1065120,I52727);
nor I_62496 (I1065154,I1065137,I52724);
not I_62497 (I1065171,I52724);
and I_62498 (I1065188,I1065171,I52730);
nand I_62499 (I1065205,I1065188,I52742);
nor I_62500 (I1065222,I1065171,I1065205);
DFFARX1 I_62501 (I1065222,I2683,I1065024,I1064989,);
not I_62502 (I1065253,I1065205);
nand I_62503 (I1065270,I1065075,I1065253);
nand I_62504 (I1065001,I1065137,I1065253);
DFFARX1 I_62505 (I1065171,I2683,I1065024,I1065016,);
not I_62506 (I1065315,I52724);
nor I_62507 (I1065332,I1065315,I52730);
nor I_62508 (I1065349,I1065332,I1065154);
DFFARX1 I_62509 (I1065349,I2683,I1065024,I1065013,);
not I_62510 (I1065380,I1065332);
DFFARX1 I_62511 (I1065380,I2683,I1065024,I1065406,);
not I_62512 (I1065414,I1065406);
nor I_62513 (I1065010,I1065414,I1065332);
nor I_62514 (I1065445,I1065315,I52727);
and I_62515 (I1065462,I1065445,I52736);
or I_62516 (I1065479,I1065462,I52739);
DFFARX1 I_62517 (I1065479,I2683,I1065024,I1065505,);
not I_62518 (I1065513,I1065505);
nand I_62519 (I1065530,I1065513,I1065253);
not I_62520 (I1065004,I1065530);
nand I_62521 (I1064998,I1065530,I1065270);
nand I_62522 (I1064995,I1065513,I1065137);
not I_62523 (I1065619,I2690);
DFFARX1 I_62524 (I674967,I2683,I1065619,I1065645,);
DFFARX1 I_62525 (I674964,I2683,I1065619,I1065662,);
not I_62526 (I1065670,I1065662);
nor I_62527 (I1065587,I1065645,I1065670);
DFFARX1 I_62528 (I1065670,I2683,I1065619,I1065602,);
nor I_62529 (I1065715,I674979,I674961);
and I_62530 (I1065732,I1065715,I674958);
nor I_62531 (I1065749,I1065732,I674979);
not I_62532 (I1065766,I674979);
and I_62533 (I1065783,I1065766,I674964);
nand I_62534 (I1065800,I1065783,I674976);
nor I_62535 (I1065817,I1065766,I1065800);
DFFARX1 I_62536 (I1065817,I2683,I1065619,I1065584,);
not I_62537 (I1065848,I1065800);
nand I_62538 (I1065865,I1065670,I1065848);
nand I_62539 (I1065596,I1065732,I1065848);
DFFARX1 I_62540 (I1065766,I2683,I1065619,I1065611,);
not I_62541 (I1065910,I674970);
nor I_62542 (I1065927,I1065910,I674964);
nor I_62543 (I1065944,I1065927,I1065749);
DFFARX1 I_62544 (I1065944,I2683,I1065619,I1065608,);
not I_62545 (I1065975,I1065927);
DFFARX1 I_62546 (I1065975,I2683,I1065619,I1066001,);
not I_62547 (I1066009,I1066001);
nor I_62548 (I1065605,I1066009,I1065927);
nor I_62549 (I1066040,I1065910,I674958);
and I_62550 (I1066057,I1066040,I674973);
or I_62551 (I1066074,I1066057,I674961);
DFFARX1 I_62552 (I1066074,I2683,I1065619,I1066100,);
not I_62553 (I1066108,I1066100);
nand I_62554 (I1066125,I1066108,I1065848);
not I_62555 (I1065599,I1066125);
nand I_62556 (I1065593,I1066125,I1065865);
nand I_62557 (I1065590,I1066108,I1065732);
not I_62558 (I1066214,I2690);
DFFARX1 I_62559 (I928771,I2683,I1066214,I1066240,);
DFFARX1 I_62560 (I928783,I2683,I1066214,I1066257,);
not I_62561 (I1066265,I1066257);
nor I_62562 (I1066182,I1066240,I1066265);
DFFARX1 I_62563 (I1066265,I2683,I1066214,I1066197,);
nor I_62564 (I1066310,I928780,I928774);
and I_62565 (I1066327,I1066310,I928768);
nor I_62566 (I1066344,I1066327,I928780);
not I_62567 (I1066361,I928780);
and I_62568 (I1066378,I1066361,I928777);
nand I_62569 (I1066395,I1066378,I928768);
nor I_62570 (I1066412,I1066361,I1066395);
DFFARX1 I_62571 (I1066412,I2683,I1066214,I1066179,);
not I_62572 (I1066443,I1066395);
nand I_62573 (I1066460,I1066265,I1066443);
nand I_62574 (I1066191,I1066327,I1066443);
DFFARX1 I_62575 (I1066361,I2683,I1066214,I1066206,);
not I_62576 (I1066505,I928792);
nor I_62577 (I1066522,I1066505,I928777);
nor I_62578 (I1066539,I1066522,I1066344);
DFFARX1 I_62579 (I1066539,I2683,I1066214,I1066203,);
not I_62580 (I1066570,I1066522);
DFFARX1 I_62581 (I1066570,I2683,I1066214,I1066596,);
not I_62582 (I1066604,I1066596);
nor I_62583 (I1066200,I1066604,I1066522);
nor I_62584 (I1066635,I1066505,I928786);
and I_62585 (I1066652,I1066635,I928789);
or I_62586 (I1066669,I1066652,I928771);
DFFARX1 I_62587 (I1066669,I2683,I1066214,I1066695,);
not I_62588 (I1066703,I1066695);
nand I_62589 (I1066720,I1066703,I1066443);
not I_62590 (I1066194,I1066720);
nand I_62591 (I1066188,I1066720,I1066460);
nand I_62592 (I1066185,I1066703,I1066327);
not I_62593 (I1066809,I2690);
DFFARX1 I_62594 (I839759,I2683,I1066809,I1066835,);
DFFARX1 I_62595 (I839771,I2683,I1066809,I1066852,);
not I_62596 (I1066860,I1066852);
nor I_62597 (I1066777,I1066835,I1066860);
DFFARX1 I_62598 (I1066860,I2683,I1066809,I1066792,);
nor I_62599 (I1066905,I839768,I839762);
and I_62600 (I1066922,I1066905,I839756);
nor I_62601 (I1066939,I1066922,I839768);
not I_62602 (I1066956,I839768);
and I_62603 (I1066973,I1066956,I839765);
nand I_62604 (I1066990,I1066973,I839756);
nor I_62605 (I1067007,I1066956,I1066990);
DFFARX1 I_62606 (I1067007,I2683,I1066809,I1066774,);
not I_62607 (I1067038,I1066990);
nand I_62608 (I1067055,I1066860,I1067038);
nand I_62609 (I1066786,I1066922,I1067038);
DFFARX1 I_62610 (I1066956,I2683,I1066809,I1066801,);
not I_62611 (I1067100,I839780);
nor I_62612 (I1067117,I1067100,I839765);
nor I_62613 (I1067134,I1067117,I1066939);
DFFARX1 I_62614 (I1067134,I2683,I1066809,I1066798,);
not I_62615 (I1067165,I1067117);
DFFARX1 I_62616 (I1067165,I2683,I1066809,I1067191,);
not I_62617 (I1067199,I1067191);
nor I_62618 (I1066795,I1067199,I1067117);
nor I_62619 (I1067230,I1067100,I839774);
and I_62620 (I1067247,I1067230,I839777);
or I_62621 (I1067264,I1067247,I839759);
DFFARX1 I_62622 (I1067264,I2683,I1066809,I1067290,);
not I_62623 (I1067298,I1067290);
nand I_62624 (I1067315,I1067298,I1067038);
not I_62625 (I1066789,I1067315);
nand I_62626 (I1066783,I1067315,I1067055);
nand I_62627 (I1066780,I1067298,I1066922);
not I_62628 (I1067404,I2690);
DFFARX1 I_62629 (I61704,I2683,I1067404,I1067430,);
DFFARX1 I_62630 (I61692,I2683,I1067404,I1067447,);
not I_62631 (I1067455,I1067447);
nor I_62632 (I1067372,I1067430,I1067455);
DFFARX1 I_62633 (I1067455,I2683,I1067404,I1067387,);
nor I_62634 (I1067500,I61683,I61707);
and I_62635 (I1067517,I1067500,I61686);
nor I_62636 (I1067534,I1067517,I61683);
not I_62637 (I1067551,I61683);
and I_62638 (I1067568,I1067551,I61689);
nand I_62639 (I1067585,I1067568,I61701);
nor I_62640 (I1067602,I1067551,I1067585);
DFFARX1 I_62641 (I1067602,I2683,I1067404,I1067369,);
not I_62642 (I1067633,I1067585);
nand I_62643 (I1067650,I1067455,I1067633);
nand I_62644 (I1067381,I1067517,I1067633);
DFFARX1 I_62645 (I1067551,I2683,I1067404,I1067396,);
not I_62646 (I1067695,I61683);
nor I_62647 (I1067712,I1067695,I61689);
nor I_62648 (I1067729,I1067712,I1067534);
DFFARX1 I_62649 (I1067729,I2683,I1067404,I1067393,);
not I_62650 (I1067760,I1067712);
DFFARX1 I_62651 (I1067760,I2683,I1067404,I1067786,);
not I_62652 (I1067794,I1067786);
nor I_62653 (I1067390,I1067794,I1067712);
nor I_62654 (I1067825,I1067695,I61686);
and I_62655 (I1067842,I1067825,I61695);
or I_62656 (I1067859,I1067842,I61698);
DFFARX1 I_62657 (I1067859,I2683,I1067404,I1067885,);
not I_62658 (I1067893,I1067885);
nand I_62659 (I1067910,I1067893,I1067633);
not I_62660 (I1067384,I1067910);
nand I_62661 (I1067378,I1067910,I1067650);
nand I_62662 (I1067375,I1067893,I1067517);
not I_62663 (I1067999,I2690);
DFFARX1 I_62664 (I694993,I2683,I1067999,I1068025,);
DFFARX1 I_62665 (I694990,I2683,I1067999,I1068042,);
not I_62666 (I1068050,I1068042);
nor I_62667 (I1067967,I1068025,I1068050);
DFFARX1 I_62668 (I1068050,I2683,I1067999,I1067982,);
nor I_62669 (I1068095,I695005,I694987);
and I_62670 (I1068112,I1068095,I694984);
nor I_62671 (I1068129,I1068112,I695005);
not I_62672 (I1068146,I695005);
and I_62673 (I1068163,I1068146,I694990);
nand I_62674 (I1068180,I1068163,I695002);
nor I_62675 (I1068197,I1068146,I1068180);
DFFARX1 I_62676 (I1068197,I2683,I1067999,I1067964,);
not I_62677 (I1068228,I1068180);
nand I_62678 (I1068245,I1068050,I1068228);
nand I_62679 (I1067976,I1068112,I1068228);
DFFARX1 I_62680 (I1068146,I2683,I1067999,I1067991,);
not I_62681 (I1068290,I694996);
nor I_62682 (I1068307,I1068290,I694990);
nor I_62683 (I1068324,I1068307,I1068129);
DFFARX1 I_62684 (I1068324,I2683,I1067999,I1067988,);
not I_62685 (I1068355,I1068307);
DFFARX1 I_62686 (I1068355,I2683,I1067999,I1068381,);
not I_62687 (I1068389,I1068381);
nor I_62688 (I1067985,I1068389,I1068307);
nor I_62689 (I1068420,I1068290,I694984);
and I_62690 (I1068437,I1068420,I694999);
or I_62691 (I1068454,I1068437,I694987);
DFFARX1 I_62692 (I1068454,I2683,I1067999,I1068480,);
not I_62693 (I1068488,I1068480);
nand I_62694 (I1068505,I1068488,I1068228);
not I_62695 (I1067979,I1068505);
nand I_62696 (I1067973,I1068505,I1068245);
nand I_62697 (I1067970,I1068488,I1068112);
not I_62698 (I1068594,I2690);
DFFARX1 I_62699 (I1708,I2683,I1068594,I1068620,);
DFFARX1 I_62700 (I1460,I2683,I1068594,I1068637,);
not I_62701 (I1068645,I1068637);
nor I_62702 (I1068562,I1068620,I1068645);
DFFARX1 I_62703 (I1068645,I2683,I1068594,I1068577,);
nor I_62704 (I1068690,I2508,I2356);
and I_62705 (I1068707,I1068690,I1524);
nor I_62706 (I1068724,I1068707,I2508);
not I_62707 (I1068741,I2508);
and I_62708 (I1068758,I1068741,I2548);
nand I_62709 (I1068775,I1068758,I2620);
nor I_62710 (I1068792,I1068741,I1068775);
DFFARX1 I_62711 (I1068792,I2683,I1068594,I1068559,);
not I_62712 (I1068823,I1068775);
nand I_62713 (I1068840,I1068645,I1068823);
nand I_62714 (I1068571,I1068707,I1068823);
DFFARX1 I_62715 (I1068741,I2683,I1068594,I1068586,);
not I_62716 (I1068885,I2364);
nor I_62717 (I1068902,I1068885,I2548);
nor I_62718 (I1068919,I1068902,I1068724);
DFFARX1 I_62719 (I1068919,I2683,I1068594,I1068583,);
not I_62720 (I1068950,I1068902);
DFFARX1 I_62721 (I1068950,I2683,I1068594,I1068976,);
not I_62722 (I1068984,I1068976);
nor I_62723 (I1068580,I1068984,I1068902);
nor I_62724 (I1069015,I1068885,I1652);
and I_62725 (I1069032,I1069015,I2140);
or I_62726 (I1069049,I1069032,I1948);
DFFARX1 I_62727 (I1069049,I2683,I1068594,I1069075,);
not I_62728 (I1069083,I1069075);
nand I_62729 (I1069100,I1069083,I1068823);
not I_62730 (I1068574,I1069100);
nand I_62731 (I1068568,I1069100,I1068840);
nand I_62732 (I1068565,I1069083,I1068707);
not I_62733 (I1069189,I2690);
DFFARX1 I_62734 (I493113,I2683,I1069189,I1069215,);
DFFARX1 I_62735 (I493107,I2683,I1069189,I1069232,);
not I_62736 (I1069240,I1069232);
nor I_62737 (I1069157,I1069215,I1069240);
DFFARX1 I_62738 (I1069240,I2683,I1069189,I1069172,);
nor I_62739 (I1069285,I493104,I493095);
and I_62740 (I1069302,I1069285,I493092);
nor I_62741 (I1069319,I1069302,I493104);
not I_62742 (I1069336,I493104);
and I_62743 (I1069353,I1069336,I493098);
nand I_62744 (I1069370,I1069353,I493110);
nor I_62745 (I1069387,I1069336,I1069370);
DFFARX1 I_62746 (I1069387,I2683,I1069189,I1069154,);
not I_62747 (I1069418,I1069370);
nand I_62748 (I1069435,I1069240,I1069418);
nand I_62749 (I1069166,I1069302,I1069418);
DFFARX1 I_62750 (I1069336,I2683,I1069189,I1069181,);
not I_62751 (I1069480,I493116);
nor I_62752 (I1069497,I1069480,I493098);
nor I_62753 (I1069514,I1069497,I1069319);
DFFARX1 I_62754 (I1069514,I2683,I1069189,I1069178,);
not I_62755 (I1069545,I1069497);
DFFARX1 I_62756 (I1069545,I2683,I1069189,I1069571,);
not I_62757 (I1069579,I1069571);
nor I_62758 (I1069175,I1069579,I1069497);
nor I_62759 (I1069610,I1069480,I493095);
and I_62760 (I1069627,I1069610,I493101);
or I_62761 (I1069644,I1069627,I493092);
DFFARX1 I_62762 (I1069644,I2683,I1069189,I1069670,);
not I_62763 (I1069678,I1069670);
nand I_62764 (I1069695,I1069678,I1069418);
not I_62765 (I1069169,I1069695);
nand I_62766 (I1069163,I1069695,I1069435);
nand I_62767 (I1069160,I1069678,I1069302);
not I_62768 (I1069784,I2690);
DFFARX1 I_62769 (I249605,I2683,I1069784,I1069810,);
DFFARX1 I_62770 (I249599,I2683,I1069784,I1069827,);
not I_62771 (I1069835,I1069827);
nor I_62772 (I1069752,I1069810,I1069835);
DFFARX1 I_62773 (I1069835,I2683,I1069784,I1069767,);
nor I_62774 (I1069880,I249587,I249608);
and I_62775 (I1069897,I1069880,I249602);
nor I_62776 (I1069914,I1069897,I249587);
not I_62777 (I1069931,I249587);
and I_62778 (I1069948,I1069931,I249584);
nand I_62779 (I1069965,I1069948,I249596);
nor I_62780 (I1069982,I1069931,I1069965);
DFFARX1 I_62781 (I1069982,I2683,I1069784,I1069749,);
not I_62782 (I1070013,I1069965);
nand I_62783 (I1070030,I1069835,I1070013);
nand I_62784 (I1069761,I1069897,I1070013);
DFFARX1 I_62785 (I1069931,I2683,I1069784,I1069776,);
not I_62786 (I1070075,I249611);
nor I_62787 (I1070092,I1070075,I249584);
nor I_62788 (I1070109,I1070092,I1069914);
DFFARX1 I_62789 (I1070109,I2683,I1069784,I1069773,);
not I_62790 (I1070140,I1070092);
DFFARX1 I_62791 (I1070140,I2683,I1069784,I1070166,);
not I_62792 (I1070174,I1070166);
nor I_62793 (I1069770,I1070174,I1070092);
nor I_62794 (I1070205,I1070075,I249593);
and I_62795 (I1070222,I1070205,I249590);
or I_62796 (I1070239,I1070222,I249584);
DFFARX1 I_62797 (I1070239,I2683,I1069784,I1070265,);
not I_62798 (I1070273,I1070265);
nand I_62799 (I1070290,I1070273,I1070013);
not I_62800 (I1069764,I1070290);
nand I_62801 (I1069758,I1070290,I1070030);
nand I_62802 (I1069755,I1070273,I1069897);
not I_62803 (I1070379,I2690);
DFFARX1 I_62804 (I502361,I2683,I1070379,I1070405,);
DFFARX1 I_62805 (I502343,I2683,I1070379,I1070422,);
not I_62806 (I1070430,I1070422);
nor I_62807 (I1070347,I1070405,I1070430);
DFFARX1 I_62808 (I1070430,I2683,I1070379,I1070362,);
nor I_62809 (I1070475,I502349,I502352);
and I_62810 (I1070492,I1070475,I502340);
nor I_62811 (I1070509,I1070492,I502349);
not I_62812 (I1070526,I502349);
and I_62813 (I1070543,I1070526,I502358);
nand I_62814 (I1070560,I1070543,I502346);
nor I_62815 (I1070577,I1070526,I1070560);
DFFARX1 I_62816 (I1070577,I2683,I1070379,I1070344,);
not I_62817 (I1070608,I1070560);
nand I_62818 (I1070625,I1070430,I1070608);
nand I_62819 (I1070356,I1070492,I1070608);
DFFARX1 I_62820 (I1070526,I2683,I1070379,I1070371,);
not I_62821 (I1070670,I502343);
nor I_62822 (I1070687,I1070670,I502358);
nor I_62823 (I1070704,I1070687,I1070509);
DFFARX1 I_62824 (I1070704,I2683,I1070379,I1070368,);
not I_62825 (I1070735,I1070687);
DFFARX1 I_62826 (I1070735,I2683,I1070379,I1070761,);
not I_62827 (I1070769,I1070761);
nor I_62828 (I1070365,I1070769,I1070687);
nor I_62829 (I1070800,I1070670,I502355);
and I_62830 (I1070817,I1070800,I502364);
or I_62831 (I1070834,I1070817,I502340);
DFFARX1 I_62832 (I1070834,I2683,I1070379,I1070860,);
not I_62833 (I1070868,I1070860);
nand I_62834 (I1070885,I1070868,I1070608);
not I_62835 (I1070359,I1070885);
nand I_62836 (I1070353,I1070885,I1070625);
nand I_62837 (I1070350,I1070868,I1070492);
not I_62838 (I1070974,I2690);
DFFARX1 I_62839 (I730333,I2683,I1070974,I1071000,);
DFFARX1 I_62840 (I730351,I2683,I1070974,I1071017,);
not I_62841 (I1071025,I1071017);
nor I_62842 (I1070942,I1071000,I1071025);
DFFARX1 I_62843 (I1071025,I2683,I1070974,I1070957,);
nor I_62844 (I1071070,I730330,I730342);
and I_62845 (I1071087,I1071070,I730327);
nor I_62846 (I1071104,I1071087,I730330);
not I_62847 (I1071121,I730330);
and I_62848 (I1071138,I1071121,I730336);
nand I_62849 (I1071155,I1071138,I730348);
nor I_62850 (I1071172,I1071121,I1071155);
DFFARX1 I_62851 (I1071172,I2683,I1070974,I1070939,);
not I_62852 (I1071203,I1071155);
nand I_62853 (I1071220,I1071025,I1071203);
nand I_62854 (I1070951,I1071087,I1071203);
DFFARX1 I_62855 (I1071121,I2683,I1070974,I1070966,);
not I_62856 (I1071265,I730339);
nor I_62857 (I1071282,I1071265,I730336);
nor I_62858 (I1071299,I1071282,I1071104);
DFFARX1 I_62859 (I1071299,I2683,I1070974,I1070963,);
not I_62860 (I1071330,I1071282);
DFFARX1 I_62861 (I1071330,I2683,I1070974,I1071356,);
not I_62862 (I1071364,I1071356);
nor I_62863 (I1070960,I1071364,I1071282);
nor I_62864 (I1071395,I1071265,I730327);
and I_62865 (I1071412,I1071395,I730354);
or I_62866 (I1071429,I1071412,I730345);
DFFARX1 I_62867 (I1071429,I2683,I1070974,I1071455,);
not I_62868 (I1071463,I1071455);
nand I_62869 (I1071480,I1071463,I1071203);
not I_62870 (I1070954,I1071480);
nand I_62871 (I1070948,I1071480,I1071220);
nand I_62872 (I1070945,I1071463,I1071087);
not I_62873 (I1071569,I2690);
DFFARX1 I_62874 (I357330,I2683,I1071569,I1071595,);
DFFARX1 I_62875 (I357336,I2683,I1071569,I1071612,);
not I_62876 (I1071620,I1071612);
nor I_62877 (I1071537,I1071595,I1071620);
DFFARX1 I_62878 (I1071620,I2683,I1071569,I1071552,);
nor I_62879 (I1071665,I357345,I357330);
and I_62880 (I1071682,I1071665,I357357);
nor I_62881 (I1071699,I1071682,I357345);
not I_62882 (I1071716,I357345);
and I_62883 (I1071733,I1071716,I357333);
nand I_62884 (I1071750,I1071733,I357354);
nor I_62885 (I1071767,I1071716,I1071750);
DFFARX1 I_62886 (I1071767,I2683,I1071569,I1071534,);
not I_62887 (I1071798,I1071750);
nand I_62888 (I1071815,I1071620,I1071798);
nand I_62889 (I1071546,I1071682,I1071798);
DFFARX1 I_62890 (I1071716,I2683,I1071569,I1071561,);
not I_62891 (I1071860,I357342);
nor I_62892 (I1071877,I1071860,I357333);
nor I_62893 (I1071894,I1071877,I1071699);
DFFARX1 I_62894 (I1071894,I2683,I1071569,I1071558,);
not I_62895 (I1071925,I1071877);
DFFARX1 I_62896 (I1071925,I2683,I1071569,I1071951,);
not I_62897 (I1071959,I1071951);
nor I_62898 (I1071555,I1071959,I1071877);
nor I_62899 (I1071990,I1071860,I357339);
and I_62900 (I1072007,I1071990,I357351);
or I_62901 (I1072024,I1072007,I357348);
DFFARX1 I_62902 (I1072024,I2683,I1071569,I1072050,);
not I_62903 (I1072058,I1072050);
nand I_62904 (I1072075,I1072058,I1071798);
not I_62905 (I1071549,I1072075);
nand I_62906 (I1071543,I1072075,I1071815);
nand I_62907 (I1071540,I1072058,I1071682);
not I_62908 (I1072164,I2690);
DFFARX1 I_62909 (I295454,I2683,I1072164,I1072190,);
DFFARX1 I_62910 (I295448,I2683,I1072164,I1072207,);
not I_62911 (I1072215,I1072207);
nor I_62912 (I1072132,I1072190,I1072215);
DFFARX1 I_62913 (I1072215,I2683,I1072164,I1072147,);
nor I_62914 (I1072260,I295436,I295457);
and I_62915 (I1072277,I1072260,I295451);
nor I_62916 (I1072294,I1072277,I295436);
not I_62917 (I1072311,I295436);
and I_62918 (I1072328,I1072311,I295433);
nand I_62919 (I1072345,I1072328,I295445);
nor I_62920 (I1072362,I1072311,I1072345);
DFFARX1 I_62921 (I1072362,I2683,I1072164,I1072129,);
not I_62922 (I1072393,I1072345);
nand I_62923 (I1072410,I1072215,I1072393);
nand I_62924 (I1072141,I1072277,I1072393);
DFFARX1 I_62925 (I1072311,I2683,I1072164,I1072156,);
not I_62926 (I1072455,I295460);
nor I_62927 (I1072472,I1072455,I295433);
nor I_62928 (I1072489,I1072472,I1072294);
DFFARX1 I_62929 (I1072489,I2683,I1072164,I1072153,);
not I_62930 (I1072520,I1072472);
DFFARX1 I_62931 (I1072520,I2683,I1072164,I1072546,);
not I_62932 (I1072554,I1072546);
nor I_62933 (I1072150,I1072554,I1072472);
nor I_62934 (I1072585,I1072455,I295442);
and I_62935 (I1072602,I1072585,I295439);
or I_62936 (I1072619,I1072602,I295433);
DFFARX1 I_62937 (I1072619,I2683,I1072164,I1072645,);
not I_62938 (I1072653,I1072645);
nand I_62939 (I1072670,I1072653,I1072393);
not I_62940 (I1072144,I1072670);
nand I_62941 (I1072138,I1072670,I1072410);
nand I_62942 (I1072135,I1072653,I1072277);
not I_62943 (I1072759,I2690);
DFFARX1 I_62944 (I50637,I2683,I1072759,I1072785,);
DFFARX1 I_62945 (I50625,I2683,I1072759,I1072802,);
not I_62946 (I1072810,I1072802);
nor I_62947 (I1072727,I1072785,I1072810);
DFFARX1 I_62948 (I1072810,I2683,I1072759,I1072742,);
nor I_62949 (I1072855,I50616,I50640);
and I_62950 (I1072872,I1072855,I50619);
nor I_62951 (I1072889,I1072872,I50616);
not I_62952 (I1072906,I50616);
and I_62953 (I1072923,I1072906,I50622);
nand I_62954 (I1072940,I1072923,I50634);
nor I_62955 (I1072957,I1072906,I1072940);
DFFARX1 I_62956 (I1072957,I2683,I1072759,I1072724,);
not I_62957 (I1072988,I1072940);
nand I_62958 (I1073005,I1072810,I1072988);
nand I_62959 (I1072736,I1072872,I1072988);
DFFARX1 I_62960 (I1072906,I2683,I1072759,I1072751,);
not I_62961 (I1073050,I50616);
nor I_62962 (I1073067,I1073050,I50622);
nor I_62963 (I1073084,I1073067,I1072889);
DFFARX1 I_62964 (I1073084,I2683,I1072759,I1072748,);
not I_62965 (I1073115,I1073067);
DFFARX1 I_62966 (I1073115,I2683,I1072759,I1073141,);
not I_62967 (I1073149,I1073141);
nor I_62968 (I1072745,I1073149,I1073067);
nor I_62969 (I1073180,I1073050,I50619);
and I_62970 (I1073197,I1073180,I50628);
or I_62971 (I1073214,I1073197,I50631);
DFFARX1 I_62972 (I1073214,I2683,I1072759,I1073240,);
not I_62973 (I1073248,I1073240);
nand I_62974 (I1073265,I1073248,I1072988);
not I_62975 (I1072739,I1073265);
nand I_62976 (I1072733,I1073265,I1073005);
nand I_62977 (I1072730,I1073248,I1072872);
not I_62978 (I1073354,I2690);
DFFARX1 I_62979 (I314953,I2683,I1073354,I1073380,);
DFFARX1 I_62980 (I314947,I2683,I1073354,I1073397,);
not I_62981 (I1073405,I1073397);
nor I_62982 (I1073322,I1073380,I1073405);
DFFARX1 I_62983 (I1073405,I2683,I1073354,I1073337,);
nor I_62984 (I1073450,I314935,I314956);
and I_62985 (I1073467,I1073450,I314950);
nor I_62986 (I1073484,I1073467,I314935);
not I_62987 (I1073501,I314935);
and I_62988 (I1073518,I1073501,I314932);
nand I_62989 (I1073535,I1073518,I314944);
nor I_62990 (I1073552,I1073501,I1073535);
DFFARX1 I_62991 (I1073552,I2683,I1073354,I1073319,);
not I_62992 (I1073583,I1073535);
nand I_62993 (I1073600,I1073405,I1073583);
nand I_62994 (I1073331,I1073467,I1073583);
DFFARX1 I_62995 (I1073501,I2683,I1073354,I1073346,);
not I_62996 (I1073645,I314959);
nor I_62997 (I1073662,I1073645,I314932);
nor I_62998 (I1073679,I1073662,I1073484);
DFFARX1 I_62999 (I1073679,I2683,I1073354,I1073343,);
not I_63000 (I1073710,I1073662);
DFFARX1 I_63001 (I1073710,I2683,I1073354,I1073736,);
not I_63002 (I1073744,I1073736);
nor I_63003 (I1073340,I1073744,I1073662);
nor I_63004 (I1073775,I1073645,I314941);
and I_63005 (I1073792,I1073775,I314938);
or I_63006 (I1073809,I1073792,I314932);
DFFARX1 I_63007 (I1073809,I2683,I1073354,I1073835,);
not I_63008 (I1073843,I1073835);
nand I_63009 (I1073860,I1073843,I1073583);
not I_63010 (I1073334,I1073860);
nand I_63011 (I1073328,I1073860,I1073600);
nand I_63012 (I1073325,I1073843,I1073467);
not I_63013 (I1073949,I2690);
DFFARX1 I_63014 (I582703,I2683,I1073949,I1073975,);
DFFARX1 I_63015 (I582685,I2683,I1073949,I1073992,);
not I_63016 (I1074000,I1073992);
nor I_63017 (I1073917,I1073975,I1074000);
DFFARX1 I_63018 (I1074000,I2683,I1073949,I1073932,);
nor I_63019 (I1074045,I582691,I582694);
and I_63020 (I1074062,I1074045,I582682);
nor I_63021 (I1074079,I1074062,I582691);
not I_63022 (I1074096,I582691);
and I_63023 (I1074113,I1074096,I582700);
nand I_63024 (I1074130,I1074113,I582688);
nor I_63025 (I1074147,I1074096,I1074130);
DFFARX1 I_63026 (I1074147,I2683,I1073949,I1073914,);
not I_63027 (I1074178,I1074130);
nand I_63028 (I1074195,I1074000,I1074178);
nand I_63029 (I1073926,I1074062,I1074178);
DFFARX1 I_63030 (I1074096,I2683,I1073949,I1073941,);
not I_63031 (I1074240,I582685);
nor I_63032 (I1074257,I1074240,I582700);
nor I_63033 (I1074274,I1074257,I1074079);
DFFARX1 I_63034 (I1074274,I2683,I1073949,I1073938,);
not I_63035 (I1074305,I1074257);
DFFARX1 I_63036 (I1074305,I2683,I1073949,I1074331,);
not I_63037 (I1074339,I1074331);
nor I_63038 (I1073935,I1074339,I1074257);
nor I_63039 (I1074370,I1074240,I582697);
and I_63040 (I1074387,I1074370,I582706);
or I_63041 (I1074404,I1074387,I582682);
DFFARX1 I_63042 (I1074404,I2683,I1073949,I1074430,);
not I_63043 (I1074438,I1074430);
nand I_63044 (I1074455,I1074438,I1074178);
not I_63045 (I1073929,I1074455);
nand I_63046 (I1073923,I1074455,I1074195);
nand I_63047 (I1073920,I1074438,I1074062);
not I_63048 (I1074544,I2690);
DFFARX1 I_63049 (I589061,I2683,I1074544,I1074570,);
DFFARX1 I_63050 (I589043,I2683,I1074544,I1074587,);
not I_63051 (I1074595,I1074587);
nor I_63052 (I1074512,I1074570,I1074595);
DFFARX1 I_63053 (I1074595,I2683,I1074544,I1074527,);
nor I_63054 (I1074640,I589049,I589052);
and I_63055 (I1074657,I1074640,I589040);
nor I_63056 (I1074674,I1074657,I589049);
not I_63057 (I1074691,I589049);
and I_63058 (I1074708,I1074691,I589058);
nand I_63059 (I1074725,I1074708,I589046);
nor I_63060 (I1074742,I1074691,I1074725);
DFFARX1 I_63061 (I1074742,I2683,I1074544,I1074509,);
not I_63062 (I1074773,I1074725);
nand I_63063 (I1074790,I1074595,I1074773);
nand I_63064 (I1074521,I1074657,I1074773);
DFFARX1 I_63065 (I1074691,I2683,I1074544,I1074536,);
not I_63066 (I1074835,I589043);
nor I_63067 (I1074852,I1074835,I589058);
nor I_63068 (I1074869,I1074852,I1074674);
DFFARX1 I_63069 (I1074869,I2683,I1074544,I1074533,);
not I_63070 (I1074900,I1074852);
DFFARX1 I_63071 (I1074900,I2683,I1074544,I1074926,);
not I_63072 (I1074934,I1074926);
nor I_63073 (I1074530,I1074934,I1074852);
nor I_63074 (I1074965,I1074835,I589055);
and I_63075 (I1074982,I1074965,I589064);
or I_63076 (I1074999,I1074982,I589040);
DFFARX1 I_63077 (I1074999,I2683,I1074544,I1075025,);
not I_63078 (I1075033,I1075025);
nand I_63079 (I1075050,I1075033,I1074773);
not I_63080 (I1074524,I1075050);
nand I_63081 (I1074518,I1075050,I1074790);
nand I_63082 (I1074515,I1075033,I1074657);
not I_63083 (I1075139,I2690);
DFFARX1 I_63084 (I800719,I2683,I1075139,I1075165,);
DFFARX1 I_63085 (I800710,I2683,I1075139,I1075182,);
not I_63086 (I1075190,I1075182);
nor I_63087 (I1075107,I1075165,I1075190);
DFFARX1 I_63088 (I1075190,I2683,I1075139,I1075122,);
nor I_63089 (I1075235,I800716,I800725);
and I_63090 (I1075252,I1075235,I800728);
nor I_63091 (I1075269,I1075252,I800716);
not I_63092 (I1075286,I800716);
and I_63093 (I1075303,I1075286,I800707);
nand I_63094 (I1075320,I1075303,I800713);
nor I_63095 (I1075337,I1075286,I1075320);
DFFARX1 I_63096 (I1075337,I2683,I1075139,I1075104,);
not I_63097 (I1075368,I1075320);
nand I_63098 (I1075385,I1075190,I1075368);
nand I_63099 (I1075116,I1075252,I1075368);
DFFARX1 I_63100 (I1075286,I2683,I1075139,I1075131,);
not I_63101 (I1075430,I800722);
nor I_63102 (I1075447,I1075430,I800707);
nor I_63103 (I1075464,I1075447,I1075269);
DFFARX1 I_63104 (I1075464,I2683,I1075139,I1075128,);
not I_63105 (I1075495,I1075447);
DFFARX1 I_63106 (I1075495,I2683,I1075139,I1075521,);
not I_63107 (I1075529,I1075521);
nor I_63108 (I1075125,I1075529,I1075447);
nor I_63109 (I1075560,I1075430,I800707);
and I_63110 (I1075577,I1075560,I800710);
or I_63111 (I1075594,I1075577,I800713);
DFFARX1 I_63112 (I1075594,I2683,I1075139,I1075620,);
not I_63113 (I1075628,I1075620);
nand I_63114 (I1075645,I1075628,I1075368);
not I_63115 (I1075119,I1075645);
nand I_63116 (I1075113,I1075645,I1075385);
nand I_63117 (I1075110,I1075628,I1075252);
not I_63118 (I1075734,I2690);
DFFARX1 I_63119 (I46421,I2683,I1075734,I1075760,);
DFFARX1 I_63120 (I46409,I2683,I1075734,I1075777,);
not I_63121 (I1075785,I1075777);
nor I_63122 (I1075702,I1075760,I1075785);
DFFARX1 I_63123 (I1075785,I2683,I1075734,I1075717,);
nor I_63124 (I1075830,I46400,I46424);
and I_63125 (I1075847,I1075830,I46403);
nor I_63126 (I1075864,I1075847,I46400);
not I_63127 (I1075881,I46400);
and I_63128 (I1075898,I1075881,I46406);
nand I_63129 (I1075915,I1075898,I46418);
nor I_63130 (I1075932,I1075881,I1075915);
DFFARX1 I_63131 (I1075932,I2683,I1075734,I1075699,);
not I_63132 (I1075963,I1075915);
nand I_63133 (I1075980,I1075785,I1075963);
nand I_63134 (I1075711,I1075847,I1075963);
DFFARX1 I_63135 (I1075881,I2683,I1075734,I1075726,);
not I_63136 (I1076025,I46400);
nor I_63137 (I1076042,I1076025,I46406);
nor I_63138 (I1076059,I1076042,I1075864);
DFFARX1 I_63139 (I1076059,I2683,I1075734,I1075723,);
not I_63140 (I1076090,I1076042);
DFFARX1 I_63141 (I1076090,I2683,I1075734,I1076116,);
not I_63142 (I1076124,I1076116);
nor I_63143 (I1075720,I1076124,I1076042);
nor I_63144 (I1076155,I1076025,I46403);
and I_63145 (I1076172,I1076155,I46412);
or I_63146 (I1076189,I1076172,I46415);
DFFARX1 I_63147 (I1076189,I2683,I1075734,I1076215,);
not I_63148 (I1076223,I1076215);
nand I_63149 (I1076240,I1076223,I1075963);
not I_63150 (I1075714,I1076240);
nand I_63151 (I1075708,I1076240,I1075980);
nand I_63152 (I1075705,I1076223,I1075847);
not I_63153 (I1076329,I2690);
DFFARX1 I_63154 (I944377,I2683,I1076329,I1076355,);
DFFARX1 I_63155 (I944389,I2683,I1076329,I1076372,);
not I_63156 (I1076380,I1076372);
nor I_63157 (I1076297,I1076355,I1076380);
DFFARX1 I_63158 (I1076380,I2683,I1076329,I1076312,);
nor I_63159 (I1076425,I944386,I944380);
and I_63160 (I1076442,I1076425,I944374);
nor I_63161 (I1076459,I1076442,I944386);
not I_63162 (I1076476,I944386);
and I_63163 (I1076493,I1076476,I944383);
nand I_63164 (I1076510,I1076493,I944374);
nor I_63165 (I1076527,I1076476,I1076510);
DFFARX1 I_63166 (I1076527,I2683,I1076329,I1076294,);
not I_63167 (I1076558,I1076510);
nand I_63168 (I1076575,I1076380,I1076558);
nand I_63169 (I1076306,I1076442,I1076558);
DFFARX1 I_63170 (I1076476,I2683,I1076329,I1076321,);
not I_63171 (I1076620,I944398);
nor I_63172 (I1076637,I1076620,I944383);
nor I_63173 (I1076654,I1076637,I1076459);
DFFARX1 I_63174 (I1076654,I2683,I1076329,I1076318,);
not I_63175 (I1076685,I1076637);
DFFARX1 I_63176 (I1076685,I2683,I1076329,I1076711,);
not I_63177 (I1076719,I1076711);
nor I_63178 (I1076315,I1076719,I1076637);
nor I_63179 (I1076750,I1076620,I944392);
and I_63180 (I1076767,I1076750,I944395);
or I_63181 (I1076784,I1076767,I944377);
DFFARX1 I_63182 (I1076784,I2683,I1076329,I1076810,);
not I_63183 (I1076818,I1076810);
nand I_63184 (I1076835,I1076818,I1076558);
not I_63185 (I1076309,I1076835);
nand I_63186 (I1076303,I1076835,I1076575);
nand I_63187 (I1076300,I1076818,I1076442);
not I_63188 (I1076924,I2690);
DFFARX1 I_63189 (I670751,I2683,I1076924,I1076950,);
DFFARX1 I_63190 (I670748,I2683,I1076924,I1076967,);
not I_63191 (I1076975,I1076967);
nor I_63192 (I1076892,I1076950,I1076975);
DFFARX1 I_63193 (I1076975,I2683,I1076924,I1076907,);
nor I_63194 (I1077020,I670763,I670745);
and I_63195 (I1077037,I1077020,I670742);
nor I_63196 (I1077054,I1077037,I670763);
not I_63197 (I1077071,I670763);
and I_63198 (I1077088,I1077071,I670748);
nand I_63199 (I1077105,I1077088,I670760);
nor I_63200 (I1077122,I1077071,I1077105);
DFFARX1 I_63201 (I1077122,I2683,I1076924,I1076889,);
not I_63202 (I1077153,I1077105);
nand I_63203 (I1077170,I1076975,I1077153);
nand I_63204 (I1076901,I1077037,I1077153);
DFFARX1 I_63205 (I1077071,I2683,I1076924,I1076916,);
not I_63206 (I1077215,I670754);
nor I_63207 (I1077232,I1077215,I670748);
nor I_63208 (I1077249,I1077232,I1077054);
DFFARX1 I_63209 (I1077249,I2683,I1076924,I1076913,);
not I_63210 (I1077280,I1077232);
DFFARX1 I_63211 (I1077280,I2683,I1076924,I1077306,);
not I_63212 (I1077314,I1077306);
nor I_63213 (I1076910,I1077314,I1077232);
nor I_63214 (I1077345,I1077215,I670742);
and I_63215 (I1077362,I1077345,I670757);
or I_63216 (I1077379,I1077362,I670745);
DFFARX1 I_63217 (I1077379,I2683,I1076924,I1077405,);
not I_63218 (I1077413,I1077405);
nand I_63219 (I1077430,I1077413,I1077153);
not I_63220 (I1076904,I1077430);
nand I_63221 (I1076898,I1077430,I1077170);
nand I_63222 (I1076895,I1077413,I1077037);
not I_63223 (I1077519,I2690);
DFFARX1 I_63224 (I159875,I2683,I1077519,I1077545,);
DFFARX1 I_63225 (I159878,I2683,I1077519,I1077562,);
not I_63226 (I1077570,I1077562);
nor I_63227 (I1077487,I1077545,I1077570);
DFFARX1 I_63228 (I1077570,I2683,I1077519,I1077502,);
nor I_63229 (I1077615,I159884,I159878);
and I_63230 (I1077632,I1077615,I159881);
nor I_63231 (I1077649,I1077632,I159884);
not I_63232 (I1077666,I159884);
and I_63233 (I1077683,I1077666,I159875);
nand I_63234 (I1077700,I1077683,I159893);
nor I_63235 (I1077717,I1077666,I1077700);
DFFARX1 I_63236 (I1077717,I2683,I1077519,I1077484,);
not I_63237 (I1077748,I1077700);
nand I_63238 (I1077765,I1077570,I1077748);
nand I_63239 (I1077496,I1077632,I1077748);
DFFARX1 I_63240 (I1077666,I2683,I1077519,I1077511,);
not I_63241 (I1077810,I159887);
nor I_63242 (I1077827,I1077810,I159875);
nor I_63243 (I1077844,I1077827,I1077649);
DFFARX1 I_63244 (I1077844,I2683,I1077519,I1077508,);
not I_63245 (I1077875,I1077827);
DFFARX1 I_63246 (I1077875,I2683,I1077519,I1077901,);
not I_63247 (I1077909,I1077901);
nor I_63248 (I1077505,I1077909,I1077827);
nor I_63249 (I1077940,I1077810,I159890);
and I_63250 (I1077957,I1077940,I159896);
or I_63251 (I1077974,I1077957,I159899);
DFFARX1 I_63252 (I1077974,I2683,I1077519,I1078000,);
not I_63253 (I1078008,I1078000);
nand I_63254 (I1078025,I1078008,I1077748);
not I_63255 (I1077499,I1078025);
nand I_63256 (I1077493,I1078025,I1077765);
nand I_63257 (I1077490,I1078008,I1077632);
not I_63258 (I1078114,I2690);
DFFARX1 I_63259 (I396107,I2683,I1078114,I1078140,);
DFFARX1 I_63260 (I396110,I2683,I1078114,I1078157,);
not I_63261 (I1078165,I1078157);
nor I_63262 (I1078082,I1078140,I1078165);
DFFARX1 I_63263 (I1078165,I2683,I1078114,I1078097,);
nor I_63264 (I1078210,I396113,I396131);
and I_63265 (I1078227,I1078210,I396116);
nor I_63266 (I1078244,I1078227,I396113);
not I_63267 (I1078261,I396113);
and I_63268 (I1078278,I1078261,I396125);
nand I_63269 (I1078295,I1078278,I396128);
nor I_63270 (I1078312,I1078261,I1078295);
DFFARX1 I_63271 (I1078312,I2683,I1078114,I1078079,);
not I_63272 (I1078343,I1078295);
nand I_63273 (I1078360,I1078165,I1078343);
nand I_63274 (I1078091,I1078227,I1078343);
DFFARX1 I_63275 (I1078261,I2683,I1078114,I1078106,);
not I_63276 (I1078405,I396119);
nor I_63277 (I1078422,I1078405,I396125);
nor I_63278 (I1078439,I1078422,I1078244);
DFFARX1 I_63279 (I1078439,I2683,I1078114,I1078103,);
not I_63280 (I1078470,I1078422);
DFFARX1 I_63281 (I1078470,I2683,I1078114,I1078496,);
not I_63282 (I1078504,I1078496);
nor I_63283 (I1078100,I1078504,I1078422);
nor I_63284 (I1078535,I1078405,I396107);
and I_63285 (I1078552,I1078535,I396122);
or I_63286 (I1078569,I1078552,I396110);
DFFARX1 I_63287 (I1078569,I2683,I1078114,I1078595,);
not I_63288 (I1078603,I1078595);
nand I_63289 (I1078620,I1078603,I1078343);
not I_63290 (I1078094,I1078620);
nand I_63291 (I1078088,I1078620,I1078360);
nand I_63292 (I1078085,I1078603,I1078227);
not I_63293 (I1078709,I2690);
DFFARX1 I_63294 (I581547,I2683,I1078709,I1078735,);
DFFARX1 I_63295 (I581529,I2683,I1078709,I1078752,);
not I_63296 (I1078760,I1078752);
nor I_63297 (I1078677,I1078735,I1078760);
DFFARX1 I_63298 (I1078760,I2683,I1078709,I1078692,);
nor I_63299 (I1078805,I581535,I581538);
and I_63300 (I1078822,I1078805,I581526);
nor I_63301 (I1078839,I1078822,I581535);
not I_63302 (I1078856,I581535);
and I_63303 (I1078873,I1078856,I581544);
nand I_63304 (I1078890,I1078873,I581532);
nor I_63305 (I1078907,I1078856,I1078890);
DFFARX1 I_63306 (I1078907,I2683,I1078709,I1078674,);
not I_63307 (I1078938,I1078890);
nand I_63308 (I1078955,I1078760,I1078938);
nand I_63309 (I1078686,I1078822,I1078938);
DFFARX1 I_63310 (I1078856,I2683,I1078709,I1078701,);
not I_63311 (I1079000,I581529);
nor I_63312 (I1079017,I1079000,I581544);
nor I_63313 (I1079034,I1079017,I1078839);
DFFARX1 I_63314 (I1079034,I2683,I1078709,I1078698,);
not I_63315 (I1079065,I1079017);
DFFARX1 I_63316 (I1079065,I2683,I1078709,I1079091,);
not I_63317 (I1079099,I1079091);
nor I_63318 (I1078695,I1079099,I1079017);
nor I_63319 (I1079130,I1079000,I581541);
and I_63320 (I1079147,I1079130,I581550);
or I_63321 (I1079164,I1079147,I581526);
DFFARX1 I_63322 (I1079164,I2683,I1078709,I1079190,);
not I_63323 (I1079198,I1079190);
nand I_63324 (I1079215,I1079198,I1078938);
not I_63325 (I1078689,I1079215);
nand I_63326 (I1078683,I1079215,I1078955);
nand I_63327 (I1078680,I1079198,I1078822);
not I_63328 (I1079304,I2690);
DFFARX1 I_63329 (I231160,I2683,I1079304,I1079330,);
DFFARX1 I_63330 (I231154,I2683,I1079304,I1079347,);
not I_63331 (I1079355,I1079347);
nor I_63332 (I1079272,I1079330,I1079355);
DFFARX1 I_63333 (I1079355,I2683,I1079304,I1079287,);
nor I_63334 (I1079400,I231142,I231163);
and I_63335 (I1079417,I1079400,I231157);
nor I_63336 (I1079434,I1079417,I231142);
not I_63337 (I1079451,I231142);
and I_63338 (I1079468,I1079451,I231139);
nand I_63339 (I1079485,I1079468,I231151);
nor I_63340 (I1079502,I1079451,I1079485);
DFFARX1 I_63341 (I1079502,I2683,I1079304,I1079269,);
not I_63342 (I1079533,I1079485);
nand I_63343 (I1079550,I1079355,I1079533);
nand I_63344 (I1079281,I1079417,I1079533);
DFFARX1 I_63345 (I1079451,I2683,I1079304,I1079296,);
not I_63346 (I1079595,I231166);
nor I_63347 (I1079612,I1079595,I231139);
nor I_63348 (I1079629,I1079612,I1079434);
DFFARX1 I_63349 (I1079629,I2683,I1079304,I1079293,);
not I_63350 (I1079660,I1079612);
DFFARX1 I_63351 (I1079660,I2683,I1079304,I1079686,);
not I_63352 (I1079694,I1079686);
nor I_63353 (I1079290,I1079694,I1079612);
nor I_63354 (I1079725,I1079595,I231148);
and I_63355 (I1079742,I1079725,I231145);
or I_63356 (I1079759,I1079742,I231139);
DFFARX1 I_63357 (I1079759,I2683,I1079304,I1079785,);
not I_63358 (I1079793,I1079785);
nand I_63359 (I1079810,I1079793,I1079533);
not I_63360 (I1079284,I1079810);
nand I_63361 (I1079278,I1079810,I1079550);
nand I_63362 (I1079275,I1079793,I1079417);
not I_63363 (I1079899,I2690);
DFFARX1 I_63364 (I409197,I2683,I1079899,I1079925,);
DFFARX1 I_63365 (I409200,I2683,I1079899,I1079942,);
not I_63366 (I1079950,I1079942);
nor I_63367 (I1079867,I1079925,I1079950);
DFFARX1 I_63368 (I1079950,I2683,I1079899,I1079882,);
nor I_63369 (I1079995,I409203,I409221);
and I_63370 (I1080012,I1079995,I409206);
nor I_63371 (I1080029,I1080012,I409203);
not I_63372 (I1080046,I409203);
and I_63373 (I1080063,I1080046,I409215);
nand I_63374 (I1080080,I1080063,I409218);
nor I_63375 (I1080097,I1080046,I1080080);
DFFARX1 I_63376 (I1080097,I2683,I1079899,I1079864,);
not I_63377 (I1080128,I1080080);
nand I_63378 (I1080145,I1079950,I1080128);
nand I_63379 (I1079876,I1080012,I1080128);
DFFARX1 I_63380 (I1080046,I2683,I1079899,I1079891,);
not I_63381 (I1080190,I409209);
nor I_63382 (I1080207,I1080190,I409215);
nor I_63383 (I1080224,I1080207,I1080029);
DFFARX1 I_63384 (I1080224,I2683,I1079899,I1079888,);
not I_63385 (I1080255,I1080207);
DFFARX1 I_63386 (I1080255,I2683,I1079899,I1080281,);
not I_63387 (I1080289,I1080281);
nor I_63388 (I1079885,I1080289,I1080207);
nor I_63389 (I1080320,I1080190,I409197);
and I_63390 (I1080337,I1080320,I409212);
or I_63391 (I1080354,I1080337,I409200);
DFFARX1 I_63392 (I1080354,I2683,I1079899,I1080380,);
not I_63393 (I1080388,I1080380);
nand I_63394 (I1080405,I1080388,I1080128);
not I_63395 (I1079879,I1080405);
nand I_63396 (I1079873,I1080405,I1080145);
nand I_63397 (I1079870,I1080388,I1080012);
not I_63398 (I1080494,I2690);
DFFARX1 I_63399 (I181295,I2683,I1080494,I1080520,);
DFFARX1 I_63400 (I181298,I2683,I1080494,I1080537,);
not I_63401 (I1080545,I1080537);
nor I_63402 (I1080462,I1080520,I1080545);
DFFARX1 I_63403 (I1080545,I2683,I1080494,I1080477,);
nor I_63404 (I1080590,I181304,I181298);
and I_63405 (I1080607,I1080590,I181301);
nor I_63406 (I1080624,I1080607,I181304);
not I_63407 (I1080641,I181304);
and I_63408 (I1080658,I1080641,I181295);
nand I_63409 (I1080675,I1080658,I181313);
nor I_63410 (I1080692,I1080641,I1080675);
DFFARX1 I_63411 (I1080692,I2683,I1080494,I1080459,);
not I_63412 (I1080723,I1080675);
nand I_63413 (I1080740,I1080545,I1080723);
nand I_63414 (I1080471,I1080607,I1080723);
DFFARX1 I_63415 (I1080641,I2683,I1080494,I1080486,);
not I_63416 (I1080785,I181307);
nor I_63417 (I1080802,I1080785,I181295);
nor I_63418 (I1080819,I1080802,I1080624);
DFFARX1 I_63419 (I1080819,I2683,I1080494,I1080483,);
not I_63420 (I1080850,I1080802);
DFFARX1 I_63421 (I1080850,I2683,I1080494,I1080876,);
not I_63422 (I1080884,I1080876);
nor I_63423 (I1080480,I1080884,I1080802);
nor I_63424 (I1080915,I1080785,I181310);
and I_63425 (I1080932,I1080915,I181316);
or I_63426 (I1080949,I1080932,I181319);
DFFARX1 I_63427 (I1080949,I2683,I1080494,I1080975,);
not I_63428 (I1080983,I1080975);
nand I_63429 (I1081000,I1080983,I1080723);
not I_63430 (I1080474,I1081000);
nand I_63431 (I1080468,I1081000,I1080740);
nand I_63432 (I1080465,I1080983,I1080607);
not I_63433 (I1081089,I2690);
DFFARX1 I_63434 (I936863,I2683,I1081089,I1081115,);
DFFARX1 I_63435 (I936875,I2683,I1081089,I1081132,);
not I_63436 (I1081140,I1081132);
nor I_63437 (I1081057,I1081115,I1081140);
DFFARX1 I_63438 (I1081140,I2683,I1081089,I1081072,);
nor I_63439 (I1081185,I936872,I936866);
and I_63440 (I1081202,I1081185,I936860);
nor I_63441 (I1081219,I1081202,I936872);
not I_63442 (I1081236,I936872);
and I_63443 (I1081253,I1081236,I936869);
nand I_63444 (I1081270,I1081253,I936860);
nor I_63445 (I1081287,I1081236,I1081270);
DFFARX1 I_63446 (I1081287,I2683,I1081089,I1081054,);
not I_63447 (I1081318,I1081270);
nand I_63448 (I1081335,I1081140,I1081318);
nand I_63449 (I1081066,I1081202,I1081318);
DFFARX1 I_63450 (I1081236,I2683,I1081089,I1081081,);
not I_63451 (I1081380,I936884);
nor I_63452 (I1081397,I1081380,I936869);
nor I_63453 (I1081414,I1081397,I1081219);
DFFARX1 I_63454 (I1081414,I2683,I1081089,I1081078,);
not I_63455 (I1081445,I1081397);
DFFARX1 I_63456 (I1081445,I2683,I1081089,I1081471,);
not I_63457 (I1081479,I1081471);
nor I_63458 (I1081075,I1081479,I1081397);
nor I_63459 (I1081510,I1081380,I936878);
and I_63460 (I1081527,I1081510,I936881);
or I_63461 (I1081544,I1081527,I936863);
DFFARX1 I_63462 (I1081544,I2683,I1081089,I1081570,);
not I_63463 (I1081578,I1081570);
nand I_63464 (I1081595,I1081578,I1081318);
not I_63465 (I1081069,I1081595);
nand I_63466 (I1081063,I1081595,I1081335);
nand I_63467 (I1081060,I1081578,I1081202);
not I_63468 (I1081684,I2690);
DFFARX1 I_63469 (I199740,I2683,I1081684,I1081710,);
DFFARX1 I_63470 (I199743,I2683,I1081684,I1081727,);
not I_63471 (I1081735,I1081727);
nor I_63472 (I1081652,I1081710,I1081735);
DFFARX1 I_63473 (I1081735,I2683,I1081684,I1081667,);
nor I_63474 (I1081780,I199749,I199743);
and I_63475 (I1081797,I1081780,I199746);
nor I_63476 (I1081814,I1081797,I199749);
not I_63477 (I1081831,I199749);
and I_63478 (I1081848,I1081831,I199740);
nand I_63479 (I1081865,I1081848,I199758);
nor I_63480 (I1081882,I1081831,I1081865);
DFFARX1 I_63481 (I1081882,I2683,I1081684,I1081649,);
not I_63482 (I1081913,I1081865);
nand I_63483 (I1081930,I1081735,I1081913);
nand I_63484 (I1081661,I1081797,I1081913);
DFFARX1 I_63485 (I1081831,I2683,I1081684,I1081676,);
not I_63486 (I1081975,I199752);
nor I_63487 (I1081992,I1081975,I199740);
nor I_63488 (I1082009,I1081992,I1081814);
DFFARX1 I_63489 (I1082009,I2683,I1081684,I1081673,);
not I_63490 (I1082040,I1081992);
DFFARX1 I_63491 (I1082040,I2683,I1081684,I1082066,);
not I_63492 (I1082074,I1082066);
nor I_63493 (I1081670,I1082074,I1081992);
nor I_63494 (I1082105,I1081975,I199755);
and I_63495 (I1082122,I1082105,I199761);
or I_63496 (I1082139,I1082122,I199764);
DFFARX1 I_63497 (I1082139,I2683,I1081684,I1082165,);
not I_63498 (I1082173,I1082165);
nand I_63499 (I1082190,I1082173,I1081913);
not I_63500 (I1081664,I1082190);
nand I_63501 (I1081658,I1082190,I1081930);
nand I_63502 (I1081655,I1082173,I1081797);
not I_63503 (I1082279,I2690);
DFFARX1 I_63504 (I20595,I2683,I1082279,I1082305,);
DFFARX1 I_63505 (I20577,I2683,I1082279,I1082322,);
not I_63506 (I1082330,I1082322);
nor I_63507 (I1082247,I1082305,I1082330);
DFFARX1 I_63508 (I1082330,I2683,I1082279,I1082262,);
nor I_63509 (I1082375,I20577,I20592);
and I_63510 (I1082392,I1082375,I20586);
nor I_63511 (I1082409,I1082392,I20577);
not I_63512 (I1082426,I20577);
and I_63513 (I1082443,I1082426,I20580);
nand I_63514 (I1082460,I1082443,I20583);
nor I_63515 (I1082477,I1082426,I1082460);
DFFARX1 I_63516 (I1082477,I2683,I1082279,I1082244,);
not I_63517 (I1082508,I1082460);
nand I_63518 (I1082525,I1082330,I1082508);
nand I_63519 (I1082256,I1082392,I1082508);
DFFARX1 I_63520 (I1082426,I2683,I1082279,I1082271,);
not I_63521 (I1082570,I20589);
nor I_63522 (I1082587,I1082570,I20580);
nor I_63523 (I1082604,I1082587,I1082409);
DFFARX1 I_63524 (I1082604,I2683,I1082279,I1082268,);
not I_63525 (I1082635,I1082587);
DFFARX1 I_63526 (I1082635,I2683,I1082279,I1082661,);
not I_63527 (I1082669,I1082661);
nor I_63528 (I1082265,I1082669,I1082587);
nor I_63529 (I1082700,I1082570,I20601);
and I_63530 (I1082717,I1082700,I20598);
or I_63531 (I1082734,I1082717,I20580);
DFFARX1 I_63532 (I1082734,I2683,I1082279,I1082760,);
not I_63533 (I1082768,I1082760);
nand I_63534 (I1082785,I1082768,I1082508);
not I_63535 (I1082259,I1082785);
nand I_63536 (I1082253,I1082785,I1082525);
nand I_63537 (I1082250,I1082768,I1082392);
not I_63538 (I1082874,I2690);
DFFARX1 I_63539 (I309156,I2683,I1082874,I1082900,);
DFFARX1 I_63540 (I309150,I2683,I1082874,I1082917,);
not I_63541 (I1082925,I1082917);
nor I_63542 (I1082842,I1082900,I1082925);
DFFARX1 I_63543 (I1082925,I2683,I1082874,I1082857,);
nor I_63544 (I1082970,I309138,I309159);
and I_63545 (I1082987,I1082970,I309153);
nor I_63546 (I1083004,I1082987,I309138);
not I_63547 (I1083021,I309138);
and I_63548 (I1083038,I1083021,I309135);
nand I_63549 (I1083055,I1083038,I309147);
nor I_63550 (I1083072,I1083021,I1083055);
DFFARX1 I_63551 (I1083072,I2683,I1082874,I1082839,);
not I_63552 (I1083103,I1083055);
nand I_63553 (I1083120,I1082925,I1083103);
nand I_63554 (I1082851,I1082987,I1083103);
DFFARX1 I_63555 (I1083021,I2683,I1082874,I1082866,);
not I_63556 (I1083165,I309162);
nor I_63557 (I1083182,I1083165,I309135);
nor I_63558 (I1083199,I1083182,I1083004);
DFFARX1 I_63559 (I1083199,I2683,I1082874,I1082863,);
not I_63560 (I1083230,I1083182);
DFFARX1 I_63561 (I1083230,I2683,I1082874,I1083256,);
not I_63562 (I1083264,I1083256);
nor I_63563 (I1082860,I1083264,I1083182);
nor I_63564 (I1083295,I1083165,I309144);
and I_63565 (I1083312,I1083295,I309141);
or I_63566 (I1083329,I1083312,I309135);
DFFARX1 I_63567 (I1083329,I2683,I1082874,I1083355,);
not I_63568 (I1083363,I1083355);
nand I_63569 (I1083380,I1083363,I1083103);
not I_63570 (I1082854,I1083380);
nand I_63571 (I1082848,I1083380,I1083120);
nand I_63572 (I1082845,I1083363,I1082987);
not I_63573 (I1083469,I2690);
DFFARX1 I_63574 (I799597,I2683,I1083469,I1083495,);
DFFARX1 I_63575 (I799588,I2683,I1083469,I1083512,);
not I_63576 (I1083520,I1083512);
nor I_63577 (I1083437,I1083495,I1083520);
DFFARX1 I_63578 (I1083520,I2683,I1083469,I1083452,);
nor I_63579 (I1083565,I799594,I799603);
and I_63580 (I1083582,I1083565,I799606);
nor I_63581 (I1083599,I1083582,I799594);
not I_63582 (I1083616,I799594);
and I_63583 (I1083633,I1083616,I799585);
nand I_63584 (I1083650,I1083633,I799591);
nor I_63585 (I1083667,I1083616,I1083650);
DFFARX1 I_63586 (I1083667,I2683,I1083469,I1083434,);
not I_63587 (I1083698,I1083650);
nand I_63588 (I1083715,I1083520,I1083698);
nand I_63589 (I1083446,I1083582,I1083698);
DFFARX1 I_63590 (I1083616,I2683,I1083469,I1083461,);
not I_63591 (I1083760,I799600);
nor I_63592 (I1083777,I1083760,I799585);
nor I_63593 (I1083794,I1083777,I1083599);
DFFARX1 I_63594 (I1083794,I2683,I1083469,I1083458,);
not I_63595 (I1083825,I1083777);
DFFARX1 I_63596 (I1083825,I2683,I1083469,I1083851,);
not I_63597 (I1083859,I1083851);
nor I_63598 (I1083455,I1083859,I1083777);
nor I_63599 (I1083890,I1083760,I799585);
and I_63600 (I1083907,I1083890,I799588);
or I_63601 (I1083924,I1083907,I799591);
DFFARX1 I_63602 (I1083924,I2683,I1083469,I1083950,);
not I_63603 (I1083958,I1083950);
nand I_63604 (I1083975,I1083958,I1083698);
not I_63605 (I1083449,I1083975);
nand I_63606 (I1083443,I1083975,I1083715);
nand I_63607 (I1083440,I1083958,I1083582);
not I_63608 (I1084064,I2690);
DFFARX1 I_63609 (I4481,I2683,I1084064,I1084090,);
DFFARX1 I_63610 (I4478,I2683,I1084064,I1084107,);
not I_63611 (I1084115,I1084107);
nor I_63612 (I1084032,I1084090,I1084115);
DFFARX1 I_63613 (I1084115,I2683,I1084064,I1084047,);
nor I_63614 (I1084160,I4496,I4493);
and I_63615 (I1084177,I1084160,I4484);
nor I_63616 (I1084194,I1084177,I4496);
not I_63617 (I1084211,I4496);
and I_63618 (I1084228,I1084211,I4481);
nand I_63619 (I1084245,I1084228,I4490);
nor I_63620 (I1084262,I1084211,I1084245);
DFFARX1 I_63621 (I1084262,I2683,I1084064,I1084029,);
not I_63622 (I1084293,I1084245);
nand I_63623 (I1084310,I1084115,I1084293);
nand I_63624 (I1084041,I1084177,I1084293);
DFFARX1 I_63625 (I1084211,I2683,I1084064,I1084056,);
not I_63626 (I1084355,I4499);
nor I_63627 (I1084372,I1084355,I4481);
nor I_63628 (I1084389,I1084372,I1084194);
DFFARX1 I_63629 (I1084389,I2683,I1084064,I1084053,);
not I_63630 (I1084420,I1084372);
DFFARX1 I_63631 (I1084420,I2683,I1084064,I1084446,);
not I_63632 (I1084454,I1084446);
nor I_63633 (I1084050,I1084454,I1084372);
nor I_63634 (I1084485,I1084355,I4478);
and I_63635 (I1084502,I1084485,I4484);
or I_63636 (I1084519,I1084502,I4487);
DFFARX1 I_63637 (I1084519,I2683,I1084064,I1084545,);
not I_63638 (I1084553,I1084545);
nand I_63639 (I1084570,I1084553,I1084293);
not I_63640 (I1084044,I1084570);
nand I_63641 (I1084038,I1084570,I1084310);
nand I_63642 (I1084035,I1084553,I1084177);
not I_63643 (I1084659,I2690);
DFFARX1 I_63644 (I911431,I2683,I1084659,I1084685,);
DFFARX1 I_63645 (I911443,I2683,I1084659,I1084702,);
not I_63646 (I1084710,I1084702);
nor I_63647 (I1084627,I1084685,I1084710);
DFFARX1 I_63648 (I1084710,I2683,I1084659,I1084642,);
nor I_63649 (I1084755,I911440,I911434);
and I_63650 (I1084772,I1084755,I911428);
nor I_63651 (I1084789,I1084772,I911440);
not I_63652 (I1084806,I911440);
and I_63653 (I1084823,I1084806,I911437);
nand I_63654 (I1084840,I1084823,I911428);
nor I_63655 (I1084857,I1084806,I1084840);
DFFARX1 I_63656 (I1084857,I2683,I1084659,I1084624,);
not I_63657 (I1084888,I1084840);
nand I_63658 (I1084905,I1084710,I1084888);
nand I_63659 (I1084636,I1084772,I1084888);
DFFARX1 I_63660 (I1084806,I2683,I1084659,I1084651,);
not I_63661 (I1084950,I911452);
nor I_63662 (I1084967,I1084950,I911437);
nor I_63663 (I1084984,I1084967,I1084789);
DFFARX1 I_63664 (I1084984,I2683,I1084659,I1084648,);
not I_63665 (I1085015,I1084967);
DFFARX1 I_63666 (I1085015,I2683,I1084659,I1085041,);
not I_63667 (I1085049,I1085041);
nor I_63668 (I1084645,I1085049,I1084967);
nor I_63669 (I1085080,I1084950,I911446);
and I_63670 (I1085097,I1085080,I911449);
or I_63671 (I1085114,I1085097,I911431);
DFFARX1 I_63672 (I1085114,I2683,I1084659,I1085140,);
not I_63673 (I1085148,I1085140);
nand I_63674 (I1085165,I1085148,I1084888);
not I_63675 (I1084639,I1085165);
nand I_63676 (I1084633,I1085165,I1084905);
nand I_63677 (I1084630,I1085148,I1084772);
not I_63678 (I1085254,I2690);
DFFARX1 I_63679 (I796792,I2683,I1085254,I1085280,);
DFFARX1 I_63680 (I796783,I2683,I1085254,I1085297,);
not I_63681 (I1085305,I1085297);
nor I_63682 (I1085222,I1085280,I1085305);
DFFARX1 I_63683 (I1085305,I2683,I1085254,I1085237,);
nor I_63684 (I1085350,I796789,I796798);
and I_63685 (I1085367,I1085350,I796801);
nor I_63686 (I1085384,I1085367,I796789);
not I_63687 (I1085401,I796789);
and I_63688 (I1085418,I1085401,I796780);
nand I_63689 (I1085435,I1085418,I796786);
nor I_63690 (I1085452,I1085401,I1085435);
DFFARX1 I_63691 (I1085452,I2683,I1085254,I1085219,);
not I_63692 (I1085483,I1085435);
nand I_63693 (I1085500,I1085305,I1085483);
nand I_63694 (I1085231,I1085367,I1085483);
DFFARX1 I_63695 (I1085401,I2683,I1085254,I1085246,);
not I_63696 (I1085545,I796795);
nor I_63697 (I1085562,I1085545,I796780);
nor I_63698 (I1085579,I1085562,I1085384);
DFFARX1 I_63699 (I1085579,I2683,I1085254,I1085243,);
not I_63700 (I1085610,I1085562);
DFFARX1 I_63701 (I1085610,I2683,I1085254,I1085636,);
not I_63702 (I1085644,I1085636);
nor I_63703 (I1085240,I1085644,I1085562);
nor I_63704 (I1085675,I1085545,I796780);
and I_63705 (I1085692,I1085675,I796783);
or I_63706 (I1085709,I1085692,I796786);
DFFARX1 I_63707 (I1085709,I2683,I1085254,I1085735,);
not I_63708 (I1085743,I1085735);
nand I_63709 (I1085760,I1085743,I1085483);
not I_63710 (I1085234,I1085760);
nand I_63711 (I1085228,I1085760,I1085500);
nand I_63712 (I1085225,I1085743,I1085367);
not I_63713 (I1085849,I2690);
DFFARX1 I_63714 (I920679,I2683,I1085849,I1085875,);
DFFARX1 I_63715 (I920691,I2683,I1085849,I1085892,);
not I_63716 (I1085900,I1085892);
nor I_63717 (I1085817,I1085875,I1085900);
DFFARX1 I_63718 (I1085900,I2683,I1085849,I1085832,);
nor I_63719 (I1085945,I920688,I920682);
and I_63720 (I1085962,I1085945,I920676);
nor I_63721 (I1085979,I1085962,I920688);
not I_63722 (I1085996,I920688);
and I_63723 (I1086013,I1085996,I920685);
nand I_63724 (I1086030,I1086013,I920676);
nor I_63725 (I1086047,I1085996,I1086030);
DFFARX1 I_63726 (I1086047,I2683,I1085849,I1085814,);
not I_63727 (I1086078,I1086030);
nand I_63728 (I1086095,I1085900,I1086078);
nand I_63729 (I1085826,I1085962,I1086078);
DFFARX1 I_63730 (I1085996,I2683,I1085849,I1085841,);
not I_63731 (I1086140,I920700);
nor I_63732 (I1086157,I1086140,I920685);
nor I_63733 (I1086174,I1086157,I1085979);
DFFARX1 I_63734 (I1086174,I2683,I1085849,I1085838,);
not I_63735 (I1086205,I1086157);
DFFARX1 I_63736 (I1086205,I2683,I1085849,I1086231,);
not I_63737 (I1086239,I1086231);
nor I_63738 (I1085835,I1086239,I1086157);
nor I_63739 (I1086270,I1086140,I920694);
and I_63740 (I1086287,I1086270,I920697);
or I_63741 (I1086304,I1086287,I920679);
DFFARX1 I_63742 (I1086304,I2683,I1085849,I1086330,);
not I_63743 (I1086338,I1086330);
nand I_63744 (I1086355,I1086338,I1086078);
not I_63745 (I1085829,I1086355);
nand I_63746 (I1085823,I1086355,I1086095);
nand I_63747 (I1085820,I1086338,I1085962);
not I_63748 (I1086444,I2690);
DFFARX1 I_63749 (I214296,I2683,I1086444,I1086470,);
DFFARX1 I_63750 (I214290,I2683,I1086444,I1086487,);
not I_63751 (I1086495,I1086487);
nor I_63752 (I1086412,I1086470,I1086495);
DFFARX1 I_63753 (I1086495,I2683,I1086444,I1086427,);
nor I_63754 (I1086540,I214278,I214299);
and I_63755 (I1086557,I1086540,I214293);
nor I_63756 (I1086574,I1086557,I214278);
not I_63757 (I1086591,I214278);
and I_63758 (I1086608,I1086591,I214275);
nand I_63759 (I1086625,I1086608,I214287);
nor I_63760 (I1086642,I1086591,I1086625);
DFFARX1 I_63761 (I1086642,I2683,I1086444,I1086409,);
not I_63762 (I1086673,I1086625);
nand I_63763 (I1086690,I1086495,I1086673);
nand I_63764 (I1086421,I1086557,I1086673);
DFFARX1 I_63765 (I1086591,I2683,I1086444,I1086436,);
not I_63766 (I1086735,I214302);
nor I_63767 (I1086752,I1086735,I214275);
nor I_63768 (I1086769,I1086752,I1086574);
DFFARX1 I_63769 (I1086769,I2683,I1086444,I1086433,);
not I_63770 (I1086800,I1086752);
DFFARX1 I_63771 (I1086800,I2683,I1086444,I1086826,);
not I_63772 (I1086834,I1086826);
nor I_63773 (I1086430,I1086834,I1086752);
nor I_63774 (I1086865,I1086735,I214284);
and I_63775 (I1086882,I1086865,I214281);
or I_63776 (I1086899,I1086882,I214275);
DFFARX1 I_63777 (I1086899,I2683,I1086444,I1086925,);
not I_63778 (I1086933,I1086925);
nand I_63779 (I1086950,I1086933,I1086673);
not I_63780 (I1086424,I1086950);
nand I_63781 (I1086418,I1086950,I1086690);
nand I_63782 (I1086415,I1086933,I1086557);
not I_63783 (I1087039,I2690);
DFFARX1 I_63784 (I677602,I2683,I1087039,I1087065,);
DFFARX1 I_63785 (I677599,I2683,I1087039,I1087082,);
not I_63786 (I1087090,I1087082);
nor I_63787 (I1087007,I1087065,I1087090);
DFFARX1 I_63788 (I1087090,I2683,I1087039,I1087022,);
nor I_63789 (I1087135,I677614,I677596);
and I_63790 (I1087152,I1087135,I677593);
nor I_63791 (I1087169,I1087152,I677614);
not I_63792 (I1087186,I677614);
and I_63793 (I1087203,I1087186,I677599);
nand I_63794 (I1087220,I1087203,I677611);
nor I_63795 (I1087237,I1087186,I1087220);
DFFARX1 I_63796 (I1087237,I2683,I1087039,I1087004,);
not I_63797 (I1087268,I1087220);
nand I_63798 (I1087285,I1087090,I1087268);
nand I_63799 (I1087016,I1087152,I1087268);
DFFARX1 I_63800 (I1087186,I2683,I1087039,I1087031,);
not I_63801 (I1087330,I677605);
nor I_63802 (I1087347,I1087330,I677599);
nor I_63803 (I1087364,I1087347,I1087169);
DFFARX1 I_63804 (I1087364,I2683,I1087039,I1087028,);
not I_63805 (I1087395,I1087347);
DFFARX1 I_63806 (I1087395,I2683,I1087039,I1087421,);
not I_63807 (I1087429,I1087421);
nor I_63808 (I1087025,I1087429,I1087347);
nor I_63809 (I1087460,I1087330,I677593);
and I_63810 (I1087477,I1087460,I677608);
or I_63811 (I1087494,I1087477,I677596);
DFFARX1 I_63812 (I1087494,I2683,I1087039,I1087520,);
not I_63813 (I1087528,I1087520);
nand I_63814 (I1087545,I1087528,I1087268);
not I_63815 (I1087019,I1087545);
nand I_63816 (I1087013,I1087545,I1087285);
nand I_63817 (I1087010,I1087528,I1087152);
not I_63818 (I1087634,I2690);
DFFARX1 I_63819 (I148570,I2683,I1087634,I1087660,);
DFFARX1 I_63820 (I148573,I2683,I1087634,I1087677,);
not I_63821 (I1087685,I1087677);
nor I_63822 (I1087602,I1087660,I1087685);
DFFARX1 I_63823 (I1087685,I2683,I1087634,I1087617,);
nor I_63824 (I1087730,I148579,I148573);
and I_63825 (I1087747,I1087730,I148576);
nor I_63826 (I1087764,I1087747,I148579);
not I_63827 (I1087781,I148579);
and I_63828 (I1087798,I1087781,I148570);
nand I_63829 (I1087815,I1087798,I148588);
nor I_63830 (I1087832,I1087781,I1087815);
DFFARX1 I_63831 (I1087832,I2683,I1087634,I1087599,);
not I_63832 (I1087863,I1087815);
nand I_63833 (I1087880,I1087685,I1087863);
nand I_63834 (I1087611,I1087747,I1087863);
DFFARX1 I_63835 (I1087781,I2683,I1087634,I1087626,);
not I_63836 (I1087925,I148582);
nor I_63837 (I1087942,I1087925,I148570);
nor I_63838 (I1087959,I1087942,I1087764);
DFFARX1 I_63839 (I1087959,I2683,I1087634,I1087623,);
not I_63840 (I1087990,I1087942);
DFFARX1 I_63841 (I1087990,I2683,I1087634,I1088016,);
not I_63842 (I1088024,I1088016);
nor I_63843 (I1087620,I1088024,I1087942);
nor I_63844 (I1088055,I1087925,I148585);
and I_63845 (I1088072,I1088055,I148591);
or I_63846 (I1088089,I1088072,I148594);
DFFARX1 I_63847 (I1088089,I2683,I1087634,I1088115,);
not I_63848 (I1088123,I1088115);
nand I_63849 (I1088140,I1088123,I1087863);
not I_63850 (I1087614,I1088140);
nand I_63851 (I1087608,I1088140,I1087880);
nand I_63852 (I1087605,I1088123,I1087747);
not I_63853 (I1088229,I2690);
DFFARX1 I_63854 (I75406,I2683,I1088229,I1088255,);
DFFARX1 I_63855 (I75394,I2683,I1088229,I1088272,);
not I_63856 (I1088280,I1088272);
nor I_63857 (I1088197,I1088255,I1088280);
DFFARX1 I_63858 (I1088280,I2683,I1088229,I1088212,);
nor I_63859 (I1088325,I75385,I75409);
and I_63860 (I1088342,I1088325,I75388);
nor I_63861 (I1088359,I1088342,I75385);
not I_63862 (I1088376,I75385);
and I_63863 (I1088393,I1088376,I75391);
nand I_63864 (I1088410,I1088393,I75403);
nor I_63865 (I1088427,I1088376,I1088410);
DFFARX1 I_63866 (I1088427,I2683,I1088229,I1088194,);
not I_63867 (I1088458,I1088410);
nand I_63868 (I1088475,I1088280,I1088458);
nand I_63869 (I1088206,I1088342,I1088458);
DFFARX1 I_63870 (I1088376,I2683,I1088229,I1088221,);
not I_63871 (I1088520,I75385);
nor I_63872 (I1088537,I1088520,I75391);
nor I_63873 (I1088554,I1088537,I1088359);
DFFARX1 I_63874 (I1088554,I2683,I1088229,I1088218,);
not I_63875 (I1088585,I1088537);
DFFARX1 I_63876 (I1088585,I2683,I1088229,I1088611,);
not I_63877 (I1088619,I1088611);
nor I_63878 (I1088215,I1088619,I1088537);
nor I_63879 (I1088650,I1088520,I75388);
and I_63880 (I1088667,I1088650,I75397);
or I_63881 (I1088684,I1088667,I75400);
DFFARX1 I_63882 (I1088684,I2683,I1088229,I1088710,);
not I_63883 (I1088718,I1088710);
nand I_63884 (I1088735,I1088718,I1088458);
not I_63885 (I1088209,I1088735);
nand I_63886 (I1088203,I1088735,I1088475);
nand I_63887 (I1088200,I1088718,I1088342);
not I_63888 (I1088824,I2690);
DFFARX1 I_63889 (I202120,I2683,I1088824,I1088850,);
DFFARX1 I_63890 (I202123,I2683,I1088824,I1088867,);
not I_63891 (I1088875,I1088867);
nor I_63892 (I1088792,I1088850,I1088875);
DFFARX1 I_63893 (I1088875,I2683,I1088824,I1088807,);
nor I_63894 (I1088920,I202129,I202123);
and I_63895 (I1088937,I1088920,I202126);
nor I_63896 (I1088954,I1088937,I202129);
not I_63897 (I1088971,I202129);
and I_63898 (I1088988,I1088971,I202120);
nand I_63899 (I1089005,I1088988,I202138);
nor I_63900 (I1089022,I1088971,I1089005);
DFFARX1 I_63901 (I1089022,I2683,I1088824,I1088789,);
not I_63902 (I1089053,I1089005);
nand I_63903 (I1089070,I1088875,I1089053);
nand I_63904 (I1088801,I1088937,I1089053);
DFFARX1 I_63905 (I1088971,I2683,I1088824,I1088816,);
not I_63906 (I1089115,I202132);
nor I_63907 (I1089132,I1089115,I202120);
nor I_63908 (I1089149,I1089132,I1088954);
DFFARX1 I_63909 (I1089149,I2683,I1088824,I1088813,);
not I_63910 (I1089180,I1089132);
DFFARX1 I_63911 (I1089180,I2683,I1088824,I1089206,);
not I_63912 (I1089214,I1089206);
nor I_63913 (I1088810,I1089214,I1089132);
nor I_63914 (I1089245,I1089115,I202135);
and I_63915 (I1089262,I1089245,I202141);
or I_63916 (I1089279,I1089262,I202144);
DFFARX1 I_63917 (I1089279,I2683,I1088824,I1089305,);
not I_63918 (I1089313,I1089305);
nand I_63919 (I1089330,I1089313,I1089053);
not I_63920 (I1088804,I1089330);
nand I_63921 (I1088798,I1089330,I1089070);
nand I_63922 (I1088795,I1089313,I1088937);
not I_63923 (I1089419,I2690);
DFFARX1 I_63924 (I385074,I2683,I1089419,I1089445,);
DFFARX1 I_63925 (I385080,I2683,I1089419,I1089462,);
not I_63926 (I1089470,I1089462);
nor I_63927 (I1089387,I1089445,I1089470);
DFFARX1 I_63928 (I1089470,I2683,I1089419,I1089402,);
nor I_63929 (I1089515,I385089,I385074);
and I_63930 (I1089532,I1089515,I385101);
nor I_63931 (I1089549,I1089532,I385089);
not I_63932 (I1089566,I385089);
and I_63933 (I1089583,I1089566,I385077);
nand I_63934 (I1089600,I1089583,I385098);
nor I_63935 (I1089617,I1089566,I1089600);
DFFARX1 I_63936 (I1089617,I2683,I1089419,I1089384,);
not I_63937 (I1089648,I1089600);
nand I_63938 (I1089665,I1089470,I1089648);
nand I_63939 (I1089396,I1089532,I1089648);
DFFARX1 I_63940 (I1089566,I2683,I1089419,I1089411,);
not I_63941 (I1089710,I385086);
nor I_63942 (I1089727,I1089710,I385077);
nor I_63943 (I1089744,I1089727,I1089549);
DFFARX1 I_63944 (I1089744,I2683,I1089419,I1089408,);
not I_63945 (I1089775,I1089727);
DFFARX1 I_63946 (I1089775,I2683,I1089419,I1089801,);
not I_63947 (I1089809,I1089801);
nor I_63948 (I1089405,I1089809,I1089727);
nor I_63949 (I1089840,I1089710,I385083);
and I_63950 (I1089857,I1089840,I385095);
or I_63951 (I1089874,I1089857,I385092);
DFFARX1 I_63952 (I1089874,I2683,I1089419,I1089900,);
not I_63953 (I1089908,I1089900);
nand I_63954 (I1089925,I1089908,I1089648);
not I_63955 (I1089399,I1089925);
nand I_63956 (I1089393,I1089925,I1089665);
nand I_63957 (I1089390,I1089908,I1089532);
not I_63958 (I1090014,I2690);
DFFARX1 I_63959 (I745191,I2683,I1090014,I1090040,);
DFFARX1 I_63960 (I745209,I2683,I1090014,I1090057,);
not I_63961 (I1090065,I1090057);
nor I_63962 (I1089982,I1090040,I1090065);
DFFARX1 I_63963 (I1090065,I2683,I1090014,I1089997,);
nor I_63964 (I1090110,I745188,I745200);
and I_63965 (I1090127,I1090110,I745185);
nor I_63966 (I1090144,I1090127,I745188);
not I_63967 (I1090161,I745188);
and I_63968 (I1090178,I1090161,I745194);
nand I_63969 (I1090195,I1090178,I745206);
nor I_63970 (I1090212,I1090161,I1090195);
DFFARX1 I_63971 (I1090212,I2683,I1090014,I1089979,);
not I_63972 (I1090243,I1090195);
nand I_63973 (I1090260,I1090065,I1090243);
nand I_63974 (I1089991,I1090127,I1090243);
DFFARX1 I_63975 (I1090161,I2683,I1090014,I1090006,);
not I_63976 (I1090305,I745197);
nor I_63977 (I1090322,I1090305,I745194);
nor I_63978 (I1090339,I1090322,I1090144);
DFFARX1 I_63979 (I1090339,I2683,I1090014,I1090003,);
not I_63980 (I1090370,I1090322);
DFFARX1 I_63981 (I1090370,I2683,I1090014,I1090396,);
not I_63982 (I1090404,I1090396);
nor I_63983 (I1090000,I1090404,I1090322);
nor I_63984 (I1090435,I1090305,I745185);
and I_63985 (I1090452,I1090435,I745212);
or I_63986 (I1090469,I1090452,I745203);
DFFARX1 I_63987 (I1090469,I2683,I1090014,I1090495,);
not I_63988 (I1090503,I1090495);
nand I_63989 (I1090520,I1090503,I1090243);
not I_63990 (I1089994,I1090520);
nand I_63991 (I1089988,I1090520,I1090260);
nand I_63992 (I1089985,I1090503,I1090127);
not I_63993 (I1090609,I2690);
DFFARX1 I_63994 (I106499,I2683,I1090609,I1090635,);
DFFARX1 I_63995 (I106487,I2683,I1090609,I1090652,);
not I_63996 (I1090660,I1090652);
nor I_63997 (I1090577,I1090635,I1090660);
DFFARX1 I_63998 (I1090660,I2683,I1090609,I1090592,);
nor I_63999 (I1090705,I106478,I106502);
and I_64000 (I1090722,I1090705,I106481);
nor I_64001 (I1090739,I1090722,I106478);
not I_64002 (I1090756,I106478);
and I_64003 (I1090773,I1090756,I106484);
nand I_64004 (I1090790,I1090773,I106496);
nor I_64005 (I1090807,I1090756,I1090790);
DFFARX1 I_64006 (I1090807,I2683,I1090609,I1090574,);
not I_64007 (I1090838,I1090790);
nand I_64008 (I1090855,I1090660,I1090838);
nand I_64009 (I1090586,I1090722,I1090838);
DFFARX1 I_64010 (I1090756,I2683,I1090609,I1090601,);
not I_64011 (I1090900,I106478);
nor I_64012 (I1090917,I1090900,I106484);
nor I_64013 (I1090934,I1090917,I1090739);
DFFARX1 I_64014 (I1090934,I2683,I1090609,I1090598,);
not I_64015 (I1090965,I1090917);
DFFARX1 I_64016 (I1090965,I2683,I1090609,I1090991,);
not I_64017 (I1090999,I1090991);
nor I_64018 (I1090595,I1090999,I1090917);
nor I_64019 (I1091030,I1090900,I106481);
and I_64020 (I1091047,I1091030,I106490);
or I_64021 (I1091064,I1091047,I106493);
DFFARX1 I_64022 (I1091064,I2683,I1090609,I1091090,);
not I_64023 (I1091098,I1091090);
nand I_64024 (I1091115,I1091098,I1090838);
not I_64025 (I1090589,I1091115);
nand I_64026 (I1090583,I1091115,I1090855);
nand I_64027 (I1090580,I1091098,I1090722);
not I_64028 (I1091204,I2690);
DFFARX1 I_64029 (I601777,I2683,I1091204,I1091230,);
DFFARX1 I_64030 (I601759,I2683,I1091204,I1091247,);
not I_64031 (I1091255,I1091247);
nor I_64032 (I1091172,I1091230,I1091255);
DFFARX1 I_64033 (I1091255,I2683,I1091204,I1091187,);
nor I_64034 (I1091300,I601765,I601768);
and I_64035 (I1091317,I1091300,I601756);
nor I_64036 (I1091334,I1091317,I601765);
not I_64037 (I1091351,I601765);
and I_64038 (I1091368,I1091351,I601774);
nand I_64039 (I1091385,I1091368,I601762);
nor I_64040 (I1091402,I1091351,I1091385);
DFFARX1 I_64041 (I1091402,I2683,I1091204,I1091169,);
not I_64042 (I1091433,I1091385);
nand I_64043 (I1091450,I1091255,I1091433);
nand I_64044 (I1091181,I1091317,I1091433);
DFFARX1 I_64045 (I1091351,I2683,I1091204,I1091196,);
not I_64046 (I1091495,I601759);
nor I_64047 (I1091512,I1091495,I601774);
nor I_64048 (I1091529,I1091512,I1091334);
DFFARX1 I_64049 (I1091529,I2683,I1091204,I1091193,);
not I_64050 (I1091560,I1091512);
DFFARX1 I_64051 (I1091560,I2683,I1091204,I1091586,);
not I_64052 (I1091594,I1091586);
nor I_64053 (I1091190,I1091594,I1091512);
nor I_64054 (I1091625,I1091495,I601771);
and I_64055 (I1091642,I1091625,I601780);
or I_64056 (I1091659,I1091642,I601756);
DFFARX1 I_64057 (I1091659,I2683,I1091204,I1091685,);
not I_64058 (I1091693,I1091685);
nand I_64059 (I1091710,I1091693,I1091433);
not I_64060 (I1091184,I1091710);
nand I_64061 (I1091178,I1091710,I1091450);
nand I_64062 (I1091175,I1091693,I1091317);
not I_64063 (I1091799,I2690);
DFFARX1 I_64064 (I804646,I2683,I1091799,I1091825,);
DFFARX1 I_64065 (I804637,I2683,I1091799,I1091842,);
not I_64066 (I1091850,I1091842);
nor I_64067 (I1091767,I1091825,I1091850);
DFFARX1 I_64068 (I1091850,I2683,I1091799,I1091782,);
nor I_64069 (I1091895,I804643,I804652);
and I_64070 (I1091912,I1091895,I804655);
nor I_64071 (I1091929,I1091912,I804643);
not I_64072 (I1091946,I804643);
and I_64073 (I1091963,I1091946,I804634);
nand I_64074 (I1091980,I1091963,I804640);
nor I_64075 (I1091997,I1091946,I1091980);
DFFARX1 I_64076 (I1091997,I2683,I1091799,I1091764,);
not I_64077 (I1092028,I1091980);
nand I_64078 (I1092045,I1091850,I1092028);
nand I_64079 (I1091776,I1091912,I1092028);
DFFARX1 I_64080 (I1091946,I2683,I1091799,I1091791,);
not I_64081 (I1092090,I804649);
nor I_64082 (I1092107,I1092090,I804634);
nor I_64083 (I1092124,I1092107,I1091929);
DFFARX1 I_64084 (I1092124,I2683,I1091799,I1091788,);
not I_64085 (I1092155,I1092107);
DFFARX1 I_64086 (I1092155,I2683,I1091799,I1092181,);
not I_64087 (I1092189,I1092181);
nor I_64088 (I1091785,I1092189,I1092107);
nor I_64089 (I1092220,I1092090,I804634);
and I_64090 (I1092237,I1092220,I804637);
or I_64091 (I1092254,I1092237,I804640);
DFFARX1 I_64092 (I1092254,I2683,I1091799,I1092280,);
not I_64093 (I1092288,I1092280);
nand I_64094 (I1092305,I1092288,I1092028);
not I_64095 (I1091779,I1092305);
nand I_64096 (I1091773,I1092305,I1092045);
nand I_64097 (I1091770,I1092288,I1091912);
not I_64098 (I1092394,I2690);
DFFARX1 I_64099 (I339922,I2683,I1092394,I1092420,);
DFFARX1 I_64100 (I339928,I2683,I1092394,I1092437,);
not I_64101 (I1092445,I1092437);
nor I_64102 (I1092362,I1092420,I1092445);
DFFARX1 I_64103 (I1092445,I2683,I1092394,I1092377,);
nor I_64104 (I1092490,I339937,I339922);
and I_64105 (I1092507,I1092490,I339949);
nor I_64106 (I1092524,I1092507,I339937);
not I_64107 (I1092541,I339937);
and I_64108 (I1092558,I1092541,I339925);
nand I_64109 (I1092575,I1092558,I339946);
nor I_64110 (I1092592,I1092541,I1092575);
DFFARX1 I_64111 (I1092592,I2683,I1092394,I1092359,);
not I_64112 (I1092623,I1092575);
nand I_64113 (I1092640,I1092445,I1092623);
nand I_64114 (I1092371,I1092507,I1092623);
DFFARX1 I_64115 (I1092541,I2683,I1092394,I1092386,);
not I_64116 (I1092685,I339934);
nor I_64117 (I1092702,I1092685,I339925);
nor I_64118 (I1092719,I1092702,I1092524);
DFFARX1 I_64119 (I1092719,I2683,I1092394,I1092383,);
not I_64120 (I1092750,I1092702);
DFFARX1 I_64121 (I1092750,I2683,I1092394,I1092776,);
not I_64122 (I1092784,I1092776);
nor I_64123 (I1092380,I1092784,I1092702);
nor I_64124 (I1092815,I1092685,I339931);
and I_64125 (I1092832,I1092815,I339943);
or I_64126 (I1092849,I1092832,I339940);
DFFARX1 I_64127 (I1092849,I2683,I1092394,I1092875,);
not I_64128 (I1092883,I1092875);
nand I_64129 (I1092900,I1092883,I1092623);
not I_64130 (I1092374,I1092900);
nand I_64131 (I1092368,I1092900,I1092640);
nand I_64132 (I1092365,I1092883,I1092507);
not I_64133 (I1092989,I2690);
DFFARX1 I_64134 (I330674,I2683,I1092989,I1093015,);
DFFARX1 I_64135 (I330680,I2683,I1092989,I1093032,);
not I_64136 (I1093040,I1093032);
nor I_64137 (I1092957,I1093015,I1093040);
DFFARX1 I_64138 (I1093040,I2683,I1092989,I1092972,);
nor I_64139 (I1093085,I330689,I330674);
and I_64140 (I1093102,I1093085,I330701);
nor I_64141 (I1093119,I1093102,I330689);
not I_64142 (I1093136,I330689);
and I_64143 (I1093153,I1093136,I330677);
nand I_64144 (I1093170,I1093153,I330698);
nor I_64145 (I1093187,I1093136,I1093170);
DFFARX1 I_64146 (I1093187,I2683,I1092989,I1092954,);
not I_64147 (I1093218,I1093170);
nand I_64148 (I1093235,I1093040,I1093218);
nand I_64149 (I1092966,I1093102,I1093218);
DFFARX1 I_64150 (I1093136,I2683,I1092989,I1092981,);
not I_64151 (I1093280,I330686);
nor I_64152 (I1093297,I1093280,I330677);
nor I_64153 (I1093314,I1093297,I1093119);
DFFARX1 I_64154 (I1093314,I2683,I1092989,I1092978,);
not I_64155 (I1093345,I1093297);
DFFARX1 I_64156 (I1093345,I2683,I1092989,I1093371,);
not I_64157 (I1093379,I1093371);
nor I_64158 (I1092975,I1093379,I1093297);
nor I_64159 (I1093410,I1093280,I330683);
and I_64160 (I1093427,I1093410,I330695);
or I_64161 (I1093444,I1093427,I330692);
DFFARX1 I_64162 (I1093444,I2683,I1092989,I1093470,);
not I_64163 (I1093478,I1093470);
nand I_64164 (I1093495,I1093478,I1093218);
not I_64165 (I1092969,I1093495);
nand I_64166 (I1092963,I1093495,I1093235);
nand I_64167 (I1092960,I1093478,I1093102);
not I_64168 (I1093584,I2690);
DFFARX1 I_64169 (I523747,I2683,I1093584,I1093610,);
DFFARX1 I_64170 (I523729,I2683,I1093584,I1093627,);
not I_64171 (I1093635,I1093627);
nor I_64172 (I1093552,I1093610,I1093635);
DFFARX1 I_64173 (I1093635,I2683,I1093584,I1093567,);
nor I_64174 (I1093680,I523735,I523738);
and I_64175 (I1093697,I1093680,I523726);
nor I_64176 (I1093714,I1093697,I523735);
not I_64177 (I1093731,I523735);
and I_64178 (I1093748,I1093731,I523744);
nand I_64179 (I1093765,I1093748,I523732);
nor I_64180 (I1093782,I1093731,I1093765);
DFFARX1 I_64181 (I1093782,I2683,I1093584,I1093549,);
not I_64182 (I1093813,I1093765);
nand I_64183 (I1093830,I1093635,I1093813);
nand I_64184 (I1093561,I1093697,I1093813);
DFFARX1 I_64185 (I1093731,I2683,I1093584,I1093576,);
not I_64186 (I1093875,I523729);
nor I_64187 (I1093892,I1093875,I523744);
nor I_64188 (I1093909,I1093892,I1093714);
DFFARX1 I_64189 (I1093909,I2683,I1093584,I1093573,);
not I_64190 (I1093940,I1093892);
DFFARX1 I_64191 (I1093940,I2683,I1093584,I1093966,);
not I_64192 (I1093974,I1093966);
nor I_64193 (I1093570,I1093974,I1093892);
nor I_64194 (I1094005,I1093875,I523741);
and I_64195 (I1094022,I1094005,I523750);
or I_64196 (I1094039,I1094022,I523726);
DFFARX1 I_64197 (I1094039,I2683,I1093584,I1094065,);
not I_64198 (I1094073,I1094065);
nand I_64199 (I1094090,I1094073,I1093813);
not I_64200 (I1093564,I1094090);
nand I_64201 (I1093558,I1094090,I1093830);
nand I_64202 (I1093555,I1094073,I1093697);
not I_64203 (I1094179,I2690);
DFFARX1 I_64204 (I814744,I2683,I1094179,I1094205,);
DFFARX1 I_64205 (I814735,I2683,I1094179,I1094222,);
not I_64206 (I1094230,I1094222);
nor I_64207 (I1094147,I1094205,I1094230);
DFFARX1 I_64208 (I1094230,I2683,I1094179,I1094162,);
nor I_64209 (I1094275,I814741,I814750);
and I_64210 (I1094292,I1094275,I814753);
nor I_64211 (I1094309,I1094292,I814741);
not I_64212 (I1094326,I814741);
and I_64213 (I1094343,I1094326,I814732);
nand I_64214 (I1094360,I1094343,I814738);
nor I_64215 (I1094377,I1094326,I1094360);
DFFARX1 I_64216 (I1094377,I2683,I1094179,I1094144,);
not I_64217 (I1094408,I1094360);
nand I_64218 (I1094425,I1094230,I1094408);
nand I_64219 (I1094156,I1094292,I1094408);
DFFARX1 I_64220 (I1094326,I2683,I1094179,I1094171,);
not I_64221 (I1094470,I814747);
nor I_64222 (I1094487,I1094470,I814732);
nor I_64223 (I1094504,I1094487,I1094309);
DFFARX1 I_64224 (I1094504,I2683,I1094179,I1094168,);
not I_64225 (I1094535,I1094487);
DFFARX1 I_64226 (I1094535,I2683,I1094179,I1094561,);
not I_64227 (I1094569,I1094561);
nor I_64228 (I1094165,I1094569,I1094487);
nor I_64229 (I1094600,I1094470,I814732);
and I_64230 (I1094617,I1094600,I814735);
or I_64231 (I1094634,I1094617,I814738);
DFFARX1 I_64232 (I1094634,I2683,I1094179,I1094660,);
not I_64233 (I1094668,I1094660);
nand I_64234 (I1094685,I1094668,I1094408);
not I_64235 (I1094159,I1094685);
nand I_64236 (I1094153,I1094685,I1094425);
nand I_64237 (I1094150,I1094668,I1094292);
not I_64238 (I1094774,I2690);
DFFARX1 I_64239 (I899293,I2683,I1094774,I1094800,);
DFFARX1 I_64240 (I899305,I2683,I1094774,I1094817,);
not I_64241 (I1094825,I1094817);
nor I_64242 (I1094742,I1094800,I1094825);
DFFARX1 I_64243 (I1094825,I2683,I1094774,I1094757,);
nor I_64244 (I1094870,I899302,I899296);
and I_64245 (I1094887,I1094870,I899290);
nor I_64246 (I1094904,I1094887,I899302);
not I_64247 (I1094921,I899302);
and I_64248 (I1094938,I1094921,I899299);
nand I_64249 (I1094955,I1094938,I899290);
nor I_64250 (I1094972,I1094921,I1094955);
DFFARX1 I_64251 (I1094972,I2683,I1094774,I1094739,);
not I_64252 (I1095003,I1094955);
nand I_64253 (I1095020,I1094825,I1095003);
nand I_64254 (I1094751,I1094887,I1095003);
DFFARX1 I_64255 (I1094921,I2683,I1094774,I1094766,);
not I_64256 (I1095065,I899314);
nor I_64257 (I1095082,I1095065,I899299);
nor I_64258 (I1095099,I1095082,I1094904);
DFFARX1 I_64259 (I1095099,I2683,I1094774,I1094763,);
not I_64260 (I1095130,I1095082);
DFFARX1 I_64261 (I1095130,I2683,I1094774,I1095156,);
not I_64262 (I1095164,I1095156);
nor I_64263 (I1094760,I1095164,I1095082);
nor I_64264 (I1095195,I1095065,I899308);
and I_64265 (I1095212,I1095195,I899311);
or I_64266 (I1095229,I1095212,I899293);
DFFARX1 I_64267 (I1095229,I2683,I1094774,I1095255,);
not I_64268 (I1095263,I1095255);
nand I_64269 (I1095280,I1095263,I1095003);
not I_64270 (I1094754,I1095280);
nand I_64271 (I1094748,I1095280,I1095020);
nand I_64272 (I1094745,I1095263,I1094887);
not I_64273 (I1095369,I2690);
DFFARX1 I_64274 (I49583,I2683,I1095369,I1095395,);
DFFARX1 I_64275 (I49571,I2683,I1095369,I1095412,);
not I_64276 (I1095420,I1095412);
nor I_64277 (I1095337,I1095395,I1095420);
DFFARX1 I_64278 (I1095420,I2683,I1095369,I1095352,);
nor I_64279 (I1095465,I49562,I49586);
and I_64280 (I1095482,I1095465,I49565);
nor I_64281 (I1095499,I1095482,I49562);
not I_64282 (I1095516,I49562);
and I_64283 (I1095533,I1095516,I49568);
nand I_64284 (I1095550,I1095533,I49580);
nor I_64285 (I1095567,I1095516,I1095550);
DFFARX1 I_64286 (I1095567,I2683,I1095369,I1095334,);
not I_64287 (I1095598,I1095550);
nand I_64288 (I1095615,I1095420,I1095598);
nand I_64289 (I1095346,I1095482,I1095598);
DFFARX1 I_64290 (I1095516,I2683,I1095369,I1095361,);
not I_64291 (I1095660,I49562);
nor I_64292 (I1095677,I1095660,I49568);
nor I_64293 (I1095694,I1095677,I1095499);
DFFARX1 I_64294 (I1095694,I2683,I1095369,I1095358,);
not I_64295 (I1095725,I1095677);
DFFARX1 I_64296 (I1095725,I2683,I1095369,I1095751,);
not I_64297 (I1095759,I1095751);
nor I_64298 (I1095355,I1095759,I1095677);
nor I_64299 (I1095790,I1095660,I49565);
and I_64300 (I1095807,I1095790,I49574);
or I_64301 (I1095824,I1095807,I49577);
DFFARX1 I_64302 (I1095824,I2683,I1095369,I1095850,);
not I_64303 (I1095858,I1095850);
nand I_64304 (I1095875,I1095858,I1095598);
not I_64305 (I1095349,I1095875);
nand I_64306 (I1095343,I1095875,I1095615);
nand I_64307 (I1095340,I1095858,I1095482);
not I_64308 (I1095964,I2690);
DFFARX1 I_64309 (I793641,I2683,I1095964,I1095990,);
DFFARX1 I_64310 (I793659,I2683,I1095964,I1096007,);
not I_64311 (I1096015,I1096007);
nor I_64312 (I1095932,I1095990,I1096015);
DFFARX1 I_64313 (I1096015,I2683,I1095964,I1095947,);
nor I_64314 (I1096060,I793638,I793650);
and I_64315 (I1096077,I1096060,I793635);
nor I_64316 (I1096094,I1096077,I793638);
not I_64317 (I1096111,I793638);
and I_64318 (I1096128,I1096111,I793644);
nand I_64319 (I1096145,I1096128,I793656);
nor I_64320 (I1096162,I1096111,I1096145);
DFFARX1 I_64321 (I1096162,I2683,I1095964,I1095929,);
not I_64322 (I1096193,I1096145);
nand I_64323 (I1096210,I1096015,I1096193);
nand I_64324 (I1095941,I1096077,I1096193);
DFFARX1 I_64325 (I1096111,I2683,I1095964,I1095956,);
not I_64326 (I1096255,I793647);
nor I_64327 (I1096272,I1096255,I793644);
nor I_64328 (I1096289,I1096272,I1096094);
DFFARX1 I_64329 (I1096289,I2683,I1095964,I1095953,);
not I_64330 (I1096320,I1096272);
DFFARX1 I_64331 (I1096320,I2683,I1095964,I1096346,);
not I_64332 (I1096354,I1096346);
nor I_64333 (I1095950,I1096354,I1096272);
nor I_64334 (I1096385,I1096255,I793635);
and I_64335 (I1096402,I1096385,I793662);
or I_64336 (I1096419,I1096402,I793653);
DFFARX1 I_64337 (I1096419,I2683,I1095964,I1096445,);
not I_64338 (I1096453,I1096445);
nand I_64339 (I1096470,I1096453,I1096193);
not I_64340 (I1095944,I1096470);
nand I_64341 (I1095938,I1096470,I1096210);
nand I_64342 (I1095935,I1096453,I1096077);
not I_64343 (I1096559,I2690);
DFFARX1 I_64344 (I553803,I2683,I1096559,I1096585,);
DFFARX1 I_64345 (I553785,I2683,I1096559,I1096602,);
not I_64346 (I1096610,I1096602);
nor I_64347 (I1096527,I1096585,I1096610);
DFFARX1 I_64348 (I1096610,I2683,I1096559,I1096542,);
nor I_64349 (I1096655,I553791,I553794);
and I_64350 (I1096672,I1096655,I553782);
nor I_64351 (I1096689,I1096672,I553791);
not I_64352 (I1096706,I553791);
and I_64353 (I1096723,I1096706,I553800);
nand I_64354 (I1096740,I1096723,I553788);
nor I_64355 (I1096757,I1096706,I1096740);
DFFARX1 I_64356 (I1096757,I2683,I1096559,I1096524,);
not I_64357 (I1096788,I1096740);
nand I_64358 (I1096805,I1096610,I1096788);
nand I_64359 (I1096536,I1096672,I1096788);
DFFARX1 I_64360 (I1096706,I2683,I1096559,I1096551,);
not I_64361 (I1096850,I553785);
nor I_64362 (I1096867,I1096850,I553800);
nor I_64363 (I1096884,I1096867,I1096689);
DFFARX1 I_64364 (I1096884,I2683,I1096559,I1096548,);
not I_64365 (I1096915,I1096867);
DFFARX1 I_64366 (I1096915,I2683,I1096559,I1096941,);
not I_64367 (I1096949,I1096941);
nor I_64368 (I1096545,I1096949,I1096867);
nor I_64369 (I1096980,I1096850,I553797);
and I_64370 (I1096997,I1096980,I553806);
or I_64371 (I1097014,I1096997,I553782);
DFFARX1 I_64372 (I1097014,I2683,I1096559,I1097040,);
not I_64373 (I1097048,I1097040);
nand I_64374 (I1097065,I1097048,I1096788);
not I_64375 (I1096539,I1097065);
nand I_64376 (I1096533,I1097065,I1096805);
nand I_64377 (I1096530,I1097048,I1096672);
not I_64378 (I1097154,I2690);
DFFARX1 I_64379 (I647563,I2683,I1097154,I1097180,);
DFFARX1 I_64380 (I647560,I2683,I1097154,I1097197,);
not I_64381 (I1097205,I1097197);
nor I_64382 (I1097122,I1097180,I1097205);
DFFARX1 I_64383 (I1097205,I2683,I1097154,I1097137,);
nor I_64384 (I1097250,I647575,I647557);
and I_64385 (I1097267,I1097250,I647554);
nor I_64386 (I1097284,I1097267,I647575);
not I_64387 (I1097301,I647575);
and I_64388 (I1097318,I1097301,I647560);
nand I_64389 (I1097335,I1097318,I647572);
nor I_64390 (I1097352,I1097301,I1097335);
DFFARX1 I_64391 (I1097352,I2683,I1097154,I1097119,);
not I_64392 (I1097383,I1097335);
nand I_64393 (I1097400,I1097205,I1097383);
nand I_64394 (I1097131,I1097267,I1097383);
DFFARX1 I_64395 (I1097301,I2683,I1097154,I1097146,);
not I_64396 (I1097445,I647566);
nor I_64397 (I1097462,I1097445,I647560);
nor I_64398 (I1097479,I1097462,I1097284);
DFFARX1 I_64399 (I1097479,I2683,I1097154,I1097143,);
not I_64400 (I1097510,I1097462);
DFFARX1 I_64401 (I1097510,I2683,I1097154,I1097536,);
not I_64402 (I1097544,I1097536);
nor I_64403 (I1097140,I1097544,I1097462);
nor I_64404 (I1097575,I1097445,I647554);
and I_64405 (I1097592,I1097575,I647569);
or I_64406 (I1097609,I1097592,I647557);
DFFARX1 I_64407 (I1097609,I2683,I1097154,I1097635,);
not I_64408 (I1097643,I1097635);
nand I_64409 (I1097660,I1097643,I1097383);
not I_64410 (I1097134,I1097660);
nand I_64411 (I1097128,I1097660,I1097400);
nand I_64412 (I1097125,I1097643,I1097267);
not I_64413 (I1097749,I2690);
DFFARX1 I_64414 (I368210,I2683,I1097749,I1097775,);
DFFARX1 I_64415 (I368216,I2683,I1097749,I1097792,);
not I_64416 (I1097800,I1097792);
nor I_64417 (I1097717,I1097775,I1097800);
DFFARX1 I_64418 (I1097800,I2683,I1097749,I1097732,);
nor I_64419 (I1097845,I368225,I368210);
and I_64420 (I1097862,I1097845,I368237);
nor I_64421 (I1097879,I1097862,I368225);
not I_64422 (I1097896,I368225);
and I_64423 (I1097913,I1097896,I368213);
nand I_64424 (I1097930,I1097913,I368234);
nor I_64425 (I1097947,I1097896,I1097930);
DFFARX1 I_64426 (I1097947,I2683,I1097749,I1097714,);
not I_64427 (I1097978,I1097930);
nand I_64428 (I1097995,I1097800,I1097978);
nand I_64429 (I1097726,I1097862,I1097978);
DFFARX1 I_64430 (I1097896,I2683,I1097749,I1097741,);
not I_64431 (I1098040,I368222);
nor I_64432 (I1098057,I1098040,I368213);
nor I_64433 (I1098074,I1098057,I1097879);
DFFARX1 I_64434 (I1098074,I2683,I1097749,I1097738,);
not I_64435 (I1098105,I1098057);
DFFARX1 I_64436 (I1098105,I2683,I1097749,I1098131,);
not I_64437 (I1098139,I1098131);
nor I_64438 (I1097735,I1098139,I1098057);
nor I_64439 (I1098170,I1098040,I368219);
and I_64440 (I1098187,I1098170,I368231);
or I_64441 (I1098204,I1098187,I368228);
DFFARX1 I_64442 (I1098204,I2683,I1097749,I1098230,);
not I_64443 (I1098238,I1098230);
nand I_64444 (I1098255,I1098238,I1097978);
not I_64445 (I1097729,I1098255);
nand I_64446 (I1097723,I1098255,I1097995);
nand I_64447 (I1097720,I1098238,I1097862);
not I_64448 (I1098344,I2690);
DFFARX1 I_64449 (I426452,I2683,I1098344,I1098370,);
DFFARX1 I_64450 (I426455,I2683,I1098344,I1098387,);
not I_64451 (I1098395,I1098387);
nor I_64452 (I1098312,I1098370,I1098395);
DFFARX1 I_64453 (I1098395,I2683,I1098344,I1098327,);
nor I_64454 (I1098440,I426458,I426476);
and I_64455 (I1098457,I1098440,I426461);
nor I_64456 (I1098474,I1098457,I426458);
not I_64457 (I1098491,I426458);
and I_64458 (I1098508,I1098491,I426470);
nand I_64459 (I1098525,I1098508,I426473);
nor I_64460 (I1098542,I1098491,I1098525);
DFFARX1 I_64461 (I1098542,I2683,I1098344,I1098309,);
not I_64462 (I1098573,I1098525);
nand I_64463 (I1098590,I1098395,I1098573);
nand I_64464 (I1098321,I1098457,I1098573);
DFFARX1 I_64465 (I1098491,I2683,I1098344,I1098336,);
not I_64466 (I1098635,I426464);
nor I_64467 (I1098652,I1098635,I426470);
nor I_64468 (I1098669,I1098652,I1098474);
DFFARX1 I_64469 (I1098669,I2683,I1098344,I1098333,);
not I_64470 (I1098700,I1098652);
DFFARX1 I_64471 (I1098700,I2683,I1098344,I1098726,);
not I_64472 (I1098734,I1098726);
nor I_64473 (I1098330,I1098734,I1098652);
nor I_64474 (I1098765,I1098635,I426452);
and I_64475 (I1098782,I1098765,I426467);
or I_64476 (I1098799,I1098782,I426455);
DFFARX1 I_64477 (I1098799,I2683,I1098344,I1098825,);
not I_64478 (I1098833,I1098825);
nand I_64479 (I1098850,I1098833,I1098573);
not I_64480 (I1098324,I1098850);
nand I_64481 (I1098318,I1098850,I1098590);
nand I_64482 (I1098315,I1098833,I1098457);
not I_64483 (I1098939,I2690);
DFFARX1 I_64484 (I97540,I2683,I1098939,I1098965,);
DFFARX1 I_64485 (I97528,I2683,I1098939,I1098982,);
not I_64486 (I1098990,I1098982);
nor I_64487 (I1098907,I1098965,I1098990);
DFFARX1 I_64488 (I1098990,I2683,I1098939,I1098922,);
nor I_64489 (I1099035,I97519,I97543);
and I_64490 (I1099052,I1099035,I97522);
nor I_64491 (I1099069,I1099052,I97519);
not I_64492 (I1099086,I97519);
and I_64493 (I1099103,I1099086,I97525);
nand I_64494 (I1099120,I1099103,I97537);
nor I_64495 (I1099137,I1099086,I1099120);
DFFARX1 I_64496 (I1099137,I2683,I1098939,I1098904,);
not I_64497 (I1099168,I1099120);
nand I_64498 (I1099185,I1098990,I1099168);
nand I_64499 (I1098916,I1099052,I1099168);
DFFARX1 I_64500 (I1099086,I2683,I1098939,I1098931,);
not I_64501 (I1099230,I97519);
nor I_64502 (I1099247,I1099230,I97525);
nor I_64503 (I1099264,I1099247,I1099069);
DFFARX1 I_64504 (I1099264,I2683,I1098939,I1098928,);
not I_64505 (I1099295,I1099247);
DFFARX1 I_64506 (I1099295,I2683,I1098939,I1099321,);
not I_64507 (I1099329,I1099321);
nor I_64508 (I1098925,I1099329,I1099247);
nor I_64509 (I1099360,I1099230,I97522);
and I_64510 (I1099377,I1099360,I97531);
or I_64511 (I1099394,I1099377,I97534);
DFFARX1 I_64512 (I1099394,I2683,I1098939,I1099420,);
not I_64513 (I1099428,I1099420);
nand I_64514 (I1099445,I1099428,I1099168);
not I_64515 (I1098919,I1099445);
nand I_64516 (I1098913,I1099445,I1099185);
nand I_64517 (I1098910,I1099428,I1099052);
not I_64518 (I1099534,I2690);
DFFARX1 I_64519 (I681818,I2683,I1099534,I1099560,);
DFFARX1 I_64520 (I681815,I2683,I1099534,I1099577,);
not I_64521 (I1099585,I1099577);
nor I_64522 (I1099502,I1099560,I1099585);
DFFARX1 I_64523 (I1099585,I2683,I1099534,I1099517,);
nor I_64524 (I1099630,I681830,I681812);
and I_64525 (I1099647,I1099630,I681809);
nor I_64526 (I1099664,I1099647,I681830);
not I_64527 (I1099681,I681830);
and I_64528 (I1099698,I1099681,I681815);
nand I_64529 (I1099715,I1099698,I681827);
nor I_64530 (I1099732,I1099681,I1099715);
DFFARX1 I_64531 (I1099732,I2683,I1099534,I1099499,);
not I_64532 (I1099763,I1099715);
nand I_64533 (I1099780,I1099585,I1099763);
nand I_64534 (I1099511,I1099647,I1099763);
DFFARX1 I_64535 (I1099681,I2683,I1099534,I1099526,);
not I_64536 (I1099825,I681821);
nor I_64537 (I1099842,I1099825,I681815);
nor I_64538 (I1099859,I1099842,I1099664);
DFFARX1 I_64539 (I1099859,I2683,I1099534,I1099523,);
not I_64540 (I1099890,I1099842);
DFFARX1 I_64541 (I1099890,I2683,I1099534,I1099916,);
not I_64542 (I1099924,I1099916);
nor I_64543 (I1099520,I1099924,I1099842);
nor I_64544 (I1099955,I1099825,I681809);
and I_64545 (I1099972,I1099955,I681824);
or I_64546 (I1099989,I1099972,I681812);
DFFARX1 I_64547 (I1099989,I2683,I1099534,I1100015,);
not I_64548 (I1100023,I1100015);
nand I_64549 (I1100040,I1100023,I1099763);
not I_64550 (I1099514,I1100040);
nand I_64551 (I1099508,I1100040,I1099780);
nand I_64552 (I1099505,I1100023,I1099647);
not I_64553 (I1100129,I2690);
DFFARX1 I_64554 (I97013,I2683,I1100129,I1100155,);
DFFARX1 I_64555 (I97001,I2683,I1100129,I1100172,);
not I_64556 (I1100180,I1100172);
nor I_64557 (I1100097,I1100155,I1100180);
DFFARX1 I_64558 (I1100180,I2683,I1100129,I1100112,);
nor I_64559 (I1100225,I96992,I97016);
and I_64560 (I1100242,I1100225,I96995);
nor I_64561 (I1100259,I1100242,I96992);
not I_64562 (I1100276,I96992);
and I_64563 (I1100293,I1100276,I96998);
nand I_64564 (I1100310,I1100293,I97010);
nor I_64565 (I1100327,I1100276,I1100310);
DFFARX1 I_64566 (I1100327,I2683,I1100129,I1100094,);
not I_64567 (I1100358,I1100310);
nand I_64568 (I1100375,I1100180,I1100358);
nand I_64569 (I1100106,I1100242,I1100358);
DFFARX1 I_64570 (I1100276,I2683,I1100129,I1100121,);
not I_64571 (I1100420,I96992);
nor I_64572 (I1100437,I1100420,I96998);
nor I_64573 (I1100454,I1100437,I1100259);
DFFARX1 I_64574 (I1100454,I2683,I1100129,I1100118,);
not I_64575 (I1100485,I1100437);
DFFARX1 I_64576 (I1100485,I2683,I1100129,I1100511,);
not I_64577 (I1100519,I1100511);
nor I_64578 (I1100115,I1100519,I1100437);
nor I_64579 (I1100550,I1100420,I96995);
and I_64580 (I1100567,I1100550,I97004);
or I_64581 (I1100584,I1100567,I97007);
DFFARX1 I_64582 (I1100584,I2683,I1100129,I1100610,);
not I_64583 (I1100618,I1100610);
nand I_64584 (I1100635,I1100618,I1100358);
not I_64585 (I1100109,I1100635);
nand I_64586 (I1100103,I1100635,I1100375);
nand I_64587 (I1100100,I1100618,I1100242);
not I_64588 (I1100724,I2690);
DFFARX1 I_64589 (I1018648,I2683,I1100724,I1100750,);
DFFARX1 I_64590 (I1018639,I2683,I1100724,I1100767,);
not I_64591 (I1100775,I1100767);
nor I_64592 (I1100692,I1100750,I1100775);
DFFARX1 I_64593 (I1100775,I2683,I1100724,I1100707,);
nor I_64594 (I1100820,I1018630,I1018645);
and I_64595 (I1100837,I1100820,I1018633);
nor I_64596 (I1100854,I1100837,I1018630);
not I_64597 (I1100871,I1018630);
and I_64598 (I1100888,I1100871,I1018636);
nand I_64599 (I1100905,I1100888,I1018654);
nor I_64600 (I1100922,I1100871,I1100905);
DFFARX1 I_64601 (I1100922,I2683,I1100724,I1100689,);
not I_64602 (I1100953,I1100905);
nand I_64603 (I1100970,I1100775,I1100953);
nand I_64604 (I1100701,I1100837,I1100953);
DFFARX1 I_64605 (I1100871,I2683,I1100724,I1100716,);
not I_64606 (I1101015,I1018630);
nor I_64607 (I1101032,I1101015,I1018636);
nor I_64608 (I1101049,I1101032,I1100854);
DFFARX1 I_64609 (I1101049,I2683,I1100724,I1100713,);
not I_64610 (I1101080,I1101032);
DFFARX1 I_64611 (I1101080,I2683,I1100724,I1101106,);
not I_64612 (I1101114,I1101106);
nor I_64613 (I1100710,I1101114,I1101032);
nor I_64614 (I1101145,I1101015,I1018633);
and I_64615 (I1101162,I1101145,I1018642);
or I_64616 (I1101179,I1101162,I1018651);
DFFARX1 I_64617 (I1101179,I2683,I1100724,I1101205,);
not I_64618 (I1101213,I1101205);
nand I_64619 (I1101230,I1101213,I1100953);
not I_64620 (I1100704,I1101230);
nand I_64621 (I1100698,I1101230,I1100970);
nand I_64622 (I1100695,I1101213,I1100837);
not I_64623 (I1101319,I2690);
DFFARX1 I_64624 (I356242,I2683,I1101319,I1101345,);
DFFARX1 I_64625 (I356248,I2683,I1101319,I1101362,);
not I_64626 (I1101370,I1101362);
nor I_64627 (I1101287,I1101345,I1101370);
DFFARX1 I_64628 (I1101370,I2683,I1101319,I1101302,);
nor I_64629 (I1101415,I356257,I356242);
and I_64630 (I1101432,I1101415,I356269);
nor I_64631 (I1101449,I1101432,I356257);
not I_64632 (I1101466,I356257);
and I_64633 (I1101483,I1101466,I356245);
nand I_64634 (I1101500,I1101483,I356266);
nor I_64635 (I1101517,I1101466,I1101500);
DFFARX1 I_64636 (I1101517,I2683,I1101319,I1101284,);
not I_64637 (I1101548,I1101500);
nand I_64638 (I1101565,I1101370,I1101548);
nand I_64639 (I1101296,I1101432,I1101548);
DFFARX1 I_64640 (I1101466,I2683,I1101319,I1101311,);
not I_64641 (I1101610,I356254);
nor I_64642 (I1101627,I1101610,I356245);
nor I_64643 (I1101644,I1101627,I1101449);
DFFARX1 I_64644 (I1101644,I2683,I1101319,I1101308,);
not I_64645 (I1101675,I1101627);
DFFARX1 I_64646 (I1101675,I2683,I1101319,I1101701,);
not I_64647 (I1101709,I1101701);
nor I_64648 (I1101305,I1101709,I1101627);
nor I_64649 (I1101740,I1101610,I356251);
and I_64650 (I1101757,I1101740,I356263);
or I_64651 (I1101774,I1101757,I356260);
DFFARX1 I_64652 (I1101774,I2683,I1101319,I1101800,);
not I_64653 (I1101808,I1101800);
nand I_64654 (I1101825,I1101808,I1101548);
not I_64655 (I1101299,I1101825);
nand I_64656 (I1101293,I1101825,I1101565);
nand I_64657 (I1101290,I1101808,I1101432);
endmodule


