module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_5_r_15,n9_15,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
and I_44(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_45(N1508_0_r_15,n55_15,N1508_0_r_10);
nor I_46(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_47(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_48(N1372_4_r_15,n39_15);
nor I_49(N1508_4_r_15,n39_15,n43_15);
nand I_50(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_51(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_52(n_576_5_r_15,n31_15,n32_15);
not I_53(n_102_5_r_15,n33_15);
nand I_54(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_55(N1507_6_r_15,n42_15,n46_15);
nand I_56(N1508_6_r_15,n39_15,n40_15);
nand I_57(n_431_5_r_15,n36_15,n37_15);
not I_58(n9_15,blif_reset_net_5_r_15);
nor I_59(n31_15,n33_15,n34_15);
nor I_60(n32_15,n44_15,N6147_2_r_10);
nor I_61(n33_15,n54_15,n55_15);
nand I_62(n34_15,n49_15,N1508_4_r_10);
nand I_63(n35_15,N1507_6_r_10,N6147_3_r_10);
not I_64(n36_15,n32_15);
nand I_65(n37_15,n34_15,n38_15);
not I_66(n38_15,n46_15);
nand I_67(n39_15,n38_15,n41_15);
nand I_68(n40_15,n41_15,n42_15);
and I_69(n41_15,n51_15,N1371_0_r_10);
and I_70(n42_15,n47_15,N6147_3_r_10);
and I_71(n43_15,n34_15,n36_15);
or I_72(n44_15,G199_8_r_10,N6147_9_r_10);
not I_73(n45_15,N1372_1_r_15);
nand I_74(n46_15,n53_15,N6147_3_r_10);
nor I_75(n47_15,n34_15,n48_15);
not I_76(n48_15,N1507_6_r_10);
and I_77(n49_15,n50_15,N1508_0_r_10);
nand I_78(n50_15,n51_15,n52_15);
nand I_79(n51_15,N6147_3_r_10,N6147_2_r_10);
not I_80(n52_15,N1371_0_r_10);
nor I_81(n53_15,n48_15,N6134_9_r_10);
nor I_82(n54_15,n_42_8_r_10,N1371_0_r_10);
not I_83(n55_15,N1508_6_r_10);
endmodule


