module test_I15228(I12930,I1477,I12653,I15160,I1470,I15228);
input I12930,I1477,I12653,I15160,I1470;
output I15228;
wire I12670,I12783,I15064,I12596,I14965,I13023,I12608,I15194,I12593,I12587,I12619,I15047,I14982,I15177,I15211,I12584;
DFFARX1 I_0(I12653,I1470,I12619,,,I12670,);
DFFARX1 I_1(I1470,I12619,,,I12783,);
nand I_2(I15064,I15047,I12587);
DFFARX1 I_3(I1470,I12619,,,I12596,);
not I_4(I14965,I1477);
DFFARX1 I_5(I1470,I12619,,,I13023,);
nor I_6(I12608,I13023,I12930);
or I_7(I15194,I15177,I12608);
nand I_8(I12593,I12670);
DFFARX1 I_9(I12670,I1470,I12619,,,I12587,);
not I_10(I12619,I1477);
nor I_11(I15047,I14982,I12584);
not I_12(I14982,I12596);
and I_13(I15177,I15160,I12593);
DFFARX1 I_14(I15194,I1470,I14965,,,I15211,);
nor I_15(I15228,I15211,I15064);
and I_16(I12584,I12670,I12783);
endmodule


