module test_I1518_rst(I1477_rst,I1518_rst);
,I1518_rst);
input I1477_rst;
output I1518_rst;
wire ;
not I_0(I1518_rst,I1477_rst);
endmodule


