module test_I7221(I5416,I1477,I5546,I1470,I7221);
input I5416,I1477,I5546,I1470;
output I7221;
wire I5659,I5450,I5073,I5625,I5088,I5433,I5563,I5512,I5105,I5642,I6924;
or I_0(I5659,I5642,I5563);
and I_1(I5450,I5416,I5433);
DFFARX1 I_2(I5450,I1470,I5105,,,I5073,);
DFFARX1 I_3(I1470,I5105,,,I5625,);
DFFARX1 I_4(I5659,I1470,I5105,,,I5088,);
nand I_5(I5433,I5416);
and I_6(I5563,I5512,I5546);
DFFARX1 I_7(I1470,I5105,,,I5512,);
nand I_8(I7221,I6924,I5088);
not I_9(I5105,I1477);
not I_10(I5642,I5625);
not I_11(I6924,I5073);
endmodule


