module test_I15576(I13761,I1477,I1470,I15863,I15576);
input I13761,I1477,I1470,I15863;
output I15576;
wire I15897,I14083,I15713,I13746,I15880,I15815,I15611,I15928,I16007;
and I_0(I15897,I15713,I15880);
DFFARX1 I_1(I1470,,,I14083,);
not I_2(I15713,I13761);
DFFARX1 I_3(I16007,I1470,I15611,,,I15576,);
not I_4(I13746,I14083);
nor I_5(I15880,I15815,I15863);
DFFARX1 I_6(I1470,I15611,,,I15815,);
not I_7(I15611,I1477);
DFFARX1 I_8(I13746,I1470,I15611,,,I15928,);
or I_9(I16007,I15928,I15897);
endmodule


