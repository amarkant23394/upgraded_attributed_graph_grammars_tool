module test_I6975(I1477,I3521,I1470,I3846,I5122,I6975);
input I1477,I3521,I1470,I3846,I5122;
output I6975;
wire I5416,I5450,I5073,I5070,I3380,I5433,I5481,I5249,I3356,I5105,I6924;
nand I_0(I5416,I5122,I3356);
and I_1(I5450,I5416,I5433);
DFFARX1 I_2(I5450,I1470,I5105,,,I5073,);
nor I_3(I6975,I6924,I5070);
and I_4(I5070,I5249,I5481);
nand I_5(I3380,I3521,I3846);
nand I_6(I5433,I5416);
DFFARX1 I_7(I5416,I1470,I5105,,,I5481,);
not I_8(I5249,I3380);
DFFARX1 I_9(I1470,,,I3356,);
not I_10(I5105,I1477);
not I_11(I6924,I5073);
endmodule


