module test_I17727(I15713,I15645,I1477,I13746,I15880,I1470,I13764,I17727);
input I15713,I15645,I1477,I13746,I15880,I1470,I13764;
output I17727;
wire I15897,I17430,I15730,I15576,I15662,I15579,I15611,I15976,I15928,I16007;
and I_0(I15897,I15713,I15880);
not I_1(I17430,I15579);
not I_2(I15730,I15713);
DFFARX1 I_3(I16007,I1470,I15611,,,I15576,);
nand I_4(I15662,I15645,I13764);
nand I_5(I15579,I15662,I15976);
not I_6(I15611,I1477);
nor I_7(I15976,I15928,I15730);
nand I_8(I17727,I17430,I15576);
DFFARX1 I_9(I13746,I1470,I15611,,,I15928,);
or I_10(I16007,I15928,I15897);
endmodule


