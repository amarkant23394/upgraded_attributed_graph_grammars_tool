module test_I9303(I5659,I1477,I1470,I9303);
input I5659,I1477,I1470;
output I9303;
wire I6875,I5073,I5088,I8862,I6907,I7221,I5105,I6924;
DFFARX1 I_0(I7221,I1470,I6907,,,I6875,);
DFFARX1 I_1(I1470,I5105,,,I5073,);
DFFARX1 I_2(I5659,I1470,I5105,,,I5088,);
DFFARX1 I_3(I6875,I1470,I8862,,,I9303,);
not I_4(I8862,I1477);
not I_5(I6907,I1477);
nand I_6(I7221,I6924,I5088);
not I_7(I5105,I1477);
not I_8(I6924,I5073);
endmodule


