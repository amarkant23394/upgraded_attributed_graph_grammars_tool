module test_I2143(I1303,I1477,I1247,I1470,I2143);
input I1303,I1477,I1247,I1470;
output I2143;
wire I2540,I2181,I2557;
DFFARX1 I_0(I1247,I1470,I2181,,,I2540,);
DFFARX1 I_1(I2557,I1470,I2181,,,I2143,);
not I_2(I2181,I1477);
and I_3(I2557,I2540,I1303);
endmodule


