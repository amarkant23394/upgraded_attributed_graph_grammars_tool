module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_7_r_16,n8_16,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
nor I_41(N1371_0_r_16,n35_16,n39_16);
nor I_42(N1508_0_r_16,n39_16,n46_16);
not I_43(N1372_1_r_16,n45_16);
nor I_44(N1508_1_r_16,n53_16,n45_16);
nor I_45(N6147_2_r_16,n37_16,n38_16);
nor I_46(N1507_6_r_16,n44_16,n49_16);
nor I_47(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_48(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_49(n_572_7_r_16,n32_16,n33_16);
nand I_50(n_573_7_r_16,n30_16,n31_16);
nand I_51(n_549_7_r_16,n47_16,N1508_0_r_1);
nand I_52(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_53(n_452_7_r_16,n34_16,n35_16);
and I_54(N3_8_l_16,n41_16,N1507_6_r_1);
not I_55(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_56(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_57(n29_16,n53_16);
nor I_58(n4_7_r_16,n35_16,n36_16);
nand I_59(n30_16,n_569_7_r_1,N6147_9_r_1);
not I_60(n31_16,n34_16);
nor I_61(n32_16,n30_16,N1507_6_r_1);
not I_62(n33_16,n_549_7_r_16);
nor I_63(n34_16,n48_16,n_549_7_r_1);
and I_64(n35_16,n50_16,G42_7_r_1);
not I_65(n36_16,n30_16);
nor I_66(n37_16,n31_16,n40_16);
nand I_67(n38_16,n29_16,n39_16);
not I_68(n39_16,n32_16);
nor I_69(n40_16,N1508_6_r_1,G42_7_r_1);
nand I_70(n41_16,N1508_0_r_1,G42_7_r_1);
nand I_71(n42_16,n35_16,n43_16);
not I_72(n43_16,n44_16);
nor I_73(n44_16,n32_16,n49_16);
nand I_74(n45_16,n36_16,n40_16);
nor I_75(n46_16,n33_16,n34_16);
nand I_76(n47_16,n_572_7_r_1,N6134_9_r_1);
or I_77(n48_16,N1508_6_r_1,n_572_7_r_1);
and I_78(n49_16,n35_16,n36_16);
and I_79(n50_16,n51_16,n_573_7_r_1);
nand I_80(n51_16,n47_16,n52_16);
not I_81(n52_16,N1508_0_r_1);
endmodule


