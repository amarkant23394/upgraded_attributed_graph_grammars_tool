module Benchmark_testing100(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294_clk,I1301_rst,I3235,I3220,I3217,I3214,I3232,I3229,I3208,I3211,I3238,I3223,I3226);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294_clk,I1301_rst;
output I3235,I3220,I3217,I3214,I3232,I3229,I3208,I3211,I3238,I3223,I3226;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294_clk,I1301_rst,I1342_rst,I1359,I1376,I1393,I1313,I1424,I1441,I1458,I1475,I1492,I1509,I1526,I1543,I1560,I1577,I1328,I1325,I1622,I1310,I1653,I1307,I1684,I1701,I1718,I1735,I1752,I1769,I1334,I1800,I1322,I1316,I1845,I1862,I1331,I1893,I1910,I1927,I1319,I1304,I2005_rst,I2022,I2039,I2056,I2073,I2090,I2107,I1976,I2138,I2155,I2172,I2189,I2206,I2223,I2240,I1973,I1967,I2285,I2302,I2319,I1994,I2350,I2367,I1985,I1979,I2412,I1982,I2443,I2460,I1997,I2491,I1991,I1988,I2536,I1970,I2600_rst,I2617,I2634,I2651,I2574,I2682,I2699,I2589,I2571,I2744,I2761,I2778,I2795,I2812,I2829,I2846,I2863,I2880,I2586,I2911,I2928,I2945,I2568,I2976,I2565,I3007,I3024,I3041,I3058,I2580,I3089,I2577,I3120,I3137,I3154,I2583,I2592,I2562,I3246_rst,I3263,I3280,I3297,I3314,I3331,I3348,I3365,I3396,I3427,I3444,I3461,I3478,I3495,I3512,I3529,I3560,I3577,I3608,I3625,I3656,I3687,I3704,I3749,I3766,I3783,I3800,I3831;
not I_0 (I1342_rst,I1301_rst);
not I_1 (I1359,I1263);
nor I_2 (I1376,I1215,I1223);
nand I_3 (I1393,I1376,I1287);
DFFARX1 I_4  ( .D(I1393), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1313) );
nor I_5 (I1424,I1359,I1215);
nand I_6 (I1441,I1424,I1247);
nand I_7 (I1458,I1441,I1393);
not I_8 (I1475,I1215);
not I_9 (I1492,I1207);
nor I_10 (I1509,I1492,I1231);
and I_11 (I1526,I1509,I1271);
or I_12 (I1543,I1526,I1255);
DFFARX1 I_13  ( .D(I1543), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1560) );
nor I_14 (I1577,I1560,I1441);
nand I_15 (I1328,I1475,I1577);
not I_16 (I1325,I1560);
and I_17 (I1622,I1560,I1458);
DFFARX1 I_18  ( .D(I1622), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1310) );
DFFARX1 I_19  ( .D(I1560), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1653) );
and I_20 (I1307,I1475,I1653);
nand I_21 (I1684,I1359,I1207);
not I_22 (I1701,I1684);
nor I_23 (I1718,I1560,I1701);
DFFARX1 I_24  ( .D(I1239), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1735) );
nand I_25 (I1752,I1735,I1684);
and I_26 (I1769,I1475,I1752);
DFFARX1 I_27  ( .D(I1769), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1334) );
not I_28 (I1800,I1735);
nand I_29 (I1322,I1735,I1718);
nand I_30 (I1316,I1735,I1701);
DFFARX1 I_31  ( .D(I1279), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1845) );
not I_32 (I1862,I1845);
nor I_33 (I1331,I1735,I1862);
nor I_34 (I1893,I1862,I1800);
and I_35 (I1910,I1441,I1893);
or I_36 (I1927,I1684,I1910);
DFFARX1 I_37  ( .D(I1927), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1319) );
DFFARX1 I_38  ( .D(I1862), .CLK(I1294_clk), .RSTB(I1342_rst), .Q(I1304) );
not I_39 (I2005_rst,I1301_rst);
nand I_40 (I2022,I1307,I1328);
and I_41 (I2039,I2022,I1313);
DFFARX1 I_42  ( .D(I2039), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I2056) );
nor I_43 (I2073,I1331,I1328);
DFFARX1 I_44  ( .D(I1334), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I2090) );
nand I_45 (I2107,I2090,I2073);
DFFARX1 I_46  ( .D(I2090), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I1976) );
nand I_47 (I2138,I1304,I1316);
and I_48 (I2155,I2138,I1325);
DFFARX1 I_49  ( .D(I2155), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I2172) );
not I_50 (I2189,I2172);
nor I_51 (I2206,I2056,I2189);
and I_52 (I2223,I2073,I2206);
and I_53 (I2240,I2172,I2107);
DFFARX1 I_54  ( .D(I2240), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I1973) );
DFFARX1 I_55  ( .D(I2172), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I1967) );
DFFARX1 I_56  ( .D(I1319), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I2285) );
and I_57 (I2302,I2285,I1322);
nand I_58 (I2319,I2302,I2172);
nor I_59 (I1994,I2302,I2073);
not I_60 (I2350,I2302);
nor I_61 (I2367,I2056,I2350);
nand I_62 (I1985,I2090,I2367);
nand I_63 (I1979,I2172,I2350);
or I_64 (I2412,I2302,I2223);
DFFARX1 I_65  ( .D(I2412), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I1982) );
DFFARX1 I_66  ( .D(I1310), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I2443) );
and I_67 (I2460,I2443,I2319);
DFFARX1 I_68  ( .D(I2460), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I1997) );
nor I_69 (I2491,I2443,I2056);
nand I_70 (I1991,I2302,I2491);
not I_71 (I1988,I2443);
DFFARX1 I_72  ( .D(I2443), .CLK(I1294_clk), .RSTB(I2005_rst), .Q(I2536) );
and I_73 (I1970,I2443,I2536);
not I_74 (I2600_rst,I1301_rst);
not I_75 (I2617,I1982);
nor I_76 (I2634,I1967,I1994);
nand I_77 (I2651,I2634,I1970);
DFFARX1 I_78  ( .D(I2651), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I2574) );
nor I_79 (I2682,I2617,I1967);
nand I_80 (I2699,I2682,I1985);
not I_81 (I2589,I2699);
DFFARX1 I_82  ( .D(I2699), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I2571) );
not I_83 (I2744,I1967);
not I_84 (I2761,I2744);
not I_85 (I2778,I1997);
nor I_86 (I2795,I2778,I1979);
and I_87 (I2812,I2795,I1988);
or I_88 (I2829,I2812,I1973);
DFFARX1 I_89  ( .D(I2829), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I2846) );
nor I_90 (I2863,I2846,I2699);
nor I_91 (I2880,I2846,I2761);
nand I_92 (I2586,I2651,I2880);
nand I_93 (I2911,I2617,I1997);
nand I_94 (I2928,I2911,I2846);
and I_95 (I2945,I2911,I2928);
DFFARX1 I_96  ( .D(I2945), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I2568) );
DFFARX1 I_97  ( .D(I2911), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I2976) );
and I_98 (I2565,I2744,I2976);
DFFARX1 I_99  ( .D(I1976), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I3007) );
not I_100 (I3024,I3007);
nor I_101 (I3041,I2699,I3024);
and I_102 (I3058,I3007,I3041);
nand I_103 (I2580,I3007,I2761);
DFFARX1 I_104  ( .D(I3007), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I3089) );
not I_105 (I2577,I3089);
DFFARX1 I_106  ( .D(I1991), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I3120) );
not I_107 (I3137,I3120);
or I_108 (I3154,I3137,I3058);
DFFARX1 I_109  ( .D(I3154), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I2583) );
nand I_110 (I2592,I3137,I2863);
DFFARX1 I_111  ( .D(I3137), .CLK(I1294_clk), .RSTB(I2600_rst), .Q(I2562) );
not I_112 (I3246_rst,I1301_rst);
not I_113 (I3263,I2568);
nor I_114 (I3280,I2565,I2589);
nand I_115 (I3297,I3280,I2586);
nor I_116 (I3314,I3263,I2565);
nand I_117 (I3331,I3314,I2592);
not I_118 (I3348,I3331);
not I_119 (I3365,I2565);
nor I_120 (I3235,I3331,I3365);
not I_121 (I3396,I3365);
nand I_122 (I3220,I3331,I3396);
not I_123 (I3427,I2583);
nor I_124 (I3444,I3427,I2574);
and I_125 (I3461,I3444,I2571);
or I_126 (I3478,I3461,I2580);
DFFARX1 I_127  ( .D(I3478), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3495) );
nor I_128 (I3512,I3495,I3348);
DFFARX1 I_129  ( .D(I3495), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3529) );
not I_130 (I3217,I3529);
nand I_131 (I3560,I3263,I2583);
and I_132 (I3577,I3560,I3512);
DFFARX1 I_133  ( .D(I3560), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3214) );
DFFARX1 I_134  ( .D(I2562), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3608) );
nor I_135 (I3625,I3608,I3331);
nand I_136 (I3232,I3495,I3625);
nor I_137 (I3656,I3608,I3396);
not I_138 (I3229,I3608);
nand I_139 (I3687,I3608,I3297);
and I_140 (I3704,I3365,I3687);
DFFARX1 I_141  ( .D(I3704), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3208) );
DFFARX1 I_142  ( .D(I3608), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3211) );
DFFARX1 I_143  ( .D(I2577), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3749) );
not I_144 (I3766,I3749);
nand I_145 (I3783,I3766,I3331);
and I_146 (I3800,I3560,I3783);
DFFARX1 I_147  ( .D(I3800), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3238) );
or I_148 (I3831,I3766,I3577);
DFFARX1 I_149  ( .D(I3831), .CLK(I1294_clk), .RSTB(I3246_rst), .Q(I3223) );
nand I_150 (I3226,I3766,I3656);
endmodule


