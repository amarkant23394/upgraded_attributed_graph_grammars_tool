module test_I10253(I7621,I7559,I1477,I10185,I7535,I1470,I10253);
input I7621,I7559,I1477,I10185,I7535,I1470;
output I10253;
wire I10086,I10219,I7570,I10236,I7541,I7544,I10052,I10202,I10103,I10069;
nor I_0(I10253,I10103,I10236);
and I_1(I10086,I10069,I7544);
DFFARX1 I_2(I10202,I1470,I10052,,,I10219,);
not I_3(I7570,I1477);
not I_4(I10236,I10219);
DFFARX1 I_5(I1470,I7570,,,I7541,);
DFFARX1 I_6(I7621,I1470,I7570,,,I7544,);
not I_7(I10052,I1477);
and I_8(I10202,I10185,I7541);
DFFARX1 I_9(I10086,I1470,I10052,,,I10103,);
nand I_10(I10069,I7559,I7535);
endmodule


