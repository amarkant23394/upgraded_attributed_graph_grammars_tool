module test_I14131(I1477,I11953,I12106,I12524,I1470,I13970,I14131);
input I1477,I11953,I12106,I12524,I1470,I13970;
output I14131;
wire I14004,I13792,I14049,I11941,I13775,I13987,I11965,I11947,I14114,I12349,I13809,I11962,I14066,I13826,I11956;
DFFARX1 I_0(I13987,I1470,I13775,,,I14004,);
nand I_1(I13792,I11953,I11965);
DFFARX1 I_2(I11962,I1470,I13775,,,I14049,);
DFFARX1 I_3(I1470,,,I11941,);
and I_4(I14131,I13826,I14114);
not I_5(I13775,I1477);
and I_6(I13987,I13970,I11941);
DFFARX1 I_7(I1470,,,I11965,);
nand I_8(I11947,I12106,I12524);
nand I_9(I14114,I14066,I14004);
DFFARX1 I_10(I1470,,,I12349,);
and I_11(I13809,I13792,I11947);
nor I_12(I11962,I12349);
and I_13(I14066,I14049,I11956);
DFFARX1 I_14(I13809,I1470,I13775,,,I13826,);
not I_15(I11956,I12349);
endmodule


