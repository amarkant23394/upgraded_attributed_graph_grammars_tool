module test_I10287(I1477,I8124,I7547,I7669,I7714,I7562,I1470,I7915,I10287);
input I1477,I8124,I7547,I7669,I7714,I7562,I1470,I7915;
output I10287;
wire I10154,I10185,I10202,I10120,I7538,I10219,I7553,I10052,I7946,I7535,I7541,I7570,I10137;
nand I_0(I10154,I10137,I10120);
nand I_1(I10185,I7547,I7562);
and I_2(I10202,I10185,I7541);
nor I_3(I10120,I7538,I7535);
DFFARX1 I_4(I7915,I1470,I7570,,,I7538,);
DFFARX1 I_5(I10202,I1470,I10052,,,I10219,);
DFFARX1 I_6(I8124,I1470,I7570,,,I7553,);
not I_7(I10052,I1477);
DFFARX1 I_8(I1470,I7570,,,I7946,);
and I_9(I7535,I7714,I7946);
DFFARX1 I_10(I7669,I1470,I7570,,,I7541,);
not I_11(I7570,I1477);
DFFARX1 I_12(I7553,I1470,I10052,,,I10137,);
and I_13(I10287,I10219,I10154);
endmodule


