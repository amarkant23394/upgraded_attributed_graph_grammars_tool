module test_I2181(I1477,I2181);
input I1477;
output I2181;
wire ;
not I_0(I2181,I1477);
endmodule


