module test_I14520(I1477,I1470,I13443,I14520);
input I1477,I1470,I13443;
output I14520;
wire I13313,I13697,I13330,I13680,I13601,I13180,I13197,I13168,I14503,I13174,I11272,I13508,I11278,I11302,I13296,I13491;
DFFARX1 I_0(I1470,I13197,,,I13313,);
or I_1(I13697,I13296,I13680);
DFFARX1 I_2(I13313,I1470,I13197,,,I13330,);
and I_3(I13680,I13601,I13443);
DFFARX1 I_4(I1470,I13197,,,I13601,);
not I_5(I13180,I13508);
not I_6(I13197,I1477);
not I_7(I13168,I13330);
nand I_8(I14503,I13180,I13168);
and I_9(I14520,I14503,I13174);
DFFARX1 I_10(I13697,I1470,I13197,,,I13174,);
DFFARX1 I_11(I1470,,,I11272,);
and I_12(I13508,I13491,I11272);
DFFARX1 I_13(I1470,,,I11278,);
DFFARX1 I_14(I1470,,,I11302,);
nor I_15(I13296,I11278,I11302);
DFFARX1 I_16(I1470,I13197,,,I13491,);
endmodule


