module test_final(IN_1_2_l_6,IN_2_2_l_6,G1_3_l_6,G2_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_5_3_l_6,IN_7_3_l_6,IN_8_3_l_6,IN_10_3_l_6,IN_11_3_l_6,blif_reset_net_0_r_8,blif_clk_net_0_r_8,ACVQN2_0_r_8,n_266_and_0_0_r_8,ACVQN1_2_r_8,P6_2_r_8,n_429_or_0_3_r_8,G78_3_r_8,n_576_3_r_8,n_102_3_r_8,n_547_3_r_8,n_42_5_r_8,G199_5_r_8);
input IN_1_2_l_6,IN_2_2_l_6,G1_3_l_6,G2_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_5_3_l_6,IN_7_3_l_6,IN_8_3_l_6,IN_10_3_l_6,IN_11_3_l_6,blif_reset_net_0_r_8,blif_clk_net_0_r_8;
output ACVQN2_0_r_8,n_266_and_0_0_r_8,ACVQN1_2_r_8,P6_2_r_8,n_429_or_0_3_r_8,G78_3_r_8,n_576_3_r_8,n_102_3_r_8,n_547_3_r_8,n_42_5_r_8,G199_5_r_8;
wire ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6,ACVQN1_2_l_6,P6_2_l_6,P6_internal_2_l_6,n_429_or_0_3_l_6,n12_3_l_6,n_431_3_l_6,G78_3_l_6,n_576_3_l_6,n11_3_l_6,n_102_3_l_6,n_547_3_l_6,n13_3_l_6,n14_3_l_6,n15_3_l_6,n16_3_l_6,ACVQN1_0_r_6,P6_internal_2_r_6,n12_3_r_6,n_431_3_r_6,n11_3_r_6,n13_3_r_6,n14_3_r_6,n15_3_r_6,n16_3_r_6,N3_5_r_6,n3_5_r_6,n1_0_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8,ACVQN1_0_l_8,N1_1_l_8,G199_1_l_8,G214_1_l_8,n3_1_l_8,n_42_5_l_8,N3_5_l_8,G199_5_l_8,n3_5_l_8,ACVQN1_0_r_8,P6_internal_2_r_8,n12_3_r_8,n_431_3_r_8,n11_3_r_8,n13_3_r_8,n14_3_r_8,n15_3_r_8,n16_3_r_8,N3_5_r_8,n3_5_r_8;
DFFARX1 I_0(G78_3_l_6,blif_clk_net_0_r_8,n1_0_r_8,ACVQN2_0_r_6,);
and I_1(n_266_and_0_0_r_6,n_429_or_0_3_l_6,ACVQN1_0_r_6);
DFFARX1 I_2(G78_3_l_6,blif_clk_net_0_r_8,n1_0_r_8,ACVQN1_2_r_6,);
not I_3(P6_2_r_6,P6_internal_2_r_6);
nand I_4(n_429_or_0_3_r_6,n_102_3_l_6,n12_3_r_6);
DFFARX1 I_5(n_431_3_r_6,blif_clk_net_0_r_8,n1_0_r_8,G78_3_r_6,);
nand I_6(n_576_3_r_6,P6_2_l_6,n11_3_r_6);
not I_7(n_102_3_r_6,ACVQN1_2_l_6);
nand I_8(n_547_3_r_6,n_576_3_l_6,n13_3_r_6);
nor I_9(n_42_5_r_6,ACVQN1_2_l_6,n_429_or_0_3_l_6);
DFFARX1 I_10(N3_5_r_6,blif_clk_net_0_r_8,n1_0_r_8,G199_5_r_6,);
DFFARX1 I_11(IN_2_2_l_6,blif_clk_net_0_r_8,n1_0_r_8,ACVQN1_2_l_6,);
not I_12(P6_2_l_6,P6_internal_2_l_6);
DFFARX1 I_13(IN_1_2_l_6,blif_clk_net_0_r_8,n1_0_r_8,P6_internal_2_l_6,);
nand I_14(n_429_or_0_3_l_6,G1_3_l_6,n12_3_l_6);
not I_15(n12_3_l_6,IN_5_3_l_6);
or I_16(n_431_3_l_6,IN_8_3_l_6,n14_3_l_6);
DFFARX1 I_17(n_431_3_l_6,blif_clk_net_0_r_8,n1_0_r_8,G78_3_l_6,);
nand I_18(n_576_3_l_6,IN_7_3_l_6,n11_3_l_6);
nor I_19(n11_3_l_6,G2_3_l_6,n12_3_l_6);
not I_20(n_102_3_l_6,G2_3_l_6);
nand I_21(n_547_3_l_6,IN_11_3_l_6,n13_3_l_6);
nor I_22(n13_3_l_6,G2_3_l_6,IN_10_3_l_6);
and I_23(n14_3_l_6,IN_2_3_l_6,n15_3_l_6);
nor I_24(n15_3_l_6,IN_4_3_l_6,n16_3_l_6);
not I_25(n16_3_l_6,G1_3_l_6);
DFFARX1 I_26(G78_3_l_6,blif_clk_net_0_r_8,n1_0_r_8,ACVQN1_0_r_6,);
DFFARX1 I_27(n_576_3_l_6,blif_clk_net_0_r_8,n1_0_r_8,P6_internal_2_r_6,);
not I_28(n12_3_r_6,P6_2_l_6);
or I_29(n_431_3_r_6,n_429_or_0_3_l_6,n14_3_r_6);
nor I_30(n11_3_r_6,ACVQN1_2_l_6,n12_3_r_6);
nor I_31(n13_3_r_6,ACVQN1_2_l_6,n_547_3_l_6);
and I_32(n14_3_r_6,ACVQN1_2_l_6,n15_3_r_6);
nor I_33(n15_3_r_6,P6_2_l_6,n16_3_r_6);
not I_34(n16_3_r_6,n_102_3_l_6);
and I_35(N3_5_r_6,n_102_3_l_6,n3_5_r_6);
nand I_36(n3_5_r_6,n_429_or_0_3_l_6,n_547_3_l_6);
DFFARX1 I_37(n_266_and_0_0_l_8,blif_clk_net_0_r_8,n1_0_r_8,ACVQN2_0_r_8,);
and I_38(n_266_and_0_0_r_8,G199_5_l_8,ACVQN1_0_r_8);
DFFARX1 I_39(G199_5_l_8,blif_clk_net_0_r_8,n1_0_r_8,ACVQN1_2_r_8,);
not I_40(P6_2_r_8,P6_internal_2_r_8);
nand I_41(n_429_or_0_3_r_8,G199_5_l_8,n12_3_r_8);
DFFARX1 I_42(n_431_3_r_8,blif_clk_net_0_r_8,n1_0_r_8,G78_3_r_8,);
nand I_43(n_576_3_r_8,n_42_5_l_8,n11_3_r_8);
not I_44(n_102_3_r_8,n_266_and_0_0_l_8);
nand I_45(n_547_3_r_8,ACVQN2_0_l_8,n13_3_r_8);
nor I_46(n_42_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8);
DFFARX1 I_47(N3_5_r_8,blif_clk_net_0_r_8,n1_0_r_8,G199_5_r_8,);
not I_48(n1_0_r_8,blif_reset_net_0_r_8);
DFFARX1 I_49(n_576_3_r_6,blif_clk_net_0_r_8,n1_0_r_8,ACVQN2_0_l_8,);
and I_50(n_266_and_0_0_l_8,ACVQN1_0_l_8,ACVQN2_0_r_6);
DFFARX1 I_51(P6_2_r_6,blif_clk_net_0_r_8,n1_0_r_8,ACVQN1_0_l_8,);
and I_52(N1_1_l_8,n3_1_l_8,G199_5_r_6);
DFFARX1 I_53(N1_1_l_8,blif_clk_net_0_r_8,n1_0_r_8,G199_1_l_8,);
DFFARX1 I_54(n_42_5_r_6,blif_clk_net_0_r_8,n1_0_r_8,G214_1_l_8,);
nand I_55(n3_1_l_8,n_266_and_0_0_r_6,ACVQN1_2_r_6);
nor I_56(n_42_5_l_8,n_429_or_0_3_r_6,n_102_3_r_6);
and I_57(N3_5_l_8,n3_5_l_8,n_547_3_r_6);
DFFARX1 I_58(N3_5_l_8,blif_clk_net_0_r_8,n1_0_r_8,G199_5_l_8,);
nand I_59(n3_5_l_8,n_429_or_0_3_r_6,G78_3_r_6);
DFFARX1 I_60(G214_1_l_8,blif_clk_net_0_r_8,n1_0_r_8,ACVQN1_0_r_8,);
DFFARX1 I_61(G214_1_l_8,blif_clk_net_0_r_8,n1_0_r_8,P6_internal_2_r_8,);
not I_62(n12_3_r_8,G199_1_l_8);
or I_63(n_431_3_r_8,n_42_5_l_8,n14_3_r_8);
nor I_64(n11_3_r_8,n_266_and_0_0_l_8,n12_3_r_8);
nor I_65(n13_3_r_8,n_266_and_0_0_l_8,G199_1_l_8);
and I_66(n14_3_r_8,ACVQN2_0_l_8,n15_3_r_8);
nor I_67(n15_3_r_8,G199_1_l_8,n16_3_r_8);
not I_68(n16_3_r_8,G199_5_l_8);
and I_69(N3_5_r_8,n_42_5_l_8,n3_5_r_8);
nand I_70(n3_5_r_8,ACVQN2_0_l_8,G214_1_l_8);
endmodule


