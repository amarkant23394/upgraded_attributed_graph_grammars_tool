module test_I3041(I2268,I2022,I1294,I2234,I1301,I3041);
input I2268,I2022,I1294,I2234,I1301;
output I3041;
wire I2203,I3024,I2583,I1902,I2039,I1908,I2634,I2617,I1929,I1937,I2945,I2702,I1926;
DFFARX1 I_0(I1294,I1937,,,I2203,);
nand I_1(I3024,I2945,I2634);
not I_2(I2583,I1301);
and I_3(I1902,I2234,I2203);
DFFARX1 I_4(I2022,I1294,I1937,,,I2039,);
and I_5(I3041,I2702,I3024);
not I_6(I1908,I2039);
nand I_7(I2634,I2617,I1929);
nor I_8(I2617,I1908,I1926);
DFFARX1 I_9(I2268,I1294,I1937,,,I1929,);
not I_10(I1937,I1301);
DFFARX1 I_11(I1902,I1294,I2583,,,I2945,);
not I_12(I2702,I1908);
nor I_13(I1926,I2234);
endmodule


