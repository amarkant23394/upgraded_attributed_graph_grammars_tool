module Benchmark_testing500(I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I251,I258,I5181,I5289,I5325,I5415,I5514,I5532,I5577,I5595,I5613,I5640,I10455,I10563,I10599,I10689,I10788,I10806,I10851,I10869,I10887,I10914);
input I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I251,I258;
output I5181,I5289,I5325,I5415,I5514,I5532,I5577,I5595,I5613,I5640,I10455,I10563,I10599,I10689,I10788,I10806,I10851,I10869,I10887,I10914;
wire I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I251,I258,I267,I294,I312,I321,I339,I366,I375,I393,I411,I429,I447,I465,I483,I501,I528,I537,I555,I573,I591,I609,I627,I645,I672,I690,I699,I717,I735,I753,I780,I789,I807,I825,I852,I861,I879,I897,I924,I942,I951,I978,I987,I1005,I1023,I1041,I1059,I1077,I1095,I1122,I1131,I1149,I1167,I1185,I1212,I1221,I1239,I1257,I1275,I1293,I1320,I1329,I1347,I1365,I1392,I1401,I1419,I1437,I1455,I1482,I1491,I1509,I1527,I1554,I1572,I1581,I1599,I1617,I1644,I1662,I1680,I1698,I1707,I1725,I1743,I1770,I1779,I1797,I1815,I1833,I1851,I1878,I1887,I1914,I1923,I1941,I1959,I1977,I1995,I2022,I2031,I2049,I2067,I2085,I2112,I2130,I2139,I2157,I2184,I2193,I2211,I2229,I2247,I2265,I2283,I2301,I2328,I2337,I2355,I2373,I2400,I2409,I2427,I2445,I2472,I2481,I2508,I2517,I2535,I2553,I2571,I2589,I2616,I2625,I2643,I2661,I2679,I2697,I2715,I2742,I2751,I2769,I2787,I2814,I2823,I2850,I2859,I2877,I2895,I2913,I2931,I2958,I2967,I2985,I3003,I3021,I3048,I3057,I3075,I3102,I3111,I3138,I3147,I3165,I3183,I3201,I3228,I3237,I3255,I3273,I3291,I3318,I3327,I3354,I3363,I3381,I3408,I3417,I3435,I3462,I3471,I3489,I3516,I3525,I3543,I3561,I3588,I3606,I3615,I3633,I3651,I3669,I3687,I3714,I3723,I3750,I3768,I3777,I3795,I3813,I3831,I3849,I3876,I3885,I3912,I3930,I3939,I3957,I3984,I3993,I4011,I4029,I4047,I4065,I4083,I4101,I4119,I4137,I4155,I4173,I4191,I4209,I4227,I4254,I4263,I4290,I4299,I4317,I4335,I4353,I4380,I4389,I4416,I4425,I4443,I4461,I4479,I4506,I4515,I4533,I4551,I4578,I4587,I4614,I4623,I4641,I4659,I4677,I4695,I4722,I4731,I4749,I4767,I4785,I4812,I4821,I4839,I4866,I4875,I4902,I4911,I4929,I4947,I4965,I4992,I5001,I5019,I5037,I5055,I5082,I5091,I5118,I5127,I5145,I5172,I5199,I5226,I5235,I5253,I5280,I5307,I5352,I5370,I5379,I5397,I5433,I5451,I5478,I5487,I5541,I5559,I5649,I5676,I5685,I5712,I5730,I5739,I5757,I5775,I5793,I5820,I5829,I5847,I5865,I5892,I5901,I5919,I5937,I5955,I5973,I6000,I6018,I6027,I6045,I6063,I6081,I6108,I6117,I6135,I6153,I6171,I6189,I6207,I6225,I6243,I6261,I6288,I6297,I6315,I6333,I6360,I6378,I6396,I6405,I6423,I6450,I6459,I6477,I6504,I6513,I6531,I6549,I6567,I6594,I6603,I6621,I6639,I6657,I6675,I6693,I6720,I6729,I6756,I6765,I6783,I6801,I6819,I6846,I6855,I6873,I6891,I6918,I6927,I6954,I6963,I6981,I6999,I7017,I7035,I7062,I7071,I7089,I7107,I7125,I7152,I7161,I7179,I7206,I7215,I7242,I7251,I7269,I7287,I7305,I7332,I7341,I7359,I7377,I7395,I7422,I7431,I7458,I7476,I7485,I7503,I7521,I7539,I7566,I7575,I7602,I7611,I7629,I7647,I7674,I7683,I7710,I7719,I7737,I7755,I7782,I7791,I7809,I7827,I7845,I7872,I7881,I7899,I7917,I7935,I7953,I7980,I7998,I8007,I8034,I8043,I8070,I8088,I8097,I8115,I8133,I8151,I8169,I8187,I8205,I8223,I8241,I8259,I8277,I8295,I8322,I8331,I8349,I8367,I8394,I8403,I8421,I8439,I8466,I8475,I8493,I8511,I8538,I8547,I8565,I8583,I8610,I8619,I8637,I8655,I8682,I8691,I8718,I8727,I8745,I8763,I8781,I8799,I8826,I8835,I8853,I8871,I8889,I8916,I8925,I8943,I8970,I8979,I9006,I9015,I9033,I9051,I9069,I9096,I9105,I9123,I9141,I9159,I9186,I9195,I9222,I9231,I9258,I9276,I9285,I9303,I9321,I9339,I9366,I9375,I9393,I9411,I9438,I9447,I9465,I9483,I9501,I9519,I9546,I9564,I9573,I9591,I9609,I9627,I9654,I9663,I9681,I9699,I9717,I9735,I9753,I9771,I9789,I9807,I9834,I9843,I9861,I9879,I9906,I9924,I9942,I9951,I9969,I9996,I10005,I10023,I10050,I10059,I10077,I10095,I10113,I10140,I10149,I10167,I10185,I10203,I10221,I10239,I10266,I10275,I10302,I10311,I10329,I10347,I10365,I10392,I10401,I10419,I10446,I10473,I10500,I10509,I10527,I10554,I10581,I10626,I10644,I10653,I10671,I10707,I10725,I10752,I10761,I10815,I10833;
not I_0 (I267,I258);
DFFARX1 I_1 (I148,I251,I267,I294,);
DFFARX1 I_2 (I294,I251,I267,I312,);
not I_3 (I321,I312);
not I_4 (I339,I294);
DFFARX1 I_5 (I132,I251,I267,I366,);
not I_6 (I375,I366);
and I_7 (I393,I339,I188);
not I_8 (I411,I204);
nand I_9 (I429,I411,I188);
not I_10 (I447,I212);
nor I_11 (I465,I447,I92);
nand I_12 (I483,I465,I124);
nor I_13 (I501,I483,I429);
DFFARX1 I_14 (I501,I251,I267,I528,);
not I_15 (I537,I483);
not I_16 (I555,I92);
nand I_17 (I573,I555,I188);
nor I_18 (I591,I92,I204);
nand I_19 (I609,I393,I591);
nand I_20 (I627,I339,I92);
nand I_21 (I645,I447,I108);
DFFARX1 I_22 (I645,I251,I267,I672,);
DFFARX1 I_23 (I645,I251,I267,I690,);
not I_24 (I699,I108);
nor I_25 (I717,I699,I164);
and I_26 (I735,I717,I220);
or I_27 (I753,I735,I156);
DFFARX1 I_28 (I753,I251,I267,I780,);
nand I_29 (I789,I780,I411);
nor I_30 (I807,I789,I573);
nor I_31 (I825,I780,I375);
DFFARX1 I_32 (I780,I251,I267,I852,);
not I_33 (I861,I852);
nor I_34 (I879,I861,I537);
not I_35 (I897,I258);
DFFARX1 I_36 (I528,I251,I897,I924,);
DFFARX1 I_37 (I924,I251,I897,I942,);
not I_38 (I951,I942);
DFFARX1 I_39 (I321,I251,I897,I978,);
not I_40 (I987,I879);
nor I_41 (I1005,I924,I987);
not I_42 (I1023,I609);
not I_43 (I1041,I807);
nand I_44 (I1059,I1041,I609);
nor I_45 (I1077,I987,I1059);
nor I_46 (I1095,I978,I1077);
DFFARX1 I_47 (I1041,I251,I897,I1122,);
nor I_48 (I1131,I807,I825);
nand I_49 (I1149,I1131,I672);
nor I_50 (I1167,I1149,I1023);
nand I_51 (I1185,I1167,I879);
DFFARX1 I_52 (I1149,I251,I897,I1212,);
nand I_53 (I1221,I1023,I807);
nor I_54 (I1239,I1023,I807);
nand I_55 (I1257,I1005,I1239);
not I_56 (I1275,I690);
nor I_57 (I1293,I1275,I1221);
DFFARX1 I_58 (I1293,I251,I897,I1320,);
nor I_59 (I1329,I1275,I528);
and I_60 (I1347,I1329,I627);
or I_61 (I1365,I1347,I825);
DFFARX1 I_62 (I1365,I251,I897,I1392,);
nor I_63 (I1401,I1392,I978);
nor I_64 (I1419,I924,I1401);
not I_65 (I1437,I1392);
nor I_66 (I1455,I1437,I1095);
DFFARX1 I_67 (I1455,I251,I897,I1482,);
nand I_68 (I1491,I1437,I1023);
nor I_69 (I1509,I1275,I1491);
not I_70 (I1527,I258);
DFFARX1 I_71 (I1419,I251,I1527,I1554,);
DFFARX1 I_72 (I1554,I251,I1527,I1572,);
not I_73 (I1581,I1572);
nand I_74 (I1599,I1482,I1509);
and I_75 (I1617,I1599,I1320);
DFFARX1 I_76 (I1617,I251,I1527,I1644,);
DFFARX1 I_77 (I1644,I251,I1527,I1662,);
DFFARX1 I_78 (I1644,I251,I1527,I1680,);
DFFARX1 I_79 (I1257,I251,I1527,I1698,);
nand I_80 (I1707,I1698,I1185);
not I_81 (I1725,I1707);
nor I_82 (I1743,I1554,I1725);
DFFARX1 I_83 (I951,I251,I1527,I1770,);
not I_84 (I1779,I1770);
nor I_85 (I1797,I1779,I1581);
nand I_86 (I1815,I1779,I1707);
nand I_87 (I1833,I1212,I1122);
and I_88 (I1851,I1833,I1509);
DFFARX1 I_89 (I1851,I251,I1527,I1878,);
nor I_90 (I1887,I1878,I1554);
DFFARX1 I_91 (I1887,I251,I1527,I1914,);
not I_92 (I1923,I1878);
nor I_93 (I1941,I1320,I1122);
not I_94 (I1959,I1941);
nor I_95 (I1977,I1707,I1959);
nor I_96 (I1995,I1923,I1977);
DFFARX1 I_97 (I1995,I251,I1527,I2022,);
nor I_98 (I2031,I1878,I1959);
nor I_99 (I2049,I1725,I2031);
nor I_100 (I2067,I1878,I1941);
not I_101 (I2085,I258);
DFFARX1 I_102 (I1797,I251,I2085,I2112,);
DFFARX1 I_103 (I1914,I251,I2085,I2130,);
not I_104 (I2139,I2130);
nor I_105 (I2157,I2112,I2139);
DFFARX1 I_106 (I2139,I251,I2085,I2184,);
nor I_107 (I2193,I1914,I1680);
and I_108 (I2211,I2193,I2049);
nor I_109 (I2229,I2211,I1914);
not I_110 (I2247,I1914);
and I_111 (I2265,I2247,I2067);
nand I_112 (I2283,I2265,I1815);
nor I_113 (I2301,I2247,I2283);
DFFARX1 I_114 (I2301,I251,I2085,I2328,);
not I_115 (I2337,I2283);
nand I_116 (I2355,I2139,I2337);
nand I_117 (I2373,I2211,I2337);
DFFARX1 I_118 (I2247,I251,I2085,I2400,);
not I_119 (I2409,I1743);
nor I_120 (I2427,I2409,I2067);
nor I_121 (I2445,I2427,I2229);
DFFARX1 I_122 (I2445,I251,I2085,I2472,);
not I_123 (I2481,I2427);
DFFARX1 I_124 (I2481,I251,I2085,I2508,);
not I_125 (I2517,I2508);
nor I_126 (I2535,I2517,I2427);
nor I_127 (I2553,I2409,I1662);
and I_128 (I2571,I2553,I2022);
or I_129 (I2589,I2571,I2067);
DFFARX1 I_130 (I2589,I251,I2085,I2616,);
not I_131 (I2625,I2616);
nand I_132 (I2643,I2625,I2337);
not I_133 (I2661,I2643);
nand I_134 (I2679,I2643,I2355);
nand I_135 (I2697,I2625,I2211);
not I_136 (I2715,I258);
DFFARX1 I_137 (I2400,I251,I2715,I2742,);
not I_138 (I2751,I2742);
nand I_139 (I2769,I2373,I2328);
and I_140 (I2787,I2769,I2661);
DFFARX1 I_141 (I2787,I251,I2715,I2814,);
not I_142 (I2823,I2328);
DFFARX1 I_143 (I2184,I251,I2715,I2850,);
not I_144 (I2859,I2850);
nor I_145 (I2877,I2859,I2751);
and I_146 (I2895,I2877,I2328);
nor I_147 (I2913,I2859,I2823);
nor I_148 (I2931,I2814,I2913);
DFFARX1 I_149 (I2697,I251,I2715,I2958,);
nor I_150 (I2967,I2958,I2814);
not I_151 (I2985,I2967);
not I_152 (I3003,I2958);
nor I_153 (I3021,I3003,I2895);
DFFARX1 I_154 (I3021,I251,I2715,I3048,);
nand I_155 (I3057,I2157,I2679);
and I_156 (I3075,I3057,I2472);
DFFARX1 I_157 (I3075,I251,I2715,I3102,);
nor I_158 (I3111,I3102,I2958);
DFFARX1 I_159 (I3111,I251,I2715,I3138,);
nand I_160 (I3147,I3102,I3003);
nand I_161 (I3165,I2985,I3147);
not I_162 (I3183,I3102);
nor I_163 (I3201,I3183,I2895);
DFFARX1 I_164 (I3201,I251,I2715,I3228,);
nor I_165 (I3237,I2535,I2679);
or I_166 (I3255,I2958,I3237);
nor I_167 (I3273,I3102,I3237);
or I_168 (I3291,I2814,I3237);
DFFARX1 I_169 (I3237,I251,I2715,I3318,);
not I_170 (I3327,I258);
DFFARX1 I_171 (I3255,I251,I3327,I3354,);
nand I_172 (I3363,I3273,I3048);
and I_173 (I3381,I3363,I3318);
DFFARX1 I_174 (I3381,I251,I3327,I3408,);
nor I_175 (I3417,I3408,I3354);
not I_176 (I3435,I3408);
DFFARX1 I_177 (I3165,I251,I3327,I3462,);
nand I_178 (I3471,I3462,I3273);
not I_179 (I3489,I3471);
DFFARX1 I_180 (I3489,I251,I3327,I3516,);
not I_181 (I3525,I3516);
nor I_182 (I3543,I3354,I3471);
nor I_183 (I3561,I3408,I3543);
DFFARX1 I_184 (I3291,I251,I3327,I3588,);
DFFARX1 I_185 (I3588,I251,I3327,I3606,);
not I_186 (I3615,I3606);
not I_187 (I3633,I3588);
nand I_188 (I3651,I3633,I3435);
nand I_189 (I3669,I3138,I2931);
and I_190 (I3687,I3669,I3138);
DFFARX1 I_191 (I3687,I251,I3327,I3714,);
nor I_192 (I3723,I3714,I3354);
DFFARX1 I_193 (I3723,I251,I3327,I3750,);
DFFARX1 I_194 (I3714,I251,I3327,I3768,);
nor I_195 (I3777,I3228,I2931);
not I_196 (I3795,I3777);
nor I_197 (I3813,I3615,I3795);
nand I_198 (I3831,I3633,I3795);
nor I_199 (I3849,I3354,I3777);
DFFARX1 I_200 (I3777,I251,I3327,I3876,);
not I_201 (I3885,I258);
DFFARX1 I_202 (I3813,I251,I3885,I3912,);
DFFARX1 I_203 (I3912,I251,I3885,I3930,);
not I_204 (I3939,I3930);
not I_205 (I3957,I3912);
DFFARX1 I_206 (I3768,I251,I3885,I3984,);
nand I_207 (I3993,I3984,I3651);
not I_208 (I4011,I3651);
not I_209 (I4029,I3561);
nand I_210 (I4047,I3417,I3750);
and I_211 (I4065,I3417,I3750);
not I_212 (I4083,I3849);
nand I_213 (I4101,I4083,I4029);
nor I_214 (I4119,I4101,I3993);
nor I_215 (I4137,I4011,I4101);
nand I_216 (I4155,I4065,I4137);
not I_217 (I4173,I3525);
nor I_218 (I4191,I4173,I3417);
nor I_219 (I4209,I4191,I3849);
nor I_220 (I4227,I3957,I4209);
DFFARX1 I_221 (I4227,I251,I3885,I4254,);
not I_222 (I4263,I4191);
DFFARX1 I_223 (I4263,I251,I3885,I4290,);
and I_224 (I4299,I3984,I4191);
nor I_225 (I4317,I4173,I3876);
and I_226 (I4335,I4317,I3750);
or I_227 (I4353,I4335,I3831);
DFFARX1 I_228 (I4353,I251,I3885,I4380,);
nor I_229 (I4389,I4380,I4083);
DFFARX1 I_230 (I4389,I251,I3885,I4416,);
nand I_231 (I4425,I4380,I3984);
nand I_232 (I4443,I4083,I4425);
nor I_233 (I4461,I4443,I4047);
not I_234 (I4479,I258);
DFFARX1 I_235 (I4155,I251,I4479,I4506,);
not I_236 (I4515,I4506);
nand I_237 (I4533,I4119,I3939);
and I_238 (I4551,I4533,I4290);
DFFARX1 I_239 (I4551,I251,I4479,I4578,);
not I_240 (I4587,I4416);
DFFARX1 I_241 (I4119,I251,I4479,I4614,);
not I_242 (I4623,I4614);
nor I_243 (I4641,I4623,I4515);
and I_244 (I4659,I4641,I4416);
nor I_245 (I4677,I4623,I4587);
nor I_246 (I4695,I4578,I4677);
DFFARX1 I_247 (I4299,I251,I4479,I4722,);
nor I_248 (I4731,I4722,I4578);
not I_249 (I4749,I4731);
not I_250 (I4767,I4722);
nor I_251 (I4785,I4767,I4659);
DFFARX1 I_252 (I4785,I251,I4479,I4812,);
nand I_253 (I4821,I4254,I4416);
and I_254 (I4839,I4821,I4155);
DFFARX1 I_255 (I4839,I251,I4479,I4866,);
nor I_256 (I4875,I4866,I4722);
DFFARX1 I_257 (I4875,I251,I4479,I4902,);
nand I_258 (I4911,I4866,I4767);
nand I_259 (I4929,I4749,I4911);
not I_260 (I4947,I4866);
nor I_261 (I4965,I4947,I4659);
DFFARX1 I_262 (I4965,I251,I4479,I4992,);
nor I_263 (I5001,I4461,I4416);
or I_264 (I5019,I4722,I5001);
nor I_265 (I5037,I4866,I5001);
or I_266 (I5055,I4578,I5001);
DFFARX1 I_267 (I5001,I251,I4479,I5082,);
not I_268 (I5091,I258);
DFFARX1 I_269 (I5019,I251,I5091,I5118,);
nand I_270 (I5127,I5037,I4812);
and I_271 (I5145,I5127,I5082);
DFFARX1 I_272 (I5145,I251,I5091,I5172,);
nor I_273 (I5181,I5172,I5118);
not I_274 (I5199,I5172);
DFFARX1 I_275 (I4929,I251,I5091,I5226,);
nand I_276 (I5235,I5226,I5037);
not I_277 (I5253,I5235);
DFFARX1 I_278 (I5253,I251,I5091,I5280,);
not I_279 (I5289,I5280);
nor I_280 (I5307,I5118,I5235);
nor I_281 (I5325,I5172,I5307);
DFFARX1 I_282 (I5055,I251,I5091,I5352,);
DFFARX1 I_283 (I5352,I251,I5091,I5370,);
not I_284 (I5379,I5370);
not I_285 (I5397,I5352);
nand I_286 (I5415,I5397,I5199);
nand I_287 (I5433,I4902,I4695);
and I_288 (I5451,I5433,I4902);
DFFARX1 I_289 (I5451,I251,I5091,I5478,);
nor I_290 (I5487,I5478,I5118);
DFFARX1 I_291 (I5487,I251,I5091,I5514,);
DFFARX1 I_292 (I5478,I251,I5091,I5532,);
nor I_293 (I5541,I4992,I4695);
not I_294 (I5559,I5541);
nor I_295 (I5577,I5379,I5559);
nand I_296 (I5595,I5397,I5559);
nor I_297 (I5613,I5118,I5541);
DFFARX1 I_298 (I5541,I251,I5091,I5640,);
not I_299 (I5649,I258);
DFFARX1 I_300 (I116,I251,I5649,I5676,);
and I_301 (I5685,I5676,I228);
DFFARX1 I_302 (I5685,I251,I5649,I5712,);
DFFARX1 I_303 (I84,I251,I5649,I5730,);
not I_304 (I5739,I100);
not I_305 (I5757,I180);
nand I_306 (I5775,I5757,I5739);
nor I_307 (I5793,I5730,I5775);
DFFARX1 I_308 (I5775,I251,I5649,I5820,);
not I_309 (I5829,I5820);
not I_310 (I5847,I244);
nand I_311 (I5865,I5757,I5847);
DFFARX1 I_312 (I5865,I251,I5649,I5892,);
not I_313 (I5901,I5892);
not I_314 (I5919,I236);
nand I_315 (I5937,I5919,I172);
and I_316 (I5955,I5739,I5937);
nor I_317 (I5973,I5865,I5955);
DFFARX1 I_318 (I5973,I251,I5649,I6000,);
DFFARX1 I_319 (I5955,I251,I5649,I6018,);
nor I_320 (I6027,I236,I76);
nor I_321 (I6045,I5865,I6027);
or I_322 (I6063,I236,I76);
nor I_323 (I6081,I140,I196);
DFFARX1 I_324 (I6081,I251,I5649,I6108,);
not I_325 (I6117,I6108);
nor I_326 (I6135,I6117,I5901);
nand I_327 (I6153,I6117,I5730);
not I_328 (I6171,I140);
nand I_329 (I6189,I6171,I5847);
nand I_330 (I6207,I6117,I6189);
nand I_331 (I6225,I6207,I6153);
nand I_332 (I6243,I6189,I6063);
not I_333 (I6261,I258);
DFFARX1 I_334 (I6135,I251,I6261,I6288,);
not I_335 (I6297,I6288);
nand I_336 (I6315,I6000,I6000);
and I_337 (I6333,I6315,I6243);
DFFARX1 I_338 (I6333,I251,I6261,I6360,);
DFFARX1 I_339 (I6360,I251,I6261,I6378,);
DFFARX1 I_340 (I5793,I251,I6261,I6396,);
nand I_341 (I6405,I6396,I6045);
not I_342 (I6423,I6405);
DFFARX1 I_343 (I6423,I251,I6261,I6450,);
not I_344 (I6459,I6450);
nor I_345 (I6477,I6297,I6459);
DFFARX1 I_346 (I5829,I251,I6261,I6504,);
nor I_347 (I6513,I6504,I6360);
nor I_348 (I6531,I6504,I6423);
nand I_349 (I6549,I5712,I6225);
and I_350 (I6567,I6549,I5793);
DFFARX1 I_351 (I6567,I251,I6261,I6594,);
not I_352 (I6603,I6594);
nand I_353 (I6621,I6603,I6504);
nand I_354 (I6639,I6603,I6405);
nor I_355 (I6657,I6018,I6225);
and I_356 (I6675,I6504,I6657);
nor I_357 (I6693,I6603,I6675);
DFFARX1 I_358 (I6693,I251,I6261,I6720,);
nor I_359 (I6729,I6288,I6657);
DFFARX1 I_360 (I6729,I251,I6261,I6756,);
nor I_361 (I6765,I6594,I6657);
not I_362 (I6783,I6765);
nand I_363 (I6801,I6783,I6621);
not I_364 (I6819,I258);
DFFARX1 I_365 (I6720,I251,I6819,I6846,);
not I_366 (I6855,I6846);
nand I_367 (I6873,I6531,I6477);
and I_368 (I6891,I6873,I6378);
DFFARX1 I_369 (I6891,I251,I6819,I6918,);
not I_370 (I6927,I6801);
DFFARX1 I_371 (I6639,I251,I6819,I6954,);
not I_372 (I6963,I6954);
nor I_373 (I6981,I6963,I6855);
and I_374 (I6999,I6981,I6801);
nor I_375 (I7017,I6963,I6927);
nor I_376 (I7035,I6918,I7017);
DFFARX1 I_377 (I6756,I251,I6819,I7062,);
nor I_378 (I7071,I7062,I6918);
not I_379 (I7089,I7071);
not I_380 (I7107,I7062);
nor I_381 (I7125,I7107,I6999);
DFFARX1 I_382 (I7125,I251,I6819,I7152,);
nand I_383 (I7161,I6756,I6531);
and I_384 (I7179,I7161,I6639);
DFFARX1 I_385 (I7179,I251,I6819,I7206,);
nor I_386 (I7215,I7206,I7062);
DFFARX1 I_387 (I7215,I251,I6819,I7242,);
nand I_388 (I7251,I7206,I7107);
nand I_389 (I7269,I7089,I7251);
not I_390 (I7287,I7206);
nor I_391 (I7305,I7287,I6999);
DFFARX1 I_392 (I7305,I251,I6819,I7332,);
nor I_393 (I7341,I6513,I6531);
or I_394 (I7359,I7062,I7341);
nor I_395 (I7377,I7206,I7341);
or I_396 (I7395,I6918,I7341);
DFFARX1 I_397 (I7341,I251,I6819,I7422,);
not I_398 (I7431,I258);
DFFARX1 I_399 (I7377,I251,I7431,I7458,);
DFFARX1 I_400 (I7458,I251,I7431,I7476,);
not I_401 (I7485,I7476);
not I_402 (I7503,I7458);
nand I_403 (I7521,I7422,I7035);
and I_404 (I7539,I7521,I7377);
DFFARX1 I_405 (I7539,I251,I7431,I7566,);
not I_406 (I7575,I7566);
DFFARX1 I_407 (I7269,I251,I7431,I7602,);
and I_408 (I7611,I7602,I7395);
nand I_409 (I7629,I7602,I7395);
nand I_410 (I7647,I7575,I7629);
DFFARX1 I_411 (I7242,I251,I7431,I7674,);
nor I_412 (I7683,I7674,I7611);
DFFARX1 I_413 (I7683,I251,I7431,I7710,);
nor I_414 (I7719,I7674,I7566);
nand I_415 (I7737,I7242,I7359);
and I_416 (I7755,I7737,I7332);
DFFARX1 I_417 (I7755,I251,I7431,I7782,);
nor I_418 (I7791,I7782,I7674);
not I_419 (I7809,I7782);
nor I_420 (I7827,I7809,I7575);
nor I_421 (I7845,I7503,I7827);
DFFARX1 I_422 (I7845,I251,I7431,I7872,);
nor I_423 (I7881,I7809,I7674);
nor I_424 (I7899,I7152,I7359);
nor I_425 (I7917,I7899,I7881);
not I_426 (I7935,I7899);
nand I_427 (I7953,I7629,I7935);
DFFARX1 I_428 (I7899,I251,I7431,I7980,);
DFFARX1 I_429 (I7899,I251,I7431,I7998,);
not I_430 (I8007,I258);
DFFARX1 I_431 (I7980,I251,I8007,I8034,);
nand I_432 (I8043,I8034,I7998);
DFFARX1 I_433 (I7710,I251,I8007,I8070,);
DFFARX1 I_434 (I8070,I251,I8007,I8088,);
not I_435 (I8097,I8088);
not I_436 (I8115,I7719);
nor I_437 (I8133,I7719,I7872);
not I_438 (I8151,I7917);
nand I_439 (I8169,I8115,I8151);
nor I_440 (I8187,I7917,I7719);
and I_441 (I8205,I8187,I8043);
not I_442 (I8223,I7647);
nand I_443 (I8241,I8223,I7485);
nor I_444 (I8259,I7647,I7791);
not I_445 (I8277,I8259);
nand I_446 (I8295,I8133,I8277);
DFFARX1 I_447 (I8259,I251,I8007,I8322,);
nor I_448 (I8331,I7953,I7917);
nor I_449 (I8349,I8331,I7872);
and I_450 (I8367,I8349,I8241);
DFFARX1 I_451 (I8367,I251,I8007,I8394,);
nor I_452 (I8403,I8331,I8169);
or I_453 (I8421,I8259,I8331);
nor I_454 (I8439,I7953,I7710);
DFFARX1 I_455 (I8439,I251,I8007,I8466,);
not I_456 (I8475,I8466);
nand I_457 (I8493,I8475,I8115);
nor I_458 (I8511,I8493,I7872);
DFFARX1 I_459 (I8511,I251,I8007,I8538,);
nor I_460 (I8547,I8475,I8169);
nor I_461 (I8565,I8331,I8547);
not I_462 (I8583,I258);
DFFARX1 I_463 (I8538,I251,I8583,I8610,);
not I_464 (I8619,I8610);
nand I_465 (I8637,I8205,I8421);
and I_466 (I8655,I8637,I8403);
DFFARX1 I_467 (I8655,I251,I8583,I8682,);
not I_468 (I8691,I8097);
DFFARX1 I_469 (I8295,I251,I8583,I8718,);
not I_470 (I8727,I8718);
nor I_471 (I8745,I8727,I8619);
and I_472 (I8763,I8745,I8097);
nor I_473 (I8781,I8727,I8691);
nor I_474 (I8799,I8682,I8781);
DFFARX1 I_475 (I8205,I251,I8583,I8826,);
nor I_476 (I8835,I8826,I8682);
not I_477 (I8853,I8835);
not I_478 (I8871,I8826);
nor I_479 (I8889,I8871,I8763);
DFFARX1 I_480 (I8889,I251,I8583,I8916,);
nand I_481 (I8925,I8322,I8538);
and I_482 (I8943,I8925,I8394);
DFFARX1 I_483 (I8943,I251,I8583,I8970,);
nor I_484 (I8979,I8970,I8826);
DFFARX1 I_485 (I8979,I251,I8583,I9006,);
nand I_486 (I9015,I8970,I8871);
nand I_487 (I9033,I8853,I9015);
not I_488 (I9051,I8970);
nor I_489 (I9069,I9051,I8763);
DFFARX1 I_490 (I9069,I251,I8583,I9096,);
nor I_491 (I9105,I8565,I8538);
or I_492 (I9123,I8826,I9105);
nor I_493 (I9141,I8970,I9105);
or I_494 (I9159,I8682,I9105);
DFFARX1 I_495 (I9105,I251,I8583,I9186,);
not I_496 (I9195,I258);
DFFARX1 I_497 (I8799,I251,I9195,I9222,);
and I_498 (I9231,I9222,I9141);
DFFARX1 I_499 (I9231,I251,I9195,I9258,);
DFFARX1 I_500 (I9159,I251,I9195,I9276,);
not I_501 (I9285,I9006);
not I_502 (I9303,I9186);
nand I_503 (I9321,I9303,I9285);
nor I_504 (I9339,I9276,I9321);
DFFARX1 I_505 (I9321,I251,I9195,I9366,);
not I_506 (I9375,I9366);
not I_507 (I9393,I9123);
nand I_508 (I9411,I9303,I9393);
DFFARX1 I_509 (I9411,I251,I9195,I9438,);
not I_510 (I9447,I9438);
not I_511 (I9465,I9096);
nand I_512 (I9483,I9465,I8916);
and I_513 (I9501,I9285,I9483);
nor I_514 (I9519,I9411,I9501);
DFFARX1 I_515 (I9519,I251,I9195,I9546,);
DFFARX1 I_516 (I9501,I251,I9195,I9564,);
nor I_517 (I9573,I9096,I9033);
nor I_518 (I9591,I9411,I9573);
or I_519 (I9609,I9096,I9033);
nor I_520 (I9627,I9006,I9141);
DFFARX1 I_521 (I9627,I251,I9195,I9654,);
not I_522 (I9663,I9654);
nor I_523 (I9681,I9663,I9447);
nand I_524 (I9699,I9663,I9276);
not I_525 (I9717,I9006);
nand I_526 (I9735,I9717,I9393);
nand I_527 (I9753,I9663,I9735);
nand I_528 (I9771,I9753,I9699);
nand I_529 (I9789,I9735,I9609);
not I_530 (I9807,I258);
DFFARX1 I_531 (I9681,I251,I9807,I9834,);
not I_532 (I9843,I9834);
nand I_533 (I9861,I9546,I9546);
and I_534 (I9879,I9861,I9789);
DFFARX1 I_535 (I9879,I251,I9807,I9906,);
DFFARX1 I_536 (I9906,I251,I9807,I9924,);
DFFARX1 I_537 (I9339,I251,I9807,I9942,);
nand I_538 (I9951,I9942,I9591);
not I_539 (I9969,I9951);
DFFARX1 I_540 (I9969,I251,I9807,I9996,);
not I_541 (I10005,I9996);
nor I_542 (I10023,I9843,I10005);
DFFARX1 I_543 (I9375,I251,I9807,I10050,);
nor I_544 (I10059,I10050,I9906);
nor I_545 (I10077,I10050,I9969);
nand I_546 (I10095,I9258,I9771);
and I_547 (I10113,I10095,I9339);
DFFARX1 I_548 (I10113,I251,I9807,I10140,);
not I_549 (I10149,I10140);
nand I_550 (I10167,I10149,I10050);
nand I_551 (I10185,I10149,I9951);
nor I_552 (I10203,I9564,I9771);
and I_553 (I10221,I10050,I10203);
nor I_554 (I10239,I10149,I10221);
DFFARX1 I_555 (I10239,I251,I9807,I10266,);
nor I_556 (I10275,I9834,I10203);
DFFARX1 I_557 (I10275,I251,I9807,I10302,);
nor I_558 (I10311,I10140,I10203);
not I_559 (I10329,I10311);
nand I_560 (I10347,I10329,I10167);
not I_561 (I10365,I258);
DFFARX1 I_562 (I10077,I251,I10365,I10392,);
nand I_563 (I10401,I10185,I10302);
and I_564 (I10419,I10401,I10059);
DFFARX1 I_565 (I10419,I251,I10365,I10446,);
nor I_566 (I10455,I10446,I10392);
not I_567 (I10473,I10446);
DFFARX1 I_568 (I10266,I251,I10365,I10500,);
nand I_569 (I10509,I10500,I10185);
not I_570 (I10527,I10509);
DFFARX1 I_571 (I10527,I251,I10365,I10554,);
not I_572 (I10563,I10554);
nor I_573 (I10581,I10392,I10509);
nor I_574 (I10599,I10446,I10581);
DFFARX1 I_575 (I9924,I251,I10365,I10626,);
DFFARX1 I_576 (I10626,I251,I10365,I10644,);
not I_577 (I10653,I10644);
not I_578 (I10671,I10626);
nand I_579 (I10689,I10671,I10473);
nand I_580 (I10707,I10302,I10347);
and I_581 (I10725,I10707,I10077);
DFFARX1 I_582 (I10725,I251,I10365,I10752,);
nor I_583 (I10761,I10752,I10392);
DFFARX1 I_584 (I10761,I251,I10365,I10788,);
DFFARX1 I_585 (I10752,I251,I10365,I10806,);
nor I_586 (I10815,I10023,I10347);
not I_587 (I10833,I10815);
nor I_588 (I10851,I10653,I10833);
nand I_589 (I10869,I10671,I10833);
nor I_590 (I10887,I10392,I10815);
DFFARX1 I_591 (I10815,I251,I10365,I10914,);
endmodule


