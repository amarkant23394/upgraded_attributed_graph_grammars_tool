module test_I10930(I9576,I1477,I10845,I1470,I9453,I10930);
input I9576,I1477,I10845,I1470,I9453;
output I10930;
wire I10879,I10647,I9462,I10862,I10896;
or I_0(I10879,I10862,I9462);
not I_1(I10647,I1477);
not I_2(I9462,I9576);
and I_3(I10862,I10845,I9453);
DFFARX1 I_4(I10879,I1470,I10647,,,I10896,);
DFFARX1 I_5(I10896,I1470,I10647,,,I10930,);
endmodule


