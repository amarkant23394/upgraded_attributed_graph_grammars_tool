module test_I3698(I2815,I1294,I1301,I3698);
input I2815,I1294,I1301;
output I3698;
wire I2554,I2866,I2583,I2832,I3246;
not I_0(I2554,I2866);
DFFARX1 I_1(I2832,I1294,I2583,,,I2866,);
not I_2(I2583,I1301);
DFFARX1 I_3(I2815,I1294,I2583,,,I2832,);
not I_4(I3246,I1301);
DFFARX1 I_5(I2554,I1294,I3246,,,I3698,);
endmodule


