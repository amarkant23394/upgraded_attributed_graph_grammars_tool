module test_final(IN_1_2_l_1,IN_2_2_l_1,G1_3_l_1,G2_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_5_3_l_1,IN_7_3_l_1,IN_8_3_l_1,IN_10_3_l_1,IN_11_3_l_1,blif_clk_net_3_r_13,blif_reset_net_3_r_13,n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13);
input IN_1_2_l_1,IN_2_2_l_1,G1_3_l_1,G2_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_5_3_l_1,IN_7_3_l_1,IN_8_3_l_1,IN_10_3_l_1,IN_11_3_l_1,blif_clk_net_3_r_13,blif_reset_net_3_r_13;
output n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13;
wire ACVQN2_0_r_1,n_266_and_0_0_r_1,G199_1_r_1,G214_1_r_1,ACVQN1_2_r_1,P6_2_r_1,n_429_or_0_3_r_1,G78_3_r_1,n_576_3_r_1,n_102_3_r_1,n_547_3_r_1,ACVQN1_2_l_1,P6_2_l_1,P6_internal_2_l_1,n_429_or_0_3_l_1,n12_3_l_1,n_431_3_l_1,G78_3_l_1,n_576_3_l_1,n11_3_l_1,n_102_3_l_1,n_547_3_l_1,n13_3_l_1,n14_3_l_1,n15_3_l_1,n16_3_l_1,ACVQN1_0_r_1,N1_1_r_1,n3_1_r_1,P6_internal_2_r_1,n12_3_r_1,n_431_3_r_1,n11_3_r_1,n13_3_r_1,n14_3_r_1,n15_3_r_1,n16_3_r_1,n2_3_r_13,ACVQN1_2_l_13,P6_2_l_13,P6_internal_2_l_13,n_429_or_0_3_l_13,n12_3_l_13,n_431_3_l_13,G78_3_l_13,n_576_3_l_13,n11_3_l_13,n_102_3_l_13,n_547_3_l_13,n13_3_l_13,n14_3_l_13,n15_3_l_13,n16_3_l_13,n12_3_r_13,n_431_3_r_13,n11_3_r_13,n13_3_r_13,n14_3_r_13,n15_3_r_13,n16_3_r_13,n4_4_r_13,n_87_4_r_13,n7_4_r_13;
DFFARX1 I_0(P6_2_l_1,blif_clk_net_3_r_13,n2_3_r_13,ACVQN2_0_r_1,);
and I_1(n_266_and_0_0_r_1,n_102_3_l_1,ACVQN1_0_r_1);
DFFARX1 I_2(N1_1_r_1,blif_clk_net_3_r_13,n2_3_r_13,G199_1_r_1,);
DFFARX1 I_3(n_576_3_l_1,blif_clk_net_3_r_13,n2_3_r_13,G214_1_r_1,);
DFFARX1 I_4(n_547_3_l_1,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_r_1,);
not I_5(P6_2_r_1,P6_internal_2_r_1);
nand I_6(n_429_or_0_3_r_1,ACVQN1_2_l_1,n12_3_r_1);
DFFARX1 I_7(n_431_3_r_1,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_1,);
nand I_8(n_576_3_r_1,n_547_3_l_1,n11_3_r_1);
not I_9(n_102_3_r_1,n_576_3_l_1);
nand I_10(n_547_3_r_1,P6_2_l_1,n13_3_r_1);
DFFARX1 I_11(IN_2_2_l_1,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_l_1,);
not I_12(P6_2_l_1,P6_internal_2_l_1);
DFFARX1 I_13(IN_1_2_l_1,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_l_1,);
nand I_14(n_429_or_0_3_l_1,G1_3_l_1,n12_3_l_1);
not I_15(n12_3_l_1,IN_5_3_l_1);
or I_16(n_431_3_l_1,IN_8_3_l_1,n14_3_l_1);
DFFARX1 I_17(n_431_3_l_1,blif_clk_net_3_r_13,n2_3_r_13,G78_3_l_1,);
nand I_18(n_576_3_l_1,IN_7_3_l_1,n11_3_l_1);
nor I_19(n11_3_l_1,G2_3_l_1,n12_3_l_1);
not I_20(n_102_3_l_1,G2_3_l_1);
nand I_21(n_547_3_l_1,IN_11_3_l_1,n13_3_l_1);
nor I_22(n13_3_l_1,G2_3_l_1,IN_10_3_l_1);
and I_23(n14_3_l_1,IN_2_3_l_1,n15_3_l_1);
nor I_24(n15_3_l_1,IN_4_3_l_1,n16_3_l_1);
not I_25(n16_3_l_1,G1_3_l_1);
DFFARX1 I_26(n_429_or_0_3_l_1,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_0_r_1,);
and I_27(N1_1_r_1,n_429_or_0_3_l_1,n3_1_r_1);
nand I_28(n3_1_r_1,n_429_or_0_3_l_1,G78_3_l_1);
DFFARX1 I_29(ACVQN1_2_l_1,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_r_1,);
not I_30(n12_3_r_1,n_102_3_l_1);
or I_31(n_431_3_r_1,P6_2_l_1,n14_3_r_1);
nor I_32(n11_3_r_1,G78_3_l_1,n12_3_r_1);
nor I_33(n13_3_r_1,G78_3_l_1,n_576_3_l_1);
and I_34(n14_3_r_1,ACVQN1_2_l_1,n15_3_r_1);
nor I_35(n15_3_r_1,n_576_3_l_1,n16_3_r_1);
not I_36(n16_3_r_1,ACVQN1_2_l_1);
nand I_37(n_429_or_0_3_r_13,n_429_or_0_3_l_13,n12_3_r_13);
DFFARX1 I_38(n_431_3_r_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_13,);
nand I_39(n_576_3_r_13,n_547_3_l_13,n11_3_r_13);
not I_40(n_102_3_r_13,ACVQN1_2_l_13);
nand I_41(n_547_3_r_13,P6_2_l_13,n13_3_r_13);
DFFARX1 I_42(n4_4_r_13,blif_clk_net_3_r_13,n2_3_r_13,G42_4_r_13,);
nor I_43(n_572_4_r_13,P6_2_l_13,n_429_or_0_3_l_13);
or I_44(n_573_4_r_13,ACVQN1_2_l_13,G78_3_l_13);
nor I_45(n_549_4_r_13,n_429_or_0_3_l_13,n7_4_r_13);
or I_46(n_569_4_r_13,n_429_or_0_3_l_13,G78_3_l_13);
nor I_47(n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13);
not I_48(n2_3_r_13,blif_reset_net_3_r_13);
DFFARX1 I_49(n_547_3_r_1,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_l_13,);
not I_50(P6_2_l_13,P6_internal_2_l_13);
DFFARX1 I_51(n_102_3_r_1,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_l_13,);
nand I_52(n_429_or_0_3_l_13,n12_3_l_13,n_429_or_0_3_r_1);
not I_53(n12_3_l_13,G199_1_r_1);
or I_54(n_431_3_l_13,n14_3_l_13,ACVQN2_0_r_1);
DFFARX1 I_55(n_431_3_l_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_l_13,);
nand I_56(n_576_3_l_13,n11_3_l_13,P6_2_r_1);
nor I_57(n11_3_l_13,n12_3_l_13,n_576_3_r_1);
not I_58(n_102_3_l_13,n_576_3_r_1);
nand I_59(n_547_3_l_13,n13_3_l_13,G78_3_r_1);
nor I_60(n13_3_l_13,n_266_and_0_0_r_1,n_576_3_r_1);
and I_61(n14_3_l_13,n15_3_l_13,G214_1_r_1);
nor I_62(n15_3_l_13,n16_3_l_13,ACVQN1_2_r_1);
not I_63(n16_3_l_13,n_429_or_0_3_r_1);
not I_64(n12_3_r_13,n_102_3_l_13);
or I_65(n_431_3_r_13,ACVQN1_2_l_13,n14_3_r_13);
nor I_66(n11_3_r_13,ACVQN1_2_l_13,n12_3_r_13);
nor I_67(n13_3_r_13,ACVQN1_2_l_13,n_576_3_l_13);
and I_68(n14_3_r_13,n_102_3_l_13,n15_3_r_13);
nor I_69(n15_3_r_13,G78_3_l_13,n16_3_r_13);
not I_70(n16_3_r_13,n_429_or_0_3_l_13);
nor I_71(n4_4_r_13,P6_2_l_13,n_547_3_l_13);
not I_72(n_87_4_r_13,P6_2_l_13);
and I_73(n7_4_r_13,n_576_3_l_13,n_87_4_r_13);
endmodule


