module test_I8462(I8394,I1477,I1470,I6144,I8462);
input I8394,I1477,I1470,I6144;
output I8462;
wire I5728,I8428,I8216,I5751,I8411,I8445,I5833,I5725,I5802,I5734;
not I_0(I5728,I5833);
and I_1(I8428,I8411,I5734);
not I_2(I8216,I1477);
not I_3(I5751,I1477);
nor I_4(I8411,I8394,I5725);
or I_5(I8445,I8428,I5728);
DFFARX1 I_6(I5802,I1470,I5751,,,I5833,);
DFFARX1 I_7(I1470,I5751,,,I5725,);
DFFARX1 I_8(I1470,I5751,,,I5802,);
DFFARX1 I_9(I6144,I1470,I5751,,,I5734,);
DFFARX1 I_10(I8445,I1470,I8216,,,I8462,);
endmodule


