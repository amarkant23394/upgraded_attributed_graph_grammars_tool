module test_I17030(I1477,I14982,I12599,I1470,I17030);
input I1477,I14982,I12599,I1470;
output I17030;
wire I12670,I12783,I15276,I14965,I12581,I17013,I15109,I14939,I15454,I15341,I14930,I15016,I12584,I14999,I14942,I15372;
DFFARX1 I_0(I1470,,,I12670,);
DFFARX1 I_1(I1470,,,I12783,);
nand I_2(I15276,I14982,I12599);
not I_3(I14965,I1477);
DFFARX1 I_4(I1470,,,I12581,);
nand I_5(I17013,I14942,I14939);
and I_6(I17030,I17013,I14930);
not I_7(I15109,I12584);
DFFARX1 I_8(I15016,I1470,I14965,,,I14939,);
DFFARX1 I_9(I15372,I1470,I14965,,,I15454,);
DFFARX1 I_10(I15276,I1470,I14965,,,I15341,);
and I_11(I14930,I15109,I15341);
nand I_12(I15016,I14999,I12581);
and I_13(I12584,I12670,I12783);
nor I_14(I14999,I12584);
not I_15(I14942,I15454);
DFFARX1 I_16(I1470,I14965,,,I15372,);
endmodule


