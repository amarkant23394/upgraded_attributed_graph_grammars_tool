module test_I17239(I1477,I16835,I15109,I14942,I1470,I15502,I17239);
input I1477,I16835,I15109,I14942,I1470,I15502;
output I17239;
wire I14927,I14965,I17047,I17013,I16852,I17030,I14957,I17222,I17205,I14939,I16818,I14930,I16869,I15341;
DFFARX1 I_0(I15502,I1470,I14965,,,I14927,);
not I_1(I14965,I1477);
DFFARX1 I_2(I17030,I1470,I16818,,,I17047,);
and I_3(I17239,I17047,I17222);
nand I_4(I17013,I14942,I14939);
and I_5(I16852,I16835,I14957);
and I_6(I17030,I17013,I14930);
nand I_7(I14957,I15502);
nand I_8(I17222,I17205,I16869);
DFFARX1 I_9(I14927,I1470,I16818,,,I17205,);
DFFARX1 I_10(I1470,I14965,,,I14939,);
not I_11(I16818,I1477);
and I_12(I14930,I15109,I15341);
DFFARX1 I_13(I16852,I1470,I16818,,,I16869,);
DFFARX1 I_14(I1470,I14965,,,I15341,);
endmodule


