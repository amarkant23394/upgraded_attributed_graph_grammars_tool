module test_I10137(I6309,I6321,I8011,I1470_clk,I1477_rst,I10137);
input I6309,I6321,I8011,I1470_clk,I1477_rst;
output I10137;
wire I8107,I8124,I7553,I8090,I7977,I10052_rst,I7570_rst,I8028;
not I_0(I8107,I8090);
or I_1(I8124,I8107,I8028);
DFFARX1 I_2 (I8124,I1470_clk,I7570_rst,I7553);
DFFARX1 I_3 (I7553,I1470_clk,I10052_rst,I10137);
DFFARX1 I_4 (I6309,I1470_clk,I7570_rst,I8090);
DFFARX1 I_5 (I6321,I1470_clk,I7570_rst,I7977);
not I_6(I10052_rst,I1477_rst);
not I_7(I7570_rst,I1477_rst);
and I_8(I8028,I7977,I8011);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule