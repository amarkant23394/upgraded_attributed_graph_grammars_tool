module test_I15211(I1477,I15143,I1470,I10636,I12882,I15211);
input I1477,I15143,I1470,I10636,I12882;
output I15211;
wire I12619,I12670,I12913,I13023,I12930,I12608,I15177,I10609,I15160,I15194,I12593,I14965,I12611;
not I_0(I12619,I1477);
DFFARX1 I_1(I1470,I12619,,,I12670,);
DFFARX1 I_2(I1470,I12619,,,I12913,);
DFFARX1 I_3(I10636,I1470,I12619,,,I13023,);
and I_4(I12930,I12913,I10609);
nor I_5(I12608,I13023,I12930);
and I_6(I15177,I15160,I12593);
DFFARX1 I_7(I1470,,,I10609,);
nor I_8(I15160,I15143,I12611);
or I_9(I15194,I15177,I12608);
nand I_10(I12593,I12670,I12882);
DFFARX1 I_11(I15194,I1470,I14965,,,I15211,);
not I_12(I14965,I1477);
DFFARX1 I_13(I1470,I12619,,,I12611,);
endmodule


