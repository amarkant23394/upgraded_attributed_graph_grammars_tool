module test_I8028(I1477,I1470,I7587,I3972,I8028);
input I1477,I1470,I7587,I3972;
output I8028;
wire I6606,I6297,I6321,I7652,I8011,I7570,I6688,I6380,I7994,I6318,I6705,I7977,I7669,I6657;
DFFARX1 I_0(I1470,,,I6606,);
DFFARX1 I_1(I1470,,,I6297,);
nand I_2(I6321,I6705,I6657);
nor I_3(I7652,I7587,I6297);
nor I_4(I8011,I7669,I7994);
not I_5(I7570,I1477);
DFFARX1 I_6(I1470,,,I6688,);
DFFARX1 I_7(I1470,,,I6380,);
and I_8(I8028,I7977,I8011);
not I_9(I7994,I7977);
not I_10(I6318,I6380);
and I_11(I6705,I6688,I3972);
DFFARX1 I_12(I6321,I1470,I7570,,,I7977,);
nand I_13(I7669,I7652,I6318);
nor I_14(I6657,I6606,I6380);
endmodule


