module test_I12041(I1477,I10397,I1470,I10202,I10120,I12041);
input I1477,I10397,I1470,I10202,I10120;
output I12041;
wire I10032,I10219,I10154,I10414,I10020,I11990,I10137,I7553,I10052,I10287,I10103;
nand I_0(I10032,I10137,I10414);
DFFARX1 I_1(I10202,I1470,I10052,,,I10219,);
nand I_2(I10154,I10137,I10120);
nor I_3(I10414,I10103,I10397);
nor I_4(I12041,I11990,I10020);
DFFARX1 I_5(I10287,I1470,I10052,,,I10020,);
not I_6(I11990,I10032);
DFFARX1 I_7(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_8(I1470,,,I7553,);
not I_9(I10052,I1477);
and I_10(I10287,I10219,I10154);
DFFARX1 I_11(I1470,I10052,,,I10103,);
endmodule


