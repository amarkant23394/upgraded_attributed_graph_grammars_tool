module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_5_r_9,n10_9,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
nor I_34(N6147_2_r_9,n62_9,n46_9);
not I_35(N1372_4_r_9,n59_9);
nor I_36(N1508_4_r_9,n58_9,n59_9);
nand I_37(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_38(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_39(n_576_5_r_9,n39_9,n40_9);
not I_40(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_41(n_547_5_r_9,n43_9,N1371_0_r_12);
and I_42(n_42_8_r_9,n44_9,n_549_7_r_12);
DFFARX1 I_43(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_44(N6147_9_r_9,n41_9,n45_9);
nor I_45(N6134_9_r_9,n45_9,n51_9);
nor I_46(I_BUFF_1_9_r_9,n41_9,N1371_0_r_12);
nor I_47(n4_7_l_9,N1508_0_r_12,n_549_7_r_12);
not I_48(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_49(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_50(N3_8_l_9,n57_9,N1508_6_r_12);
DFFARX1 I_51(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_52(n38_9,n63_9);
nor I_53(n_431_5_r_9,G42_7_r_12,n_572_7_r_12);
nor I_54(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_55(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_56(n40_9,n41_9);
nand I_57(n41_9,n_572_7_r_12,n_549_7_r_12);
nor I_58(n42_9,N1507_6_r_12,N6147_9_r_12);
nor I_59(n43_9,n63_9,n41_9);
nor I_60(n44_9,n_569_7_r_12,N6147_9_r_12);
and I_61(n45_9,n52_9,N1371_0_r_12);
nor I_62(n46_9,n47_9,n48_9);
nor I_63(n47_9,n49_9,n50_9);
not I_64(n48_9,n_429_or_0_5_r_9);
not I_65(n49_9,n42_9);
or I_66(n50_9,n63_9,n51_9);
nor I_67(n51_9,N1508_0_r_12,N1507_6_r_12);
nor I_68(n52_9,n49_9,n_572_7_r_12);
nor I_69(n53_9,n54_9,n55_9);
nor I_70(n54_9,n56_9,n_572_7_r_12);
or I_71(n55_9,n44_9,N1507_6_r_12);
not I_72(n56_9,N1371_0_r_12);
nand I_73(n57_9,N1507_6_r_12,N1508_6_r_12);
nor I_74(n58_9,n62_9,n60_9);
nand I_75(n59_9,n51_9,n61_9);
nor I_76(n60_9,n38_9,n44_9);
nor I_77(n61_9,n_569_7_r_12,n_549_7_r_12);
endmodule


