module test_I4773(I1477,I1470,I2146,I4773);
input I1477,I1470,I2146;
output I4773;
wire I4544,I4708,I4725,I4742,I2164,I2263,I2158;
not I_0(I4544,I1477);
nand I_1(I4708,I2146,I2164);
and I_2(I4725,I4708,I2158);
DFFARX1 I_3(I4725,I1470,I4544,,,I4742,);
DFFARX1 I_4(I1470,,,I2164,);
not I_5(I4773,I4742);
DFFARX1 I_6(I1470,,,I2263,);
not I_7(I2158,I2263);
endmodule


