module test_I9771(I1477,I1470,I8298,I5740,I5731,I9771);
input I1477,I1470,I8298,I5740,I5731;
output I9771;
wire I8187,I8216,I8753,I9754,I8178,I8315,I8736,I9491;
DFFARX1 I_0(I8315,I1470,I8216,,,I8187,);
not I_1(I8216,I1477);
not I_2(I8753,I8736);
DFFARX1 I_3(I8187,I1470,I9491,,,I9754,);
and I_4(I9771,I9754,I8178);
DFFARX1 I_5(I8753,I1470,I8216,,,I8178,);
nand I_6(I8315,I8298,I5740);
DFFARX1 I_7(I5731,I1470,I8216,,,I8736,);
not I_8(I9491,I1477);
endmodule


