module test_I15781(I1477,I1470,I13970,I11959,I15781);
input I1477,I1470,I13970,I11959;
output I15781;
wire I13908,I14004,I13749,I13891,I11941,I14131,I13737,I13775,I13987,I13843,I11965,I13755,I15747,I14114,I13826,I15764,I14162,I13925;
not I_0(I13908,I13891);
DFFARX1 I_1(I13987,I1470,I13775,,,I14004,);
nand I_2(I13749,I14162,I13908);
DFFARX1 I_3(I1470,I13775,,,I13891,);
and I_4(I15781,I15764,I13755);
DFFARX1 I_5(I1470,,,I11941,);
and I_6(I14131,I13826,I14114);
DFFARX1 I_7(I14131,I1470,I13775,,,I13737,);
not I_8(I13775,I1477);
and I_9(I13987,I13970,I11941);
nor I_10(I13843,I11959,I11965);
DFFARX1 I_11(I1470,,,I11965,);
nand I_12(I13755,I14004,I13925);
not I_13(I15747,I13749);
nand I_14(I14114,I14004);
DFFARX1 I_15(I1470,I13775,,,I13826,);
nor I_16(I15764,I15747,I13737);
DFFARX1 I_17(I1470,I13775,,,I14162,);
nor I_18(I13925,I13843,I13908);
endmodule


