module test_I10647(I1477_rst,I10647);
input I1477_rst;
output I10647;
wire ;
not I_0(I10647,I1477_rst);
endmodule


