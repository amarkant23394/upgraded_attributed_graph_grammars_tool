module test_I3024(I1294,I2070,I1954,I1301,I3024);
input I1294,I2070,I1954,I1301;
output I3024;
wire I2583,I2313,I1902,I2945,I2268,I2234,I1908,I2634,I1929,I2039,I2203,I1926,I2172,I2251,I1937,I2617,I1304;
nand I_0(I3024,I2945,I2634);
not I_1(I2583,I1301);
DFFARX1 I_2(I1294,I1937,,,I2313,);
and I_3(I1902,I2234,I2203);
DFFARX1 I_4(I1902,I1294,I2583,,,I2945,);
and I_5(I2268,I2070,I2251);
nand I_6(I2234,I1954,I1304);
not I_7(I1908,I2039);
nand I_8(I2634,I2617,I1929);
DFFARX1 I_9(I2268,I1294,I1937,,,I1929,);
DFFARX1 I_10(I1294,I1937,,,I2039,);
DFFARX1 I_11(I2172,I1294,I1937,,,I2203,);
nor I_12(I1926,I2313,I2234);
DFFARX1 I_13(I1294,I1937,,,I2172,);
nand I_14(I2251,I2234);
not I_15(I1937,I1301);
nor I_16(I2617,I1908,I1926);
DFFARX1 I_17(I1294,,,I1304,);
endmodule


