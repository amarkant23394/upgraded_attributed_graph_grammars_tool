module test_I9066(I8998,I1477,I7026,I1470,I9066);
input I8998,I1477,I7026,I1470;
output I9066;
wire I9032,I9049,I7365,I8862,I9015,I6907,I7269,I7348,I6890,I6899,I6869;
DFFARX1 I_0(I9049,I1470,I8862,,,I9066,);
and I_1(I9032,I9015,I6890);
or I_2(I9049,I9032,I6869);
and I_3(I7365,I7026,I7348);
not I_4(I8862,I1477);
nor I_5(I9015,I8998,I6899);
not I_6(I6907,I1477);
DFFARX1 I_7(I1470,I6907,,,I7269,);
nand I_8(I7348,I7269);
not I_9(I6890,I7269);
DFFARX1 I_10(I1470,I6907,,,I6899,);
DFFARX1 I_11(I7365,I1470,I6907,,,I6869,);
endmodule


