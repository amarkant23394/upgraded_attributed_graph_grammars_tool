module test_I15662(I1477,I13792,I13843,I11944,I11947,I11938,I1470,I13970,I15662);
input I1477,I13792,I13843,I11944,I11947,I11938,I1470,I13970;
output I15662;
wire I15645,I14004,I13860,I13891,I11941,I13775,I13987,I13761,I13809,I13740,I13764,I13826,I14162;
nor I_0(I15645,I13761,I13740);
DFFARX1 I_1(I13987,I1470,I13775,,,I14004,);
nor I_2(I13860,I13843,I13826);
nand I_3(I15662,I15645,I13764);
DFFARX1 I_4(I11944,I1470,I13775,,,I13891,);
DFFARX1 I_5(I1470,,,I11941,);
not I_6(I13775,I1477);
and I_7(I13987,I13970,I11941);
nand I_8(I13761,I13891,I13860);
and I_9(I13809,I13792,I11947);
DFFARX1 I_10(I14162,I1470,I13775,,,I13740,);
nor I_11(I13764,I14004,I13826);
DFFARX1 I_12(I13809,I1470,I13775,,,I13826,);
DFFARX1 I_13(I11938,I1470,I13775,,,I14162,);
endmodule


