module test_I8640(I1477,I4533,I1470,I8640);
input I1477,I4533,I1470;
output I8640;
wire I8216,I6110,I8623,I5743,I6028,I6127,I6079,I5802;
not I_0(I8640,I8623);
not I_1(I8216,I1477);
DFFARX1 I_2(I1470,,,I6110,);
DFFARX1 I_3(I5743,I1470,I8216,,,I8623,);
nand I_4(I5743,I6127,I6079);
DFFARX1 I_5(I1470,,,I6028,);
and I_6(I6127,I6110,I4533);
nor I_7(I6079,I6028,I5802);
DFFARX1 I_8(I1470,,,I5802,);
endmodule


