module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_3,n9_3,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_3,n9_3,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_3,n9_3,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_3,n9_3,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_3,n9_3,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_3,n9_3,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_3,n9_3,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_3,n9_3,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_31(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_32(n_573_1_r_3,n26_3,n27_3);
nor I_33(n_549_1_r_3,n40_3,n32_3);
nand I_34(n_569_1_r_3,n27_3,n31_3);
and I_35(n_452_1_r_3,n26_3,n_549_1_r_10);
nor I_36(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_37(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_38(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_39(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_40(n4_1_l_3,n_572_1_r_10,n_549_1_r_10);
not I_41(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_42(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_43(n22_3,G42_1_l_3);
DFFARX1 I_44(G42_1_r_10,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_45(ACVQN2_3_r_10,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_46(n25_3,n25_internal_3);
nor I_47(n4_1_r_3,n40_3,n36_3);
nor I_48(N3_2_r_3,n26_3,n37_3);
nor I_49(n_572_1_l_3,G42_1_r_10,n_42_2_r_10);
DFFARX1 I_50(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_51(n26_3,G199_2_r_10,n_573_1_r_10);
not I_52(n27_3,n_572_1_r_10);
nor I_53(n28_3,n29_3,n_572_1_r_10);
nor I_54(n29_3,n30_3,n_42_2_r_10);
not I_55(n30_3,n_573_1_r_10);
nor I_56(n31_3,n40_3,n_573_1_r_10);
nor I_57(n32_3,n25_3,n33_3);
nand I_58(n33_3,n22_3,n_266_and_0_3_r_10);
or I_59(n34_3,n_572_1_r_10,n_573_1_r_10);
nand I_60(n35_3,ACVQN1_3_r_3,n_266_and_0_3_r_10);
nor I_61(n36_3,n_549_1_r_10,G199_2_r_10);
nor I_62(n37_3,n38_3,n39_3);
not I_63(n38_3,n_572_1_l_3);
nand I_64(n39_3,n27_3,n30_3);
endmodule


