module test_I9960(I8496,I1477,I8315,I9672,I8360,I8267,I1470,I9960);
input I8496,I1477,I8315,I9672,I8360,I8267,I1470;
output I9960;
wire I8202,I8753,I8216,I9816,I9771,I8178,I9909,I9491,I8181,I9754,I8592,I9943,I8736,I9926,I8187,I9576,I9689;
nand I_0(I8202,I8267,I8496);
not I_1(I8753,I8736);
not I_2(I8216,I1477);
DFFARX1 I_3(I1470,I9491,,,I9816,);
and I_4(I9771,I9754,I8178);
DFFARX1 I_5(I8753,I1470,I8216,,,I8178,);
not I_6(I9909,I9816);
not I_7(I9491,I1477);
and I_8(I8181,I8360,I8592);
DFFARX1 I_9(I8187,I1470,I9491,,,I9754,);
DFFARX1 I_10(I1470,I8216,,,I8592,);
and I_11(I9943,I9576,I9926);
DFFARX1 I_12(I1470,I8216,,,I8736,);
nor I_13(I9926,I9689,I9909);
DFFARX1 I_14(I8315,I1470,I8216,,,I8187,);
nor I_15(I9576,I8181,I8202);
or I_16(I9960,I9771,I9943);
DFFARX1 I_17(I9672,I1470,I9491,,,I9689,);
endmodule


