module test_I14347(I14554,I1477,I13186,I1470,I13635,I14347);
input I14554,I1477,I13186,I1470,I13635;
output I14347;
wire I14667,I13189,I14777,I14571,I13197,I14650,I14588,I13165,I14421,I13159,I14438,I14370;
and I_0(I14667,I14650,I13189);
DFFARX1 I_1(I13635,I1470,I13197,,,I13189,);
or I_2(I14777,I14667,I14588);
nor I_3(I14571,I14421,I14554);
not I_4(I13197,I1477);
DFFARX1 I_5(I14777,I1470,I14370,,,I14347,);
DFFARX1 I_6(I13165,I1470,I14370,,,I14650,);
and I_7(I14588,I14438,I14571);
DFFARX1 I_8(I1470,I13197,,,I13165,);
DFFARX1 I_9(I1470,I14370,,,I14421,);
DFFARX1 I_10(I1470,I13197,,,I13159,);
nor I_11(I14438,I13159,I13186);
not I_12(I14370,I1477);
endmodule


