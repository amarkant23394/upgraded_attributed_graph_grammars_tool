module test_I12718(I1477,I11167,I9771,I1470,I9737,I10732,I9471,I12718);
input I1477,I11167,I9771,I1470,I9737,I10732,I9471;
output I12718;
wire I10647,I10615,I10961,I10664,I11184,I10639,I9459,I11201;
not I_0(I10647,I1477);
nor I_1(I12718,I10615,I10639);
DFFARX1 I_2(I10961,I1470,I10647,,,I10615,);
nand I_3(I10961,I10664,I9459);
not I_4(I10664,I9471);
nand I_5(I11184,I11167,I10732);
DFFARX1 I_6(I11201,I1470,I10647,,,I10639,);
nand I_7(I9459,I9771,I9737);
and I_8(I11201,I10961,I11184);
endmodule


