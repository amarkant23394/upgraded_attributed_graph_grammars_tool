module test_I14503(I11296,I1477,I11768,I11293,I1470,I14503);
input I11296,I1477,I11768,I11293,I1470;
output I14503;
wire I13313,I13330,I13180,I13197,I13168,I11272,I13508,I13491,I11310;
DFFARX1 I_0(I11293,I1470,I13197,,,I13313,);
DFFARX1 I_1(I13313,I1470,I13197,,,I13330,);
not I_2(I13180,I13508);
not I_3(I13197,I1477);
not I_4(I13168,I13330);
nand I_5(I14503,I13180,I13168);
DFFARX1 I_6(I11768,I1470,I11310,,,I11272,);
and I_7(I13508,I13491,I11272);
DFFARX1 I_8(I11296,I1470,I13197,,,I13491,);
not I_9(I11310,I1477);
endmodule


