module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_6,blif_reset_net_1_r_6,G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_6,blif_reset_net_1_r_6;
output G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,N3_2_l_6,n4_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_6,n4_6,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_6,n4_6,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_6,n4_6,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_6,n4_6,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_6,n4_6,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_6,n4_6,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_6,n4_6,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_6,n4_6,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_6,n4_6,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_6,blif_clk_net_1_r_6,n4_6,G42_1_r_6,);
nor I_34(n_572_1_r_6,n27_6,n28_6);
nand I_35(n_573_1_r_6,n18_6,n19_6);
nor I_36(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_37(n_569_1_r_6,n19_6,n20_6);
nor I_38(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_39(N1_4_r_6,blif_clk_net_1_r_6,n4_6,G199_4_r_6,);
DFFARX1 I_40(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,G214_4_r_6,);
DFFARX1 I_41(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_6,);
not I_42(P6_5_r_6,P6_5_r_internal_6);
and I_43(N3_2_l_6,n23_6,n_572_1_r_9);
not I_44(n4_6,blif_reset_net_1_r_6);
DFFARX1 I_45(N3_2_l_6,blif_clk_net_1_r_6,n4_6,n27_6,);
not I_46(n17_6,n27_6);
DFFARX1 I_47(G42_1_r_9,blif_clk_net_1_r_6,n4_6,n28_6,);
DFFARX1 I_48(n_572_1_r_9,blif_clk_net_1_r_6,n4_6,n26_6,);
and I_49(N1_4_l_6,n25_6,G42_1_r_9);
DFFARX1 I_50(N1_4_l_6,blif_clk_net_1_r_6,n4_6,n29_6,);
not I_51(n18_6,n29_6);
DFFARX1 I_52(G199_4_r_9,blif_clk_net_1_r_6,n4_6,G214_4_l_6,);
not I_53(n12_6,G214_4_l_6);
nor I_54(n4_1_r_6,n28_6,n22_6);
nor I_55(N1_4_r_6,n12_6,n24_6);
nor I_56(n_42_2_l_6,n_569_1_r_9,n_42_2_r_9);
DFFARX1 I_57(G214_4_l_6,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_6,);
nand I_58(n19_6,n26_6,n_573_1_r_9);
not I_59(n20_6,n_42_2_l_6);
nor I_60(n21_6,n17_6,n28_6);
and I_61(n22_6,n26_6,n_573_1_r_9);
nand I_62(n23_6,n_569_1_r_9,G214_4_r_9);
nor I_63(n24_6,n17_6,n18_6);
nand I_64(n25_6,n_549_1_r_9,G199_2_r_9);
endmodule


