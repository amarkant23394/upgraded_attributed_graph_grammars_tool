module test_I2563(I1301,I2234,I1908,I1294,I2563);
input I1301,I2234,I1908,I1294;
output I2563;
wire I2733,I2583,I2313,I1902,I2203,I2993,I2945,I2702,I3086,I3103,I1920;
nand I_0(I2563,I3103,I2993);
not I_1(I2733,I2702);
not I_2(I2583,I1301);
DFFARX1 I_3(I1294,,,I2313,);
and I_4(I1902,I2234,I2203);
DFFARX1 I_5(I1294,,,I2203,);
nor I_6(I2993,I2945,I2733);
DFFARX1 I_7(I1902,I1294,I2583,,,I2945,);
not I_8(I2702,I1908);
DFFARX1 I_9(I1920,I1294,I2583,,,I3086,);
not I_10(I3103,I3086);
not I_11(I1920,I2313);
endmodule


