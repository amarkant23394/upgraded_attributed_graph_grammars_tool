module test_I17378(I15696,I1477,I1470,I17378);
input I15696,I1477,I1470;
output I17378;
wire I17413,I15959,I17775,I16052,I15585,I15928,I16069;
not I_0(I17413,I1477);
nor I_1(I15959,I15928,I15696);
DFFARX1 I_2(I15585,I1470,I17413,,,I17775,);
DFFARX1 I_3(I1470,,,I16052,);
nand I_4(I15585,I16069,I15959);
DFFARX1 I_5(I17775,I1470,I17413,,,I17378,);
DFFARX1 I_6(I1470,,,I15928,);
not I_7(I16069,I16052);
endmodule


