module test_final(IN_1_1_l,IN_2_1_l,IN_3_1_l,blif_clk_net_8_l,blif_reset_net_8_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,N1372_1_r,N1508_1_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,N1372_10_r,N1508_10_r);
input IN_1_1_l,IN_2_1_l,IN_3_1_l,blif_clk_net_8_l,blif_reset_net_8_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l;
output N1372_1_r,N1508_1_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,N1372_10_r,N1508_10_r;
wire N1372_1_l,N1508_1_l,n4_1_l,n_42_8_l,G199_8_l,N3_8_l,n1_8_l,n3_8_l,N1372_10_l,N1508_10_l,n5_10_l,n6_10_l,n4_1_r,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n6_4_r,n7_4_r,n8_4_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,n5_10_r,n6_10_r;
not I_0(N1372_1_l,n4_1_l);
nor I_1(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_2(n4_1_l,IN_1_1_l,IN_2_1_l);
nor I_3(n_42_8_l,IN_1_8_l,IN_3_8_l);
DFFARX1 I_4(N3_8_l,blif_clk_net_8_l,n1_8_l,G199_8_l,);
and I_5(N3_8_l,IN_6_8_l,n3_8_l);
not I_6(n1_8_l,blif_reset_net_8_l);
nand I_7(n3_8_l,IN_2_8_l,IN_3_8_l);
not I_8(N1372_10_l,n6_10_l);
nor I_9(N1508_10_l,n5_10_l,n6_10_l);
nor I_10(n5_10_l,IN_3_10_l,IN_4_10_l);
nand I_11(n6_10_l,IN_1_10_l,IN_2_10_l);
not I_12(N1372_1_r,n4_1_r);
nor I_13(N1508_1_r,n4_1_r,G199_8_l);
nand I_14(n4_1_r,N1508_1_l,n_42_8_l);
nor I_15(N6147_2_r,n5_2_r,n6_2_r);
nor I_16(n5_2_r,n7_2_r,N1508_10_l);
not I_17(n6_2_r,N6138_2_r);
nor I_18(N6138_2_r,N1508_10_l,G199_8_l);
nor I_19(n7_2_r,N1372_1_l,N1372_10_l);
nor I_20(N6147_3_r,n3_3_r,N1508_1_l);
not I_21(n3_3_r,N6138_3_r);
nor I_22(N6138_3_r,N1508_1_l,N1508_10_l);
not I_23(N1372_4_r,n7_4_r);
nor I_24(N1508_4_r,n6_4_r,n7_4_r);
nor I_25(n6_4_r,n8_4_r,N1372_10_l);
nand I_26(n7_4_r,N1372_10_l,N1508_10_l);
and I_27(n8_4_r,n_42_8_l,G199_8_l);
nor I_28(N1507_6_r,n8_6_r,n9_6_r);
and I_29(N1508_6_r,n6_6_r,N1372_10_l);
nor I_30(n6_6_r,n7_6_r,n8_6_r);
not I_31(n7_6_r,n_42_8_l);
nor I_32(n8_6_r,n9_6_r,N1372_1_l);
and I_33(n9_6_r,N1372_1_l,N1508_1_l);
not I_34(N1372_10_r,n6_10_r);
nor I_35(N1508_10_r,n5_10_r,n6_10_r);
nor I_36(n5_10_r,N1372_1_l,G199_8_l);
nand I_37(n6_10_r,G199_8_l,n_42_8_l);
endmodule


