module test_I7461(I1477,I5368,I5563,I5070,I5642,I5450,I1470,I5082,I7461);
input I1477,I5368,I5563,I5070,I5642,I5450,I1470,I5082;
output I7461;
wire I5659,I5088,I6907,I7221,I5097,I7444,I6975,I7410,I5073,I6992,I5105,I6924,I7427;
or I_0(I5659,I5642,I5563);
DFFARX1 I_1(I5659,I1470,I5105,,,I5088,);
not I_2(I6907,I1477);
nand I_3(I7221,I6924,I5088);
nand I_4(I5097,I5642,I5368);
nand I_5(I7444,I7427,I6992);
nor I_6(I6975,I6924,I5070);
and I_7(I7461,I7221,I7444);
DFFARX1 I_8(I5082,I1470,I6907,,,I7410,);
DFFARX1 I_9(I5450,I1470,I5105,,,I5073,);
nand I_10(I6992,I6975,I5097);
not I_11(I5105,I1477);
not I_12(I6924,I5073);
not I_13(I7427,I7410);
endmodule


