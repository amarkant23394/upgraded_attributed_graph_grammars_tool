module Benchmark_testing5000(I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I252,I260,I268,I276,I284,I292,I300,I308,I316,I324,I332,I340,I348,I356,I364,I372,I380,I388,I396,I404,I412,I420,I428,I436,I444,I452,I460,I468,I476,I484,I492,I500,I508,I515,I522,I17352,I17433,I17469,I17640,I17658,I17685,I17775,I17865,I17883,I35163,I35280,I35370,I35397,I35460,I35487,I35505,I35523,I35550,I52614,I52677,I52731,I52785,I52884,I52920,I52974,I53001,I53019,I70002,I70047,I70092,I70173,I70209,I70308,I70335,I70353,I70371,I87246,I87264,I87327,I87381,I87399,I87498,I87606,I87633,I87651);
input I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I252,I260,I268,I276,I284,I292,I300,I308,I316,I324,I332,I340,I348,I356,I364,I372,I380,I388,I396,I404,I412,I420,I428,I436,I444,I452,I460,I468,I476,I484,I492,I500,I508,I515,I522;
output I17352,I17433,I17469,I17640,I17658,I17685,I17775,I17865,I17883,I35163,I35280,I35370,I35397,I35460,I35487,I35505,I35523,I35550,I52614,I52677,I52731,I52785,I52884,I52920,I52974,I53001,I53019,I70002,I70047,I70092,I70173,I70209,I70308,I70335,I70353,I70371,I87246,I87264,I87327,I87381,I87399,I87498,I87606,I87633,I87651;
wire I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I252,I260,I268,I276,I284,I292,I300,I308,I316,I324,I332,I340,I348,I356,I364,I372,I380,I388,I396,I404,I412,I420,I428,I436,I444,I452,I460,I468,I476,I484,I492,I500,I508,I515,I522,I531,I558,I567,I594,I612,I621,I639,I657,I675,I702,I711,I729,I747,I774,I783,I801,I819,I837,I855,I882,I900,I909,I927,I945,I963,I990,I999,I1017,I1035,I1053,I1071,I1089,I1107,I1125,I1143,I1170,I1188,I1197,I1215,I1242,I1251,I1269,I1287,I1305,I1323,I1341,I1359,I1386,I1395,I1413,I1431,I1458,I1467,I1485,I1503,I1530,I1539,I1566,I1575,I1593,I1611,I1629,I1647,I1674,I1683,I1701,I1719,I1737,I1755,I1773,I1800,I1809,I1827,I1854,I1863,I1881,I1908,I1917,I1935,I1962,I1971,I1989,I2007,I2034,I2052,I2061,I2079,I2097,I2115,I2133,I2160,I2169,I2196,I2214,I2223,I2241,I2259,I2277,I2295,I2322,I2331,I2358,I2367,I2394,I2412,I2421,I2439,I2457,I2475,I2493,I2511,I2529,I2547,I2565,I2583,I2601,I2619,I2646,I2655,I2673,I2691,I2718,I2727,I2745,I2763,I2790,I2799,I2817,I2835,I2862,I2871,I2889,I2907,I2934,I2952,I2961,I2979,I2997,I3015,I3033,I3051,I3078,I3087,I3105,I3132,I3141,I3159,I3177,I3204,I3213,I3231,I3258,I3267,I3285,I3303,I3321,I3339,I3357,I3375,I3393,I3420,I3429,I3447,I3465,I3483,I3501,I3519,I3537,I3555,I3573,I3591,I3618,I3627,I3654,I3672,I3681,I3699,I3717,I3735,I3762,I3771,I3789,I3807,I3834,I3843,I3861,I3879,I3897,I3915,I3942,I3960,I3969,I3987,I4005,I4023,I4050,I4059,I4077,I4095,I4113,I4131,I4149,I4167,I4185,I4203,I4230,I4248,I4257,I4275,I4293,I4311,I4338,I4347,I4374,I4383,I4401,I4419,I4446,I4455,I4482,I4491,I4509,I4527,I4554,I4563,I4581,I4599,I4617,I4644,I4653,I4671,I4689,I4707,I4725,I4752,I4770,I4779,I4806,I4815,I4842,I4860,I4869,I4887,I4905,I4923,I4950,I4959,I4977,I4995,I5022,I5031,I5049,I5067,I5085,I5103,I5130,I5148,I5157,I5175,I5193,I5211,I5238,I5247,I5265,I5283,I5301,I5319,I5337,I5355,I5373,I5391,I5418,I5427,I5445,I5463,I5490,I5499,I5526,I5535,I5553,I5571,I5589,I5607,I5634,I5643,I5661,I5679,I5697,I5724,I5733,I5751,I5778,I5787,I5814,I5823,I5841,I5859,I5877,I5904,I5913,I5931,I5949,I5967,I5994,I6003,I6030,I6039,I6057,I6075,I6102,I6120,I6129,I6147,I6174,I6183,I6201,I6219,I6246,I6264,I6273,I6291,I6318,I6336,I6345,I6363,I6381,I6399,I6417,I6435,I6453,I6480,I6489,I6507,I6525,I6543,I6561,I6588,I6606,I6615,I6633,I6651,I6669,I6696,I6705,I6732,I6741,I6759,I6777,I6804,I6813,I6840,I6849,I6867,I6885,I6912,I6921,I6939,I6957,I6975,I7002,I7011,I7029,I7047,I7065,I7083,I7110,I7128,I7137,I7164,I7173,I7191,I7209,I7236,I7245,I7272,I7281,I7299,I7317,I7335,I7353,I7380,I7389,I7407,I7425,I7443,I7470,I7479,I7497,I7524,I7533,I7560,I7569,I7587,I7605,I7623,I7650,I7659,I7677,I7695,I7713,I7740,I7749,I7776,I7794,I7803,I7821,I7839,I7857,I7884,I7893,I7920,I7929,I7947,I7965,I7992,I8001,I8028,I8037,I8055,I8073,I8100,I8109,I8127,I8145,I8163,I8190,I8199,I8217,I8235,I8253,I8271,I8298,I8316,I8325,I8352,I8361,I8379,I8406,I8415,I8433,I8460,I8469,I8487,I8514,I8523,I8541,I8559,I8586,I8604,I8613,I8631,I8649,I8667,I8685,I8712,I8721,I8748,I8766,I8775,I8793,I8811,I8829,I8847,I8874,I8883,I8910,I8919,I8937,I8955,I8982,I8991,I9018,I9027,I9045,I9063,I9081,I9099,I9126,I9135,I9153,I9171,I9189,I9216,I9225,I9243,I9270,I9279,I9306,I9315,I9333,I9351,I9369,I9396,I9405,I9423,I9441,I9459,I9486,I9495,I9522,I9531,I9549,I9576,I9585,I9603,I9630,I9639,I9657,I9684,I9693,I9711,I9729,I9756,I9774,I9783,I9801,I9819,I9837,I9855,I9882,I9891,I9918,I9936,I9945,I9963,I9981,I9999,I10017,I10044,I10053,I10080,I10098,I10107,I10125,I10152,I10161,I10179,I10197,I10215,I10233,I10251,I10269,I10287,I10314,I10323,I10341,I10359,I10377,I10395,I10413,I10431,I10458,I10476,I10485,I10503,I10521,I10539,I10566,I10575,I10593,I10611,I10638,I10647,I10665,I10683,I10710,I10719,I10746,I10764,I10773,I10791,I10809,I10827,I10845,I10863,I10881,I10899,I10917,I10935,I10953,I10971,I10998,I11007,I11025,I11043,I11070,I11079,I11097,I11115,I11142,I11151,I11169,I11187,I11214,I11223,I11241,I11259,I11286,I11295,I11313,I11331,I11358,I11367,I11394,I11403,I11421,I11439,I11457,I11475,I11502,I11511,I11529,I11547,I11565,I11592,I11601,I11619,I11646,I11655,I11682,I11691,I11709,I11727,I11745,I11772,I11781,I11799,I11817,I11835,I11862,I11871,I11898,I11916,I11925,I11943,I11970,I11979,I11997,I12015,I12033,I12051,I12069,I12087,I12105,I12123,I12141,I12159,I12177,I12195,I12213,I12240,I12249,I12276,I12285,I12303,I12321,I12339,I12366,I12375,I12402,I12411,I12429,I12447,I12465,I12492,I12510,I12519,I12537,I12564,I12573,I12591,I12609,I12627,I12645,I12663,I12681,I12708,I12717,I12735,I12753,I12780,I12789,I12807,I12825,I12852,I12861,I12888,I12897,I12915,I12933,I12951,I12969,I12996,I13005,I13023,I13041,I13059,I13077,I13095,I13122,I13131,I13158,I13176,I13185,I13203,I13221,I13239,I13266,I13275,I13293,I13311,I13338,I13347,I13365,I13383,I13401,I13419,I13446,I13464,I13473,I13491,I13509,I13527,I13554,I13563,I13581,I13599,I13617,I13635,I13653,I13671,I13689,I13707,I13734,I13743,I13761,I13779,I13806,I13815,I13842,I13851,I13869,I13887,I13905,I13923,I13950,I13959,I13977,I13995,I14013,I14040,I14049,I14067,I14094,I14103,I14130,I14139,I14157,I14175,I14193,I14220,I14229,I14247,I14265,I14283,I14310,I14319,I14346,I14364,I14373,I14400,I14409,I14427,I14445,I14463,I14481,I14499,I14517,I14544,I14553,I14571,I14589,I14607,I14634,I14643,I14661,I14679,I14697,I14715,I14742,I14751,I14769,I14787,I14814,I14823,I14841,I14859,I14877,I14904,I14913,I14931,I14949,I14976,I14994,I15003,I15021,I15039,I15066,I15084,I15102,I15120,I15129,I15147,I15165,I15192,I15201,I15219,I15237,I15255,I15273,I15300,I15309,I15336,I15345,I15363,I15381,I15399,I15417,I15444,I15453,I15471,I15489,I15507,I15534,I15543,I15561,I15588,I15597,I15615,I15642,I15651,I15669,I15696,I15705,I15723,I15741,I15768,I15786,I15795,I15813,I15831,I15849,I15867,I15894,I15903,I15930,I15948,I15957,I15975,I15993,I16011,I16029,I16056,I16065,I16092,I16101,I16128,I16137,I16155,I16173,I16191,I16209,I16236,I16245,I16263,I16281,I16299,I16317,I16335,I16353,I16371,I16389,I16407,I16425,I16443,I16461,I16479,I16497,I16515,I16542,I16551,I16578,I16596,I16605,I16623,I16641,I16668,I16677,I16704,I16713,I16731,I16749,I16776,I16785,I16812,I16821,I16839,I16857,I16875,I16893,I16920,I16929,I16947,I16965,I16983,I17010,I17019,I17037,I17064,I17073,I17100,I17109,I17127,I17145,I17163,I17190,I17199,I17217,I17235,I17253,I17280,I17289,I17316,I17325,I17370,I17379,I17397,I17415,I17460,I17487,I17505,I17532,I17541,I17559,I17577,I17595,I17613,I17667,I17703,I17721,I17748,I17757,I17793,I17811,I17829,I17847,I17901,I17928,I17946,I17955,I17973,I17991,I18009,I18036,I18045,I18072,I18081,I18099,I18117,I18144,I18153,I18180,I18189,I18207,I18225,I18252,I18261,I18279,I18297,I18315,I18342,I18351,I18369,I18387,I18405,I18423,I18450,I18468,I18477,I18504,I18513,I18531,I18549,I18576,I18594,I18603,I18621,I18648,I18657,I18675,I18693,I18720,I18738,I18747,I18765,I18792,I18810,I18819,I18837,I18855,I18873,I18891,I18909,I18927,I18954,I18963,I18981,I18999,I19017,I19035,I19062,I19071,I19098,I19116,I19125,I19143,I19161,I19179,I19206,I19215,I19233,I19251,I19278,I19287,I19305,I19323,I19341,I19359,I19386,I19404,I19413,I19431,I19449,I19467,I19494,I19503,I19521,I19539,I19557,I19575,I19593,I19611,I19629,I19647,I19674,I19692,I19701,I19728,I19737,I19755,I19773,I19791,I19809,I19827,I19845,I19872,I19881,I19899,I19917,I19935,I19962,I19971,I19989,I20007,I20025,I20043,I20070,I20079,I20097,I20115,I20142,I20151,I20169,I20187,I20205,I20232,I20241,I20259,I20277,I20304,I20313,I20331,I20358,I20367,I20385,I20412,I20421,I20439,I20466,I20475,I20493,I20511,I20538,I20556,I20565,I20583,I20601,I20619,I20637,I20664,I20673,I20700,I20718,I20727,I20745,I20763,I20781,I20799,I20826,I20835,I20862,I20880,I20889,I20907,I20925,I20943,I20961,I20979,I21006,I21015,I21033,I21060,I21069,I21087,I21105,I21132,I21141,I21159,I21186,I21195,I21213,I21231,I21249,I21267,I21285,I21303,I21321,I21348,I21357,I21375,I21393,I21411,I21429,I21447,I21465,I21483,I21501,I21519,I21546,I21555,I21573,I21591,I21618,I21627,I21654,I21663,I21681,I21699,I21717,I21735,I21762,I21771,I21789,I21807,I21825,I21852,I21861,I21879,I21906,I21915,I21942,I21951,I21969,I21987,I22005,I22032,I22041,I22059,I22077,I22095,I22122,I22131,I22158,I22167,I22194,I22212,I22221,I22239,I22257,I22275,I22302,I22311,I22329,I22347,I22374,I22383,I22401,I22419,I22437,I22455,I22482,I22500,I22509,I22527,I22545,I22563,I22590,I22599,I22617,I22635,I22653,I22671,I22689,I22707,I22725,I22743,I22770,I22779,I22797,I22824,I22833,I22851,I22869,I22887,I22905,I22932,I22941,I22959,I22977,I22995,I23013,I23031,I23049,I23076,I23085,I23103,I23121,I23139,I23157,I23175,I23202,I23211,I23238,I23247,I23274,I23292,I23301,I23319,I23337,I23355,I23382,I23391,I23418,I23436,I23445,I23463,I23481,I23499,I23526,I23535,I23553,I23571,I23598,I23607,I23625,I23643,I23661,I23679,I23706,I23724,I23733,I23751,I23769,I23787,I23814,I23823,I23841,I23859,I23877,I23895,I23913,I23931,I23949,I23967,I23994,I24012,I24021,I24039,I24057,I24084,I24102,I24120,I24138,I24147,I24165,I24183,I24210,I24219,I24237,I24255,I24273,I24291,I24318,I24327,I24354,I24363,I24381,I24399,I24417,I24435,I24462,I24471,I24489,I24507,I24525,I24552,I24561,I24588,I24606,I24615,I24633,I24651,I24669,I24696,I24705,I24723,I24741,I24768,I24777,I24795,I24813,I24831,I24849,I24876,I24894,I24903,I24921,I24939,I24957,I24984,I24993,I25011,I25029,I25047,I25065,I25083,I25101,I25119,I25137,I25164,I25182,I25191,I25218,I25227,I25245,I25263,I25281,I25299,I25317,I25335,I25362,I25371,I25389,I25407,I25425,I25452,I25461,I25479,I25497,I25515,I25533,I25560,I25569,I25587,I25605,I25632,I25641,I25659,I25677,I25695,I25722,I25731,I25749,I25767,I25794,I25812,I25821,I25839,I25866,I25875,I25893,I25911,I25929,I25947,I25965,I25983,I26001,I26028,I26037,I26055,I26073,I26091,I26109,I26127,I26145,I26172,I26190,I26199,I26217,I26235,I26253,I26280,I26289,I26307,I26325,I26352,I26361,I26379,I26397,I26424,I26433,I26460,I26478,I26487,I26505,I26523,I26541,I26568,I26577,I26595,I26613,I26640,I26649,I26667,I26685,I26703,I26721,I26748,I26766,I26775,I26793,I26811,I26829,I26856,I26865,I26883,I26901,I26919,I26937,I26955,I26973,I26991,I27009,I27036,I27045,I27063,I27081,I27108,I27117,I27144,I27153,I27171,I27189,I27207,I27225,I27252,I27261,I27279,I27297,I27315,I27342,I27351,I27369,I27396,I27405,I27432,I27441,I27459,I27477,I27495,I27522,I27531,I27549,I27567,I27585,I27612,I27621,I27648,I27657,I27684,I27693,I27711,I27729,I27747,I27765,I27792,I27801,I27819,I27837,I27855,I27873,I27891,I27909,I27927,I27945,I27963,I27981,I27999,I28017,I28035,I28053,I28071,I28098,I28107,I28134,I28152,I28161,I28179,I28197,I28224,I28233,I28260,I28269,I28287,I28314,I28323,I28341,I28368,I28377,I28395,I28422,I28431,I28449,I28467,I28494,I28512,I28521,I28539,I28557,I28575,I28593,I28620,I28629,I28656,I28674,I28683,I28701,I28719,I28737,I28755,I28782,I28791,I28818,I28836,I28845,I28863,I28881,I28899,I28917,I28935,I28962,I28971,I28989,I29016,I29025,I29043,I29061,I29088,I29097,I29115,I29142,I29151,I29169,I29187,I29205,I29223,I29241,I29259,I29277,I29304,I29313,I29331,I29349,I29367,I29385,I29403,I29421,I29439,I29457,I29475,I29502,I29511,I29538,I29556,I29565,I29583,I29601,I29619,I29646,I29655,I29673,I29691,I29718,I29727,I29745,I29763,I29781,I29799,I29826,I29844,I29853,I29871,I29889,I29907,I29934,I29943,I29961,I29979,I29997,I30015,I30033,I30051,I30069,I30087,I30114,I30132,I30141,I30168,I30177,I30195,I30213,I30231,I30249,I30267,I30285,I30312,I30321,I30339,I30357,I30375,I30402,I30411,I30429,I30447,I30465,I30483,I30510,I30519,I30537,I30555,I30582,I30591,I30609,I30627,I30645,I30672,I30681,I30699,I30717,I30744,I30753,I30780,I30798,I30807,I30825,I30843,I30861,I30888,I30897,I30915,I30933,I30960,I30969,I30987,I31005,I31023,I31041,I31068,I31086,I31095,I31113,I31131,I31149,I31176,I31185,I31203,I31221,I31239,I31257,I31275,I31293,I31311,I31329,I31356,I31365,I31392,I31410,I31419,I31437,I31455,I31473,I31491,I31509,I31527,I31545,I31563,I31581,I31599,I31617,I31644,I31653,I31671,I31689,I31716,I31725,I31743,I31761,I31788,I31797,I31815,I31833,I31860,I31869,I31887,I31905,I31932,I31941,I31968,I31986,I31995,I32013,I32031,I32049,I32076,I32085,I32103,I32121,I32148,I32157,I32175,I32193,I32211,I32229,I32256,I32274,I32283,I32301,I32319,I32337,I32364,I32373,I32391,I32409,I32427,I32445,I32463,I32481,I32499,I32517,I32544,I32562,I32571,I32589,I32607,I32625,I32643,I32661,I32688,I32697,I32715,I32742,I32751,I32769,I32787,I32814,I32823,I32841,I32868,I32877,I32895,I32913,I32931,I32949,I32967,I32985,I33003,I33030,I33039,I33057,I33075,I33093,I33111,I33129,I33147,I33165,I33183,I33201,I33228,I33246,I33255,I33273,I33291,I33318,I33336,I33354,I33372,I33381,I33399,I33417,I33444,I33453,I33471,I33489,I33507,I33525,I33552,I33561,I33588,I33597,I33615,I33633,I33651,I33669,I33696,I33705,I33723,I33741,I33759,I33786,I33795,I33822,I33840,I33849,I33867,I33885,I33903,I33921,I33939,I33957,I33975,I33993,I34011,I34029,I34047,I34074,I34083,I34101,I34119,I34146,I34155,I34173,I34191,I34218,I34227,I34245,I34263,I34290,I34299,I34317,I34335,I34362,I34371,I34398,I34416,I34425,I34443,I34461,I34479,I34506,I34515,I34533,I34551,I34578,I34587,I34605,I34623,I34641,I34659,I34686,I34704,I34713,I34731,I34749,I34767,I34794,I34803,I34821,I34839,I34857,I34875,I34893,I34911,I34929,I34947,I34974,I34983,I35001,I35019,I35046,I35055,I35082,I35091,I35109,I35127,I35145,I35190,I35199,I35217,I35235,I35253,I35289,I35307,I35334,I35343,I35379,I35415,I35433,I35469,I35559,I35586,I35595,I35613,I35631,I35658,I35667,I35694,I35703,I35721,I35739,I35757,I35775,I35802,I35811,I35829,I35847,I35865,I35892,I35901,I35919,I35946,I35955,I35982,I35991,I36009,I36027,I36045,I36072,I36081,I36099,I36117,I36135,I36162,I36171,I36198,I36216,I36225,I36243,I36261,I36279,I36297,I36315,I36342,I36351,I36369,I36396,I36405,I36423,I36441,I36468,I36477,I36495,I36522,I36531,I36549,I36567,I36585,I36603,I36621,I36639,I36657,I36684,I36693,I36711,I36729,I36747,I36765,I36783,I36801,I36819,I36837,I36855,I36882,I36900,I36909,I36936,I36945,I36963,I36981,I36999,I37017,I37035,I37053,I37080,I37089,I37107,I37125,I37143,I37170,I37179,I37197,I37215,I37233,I37251,I37278,I37287,I37305,I37323,I37350,I37359,I37377,I37395,I37413,I37440,I37449,I37467,I37485,I37512,I37521,I37539,I37566,I37575,I37593,I37620,I37629,I37647,I37674,I37683,I37701,I37719,I37746,I37764,I37773,I37791,I37809,I37827,I37845,I37872,I37881,I37908,I37926,I37935,I37953,I37971,I37989,I38007,I38034,I38043,I38070,I38088,I38097,I38115,I38142,I38151,I38169,I38187,I38205,I38223,I38241,I38259,I38286,I38295,I38313,I38331,I38358,I38367,I38385,I38403,I38430,I38439,I38466,I38475,I38493,I38511,I38529,I38547,I38574,I38583,I38601,I38619,I38637,I38655,I38673,I38700,I38709,I38727,I38745,I38772,I38790,I38799,I38817,I38844,I38853,I38871,I38889,I38916,I38934,I38943,I38961,I38988,I39006,I39015,I39033,I39051,I39069,I39087,I39105,I39123,I39150,I39159,I39177,I39195,I39213,I39231,I39258,I39267,I39294,I39312,I39321,I39339,I39357,I39375,I39402,I39411,I39429,I39447,I39474,I39483,I39501,I39519,I39537,I39555,I39582,I39600,I39609,I39627,I39645,I39663,I39690,I39699,I39717,I39735,I39753,I39771,I39789,I39807,I39825,I39843,I39870,I39879,I39897,I39924,I39933,I39951,I39978,I39987,I40005,I40032,I40041,I40059,I40077,I40104,I40122,I40131,I40149,I40167,I40185,I40203,I40230,I40239,I40266,I40284,I40293,I40311,I40329,I40347,I40365,I40392,I40401,I40428,I40437,I40464,I40482,I40491,I40509,I40527,I40545,I40572,I40581,I40599,I40617,I40644,I40653,I40671,I40689,I40707,I40725,I40752,I40770,I40779,I40797,I40815,I40833,I40860,I40869,I40887,I40905,I40923,I40941,I40959,I40977,I40995,I41013,I41040,I41049,I41067,I41094,I41103,I41121,I41148,I41157,I41175,I41202,I41211,I41229,I41247,I41274,I41292,I41301,I41319,I41337,I41355,I41373,I41400,I41409,I41436,I41454,I41463,I41481,I41499,I41517,I41535,I41562,I41571,I41598,I41607,I41625,I41643,I41670,I41679,I41706,I41715,I41733,I41751,I41769,I41787,I41814,I41823,I41841,I41859,I41877,I41904,I41913,I41931,I41958,I41967,I41994,I42003,I42021,I42039,I42057,I42084,I42093,I42111,I42129,I42147,I42174,I42183,I42210,I42219,I42237,I42264,I42273,I42291,I42318,I42327,I42345,I42372,I42381,I42399,I42417,I42444,I42462,I42471,I42489,I42507,I42525,I42543,I42570,I42579,I42606,I42624,I42633,I42651,I42669,I42687,I42705,I42732,I42741,I42768,I42786,I42795,I42813,I42840,I42849,I42867,I42885,I42903,I42921,I42939,I42957,I42975,I43002,I43011,I43029,I43047,I43065,I43083,I43101,I43119,I43146,I43164,I43173,I43191,I43209,I43227,I43254,I43263,I43281,I43299,I43326,I43335,I43353,I43371,I43398,I43407,I43425,I43443,I43470,I43479,I43506,I43515,I43533,I43551,I43569,I43587,I43614,I43623,I43641,I43659,I43677,I43704,I43713,I43731,I43758,I43767,I43794,I43803,I43821,I43839,I43857,I43884,I43893,I43911,I43929,I43947,I43974,I43983,I44010,I44019,I44046,I44064,I44073,I44091,I44109,I44127,I44154,I44163,I44181,I44199,I44226,I44235,I44253,I44271,I44289,I44307,I44334,I44352,I44361,I44379,I44397,I44415,I44442,I44451,I44469,I44487,I44505,I44523,I44541,I44559,I44577,I44595,I44622,I44640,I44649,I44676,I44685,I44703,I44721,I44739,I44757,I44775,I44793,I44820,I44829,I44847,I44865,I44883,I44910,I44919,I44937,I44955,I44973,I44991,I45018,I45027,I45045,I45063,I45090,I45099,I45117,I45135,I45153,I45180,I45189,I45207,I45225,I45252,I45270,I45279,I45297,I45315,I45342,I45360,I45378,I45396,I45405,I45423,I45441,I45468,I45477,I45495,I45513,I45531,I45549,I45576,I45585,I45612,I45621,I45639,I45657,I45675,I45693,I45720,I45729,I45747,I45765,I45783,I45810,I45819,I45837,I45855,I45882,I45891,I45918,I45927,I45945,I45963,I45981,I45999,I46026,I46035,I46053,I46071,I46089,I46116,I46125,I46143,I46170,I46179,I46206,I46215,I46233,I46251,I46269,I46296,I46305,I46323,I46341,I46359,I46386,I46395,I46422,I46440,I46449,I46467,I46485,I46503,I46521,I46539,I46566,I46575,I46593,I46620,I46629,I46647,I46665,I46692,I46701,I46719,I46746,I46755,I46773,I46791,I46809,I46827,I46845,I46863,I46881,I46908,I46917,I46935,I46953,I46971,I46989,I47007,I47025,I47043,I47061,I47079,I47106,I47115,I47133,I47160,I47169,I47187,I47214,I47223,I47241,I47268,I47277,I47295,I47313,I47340,I47358,I47367,I47385,I47403,I47421,I47439,I47466,I47475,I47502,I47520,I47529,I47547,I47565,I47583,I47601,I47628,I47637,I47664,I47673,I47691,I47718,I47727,I47745,I47763,I47781,I47799,I47826,I47835,I47853,I47871,I47889,I47907,I47925,I47943,I47970,I47979,I47997,I48015,I48033,I48051,I48069,I48096,I48105,I48132,I48141,I48168,I48186,I48195,I48213,I48231,I48249,I48276,I48294,I48303,I48321,I48348,I48357,I48375,I48393,I48411,I48429,I48447,I48465,I48492,I48501,I48519,I48537,I48564,I48573,I48591,I48609,I48636,I48645,I48672,I48681,I48699,I48717,I48735,I48753,I48780,I48789,I48807,I48825,I48843,I48861,I48879,I48906,I48924,I48933,I48951,I48969,I48996,I49014,I49032,I49050,I49059,I49077,I49095,I49122,I49131,I49149,I49167,I49185,I49203,I49230,I49239,I49266,I49275,I49293,I49311,I49329,I49347,I49374,I49383,I49401,I49419,I49437,I49464,I49482,I49491,I49509,I49527,I49545,I49572,I49581,I49608,I49617,I49635,I49653,I49680,I49689,I49716,I49725,I49743,I49761,I49788,I49797,I49815,I49833,I49851,I49878,I49887,I49905,I49923,I49941,I49959,I49986,I50004,I50013,I50040,I50049,I50076,I50094,I50103,I50121,I50139,I50157,I50184,I50193,I50211,I50229,I50256,I50265,I50283,I50301,I50319,I50337,I50364,I50382,I50391,I50409,I50427,I50445,I50472,I50481,I50499,I50517,I50535,I50553,I50571,I50589,I50607,I50625,I50652,I50670,I50679,I50697,I50724,I50733,I50751,I50769,I50787,I50805,I50823,I50841,I50859,I50886,I50895,I50913,I50931,I50949,I50967,I50985,I51003,I51030,I51048,I51057,I51075,I51093,I51111,I51138,I51147,I51165,I51183,I51210,I51219,I51237,I51255,I51282,I51291,I51309,I51327,I51354,I51363,I51390,I51399,I51417,I51435,I51453,I51471,I51498,I51507,I51525,I51543,I51561,I51588,I51597,I51615,I51642,I51651,I51678,I51687,I51705,I51723,I51741,I51768,I51777,I51795,I51813,I51831,I51858,I51867,I51894,I51912,I51921,I51939,I51957,I51984,I52002,I52020,I52038,I52047,I52065,I52083,I52110,I52119,I52137,I52155,I52173,I52191,I52218,I52227,I52254,I52263,I52281,I52299,I52317,I52335,I52362,I52371,I52389,I52407,I52425,I52452,I52461,I52479,I52506,I52515,I52533,I52551,I52569,I52587,I52623,I52641,I52659,I52695,I52713,I52758,I52767,I52803,I52821,I52839,I52857,I52893,I52929,I52956,I52983,I53037,I53064,I53073,I53100,I53118,I53127,I53145,I53163,I53181,I53199,I53217,I53235,I53253,I53271,I53289,I53307,I53325,I53352,I53361,I53379,I53397,I53424,I53433,I53451,I53469,I53496,I53505,I53523,I53541,I53568,I53577,I53595,I53613,I53640,I53649,I53667,I53685,I53712,I53730,I53739,I53757,I53784,I53793,I53811,I53829,I53856,I53874,I53883,I53901,I53928,I53946,I53955,I53973,I53991,I54009,I54027,I54045,I54063,I54090,I54099,I54117,I54135,I54153,I54171,I54198,I54207,I54225,I54243,I54270,I54279,I54306,I54315,I54333,I54351,I54369,I54387,I54414,I54423,I54441,I54459,I54477,I54504,I54513,I54531,I54558,I54567,I54594,I54603,I54621,I54639,I54657,I54684,I54693,I54711,I54729,I54747,I54774,I54783,I54810,I54828,I54837,I54855,I54873,I54891,I54909,I54927,I54954,I54963,I54981,I55008,I55017,I55035,I55053,I55080,I55089,I55107,I55134,I55143,I55161,I55179,I55197,I55215,I55233,I55251,I55269,I55296,I55305,I55323,I55341,I55359,I55377,I55395,I55413,I55431,I55449,I55467,I55494,I55512,I55521,I55539,I55566,I55575,I55593,I55611,I55629,I55647,I55665,I55683,I55701,I55728,I55737,I55755,I55773,I55791,I55809,I55827,I55845,I55872,I55890,I55899,I55917,I55935,I55953,I55980,I55989,I56007,I56025,I56052,I56061,I56079,I56097,I56124,I56142,I56151,I56178,I56187,I56205,I56223,I56241,I56259,I56277,I56295,I56322,I56331,I56349,I56367,I56385,I56412,I56421,I56439,I56457,I56475,I56493,I56520,I56529,I56547,I56565,I56592,I56601,I56619,I56637,I56655,I56682,I56691,I56709,I56727,I56754,I56763,I56781,I56799,I56826,I56835,I56862,I56871,I56889,I56907,I56925,I56943,I56970,I56979,I56997,I57015,I57033,I57060,I57069,I57087,I57114,I57123,I57150,I57159,I57177,I57195,I57213,I57240,I57249,I57267,I57285,I57303,I57330,I57339,I57366,I57375,I57393,I57420,I57429,I57447,I57474,I57483,I57501,I57528,I57537,I57555,I57573,I57600,I57618,I57627,I57645,I57663,I57681,I57699,I57726,I57735,I57762,I57780,I57789,I57807,I57825,I57843,I57861,I57888,I57897,I57924,I57933,I57960,I57969,I57987,I58005,I58023,I58041,I58068,I58077,I58095,I58113,I58131,I58149,I58167,I58185,I58203,I58221,I58239,I58257,I58275,I58293,I58311,I58329,I58347,I58374,I58383,I58410,I58428,I58437,I58455,I58473,I58500,I58509,I58536,I58554,I58563,I58581,I58599,I58617,I58644,I58653,I58680,I58689,I58707,I58725,I58752,I58761,I58788,I58797,I58815,I58833,I58860,I58869,I58887,I58905,I58923,I58950,I58959,I58977,I58995,I59013,I59031,I59058,I59076,I59085,I59112,I59121,I59148,I59166,I59175,I59193,I59211,I59229,I59247,I59265,I59283,I59301,I59319,I59337,I59355,I59373,I59400,I59409,I59427,I59445,I59472,I59481,I59499,I59517,I59544,I59553,I59571,I59589,I59616,I59625,I59643,I59661,I59688,I59706,I59715,I59733,I59760,I59769,I59787,I59805,I59823,I59841,I59859,I59877,I59895,I59922,I59931,I59949,I59967,I59985,I60003,I60021,I60039,I60066,I60084,I60093,I60111,I60129,I60147,I60174,I60183,I60201,I60219,I60246,I60255,I60273,I60291,I60318,I60327,I60345,I60363,I60390,I60408,I60426,I60435,I60453,I60480,I60489,I60507,I60534,I60543,I60561,I60579,I60597,I60624,I60633,I60651,I60669,I60687,I60705,I60723,I60750,I60759,I60786,I60795,I60813,I60831,I60849,I60876,I60885,I60912,I60921,I60939,I60957,I60975,I60993,I61020,I61029,I61047,I61065,I61083,I61101,I61119,I61137,I61155,I61173,I61191,I61209,I61227,I61245,I61263,I61281,I61299,I61326,I61335,I61362,I61380,I61389,I61407,I61425,I61452,I61461,I61488,I61497,I61515,I61533,I61560,I61578,I61587,I61605,I61632,I61641,I61659,I61677,I61704,I61722,I61731,I61749,I61776,I61794,I61803,I61821,I61839,I61857,I61875,I61893,I61911,I61938,I61947,I61965,I61983,I62001,I62019,I62046,I62064,I62073,I62091,I62118,I62127,I62145,I62163,I62181,I62199,I62217,I62235,I62253,I62280,I62289,I62307,I62325,I62343,I62361,I62379,I62397,I62424,I62442,I62451,I62469,I62487,I62505,I62532,I62541,I62559,I62577,I62604,I62613,I62631,I62649,I62676,I62685,I62712,I62730,I62739,I62757,I62775,I62793,I62811,I62829,I62847,I62865,I62883,I62901,I62919,I62937,I62964,I62973,I62991,I63009,I63036,I63045,I63063,I63081,I63108,I63117,I63135,I63153,I63180,I63189,I63207,I63225,I63252,I63261,I63279,I63297,I63324,I63333,I63360,I63369,I63387,I63405,I63423,I63441,I63468,I63477,I63495,I63513,I63531,I63558,I63567,I63585,I63612,I63621,I63648,I63657,I63675,I63693,I63711,I63738,I63747,I63765,I63783,I63801,I63828,I63837,I63864,I63873,I63891,I63918,I63927,I63945,I63972,I63981,I63999,I64026,I64035,I64053,I64071,I64098,I64116,I64125,I64143,I64161,I64179,I64197,I64224,I64233,I64260,I64278,I64287,I64305,I64323,I64341,I64359,I64386,I64395,I64422,I64440,I64449,I64467,I64494,I64503,I64521,I64539,I64557,I64575,I64593,I64611,I64629,I64647,I64665,I64683,I64701,I64719,I64737,I64764,I64773,I64800,I64809,I64827,I64845,I64863,I64890,I64899,I64926,I64935,I64953,I64971,I64989,I65016,I65025,I65043,I65061,I65088,I65106,I65124,I65133,I65151,I65178,I65187,I65205,I65232,I65241,I65259,I65277,I65295,I65322,I65331,I65349,I65367,I65385,I65403,I65421,I65448,I65457,I65484,I65493,I65511,I65529,I65547,I65574,I65592,I65601,I65619,I65637,I65664,I65682,I65700,I65718,I65727,I65745,I65763,I65790,I65799,I65817,I65835,I65853,I65871,I65898,I65907,I65934,I65943,I65961,I65979,I65997,I66015,I66042,I66051,I66069,I66087,I66105,I66132,I66150,I66159,I66177,I66195,I66213,I66231,I66249,I66276,I66285,I66303,I66330,I66339,I66357,I66375,I66402,I66411,I66429,I66456,I66465,I66483,I66501,I66519,I66537,I66555,I66573,I66591,I66618,I66627,I66645,I66663,I66681,I66699,I66717,I66735,I66753,I66771,I66789,I66816,I66834,I66843,I66861,I66888,I66897,I66915,I66933,I66951,I66969,I66987,I67005,I67023,I67050,I67059,I67077,I67095,I67113,I67131,I67149,I67167,I67194,I67212,I67221,I67239,I67257,I67275,I67302,I67311,I67329,I67347,I67374,I67383,I67401,I67419,I67446,I67455,I67473,I67491,I67518,I67536,I67554,I67563,I67581,I67608,I67617,I67635,I67662,I67671,I67689,I67707,I67725,I67752,I67761,I67779,I67797,I67815,I67833,I67851,I67878,I67887,I67914,I67923,I67941,I67959,I67977,I68004,I68013,I68040,I68058,I68067,I68085,I68103,I68121,I68148,I68157,I68175,I68193,I68220,I68229,I68247,I68265,I68283,I68301,I68328,I68346,I68355,I68373,I68391,I68409,I68436,I68445,I68463,I68481,I68499,I68517,I68535,I68553,I68571,I68589,I68616,I68634,I68643,I68661,I68688,I68697,I68715,I68733,I68751,I68769,I68787,I68805,I68832,I68841,I68859,I68877,I68904,I68913,I68931,I68949,I68976,I68985,I69012,I69021,I69039,I69057,I69075,I69093,I69120,I69129,I69147,I69165,I69183,I69201,I69219,I69246,I69255,I69282,I69300,I69309,I69327,I69345,I69363,I69390,I69399,I69417,I69435,I69462,I69471,I69489,I69507,I69525,I69543,I69570,I69588,I69597,I69615,I69633,I69651,I69678,I69687,I69705,I69723,I69741,I69759,I69777,I69795,I69813,I69831,I69858,I69867,I69885,I69903,I69930,I69948,I69957,I69975,I70011,I70029,I70074,I70101,I70119,I70146,I70164,I70191,I70227,I70245,I70263,I70281,I70317,I70389,I70416,I70425,I70452,I70470,I70479,I70497,I70515,I70533,I70560,I70569,I70587,I70605,I70632,I70641,I70659,I70677,I70695,I70713,I70740,I70758,I70767,I70785,I70803,I70821,I70848,I70857,I70875,I70893,I70911,I70929,I70947,I70965,I70983,I71001,I71028,I71046,I71055,I71073,I71100,I71109,I71127,I71145,I71163,I71181,I71199,I71217,I71244,I71253,I71271,I71289,I71316,I71325,I71343,I71361,I71388,I71397,I71424,I71433,I71451,I71469,I71487,I71505,I71532,I71541,I71559,I71577,I71595,I71613,I71631,I71658,I71667,I71685,I71703,I71730,I71748,I71757,I71775,I71802,I71811,I71829,I71847,I71874,I71892,I71901,I71919,I71946,I71964,I71973,I71991,I72009,I72027,I72045,I72063,I72081,I72108,I72117,I72135,I72153,I72171,I72189,I72216,I72234,I72243,I72261,I72288,I72297,I72315,I72333,I72351,I72369,I72387,I72405,I72423,I72450,I72459,I72477,I72495,I72513,I72531,I72549,I72567,I72594,I72612,I72621,I72639,I72657,I72675,I72702,I72711,I72729,I72747,I72774,I72783,I72801,I72819,I72846,I72855,I72882,I72900,I72909,I72927,I72945,I72963,I72981,I72999,I73017,I73035,I73053,I73071,I73089,I73107,I73134,I73143,I73161,I73179,I73206,I73215,I73233,I73251,I73278,I73287,I73305,I73323,I73350,I73359,I73377,I73395,I73422,I73431,I73449,I73467,I73494,I73512,I73521,I73539,I73566,I73575,I73593,I73611,I73638,I73656,I73665,I73683,I73710,I73728,I73737,I73755,I73773,I73791,I73809,I73827,I73845,I73872,I73881,I73899,I73917,I73935,I73953,I73980,I73989,I74007,I74025,I74052,I74070,I74088,I74097,I74115,I74142,I74151,I74169,I74196,I74205,I74223,I74241,I74259,I74286,I74295,I74313,I74331,I74349,I74367,I74385,I74412,I74421,I74448,I74457,I74475,I74493,I74511,I74538,I74547,I74565,I74583,I74610,I74619,I74646,I74655,I74673,I74691,I74709,I74727,I74754,I74763,I74781,I74799,I74817,I74844,I74853,I74871,I74898,I74907,I74934,I74943,I74961,I74979,I74997,I75024,I75033,I75051,I75069,I75087,I75114,I75123,I75150,I75168,I75177,I75195,I75222,I75231,I75249,I75267,I75285,I75303,I75321,I75339,I75357,I75375,I75393,I75411,I75429,I75447,I75465,I75492,I75501,I75528,I75537,I75555,I75573,I75591,I75618,I75627,I75654,I75663,I75681,I75699,I75717,I75744,I75753,I75780,I75798,I75807,I75825,I75843,I75861,I75888,I75897,I75915,I75933,I75960,I75969,I75987,I76005,I76023,I76041,I76068,I76086,I76095,I76113,I76131,I76149,I76176,I76185,I76203,I76221,I76239,I76257,I76275,I76293,I76311,I76329,I76356,I76365,I76392,I76401,I76419,I76437,I76455,I76473,I76500,I76509,I76527,I76545,I76563,I76581,I76599,I76617,I76635,I76653,I76671,I76689,I76707,I76725,I76743,I76761,I76779,I76806,I76815,I76842,I76860,I76869,I76887,I76905,I76932,I76941,I76968,I76977,I76995,I77013,I77040,I77058,I77067,I77085,I77112,I77121,I77139,I77157,I77184,I77202,I77211,I77229,I77256,I77274,I77283,I77301,I77319,I77337,I77355,I77373,I77391,I77418,I77427,I77445,I77463,I77481,I77499,I77526,I77535,I77562,I77580,I77589,I77607,I77625,I77643,I77670,I77679,I77697,I77715,I77742,I77751,I77769,I77787,I77805,I77823,I77850,I77868,I77877,I77895,I77913,I77931,I77958,I77967,I77985,I78003,I78021,I78039,I78057,I78075,I78093,I78111,I78138,I78156,I78165,I78183,I78210,I78219,I78237,I78255,I78273,I78291,I78309,I78327,I78345,I78372,I78381,I78399,I78417,I78435,I78453,I78471,I78489,I78516,I78534,I78543,I78561,I78579,I78597,I78624,I78633,I78651,I78669,I78696,I78705,I78723,I78741,I78768,I78777,I78795,I78822,I78831,I78849,I78876,I78885,I78903,I78930,I78939,I78957,I78975,I79002,I79020,I79029,I79047,I79065,I79083,I79101,I79128,I79137,I79164,I79182,I79191,I79209,I79227,I79245,I79263,I79290,I79299,I79326,I79344,I79353,I79371,I79398,I79407,I79425,I79443,I79461,I79479,I79497,I79515,I79533,I79560,I79569,I79587,I79605,I79623,I79641,I79659,I79677,I79704,I79722,I79731,I79749,I79767,I79785,I79812,I79821,I79839,I79857,I79884,I79893,I79911,I79929,I79956,I79965,I79983,I80001,I80028,I80037,I80064,I80073,I80091,I80109,I80127,I80145,I80172,I80181,I80199,I80217,I80235,I80262,I80271,I80289,I80316,I80325,I80352,I80361,I80379,I80397,I80415,I80442,I80451,I80469,I80487,I80505,I80532,I80541,I80568,I80577,I80604,I80622,I80631,I80649,I80667,I80685,I80703,I80721,I80739,I80757,I80775,I80793,I80811,I80829,I80856,I80865,I80883,I80901,I80928,I80937,I80955,I80973,I81000,I81009,I81027,I81045,I81072,I81081,I81099,I81117,I81144,I81153,I81171,I81189,I81216,I81234,I81252,I81261,I81279,I81306,I81315,I81333,I81360,I81369,I81387,I81405,I81423,I81450,I81459,I81477,I81495,I81513,I81531,I81549,I81576,I81585,I81612,I81621,I81639,I81657,I81675,I81702,I81711,I81738,I81747,I81765,I81783,I81801,I81819,I81846,I81855,I81873,I81891,I81909,I81927,I81945,I81963,I81981,I81999,I82017,I82035,I82053,I82071,I82089,I82107,I82125,I82152,I82161,I82188,I82206,I82215,I82233,I82251,I82278,I82287,I82314,I82332,I82341,I82359,I82386,I82395,I82413,I82431,I82449,I82467,I82485,I82503,I82530,I82539,I82557,I82575,I82602,I82611,I82629,I82647,I82674,I82683,I82710,I82719,I82737,I82755,I82773,I82791,I82818,I82827,I82845,I82863,I82881,I82899,I82917,I82944,I82953,I82971,I82989,I83016,I83034,I83043,I83061,I83088,I83097,I83115,I83133,I83160,I83178,I83187,I83205,I83232,I83250,I83259,I83277,I83295,I83313,I83331,I83349,I83367,I83394,I83403,I83421,I83439,I83457,I83475,I83502,I83520,I83529,I83547,I83574,I83583,I83601,I83619,I83637,I83655,I83673,I83691,I83709,I83736,I83745,I83763,I83781,I83799,I83817,I83835,I83853,I83880,I83898,I83907,I83925,I83943,I83961,I83988,I83997,I84015,I84033,I84060,I84069,I84087,I84105,I84132,I84141,I84159,I84177,I84204,I84213,I84240,I84249,I84267,I84285,I84303,I84321,I84348,I84357,I84375,I84393,I84411,I84438,I84447,I84465,I84492,I84501,I84528,I84537,I84555,I84573,I84591,I84618,I84627,I84645,I84663,I84681,I84708,I84717,I84744,I84753,I84780,I84789,I84807,I84825,I84843,I84861,I84888,I84897,I84915,I84933,I84951,I84969,I84987,I85005,I85023,I85041,I85059,I85077,I85095,I85113,I85131,I85149,I85167,I85194,I85203,I85230,I85248,I85257,I85275,I85293,I85320,I85329,I85356,I85365,I85392,I85410,I85419,I85437,I85455,I85473,I85500,I85509,I85527,I85545,I85572,I85581,I85599,I85617,I85635,I85653,I85680,I85698,I85707,I85725,I85743,I85761,I85788,I85797,I85815,I85833,I85851,I85869,I85887,I85905,I85923,I85941,I85968,I85977,I85995,I86013,I86040,I86049,I86076,I86085,I86103,I86121,I86139,I86157,I86184,I86193,I86211,I86229,I86247,I86274,I86283,I86301,I86328,I86337,I86364,I86373,I86391,I86409,I86427,I86454,I86463,I86481,I86499,I86517,I86544,I86553,I86580,I86589,I86607,I86625,I86652,I86670,I86688,I86697,I86715,I86742,I86751,I86769,I86796,I86805,I86823,I86841,I86859,I86886,I86895,I86913,I86931,I86949,I86967,I86985,I87012,I87021,I87048,I87057,I87075,I87093,I87111,I87138,I87156,I87165,I87183,I87201,I87228,I87282,I87291,I87309,I87354,I87363,I87417,I87435,I87462,I87471,I87507,I87525,I87543,I87561,I87579,I87615;
not I_0 (I531,I522);
DFFARX1 I_1 (I108,I515,I531,I558,);
and I_2 (I567,I558,I140);
DFFARX1 I_3 (I567,I515,I531,I594,);
DFFARX1 I_4 (I148,I515,I531,I612,);
not I_5 (I621,I492);
not I_6 (I639,I340);
nand I_7 (I657,I639,I621);
nor I_8 (I675,I612,I657);
DFFARX1 I_9 (I657,I515,I531,I702,);
not I_10 (I711,I702);
not I_11 (I729,I316);
nand I_12 (I747,I639,I729);
DFFARX1 I_13 (I747,I515,I531,I774,);
not I_14 (I783,I774);
not I_15 (I801,I292);
nand I_16 (I819,I801,I156);
and I_17 (I837,I621,I819);
nor I_18 (I855,I747,I837);
DFFARX1 I_19 (I855,I515,I531,I882,);
DFFARX1 I_20 (I837,I515,I531,I900,);
nor I_21 (I909,I292,I300);
nor I_22 (I927,I747,I909);
or I_23 (I945,I292,I300);
nor I_24 (I963,I124,I188);
DFFARX1 I_25 (I963,I515,I531,I990,);
not I_26 (I999,I990);
nor I_27 (I1017,I999,I783);
nand I_28 (I1035,I999,I612);
not I_29 (I1053,I124);
nand I_30 (I1071,I1053,I729);
nand I_31 (I1089,I999,I1071);
nand I_32 (I1107,I1089,I1035);
nand I_33 (I1125,I1071,I945);
not I_34 (I1143,I522);
DFFARX1 I_35 (I675,I515,I1143,I1170,);
DFFARX1 I_36 (I594,I515,I1143,I1188,);
not I_37 (I1197,I1188);
nor I_38 (I1215,I1170,I1197);
DFFARX1 I_39 (I1197,I515,I1143,I1242,);
nor I_40 (I1251,I927,I1125);
and I_41 (I1269,I1251,I882);
nor I_42 (I1287,I1269,I927);
not I_43 (I1305,I927);
and I_44 (I1323,I1305,I1107);
nand I_45 (I1341,I1323,I882);
nor I_46 (I1359,I1305,I1341);
DFFARX1 I_47 (I1359,I515,I1143,I1386,);
not I_48 (I1395,I1341);
nand I_49 (I1413,I1197,I1395);
nand I_50 (I1431,I1269,I1395);
DFFARX1 I_51 (I1305,I515,I1143,I1458,);
not I_52 (I1467,I711);
nor I_53 (I1485,I1467,I1107);
nor I_54 (I1503,I1485,I1287);
DFFARX1 I_55 (I1503,I515,I1143,I1530,);
not I_56 (I1539,I1485);
DFFARX1 I_57 (I1539,I515,I1143,I1566,);
not I_58 (I1575,I1566);
nor I_59 (I1593,I1575,I1485);
nor I_60 (I1611,I1467,I1017);
and I_61 (I1629,I1611,I900);
or I_62 (I1647,I1629,I675);
DFFARX1 I_63 (I1647,I515,I1143,I1674,);
not I_64 (I1683,I1674);
nand I_65 (I1701,I1683,I1395);
not I_66 (I1719,I1701);
nand I_67 (I1737,I1701,I1413);
nand I_68 (I1755,I1683,I1269);
not I_69 (I1773,I522);
DFFARX1 I_70 (I1593,I515,I1773,I1800,);
nand I_71 (I1809,I1386,I1386);
and I_72 (I1827,I1809,I1458);
DFFARX1 I_73 (I1827,I515,I1773,I1854,);
nor I_74 (I1863,I1854,I1800);
not I_75 (I1881,I1854);
DFFARX1 I_76 (I1719,I515,I1773,I1908,);
nand I_77 (I1917,I1908,I1242);
not I_78 (I1935,I1917);
DFFARX1 I_79 (I1935,I515,I1773,I1962,);
not I_80 (I1971,I1962);
nor I_81 (I1989,I1800,I1917);
nor I_82 (I2007,I1854,I1989);
DFFARX1 I_83 (I1737,I515,I1773,I2034,);
DFFARX1 I_84 (I2034,I515,I1773,I2052,);
not I_85 (I2061,I2052);
not I_86 (I2079,I2034);
nand I_87 (I2097,I2079,I1881);
nand I_88 (I2115,I1755,I1215);
and I_89 (I2133,I2115,I1530);
DFFARX1 I_90 (I2133,I515,I1773,I2160,);
nor I_91 (I2169,I2160,I1800);
DFFARX1 I_92 (I2169,I515,I1773,I2196,);
DFFARX1 I_93 (I2160,I515,I1773,I2214,);
nor I_94 (I2223,I1431,I1215);
not I_95 (I2241,I2223);
nor I_96 (I2259,I2061,I2241);
nand I_97 (I2277,I2079,I2241);
nor I_98 (I2295,I1800,I2223);
DFFARX1 I_99 (I2223,I515,I1773,I2322,);
not I_100 (I2331,I522);
DFFARX1 I_101 (I2097,I515,I2331,I2358,);
nand I_102 (I2367,I2358,I2295);
DFFARX1 I_103 (I2007,I515,I2331,I2394,);
DFFARX1 I_104 (I2394,I515,I2331,I2412,);
not I_105 (I2421,I2412);
not I_106 (I2439,I2214);
nor I_107 (I2457,I2214,I1863);
not I_108 (I2475,I1971);
nand I_109 (I2493,I2439,I2475);
nor I_110 (I2511,I1971,I2214);
and I_111 (I2529,I2511,I2367);
not I_112 (I2547,I2277);
nand I_113 (I2565,I2547,I2322);
nor I_114 (I2583,I2277,I2196);
not I_115 (I2601,I2583);
nand I_116 (I2619,I2457,I2601);
DFFARX1 I_117 (I2583,I515,I2331,I2646,);
nor I_118 (I2655,I2259,I1971);
nor I_119 (I2673,I2655,I1863);
and I_120 (I2691,I2673,I2565);
DFFARX1 I_121 (I2691,I515,I2331,I2718,);
nor I_122 (I2727,I2655,I2493);
or I_123 (I2745,I2583,I2655);
nor I_124 (I2763,I2259,I2196);
DFFARX1 I_125 (I2763,I515,I2331,I2790,);
not I_126 (I2799,I2790);
nand I_127 (I2817,I2799,I2439);
nor I_128 (I2835,I2817,I1863);
DFFARX1 I_129 (I2835,I515,I2331,I2862,);
nor I_130 (I2871,I2799,I2493);
nor I_131 (I2889,I2655,I2871);
not I_132 (I2907,I522);
DFFARX1 I_133 (I2718,I515,I2907,I2934,);
DFFARX1 I_134 (I2421,I515,I2907,I2952,);
not I_135 (I2961,I2952);
not I_136 (I2979,I2646);
nor I_137 (I2997,I2979,I2862);
not I_138 (I3015,I2529);
nor I_139 (I3033,I2997,I2889);
nor I_140 (I3051,I2952,I3033);
DFFARX1 I_141 (I3051,I515,I2907,I3078,);
nor I_142 (I3087,I2889,I2862);
nand I_143 (I3105,I3087,I2646);
DFFARX1 I_144 (I3105,I515,I2907,I3132,);
nor I_145 (I3141,I3015,I2889);
nand I_146 (I3159,I3141,I2529);
nor I_147 (I3177,I2934,I3159);
DFFARX1 I_148 (I3177,I515,I2907,I3204,);
not I_149 (I3213,I3159);
nand I_150 (I3231,I2952,I3213);
DFFARX1 I_151 (I3159,I515,I2907,I3258,);
not I_152 (I3267,I3258);
not I_153 (I3285,I2889);
not I_154 (I3303,I2745);
nor I_155 (I3321,I3303,I2529);
nor I_156 (I3339,I3267,I3321);
nor I_157 (I3357,I3303,I2862);
and I_158 (I3375,I3357,I2619);
or I_159 (I3393,I3375,I2727);
DFFARX1 I_160 (I3393,I515,I2907,I3420,);
nor I_161 (I3429,I3420,I2934);
not I_162 (I3447,I3420);
and I_163 (I3465,I3447,I2934);
nor I_164 (I3483,I2961,I3465);
nand I_165 (I3501,I3447,I3015);
nor I_166 (I3519,I3303,I3501);
nand I_167 (I3537,I3447,I3213);
nand I_168 (I3555,I3015,I2745);
nor I_169 (I3573,I3285,I3555);
not I_170 (I3591,I522);
DFFARX1 I_171 (I3537,I515,I3591,I3618,);
and I_172 (I3627,I3618,I3204);
DFFARX1 I_173 (I3627,I515,I3591,I3654,);
DFFARX1 I_174 (I3573,I515,I3591,I3672,);
not I_175 (I3681,I3483);
not I_176 (I3699,I3078);
nand I_177 (I3717,I3699,I3681);
nor I_178 (I3735,I3672,I3717);
DFFARX1 I_179 (I3717,I515,I3591,I3762,);
not I_180 (I3771,I3762);
not I_181 (I3789,I3339);
nand I_182 (I3807,I3699,I3789);
DFFARX1 I_183 (I3807,I515,I3591,I3834,);
not I_184 (I3843,I3834);
not I_185 (I3861,I3519);
nand I_186 (I3879,I3861,I3132);
and I_187 (I3897,I3681,I3879);
nor I_188 (I3915,I3807,I3897);
DFFARX1 I_189 (I3915,I515,I3591,I3942,);
DFFARX1 I_190 (I3897,I515,I3591,I3960,);
nor I_191 (I3969,I3519,I3429);
nor I_192 (I3987,I3807,I3969);
or I_193 (I4005,I3519,I3429);
nor I_194 (I4023,I3204,I3231);
DFFARX1 I_195 (I4023,I515,I3591,I4050,);
not I_196 (I4059,I4050);
nor I_197 (I4077,I4059,I3843);
nand I_198 (I4095,I4059,I3672);
not I_199 (I4113,I3204);
nand I_200 (I4131,I4113,I3789);
nand I_201 (I4149,I4059,I4131);
nand I_202 (I4167,I4149,I4095);
nand I_203 (I4185,I4131,I4005);
not I_204 (I4203,I522);
DFFARX1 I_205 (I3735,I515,I4203,I4230,);
DFFARX1 I_206 (I4230,I515,I4203,I4248,);
not I_207 (I4257,I4248);
not I_208 (I4275,I4230);
nand I_209 (I4293,I3654,I3735);
and I_210 (I4311,I4293,I4185);
DFFARX1 I_211 (I4311,I515,I4203,I4338,);
not I_212 (I4347,I4338);
DFFARX1 I_213 (I3771,I515,I4203,I4374,);
and I_214 (I4383,I4374,I3942);
nand I_215 (I4401,I4374,I3942);
nand I_216 (I4419,I4347,I4401);
DFFARX1 I_217 (I4077,I515,I4203,I4446,);
nor I_218 (I4455,I4446,I4383);
DFFARX1 I_219 (I4455,I515,I4203,I4482,);
nor I_220 (I4491,I4446,I4338);
nand I_221 (I4509,I3987,I4167);
and I_222 (I4527,I4509,I3960);
DFFARX1 I_223 (I4527,I515,I4203,I4554,);
nor I_224 (I4563,I4554,I4446);
not I_225 (I4581,I4554);
nor I_226 (I4599,I4581,I4347);
nor I_227 (I4617,I4275,I4599);
DFFARX1 I_228 (I4617,I515,I4203,I4644,);
nor I_229 (I4653,I4581,I4446);
nor I_230 (I4671,I3942,I4167);
nor I_231 (I4689,I4671,I4653);
not I_232 (I4707,I4671);
nand I_233 (I4725,I4401,I4707);
DFFARX1 I_234 (I4671,I515,I4203,I4752,);
DFFARX1 I_235 (I4671,I515,I4203,I4770,);
not I_236 (I4779,I522);
DFFARX1 I_237 (I4482,I515,I4779,I4806,);
and I_238 (I4815,I4806,I4491);
DFFARX1 I_239 (I4815,I515,I4779,I4842,);
DFFARX1 I_240 (I4644,I515,I4779,I4860,);
not I_241 (I4869,I4725);
not I_242 (I4887,I4257);
nand I_243 (I4905,I4887,I4869);
nor I_244 (I4923,I4860,I4905);
DFFARX1 I_245 (I4905,I515,I4779,I4950,);
not I_246 (I4959,I4950);
not I_247 (I4977,I4563);
nand I_248 (I4995,I4887,I4977);
DFFARX1 I_249 (I4995,I515,I4779,I5022,);
not I_250 (I5031,I5022);
not I_251 (I5049,I4419);
nand I_252 (I5067,I5049,I4482);
and I_253 (I5085,I4869,I5067);
nor I_254 (I5103,I4995,I5085);
DFFARX1 I_255 (I5103,I515,I4779,I5130,);
DFFARX1 I_256 (I5085,I515,I4779,I5148,);
nor I_257 (I5157,I4419,I4689);
nor I_258 (I5175,I4995,I5157);
or I_259 (I5193,I4419,I4689);
nor I_260 (I5211,I4752,I4770);
DFFARX1 I_261 (I5211,I515,I4779,I5238,);
not I_262 (I5247,I5238);
nor I_263 (I5265,I5247,I5031);
nand I_264 (I5283,I5247,I4860);
not I_265 (I5301,I4752);
nand I_266 (I5319,I5301,I4977);
nand I_267 (I5337,I5247,I5319);
nand I_268 (I5355,I5337,I5283);
nand I_269 (I5373,I5319,I5193);
not I_270 (I5391,I522);
DFFARX1 I_271 (I5265,I515,I5391,I5418,);
not I_272 (I5427,I5418);
nand I_273 (I5445,I5130,I5175);
and I_274 (I5463,I5445,I4842);
DFFARX1 I_275 (I5463,I515,I5391,I5490,);
not I_276 (I5499,I5355);
DFFARX1 I_277 (I5373,I515,I5391,I5526,);
not I_278 (I5535,I5526);
nor I_279 (I5553,I5535,I5427);
and I_280 (I5571,I5553,I5355);
nor I_281 (I5589,I5535,I5499);
nor I_282 (I5607,I5490,I5589);
DFFARX1 I_283 (I4959,I515,I5391,I5634,);
nor I_284 (I5643,I5634,I5490);
not I_285 (I5661,I5643);
not I_286 (I5679,I5634);
nor I_287 (I5697,I5679,I5571);
DFFARX1 I_288 (I5697,I515,I5391,I5724,);
nand I_289 (I5733,I4923,I4923);
and I_290 (I5751,I5733,I5130);
DFFARX1 I_291 (I5751,I515,I5391,I5778,);
nor I_292 (I5787,I5778,I5634);
DFFARX1 I_293 (I5787,I515,I5391,I5814,);
nand I_294 (I5823,I5778,I5679);
nand I_295 (I5841,I5661,I5823);
not I_296 (I5859,I5778);
nor I_297 (I5877,I5859,I5571);
DFFARX1 I_298 (I5877,I515,I5391,I5904,);
nor I_299 (I5913,I5148,I4923);
or I_300 (I5931,I5634,I5913);
nor I_301 (I5949,I5778,I5913);
or I_302 (I5967,I5490,I5913);
DFFARX1 I_303 (I5913,I515,I5391,I5994,);
not I_304 (I6003,I522);
DFFARX1 I_305 (I5931,I515,I6003,I6030,);
not I_306 (I6039,I6030);
nand I_307 (I6057,I5949,I5904);
and I_308 (I6075,I6057,I5814);
DFFARX1 I_309 (I6075,I515,I6003,I6102,);
DFFARX1 I_310 (I5949,I515,I6003,I6120,);
and I_311 (I6129,I6120,I5967);
nor I_312 (I6147,I6102,I6129);
DFFARX1 I_313 (I6147,I515,I6003,I6174,);
nand I_314 (I6183,I6120,I5967);
nand I_315 (I6201,I6039,I6183);
not I_316 (I6219,I6201);
DFFARX1 I_317 (I5814,I515,I6003,I6246,);
DFFARX1 I_318 (I6246,I515,I6003,I6264,);
nand I_319 (I6273,I5724,I5841);
and I_320 (I6291,I6273,I5994);
DFFARX1 I_321 (I6291,I515,I6003,I6318,);
DFFARX1 I_322 (I6318,I515,I6003,I6336,);
not I_323 (I6345,I6336);
not I_324 (I6363,I6318);
nand I_325 (I6381,I6363,I6183);
nor I_326 (I6399,I5607,I5841);
not I_327 (I6417,I6399);
nor I_328 (I6435,I6363,I6417);
nor I_329 (I6453,I6039,I6435);
DFFARX1 I_330 (I6453,I515,I6003,I6480,);
nor I_331 (I6489,I6102,I6417);
nor I_332 (I6507,I6318,I6489);
nor I_333 (I6525,I6246,I6399);
nor I_334 (I6543,I6102,I6399);
not I_335 (I6561,I522);
DFFARX1 I_336 (I6507,I515,I6561,I6588,);
DFFARX1 I_337 (I6588,I515,I6561,I6606,);
not I_338 (I6615,I6606);
not I_339 (I6633,I6588);
nand I_340 (I6651,I6264,I6174);
and I_341 (I6669,I6651,I6543);
DFFARX1 I_342 (I6669,I515,I6561,I6696,);
not I_343 (I6705,I6696);
DFFARX1 I_344 (I6381,I515,I6561,I6732,);
and I_345 (I6741,I6732,I6543);
nand I_346 (I6759,I6732,I6543);
nand I_347 (I6777,I6705,I6759);
DFFARX1 I_348 (I6480,I515,I6561,I6804,);
nor I_349 (I6813,I6804,I6741);
DFFARX1 I_350 (I6813,I515,I6561,I6840,);
nor I_351 (I6849,I6804,I6696);
nand I_352 (I6867,I6174,I6525);
and I_353 (I6885,I6867,I6219);
DFFARX1 I_354 (I6885,I515,I6561,I6912,);
nor I_355 (I6921,I6912,I6804);
not I_356 (I6939,I6912);
nor I_357 (I6957,I6939,I6705);
nor I_358 (I6975,I6633,I6957);
DFFARX1 I_359 (I6975,I515,I6561,I7002,);
nor I_360 (I7011,I6939,I6804);
nor I_361 (I7029,I6345,I6525);
nor I_362 (I7047,I7029,I7011);
not I_363 (I7065,I7029);
nand I_364 (I7083,I6759,I7065);
DFFARX1 I_365 (I7029,I515,I6561,I7110,);
DFFARX1 I_366 (I7029,I515,I6561,I7128,);
not I_367 (I7137,I522);
DFFARX1 I_368 (I7047,I515,I7137,I7164,);
not I_369 (I7173,I7164);
nand I_370 (I7191,I6840,I7002);
and I_371 (I7209,I7191,I7128);
DFFARX1 I_372 (I7209,I515,I7137,I7236,);
not I_373 (I7245,I6849);
DFFARX1 I_374 (I6921,I515,I7137,I7272,);
not I_375 (I7281,I7272);
nor I_376 (I7299,I7281,I7173);
and I_377 (I7317,I7299,I6849);
nor I_378 (I7335,I7281,I7245);
nor I_379 (I7353,I7236,I7335);
DFFARX1 I_380 (I7083,I515,I7137,I7380,);
nor I_381 (I7389,I7380,I7236);
not I_382 (I7407,I7389);
not I_383 (I7425,I7380);
nor I_384 (I7443,I7425,I7317);
DFFARX1 I_385 (I7443,I515,I7137,I7470,);
nand I_386 (I7479,I6615,I7110);
and I_387 (I7497,I7479,I6777);
DFFARX1 I_388 (I7497,I515,I7137,I7524,);
nor I_389 (I7533,I7524,I7380);
DFFARX1 I_390 (I7533,I515,I7137,I7560,);
nand I_391 (I7569,I7524,I7425);
nand I_392 (I7587,I7407,I7569);
not I_393 (I7605,I7524);
nor I_394 (I7623,I7605,I7317);
DFFARX1 I_395 (I7623,I515,I7137,I7650,);
nor I_396 (I7659,I6840,I7110);
or I_397 (I7677,I7380,I7659);
nor I_398 (I7695,I7524,I7659);
or I_399 (I7713,I7236,I7659);
DFFARX1 I_400 (I7659,I515,I7137,I7740,);
not I_401 (I7749,I522);
DFFARX1 I_402 (I7695,I515,I7749,I7776,);
DFFARX1 I_403 (I7776,I515,I7749,I7794,);
not I_404 (I7803,I7794);
not I_405 (I7821,I7776);
nand I_406 (I7839,I7740,I7353);
and I_407 (I7857,I7839,I7695);
DFFARX1 I_408 (I7857,I515,I7749,I7884,);
not I_409 (I7893,I7884);
DFFARX1 I_410 (I7587,I515,I7749,I7920,);
and I_411 (I7929,I7920,I7713);
nand I_412 (I7947,I7920,I7713);
nand I_413 (I7965,I7893,I7947);
DFFARX1 I_414 (I7560,I515,I7749,I7992,);
nor I_415 (I8001,I7992,I7929);
DFFARX1 I_416 (I8001,I515,I7749,I8028,);
nor I_417 (I8037,I7992,I7884);
nand I_418 (I8055,I7560,I7677);
and I_419 (I8073,I8055,I7650);
DFFARX1 I_420 (I8073,I515,I7749,I8100,);
nor I_421 (I8109,I8100,I7992);
not I_422 (I8127,I8100);
nor I_423 (I8145,I8127,I7893);
nor I_424 (I8163,I7821,I8145);
DFFARX1 I_425 (I8163,I515,I7749,I8190,);
nor I_426 (I8199,I8127,I7992);
nor I_427 (I8217,I7470,I7677);
nor I_428 (I8235,I8217,I8199);
not I_429 (I8253,I8217);
nand I_430 (I8271,I7947,I8253);
DFFARX1 I_431 (I8217,I515,I7749,I8298,);
DFFARX1 I_432 (I8217,I515,I7749,I8316,);
not I_433 (I8325,I522);
DFFARX1 I_434 (I8271,I515,I8325,I8352,);
nand I_435 (I8361,I8298,I8109);
and I_436 (I8379,I8361,I7803);
DFFARX1 I_437 (I8379,I515,I8325,I8406,);
nor I_438 (I8415,I8406,I8352);
not I_439 (I8433,I8406);
DFFARX1 I_440 (I8190,I515,I8325,I8460,);
nand I_441 (I8469,I8460,I8028);
not I_442 (I8487,I8469);
DFFARX1 I_443 (I8487,I515,I8325,I8514,);
not I_444 (I8523,I8514);
nor I_445 (I8541,I8352,I8469);
nor I_446 (I8559,I8406,I8541);
DFFARX1 I_447 (I8037,I515,I8325,I8586,);
DFFARX1 I_448 (I8586,I515,I8325,I8604,);
not I_449 (I8613,I8604);
not I_450 (I8631,I8586);
nand I_451 (I8649,I8631,I8433);
nand I_452 (I8667,I8028,I7965);
and I_453 (I8685,I8667,I8235);
DFFARX1 I_454 (I8685,I515,I8325,I8712,);
nor I_455 (I8721,I8712,I8352);
DFFARX1 I_456 (I8721,I515,I8325,I8748,);
DFFARX1 I_457 (I8712,I515,I8325,I8766,);
nor I_458 (I8775,I8316,I7965);
not I_459 (I8793,I8775);
nor I_460 (I8811,I8613,I8793);
nand I_461 (I8829,I8631,I8793);
nor I_462 (I8847,I8352,I8775);
DFFARX1 I_463 (I8775,I515,I8325,I8874,);
not I_464 (I8883,I522);
DFFARX1 I_465 (I8874,I515,I8883,I8910,);
not I_466 (I8919,I8910);
nand I_467 (I8937,I8523,I8415);
and I_468 (I8955,I8937,I8748);
DFFARX1 I_469 (I8955,I515,I8883,I8982,);
not I_470 (I8991,I8829);
DFFARX1 I_471 (I8748,I515,I8883,I9018,);
not I_472 (I9027,I9018);
nor I_473 (I9045,I9027,I8919);
and I_474 (I9063,I9045,I8829);
nor I_475 (I9081,I9027,I8991);
nor I_476 (I9099,I8982,I9081);
DFFARX1 I_477 (I8559,I515,I8883,I9126,);
nor I_478 (I9135,I9126,I8982);
not I_479 (I9153,I9135);
not I_480 (I9171,I9126);
nor I_481 (I9189,I9171,I9063);
DFFARX1 I_482 (I9189,I515,I8883,I9216,);
nand I_483 (I9225,I8649,I8811);
and I_484 (I9243,I9225,I8766);
DFFARX1 I_485 (I9243,I515,I8883,I9270,);
nor I_486 (I9279,I9270,I9126);
DFFARX1 I_487 (I9279,I515,I8883,I9306,);
nand I_488 (I9315,I9270,I9171);
nand I_489 (I9333,I9153,I9315);
not I_490 (I9351,I9270);
nor I_491 (I9369,I9351,I9063);
DFFARX1 I_492 (I9369,I515,I8883,I9396,);
nor I_493 (I9405,I8847,I8811);
or I_494 (I9423,I9126,I9405);
nor I_495 (I9441,I9270,I9405);
or I_496 (I9459,I8982,I9405);
DFFARX1 I_497 (I9405,I515,I8883,I9486,);
not I_498 (I9495,I522);
DFFARX1 I_499 (I9423,I515,I9495,I9522,);
nand I_500 (I9531,I9441,I9216);
and I_501 (I9549,I9531,I9486);
DFFARX1 I_502 (I9549,I515,I9495,I9576,);
nor I_503 (I9585,I9576,I9522);
not I_504 (I9603,I9576);
DFFARX1 I_505 (I9333,I515,I9495,I9630,);
nand I_506 (I9639,I9630,I9441);
not I_507 (I9657,I9639);
DFFARX1 I_508 (I9657,I515,I9495,I9684,);
not I_509 (I9693,I9684);
nor I_510 (I9711,I9522,I9639);
nor I_511 (I9729,I9576,I9711);
DFFARX1 I_512 (I9459,I515,I9495,I9756,);
DFFARX1 I_513 (I9756,I515,I9495,I9774,);
not I_514 (I9783,I9774);
not I_515 (I9801,I9756);
nand I_516 (I9819,I9801,I9603);
nand I_517 (I9837,I9306,I9099);
and I_518 (I9855,I9837,I9306);
DFFARX1 I_519 (I9855,I515,I9495,I9882,);
nor I_520 (I9891,I9882,I9522);
DFFARX1 I_521 (I9891,I515,I9495,I9918,);
DFFARX1 I_522 (I9882,I515,I9495,I9936,);
nor I_523 (I9945,I9396,I9099);
not I_524 (I9963,I9945);
nor I_525 (I9981,I9783,I9963);
nand I_526 (I9999,I9801,I9963);
nor I_527 (I10017,I9522,I9945);
DFFARX1 I_528 (I9945,I515,I9495,I10044,);
not I_529 (I10053,I522);
DFFARX1 I_530 (I9918,I515,I10053,I10080,);
DFFARX1 I_531 (I10080,I515,I10053,I10098,);
not I_532 (I10107,I10098);
not I_533 (I10125,I10080);
DFFARX1 I_534 (I10017,I515,I10053,I10152,);
not I_535 (I10161,I10152);
and I_536 (I10179,I10125,I9819);
not I_537 (I10197,I9918);
nand I_538 (I10215,I10197,I9819);
not I_539 (I10233,I9729);
nor I_540 (I10251,I10233,I10044);
nand I_541 (I10269,I10251,I9981);
nor I_542 (I10287,I10269,I10215);
DFFARX1 I_543 (I10287,I515,I10053,I10314,);
not I_544 (I10323,I10269);
not I_545 (I10341,I10044);
nand I_546 (I10359,I10341,I9819);
nor I_547 (I10377,I10044,I9918);
nand I_548 (I10395,I10179,I10377);
nand I_549 (I10413,I10125,I10044);
nand I_550 (I10431,I10233,I9936);
DFFARX1 I_551 (I10431,I515,I10053,I10458,);
DFFARX1 I_552 (I10431,I515,I10053,I10476,);
not I_553 (I10485,I9936);
nor I_554 (I10503,I10485,I9999);
and I_555 (I10521,I10503,I9693);
or I_556 (I10539,I10521,I9585);
DFFARX1 I_557 (I10539,I515,I10053,I10566,);
nand I_558 (I10575,I10566,I10197);
nor I_559 (I10593,I10575,I10359);
nor I_560 (I10611,I10566,I10161);
DFFARX1 I_561 (I10566,I515,I10053,I10638,);
not I_562 (I10647,I10638);
nor I_563 (I10665,I10647,I10323);
not I_564 (I10683,I522);
DFFARX1 I_565 (I10593,I515,I10683,I10710,);
nand I_566 (I10719,I10710,I10107);
DFFARX1 I_567 (I10476,I515,I10683,I10746,);
DFFARX1 I_568 (I10746,I515,I10683,I10764,);
not I_569 (I10773,I10764);
not I_570 (I10791,I10314);
nor I_571 (I10809,I10314,I10413);
not I_572 (I10827,I10395);
nand I_573 (I10845,I10791,I10827);
nor I_574 (I10863,I10395,I10314);
and I_575 (I10881,I10863,I10719);
not I_576 (I10899,I10665);
nand I_577 (I10917,I10899,I10314);
nor I_578 (I10935,I10665,I10611);
not I_579 (I10953,I10935);
nand I_580 (I10971,I10809,I10953);
DFFARX1 I_581 (I10935,I515,I10683,I10998,);
nor I_582 (I11007,I10611,I10395);
nor I_583 (I11025,I11007,I10413);
and I_584 (I11043,I11025,I10917);
DFFARX1 I_585 (I11043,I515,I10683,I11070,);
nor I_586 (I11079,I11007,I10845);
or I_587 (I11097,I10935,I11007);
nor I_588 (I11115,I10611,I10458);
DFFARX1 I_589 (I11115,I515,I10683,I11142,);
not I_590 (I11151,I11142);
nand I_591 (I11169,I11151,I10791);
nor I_592 (I11187,I11169,I10413);
DFFARX1 I_593 (I11187,I515,I10683,I11214,);
nor I_594 (I11223,I11151,I10845);
nor I_595 (I11241,I11007,I11223);
not I_596 (I11259,I522);
DFFARX1 I_597 (I11214,I515,I11259,I11286,);
not I_598 (I11295,I11286);
nand I_599 (I11313,I10881,I11097);
and I_600 (I11331,I11313,I11079);
DFFARX1 I_601 (I11331,I515,I11259,I11358,);
not I_602 (I11367,I10773);
DFFARX1 I_603 (I10971,I515,I11259,I11394,);
not I_604 (I11403,I11394);
nor I_605 (I11421,I11403,I11295);
and I_606 (I11439,I11421,I10773);
nor I_607 (I11457,I11403,I11367);
nor I_608 (I11475,I11358,I11457);
DFFARX1 I_609 (I10881,I515,I11259,I11502,);
nor I_610 (I11511,I11502,I11358);
not I_611 (I11529,I11511);
not I_612 (I11547,I11502);
nor I_613 (I11565,I11547,I11439);
DFFARX1 I_614 (I11565,I515,I11259,I11592,);
nand I_615 (I11601,I10998,I11214);
and I_616 (I11619,I11601,I11070);
DFFARX1 I_617 (I11619,I515,I11259,I11646,);
nor I_618 (I11655,I11646,I11502);
DFFARX1 I_619 (I11655,I515,I11259,I11682,);
nand I_620 (I11691,I11646,I11547);
nand I_621 (I11709,I11529,I11691);
not I_622 (I11727,I11646);
nor I_623 (I11745,I11727,I11439);
DFFARX1 I_624 (I11745,I515,I11259,I11772,);
nor I_625 (I11781,I11241,I11214);
or I_626 (I11799,I11502,I11781);
nor I_627 (I11817,I11646,I11781);
or I_628 (I11835,I11358,I11781);
DFFARX1 I_629 (I11781,I515,I11259,I11862,);
not I_630 (I11871,I522);
DFFARX1 I_631 (I11817,I515,I11871,I11898,);
DFFARX1 I_632 (I11898,I515,I11871,I11916,);
not I_633 (I11925,I11916);
not I_634 (I11943,I11898);
DFFARX1 I_635 (I11475,I515,I11871,I11970,);
nand I_636 (I11979,I11970,I11862);
not I_637 (I11997,I11862);
not I_638 (I12015,I11835);
nand I_639 (I12033,I11709,I11682);
and I_640 (I12051,I11709,I11682);
not I_641 (I12069,I11592);
nand I_642 (I12087,I12069,I12015);
nor I_643 (I12105,I12087,I11979);
nor I_644 (I12123,I11997,I12087);
nand I_645 (I12141,I12051,I12123);
not I_646 (I12159,I11772);
nor I_647 (I12177,I12159,I11709);
nor I_648 (I12195,I12177,I11592);
nor I_649 (I12213,I11943,I12195);
DFFARX1 I_650 (I12213,I515,I11871,I12240,);
not I_651 (I12249,I12177);
DFFARX1 I_652 (I12249,I515,I11871,I12276,);
and I_653 (I12285,I11970,I12177);
nor I_654 (I12303,I12159,I11682);
and I_655 (I12321,I12303,I11799);
or I_656 (I12339,I12321,I11817);
DFFARX1 I_657 (I12339,I515,I11871,I12366,);
nor I_658 (I12375,I12366,I12069);
DFFARX1 I_659 (I12375,I515,I11871,I12402,);
nand I_660 (I12411,I12366,I11970);
nand I_661 (I12429,I12069,I12411);
nor I_662 (I12447,I12429,I12033);
not I_663 (I12465,I522);
DFFARX1 I_664 (I12285,I515,I12465,I12492,);
DFFARX1 I_665 (I12105,I515,I12465,I12510,);
not I_666 (I12519,I12510);
nor I_667 (I12537,I12492,I12519);
DFFARX1 I_668 (I12519,I515,I12465,I12564,);
nor I_669 (I12573,I12447,I12276);
and I_670 (I12591,I12573,I11925);
nor I_671 (I12609,I12591,I12447);
not I_672 (I12627,I12447);
and I_673 (I12645,I12627,I12402);
nand I_674 (I12663,I12645,I12141);
nor I_675 (I12681,I12627,I12663);
DFFARX1 I_676 (I12681,I515,I12465,I12708,);
not I_677 (I12717,I12663);
nand I_678 (I12735,I12519,I12717);
nand I_679 (I12753,I12591,I12717);
DFFARX1 I_680 (I12627,I515,I12465,I12780,);
not I_681 (I12789,I12240);
nor I_682 (I12807,I12789,I12402);
nor I_683 (I12825,I12807,I12609);
DFFARX1 I_684 (I12825,I515,I12465,I12852,);
not I_685 (I12861,I12807);
DFFARX1 I_686 (I12861,I515,I12465,I12888,);
not I_687 (I12897,I12888);
nor I_688 (I12915,I12897,I12807);
nor I_689 (I12933,I12789,I12402);
and I_690 (I12951,I12933,I12105);
or I_691 (I12969,I12951,I12141);
DFFARX1 I_692 (I12969,I515,I12465,I12996,);
not I_693 (I13005,I12996);
nand I_694 (I13023,I13005,I12717);
not I_695 (I13041,I13023);
nand I_696 (I13059,I13023,I12735);
nand I_697 (I13077,I13005,I12591);
not I_698 (I13095,I522);
DFFARX1 I_699 (I12780,I515,I13095,I13122,);
and I_700 (I13131,I13122,I13059);
DFFARX1 I_701 (I13131,I515,I13095,I13158,);
DFFARX1 I_702 (I12708,I515,I13095,I13176,);
not I_703 (I13185,I13041);
not I_704 (I13203,I12537);
nand I_705 (I13221,I13203,I13185);
nor I_706 (I13239,I13176,I13221);
DFFARX1 I_707 (I13221,I515,I13095,I13266,);
not I_708 (I13275,I13266);
not I_709 (I13293,I12753);
nand I_710 (I13311,I13203,I13293);
DFFARX1 I_711 (I13311,I515,I13095,I13338,);
not I_712 (I13347,I13338);
not I_713 (I13365,I12915);
nand I_714 (I13383,I13365,I12708);
and I_715 (I13401,I13185,I13383);
nor I_716 (I13419,I13311,I13401);
DFFARX1 I_717 (I13419,I515,I13095,I13446,);
DFFARX1 I_718 (I13401,I515,I13095,I13464,);
nor I_719 (I13473,I12915,I12852);
nor I_720 (I13491,I13311,I13473);
or I_721 (I13509,I12915,I12852);
nor I_722 (I13527,I12564,I13077);
DFFARX1 I_723 (I13527,I515,I13095,I13554,);
not I_724 (I13563,I13554);
nor I_725 (I13581,I13563,I13347);
nand I_726 (I13599,I13563,I13176);
not I_727 (I13617,I12564);
nand I_728 (I13635,I13617,I13293);
nand I_729 (I13653,I13563,I13635);
nand I_730 (I13671,I13653,I13599);
nand I_731 (I13689,I13635,I13509);
not I_732 (I13707,I522);
DFFARX1 I_733 (I13581,I515,I13707,I13734,);
not I_734 (I13743,I13734);
nand I_735 (I13761,I13446,I13491);
and I_736 (I13779,I13761,I13158);
DFFARX1 I_737 (I13779,I515,I13707,I13806,);
not I_738 (I13815,I13671);
DFFARX1 I_739 (I13689,I515,I13707,I13842,);
not I_740 (I13851,I13842);
nor I_741 (I13869,I13851,I13743);
and I_742 (I13887,I13869,I13671);
nor I_743 (I13905,I13851,I13815);
nor I_744 (I13923,I13806,I13905);
DFFARX1 I_745 (I13275,I515,I13707,I13950,);
nor I_746 (I13959,I13950,I13806);
not I_747 (I13977,I13959);
not I_748 (I13995,I13950);
nor I_749 (I14013,I13995,I13887);
DFFARX1 I_750 (I14013,I515,I13707,I14040,);
nand I_751 (I14049,I13239,I13239);
and I_752 (I14067,I14049,I13446);
DFFARX1 I_753 (I14067,I515,I13707,I14094,);
nor I_754 (I14103,I14094,I13950);
DFFARX1 I_755 (I14103,I515,I13707,I14130,);
nand I_756 (I14139,I14094,I13995);
nand I_757 (I14157,I13977,I14139);
not I_758 (I14175,I14094);
nor I_759 (I14193,I14175,I13887);
DFFARX1 I_760 (I14193,I515,I13707,I14220,);
nor I_761 (I14229,I13464,I13239);
or I_762 (I14247,I13950,I14229);
nor I_763 (I14265,I14094,I14229);
or I_764 (I14283,I13806,I14229);
DFFARX1 I_765 (I14229,I515,I13707,I14310,);
not I_766 (I14319,I522);
DFFARX1 I_767 (I14157,I515,I14319,I14346,);
DFFARX1 I_768 (I14346,I515,I14319,I14364,);
not I_769 (I14373,I14364);
DFFARX1 I_770 (I14265,I515,I14319,I14400,);
not I_771 (I14409,I14130);
nor I_772 (I14427,I14346,I14409);
not I_773 (I14445,I14247);
not I_774 (I14463,I13923);
nand I_775 (I14481,I14463,I14247);
nor I_776 (I14499,I14409,I14481);
nor I_777 (I14517,I14400,I14499);
DFFARX1 I_778 (I14463,I515,I14319,I14544,);
nor I_779 (I14553,I13923,I14310);
nand I_780 (I14571,I14553,I14040);
nor I_781 (I14589,I14571,I14445);
nand I_782 (I14607,I14589,I14130);
DFFARX1 I_783 (I14571,I515,I14319,I14634,);
nand I_784 (I14643,I14445,I13923);
nor I_785 (I14661,I14445,I13923);
nand I_786 (I14679,I14427,I14661);
not I_787 (I14697,I14283);
nor I_788 (I14715,I14697,I14643);
DFFARX1 I_789 (I14715,I515,I14319,I14742,);
nor I_790 (I14751,I14697,I14220);
and I_791 (I14769,I14751,I14130);
or I_792 (I14787,I14769,I14265);
DFFARX1 I_793 (I14787,I515,I14319,I14814,);
nor I_794 (I14823,I14814,I14400);
nor I_795 (I14841,I14346,I14823);
not I_796 (I14859,I14814);
nor I_797 (I14877,I14859,I14517);
DFFARX1 I_798 (I14877,I515,I14319,I14904,);
nand I_799 (I14913,I14859,I14445);
nor I_800 (I14931,I14697,I14913);
not I_801 (I14949,I522);
DFFARX1 I_802 (I14841,I515,I14949,I14976,);
DFFARX1 I_803 (I14976,I515,I14949,I14994,);
not I_804 (I15003,I14994);
nand I_805 (I15021,I14904,I14931);
and I_806 (I15039,I15021,I14742);
DFFARX1 I_807 (I15039,I515,I14949,I15066,);
DFFARX1 I_808 (I15066,I515,I14949,I15084,);
DFFARX1 I_809 (I15066,I515,I14949,I15102,);
DFFARX1 I_810 (I14679,I515,I14949,I15120,);
nand I_811 (I15129,I15120,I14607);
not I_812 (I15147,I15129);
nor I_813 (I15165,I14976,I15147);
DFFARX1 I_814 (I14373,I515,I14949,I15192,);
not I_815 (I15201,I15192);
nor I_816 (I15219,I15201,I15003);
nand I_817 (I15237,I15201,I15129);
nand I_818 (I15255,I14634,I14544);
and I_819 (I15273,I15255,I14931);
DFFARX1 I_820 (I15273,I515,I14949,I15300,);
nor I_821 (I15309,I15300,I14976);
DFFARX1 I_822 (I15309,I515,I14949,I15336,);
not I_823 (I15345,I15300);
nor I_824 (I15363,I14742,I14544);
not I_825 (I15381,I15363);
nor I_826 (I15399,I15129,I15381);
nor I_827 (I15417,I15345,I15399);
DFFARX1 I_828 (I15417,I515,I14949,I15444,);
nor I_829 (I15453,I15300,I15381);
nor I_830 (I15471,I15147,I15453);
nor I_831 (I15489,I15300,I15363);
not I_832 (I15507,I522);
DFFARX1 I_833 (I15336,I515,I15507,I15534,);
nand I_834 (I15543,I15102,I15489);
and I_835 (I15561,I15543,I15336);
DFFARX1 I_836 (I15561,I515,I15507,I15588,);
nor I_837 (I15597,I15588,I15534);
not I_838 (I15615,I15588);
DFFARX1 I_839 (I15237,I515,I15507,I15642,);
nand I_840 (I15651,I15642,I15084);
not I_841 (I15669,I15651);
DFFARX1 I_842 (I15669,I515,I15507,I15696,);
not I_843 (I15705,I15696);
nor I_844 (I15723,I15534,I15651);
nor I_845 (I15741,I15588,I15723);
DFFARX1 I_846 (I15471,I515,I15507,I15768,);
DFFARX1 I_847 (I15768,I515,I15507,I15786,);
not I_848 (I15795,I15786);
not I_849 (I15813,I15768);
nand I_850 (I15831,I15813,I15615);
nand I_851 (I15849,I15444,I15489);
and I_852 (I15867,I15849,I15165);
DFFARX1 I_853 (I15867,I515,I15507,I15894,);
nor I_854 (I15903,I15894,I15534);
DFFARX1 I_855 (I15903,I515,I15507,I15930,);
DFFARX1 I_856 (I15894,I515,I15507,I15948,);
nor I_857 (I15957,I15219,I15489);
not I_858 (I15975,I15957);
nor I_859 (I15993,I15795,I15975);
nand I_860 (I16011,I15813,I15975);
nor I_861 (I16029,I15534,I15957);
DFFARX1 I_862 (I15957,I515,I15507,I16056,);
not I_863 (I16065,I522);
DFFARX1 I_864 (I16011,I515,I16065,I16092,);
not I_865 (I16101,I16092);
DFFARX1 I_866 (I15993,I515,I16065,I16128,);
not I_867 (I16137,I16056);
nand I_868 (I16155,I16137,I15597);
not I_869 (I16173,I16155);
nor I_870 (I16191,I16173,I15705);
nor I_871 (I16209,I16101,I16191);
DFFARX1 I_872 (I16209,I515,I16065,I16236,);
not I_873 (I16245,I15705);
nand I_874 (I16263,I16245,I16173);
and I_875 (I16281,I16245,I15741);
nand I_876 (I16299,I16281,I15930);
nor I_877 (I16317,I16299,I16245);
and I_878 (I16335,I16128,I16299);
not I_879 (I16353,I16299);
nand I_880 (I16371,I16128,I16353);
nor I_881 (I16389,I16092,I16299);
not I_882 (I16407,I15930);
nor I_883 (I16425,I16407,I15741);
nand I_884 (I16443,I16425,I16245);
nor I_885 (I16461,I16155,I16443);
nor I_886 (I16479,I16407,I16029);
and I_887 (I16497,I16479,I15948);
or I_888 (I16515,I16497,I15831);
DFFARX1 I_889 (I16515,I515,I16065,I16542,);
nor I_890 (I16551,I16542,I16263);
DFFARX1 I_891 (I16551,I515,I16065,I16578,);
DFFARX1 I_892 (I16542,I515,I16065,I16596,);
not I_893 (I16605,I16542);
nor I_894 (I16623,I16605,I16128);
nor I_895 (I16641,I16425,I16623);
DFFARX1 I_896 (I16641,I515,I16065,I16668,);
not I_897 (I16677,I522);
DFFARX1 I_898 (I16578,I515,I16677,I16704,);
not I_899 (I16713,I16704);
nand I_900 (I16731,I16371,I16236);
and I_901 (I16749,I16731,I16596);
DFFARX1 I_902 (I16749,I515,I16677,I16776,);
not I_903 (I16785,I16668);
DFFARX1 I_904 (I16335,I515,I16677,I16812,);
not I_905 (I16821,I16812);
nor I_906 (I16839,I16821,I16713);
and I_907 (I16857,I16839,I16668);
nor I_908 (I16875,I16821,I16785);
nor I_909 (I16893,I16776,I16875);
DFFARX1 I_910 (I16317,I515,I16677,I16920,);
nor I_911 (I16929,I16920,I16776);
not I_912 (I16947,I16929);
not I_913 (I16965,I16920);
nor I_914 (I16983,I16965,I16857);
DFFARX1 I_915 (I16983,I515,I16677,I17010,);
nand I_916 (I17019,I16461,I16389);
and I_917 (I17037,I17019,I16578);
DFFARX1 I_918 (I17037,I515,I16677,I17064,);
nor I_919 (I17073,I17064,I16920);
DFFARX1 I_920 (I17073,I515,I16677,I17100,);
nand I_921 (I17109,I17064,I16965);
nand I_922 (I17127,I16947,I17109);
not I_923 (I17145,I17064);
nor I_924 (I17163,I17145,I16857);
DFFARX1 I_925 (I17163,I515,I16677,I17190,);
nor I_926 (I17199,I16389,I16389);
or I_927 (I17217,I16920,I17199);
nor I_928 (I17235,I17064,I17199);
or I_929 (I17253,I16776,I17199);
DFFARX1 I_930 (I17199,I515,I16677,I17280,);
not I_931 (I17289,I522);
DFFARX1 I_932 (I16893,I515,I17289,I17316,);
and I_933 (I17325,I17316,I17235);
DFFARX1 I_934 (I17325,I515,I17289,I17352,);
DFFARX1 I_935 (I17253,I515,I17289,I17370,);
not I_936 (I17379,I17100);
not I_937 (I17397,I17280);
nand I_938 (I17415,I17397,I17379);
nor I_939 (I17433,I17370,I17415);
DFFARX1 I_940 (I17415,I515,I17289,I17460,);
not I_941 (I17469,I17460);
not I_942 (I17487,I17217);
nand I_943 (I17505,I17397,I17487);
DFFARX1 I_944 (I17505,I515,I17289,I17532,);
not I_945 (I17541,I17532);
not I_946 (I17559,I17190);
nand I_947 (I17577,I17559,I17010);
and I_948 (I17595,I17379,I17577);
nor I_949 (I17613,I17505,I17595);
DFFARX1 I_950 (I17613,I515,I17289,I17640,);
DFFARX1 I_951 (I17595,I515,I17289,I17658,);
nor I_952 (I17667,I17190,I17127);
nor I_953 (I17685,I17505,I17667);
or I_954 (I17703,I17190,I17127);
nor I_955 (I17721,I17100,I17235);
DFFARX1 I_956 (I17721,I515,I17289,I17748,);
not I_957 (I17757,I17748);
nor I_958 (I17775,I17757,I17541);
nand I_959 (I17793,I17757,I17370);
not I_960 (I17811,I17100);
nand I_961 (I17829,I17811,I17487);
nand I_962 (I17847,I17757,I17829);
nand I_963 (I17865,I17847,I17793);
nand I_964 (I17883,I17829,I17703);
not I_965 (I17901,I522);
DFFARX1 I_966 (I348,I515,I17901,I17928,);
DFFARX1 I_967 (I17928,I515,I17901,I17946,);
not I_968 (I17955,I17946);
not I_969 (I17973,I17928);
nand I_970 (I17991,I252,I92);
and I_971 (I18009,I17991,I308);
DFFARX1 I_972 (I18009,I515,I17901,I18036,);
not I_973 (I18045,I18036);
DFFARX1 I_974 (I484,I515,I17901,I18072,);
and I_975 (I18081,I18072,I380);
nand I_976 (I18099,I18072,I380);
nand I_977 (I18117,I18045,I18099);
DFFARX1 I_978 (I76,I515,I17901,I18144,);
nor I_979 (I18153,I18144,I18081);
DFFARX1 I_980 (I18153,I515,I17901,I18180,);
nor I_981 (I18189,I18144,I18036);
nand I_982 (I18207,I460,I500);
and I_983 (I18225,I18207,I276);
DFFARX1 I_984 (I18225,I515,I17901,I18252,);
nor I_985 (I18261,I18252,I18144);
not I_986 (I18279,I18252);
nor I_987 (I18297,I18279,I18045);
nor I_988 (I18315,I17973,I18297);
DFFARX1 I_989 (I18315,I515,I17901,I18342,);
nor I_990 (I18351,I18279,I18144);
nor I_991 (I18369,I508,I500);
nor I_992 (I18387,I18369,I18351);
not I_993 (I18405,I18369);
nand I_994 (I18423,I18099,I18405);
DFFARX1 I_995 (I18369,I515,I17901,I18450,);
DFFARX1 I_996 (I18369,I515,I17901,I18468,);
not I_997 (I18477,I522);
DFFARX1 I_998 (I18342,I515,I18477,I18504,);
not I_999 (I18513,I18504);
nand I_1000 (I18531,I18423,I18261);
and I_1001 (I18549,I18531,I18450);
DFFARX1 I_1002 (I18549,I515,I18477,I18576,);
DFFARX1 I_1003 (I18117,I515,I18477,I18594,);
and I_1004 (I18603,I18594,I18180);
nor I_1005 (I18621,I18576,I18603);
DFFARX1 I_1006 (I18621,I515,I18477,I18648,);
nand I_1007 (I18657,I18594,I18180);
nand I_1008 (I18675,I18513,I18657);
not I_1009 (I18693,I18675);
DFFARX1 I_1010 (I18180,I515,I18477,I18720,);
DFFARX1 I_1011 (I18720,I515,I18477,I18738,);
nand I_1012 (I18747,I17955,I18387);
and I_1013 (I18765,I18747,I18189);
DFFARX1 I_1014 (I18765,I515,I18477,I18792,);
DFFARX1 I_1015 (I18792,I515,I18477,I18810,);
not I_1016 (I18819,I18810);
not I_1017 (I18837,I18792);
nand I_1018 (I18855,I18837,I18657);
nor I_1019 (I18873,I18468,I18387);
not I_1020 (I18891,I18873);
nor I_1021 (I18909,I18837,I18891);
nor I_1022 (I18927,I18513,I18909);
DFFARX1 I_1023 (I18927,I515,I18477,I18954,);
nor I_1024 (I18963,I18576,I18891);
nor I_1025 (I18981,I18792,I18963);
nor I_1026 (I18999,I18720,I18873);
nor I_1027 (I19017,I18576,I18873);
not I_1028 (I19035,I522);
DFFARX1 I_1029 (I18819,I515,I19035,I19062,);
and I_1030 (I19071,I19062,I18648);
DFFARX1 I_1031 (I19071,I515,I19035,I19098,);
DFFARX1 I_1032 (I18954,I515,I19035,I19116,);
not I_1033 (I19125,I18981);
not I_1034 (I19143,I19017);
nand I_1035 (I19161,I19143,I19125);
nor I_1036 (I19179,I19116,I19161);
DFFARX1 I_1037 (I19161,I515,I19035,I19206,);
not I_1038 (I19215,I19206);
not I_1039 (I19233,I18693);
nand I_1040 (I19251,I19143,I19233);
DFFARX1 I_1041 (I19251,I515,I19035,I19278,);
not I_1042 (I19287,I19278);
not I_1043 (I19305,I19017);
nand I_1044 (I19323,I19305,I18738);
and I_1045 (I19341,I19125,I19323);
nor I_1046 (I19359,I19251,I19341);
DFFARX1 I_1047 (I19359,I515,I19035,I19386,);
DFFARX1 I_1048 (I19341,I515,I19035,I19404,);
nor I_1049 (I19413,I19017,I18999);
nor I_1050 (I19431,I19251,I19413);
or I_1051 (I19449,I19017,I18999);
nor I_1052 (I19467,I18855,I18648);
DFFARX1 I_1053 (I19467,I515,I19035,I19494,);
not I_1054 (I19503,I19494);
nor I_1055 (I19521,I19503,I19287);
nand I_1056 (I19539,I19503,I19116);
not I_1057 (I19557,I18855);
nand I_1058 (I19575,I19557,I19233);
nand I_1059 (I19593,I19503,I19575);
nand I_1060 (I19611,I19593,I19539);
nand I_1061 (I19629,I19575,I19449);
not I_1062 (I19647,I522);
DFFARX1 I_1063 (I19521,I515,I19647,I19674,);
DFFARX1 I_1064 (I19674,I515,I19647,I19692,);
not I_1065 (I19701,I19692);
DFFARX1 I_1066 (I19386,I515,I19647,I19728,);
not I_1067 (I19737,I19629);
nor I_1068 (I19755,I19674,I19737);
not I_1069 (I19773,I19404);
not I_1070 (I19791,I19431);
nand I_1071 (I19809,I19791,I19404);
nor I_1072 (I19827,I19737,I19809);
nor I_1073 (I19845,I19728,I19827);
DFFARX1 I_1074 (I19791,I515,I19647,I19872,);
nor I_1075 (I19881,I19431,I19215);
nand I_1076 (I19899,I19881,I19179);
nor I_1077 (I19917,I19899,I19773);
nand I_1078 (I19935,I19917,I19629);
DFFARX1 I_1079 (I19899,I515,I19647,I19962,);
nand I_1080 (I19971,I19773,I19431);
nor I_1081 (I19989,I19773,I19431);
nand I_1082 (I20007,I19755,I19989);
not I_1083 (I20025,I19611);
nor I_1084 (I20043,I20025,I19971);
DFFARX1 I_1085 (I20043,I515,I19647,I20070,);
nor I_1086 (I20079,I20025,I19098);
and I_1087 (I20097,I20079,I19386);
or I_1088 (I20115,I20097,I19179);
DFFARX1 I_1089 (I20115,I515,I19647,I20142,);
nor I_1090 (I20151,I20142,I19728);
nor I_1091 (I20169,I19674,I20151);
not I_1092 (I20187,I20142);
nor I_1093 (I20205,I20187,I19845);
DFFARX1 I_1094 (I20205,I515,I19647,I20232,);
nand I_1095 (I20241,I20187,I19773);
nor I_1096 (I20259,I20025,I20241);
not I_1097 (I20277,I522);
DFFARX1 I_1098 (I20259,I515,I20277,I20304,);
nand I_1099 (I20313,I20259,I20232);
and I_1100 (I20331,I20313,I20070);
DFFARX1 I_1101 (I20331,I515,I20277,I20358,);
nor I_1102 (I20367,I20358,I20304);
not I_1103 (I20385,I20358);
DFFARX1 I_1104 (I19701,I515,I20277,I20412,);
nand I_1105 (I20421,I20412,I19872);
not I_1106 (I20439,I20421);
DFFARX1 I_1107 (I20439,I515,I20277,I20466,);
not I_1108 (I20475,I20466);
nor I_1109 (I20493,I20304,I20421);
nor I_1110 (I20511,I20358,I20493);
DFFARX1 I_1111 (I20007,I515,I20277,I20538,);
DFFARX1 I_1112 (I20538,I515,I20277,I20556,);
not I_1113 (I20565,I20556);
not I_1114 (I20583,I20538);
nand I_1115 (I20601,I20583,I20385);
nand I_1116 (I20619,I20070,I20169);
and I_1117 (I20637,I20619,I19962);
DFFARX1 I_1118 (I20637,I515,I20277,I20664,);
nor I_1119 (I20673,I20664,I20304);
DFFARX1 I_1120 (I20673,I515,I20277,I20700,);
DFFARX1 I_1121 (I20664,I515,I20277,I20718,);
nor I_1122 (I20727,I19935,I20169);
not I_1123 (I20745,I20727);
nor I_1124 (I20763,I20565,I20745);
nand I_1125 (I20781,I20583,I20745);
nor I_1126 (I20799,I20304,I20727);
DFFARX1 I_1127 (I20727,I515,I20277,I20826,);
not I_1128 (I20835,I522);
DFFARX1 I_1129 (I20700,I515,I20835,I20862,);
DFFARX1 I_1130 (I20781,I515,I20835,I20880,);
not I_1131 (I20889,I20880);
not I_1132 (I20907,I20475);
nor I_1133 (I20925,I20907,I20799);
not I_1134 (I20943,I20826);
nor I_1135 (I20961,I20925,I20511);
nor I_1136 (I20979,I20880,I20961);
DFFARX1 I_1137 (I20979,I515,I20835,I21006,);
nor I_1138 (I21015,I20511,I20799);
nand I_1139 (I21033,I21015,I20475);
DFFARX1 I_1140 (I21033,I515,I20835,I21060,);
nor I_1141 (I21069,I20943,I20511);
nand I_1142 (I21087,I21069,I20700);
nor I_1143 (I21105,I20862,I21087);
DFFARX1 I_1144 (I21105,I515,I20835,I21132,);
not I_1145 (I21141,I21087);
nand I_1146 (I21159,I20880,I21141);
DFFARX1 I_1147 (I21087,I515,I20835,I21186,);
not I_1148 (I21195,I21186);
not I_1149 (I21213,I20511);
not I_1150 (I21231,I20601);
nor I_1151 (I21249,I21231,I20826);
nor I_1152 (I21267,I21195,I21249);
nor I_1153 (I21285,I21231,I20763);
and I_1154 (I21303,I21285,I20367);
or I_1155 (I21321,I21303,I20718);
DFFARX1 I_1156 (I21321,I515,I20835,I21348,);
nor I_1157 (I21357,I21348,I20862);
not I_1158 (I21375,I21348);
and I_1159 (I21393,I21375,I20862);
nor I_1160 (I21411,I20889,I21393);
nand I_1161 (I21429,I21375,I20943);
nor I_1162 (I21447,I21231,I21429);
nand I_1163 (I21465,I21375,I21141);
nand I_1164 (I21483,I20943,I20601);
nor I_1165 (I21501,I21213,I21483);
not I_1166 (I21519,I522);
DFFARX1 I_1167 (I21060,I515,I21519,I21546,);
not I_1168 (I21555,I21546);
nand I_1169 (I21573,I21132,I21357);
and I_1170 (I21591,I21573,I21267);
DFFARX1 I_1171 (I21591,I515,I21519,I21618,);
not I_1172 (I21627,I21159);
DFFARX1 I_1173 (I21447,I515,I21519,I21654,);
not I_1174 (I21663,I21654);
nor I_1175 (I21681,I21663,I21555);
and I_1176 (I21699,I21681,I21159);
nor I_1177 (I21717,I21663,I21627);
nor I_1178 (I21735,I21618,I21717);
DFFARX1 I_1179 (I21132,I515,I21519,I21762,);
nor I_1180 (I21771,I21762,I21618);
not I_1181 (I21789,I21771);
not I_1182 (I21807,I21762);
nor I_1183 (I21825,I21807,I21699);
DFFARX1 I_1184 (I21825,I515,I21519,I21852,);
nand I_1185 (I21861,I21501,I21411);
and I_1186 (I21879,I21861,I21006);
DFFARX1 I_1187 (I21879,I515,I21519,I21906,);
nor I_1188 (I21915,I21906,I21762);
DFFARX1 I_1189 (I21915,I515,I21519,I21942,);
nand I_1190 (I21951,I21906,I21807);
nand I_1191 (I21969,I21789,I21951);
not I_1192 (I21987,I21906);
nor I_1193 (I22005,I21987,I21699);
DFFARX1 I_1194 (I22005,I515,I21519,I22032,);
nor I_1195 (I22041,I21465,I21411);
or I_1196 (I22059,I21762,I22041);
nor I_1197 (I22077,I21906,I22041);
or I_1198 (I22095,I21618,I22041);
DFFARX1 I_1199 (I22041,I515,I21519,I22122,);
not I_1200 (I22131,I522);
DFFARX1 I_1201 (I21735,I515,I22131,I22158,);
and I_1202 (I22167,I22158,I22077);
DFFARX1 I_1203 (I22167,I515,I22131,I22194,);
DFFARX1 I_1204 (I22095,I515,I22131,I22212,);
not I_1205 (I22221,I21942);
not I_1206 (I22239,I22122);
nand I_1207 (I22257,I22239,I22221);
nor I_1208 (I22275,I22212,I22257);
DFFARX1 I_1209 (I22257,I515,I22131,I22302,);
not I_1210 (I22311,I22302);
not I_1211 (I22329,I22059);
nand I_1212 (I22347,I22239,I22329);
DFFARX1 I_1213 (I22347,I515,I22131,I22374,);
not I_1214 (I22383,I22374);
not I_1215 (I22401,I22032);
nand I_1216 (I22419,I22401,I21852);
and I_1217 (I22437,I22221,I22419);
nor I_1218 (I22455,I22347,I22437);
DFFARX1 I_1219 (I22455,I515,I22131,I22482,);
DFFARX1 I_1220 (I22437,I515,I22131,I22500,);
nor I_1221 (I22509,I22032,I21969);
nor I_1222 (I22527,I22347,I22509);
or I_1223 (I22545,I22032,I21969);
nor I_1224 (I22563,I21942,I22077);
DFFARX1 I_1225 (I22563,I515,I22131,I22590,);
not I_1226 (I22599,I22590);
nor I_1227 (I22617,I22599,I22383);
nand I_1228 (I22635,I22599,I22212);
not I_1229 (I22653,I21942);
nand I_1230 (I22671,I22653,I22329);
nand I_1231 (I22689,I22599,I22671);
nand I_1232 (I22707,I22689,I22635);
nand I_1233 (I22725,I22671,I22545);
not I_1234 (I22743,I522);
DFFARX1 I_1235 (I22617,I515,I22743,I22770,);
nand I_1236 (I22779,I22770,I22275);
not I_1237 (I22797,I22779);
DFFARX1 I_1238 (I22725,I515,I22743,I22824,);
not I_1239 (I22833,I22824);
not I_1240 (I22851,I22500);
or I_1241 (I22869,I22311,I22500);
nor I_1242 (I22887,I22311,I22500);
or I_1243 (I22905,I22482,I22311);
DFFARX1 I_1244 (I22905,I515,I22743,I22932,);
not I_1245 (I22941,I22527);
nand I_1246 (I22959,I22941,I22194);
nand I_1247 (I22977,I22851,I22959);
and I_1248 (I22995,I22833,I22977);
nor I_1249 (I23013,I22527,I22707);
and I_1250 (I23031,I22833,I23013);
nor I_1251 (I23049,I22797,I23031);
DFFARX1 I_1252 (I23013,I515,I22743,I23076,);
not I_1253 (I23085,I23076);
nor I_1254 (I23103,I22833,I23085);
or I_1255 (I23121,I22905,I22482);
nor I_1256 (I23139,I22482,I22482);
nand I_1257 (I23157,I22977,I23139);
nand I_1258 (I23175,I23121,I23157);
DFFARX1 I_1259 (I23175,I515,I22743,I23202,);
nor I_1260 (I23211,I23139,I22869);
DFFARX1 I_1261 (I23211,I515,I22743,I23238,);
nor I_1262 (I23247,I22482,I22275);
DFFARX1 I_1263 (I23247,I515,I22743,I23274,);
DFFARX1 I_1264 (I23274,I515,I22743,I23292,);
not I_1265 (I23301,I23274);
nand I_1266 (I23319,I23301,I22779);
nand I_1267 (I23337,I23301,I22887);
not I_1268 (I23355,I522);
DFFARX1 I_1269 (I22932,I515,I23355,I23382,);
and I_1270 (I23391,I23382,I23337);
DFFARX1 I_1271 (I23391,I515,I23355,I23418,);
DFFARX1 I_1272 (I23292,I515,I23355,I23436,);
not I_1273 (I23445,I23238);
not I_1274 (I23463,I23319);
nand I_1275 (I23481,I23463,I23445);
nor I_1276 (I23499,I23436,I23481);
DFFARX1 I_1277 (I23481,I515,I23355,I23526,);
not I_1278 (I23535,I23526);
not I_1279 (I23553,I22995);
nand I_1280 (I23571,I23463,I23553);
DFFARX1 I_1281 (I23571,I515,I23355,I23598,);
not I_1282 (I23607,I23598);
not I_1283 (I23625,I23238);
nand I_1284 (I23643,I23625,I22995);
and I_1285 (I23661,I23445,I23643);
nor I_1286 (I23679,I23571,I23661);
DFFARX1 I_1287 (I23679,I515,I23355,I23706,);
DFFARX1 I_1288 (I23661,I515,I23355,I23724,);
nor I_1289 (I23733,I23238,I23202);
nor I_1290 (I23751,I23571,I23733);
or I_1291 (I23769,I23238,I23202);
nor I_1292 (I23787,I23049,I23103);
DFFARX1 I_1293 (I23787,I515,I23355,I23814,);
not I_1294 (I23823,I23814);
nor I_1295 (I23841,I23823,I23607);
nand I_1296 (I23859,I23823,I23436);
not I_1297 (I23877,I23049);
nand I_1298 (I23895,I23877,I23553);
nand I_1299 (I23913,I23823,I23895);
nand I_1300 (I23931,I23913,I23859);
nand I_1301 (I23949,I23895,I23769);
not I_1302 (I23967,I522);
DFFARX1 I_1303 (I23535,I515,I23967,I23994,);
DFFARX1 I_1304 (I23994,I515,I23967,I24012,);
not I_1305 (I24021,I24012);
nand I_1306 (I24039,I23751,I23499);
and I_1307 (I24057,I24039,I23706);
DFFARX1 I_1308 (I24057,I515,I23967,I24084,);
DFFARX1 I_1309 (I24084,I515,I23967,I24102,);
DFFARX1 I_1310 (I24084,I515,I23967,I24120,);
DFFARX1 I_1311 (I23949,I515,I23967,I24138,);
nand I_1312 (I24147,I24138,I23841);
not I_1313 (I24165,I24147);
nor I_1314 (I24183,I23994,I24165);
DFFARX1 I_1315 (I23418,I515,I23967,I24210,);
not I_1316 (I24219,I24210);
nor I_1317 (I24237,I24219,I24021);
nand I_1318 (I24255,I24219,I24147);
nand I_1319 (I24273,I23931,I23499);
and I_1320 (I24291,I24273,I23724);
DFFARX1 I_1321 (I24291,I515,I23967,I24318,);
nor I_1322 (I24327,I24318,I23994);
DFFARX1 I_1323 (I24327,I515,I23967,I24354,);
not I_1324 (I24363,I24318);
nor I_1325 (I24381,I23706,I23499);
not I_1326 (I24399,I24381);
nor I_1327 (I24417,I24147,I24399);
nor I_1328 (I24435,I24363,I24417);
DFFARX1 I_1329 (I24435,I515,I23967,I24462,);
nor I_1330 (I24471,I24318,I24399);
nor I_1331 (I24489,I24165,I24471);
nor I_1332 (I24507,I24318,I24381);
not I_1333 (I24525,I522);
DFFARX1 I_1334 (I24354,I515,I24525,I24552,);
and I_1335 (I24561,I24552,I24507);
DFFARX1 I_1336 (I24561,I515,I24525,I24588,);
DFFARX1 I_1337 (I24507,I515,I24525,I24606,);
not I_1338 (I24615,I24255);
not I_1339 (I24633,I24462);
nand I_1340 (I24651,I24633,I24615);
nor I_1341 (I24669,I24606,I24651);
DFFARX1 I_1342 (I24651,I515,I24525,I24696,);
not I_1343 (I24705,I24696);
not I_1344 (I24723,I24120);
nand I_1345 (I24741,I24633,I24723);
DFFARX1 I_1346 (I24741,I515,I24525,I24768,);
not I_1347 (I24777,I24768);
not I_1348 (I24795,I24237);
nand I_1349 (I24813,I24795,I24354);
and I_1350 (I24831,I24615,I24813);
nor I_1351 (I24849,I24741,I24831);
DFFARX1 I_1352 (I24849,I515,I24525,I24876,);
DFFARX1 I_1353 (I24831,I515,I24525,I24894,);
nor I_1354 (I24903,I24237,I24183);
nor I_1355 (I24921,I24741,I24903);
or I_1356 (I24939,I24237,I24183);
nor I_1357 (I24957,I24489,I24102);
DFFARX1 I_1358 (I24957,I515,I24525,I24984,);
not I_1359 (I24993,I24984);
nor I_1360 (I25011,I24993,I24777);
nand I_1361 (I25029,I24993,I24606);
not I_1362 (I25047,I24489);
nand I_1363 (I25065,I25047,I24723);
nand I_1364 (I25083,I24993,I25065);
nand I_1365 (I25101,I25083,I25029);
nand I_1366 (I25119,I25065,I24939);
not I_1367 (I25137,I522);
DFFARX1 I_1368 (I25011,I515,I25137,I25164,);
DFFARX1 I_1369 (I25164,I515,I25137,I25182,);
not I_1370 (I25191,I25182);
DFFARX1 I_1371 (I24876,I515,I25137,I25218,);
not I_1372 (I25227,I25119);
nor I_1373 (I25245,I25164,I25227);
not I_1374 (I25263,I24894);
not I_1375 (I25281,I24921);
nand I_1376 (I25299,I25281,I24894);
nor I_1377 (I25317,I25227,I25299);
nor I_1378 (I25335,I25218,I25317);
DFFARX1 I_1379 (I25281,I515,I25137,I25362,);
nor I_1380 (I25371,I24921,I24705);
nand I_1381 (I25389,I25371,I24669);
nor I_1382 (I25407,I25389,I25263);
nand I_1383 (I25425,I25407,I25119);
DFFARX1 I_1384 (I25389,I515,I25137,I25452,);
nand I_1385 (I25461,I25263,I24921);
nor I_1386 (I25479,I25263,I24921);
nand I_1387 (I25497,I25245,I25479);
not I_1388 (I25515,I25101);
nor I_1389 (I25533,I25515,I25461);
DFFARX1 I_1390 (I25533,I515,I25137,I25560,);
nor I_1391 (I25569,I25515,I24588);
and I_1392 (I25587,I25569,I24876);
or I_1393 (I25605,I25587,I24669);
DFFARX1 I_1394 (I25605,I515,I25137,I25632,);
nor I_1395 (I25641,I25632,I25218);
nor I_1396 (I25659,I25164,I25641);
not I_1397 (I25677,I25632);
nor I_1398 (I25695,I25677,I25335);
DFFARX1 I_1399 (I25695,I515,I25137,I25722,);
nand I_1400 (I25731,I25677,I25263);
nor I_1401 (I25749,I25515,I25731);
not I_1402 (I25767,I522);
DFFARX1 I_1403 (I25497,I515,I25767,I25794,);
DFFARX1 I_1404 (I25794,I515,I25767,I25812,);
not I_1405 (I25821,I25812);
not I_1406 (I25839,I25794);
DFFARX1 I_1407 (I25425,I515,I25767,I25866,);
not I_1408 (I25875,I25866);
and I_1409 (I25893,I25839,I25362);
not I_1410 (I25911,I25452);
nand I_1411 (I25929,I25911,I25362);
not I_1412 (I25947,I25659);
nor I_1413 (I25965,I25947,I25560);
nand I_1414 (I25983,I25965,I25749);
nor I_1415 (I26001,I25983,I25929);
DFFARX1 I_1416 (I26001,I515,I25767,I26028,);
not I_1417 (I26037,I25983);
not I_1418 (I26055,I25560);
nand I_1419 (I26073,I26055,I25362);
nor I_1420 (I26091,I25560,I25452);
nand I_1421 (I26109,I25893,I26091);
nand I_1422 (I26127,I25839,I25560);
nand I_1423 (I26145,I25947,I25191);
DFFARX1 I_1424 (I26145,I515,I25767,I26172,);
DFFARX1 I_1425 (I26145,I515,I25767,I26190,);
not I_1426 (I26199,I25191);
nor I_1427 (I26217,I26199,I25722);
and I_1428 (I26235,I26217,I25560);
or I_1429 (I26253,I26235,I25749);
DFFARX1 I_1430 (I26253,I515,I25767,I26280,);
nand I_1431 (I26289,I26280,I25911);
nor I_1432 (I26307,I26289,I26073);
nor I_1433 (I26325,I26280,I25875);
DFFARX1 I_1434 (I26280,I515,I25767,I26352,);
not I_1435 (I26361,I26352);
nor I_1436 (I26379,I26361,I26037);
not I_1437 (I26397,I522);
DFFARX1 I_1438 (I26028,I515,I26397,I26424,);
and I_1439 (I26433,I26424,I26325);
DFFARX1 I_1440 (I26433,I515,I26397,I26460,);
DFFARX1 I_1441 (I26325,I515,I26397,I26478,);
not I_1442 (I26487,I26379);
not I_1443 (I26505,I25821);
nand I_1444 (I26523,I26505,I26487);
nor I_1445 (I26541,I26478,I26523);
DFFARX1 I_1446 (I26523,I515,I26397,I26568,);
not I_1447 (I26577,I26568);
not I_1448 (I26595,I26109);
nand I_1449 (I26613,I26505,I26595);
DFFARX1 I_1450 (I26613,I515,I26397,I26640,);
not I_1451 (I26649,I26640);
not I_1452 (I26667,I26307);
nand I_1453 (I26685,I26667,I26127);
and I_1454 (I26703,I26487,I26685);
nor I_1455 (I26721,I26613,I26703);
DFFARX1 I_1456 (I26721,I515,I26397,I26748,);
DFFARX1 I_1457 (I26703,I515,I26397,I26766,);
nor I_1458 (I26775,I26307,I26028);
nor I_1459 (I26793,I26613,I26775);
or I_1460 (I26811,I26307,I26028);
nor I_1461 (I26829,I26190,I26172);
DFFARX1 I_1462 (I26829,I515,I26397,I26856,);
not I_1463 (I26865,I26856);
nor I_1464 (I26883,I26865,I26649);
nand I_1465 (I26901,I26865,I26478);
not I_1466 (I26919,I26190);
nand I_1467 (I26937,I26919,I26595);
nand I_1468 (I26955,I26865,I26937);
nand I_1469 (I26973,I26955,I26901);
nand I_1470 (I26991,I26937,I26811);
not I_1471 (I27009,I522);
DFFARX1 I_1472 (I26883,I515,I27009,I27036,);
not I_1473 (I27045,I27036);
nand I_1474 (I27063,I26748,I26793);
and I_1475 (I27081,I27063,I26460);
DFFARX1 I_1476 (I27081,I515,I27009,I27108,);
not I_1477 (I27117,I26973);
DFFARX1 I_1478 (I26991,I515,I27009,I27144,);
not I_1479 (I27153,I27144);
nor I_1480 (I27171,I27153,I27045);
and I_1481 (I27189,I27171,I26973);
nor I_1482 (I27207,I27153,I27117);
nor I_1483 (I27225,I27108,I27207);
DFFARX1 I_1484 (I26577,I515,I27009,I27252,);
nor I_1485 (I27261,I27252,I27108);
not I_1486 (I27279,I27261);
not I_1487 (I27297,I27252);
nor I_1488 (I27315,I27297,I27189);
DFFARX1 I_1489 (I27315,I515,I27009,I27342,);
nand I_1490 (I27351,I26541,I26541);
and I_1491 (I27369,I27351,I26748);
DFFARX1 I_1492 (I27369,I515,I27009,I27396,);
nor I_1493 (I27405,I27396,I27252);
DFFARX1 I_1494 (I27405,I515,I27009,I27432,);
nand I_1495 (I27441,I27396,I27297);
nand I_1496 (I27459,I27279,I27441);
not I_1497 (I27477,I27396);
nor I_1498 (I27495,I27477,I27189);
DFFARX1 I_1499 (I27495,I515,I27009,I27522,);
nor I_1500 (I27531,I26766,I26541);
or I_1501 (I27549,I27252,I27531);
nor I_1502 (I27567,I27396,I27531);
or I_1503 (I27585,I27108,I27531);
DFFARX1 I_1504 (I27531,I515,I27009,I27612,);
not I_1505 (I27621,I522);
DFFARX1 I_1506 (I27432,I515,I27621,I27648,);
not I_1507 (I27657,I27648);
DFFARX1 I_1508 (I27549,I515,I27621,I27684,);
not I_1509 (I27693,I27567);
nand I_1510 (I27711,I27693,I27585);
not I_1511 (I27729,I27711);
nor I_1512 (I27747,I27729,I27459);
nor I_1513 (I27765,I27657,I27747);
DFFARX1 I_1514 (I27765,I515,I27621,I27792,);
not I_1515 (I27801,I27459);
nand I_1516 (I27819,I27801,I27729);
and I_1517 (I27837,I27801,I27567);
nand I_1518 (I27855,I27837,I27225);
nor I_1519 (I27873,I27855,I27801);
and I_1520 (I27891,I27684,I27855);
not I_1521 (I27909,I27855);
nand I_1522 (I27927,I27684,I27909);
nor I_1523 (I27945,I27648,I27855);
not I_1524 (I27963,I27522);
nor I_1525 (I27981,I27963,I27567);
nand I_1526 (I27999,I27981,I27801);
nor I_1527 (I28017,I27711,I27999);
nor I_1528 (I28035,I27963,I27432);
and I_1529 (I28053,I28035,I27342);
or I_1530 (I28071,I28053,I27612);
DFFARX1 I_1531 (I28071,I515,I27621,I28098,);
nor I_1532 (I28107,I28098,I27819);
DFFARX1 I_1533 (I28107,I515,I27621,I28134,);
DFFARX1 I_1534 (I28098,I515,I27621,I28152,);
not I_1535 (I28161,I28098);
nor I_1536 (I28179,I28161,I27684);
nor I_1537 (I28197,I27981,I28179);
DFFARX1 I_1538 (I28197,I515,I27621,I28224,);
not I_1539 (I28233,I522);
DFFARX1 I_1540 (I27873,I515,I28233,I28260,);
nand I_1541 (I28269,I28134,I27945);
and I_1542 (I28287,I28269,I27792);
DFFARX1 I_1543 (I28287,I515,I28233,I28314,);
nor I_1544 (I28323,I28314,I28260);
not I_1545 (I28341,I28314);
DFFARX1 I_1546 (I28017,I515,I28233,I28368,);
nand I_1547 (I28377,I28368,I27945);
not I_1548 (I28395,I28377);
DFFARX1 I_1549 (I28395,I515,I28233,I28422,);
not I_1550 (I28431,I28422);
nor I_1551 (I28449,I28260,I28377);
nor I_1552 (I28467,I28314,I28449);
DFFARX1 I_1553 (I27927,I515,I28233,I28494,);
DFFARX1 I_1554 (I28494,I515,I28233,I28512,);
not I_1555 (I28521,I28512);
not I_1556 (I28539,I28494);
nand I_1557 (I28557,I28539,I28341);
nand I_1558 (I28575,I28152,I28134);
and I_1559 (I28593,I28575,I28224);
DFFARX1 I_1560 (I28593,I515,I28233,I28620,);
nor I_1561 (I28629,I28620,I28260);
DFFARX1 I_1562 (I28629,I515,I28233,I28656,);
DFFARX1 I_1563 (I28620,I515,I28233,I28674,);
nor I_1564 (I28683,I27891,I28134);
not I_1565 (I28701,I28683);
nor I_1566 (I28719,I28521,I28701);
nand I_1567 (I28737,I28539,I28701);
nor I_1568 (I28755,I28260,I28683);
DFFARX1 I_1569 (I28683,I515,I28233,I28782,);
not I_1570 (I28791,I522);
DFFARX1 I_1571 (I28656,I515,I28791,I28818,);
DFFARX1 I_1572 (I28737,I515,I28791,I28836,);
not I_1573 (I28845,I28836);
not I_1574 (I28863,I28431);
nor I_1575 (I28881,I28863,I28755);
not I_1576 (I28899,I28782);
nor I_1577 (I28917,I28881,I28467);
nor I_1578 (I28935,I28836,I28917);
DFFARX1 I_1579 (I28935,I515,I28791,I28962,);
nor I_1580 (I28971,I28467,I28755);
nand I_1581 (I28989,I28971,I28431);
DFFARX1 I_1582 (I28989,I515,I28791,I29016,);
nor I_1583 (I29025,I28899,I28467);
nand I_1584 (I29043,I29025,I28656);
nor I_1585 (I29061,I28818,I29043);
DFFARX1 I_1586 (I29061,I515,I28791,I29088,);
not I_1587 (I29097,I29043);
nand I_1588 (I29115,I28836,I29097);
DFFARX1 I_1589 (I29043,I515,I28791,I29142,);
not I_1590 (I29151,I29142);
not I_1591 (I29169,I28467);
not I_1592 (I29187,I28557);
nor I_1593 (I29205,I29187,I28782);
nor I_1594 (I29223,I29151,I29205);
nor I_1595 (I29241,I29187,I28719);
and I_1596 (I29259,I29241,I28323);
or I_1597 (I29277,I29259,I28674);
DFFARX1 I_1598 (I29277,I515,I28791,I29304,);
nor I_1599 (I29313,I29304,I28818);
not I_1600 (I29331,I29304);
and I_1601 (I29349,I29331,I28818);
nor I_1602 (I29367,I28845,I29349);
nand I_1603 (I29385,I29331,I28899);
nor I_1604 (I29403,I29187,I29385);
nand I_1605 (I29421,I29331,I29097);
nand I_1606 (I29439,I28899,I28557);
nor I_1607 (I29457,I29169,I29439);
not I_1608 (I29475,I522);
DFFARX1 I_1609 (I29421,I515,I29475,I29502,);
and I_1610 (I29511,I29502,I29088);
DFFARX1 I_1611 (I29511,I515,I29475,I29538,);
DFFARX1 I_1612 (I29457,I515,I29475,I29556,);
not I_1613 (I29565,I29367);
not I_1614 (I29583,I28962);
nand I_1615 (I29601,I29583,I29565);
nor I_1616 (I29619,I29556,I29601);
DFFARX1 I_1617 (I29601,I515,I29475,I29646,);
not I_1618 (I29655,I29646);
not I_1619 (I29673,I29223);
nand I_1620 (I29691,I29583,I29673);
DFFARX1 I_1621 (I29691,I515,I29475,I29718,);
not I_1622 (I29727,I29718);
not I_1623 (I29745,I29403);
nand I_1624 (I29763,I29745,I29016);
and I_1625 (I29781,I29565,I29763);
nor I_1626 (I29799,I29691,I29781);
DFFARX1 I_1627 (I29799,I515,I29475,I29826,);
DFFARX1 I_1628 (I29781,I515,I29475,I29844,);
nor I_1629 (I29853,I29403,I29313);
nor I_1630 (I29871,I29691,I29853);
or I_1631 (I29889,I29403,I29313);
nor I_1632 (I29907,I29088,I29115);
DFFARX1 I_1633 (I29907,I515,I29475,I29934,);
not I_1634 (I29943,I29934);
nor I_1635 (I29961,I29943,I29727);
nand I_1636 (I29979,I29943,I29556);
not I_1637 (I29997,I29088);
nand I_1638 (I30015,I29997,I29673);
nand I_1639 (I30033,I29943,I30015);
nand I_1640 (I30051,I30033,I29979);
nand I_1641 (I30069,I30015,I29889);
not I_1642 (I30087,I522);
DFFARX1 I_1643 (I29961,I515,I30087,I30114,);
DFFARX1 I_1644 (I30114,I515,I30087,I30132,);
not I_1645 (I30141,I30132);
DFFARX1 I_1646 (I29826,I515,I30087,I30168,);
not I_1647 (I30177,I30069);
nor I_1648 (I30195,I30114,I30177);
not I_1649 (I30213,I29844);
not I_1650 (I30231,I29871);
nand I_1651 (I30249,I30231,I29844);
nor I_1652 (I30267,I30177,I30249);
nor I_1653 (I30285,I30168,I30267);
DFFARX1 I_1654 (I30231,I515,I30087,I30312,);
nor I_1655 (I30321,I29871,I29655);
nand I_1656 (I30339,I30321,I29619);
nor I_1657 (I30357,I30339,I30213);
nand I_1658 (I30375,I30357,I30069);
DFFARX1 I_1659 (I30339,I515,I30087,I30402,);
nand I_1660 (I30411,I30213,I29871);
nor I_1661 (I30429,I30213,I29871);
nand I_1662 (I30447,I30195,I30429);
not I_1663 (I30465,I30051);
nor I_1664 (I30483,I30465,I30411);
DFFARX1 I_1665 (I30483,I515,I30087,I30510,);
nor I_1666 (I30519,I30465,I29538);
and I_1667 (I30537,I30519,I29826);
or I_1668 (I30555,I30537,I29619);
DFFARX1 I_1669 (I30555,I515,I30087,I30582,);
nor I_1670 (I30591,I30582,I30168);
nor I_1671 (I30609,I30114,I30591);
not I_1672 (I30627,I30582);
nor I_1673 (I30645,I30627,I30285);
DFFARX1 I_1674 (I30645,I515,I30087,I30672,);
nand I_1675 (I30681,I30627,I30213);
nor I_1676 (I30699,I30465,I30681);
not I_1677 (I30717,I522);
DFFARX1 I_1678 (I30699,I515,I30717,I30744,);
and I_1679 (I30753,I30744,I30402);
DFFARX1 I_1680 (I30753,I515,I30717,I30780,);
DFFARX1 I_1681 (I30609,I515,I30717,I30798,);
not I_1682 (I30807,I30699);
not I_1683 (I30825,I30312);
nand I_1684 (I30843,I30825,I30807);
nor I_1685 (I30861,I30798,I30843);
DFFARX1 I_1686 (I30843,I515,I30717,I30888,);
not I_1687 (I30897,I30888);
not I_1688 (I30915,I30447);
nand I_1689 (I30933,I30825,I30915);
DFFARX1 I_1690 (I30933,I515,I30717,I30960,);
not I_1691 (I30969,I30960);
not I_1692 (I30987,I30141);
nand I_1693 (I31005,I30987,I30510);
and I_1694 (I31023,I30807,I31005);
nor I_1695 (I31041,I30933,I31023);
DFFARX1 I_1696 (I31041,I515,I30717,I31068,);
DFFARX1 I_1697 (I31023,I515,I30717,I31086,);
nor I_1698 (I31095,I30141,I30510);
nor I_1699 (I31113,I30933,I31095);
or I_1700 (I31131,I30141,I30510);
nor I_1701 (I31149,I30375,I30672);
DFFARX1 I_1702 (I31149,I515,I30717,I31176,);
not I_1703 (I31185,I31176);
nor I_1704 (I31203,I31185,I30969);
nand I_1705 (I31221,I31185,I30798);
not I_1706 (I31239,I30375);
nand I_1707 (I31257,I31239,I30915);
nand I_1708 (I31275,I31185,I31257);
nand I_1709 (I31293,I31275,I31221);
nand I_1710 (I31311,I31257,I31131);
not I_1711 (I31329,I522);
DFFARX1 I_1712 (I30897,I515,I31329,I31356,);
nand I_1713 (I31365,I31356,I30861);
DFFARX1 I_1714 (I31068,I515,I31329,I31392,);
DFFARX1 I_1715 (I31392,I515,I31329,I31410,);
not I_1716 (I31419,I31410);
not I_1717 (I31437,I31113);
nor I_1718 (I31455,I31113,I31086);
not I_1719 (I31473,I31293);
nand I_1720 (I31491,I31437,I31473);
nor I_1721 (I31509,I31293,I31113);
and I_1722 (I31527,I31509,I31365);
not I_1723 (I31545,I31203);
nand I_1724 (I31563,I31545,I30780);
nor I_1725 (I31581,I31203,I31068);
not I_1726 (I31599,I31581);
nand I_1727 (I31617,I31455,I31599);
DFFARX1 I_1728 (I31581,I515,I31329,I31644,);
nor I_1729 (I31653,I30861,I31293);
nor I_1730 (I31671,I31653,I31086);
and I_1731 (I31689,I31671,I31563);
DFFARX1 I_1732 (I31689,I515,I31329,I31716,);
nor I_1733 (I31725,I31653,I31491);
or I_1734 (I31743,I31581,I31653);
nor I_1735 (I31761,I30861,I31311);
DFFARX1 I_1736 (I31761,I515,I31329,I31788,);
not I_1737 (I31797,I31788);
nand I_1738 (I31815,I31797,I31437);
nor I_1739 (I31833,I31815,I31086);
DFFARX1 I_1740 (I31833,I515,I31329,I31860,);
nor I_1741 (I31869,I31797,I31491);
nor I_1742 (I31887,I31653,I31869);
not I_1743 (I31905,I522);
DFFARX1 I_1744 (I31644,I515,I31905,I31932,);
and I_1745 (I31941,I31932,I31725);
DFFARX1 I_1746 (I31941,I515,I31905,I31968,);
DFFARX1 I_1747 (I31860,I515,I31905,I31986,);
not I_1748 (I31995,I31617);
not I_1749 (I32013,I31716);
nand I_1750 (I32031,I32013,I31995);
nor I_1751 (I32049,I31986,I32031);
DFFARX1 I_1752 (I32031,I515,I31905,I32076,);
not I_1753 (I32085,I32076);
not I_1754 (I32103,I31860);
nand I_1755 (I32121,I32013,I32103);
DFFARX1 I_1756 (I32121,I515,I31905,I32148,);
not I_1757 (I32157,I32148);
not I_1758 (I32175,I31419);
nand I_1759 (I32193,I32175,I31743);
and I_1760 (I32211,I31995,I32193);
nor I_1761 (I32229,I32121,I32211);
DFFARX1 I_1762 (I32229,I515,I31905,I32256,);
DFFARX1 I_1763 (I32211,I515,I31905,I32274,);
nor I_1764 (I32283,I31419,I31527);
nor I_1765 (I32301,I32121,I32283);
or I_1766 (I32319,I31419,I31527);
nor I_1767 (I32337,I31887,I31527);
DFFARX1 I_1768 (I32337,I515,I31905,I32364,);
not I_1769 (I32373,I32364);
nor I_1770 (I32391,I32373,I32157);
nand I_1771 (I32409,I32373,I31986);
not I_1772 (I32427,I31887);
nand I_1773 (I32445,I32427,I32103);
nand I_1774 (I32463,I32373,I32445);
nand I_1775 (I32481,I32463,I32409);
nand I_1776 (I32499,I32445,I32319);
not I_1777 (I32517,I522);
DFFARX1 I_1778 (I32391,I515,I32517,I32544,);
DFFARX1 I_1779 (I32256,I515,I32517,I32562,);
not I_1780 (I32571,I32562);
not I_1781 (I32589,I32481);
nor I_1782 (I32607,I32589,I32274);
not I_1783 (I32625,I32049);
nor I_1784 (I32643,I32607,I32301);
nor I_1785 (I32661,I32562,I32643);
DFFARX1 I_1786 (I32661,I515,I32517,I32688,);
nor I_1787 (I32697,I32301,I32274);
nand I_1788 (I32715,I32697,I32481);
DFFARX1 I_1789 (I32715,I515,I32517,I32742,);
nor I_1790 (I32751,I32625,I32301);
nand I_1791 (I32769,I32751,I32085);
nor I_1792 (I32787,I32544,I32769);
DFFARX1 I_1793 (I32787,I515,I32517,I32814,);
not I_1794 (I32823,I32769);
nand I_1795 (I32841,I32562,I32823);
DFFARX1 I_1796 (I32769,I515,I32517,I32868,);
not I_1797 (I32877,I32868);
not I_1798 (I32895,I32301);
not I_1799 (I32913,I32256);
nor I_1800 (I32931,I32913,I32049);
nor I_1801 (I32949,I32877,I32931);
nor I_1802 (I32967,I32913,I32499);
and I_1803 (I32985,I32967,I31968);
or I_1804 (I33003,I32985,I32049);
DFFARX1 I_1805 (I33003,I515,I32517,I33030,);
nor I_1806 (I33039,I33030,I32544);
not I_1807 (I33057,I33030);
and I_1808 (I33075,I33057,I32544);
nor I_1809 (I33093,I32571,I33075);
nand I_1810 (I33111,I33057,I32625);
nor I_1811 (I33129,I32913,I33111);
nand I_1812 (I33147,I33057,I32823);
nand I_1813 (I33165,I32625,I32256);
nor I_1814 (I33183,I32895,I33165);
not I_1815 (I33201,I522);
DFFARX1 I_1816 (I32742,I515,I33201,I33228,);
DFFARX1 I_1817 (I33228,I515,I33201,I33246,);
not I_1818 (I33255,I33246);
nand I_1819 (I33273,I32814,I32949);
and I_1820 (I33291,I33273,I32841);
DFFARX1 I_1821 (I33291,I515,I33201,I33318,);
DFFARX1 I_1822 (I33318,I515,I33201,I33336,);
DFFARX1 I_1823 (I33318,I515,I33201,I33354,);
DFFARX1 I_1824 (I33183,I515,I33201,I33372,);
nand I_1825 (I33381,I33372,I33129);
not I_1826 (I33399,I33381);
nor I_1827 (I33417,I33228,I33399);
DFFARX1 I_1828 (I32688,I515,I33201,I33444,);
not I_1829 (I33453,I33444);
nor I_1830 (I33471,I33453,I33255);
nand I_1831 (I33489,I33453,I33381);
nand I_1832 (I33507,I33147,I33093);
and I_1833 (I33525,I33507,I32814);
DFFARX1 I_1834 (I33525,I515,I33201,I33552,);
nor I_1835 (I33561,I33552,I33228);
DFFARX1 I_1836 (I33561,I515,I33201,I33588,);
not I_1837 (I33597,I33552);
nor I_1838 (I33615,I33039,I33093);
not I_1839 (I33633,I33615);
nor I_1840 (I33651,I33381,I33633);
nor I_1841 (I33669,I33597,I33651);
DFFARX1 I_1842 (I33669,I515,I33201,I33696,);
nor I_1843 (I33705,I33552,I33633);
nor I_1844 (I33723,I33399,I33705);
nor I_1845 (I33741,I33552,I33615);
not I_1846 (I33759,I522);
DFFARX1 I_1847 (I33723,I515,I33759,I33786,);
nand I_1848 (I33795,I33786,I33741);
DFFARX1 I_1849 (I33354,I515,I33759,I33822,);
DFFARX1 I_1850 (I33822,I515,I33759,I33840,);
not I_1851 (I33849,I33840);
not I_1852 (I33867,I33417);
nor I_1853 (I33885,I33417,I33696);
not I_1854 (I33903,I33588);
nand I_1855 (I33921,I33867,I33903);
nor I_1856 (I33939,I33588,I33417);
and I_1857 (I33957,I33939,I33795);
not I_1858 (I33975,I33471);
nand I_1859 (I33993,I33975,I33489);
nor I_1860 (I34011,I33471,I33588);
not I_1861 (I34029,I34011);
nand I_1862 (I34047,I33885,I34029);
DFFARX1 I_1863 (I34011,I515,I33759,I34074,);
nor I_1864 (I34083,I33741,I33588);
nor I_1865 (I34101,I34083,I33696);
and I_1866 (I34119,I34101,I33993);
DFFARX1 I_1867 (I34119,I515,I33759,I34146,);
nor I_1868 (I34155,I34083,I33921);
or I_1869 (I34173,I34011,I34083);
nor I_1870 (I34191,I33741,I33336);
DFFARX1 I_1871 (I34191,I515,I33759,I34218,);
not I_1872 (I34227,I34218);
nand I_1873 (I34245,I34227,I33867);
nor I_1874 (I34263,I34245,I33696);
DFFARX1 I_1875 (I34263,I515,I33759,I34290,);
nor I_1876 (I34299,I34227,I33921);
nor I_1877 (I34317,I34083,I34299);
not I_1878 (I34335,I522);
DFFARX1 I_1879 (I34074,I515,I34335,I34362,);
and I_1880 (I34371,I34362,I34155);
DFFARX1 I_1881 (I34371,I515,I34335,I34398,);
DFFARX1 I_1882 (I34290,I515,I34335,I34416,);
not I_1883 (I34425,I34047);
not I_1884 (I34443,I34146);
nand I_1885 (I34461,I34443,I34425);
nor I_1886 (I34479,I34416,I34461);
DFFARX1 I_1887 (I34461,I515,I34335,I34506,);
not I_1888 (I34515,I34506);
not I_1889 (I34533,I34290);
nand I_1890 (I34551,I34443,I34533);
DFFARX1 I_1891 (I34551,I515,I34335,I34578,);
not I_1892 (I34587,I34578);
not I_1893 (I34605,I33849);
nand I_1894 (I34623,I34605,I34173);
and I_1895 (I34641,I34425,I34623);
nor I_1896 (I34659,I34551,I34641);
DFFARX1 I_1897 (I34659,I515,I34335,I34686,);
DFFARX1 I_1898 (I34641,I515,I34335,I34704,);
nor I_1899 (I34713,I33849,I33957);
nor I_1900 (I34731,I34551,I34713);
or I_1901 (I34749,I33849,I33957);
nor I_1902 (I34767,I34317,I33957);
DFFARX1 I_1903 (I34767,I515,I34335,I34794,);
not I_1904 (I34803,I34794);
nor I_1905 (I34821,I34803,I34587);
nand I_1906 (I34839,I34803,I34416);
not I_1907 (I34857,I34317);
nand I_1908 (I34875,I34857,I34533);
nand I_1909 (I34893,I34803,I34875);
nand I_1910 (I34911,I34893,I34839);
nand I_1911 (I34929,I34875,I34749);
not I_1912 (I34947,I522);
DFFARX1 I_1913 (I34821,I515,I34947,I34974,);
not I_1914 (I34983,I34974);
nand I_1915 (I35001,I34686,I34731);
and I_1916 (I35019,I35001,I34398);
DFFARX1 I_1917 (I35019,I515,I34947,I35046,);
not I_1918 (I35055,I34911);
DFFARX1 I_1919 (I34929,I515,I34947,I35082,);
not I_1920 (I35091,I35082);
nor I_1921 (I35109,I35091,I34983);
and I_1922 (I35127,I35109,I34911);
nor I_1923 (I35145,I35091,I35055);
nor I_1924 (I35163,I35046,I35145);
DFFARX1 I_1925 (I34515,I515,I34947,I35190,);
nor I_1926 (I35199,I35190,I35046);
not I_1927 (I35217,I35199);
not I_1928 (I35235,I35190);
nor I_1929 (I35253,I35235,I35127);
DFFARX1 I_1930 (I35253,I515,I34947,I35280,);
nand I_1931 (I35289,I34479,I34479);
and I_1932 (I35307,I35289,I34686);
DFFARX1 I_1933 (I35307,I515,I34947,I35334,);
nor I_1934 (I35343,I35334,I35190);
DFFARX1 I_1935 (I35343,I515,I34947,I35370,);
nand I_1936 (I35379,I35334,I35235);
nand I_1937 (I35397,I35217,I35379);
not I_1938 (I35415,I35334);
nor I_1939 (I35433,I35415,I35127);
DFFARX1 I_1940 (I35433,I515,I34947,I35460,);
nor I_1941 (I35469,I34704,I34479);
or I_1942 (I35487,I35190,I35469);
nor I_1943 (I35505,I35334,I35469);
or I_1944 (I35523,I35046,I35469);
DFFARX1 I_1945 (I35469,I515,I34947,I35550,);
not I_1946 (I35559,I522);
DFFARX1 I_1947 (I396,I515,I35559,I35586,);
not I_1948 (I35595,I35586);
nand I_1949 (I35613,I356,I412);
and I_1950 (I35631,I35613,I468);
DFFARX1 I_1951 (I35631,I515,I35559,I35658,);
not I_1952 (I35667,I84);
DFFARX1 I_1953 (I172,I515,I35559,I35694,);
not I_1954 (I35703,I35694);
nor I_1955 (I35721,I35703,I35595);
and I_1956 (I35739,I35721,I84);
nor I_1957 (I35757,I35703,I35667);
nor I_1958 (I35775,I35658,I35757);
DFFARX1 I_1959 (I324,I515,I35559,I35802,);
nor I_1960 (I35811,I35802,I35658);
not I_1961 (I35829,I35811);
not I_1962 (I35847,I35802);
nor I_1963 (I35865,I35847,I35739);
DFFARX1 I_1964 (I35865,I515,I35559,I35892,);
nand I_1965 (I35901,I332,I420);
and I_1966 (I35919,I35901,I268);
DFFARX1 I_1967 (I35919,I515,I35559,I35946,);
nor I_1968 (I35955,I35946,I35802);
DFFARX1 I_1969 (I35955,I515,I35559,I35982,);
nand I_1970 (I35991,I35946,I35847);
nand I_1971 (I36009,I35829,I35991);
not I_1972 (I36027,I35946);
nor I_1973 (I36045,I36027,I35739);
DFFARX1 I_1974 (I36045,I515,I35559,I36072,);
nor I_1975 (I36081,I196,I420);
or I_1976 (I36099,I35802,I36081);
nor I_1977 (I36117,I35946,I36081);
or I_1978 (I36135,I35658,I36081);
DFFARX1 I_1979 (I36081,I515,I35559,I36162,);
not I_1980 (I36171,I522);
DFFARX1 I_1981 (I36135,I515,I36171,I36198,);
DFFARX1 I_1982 (I35982,I515,I36171,I36216,);
not I_1983 (I36225,I36216);
not I_1984 (I36243,I35775);
nor I_1985 (I36261,I36243,I35982);
not I_1986 (I36279,I36009);
nor I_1987 (I36297,I36261,I35892);
nor I_1988 (I36315,I36216,I36297);
DFFARX1 I_1989 (I36315,I515,I36171,I36342,);
nor I_1990 (I36351,I35892,I35982);
nand I_1991 (I36369,I36351,I35775);
DFFARX1 I_1992 (I36369,I515,I36171,I36396,);
nor I_1993 (I36405,I36279,I35892);
nand I_1994 (I36423,I36405,I36117);
nor I_1995 (I36441,I36198,I36423);
DFFARX1 I_1996 (I36441,I515,I36171,I36468,);
not I_1997 (I36477,I36423);
nand I_1998 (I36495,I36216,I36477);
DFFARX1 I_1999 (I36423,I515,I36171,I36522,);
not I_2000 (I36531,I36522);
not I_2001 (I36549,I35892);
not I_2002 (I36567,I36099);
nor I_2003 (I36585,I36567,I36009);
nor I_2004 (I36603,I36531,I36585);
nor I_2005 (I36621,I36567,I36072);
and I_2006 (I36639,I36621,I36162);
or I_2007 (I36657,I36639,I36117);
DFFARX1 I_2008 (I36657,I515,I36171,I36684,);
nor I_2009 (I36693,I36684,I36198);
not I_2010 (I36711,I36684);
and I_2011 (I36729,I36711,I36198);
nor I_2012 (I36747,I36225,I36729);
nand I_2013 (I36765,I36711,I36279);
nor I_2014 (I36783,I36567,I36765);
nand I_2015 (I36801,I36711,I36477);
nand I_2016 (I36819,I36279,I36099);
nor I_2017 (I36837,I36549,I36819);
not I_2018 (I36855,I522);
DFFARX1 I_2019 (I36693,I515,I36855,I36882,);
DFFARX1 I_2020 (I36882,I515,I36855,I36900,);
not I_2021 (I36909,I36900);
DFFARX1 I_2022 (I36783,I515,I36855,I36936,);
not I_2023 (I36945,I36468);
nor I_2024 (I36963,I36882,I36945);
not I_2025 (I36981,I36495);
not I_2026 (I36999,I36747);
nand I_2027 (I37017,I36999,I36495);
nor I_2028 (I37035,I36945,I37017);
nor I_2029 (I37053,I36936,I37035);
DFFARX1 I_2030 (I36999,I515,I36855,I37080,);
nor I_2031 (I37089,I36747,I36837);
nand I_2032 (I37107,I37089,I36342);
nor I_2033 (I37125,I37107,I36981);
nand I_2034 (I37143,I37125,I36468);
DFFARX1 I_2035 (I37107,I515,I36855,I37170,);
nand I_2036 (I37179,I36981,I36747);
nor I_2037 (I37197,I36981,I36747);
nand I_2038 (I37215,I36963,I37197);
not I_2039 (I37233,I36396);
nor I_2040 (I37251,I37233,I37179);
DFFARX1 I_2041 (I37251,I515,I36855,I37278,);
nor I_2042 (I37287,I37233,I36603);
and I_2043 (I37305,I37287,I36801);
or I_2044 (I37323,I37305,I36468);
DFFARX1 I_2045 (I37323,I515,I36855,I37350,);
nor I_2046 (I37359,I37350,I36936);
nor I_2047 (I37377,I36882,I37359);
not I_2048 (I37395,I37350);
nor I_2049 (I37413,I37395,I37053);
DFFARX1 I_2050 (I37413,I515,I36855,I37440,);
nand I_2051 (I37449,I37395,I36981);
nor I_2052 (I37467,I37233,I37449);
not I_2053 (I37485,I522);
DFFARX1 I_2054 (I37467,I515,I37485,I37512,);
nand I_2055 (I37521,I37467,I37440);
and I_2056 (I37539,I37521,I37278);
DFFARX1 I_2057 (I37539,I515,I37485,I37566,);
nor I_2058 (I37575,I37566,I37512);
not I_2059 (I37593,I37566);
DFFARX1 I_2060 (I36909,I515,I37485,I37620,);
nand I_2061 (I37629,I37620,I37080);
not I_2062 (I37647,I37629);
DFFARX1 I_2063 (I37647,I515,I37485,I37674,);
not I_2064 (I37683,I37674);
nor I_2065 (I37701,I37512,I37629);
nor I_2066 (I37719,I37566,I37701);
DFFARX1 I_2067 (I37215,I515,I37485,I37746,);
DFFARX1 I_2068 (I37746,I515,I37485,I37764,);
not I_2069 (I37773,I37764);
not I_2070 (I37791,I37746);
nand I_2071 (I37809,I37791,I37593);
nand I_2072 (I37827,I37278,I37377);
and I_2073 (I37845,I37827,I37170);
DFFARX1 I_2074 (I37845,I515,I37485,I37872,);
nor I_2075 (I37881,I37872,I37512);
DFFARX1 I_2076 (I37881,I515,I37485,I37908,);
DFFARX1 I_2077 (I37872,I515,I37485,I37926,);
nor I_2078 (I37935,I37143,I37377);
not I_2079 (I37953,I37935);
nor I_2080 (I37971,I37773,I37953);
nand I_2081 (I37989,I37791,I37953);
nor I_2082 (I38007,I37512,I37935);
DFFARX1 I_2083 (I37935,I515,I37485,I38034,);
not I_2084 (I38043,I522);
DFFARX1 I_2085 (I37971,I515,I38043,I38070,);
DFFARX1 I_2086 (I38007,I515,I38043,I38088,);
not I_2087 (I38097,I38088);
nor I_2088 (I38115,I38070,I38097);
DFFARX1 I_2089 (I38097,I515,I38043,I38142,);
nor I_2090 (I38151,I37575,I38034);
and I_2091 (I38169,I38151,I37926);
nor I_2092 (I38187,I38169,I37575);
not I_2093 (I38205,I37575);
and I_2094 (I38223,I38205,I37908);
nand I_2095 (I38241,I38223,I37809);
nor I_2096 (I38259,I38205,I38241);
DFFARX1 I_2097 (I38259,I515,I38043,I38286,);
not I_2098 (I38295,I38241);
nand I_2099 (I38313,I38097,I38295);
nand I_2100 (I38331,I38169,I38295);
DFFARX1 I_2101 (I38205,I515,I38043,I38358,);
not I_2102 (I38367,I37683);
nor I_2103 (I38385,I38367,I37908);
nor I_2104 (I38403,I38385,I38187);
DFFARX1 I_2105 (I38403,I515,I38043,I38430,);
not I_2106 (I38439,I38385);
DFFARX1 I_2107 (I38439,I515,I38043,I38466,);
not I_2108 (I38475,I38466);
nor I_2109 (I38493,I38475,I38385);
nor I_2110 (I38511,I38367,I37719);
and I_2111 (I38529,I38511,I37989);
or I_2112 (I38547,I38529,I37908);
DFFARX1 I_2113 (I38547,I515,I38043,I38574,);
not I_2114 (I38583,I38574);
nand I_2115 (I38601,I38583,I38295);
not I_2116 (I38619,I38601);
nand I_2117 (I38637,I38601,I38313);
nand I_2118 (I38655,I38583,I38169);
not I_2119 (I38673,I522);
DFFARX1 I_2120 (I38331,I515,I38673,I38700,);
not I_2121 (I38709,I38700);
nand I_2122 (I38727,I38655,I38358);
and I_2123 (I38745,I38727,I38115);
DFFARX1 I_2124 (I38745,I515,I38673,I38772,);
DFFARX1 I_2125 (I38430,I515,I38673,I38790,);
and I_2126 (I38799,I38790,I38493);
nor I_2127 (I38817,I38772,I38799);
DFFARX1 I_2128 (I38817,I515,I38673,I38844,);
nand I_2129 (I38853,I38790,I38493);
nand I_2130 (I38871,I38709,I38853);
not I_2131 (I38889,I38871);
DFFARX1 I_2132 (I38637,I515,I38673,I38916,);
DFFARX1 I_2133 (I38916,I515,I38673,I38934,);
nand I_2134 (I38943,I38142,I38619);
and I_2135 (I38961,I38943,I38286);
DFFARX1 I_2136 (I38961,I515,I38673,I38988,);
DFFARX1 I_2137 (I38988,I515,I38673,I39006,);
not I_2138 (I39015,I39006);
not I_2139 (I39033,I38988);
nand I_2140 (I39051,I39033,I38853);
nor I_2141 (I39069,I38286,I38619);
not I_2142 (I39087,I39069);
nor I_2143 (I39105,I39033,I39087);
nor I_2144 (I39123,I38709,I39105);
DFFARX1 I_2145 (I39123,I515,I38673,I39150,);
nor I_2146 (I39159,I38772,I39087);
nor I_2147 (I39177,I38988,I39159);
nor I_2148 (I39195,I38916,I39069);
nor I_2149 (I39213,I38772,I39069);
not I_2150 (I39231,I522);
DFFARX1 I_2151 (I39015,I515,I39231,I39258,);
and I_2152 (I39267,I39258,I38844);
DFFARX1 I_2153 (I39267,I515,I39231,I39294,);
DFFARX1 I_2154 (I39150,I515,I39231,I39312,);
not I_2155 (I39321,I39177);
not I_2156 (I39339,I39213);
nand I_2157 (I39357,I39339,I39321);
nor I_2158 (I39375,I39312,I39357);
DFFARX1 I_2159 (I39357,I515,I39231,I39402,);
not I_2160 (I39411,I39402);
not I_2161 (I39429,I38889);
nand I_2162 (I39447,I39339,I39429);
DFFARX1 I_2163 (I39447,I515,I39231,I39474,);
not I_2164 (I39483,I39474);
not I_2165 (I39501,I39213);
nand I_2166 (I39519,I39501,I38934);
and I_2167 (I39537,I39321,I39519);
nor I_2168 (I39555,I39447,I39537);
DFFARX1 I_2169 (I39555,I515,I39231,I39582,);
DFFARX1 I_2170 (I39537,I515,I39231,I39600,);
nor I_2171 (I39609,I39213,I39195);
nor I_2172 (I39627,I39447,I39609);
or I_2173 (I39645,I39213,I39195);
nor I_2174 (I39663,I39051,I38844);
DFFARX1 I_2175 (I39663,I515,I39231,I39690,);
not I_2176 (I39699,I39690);
nor I_2177 (I39717,I39699,I39483);
nand I_2178 (I39735,I39699,I39312);
not I_2179 (I39753,I39051);
nand I_2180 (I39771,I39753,I39429);
nand I_2181 (I39789,I39699,I39771);
nand I_2182 (I39807,I39789,I39735);
nand I_2183 (I39825,I39771,I39645);
not I_2184 (I39843,I522);
DFFARX1 I_2185 (I39582,I515,I39843,I39870,);
nand I_2186 (I39879,I39294,I39582);
and I_2187 (I39897,I39879,I39717);
DFFARX1 I_2188 (I39897,I515,I39843,I39924,);
nor I_2189 (I39933,I39924,I39870);
not I_2190 (I39951,I39924);
DFFARX1 I_2191 (I39411,I515,I39843,I39978,);
nand I_2192 (I39987,I39978,I39825);
not I_2193 (I40005,I39987);
DFFARX1 I_2194 (I40005,I515,I39843,I40032,);
not I_2195 (I40041,I40032);
nor I_2196 (I40059,I39870,I39987);
nor I_2197 (I40077,I39924,I40059);
DFFARX1 I_2198 (I39375,I515,I39843,I40104,);
DFFARX1 I_2199 (I40104,I515,I39843,I40122,);
not I_2200 (I40131,I40122);
not I_2201 (I40149,I40104);
nand I_2202 (I40167,I40149,I39951);
nand I_2203 (I40185,I39375,I39807);
and I_2204 (I40203,I40185,I39600);
DFFARX1 I_2205 (I40203,I515,I39843,I40230,);
nor I_2206 (I40239,I40230,I39870);
DFFARX1 I_2207 (I40239,I515,I39843,I40266,);
DFFARX1 I_2208 (I40230,I515,I39843,I40284,);
nor I_2209 (I40293,I39627,I39807);
not I_2210 (I40311,I40293);
nor I_2211 (I40329,I40131,I40311);
nand I_2212 (I40347,I40149,I40311);
nor I_2213 (I40365,I39870,I40293);
DFFARX1 I_2214 (I40293,I515,I39843,I40392,);
not I_2215 (I40401,I522);
DFFARX1 I_2216 (I40041,I515,I40401,I40428,);
and I_2217 (I40437,I40428,I40167);
DFFARX1 I_2218 (I40437,I515,I40401,I40464,);
DFFARX1 I_2219 (I40284,I515,I40401,I40482,);
not I_2220 (I40491,I40266);
not I_2221 (I40509,I40329);
nand I_2222 (I40527,I40509,I40491);
nor I_2223 (I40545,I40482,I40527);
DFFARX1 I_2224 (I40527,I515,I40401,I40572,);
not I_2225 (I40581,I40572);
not I_2226 (I40599,I40392);
nand I_2227 (I40617,I40509,I40599);
DFFARX1 I_2228 (I40617,I515,I40401,I40644,);
not I_2229 (I40653,I40644);
not I_2230 (I40671,I40365);
nand I_2231 (I40689,I40671,I39933);
and I_2232 (I40707,I40491,I40689);
nor I_2233 (I40725,I40617,I40707);
DFFARX1 I_2234 (I40725,I515,I40401,I40752,);
DFFARX1 I_2235 (I40707,I515,I40401,I40770,);
nor I_2236 (I40779,I40365,I40077);
nor I_2237 (I40797,I40617,I40779);
or I_2238 (I40815,I40365,I40077);
nor I_2239 (I40833,I40347,I40266);
DFFARX1 I_2240 (I40833,I515,I40401,I40860,);
not I_2241 (I40869,I40860);
nor I_2242 (I40887,I40869,I40653);
nand I_2243 (I40905,I40869,I40482);
not I_2244 (I40923,I40347);
nand I_2245 (I40941,I40923,I40599);
nand I_2246 (I40959,I40869,I40941);
nand I_2247 (I40977,I40959,I40905);
nand I_2248 (I40995,I40941,I40815);
not I_2249 (I41013,I522);
DFFARX1 I_2250 (I40752,I515,I41013,I41040,);
nand I_2251 (I41049,I40464,I40752);
and I_2252 (I41067,I41049,I40887);
DFFARX1 I_2253 (I41067,I515,I41013,I41094,);
nor I_2254 (I41103,I41094,I41040);
not I_2255 (I41121,I41094);
DFFARX1 I_2256 (I40581,I515,I41013,I41148,);
nand I_2257 (I41157,I41148,I40995);
not I_2258 (I41175,I41157);
DFFARX1 I_2259 (I41175,I515,I41013,I41202,);
not I_2260 (I41211,I41202);
nor I_2261 (I41229,I41040,I41157);
nor I_2262 (I41247,I41094,I41229);
DFFARX1 I_2263 (I40545,I515,I41013,I41274,);
DFFARX1 I_2264 (I41274,I515,I41013,I41292,);
not I_2265 (I41301,I41292);
not I_2266 (I41319,I41274);
nand I_2267 (I41337,I41319,I41121);
nand I_2268 (I41355,I40545,I40977);
and I_2269 (I41373,I41355,I40770);
DFFARX1 I_2270 (I41373,I515,I41013,I41400,);
nor I_2271 (I41409,I41400,I41040);
DFFARX1 I_2272 (I41409,I515,I41013,I41436,);
DFFARX1 I_2273 (I41400,I515,I41013,I41454,);
nor I_2274 (I41463,I40797,I40977);
not I_2275 (I41481,I41463);
nor I_2276 (I41499,I41301,I41481);
nand I_2277 (I41517,I41319,I41481);
nor I_2278 (I41535,I41040,I41463);
DFFARX1 I_2279 (I41463,I515,I41013,I41562,);
not I_2280 (I41571,I522);
DFFARX1 I_2281 (I41562,I515,I41571,I41598,);
not I_2282 (I41607,I41598);
nand I_2283 (I41625,I41211,I41103);
and I_2284 (I41643,I41625,I41436);
DFFARX1 I_2285 (I41643,I515,I41571,I41670,);
not I_2286 (I41679,I41517);
DFFARX1 I_2287 (I41436,I515,I41571,I41706,);
not I_2288 (I41715,I41706);
nor I_2289 (I41733,I41715,I41607);
and I_2290 (I41751,I41733,I41517);
nor I_2291 (I41769,I41715,I41679);
nor I_2292 (I41787,I41670,I41769);
DFFARX1 I_2293 (I41247,I515,I41571,I41814,);
nor I_2294 (I41823,I41814,I41670);
not I_2295 (I41841,I41823);
not I_2296 (I41859,I41814);
nor I_2297 (I41877,I41859,I41751);
DFFARX1 I_2298 (I41877,I515,I41571,I41904,);
nand I_2299 (I41913,I41337,I41499);
and I_2300 (I41931,I41913,I41454);
DFFARX1 I_2301 (I41931,I515,I41571,I41958,);
nor I_2302 (I41967,I41958,I41814);
DFFARX1 I_2303 (I41967,I515,I41571,I41994,);
nand I_2304 (I42003,I41958,I41859);
nand I_2305 (I42021,I41841,I42003);
not I_2306 (I42039,I41958);
nor I_2307 (I42057,I42039,I41751);
DFFARX1 I_2308 (I42057,I515,I41571,I42084,);
nor I_2309 (I42093,I41535,I41499);
or I_2310 (I42111,I41814,I42093);
nor I_2311 (I42129,I41958,I42093);
or I_2312 (I42147,I41670,I42093);
DFFARX1 I_2313 (I42093,I515,I41571,I42174,);
not I_2314 (I42183,I522);
DFFARX1 I_2315 (I42111,I515,I42183,I42210,);
nand I_2316 (I42219,I42129,I41904);
and I_2317 (I42237,I42219,I42174);
DFFARX1 I_2318 (I42237,I515,I42183,I42264,);
nor I_2319 (I42273,I42264,I42210);
not I_2320 (I42291,I42264);
DFFARX1 I_2321 (I42021,I515,I42183,I42318,);
nand I_2322 (I42327,I42318,I42129);
not I_2323 (I42345,I42327);
DFFARX1 I_2324 (I42345,I515,I42183,I42372,);
not I_2325 (I42381,I42372);
nor I_2326 (I42399,I42210,I42327);
nor I_2327 (I42417,I42264,I42399);
DFFARX1 I_2328 (I42147,I515,I42183,I42444,);
DFFARX1 I_2329 (I42444,I515,I42183,I42462,);
not I_2330 (I42471,I42462);
not I_2331 (I42489,I42444);
nand I_2332 (I42507,I42489,I42291);
nand I_2333 (I42525,I41994,I41787);
and I_2334 (I42543,I42525,I41994);
DFFARX1 I_2335 (I42543,I515,I42183,I42570,);
nor I_2336 (I42579,I42570,I42210);
DFFARX1 I_2337 (I42579,I515,I42183,I42606,);
DFFARX1 I_2338 (I42570,I515,I42183,I42624,);
nor I_2339 (I42633,I42084,I41787);
not I_2340 (I42651,I42633);
nor I_2341 (I42669,I42471,I42651);
nand I_2342 (I42687,I42489,I42651);
nor I_2343 (I42705,I42210,I42633);
DFFARX1 I_2344 (I42633,I515,I42183,I42732,);
not I_2345 (I42741,I522);
DFFARX1 I_2346 (I42606,I515,I42741,I42768,);
DFFARX1 I_2347 (I42768,I515,I42741,I42786,);
not I_2348 (I42795,I42786);
not I_2349 (I42813,I42768);
DFFARX1 I_2350 (I42705,I515,I42741,I42840,);
not I_2351 (I42849,I42840);
and I_2352 (I42867,I42813,I42507);
not I_2353 (I42885,I42606);
nand I_2354 (I42903,I42885,I42507);
not I_2355 (I42921,I42417);
nor I_2356 (I42939,I42921,I42732);
nand I_2357 (I42957,I42939,I42669);
nor I_2358 (I42975,I42957,I42903);
DFFARX1 I_2359 (I42975,I515,I42741,I43002,);
not I_2360 (I43011,I42957);
not I_2361 (I43029,I42732);
nand I_2362 (I43047,I43029,I42507);
nor I_2363 (I43065,I42732,I42606);
nand I_2364 (I43083,I42867,I43065);
nand I_2365 (I43101,I42813,I42732);
nand I_2366 (I43119,I42921,I42624);
DFFARX1 I_2367 (I43119,I515,I42741,I43146,);
DFFARX1 I_2368 (I43119,I515,I42741,I43164,);
not I_2369 (I43173,I42624);
nor I_2370 (I43191,I43173,I42687);
and I_2371 (I43209,I43191,I42381);
or I_2372 (I43227,I43209,I42273);
DFFARX1 I_2373 (I43227,I515,I42741,I43254,);
nand I_2374 (I43263,I43254,I42885);
nor I_2375 (I43281,I43263,I43047);
nor I_2376 (I43299,I43254,I42849);
DFFARX1 I_2377 (I43254,I515,I42741,I43326,);
not I_2378 (I43335,I43326);
nor I_2379 (I43353,I43335,I43011);
not I_2380 (I43371,I522);
DFFARX1 I_2381 (I43002,I515,I43371,I43398,);
not I_2382 (I43407,I43398);
nand I_2383 (I43425,I43299,I42795);
and I_2384 (I43443,I43425,I43083);
DFFARX1 I_2385 (I43443,I515,I43371,I43470,);
not I_2386 (I43479,I43281);
DFFARX1 I_2387 (I43002,I515,I43371,I43506,);
not I_2388 (I43515,I43506);
nor I_2389 (I43533,I43515,I43407);
and I_2390 (I43551,I43533,I43281);
nor I_2391 (I43569,I43515,I43479);
nor I_2392 (I43587,I43470,I43569);
DFFARX1 I_2393 (I43353,I515,I43371,I43614,);
nor I_2394 (I43623,I43614,I43470);
not I_2395 (I43641,I43623);
not I_2396 (I43659,I43614);
nor I_2397 (I43677,I43659,I43551);
DFFARX1 I_2398 (I43677,I515,I43371,I43704,);
nand I_2399 (I43713,I43299,I43101);
and I_2400 (I43731,I43713,I43164);
DFFARX1 I_2401 (I43731,I515,I43371,I43758,);
nor I_2402 (I43767,I43758,I43614);
DFFARX1 I_2403 (I43767,I515,I43371,I43794,);
nand I_2404 (I43803,I43758,I43659);
nand I_2405 (I43821,I43641,I43803);
not I_2406 (I43839,I43758);
nor I_2407 (I43857,I43839,I43551);
DFFARX1 I_2408 (I43857,I515,I43371,I43884,);
nor I_2409 (I43893,I43146,I43101);
or I_2410 (I43911,I43614,I43893);
nor I_2411 (I43929,I43758,I43893);
or I_2412 (I43947,I43470,I43893);
DFFARX1 I_2413 (I43893,I515,I43371,I43974,);
not I_2414 (I43983,I522);
DFFARX1 I_2415 (I43587,I515,I43983,I44010,);
and I_2416 (I44019,I44010,I43929);
DFFARX1 I_2417 (I44019,I515,I43983,I44046,);
DFFARX1 I_2418 (I43947,I515,I43983,I44064,);
not I_2419 (I44073,I43794);
not I_2420 (I44091,I43974);
nand I_2421 (I44109,I44091,I44073);
nor I_2422 (I44127,I44064,I44109);
DFFARX1 I_2423 (I44109,I515,I43983,I44154,);
not I_2424 (I44163,I44154);
not I_2425 (I44181,I43911);
nand I_2426 (I44199,I44091,I44181);
DFFARX1 I_2427 (I44199,I515,I43983,I44226,);
not I_2428 (I44235,I44226);
not I_2429 (I44253,I43884);
nand I_2430 (I44271,I44253,I43704);
and I_2431 (I44289,I44073,I44271);
nor I_2432 (I44307,I44199,I44289);
DFFARX1 I_2433 (I44307,I515,I43983,I44334,);
DFFARX1 I_2434 (I44289,I515,I43983,I44352,);
nor I_2435 (I44361,I43884,I43821);
nor I_2436 (I44379,I44199,I44361);
or I_2437 (I44397,I43884,I43821);
nor I_2438 (I44415,I43794,I43929);
DFFARX1 I_2439 (I44415,I515,I43983,I44442,);
not I_2440 (I44451,I44442);
nor I_2441 (I44469,I44451,I44235);
nand I_2442 (I44487,I44451,I44064);
not I_2443 (I44505,I43794);
nand I_2444 (I44523,I44505,I44181);
nand I_2445 (I44541,I44451,I44523);
nand I_2446 (I44559,I44541,I44487);
nand I_2447 (I44577,I44523,I44397);
not I_2448 (I44595,I522);
DFFARX1 I_2449 (I44469,I515,I44595,I44622,);
DFFARX1 I_2450 (I44622,I515,I44595,I44640,);
not I_2451 (I44649,I44640);
DFFARX1 I_2452 (I44334,I515,I44595,I44676,);
not I_2453 (I44685,I44577);
nor I_2454 (I44703,I44622,I44685);
not I_2455 (I44721,I44352);
not I_2456 (I44739,I44379);
nand I_2457 (I44757,I44739,I44352);
nor I_2458 (I44775,I44685,I44757);
nor I_2459 (I44793,I44676,I44775);
DFFARX1 I_2460 (I44739,I515,I44595,I44820,);
nor I_2461 (I44829,I44379,I44163);
nand I_2462 (I44847,I44829,I44127);
nor I_2463 (I44865,I44847,I44721);
nand I_2464 (I44883,I44865,I44577);
DFFARX1 I_2465 (I44847,I515,I44595,I44910,);
nand I_2466 (I44919,I44721,I44379);
nor I_2467 (I44937,I44721,I44379);
nand I_2468 (I44955,I44703,I44937);
not I_2469 (I44973,I44559);
nor I_2470 (I44991,I44973,I44919);
DFFARX1 I_2471 (I44991,I515,I44595,I45018,);
nor I_2472 (I45027,I44973,I44046);
and I_2473 (I45045,I45027,I44334);
or I_2474 (I45063,I45045,I44127);
DFFARX1 I_2475 (I45063,I515,I44595,I45090,);
nor I_2476 (I45099,I45090,I44676);
nor I_2477 (I45117,I44622,I45099);
not I_2478 (I45135,I45090);
nor I_2479 (I45153,I45135,I44793);
DFFARX1 I_2480 (I45153,I515,I44595,I45180,);
nand I_2481 (I45189,I45135,I44721);
nor I_2482 (I45207,I44973,I45189);
not I_2483 (I45225,I522);
DFFARX1 I_2484 (I45117,I515,I45225,I45252,);
DFFARX1 I_2485 (I45252,I515,I45225,I45270,);
not I_2486 (I45279,I45270);
nand I_2487 (I45297,I45180,I45207);
and I_2488 (I45315,I45297,I45018);
DFFARX1 I_2489 (I45315,I515,I45225,I45342,);
DFFARX1 I_2490 (I45342,I515,I45225,I45360,);
DFFARX1 I_2491 (I45342,I515,I45225,I45378,);
DFFARX1 I_2492 (I44955,I515,I45225,I45396,);
nand I_2493 (I45405,I45396,I44883);
not I_2494 (I45423,I45405);
nor I_2495 (I45441,I45252,I45423);
DFFARX1 I_2496 (I44649,I515,I45225,I45468,);
not I_2497 (I45477,I45468);
nor I_2498 (I45495,I45477,I45279);
nand I_2499 (I45513,I45477,I45405);
nand I_2500 (I45531,I44910,I44820);
and I_2501 (I45549,I45531,I45207);
DFFARX1 I_2502 (I45549,I515,I45225,I45576,);
nor I_2503 (I45585,I45576,I45252);
DFFARX1 I_2504 (I45585,I515,I45225,I45612,);
not I_2505 (I45621,I45576);
nor I_2506 (I45639,I45018,I44820);
not I_2507 (I45657,I45639);
nor I_2508 (I45675,I45405,I45657);
nor I_2509 (I45693,I45621,I45675);
DFFARX1 I_2510 (I45693,I515,I45225,I45720,);
nor I_2511 (I45729,I45576,I45657);
nor I_2512 (I45747,I45423,I45729);
nor I_2513 (I45765,I45576,I45639);
not I_2514 (I45783,I522);
DFFARX1 I_2515 (I45441,I515,I45783,I45810,);
not I_2516 (I45819,I45810);
nand I_2517 (I45837,I45747,I45612);
and I_2518 (I45855,I45837,I45612);
DFFARX1 I_2519 (I45855,I515,I45783,I45882,);
not I_2520 (I45891,I45765);
DFFARX1 I_2521 (I45495,I515,I45783,I45918,);
not I_2522 (I45927,I45918);
nor I_2523 (I45945,I45927,I45819);
and I_2524 (I45963,I45945,I45765);
nor I_2525 (I45981,I45927,I45891);
nor I_2526 (I45999,I45882,I45981);
DFFARX1 I_2527 (I45765,I515,I45783,I46026,);
nor I_2528 (I46035,I46026,I45882);
not I_2529 (I46053,I46035);
not I_2530 (I46071,I46026);
nor I_2531 (I46089,I46071,I45963);
DFFARX1 I_2532 (I46089,I515,I45783,I46116,);
nand I_2533 (I46125,I45720,I45513);
and I_2534 (I46143,I46125,I45378);
DFFARX1 I_2535 (I46143,I515,I45783,I46170,);
nor I_2536 (I46179,I46170,I46026);
DFFARX1 I_2537 (I46179,I515,I45783,I46206,);
nand I_2538 (I46215,I46170,I46071);
nand I_2539 (I46233,I46053,I46215);
not I_2540 (I46251,I46170);
nor I_2541 (I46269,I46251,I45963);
DFFARX1 I_2542 (I46269,I515,I45783,I46296,);
nor I_2543 (I46305,I45360,I45513);
or I_2544 (I46323,I46026,I46305);
nor I_2545 (I46341,I46170,I46305);
or I_2546 (I46359,I45882,I46305);
DFFARX1 I_2547 (I46305,I515,I45783,I46386,);
not I_2548 (I46395,I522);
DFFARX1 I_2549 (I46359,I515,I46395,I46422,);
DFFARX1 I_2550 (I46206,I515,I46395,I46440,);
not I_2551 (I46449,I46440);
not I_2552 (I46467,I45999);
nor I_2553 (I46485,I46467,I46206);
not I_2554 (I46503,I46233);
nor I_2555 (I46521,I46485,I46116);
nor I_2556 (I46539,I46440,I46521);
DFFARX1 I_2557 (I46539,I515,I46395,I46566,);
nor I_2558 (I46575,I46116,I46206);
nand I_2559 (I46593,I46575,I45999);
DFFARX1 I_2560 (I46593,I515,I46395,I46620,);
nor I_2561 (I46629,I46503,I46116);
nand I_2562 (I46647,I46629,I46341);
nor I_2563 (I46665,I46422,I46647);
DFFARX1 I_2564 (I46665,I515,I46395,I46692,);
not I_2565 (I46701,I46647);
nand I_2566 (I46719,I46440,I46701);
DFFARX1 I_2567 (I46647,I515,I46395,I46746,);
not I_2568 (I46755,I46746);
not I_2569 (I46773,I46116);
not I_2570 (I46791,I46323);
nor I_2571 (I46809,I46791,I46233);
nor I_2572 (I46827,I46755,I46809);
nor I_2573 (I46845,I46791,I46296);
and I_2574 (I46863,I46845,I46386);
or I_2575 (I46881,I46863,I46341);
DFFARX1 I_2576 (I46881,I515,I46395,I46908,);
nor I_2577 (I46917,I46908,I46422);
not I_2578 (I46935,I46908);
and I_2579 (I46953,I46935,I46422);
nor I_2580 (I46971,I46449,I46953);
nand I_2581 (I46989,I46935,I46503);
nor I_2582 (I47007,I46791,I46989);
nand I_2583 (I47025,I46935,I46701);
nand I_2584 (I47043,I46503,I46323);
nor I_2585 (I47061,I46773,I47043);
not I_2586 (I47079,I522);
DFFARX1 I_2587 (I47007,I515,I47079,I47106,);
nand I_2588 (I47115,I46692,I47061);
and I_2589 (I47133,I47115,I46971);
DFFARX1 I_2590 (I47133,I515,I47079,I47160,);
nor I_2591 (I47169,I47160,I47106);
not I_2592 (I47187,I47160);
DFFARX1 I_2593 (I46620,I515,I47079,I47214,);
nand I_2594 (I47223,I47214,I47025);
not I_2595 (I47241,I47223);
DFFARX1 I_2596 (I47241,I515,I47079,I47268,);
not I_2597 (I47277,I47268);
nor I_2598 (I47295,I47106,I47223);
nor I_2599 (I47313,I47160,I47295);
DFFARX1 I_2600 (I46719,I515,I47079,I47340,);
DFFARX1 I_2601 (I47340,I515,I47079,I47358,);
not I_2602 (I47367,I47358);
not I_2603 (I47385,I47340);
nand I_2604 (I47403,I47385,I47187);
nand I_2605 (I47421,I46692,I46827);
and I_2606 (I47439,I47421,I46917);
DFFARX1 I_2607 (I47439,I515,I47079,I47466,);
nor I_2608 (I47475,I47466,I47106);
DFFARX1 I_2609 (I47475,I515,I47079,I47502,);
DFFARX1 I_2610 (I47466,I515,I47079,I47520,);
nor I_2611 (I47529,I46566,I46827);
not I_2612 (I47547,I47529);
nor I_2613 (I47565,I47367,I47547);
nand I_2614 (I47583,I47385,I47547);
nor I_2615 (I47601,I47106,I47529);
DFFARX1 I_2616 (I47529,I515,I47079,I47628,);
not I_2617 (I47637,I522);
DFFARX1 I_2618 (I47583,I515,I47637,I47664,);
nand I_2619 (I47673,I47664,I47277);
not I_2620 (I47691,I47673);
DFFARX1 I_2621 (I47565,I515,I47637,I47718,);
not I_2622 (I47727,I47718);
not I_2623 (I47745,I47313);
or I_2624 (I47763,I47628,I47313);
nor I_2625 (I47781,I47628,I47313);
or I_2626 (I47799,I47601,I47628);
DFFARX1 I_2627 (I47799,I515,I47637,I47826,);
not I_2628 (I47835,I47169);
nand I_2629 (I47853,I47835,I47502);
nand I_2630 (I47871,I47745,I47853);
and I_2631 (I47889,I47727,I47871);
nor I_2632 (I47907,I47169,I47403);
and I_2633 (I47925,I47727,I47907);
nor I_2634 (I47943,I47691,I47925);
DFFARX1 I_2635 (I47907,I515,I47637,I47970,);
not I_2636 (I47979,I47970);
nor I_2637 (I47997,I47727,I47979);
or I_2638 (I48015,I47799,I47520);
nor I_2639 (I48033,I47520,I47601);
nand I_2640 (I48051,I47871,I48033);
nand I_2641 (I48069,I48015,I48051);
DFFARX1 I_2642 (I48069,I515,I47637,I48096,);
nor I_2643 (I48105,I48033,I47763);
DFFARX1 I_2644 (I48105,I515,I47637,I48132,);
nor I_2645 (I48141,I47520,I47502);
DFFARX1 I_2646 (I48141,I515,I47637,I48168,);
DFFARX1 I_2647 (I48168,I515,I47637,I48186,);
not I_2648 (I48195,I48168);
nand I_2649 (I48213,I48195,I47673);
nand I_2650 (I48231,I48195,I47781);
not I_2651 (I48249,I522);
DFFARX1 I_2652 (I47997,I515,I48249,I48276,);
DFFARX1 I_2653 (I47943,I515,I48249,I48294,);
not I_2654 (I48303,I48294);
nor I_2655 (I48321,I48276,I48303);
DFFARX1 I_2656 (I48303,I515,I48249,I48348,);
nor I_2657 (I48357,I48132,I48186);
and I_2658 (I48375,I48357,I47889);
nor I_2659 (I48393,I48375,I48132);
not I_2660 (I48411,I48132);
and I_2661 (I48429,I48411,I48231);
nand I_2662 (I48447,I48429,I47826);
nor I_2663 (I48465,I48411,I48447);
DFFARX1 I_2664 (I48465,I515,I48249,I48492,);
not I_2665 (I48501,I48447);
nand I_2666 (I48519,I48303,I48501);
nand I_2667 (I48537,I48375,I48501);
DFFARX1 I_2668 (I48411,I515,I48249,I48564,);
not I_2669 (I48573,I48132);
nor I_2670 (I48591,I48573,I48231);
nor I_2671 (I48609,I48591,I48393);
DFFARX1 I_2672 (I48609,I515,I48249,I48636,);
not I_2673 (I48645,I48591);
DFFARX1 I_2674 (I48645,I515,I48249,I48672,);
not I_2675 (I48681,I48672);
nor I_2676 (I48699,I48681,I48591);
nor I_2677 (I48717,I48573,I47889);
and I_2678 (I48735,I48717,I48213);
or I_2679 (I48753,I48735,I48096);
DFFARX1 I_2680 (I48753,I515,I48249,I48780,);
not I_2681 (I48789,I48780);
nand I_2682 (I48807,I48789,I48501);
not I_2683 (I48825,I48807);
nand I_2684 (I48843,I48807,I48519);
nand I_2685 (I48861,I48789,I48375);
not I_2686 (I48879,I522);
DFFARX1 I_2687 (I48492,I515,I48879,I48906,);
DFFARX1 I_2688 (I48906,I515,I48879,I48924,);
not I_2689 (I48933,I48924);
nand I_2690 (I48951,I48321,I48843);
and I_2691 (I48969,I48951,I48348);
DFFARX1 I_2692 (I48969,I515,I48879,I48996,);
DFFARX1 I_2693 (I48996,I515,I48879,I49014,);
DFFARX1 I_2694 (I48996,I515,I48879,I49032,);
DFFARX1 I_2695 (I48699,I515,I48879,I49050,);
nand I_2696 (I49059,I49050,I48537);
not I_2697 (I49077,I49059);
nor I_2698 (I49095,I48906,I49077);
DFFARX1 I_2699 (I48492,I515,I48879,I49122,);
not I_2700 (I49131,I49122);
nor I_2701 (I49149,I49131,I48933);
nand I_2702 (I49167,I49131,I49059);
nand I_2703 (I49185,I48564,I48861);
and I_2704 (I49203,I49185,I48825);
DFFARX1 I_2705 (I49203,I515,I48879,I49230,);
nor I_2706 (I49239,I49230,I48906);
DFFARX1 I_2707 (I49239,I515,I48879,I49266,);
not I_2708 (I49275,I49230);
nor I_2709 (I49293,I48636,I48861);
not I_2710 (I49311,I49293);
nor I_2711 (I49329,I49059,I49311);
nor I_2712 (I49347,I49275,I49329);
DFFARX1 I_2713 (I49347,I515,I48879,I49374,);
nor I_2714 (I49383,I49230,I49311);
nor I_2715 (I49401,I49077,I49383);
nor I_2716 (I49419,I49230,I49293);
not I_2717 (I49437,I522);
DFFARX1 I_2718 (I49095,I515,I49437,I49464,);
DFFARX1 I_2719 (I49464,I515,I49437,I49482,);
not I_2720 (I49491,I49482);
not I_2721 (I49509,I49464);
nand I_2722 (I49527,I49266,I49032);
and I_2723 (I49545,I49527,I49419);
DFFARX1 I_2724 (I49545,I515,I49437,I49572,);
not I_2725 (I49581,I49572);
DFFARX1 I_2726 (I49014,I515,I49437,I49608,);
and I_2727 (I49617,I49608,I49149);
nand I_2728 (I49635,I49608,I49149);
nand I_2729 (I49653,I49581,I49635);
DFFARX1 I_2730 (I49374,I515,I49437,I49680,);
nor I_2731 (I49689,I49680,I49617);
DFFARX1 I_2732 (I49689,I515,I49437,I49716,);
nor I_2733 (I49725,I49680,I49572);
nand I_2734 (I49743,I49266,I49419);
and I_2735 (I49761,I49743,I49167);
DFFARX1 I_2736 (I49761,I515,I49437,I49788,);
nor I_2737 (I49797,I49788,I49680);
not I_2738 (I49815,I49788);
nor I_2739 (I49833,I49815,I49581);
nor I_2740 (I49851,I49509,I49833);
DFFARX1 I_2741 (I49851,I515,I49437,I49878,);
nor I_2742 (I49887,I49815,I49680);
nor I_2743 (I49905,I49401,I49419);
nor I_2744 (I49923,I49905,I49887);
not I_2745 (I49941,I49905);
nand I_2746 (I49959,I49635,I49941);
DFFARX1 I_2747 (I49905,I515,I49437,I49986,);
DFFARX1 I_2748 (I49905,I515,I49437,I50004,);
not I_2749 (I50013,I522);
DFFARX1 I_2750 (I49716,I515,I50013,I50040,);
and I_2751 (I50049,I50040,I49725);
DFFARX1 I_2752 (I50049,I515,I50013,I50076,);
DFFARX1 I_2753 (I49878,I515,I50013,I50094,);
not I_2754 (I50103,I49959);
not I_2755 (I50121,I49491);
nand I_2756 (I50139,I50121,I50103);
nor I_2757 (I50157,I50094,I50139);
DFFARX1 I_2758 (I50139,I515,I50013,I50184,);
not I_2759 (I50193,I50184);
not I_2760 (I50211,I49797);
nand I_2761 (I50229,I50121,I50211);
DFFARX1 I_2762 (I50229,I515,I50013,I50256,);
not I_2763 (I50265,I50256);
not I_2764 (I50283,I49653);
nand I_2765 (I50301,I50283,I49716);
and I_2766 (I50319,I50103,I50301);
nor I_2767 (I50337,I50229,I50319);
DFFARX1 I_2768 (I50337,I515,I50013,I50364,);
DFFARX1 I_2769 (I50319,I515,I50013,I50382,);
nor I_2770 (I50391,I49653,I49923);
nor I_2771 (I50409,I50229,I50391);
or I_2772 (I50427,I49653,I49923);
nor I_2773 (I50445,I49986,I50004);
DFFARX1 I_2774 (I50445,I515,I50013,I50472,);
not I_2775 (I50481,I50472);
nor I_2776 (I50499,I50481,I50265);
nand I_2777 (I50517,I50481,I50094);
not I_2778 (I50535,I49986);
nand I_2779 (I50553,I50535,I50211);
nand I_2780 (I50571,I50481,I50553);
nand I_2781 (I50589,I50571,I50517);
nand I_2782 (I50607,I50553,I50427);
not I_2783 (I50625,I522);
DFFARX1 I_2784 (I50364,I515,I50625,I50652,);
DFFARX1 I_2785 (I50652,I515,I50625,I50670,);
not I_2786 (I50679,I50670);
not I_2787 (I50697,I50652);
DFFARX1 I_2788 (I50364,I515,I50625,I50724,);
not I_2789 (I50733,I50724);
and I_2790 (I50751,I50697,I50157);
not I_2791 (I50769,I50076);
nand I_2792 (I50787,I50769,I50157);
not I_2793 (I50805,I50382);
nor I_2794 (I50823,I50805,I50409);
nand I_2795 (I50841,I50823,I50499);
nor I_2796 (I50859,I50841,I50787);
DFFARX1 I_2797 (I50859,I515,I50625,I50886,);
not I_2798 (I50895,I50841);
not I_2799 (I50913,I50409);
nand I_2800 (I50931,I50913,I50157);
nor I_2801 (I50949,I50409,I50076);
nand I_2802 (I50967,I50751,I50949);
nand I_2803 (I50985,I50697,I50409);
nand I_2804 (I51003,I50805,I50589);
DFFARX1 I_2805 (I51003,I515,I50625,I51030,);
DFFARX1 I_2806 (I51003,I515,I50625,I51048,);
not I_2807 (I51057,I50589);
nor I_2808 (I51075,I51057,I50607);
and I_2809 (I51093,I51075,I50193);
or I_2810 (I51111,I51093,I50157);
DFFARX1 I_2811 (I51111,I515,I50625,I51138,);
nand I_2812 (I51147,I51138,I50769);
nor I_2813 (I51165,I51147,I50931);
nor I_2814 (I51183,I51138,I50733);
DFFARX1 I_2815 (I51138,I515,I50625,I51210,);
not I_2816 (I51219,I51210);
nor I_2817 (I51237,I51219,I50895);
not I_2818 (I51255,I522);
DFFARX1 I_2819 (I50886,I515,I51255,I51282,);
not I_2820 (I51291,I51282);
nand I_2821 (I51309,I51183,I50679);
and I_2822 (I51327,I51309,I50967);
DFFARX1 I_2823 (I51327,I515,I51255,I51354,);
not I_2824 (I51363,I51165);
DFFARX1 I_2825 (I50886,I515,I51255,I51390,);
not I_2826 (I51399,I51390);
nor I_2827 (I51417,I51399,I51291);
and I_2828 (I51435,I51417,I51165);
nor I_2829 (I51453,I51399,I51363);
nor I_2830 (I51471,I51354,I51453);
DFFARX1 I_2831 (I51237,I515,I51255,I51498,);
nor I_2832 (I51507,I51498,I51354);
not I_2833 (I51525,I51507);
not I_2834 (I51543,I51498);
nor I_2835 (I51561,I51543,I51435);
DFFARX1 I_2836 (I51561,I515,I51255,I51588,);
nand I_2837 (I51597,I51183,I50985);
and I_2838 (I51615,I51597,I51048);
DFFARX1 I_2839 (I51615,I515,I51255,I51642,);
nor I_2840 (I51651,I51642,I51498);
DFFARX1 I_2841 (I51651,I515,I51255,I51678,);
nand I_2842 (I51687,I51642,I51543);
nand I_2843 (I51705,I51525,I51687);
not I_2844 (I51723,I51642);
nor I_2845 (I51741,I51723,I51435);
DFFARX1 I_2846 (I51741,I515,I51255,I51768,);
nor I_2847 (I51777,I51030,I50985);
or I_2848 (I51795,I51498,I51777);
nor I_2849 (I51813,I51642,I51777);
or I_2850 (I51831,I51354,I51777);
DFFARX1 I_2851 (I51777,I515,I51255,I51858,);
not I_2852 (I51867,I522);
DFFARX1 I_2853 (I51831,I515,I51867,I51894,);
DFFARX1 I_2854 (I51894,I515,I51867,I51912,);
not I_2855 (I51921,I51912);
nand I_2856 (I51939,I51768,I51858);
and I_2857 (I51957,I51939,I51813);
DFFARX1 I_2858 (I51957,I515,I51867,I51984,);
DFFARX1 I_2859 (I51984,I515,I51867,I52002,);
DFFARX1 I_2860 (I51984,I515,I51867,I52020,);
DFFARX1 I_2861 (I51705,I515,I51867,I52038,);
nand I_2862 (I52047,I52038,I51471);
not I_2863 (I52065,I52047);
nor I_2864 (I52083,I51894,I52065);
DFFARX1 I_2865 (I51813,I515,I51867,I52110,);
not I_2866 (I52119,I52110);
nor I_2867 (I52137,I52119,I51921);
nand I_2868 (I52155,I52119,I52047);
nand I_2869 (I52173,I51588,I51678);
and I_2870 (I52191,I52173,I51795);
DFFARX1 I_2871 (I52191,I515,I51867,I52218,);
nor I_2872 (I52227,I52218,I51894);
DFFARX1 I_2873 (I52227,I515,I51867,I52254,);
not I_2874 (I52263,I52218);
nor I_2875 (I52281,I51678,I51678);
not I_2876 (I52299,I52281);
nor I_2877 (I52317,I52047,I52299);
nor I_2878 (I52335,I52263,I52317);
DFFARX1 I_2879 (I52335,I515,I51867,I52362,);
nor I_2880 (I52371,I52218,I52299);
nor I_2881 (I52389,I52065,I52371);
nor I_2882 (I52407,I52218,I52281);
not I_2883 (I52425,I522);
DFFARX1 I_2884 (I52155,I515,I52425,I52452,);
nand I_2885 (I52461,I52452,I52254);
not I_2886 (I52479,I52461);
DFFARX1 I_2887 (I52137,I515,I52425,I52506,);
not I_2888 (I52515,I52506);
not I_2889 (I52533,I52362);
or I_2890 (I52551,I52020,I52362);
nor I_2891 (I52569,I52020,I52362);
or I_2892 (I52587,I52389,I52020);
DFFARX1 I_2893 (I52587,I515,I52425,I52614,);
not I_2894 (I52623,I52083);
nand I_2895 (I52641,I52623,I52002);
nand I_2896 (I52659,I52533,I52641);
and I_2897 (I52677,I52515,I52659);
nor I_2898 (I52695,I52083,I52407);
and I_2899 (I52713,I52515,I52695);
nor I_2900 (I52731,I52479,I52713);
DFFARX1 I_2901 (I52695,I515,I52425,I52758,);
not I_2902 (I52767,I52758);
nor I_2903 (I52785,I52515,I52767);
or I_2904 (I52803,I52587,I52407);
nor I_2905 (I52821,I52407,I52389);
nand I_2906 (I52839,I52659,I52821);
nand I_2907 (I52857,I52803,I52839);
DFFARX1 I_2908 (I52857,I515,I52425,I52884,);
nor I_2909 (I52893,I52821,I52551);
DFFARX1 I_2910 (I52893,I515,I52425,I52920,);
nor I_2911 (I52929,I52407,I52254);
DFFARX1 I_2912 (I52929,I515,I52425,I52956,);
DFFARX1 I_2913 (I52956,I515,I52425,I52974,);
not I_2914 (I52983,I52956);
nand I_2915 (I53001,I52983,I52461);
nand I_2916 (I53019,I52983,I52569);
not I_2917 (I53037,I522);
DFFARX1 I_2918 (I428,I515,I53037,I53064,);
nand I_2919 (I53073,I53064,I204);
DFFARX1 I_2920 (I132,I515,I53037,I53100,);
DFFARX1 I_2921 (I53100,I515,I53037,I53118,);
not I_2922 (I53127,I53118);
not I_2923 (I53145,I212);
nor I_2924 (I53163,I212,I244);
not I_2925 (I53181,I236);
nand I_2926 (I53199,I53145,I53181);
nor I_2927 (I53217,I236,I212);
and I_2928 (I53235,I53217,I53073);
not I_2929 (I53253,I364);
nand I_2930 (I53271,I53253,I452);
nor I_2931 (I53289,I364,I284);
not I_2932 (I53307,I53289);
nand I_2933 (I53325,I53163,I53307);
DFFARX1 I_2934 (I53289,I515,I53037,I53352,);
nor I_2935 (I53361,I100,I236);
nor I_2936 (I53379,I53361,I244);
and I_2937 (I53397,I53379,I53271);
DFFARX1 I_2938 (I53397,I515,I53037,I53424,);
nor I_2939 (I53433,I53361,I53199);
or I_2940 (I53451,I53289,I53361);
nor I_2941 (I53469,I100,I164);
DFFARX1 I_2942 (I53469,I515,I53037,I53496,);
not I_2943 (I53505,I53496);
nand I_2944 (I53523,I53505,I53145);
nor I_2945 (I53541,I53523,I244);
DFFARX1 I_2946 (I53541,I515,I53037,I53568,);
nor I_2947 (I53577,I53505,I53199);
nor I_2948 (I53595,I53361,I53577);
not I_2949 (I53613,I522);
DFFARX1 I_2950 (I53325,I515,I53613,I53640,);
not I_2951 (I53649,I53640);
nand I_2952 (I53667,I53568,I53352);
and I_2953 (I53685,I53667,I53451);
DFFARX1 I_2954 (I53685,I515,I53613,I53712,);
DFFARX1 I_2955 (I53235,I515,I53613,I53730,);
and I_2956 (I53739,I53730,I53433);
nor I_2957 (I53757,I53712,I53739);
DFFARX1 I_2958 (I53757,I515,I53613,I53784,);
nand I_2959 (I53793,I53730,I53433);
nand I_2960 (I53811,I53649,I53793);
not I_2961 (I53829,I53811);
DFFARX1 I_2962 (I53235,I515,I53613,I53856,);
DFFARX1 I_2963 (I53856,I515,I53613,I53874,);
nand I_2964 (I53883,I53127,I53595);
and I_2965 (I53901,I53883,I53568);
DFFARX1 I_2966 (I53901,I515,I53613,I53928,);
DFFARX1 I_2967 (I53928,I515,I53613,I53946,);
not I_2968 (I53955,I53946);
not I_2969 (I53973,I53928);
nand I_2970 (I53991,I53973,I53793);
nor I_2971 (I54009,I53424,I53595);
not I_2972 (I54027,I54009);
nor I_2973 (I54045,I53973,I54027);
nor I_2974 (I54063,I53649,I54045);
DFFARX1 I_2975 (I54063,I515,I53613,I54090,);
nor I_2976 (I54099,I53712,I54027);
nor I_2977 (I54117,I53928,I54099);
nor I_2978 (I54135,I53856,I54009);
nor I_2979 (I54153,I53712,I54009);
not I_2980 (I54171,I522);
DFFARX1 I_2981 (I54153,I515,I54171,I54198,);
not I_2982 (I54207,I54198);
nand I_2983 (I54225,I53829,I53874);
and I_2984 (I54243,I54225,I53784);
DFFARX1 I_2985 (I54243,I515,I54171,I54270,);
not I_2986 (I54279,I54153);
DFFARX1 I_2987 (I54090,I515,I54171,I54306,);
not I_2988 (I54315,I54306);
nor I_2989 (I54333,I54315,I54207);
and I_2990 (I54351,I54333,I54153);
nor I_2991 (I54369,I54315,I54279);
nor I_2992 (I54387,I54270,I54369);
DFFARX1 I_2993 (I53991,I515,I54171,I54414,);
nor I_2994 (I54423,I54414,I54270);
not I_2995 (I54441,I54423);
not I_2996 (I54459,I54414);
nor I_2997 (I54477,I54459,I54351);
DFFARX1 I_2998 (I54477,I515,I54171,I54504,);
nand I_2999 (I54513,I53955,I53784);
and I_3000 (I54531,I54513,I54117);
DFFARX1 I_3001 (I54531,I515,I54171,I54558,);
nor I_3002 (I54567,I54558,I54414);
DFFARX1 I_3003 (I54567,I515,I54171,I54594,);
nand I_3004 (I54603,I54558,I54459);
nand I_3005 (I54621,I54441,I54603);
not I_3006 (I54639,I54558);
nor I_3007 (I54657,I54639,I54351);
DFFARX1 I_3008 (I54657,I515,I54171,I54684,);
nor I_3009 (I54693,I54135,I53784);
or I_3010 (I54711,I54414,I54693);
nor I_3011 (I54729,I54558,I54693);
or I_3012 (I54747,I54270,I54693);
DFFARX1 I_3013 (I54693,I515,I54171,I54774,);
not I_3014 (I54783,I522);
DFFARX1 I_3015 (I54747,I515,I54783,I54810,);
DFFARX1 I_3016 (I54594,I515,I54783,I54828,);
not I_3017 (I54837,I54828);
not I_3018 (I54855,I54387);
nor I_3019 (I54873,I54855,I54594);
not I_3020 (I54891,I54621);
nor I_3021 (I54909,I54873,I54504);
nor I_3022 (I54927,I54828,I54909);
DFFARX1 I_3023 (I54927,I515,I54783,I54954,);
nor I_3024 (I54963,I54504,I54594);
nand I_3025 (I54981,I54963,I54387);
DFFARX1 I_3026 (I54981,I515,I54783,I55008,);
nor I_3027 (I55017,I54891,I54504);
nand I_3028 (I55035,I55017,I54729);
nor I_3029 (I55053,I54810,I55035);
DFFARX1 I_3030 (I55053,I515,I54783,I55080,);
not I_3031 (I55089,I55035);
nand I_3032 (I55107,I54828,I55089);
DFFARX1 I_3033 (I55035,I515,I54783,I55134,);
not I_3034 (I55143,I55134);
not I_3035 (I55161,I54504);
not I_3036 (I55179,I54711);
nor I_3037 (I55197,I55179,I54621);
nor I_3038 (I55215,I55143,I55197);
nor I_3039 (I55233,I55179,I54684);
and I_3040 (I55251,I55233,I54774);
or I_3041 (I55269,I55251,I54729);
DFFARX1 I_3042 (I55269,I515,I54783,I55296,);
nor I_3043 (I55305,I55296,I54810);
not I_3044 (I55323,I55296);
and I_3045 (I55341,I55323,I54810);
nor I_3046 (I55359,I54837,I55341);
nand I_3047 (I55377,I55323,I54891);
nor I_3048 (I55395,I55179,I55377);
nand I_3049 (I55413,I55323,I55089);
nand I_3050 (I55431,I54891,I54711);
nor I_3051 (I55449,I55161,I55431);
not I_3052 (I55467,I522);
DFFARX1 I_3053 (I55305,I515,I55467,I55494,);
DFFARX1 I_3054 (I55494,I515,I55467,I55512,);
not I_3055 (I55521,I55512);
not I_3056 (I55539,I55494);
DFFARX1 I_3057 (I55008,I515,I55467,I55566,);
not I_3058 (I55575,I55566);
and I_3059 (I55593,I55539,I55107);
not I_3060 (I55611,I55395);
nand I_3061 (I55629,I55611,I55107);
not I_3062 (I55647,I55359);
nor I_3063 (I55665,I55647,I55215);
nand I_3064 (I55683,I55665,I55080);
nor I_3065 (I55701,I55683,I55629);
DFFARX1 I_3066 (I55701,I515,I55467,I55728,);
not I_3067 (I55737,I55683);
not I_3068 (I55755,I55215);
nand I_3069 (I55773,I55755,I55107);
nor I_3070 (I55791,I55215,I55395);
nand I_3071 (I55809,I55593,I55791);
nand I_3072 (I55827,I55539,I55215);
nand I_3073 (I55845,I55647,I55413);
DFFARX1 I_3074 (I55845,I515,I55467,I55872,);
DFFARX1 I_3075 (I55845,I515,I55467,I55890,);
not I_3076 (I55899,I55413);
nor I_3077 (I55917,I55899,I55449);
and I_3078 (I55935,I55917,I55080);
or I_3079 (I55953,I55935,I54954);
DFFARX1 I_3080 (I55953,I515,I55467,I55980,);
nand I_3081 (I55989,I55980,I55611);
nor I_3082 (I56007,I55989,I55773);
nor I_3083 (I56025,I55980,I55575);
DFFARX1 I_3084 (I55980,I515,I55467,I56052,);
not I_3085 (I56061,I56052);
nor I_3086 (I56079,I56061,I55737);
not I_3087 (I56097,I522);
DFFARX1 I_3088 (I55728,I515,I56097,I56124,);
DFFARX1 I_3089 (I56124,I515,I56097,I56142,);
not I_3090 (I56151,I56142);
DFFARX1 I_3091 (I55521,I515,I56097,I56178,);
not I_3092 (I56187,I56079);
nor I_3093 (I56205,I56124,I56187);
not I_3094 (I56223,I55809);
not I_3095 (I56241,I56007);
nand I_3096 (I56259,I56241,I55809);
nor I_3097 (I56277,I56187,I56259);
nor I_3098 (I56295,I56178,I56277);
DFFARX1 I_3099 (I56241,I515,I56097,I56322,);
nor I_3100 (I56331,I56007,I56025);
nand I_3101 (I56349,I56331,I55872);
nor I_3102 (I56367,I56349,I56223);
nand I_3103 (I56385,I56367,I56079);
DFFARX1 I_3104 (I56349,I515,I56097,I56412,);
nand I_3105 (I56421,I56223,I56007);
nor I_3106 (I56439,I56223,I56007);
nand I_3107 (I56457,I56205,I56439);
not I_3108 (I56475,I55890);
nor I_3109 (I56493,I56475,I56421);
DFFARX1 I_3110 (I56493,I515,I56097,I56520,);
nor I_3111 (I56529,I56475,I55728);
and I_3112 (I56547,I56529,I55827);
or I_3113 (I56565,I56547,I56025);
DFFARX1 I_3114 (I56565,I515,I56097,I56592,);
nor I_3115 (I56601,I56592,I56178);
nor I_3116 (I56619,I56124,I56601);
not I_3117 (I56637,I56592);
nor I_3118 (I56655,I56637,I56295);
DFFARX1 I_3119 (I56655,I515,I56097,I56682,);
nand I_3120 (I56691,I56637,I56223);
nor I_3121 (I56709,I56475,I56691);
not I_3122 (I56727,I522);
DFFARX1 I_3123 (I56520,I515,I56727,I56754,);
not I_3124 (I56763,I56754);
nand I_3125 (I56781,I56682,I56520);
and I_3126 (I56799,I56781,I56709);
DFFARX1 I_3127 (I56799,I515,I56727,I56826,);
not I_3128 (I56835,I56709);
DFFARX1 I_3129 (I56457,I515,I56727,I56862,);
not I_3130 (I56871,I56862);
nor I_3131 (I56889,I56871,I56763);
and I_3132 (I56907,I56889,I56709);
nor I_3133 (I56925,I56871,I56835);
nor I_3134 (I56943,I56826,I56925);
DFFARX1 I_3135 (I56385,I515,I56727,I56970,);
nor I_3136 (I56979,I56970,I56826);
not I_3137 (I56997,I56979);
not I_3138 (I57015,I56970);
nor I_3139 (I57033,I57015,I56907);
DFFARX1 I_3140 (I57033,I515,I56727,I57060,);
nand I_3141 (I57069,I56619,I56412);
and I_3142 (I57087,I57069,I56151);
DFFARX1 I_3143 (I57087,I515,I56727,I57114,);
nor I_3144 (I57123,I57114,I56970);
DFFARX1 I_3145 (I57123,I515,I56727,I57150,);
nand I_3146 (I57159,I57114,I57015);
nand I_3147 (I57177,I56997,I57159);
not I_3148 (I57195,I57114);
nor I_3149 (I57213,I57195,I56907);
DFFARX1 I_3150 (I57213,I515,I56727,I57240,);
nor I_3151 (I57249,I56322,I56412);
or I_3152 (I57267,I56970,I57249);
nor I_3153 (I57285,I57114,I57249);
or I_3154 (I57303,I56826,I57249);
DFFARX1 I_3155 (I57249,I515,I56727,I57330,);
not I_3156 (I57339,I522);
DFFARX1 I_3157 (I57267,I515,I57339,I57366,);
nand I_3158 (I57375,I57285,I57060);
and I_3159 (I57393,I57375,I57330);
DFFARX1 I_3160 (I57393,I515,I57339,I57420,);
nor I_3161 (I57429,I57420,I57366);
not I_3162 (I57447,I57420);
DFFARX1 I_3163 (I57177,I515,I57339,I57474,);
nand I_3164 (I57483,I57474,I57285);
not I_3165 (I57501,I57483);
DFFARX1 I_3166 (I57501,I515,I57339,I57528,);
not I_3167 (I57537,I57528);
nor I_3168 (I57555,I57366,I57483);
nor I_3169 (I57573,I57420,I57555);
DFFARX1 I_3170 (I57303,I515,I57339,I57600,);
DFFARX1 I_3171 (I57600,I515,I57339,I57618,);
not I_3172 (I57627,I57618);
not I_3173 (I57645,I57600);
nand I_3174 (I57663,I57645,I57447);
nand I_3175 (I57681,I57150,I56943);
and I_3176 (I57699,I57681,I57150);
DFFARX1 I_3177 (I57699,I515,I57339,I57726,);
nor I_3178 (I57735,I57726,I57366);
DFFARX1 I_3179 (I57735,I515,I57339,I57762,);
DFFARX1 I_3180 (I57726,I515,I57339,I57780,);
nor I_3181 (I57789,I57240,I56943);
not I_3182 (I57807,I57789);
nor I_3183 (I57825,I57627,I57807);
nand I_3184 (I57843,I57645,I57807);
nor I_3185 (I57861,I57366,I57789);
DFFARX1 I_3186 (I57789,I515,I57339,I57888,);
not I_3187 (I57897,I522);
DFFARX1 I_3188 (I57843,I515,I57897,I57924,);
not I_3189 (I57933,I57924);
DFFARX1 I_3190 (I57825,I515,I57897,I57960,);
not I_3191 (I57969,I57888);
nand I_3192 (I57987,I57969,I57429);
not I_3193 (I58005,I57987);
nor I_3194 (I58023,I58005,I57537);
nor I_3195 (I58041,I57933,I58023);
DFFARX1 I_3196 (I58041,I515,I57897,I58068,);
not I_3197 (I58077,I57537);
nand I_3198 (I58095,I58077,I58005);
and I_3199 (I58113,I58077,I57573);
nand I_3200 (I58131,I58113,I57762);
nor I_3201 (I58149,I58131,I58077);
and I_3202 (I58167,I57960,I58131);
not I_3203 (I58185,I58131);
nand I_3204 (I58203,I57960,I58185);
nor I_3205 (I58221,I57924,I58131);
not I_3206 (I58239,I57762);
nor I_3207 (I58257,I58239,I57573);
nand I_3208 (I58275,I58257,I58077);
nor I_3209 (I58293,I57987,I58275);
nor I_3210 (I58311,I58239,I57861);
and I_3211 (I58329,I58311,I57780);
or I_3212 (I58347,I58329,I57663);
DFFARX1 I_3213 (I58347,I515,I57897,I58374,);
nor I_3214 (I58383,I58374,I58095);
DFFARX1 I_3215 (I58383,I515,I57897,I58410,);
DFFARX1 I_3216 (I58374,I515,I57897,I58428,);
not I_3217 (I58437,I58374);
nor I_3218 (I58455,I58437,I57960);
nor I_3219 (I58473,I58257,I58455);
DFFARX1 I_3220 (I58473,I515,I57897,I58500,);
not I_3221 (I58509,I522);
DFFARX1 I_3222 (I58221,I515,I58509,I58536,);
DFFARX1 I_3223 (I58536,I515,I58509,I58554,);
not I_3224 (I58563,I58554);
not I_3225 (I58581,I58536);
nand I_3226 (I58599,I58410,I58500);
and I_3227 (I58617,I58599,I58428);
DFFARX1 I_3228 (I58617,I515,I58509,I58644,);
not I_3229 (I58653,I58644);
DFFARX1 I_3230 (I58203,I515,I58509,I58680,);
and I_3231 (I58689,I58680,I58293);
nand I_3232 (I58707,I58680,I58293);
nand I_3233 (I58725,I58653,I58707);
DFFARX1 I_3234 (I58149,I515,I58509,I58752,);
nor I_3235 (I58761,I58752,I58689);
DFFARX1 I_3236 (I58761,I515,I58509,I58788,);
nor I_3237 (I58797,I58752,I58644);
nand I_3238 (I58815,I58410,I58167);
and I_3239 (I58833,I58815,I58068);
DFFARX1 I_3240 (I58833,I515,I58509,I58860,);
nor I_3241 (I58869,I58860,I58752);
not I_3242 (I58887,I58860);
nor I_3243 (I58905,I58887,I58653);
nor I_3244 (I58923,I58581,I58905);
DFFARX1 I_3245 (I58923,I515,I58509,I58950,);
nor I_3246 (I58959,I58887,I58752);
nor I_3247 (I58977,I58221,I58167);
nor I_3248 (I58995,I58977,I58959);
not I_3249 (I59013,I58977);
nand I_3250 (I59031,I58707,I59013);
DFFARX1 I_3251 (I58977,I515,I58509,I59058,);
DFFARX1 I_3252 (I58977,I515,I58509,I59076,);
not I_3253 (I59085,I522);
DFFARX1 I_3254 (I59058,I515,I59085,I59112,);
nand I_3255 (I59121,I59112,I59076);
DFFARX1 I_3256 (I58788,I515,I59085,I59148,);
DFFARX1 I_3257 (I59148,I515,I59085,I59166,);
not I_3258 (I59175,I59166);
not I_3259 (I59193,I58797);
nor I_3260 (I59211,I58797,I58950);
not I_3261 (I59229,I58995);
nand I_3262 (I59247,I59193,I59229);
nor I_3263 (I59265,I58995,I58797);
and I_3264 (I59283,I59265,I59121);
not I_3265 (I59301,I58725);
nand I_3266 (I59319,I59301,I58563);
nor I_3267 (I59337,I58725,I58869);
not I_3268 (I59355,I59337);
nand I_3269 (I59373,I59211,I59355);
DFFARX1 I_3270 (I59337,I515,I59085,I59400,);
nor I_3271 (I59409,I59031,I58995);
nor I_3272 (I59427,I59409,I58950);
and I_3273 (I59445,I59427,I59319);
DFFARX1 I_3274 (I59445,I515,I59085,I59472,);
nor I_3275 (I59481,I59409,I59247);
or I_3276 (I59499,I59337,I59409);
nor I_3277 (I59517,I59031,I58788);
DFFARX1 I_3278 (I59517,I515,I59085,I59544,);
not I_3279 (I59553,I59544);
nand I_3280 (I59571,I59553,I59193);
nor I_3281 (I59589,I59571,I58950);
DFFARX1 I_3282 (I59589,I515,I59085,I59616,);
nor I_3283 (I59625,I59553,I59247);
nor I_3284 (I59643,I59409,I59625);
not I_3285 (I59661,I522);
DFFARX1 I_3286 (I59472,I515,I59661,I59688,);
DFFARX1 I_3287 (I59688,I515,I59661,I59706,);
not I_3288 (I59715,I59706);
not I_3289 (I59733,I59688);
DFFARX1 I_3290 (I59283,I515,I59661,I59760,);
not I_3291 (I59769,I59760);
and I_3292 (I59787,I59733,I59400);
not I_3293 (I59805,I59283);
nand I_3294 (I59823,I59805,I59400);
not I_3295 (I59841,I59175);
nor I_3296 (I59859,I59841,I59481);
nand I_3297 (I59877,I59859,I59499);
nor I_3298 (I59895,I59877,I59823);
DFFARX1 I_3299 (I59895,I515,I59661,I59922,);
not I_3300 (I59931,I59877);
not I_3301 (I59949,I59481);
nand I_3302 (I59967,I59949,I59400);
nor I_3303 (I59985,I59481,I59283);
nand I_3304 (I60003,I59787,I59985);
nand I_3305 (I60021,I59733,I59481);
nand I_3306 (I60039,I59841,I59643);
DFFARX1 I_3307 (I60039,I515,I59661,I60066,);
DFFARX1 I_3308 (I60039,I515,I59661,I60084,);
not I_3309 (I60093,I59643);
nor I_3310 (I60111,I60093,I59616);
and I_3311 (I60129,I60111,I59373);
or I_3312 (I60147,I60129,I59616);
DFFARX1 I_3313 (I60147,I515,I59661,I60174,);
nand I_3314 (I60183,I60174,I59805);
nor I_3315 (I60201,I60183,I59967);
nor I_3316 (I60219,I60174,I59769);
DFFARX1 I_3317 (I60174,I515,I59661,I60246,);
not I_3318 (I60255,I60246);
nor I_3319 (I60273,I60255,I59931);
not I_3320 (I60291,I522);
DFFARX1 I_3321 (I60021,I515,I60291,I60318,);
not I_3322 (I60327,I60318);
nand I_3323 (I60345,I60219,I60066);
and I_3324 (I60363,I60345,I60003);
DFFARX1 I_3325 (I60363,I515,I60291,I60390,);
DFFARX1 I_3326 (I60390,I515,I60291,I60408,);
DFFARX1 I_3327 (I60273,I515,I60291,I60426,);
nand I_3328 (I60435,I60426,I60084);
not I_3329 (I60453,I60435);
DFFARX1 I_3330 (I60453,I515,I60291,I60480,);
not I_3331 (I60489,I60480);
nor I_3332 (I60507,I60327,I60489);
DFFARX1 I_3333 (I60201,I515,I60291,I60534,);
nor I_3334 (I60543,I60534,I60390);
nor I_3335 (I60561,I60534,I60453);
nand I_3336 (I60579,I59922,I59715);
and I_3337 (I60597,I60579,I60219);
DFFARX1 I_3338 (I60597,I515,I60291,I60624,);
not I_3339 (I60633,I60624);
nand I_3340 (I60651,I60633,I60534);
nand I_3341 (I60669,I60633,I60435);
nor I_3342 (I60687,I59922,I59715);
and I_3343 (I60705,I60534,I60687);
nor I_3344 (I60723,I60633,I60705);
DFFARX1 I_3345 (I60723,I515,I60291,I60750,);
nor I_3346 (I60759,I60318,I60687);
DFFARX1 I_3347 (I60759,I515,I60291,I60786,);
nor I_3348 (I60795,I60624,I60687);
not I_3349 (I60813,I60795);
nand I_3350 (I60831,I60813,I60651);
not I_3351 (I60849,I522);
DFFARX1 I_3352 (I60669,I515,I60849,I60876,);
not I_3353 (I60885,I60876);
DFFARX1 I_3354 (I60669,I515,I60849,I60912,);
not I_3355 (I60921,I60561);
nand I_3356 (I60939,I60921,I60408);
not I_3357 (I60957,I60939);
nor I_3358 (I60975,I60957,I60543);
nor I_3359 (I60993,I60885,I60975);
DFFARX1 I_3360 (I60993,I515,I60849,I61020,);
not I_3361 (I61029,I60543);
nand I_3362 (I61047,I61029,I60957);
and I_3363 (I61065,I61029,I60831);
nand I_3364 (I61083,I61065,I60786);
nor I_3365 (I61101,I61083,I61029);
and I_3366 (I61119,I60912,I61083);
not I_3367 (I61137,I61083);
nand I_3368 (I61155,I60912,I61137);
nor I_3369 (I61173,I60876,I61083);
not I_3370 (I61191,I60507);
nor I_3371 (I61209,I61191,I60831);
nand I_3372 (I61227,I61209,I61029);
nor I_3373 (I61245,I60939,I61227);
nor I_3374 (I61263,I61191,I60786);
and I_3375 (I61281,I61263,I60561);
or I_3376 (I61299,I61281,I60750);
DFFARX1 I_3377 (I61299,I515,I60849,I61326,);
nor I_3378 (I61335,I61326,I61047);
DFFARX1 I_3379 (I61335,I515,I60849,I61362,);
DFFARX1 I_3380 (I61326,I515,I60849,I61380,);
not I_3381 (I61389,I61326);
nor I_3382 (I61407,I61389,I60912);
nor I_3383 (I61425,I61209,I61407);
DFFARX1 I_3384 (I61425,I515,I60849,I61452,);
not I_3385 (I61461,I522);
DFFARX1 I_3386 (I61155,I515,I61461,I61488,);
not I_3387 (I61497,I61488);
nand I_3388 (I61515,I61452,I61119);
and I_3389 (I61533,I61515,I61362);
DFFARX1 I_3390 (I61533,I515,I61461,I61560,);
DFFARX1 I_3391 (I61101,I515,I61461,I61578,);
and I_3392 (I61587,I61578,I61173);
nor I_3393 (I61605,I61560,I61587);
DFFARX1 I_3394 (I61605,I515,I61461,I61632,);
nand I_3395 (I61641,I61578,I61173);
nand I_3396 (I61659,I61497,I61641);
not I_3397 (I61677,I61659);
DFFARX1 I_3398 (I61245,I515,I61461,I61704,);
DFFARX1 I_3399 (I61704,I515,I61461,I61722,);
nand I_3400 (I61731,I61020,I61380);
and I_3401 (I61749,I61731,I61362);
DFFARX1 I_3402 (I61749,I515,I61461,I61776,);
DFFARX1 I_3403 (I61776,I515,I61461,I61794,);
not I_3404 (I61803,I61794);
not I_3405 (I61821,I61776);
nand I_3406 (I61839,I61821,I61641);
nor I_3407 (I61857,I61173,I61380);
not I_3408 (I61875,I61857);
nor I_3409 (I61893,I61821,I61875);
nor I_3410 (I61911,I61497,I61893);
DFFARX1 I_3411 (I61911,I515,I61461,I61938,);
nor I_3412 (I61947,I61560,I61875);
nor I_3413 (I61965,I61776,I61947);
nor I_3414 (I61983,I61704,I61857);
nor I_3415 (I62001,I61560,I61857);
not I_3416 (I62019,I522);
DFFARX1 I_3417 (I61839,I515,I62019,I62046,);
DFFARX1 I_3418 (I62046,I515,I62019,I62064,);
not I_3419 (I62073,I62064);
not I_3420 (I62091,I62046);
DFFARX1 I_3421 (I62001,I515,I62019,I62118,);
not I_3422 (I62127,I62118);
and I_3423 (I62145,I62091,I61632);
not I_3424 (I62163,I61722);
nand I_3425 (I62181,I62163,I61632);
not I_3426 (I62199,I61983);
nor I_3427 (I62217,I62199,I61965);
nand I_3428 (I62235,I62217,I61677);
nor I_3429 (I62253,I62235,I62181);
DFFARX1 I_3430 (I62253,I515,I62019,I62280,);
not I_3431 (I62289,I62235);
not I_3432 (I62307,I61965);
nand I_3433 (I62325,I62307,I61632);
nor I_3434 (I62343,I61965,I61722);
nand I_3435 (I62361,I62145,I62343);
nand I_3436 (I62379,I62091,I61965);
nand I_3437 (I62397,I62199,I61632);
DFFARX1 I_3438 (I62397,I515,I62019,I62424,);
DFFARX1 I_3439 (I62397,I515,I62019,I62442,);
not I_3440 (I62451,I61632);
nor I_3441 (I62469,I62451,I61938);
and I_3442 (I62487,I62469,I61803);
or I_3443 (I62505,I62487,I62001);
DFFARX1 I_3444 (I62505,I515,I62019,I62532,);
nand I_3445 (I62541,I62532,I62163);
nor I_3446 (I62559,I62541,I62325);
nor I_3447 (I62577,I62532,I62127);
DFFARX1 I_3448 (I62532,I515,I62019,I62604,);
not I_3449 (I62613,I62604);
nor I_3450 (I62631,I62613,I62289);
not I_3451 (I62649,I522);
DFFARX1 I_3452 (I62559,I515,I62649,I62676,);
nand I_3453 (I62685,I62676,I62073);
DFFARX1 I_3454 (I62442,I515,I62649,I62712,);
DFFARX1 I_3455 (I62712,I515,I62649,I62730,);
not I_3456 (I62739,I62730);
not I_3457 (I62757,I62280);
nor I_3458 (I62775,I62280,I62379);
not I_3459 (I62793,I62361);
nand I_3460 (I62811,I62757,I62793);
nor I_3461 (I62829,I62361,I62280);
and I_3462 (I62847,I62829,I62685);
not I_3463 (I62865,I62631);
nand I_3464 (I62883,I62865,I62280);
nor I_3465 (I62901,I62631,I62577);
not I_3466 (I62919,I62901);
nand I_3467 (I62937,I62775,I62919);
DFFARX1 I_3468 (I62901,I515,I62649,I62964,);
nor I_3469 (I62973,I62577,I62361);
nor I_3470 (I62991,I62973,I62379);
and I_3471 (I63009,I62991,I62883);
DFFARX1 I_3472 (I63009,I515,I62649,I63036,);
nor I_3473 (I63045,I62973,I62811);
or I_3474 (I63063,I62901,I62973);
nor I_3475 (I63081,I62577,I62424);
DFFARX1 I_3476 (I63081,I515,I62649,I63108,);
not I_3477 (I63117,I63108);
nand I_3478 (I63135,I63117,I62757);
nor I_3479 (I63153,I63135,I62379);
DFFARX1 I_3480 (I63153,I515,I62649,I63180,);
nor I_3481 (I63189,I63117,I62811);
nor I_3482 (I63207,I62973,I63189);
not I_3483 (I63225,I522);
DFFARX1 I_3484 (I63180,I515,I63225,I63252,);
not I_3485 (I63261,I63252);
nand I_3486 (I63279,I62847,I63063);
and I_3487 (I63297,I63279,I63045);
DFFARX1 I_3488 (I63297,I515,I63225,I63324,);
not I_3489 (I63333,I62739);
DFFARX1 I_3490 (I62937,I515,I63225,I63360,);
not I_3491 (I63369,I63360);
nor I_3492 (I63387,I63369,I63261);
and I_3493 (I63405,I63387,I62739);
nor I_3494 (I63423,I63369,I63333);
nor I_3495 (I63441,I63324,I63423);
DFFARX1 I_3496 (I62847,I515,I63225,I63468,);
nor I_3497 (I63477,I63468,I63324);
not I_3498 (I63495,I63477);
not I_3499 (I63513,I63468);
nor I_3500 (I63531,I63513,I63405);
DFFARX1 I_3501 (I63531,I515,I63225,I63558,);
nand I_3502 (I63567,I62964,I63180);
and I_3503 (I63585,I63567,I63036);
DFFARX1 I_3504 (I63585,I515,I63225,I63612,);
nor I_3505 (I63621,I63612,I63468);
DFFARX1 I_3506 (I63621,I515,I63225,I63648,);
nand I_3507 (I63657,I63612,I63513);
nand I_3508 (I63675,I63495,I63657);
not I_3509 (I63693,I63612);
nor I_3510 (I63711,I63693,I63405);
DFFARX1 I_3511 (I63711,I515,I63225,I63738,);
nor I_3512 (I63747,I63207,I63180);
or I_3513 (I63765,I63468,I63747);
nor I_3514 (I63783,I63612,I63747);
or I_3515 (I63801,I63324,I63747);
DFFARX1 I_3516 (I63747,I515,I63225,I63828,);
not I_3517 (I63837,I522);
DFFARX1 I_3518 (I63765,I515,I63837,I63864,);
nand I_3519 (I63873,I63783,I63558);
and I_3520 (I63891,I63873,I63828);
DFFARX1 I_3521 (I63891,I515,I63837,I63918,);
nor I_3522 (I63927,I63918,I63864);
not I_3523 (I63945,I63918);
DFFARX1 I_3524 (I63675,I515,I63837,I63972,);
nand I_3525 (I63981,I63972,I63783);
not I_3526 (I63999,I63981);
DFFARX1 I_3527 (I63999,I515,I63837,I64026,);
not I_3528 (I64035,I64026);
nor I_3529 (I64053,I63864,I63981);
nor I_3530 (I64071,I63918,I64053);
DFFARX1 I_3531 (I63801,I515,I63837,I64098,);
DFFARX1 I_3532 (I64098,I515,I63837,I64116,);
not I_3533 (I64125,I64116);
not I_3534 (I64143,I64098);
nand I_3535 (I64161,I64143,I63945);
nand I_3536 (I64179,I63648,I63441);
and I_3537 (I64197,I64179,I63648);
DFFARX1 I_3538 (I64197,I515,I63837,I64224,);
nor I_3539 (I64233,I64224,I63864);
DFFARX1 I_3540 (I64233,I515,I63837,I64260,);
DFFARX1 I_3541 (I64224,I515,I63837,I64278,);
nor I_3542 (I64287,I63738,I63441);
not I_3543 (I64305,I64287);
nor I_3544 (I64323,I64125,I64305);
nand I_3545 (I64341,I64143,I64305);
nor I_3546 (I64359,I63864,I64287);
DFFARX1 I_3547 (I64287,I515,I63837,I64386,);
not I_3548 (I64395,I522);
DFFARX1 I_3549 (I64323,I515,I64395,I64422,);
DFFARX1 I_3550 (I64422,I515,I64395,I64440,);
not I_3551 (I64449,I64440);
not I_3552 (I64467,I64422);
DFFARX1 I_3553 (I64278,I515,I64395,I64494,);
nand I_3554 (I64503,I64494,I64161);
not I_3555 (I64521,I64161);
not I_3556 (I64539,I64071);
nand I_3557 (I64557,I63927,I64260);
and I_3558 (I64575,I63927,I64260);
not I_3559 (I64593,I64359);
nand I_3560 (I64611,I64593,I64539);
nor I_3561 (I64629,I64611,I64503);
nor I_3562 (I64647,I64521,I64611);
nand I_3563 (I64665,I64575,I64647);
not I_3564 (I64683,I64035);
nor I_3565 (I64701,I64683,I63927);
nor I_3566 (I64719,I64701,I64359);
nor I_3567 (I64737,I64467,I64719);
DFFARX1 I_3568 (I64737,I515,I64395,I64764,);
not I_3569 (I64773,I64701);
DFFARX1 I_3570 (I64773,I515,I64395,I64800,);
and I_3571 (I64809,I64494,I64701);
nor I_3572 (I64827,I64683,I64386);
and I_3573 (I64845,I64827,I64260);
or I_3574 (I64863,I64845,I64341);
DFFARX1 I_3575 (I64863,I515,I64395,I64890,);
nor I_3576 (I64899,I64890,I64593);
DFFARX1 I_3577 (I64899,I515,I64395,I64926,);
nand I_3578 (I64935,I64890,I64494);
nand I_3579 (I64953,I64593,I64935);
nor I_3580 (I64971,I64953,I64557);
not I_3581 (I64989,I522);
DFFARX1 I_3582 (I64971,I515,I64989,I65016,);
not I_3583 (I65025,I65016);
nand I_3584 (I65043,I64800,I64665);
and I_3585 (I65061,I65043,I64629);
DFFARX1 I_3586 (I65061,I515,I64989,I65088,);
DFFARX1 I_3587 (I65088,I515,I64989,I65106,);
DFFARX1 I_3588 (I64629,I515,I64989,I65124,);
nand I_3589 (I65133,I65124,I64926);
not I_3590 (I65151,I65133);
DFFARX1 I_3591 (I65151,I515,I64989,I65178,);
not I_3592 (I65187,I65178);
nor I_3593 (I65205,I65025,I65187);
DFFARX1 I_3594 (I64665,I515,I64989,I65232,);
nor I_3595 (I65241,I65232,I65088);
nor I_3596 (I65259,I65232,I65151);
nand I_3597 (I65277,I64449,I64809);
and I_3598 (I65295,I65277,I64764);
DFFARX1 I_3599 (I65295,I515,I64989,I65322,);
not I_3600 (I65331,I65322);
nand I_3601 (I65349,I65331,I65232);
nand I_3602 (I65367,I65331,I65133);
nor I_3603 (I65385,I64926,I64809);
and I_3604 (I65403,I65232,I65385);
nor I_3605 (I65421,I65331,I65403);
DFFARX1 I_3606 (I65421,I515,I64989,I65448,);
nor I_3607 (I65457,I65016,I65385);
DFFARX1 I_3608 (I65457,I515,I64989,I65484,);
nor I_3609 (I65493,I65322,I65385);
not I_3610 (I65511,I65493);
nand I_3611 (I65529,I65511,I65349);
not I_3612 (I65547,I522);
DFFARX1 I_3613 (I65529,I515,I65547,I65574,);
DFFARX1 I_3614 (I65574,I515,I65547,I65592,);
not I_3615 (I65601,I65592);
nand I_3616 (I65619,I65484,I65205);
and I_3617 (I65637,I65619,I65259);
DFFARX1 I_3618 (I65637,I515,I65547,I65664,);
DFFARX1 I_3619 (I65664,I515,I65547,I65682,);
DFFARX1 I_3620 (I65664,I515,I65547,I65700,);
DFFARX1 I_3621 (I65259,I515,I65547,I65718,);
nand I_3622 (I65727,I65718,I65106);
not I_3623 (I65745,I65727);
nor I_3624 (I65763,I65574,I65745);
DFFARX1 I_3625 (I65241,I515,I65547,I65790,);
not I_3626 (I65799,I65790);
nor I_3627 (I65817,I65799,I65601);
nand I_3628 (I65835,I65799,I65727);
nand I_3629 (I65853,I65367,I65448);
and I_3630 (I65871,I65853,I65484);
DFFARX1 I_3631 (I65871,I515,I65547,I65898,);
nor I_3632 (I65907,I65898,I65574);
DFFARX1 I_3633 (I65907,I515,I65547,I65934,);
not I_3634 (I65943,I65898);
nor I_3635 (I65961,I65367,I65448);
not I_3636 (I65979,I65961);
nor I_3637 (I65997,I65727,I65979);
nor I_3638 (I66015,I65943,I65997);
DFFARX1 I_3639 (I66015,I515,I65547,I66042,);
nor I_3640 (I66051,I65898,I65979);
nor I_3641 (I66069,I65745,I66051);
nor I_3642 (I66087,I65898,I65961);
not I_3643 (I66105,I522);
DFFARX1 I_3644 (I65934,I515,I66105,I66132,);
DFFARX1 I_3645 (I65835,I515,I66105,I66150,);
not I_3646 (I66159,I66150);
not I_3647 (I66177,I65934);
nor I_3648 (I66195,I66177,I65763);
not I_3649 (I66213,I65700);
nor I_3650 (I66231,I66195,I65817);
nor I_3651 (I66249,I66150,I66231);
DFFARX1 I_3652 (I66249,I515,I66105,I66276,);
nor I_3653 (I66285,I65817,I65763);
nand I_3654 (I66303,I66285,I65934);
DFFARX1 I_3655 (I66303,I515,I66105,I66330,);
nor I_3656 (I66339,I66213,I65817);
nand I_3657 (I66357,I66339,I66087);
nor I_3658 (I66375,I66132,I66357);
DFFARX1 I_3659 (I66375,I515,I66105,I66402,);
not I_3660 (I66411,I66357);
nand I_3661 (I66429,I66150,I66411);
DFFARX1 I_3662 (I66357,I515,I66105,I66456,);
not I_3663 (I66465,I66456);
not I_3664 (I66483,I65817);
not I_3665 (I66501,I66087);
nor I_3666 (I66519,I66501,I65700);
nor I_3667 (I66537,I66465,I66519);
nor I_3668 (I66555,I66501,I66042);
and I_3669 (I66573,I66555,I65682);
or I_3670 (I66591,I66573,I66069);
DFFARX1 I_3671 (I66591,I515,I66105,I66618,);
nor I_3672 (I66627,I66618,I66132);
not I_3673 (I66645,I66618);
and I_3674 (I66663,I66645,I66132);
nor I_3675 (I66681,I66159,I66663);
nand I_3676 (I66699,I66645,I66213);
nor I_3677 (I66717,I66501,I66699);
nand I_3678 (I66735,I66645,I66411);
nand I_3679 (I66753,I66213,I66087);
nor I_3680 (I66771,I66483,I66753);
not I_3681 (I66789,I522);
DFFARX1 I_3682 (I66627,I515,I66789,I66816,);
DFFARX1 I_3683 (I66816,I515,I66789,I66834,);
not I_3684 (I66843,I66834);
not I_3685 (I66861,I66816);
DFFARX1 I_3686 (I66330,I515,I66789,I66888,);
not I_3687 (I66897,I66888);
and I_3688 (I66915,I66861,I66429);
not I_3689 (I66933,I66717);
nand I_3690 (I66951,I66933,I66429);
not I_3691 (I66969,I66681);
nor I_3692 (I66987,I66969,I66537);
nand I_3693 (I67005,I66987,I66402);
nor I_3694 (I67023,I67005,I66951);
DFFARX1 I_3695 (I67023,I515,I66789,I67050,);
not I_3696 (I67059,I67005);
not I_3697 (I67077,I66537);
nand I_3698 (I67095,I67077,I66429);
nor I_3699 (I67113,I66537,I66717);
nand I_3700 (I67131,I66915,I67113);
nand I_3701 (I67149,I66861,I66537);
nand I_3702 (I67167,I66969,I66735);
DFFARX1 I_3703 (I67167,I515,I66789,I67194,);
DFFARX1 I_3704 (I67167,I515,I66789,I67212,);
not I_3705 (I67221,I66735);
nor I_3706 (I67239,I67221,I66771);
and I_3707 (I67257,I67239,I66402);
or I_3708 (I67275,I67257,I66276);
DFFARX1 I_3709 (I67275,I515,I66789,I67302,);
nand I_3710 (I67311,I67302,I66933);
nor I_3711 (I67329,I67311,I67095);
nor I_3712 (I67347,I67302,I66897);
DFFARX1 I_3713 (I67302,I515,I66789,I67374,);
not I_3714 (I67383,I67374);
nor I_3715 (I67401,I67383,I67059);
not I_3716 (I67419,I522);
DFFARX1 I_3717 (I67149,I515,I67419,I67446,);
not I_3718 (I67455,I67446);
nand I_3719 (I67473,I67347,I67194);
and I_3720 (I67491,I67473,I67131);
DFFARX1 I_3721 (I67491,I515,I67419,I67518,);
DFFARX1 I_3722 (I67518,I515,I67419,I67536,);
DFFARX1 I_3723 (I67401,I515,I67419,I67554,);
nand I_3724 (I67563,I67554,I67212);
not I_3725 (I67581,I67563);
DFFARX1 I_3726 (I67581,I515,I67419,I67608,);
not I_3727 (I67617,I67608);
nor I_3728 (I67635,I67455,I67617);
DFFARX1 I_3729 (I67329,I515,I67419,I67662,);
nor I_3730 (I67671,I67662,I67518);
nor I_3731 (I67689,I67662,I67581);
nand I_3732 (I67707,I67050,I66843);
and I_3733 (I67725,I67707,I67347);
DFFARX1 I_3734 (I67725,I515,I67419,I67752,);
not I_3735 (I67761,I67752);
nand I_3736 (I67779,I67761,I67662);
nand I_3737 (I67797,I67761,I67563);
nor I_3738 (I67815,I67050,I66843);
and I_3739 (I67833,I67662,I67815);
nor I_3740 (I67851,I67761,I67833);
DFFARX1 I_3741 (I67851,I515,I67419,I67878,);
nor I_3742 (I67887,I67446,I67815);
DFFARX1 I_3743 (I67887,I515,I67419,I67914,);
nor I_3744 (I67923,I67752,I67815);
not I_3745 (I67941,I67923);
nand I_3746 (I67959,I67941,I67779);
not I_3747 (I67977,I522);
DFFARX1 I_3748 (I67689,I515,I67977,I68004,);
and I_3749 (I68013,I68004,I67959);
DFFARX1 I_3750 (I68013,I515,I67977,I68040,);
DFFARX1 I_3751 (I67878,I515,I67977,I68058,);
not I_3752 (I68067,I67914);
not I_3753 (I68085,I67914);
nand I_3754 (I68103,I68085,I68067);
nor I_3755 (I68121,I68058,I68103);
DFFARX1 I_3756 (I68103,I515,I67977,I68148,);
not I_3757 (I68157,I68148);
not I_3758 (I68175,I67536);
nand I_3759 (I68193,I68085,I68175);
DFFARX1 I_3760 (I68193,I515,I67977,I68220,);
not I_3761 (I68229,I68220);
not I_3762 (I68247,I67671);
nand I_3763 (I68265,I68247,I67689);
and I_3764 (I68283,I68067,I68265);
nor I_3765 (I68301,I68193,I68283);
DFFARX1 I_3766 (I68301,I515,I67977,I68328,);
DFFARX1 I_3767 (I68283,I515,I67977,I68346,);
nor I_3768 (I68355,I67671,I67635);
nor I_3769 (I68373,I68193,I68355);
or I_3770 (I68391,I67671,I67635);
nor I_3771 (I68409,I67797,I67797);
DFFARX1 I_3772 (I68409,I515,I67977,I68436,);
not I_3773 (I68445,I68436);
nor I_3774 (I68463,I68445,I68229);
nand I_3775 (I68481,I68445,I68058);
not I_3776 (I68499,I67797);
nand I_3777 (I68517,I68499,I68175);
nand I_3778 (I68535,I68445,I68517);
nand I_3779 (I68553,I68535,I68481);
nand I_3780 (I68571,I68517,I68391);
not I_3781 (I68589,I522);
DFFARX1 I_3782 (I68121,I515,I68589,I68616,);
DFFARX1 I_3783 (I68040,I515,I68589,I68634,);
not I_3784 (I68643,I68634);
nor I_3785 (I68661,I68616,I68643);
DFFARX1 I_3786 (I68643,I515,I68589,I68688,);
nor I_3787 (I68697,I68373,I68571);
and I_3788 (I68715,I68697,I68328);
nor I_3789 (I68733,I68715,I68373);
not I_3790 (I68751,I68373);
and I_3791 (I68769,I68751,I68553);
nand I_3792 (I68787,I68769,I68328);
nor I_3793 (I68805,I68751,I68787);
DFFARX1 I_3794 (I68805,I515,I68589,I68832,);
not I_3795 (I68841,I68787);
nand I_3796 (I68859,I68643,I68841);
nand I_3797 (I68877,I68715,I68841);
DFFARX1 I_3798 (I68751,I515,I68589,I68904,);
not I_3799 (I68913,I68157);
nor I_3800 (I68931,I68913,I68553);
nor I_3801 (I68949,I68931,I68733);
DFFARX1 I_3802 (I68949,I515,I68589,I68976,);
not I_3803 (I68985,I68931);
DFFARX1 I_3804 (I68985,I515,I68589,I69012,);
not I_3805 (I69021,I69012);
nor I_3806 (I69039,I69021,I68931);
nor I_3807 (I69057,I68913,I68463);
and I_3808 (I69075,I69057,I68346);
or I_3809 (I69093,I69075,I68121);
DFFARX1 I_3810 (I69093,I515,I68589,I69120,);
not I_3811 (I69129,I69120);
nand I_3812 (I69147,I69129,I68841);
not I_3813 (I69165,I69147);
nand I_3814 (I69183,I69147,I68859);
nand I_3815 (I69201,I69129,I68715);
not I_3816 (I69219,I522);
DFFARX1 I_3817 (I68904,I515,I69219,I69246,);
and I_3818 (I69255,I69246,I69183);
DFFARX1 I_3819 (I69255,I515,I69219,I69282,);
DFFARX1 I_3820 (I68832,I515,I69219,I69300,);
not I_3821 (I69309,I69165);
not I_3822 (I69327,I68661);
nand I_3823 (I69345,I69327,I69309);
nor I_3824 (I69363,I69300,I69345);
DFFARX1 I_3825 (I69345,I515,I69219,I69390,);
not I_3826 (I69399,I69390);
not I_3827 (I69417,I68877);
nand I_3828 (I69435,I69327,I69417);
DFFARX1 I_3829 (I69435,I515,I69219,I69462,);
not I_3830 (I69471,I69462);
not I_3831 (I69489,I69039);
nand I_3832 (I69507,I69489,I68832);
and I_3833 (I69525,I69309,I69507);
nor I_3834 (I69543,I69435,I69525);
DFFARX1 I_3835 (I69543,I515,I69219,I69570,);
DFFARX1 I_3836 (I69525,I515,I69219,I69588,);
nor I_3837 (I69597,I69039,I68976);
nor I_3838 (I69615,I69435,I69597);
or I_3839 (I69633,I69039,I68976);
nor I_3840 (I69651,I68688,I69201);
DFFARX1 I_3841 (I69651,I515,I69219,I69678,);
not I_3842 (I69687,I69678);
nor I_3843 (I69705,I69687,I69471);
nand I_3844 (I69723,I69687,I69300);
not I_3845 (I69741,I68688);
nand I_3846 (I69759,I69741,I69417);
nand I_3847 (I69777,I69687,I69759);
nand I_3848 (I69795,I69777,I69723);
nand I_3849 (I69813,I69759,I69633);
not I_3850 (I69831,I522);
DFFARX1 I_3851 (I69813,I515,I69831,I69858,);
not I_3852 (I69867,I69858);
nand I_3853 (I69885,I69588,I69570);
and I_3854 (I69903,I69885,I69363);
DFFARX1 I_3855 (I69903,I515,I69831,I69930,);
DFFARX1 I_3856 (I69399,I515,I69831,I69948,);
and I_3857 (I69957,I69948,I69363);
nor I_3858 (I69975,I69930,I69957);
DFFARX1 I_3859 (I69975,I515,I69831,I70002,);
nand I_3860 (I70011,I69948,I69363);
nand I_3861 (I70029,I69867,I70011);
not I_3862 (I70047,I70029);
DFFARX1 I_3863 (I69570,I515,I69831,I70074,);
DFFARX1 I_3864 (I70074,I515,I69831,I70092,);
nand I_3865 (I70101,I69615,I69795);
and I_3866 (I70119,I70101,I69282);
DFFARX1 I_3867 (I70119,I515,I69831,I70146,);
DFFARX1 I_3868 (I70146,I515,I69831,I70164,);
not I_3869 (I70173,I70164);
not I_3870 (I70191,I70146);
nand I_3871 (I70209,I70191,I70011);
nor I_3872 (I70227,I69705,I69795);
not I_3873 (I70245,I70227);
nor I_3874 (I70263,I70191,I70245);
nor I_3875 (I70281,I69867,I70263);
DFFARX1 I_3876 (I70281,I515,I69831,I70308,);
nor I_3877 (I70317,I69930,I70245);
nor I_3878 (I70335,I70146,I70317);
nor I_3879 (I70353,I70074,I70227);
nor I_3880 (I70371,I69930,I70227);
not I_3881 (I70389,I522);
DFFARX1 I_3882 (I116,I515,I70389,I70416,);
and I_3883 (I70425,I70416,I260);
DFFARX1 I_3884 (I70425,I515,I70389,I70452,);
DFFARX1 I_3885 (I372,I515,I70389,I70470,);
not I_3886 (I70479,I436);
not I_3887 (I70497,I228);
nand I_3888 (I70515,I70497,I70479);
nor I_3889 (I70533,I70470,I70515);
DFFARX1 I_3890 (I70515,I515,I70389,I70560,);
not I_3891 (I70569,I70560);
not I_3892 (I70587,I220);
nand I_3893 (I70605,I70497,I70587);
DFFARX1 I_3894 (I70605,I515,I70389,I70632,);
not I_3895 (I70641,I70632);
not I_3896 (I70659,I388);
nand I_3897 (I70677,I70659,I180);
and I_3898 (I70695,I70479,I70677);
nor I_3899 (I70713,I70605,I70695);
DFFARX1 I_3900 (I70713,I515,I70389,I70740,);
DFFARX1 I_3901 (I70695,I515,I70389,I70758,);
nor I_3902 (I70767,I388,I444);
nor I_3903 (I70785,I70605,I70767);
or I_3904 (I70803,I388,I444);
nor I_3905 (I70821,I404,I476);
DFFARX1 I_3906 (I70821,I515,I70389,I70848,);
not I_3907 (I70857,I70848);
nor I_3908 (I70875,I70857,I70641);
nand I_3909 (I70893,I70857,I70470);
not I_3910 (I70911,I404);
nand I_3911 (I70929,I70911,I70587);
nand I_3912 (I70947,I70857,I70929);
nand I_3913 (I70965,I70947,I70893);
nand I_3914 (I70983,I70929,I70803);
not I_3915 (I71001,I522);
DFFARX1 I_3916 (I70533,I515,I71001,I71028,);
DFFARX1 I_3917 (I70452,I515,I71001,I71046,);
not I_3918 (I71055,I71046);
nor I_3919 (I71073,I71028,I71055);
DFFARX1 I_3920 (I71055,I515,I71001,I71100,);
nor I_3921 (I71109,I70785,I70983);
and I_3922 (I71127,I71109,I70740);
nor I_3923 (I71145,I71127,I70785);
not I_3924 (I71163,I70785);
and I_3925 (I71181,I71163,I70965);
nand I_3926 (I71199,I71181,I70740);
nor I_3927 (I71217,I71163,I71199);
DFFARX1 I_3928 (I71217,I515,I71001,I71244,);
not I_3929 (I71253,I71199);
nand I_3930 (I71271,I71055,I71253);
nand I_3931 (I71289,I71127,I71253);
DFFARX1 I_3932 (I71163,I515,I71001,I71316,);
not I_3933 (I71325,I70569);
nor I_3934 (I71343,I71325,I70965);
nor I_3935 (I71361,I71343,I71145);
DFFARX1 I_3936 (I71361,I515,I71001,I71388,);
not I_3937 (I71397,I71343);
DFFARX1 I_3938 (I71397,I515,I71001,I71424,);
not I_3939 (I71433,I71424);
nor I_3940 (I71451,I71433,I71343);
nor I_3941 (I71469,I71325,I70875);
and I_3942 (I71487,I71469,I70758);
or I_3943 (I71505,I71487,I70533);
DFFARX1 I_3944 (I71505,I515,I71001,I71532,);
not I_3945 (I71541,I71532);
nand I_3946 (I71559,I71541,I71253);
not I_3947 (I71577,I71559);
nand I_3948 (I71595,I71559,I71271);
nand I_3949 (I71613,I71541,I71127);
not I_3950 (I71631,I522);
DFFARX1 I_3951 (I71289,I515,I71631,I71658,);
not I_3952 (I71667,I71658);
nand I_3953 (I71685,I71613,I71316);
and I_3954 (I71703,I71685,I71073);
DFFARX1 I_3955 (I71703,I515,I71631,I71730,);
DFFARX1 I_3956 (I71388,I515,I71631,I71748,);
and I_3957 (I71757,I71748,I71451);
nor I_3958 (I71775,I71730,I71757);
DFFARX1 I_3959 (I71775,I515,I71631,I71802,);
nand I_3960 (I71811,I71748,I71451);
nand I_3961 (I71829,I71667,I71811);
not I_3962 (I71847,I71829);
DFFARX1 I_3963 (I71595,I515,I71631,I71874,);
DFFARX1 I_3964 (I71874,I515,I71631,I71892,);
nand I_3965 (I71901,I71100,I71577);
and I_3966 (I71919,I71901,I71244);
DFFARX1 I_3967 (I71919,I515,I71631,I71946,);
DFFARX1 I_3968 (I71946,I515,I71631,I71964,);
not I_3969 (I71973,I71964);
not I_3970 (I71991,I71946);
nand I_3971 (I72009,I71991,I71811);
nor I_3972 (I72027,I71244,I71577);
not I_3973 (I72045,I72027);
nor I_3974 (I72063,I71991,I72045);
nor I_3975 (I72081,I71667,I72063);
DFFARX1 I_3976 (I72081,I515,I71631,I72108,);
nor I_3977 (I72117,I71730,I72045);
nor I_3978 (I72135,I71946,I72117);
nor I_3979 (I72153,I71874,I72027);
nor I_3980 (I72171,I71730,I72027);
not I_3981 (I72189,I522);
DFFARX1 I_3982 (I72009,I515,I72189,I72216,);
DFFARX1 I_3983 (I72216,I515,I72189,I72234,);
not I_3984 (I72243,I72234);
not I_3985 (I72261,I72216);
DFFARX1 I_3986 (I72171,I515,I72189,I72288,);
not I_3987 (I72297,I72288);
and I_3988 (I72315,I72261,I71802);
not I_3989 (I72333,I71892);
nand I_3990 (I72351,I72333,I71802);
not I_3991 (I72369,I72153);
nor I_3992 (I72387,I72369,I72135);
nand I_3993 (I72405,I72387,I71847);
nor I_3994 (I72423,I72405,I72351);
DFFARX1 I_3995 (I72423,I515,I72189,I72450,);
not I_3996 (I72459,I72405);
not I_3997 (I72477,I72135);
nand I_3998 (I72495,I72477,I71802);
nor I_3999 (I72513,I72135,I71892);
nand I_4000 (I72531,I72315,I72513);
nand I_4001 (I72549,I72261,I72135);
nand I_4002 (I72567,I72369,I71802);
DFFARX1 I_4003 (I72567,I515,I72189,I72594,);
DFFARX1 I_4004 (I72567,I515,I72189,I72612,);
not I_4005 (I72621,I71802);
nor I_4006 (I72639,I72621,I72108);
and I_4007 (I72657,I72639,I71973);
or I_4008 (I72675,I72657,I72171);
DFFARX1 I_4009 (I72675,I515,I72189,I72702,);
nand I_4010 (I72711,I72702,I72333);
nor I_4011 (I72729,I72711,I72495);
nor I_4012 (I72747,I72702,I72297);
DFFARX1 I_4013 (I72702,I515,I72189,I72774,);
not I_4014 (I72783,I72774);
nor I_4015 (I72801,I72783,I72459);
not I_4016 (I72819,I522);
DFFARX1 I_4017 (I72729,I515,I72819,I72846,);
nand I_4018 (I72855,I72846,I72243);
DFFARX1 I_4019 (I72612,I515,I72819,I72882,);
DFFARX1 I_4020 (I72882,I515,I72819,I72900,);
not I_4021 (I72909,I72900);
not I_4022 (I72927,I72450);
nor I_4023 (I72945,I72450,I72549);
not I_4024 (I72963,I72531);
nand I_4025 (I72981,I72927,I72963);
nor I_4026 (I72999,I72531,I72450);
and I_4027 (I73017,I72999,I72855);
not I_4028 (I73035,I72801);
nand I_4029 (I73053,I73035,I72450);
nor I_4030 (I73071,I72801,I72747);
not I_4031 (I73089,I73071);
nand I_4032 (I73107,I72945,I73089);
DFFARX1 I_4033 (I73071,I515,I72819,I73134,);
nor I_4034 (I73143,I72747,I72531);
nor I_4035 (I73161,I73143,I72549);
and I_4036 (I73179,I73161,I73053);
DFFARX1 I_4037 (I73179,I515,I72819,I73206,);
nor I_4038 (I73215,I73143,I72981);
or I_4039 (I73233,I73071,I73143);
nor I_4040 (I73251,I72747,I72594);
DFFARX1 I_4041 (I73251,I515,I72819,I73278,);
not I_4042 (I73287,I73278);
nand I_4043 (I73305,I73287,I72927);
nor I_4044 (I73323,I73305,I72549);
DFFARX1 I_4045 (I73323,I515,I72819,I73350,);
nor I_4046 (I73359,I73287,I72981);
nor I_4047 (I73377,I73143,I73359);
not I_4048 (I73395,I522);
DFFARX1 I_4049 (I73107,I515,I73395,I73422,);
not I_4050 (I73431,I73422);
nand I_4051 (I73449,I73350,I73134);
and I_4052 (I73467,I73449,I73233);
DFFARX1 I_4053 (I73467,I515,I73395,I73494,);
DFFARX1 I_4054 (I73017,I515,I73395,I73512,);
and I_4055 (I73521,I73512,I73215);
nor I_4056 (I73539,I73494,I73521);
DFFARX1 I_4057 (I73539,I515,I73395,I73566,);
nand I_4058 (I73575,I73512,I73215);
nand I_4059 (I73593,I73431,I73575);
not I_4060 (I73611,I73593);
DFFARX1 I_4061 (I73017,I515,I73395,I73638,);
DFFARX1 I_4062 (I73638,I515,I73395,I73656,);
nand I_4063 (I73665,I72909,I73377);
and I_4064 (I73683,I73665,I73350);
DFFARX1 I_4065 (I73683,I515,I73395,I73710,);
DFFARX1 I_4066 (I73710,I515,I73395,I73728,);
not I_4067 (I73737,I73728);
not I_4068 (I73755,I73710);
nand I_4069 (I73773,I73755,I73575);
nor I_4070 (I73791,I73206,I73377);
not I_4071 (I73809,I73791);
nor I_4072 (I73827,I73755,I73809);
nor I_4073 (I73845,I73431,I73827);
DFFARX1 I_4074 (I73845,I515,I73395,I73872,);
nor I_4075 (I73881,I73494,I73809);
nor I_4076 (I73899,I73710,I73881);
nor I_4077 (I73917,I73638,I73791);
nor I_4078 (I73935,I73494,I73791);
not I_4079 (I73953,I522);
DFFARX1 I_4080 (I73737,I515,I73953,I73980,);
not I_4081 (I73989,I73980);
nand I_4082 (I74007,I73566,I73773);
and I_4083 (I74025,I74007,I73935);
DFFARX1 I_4084 (I74025,I515,I73953,I74052,);
DFFARX1 I_4085 (I74052,I515,I73953,I74070,);
DFFARX1 I_4086 (I73656,I515,I73953,I74088,);
nand I_4087 (I74097,I74088,I73611);
not I_4088 (I74115,I74097);
DFFARX1 I_4089 (I74115,I515,I73953,I74142,);
not I_4090 (I74151,I74142);
nor I_4091 (I74169,I73989,I74151);
DFFARX1 I_4092 (I73899,I515,I73953,I74196,);
nor I_4093 (I74205,I74196,I74052);
nor I_4094 (I74223,I74196,I74115);
nand I_4095 (I74241,I73872,I73917);
and I_4096 (I74259,I74241,I73935);
DFFARX1 I_4097 (I74259,I515,I73953,I74286,);
not I_4098 (I74295,I74286);
nand I_4099 (I74313,I74295,I74196);
nand I_4100 (I74331,I74295,I74097);
nor I_4101 (I74349,I73566,I73917);
and I_4102 (I74367,I74196,I74349);
nor I_4103 (I74385,I74295,I74367);
DFFARX1 I_4104 (I74385,I515,I73953,I74412,);
nor I_4105 (I74421,I73980,I74349);
DFFARX1 I_4106 (I74421,I515,I73953,I74448,);
nor I_4107 (I74457,I74286,I74349);
not I_4108 (I74475,I74457);
nand I_4109 (I74493,I74475,I74313);
not I_4110 (I74511,I522);
DFFARX1 I_4111 (I74412,I515,I74511,I74538,);
not I_4112 (I74547,I74538);
nand I_4113 (I74565,I74223,I74169);
and I_4114 (I74583,I74565,I74070);
DFFARX1 I_4115 (I74583,I515,I74511,I74610,);
not I_4116 (I74619,I74493);
DFFARX1 I_4117 (I74331,I515,I74511,I74646,);
not I_4118 (I74655,I74646);
nor I_4119 (I74673,I74655,I74547);
and I_4120 (I74691,I74673,I74493);
nor I_4121 (I74709,I74655,I74619);
nor I_4122 (I74727,I74610,I74709);
DFFARX1 I_4123 (I74448,I515,I74511,I74754,);
nor I_4124 (I74763,I74754,I74610);
not I_4125 (I74781,I74763);
not I_4126 (I74799,I74754);
nor I_4127 (I74817,I74799,I74691);
DFFARX1 I_4128 (I74817,I515,I74511,I74844,);
nand I_4129 (I74853,I74448,I74223);
and I_4130 (I74871,I74853,I74331);
DFFARX1 I_4131 (I74871,I515,I74511,I74898,);
nor I_4132 (I74907,I74898,I74754);
DFFARX1 I_4133 (I74907,I515,I74511,I74934,);
nand I_4134 (I74943,I74898,I74799);
nand I_4135 (I74961,I74781,I74943);
not I_4136 (I74979,I74898);
nor I_4137 (I74997,I74979,I74691);
DFFARX1 I_4138 (I74997,I515,I74511,I75024,);
nor I_4139 (I75033,I74205,I74223);
or I_4140 (I75051,I74754,I75033);
nor I_4141 (I75069,I74898,I75033);
or I_4142 (I75087,I74610,I75033);
DFFARX1 I_4143 (I75033,I515,I74511,I75114,);
not I_4144 (I75123,I522);
DFFARX1 I_4145 (I75069,I515,I75123,I75150,);
DFFARX1 I_4146 (I75150,I515,I75123,I75168,);
not I_4147 (I75177,I75168);
not I_4148 (I75195,I75150);
DFFARX1 I_4149 (I74727,I515,I75123,I75222,);
nand I_4150 (I75231,I75222,I75114);
not I_4151 (I75249,I75114);
not I_4152 (I75267,I75087);
nand I_4153 (I75285,I74961,I74934);
and I_4154 (I75303,I74961,I74934);
not I_4155 (I75321,I74844);
nand I_4156 (I75339,I75321,I75267);
nor I_4157 (I75357,I75339,I75231);
nor I_4158 (I75375,I75249,I75339);
nand I_4159 (I75393,I75303,I75375);
not I_4160 (I75411,I75024);
nor I_4161 (I75429,I75411,I74961);
nor I_4162 (I75447,I75429,I74844);
nor I_4163 (I75465,I75195,I75447);
DFFARX1 I_4164 (I75465,I515,I75123,I75492,);
not I_4165 (I75501,I75429);
DFFARX1 I_4166 (I75501,I515,I75123,I75528,);
and I_4167 (I75537,I75222,I75429);
nor I_4168 (I75555,I75411,I74934);
and I_4169 (I75573,I75555,I75051);
or I_4170 (I75591,I75573,I75069);
DFFARX1 I_4171 (I75591,I515,I75123,I75618,);
nor I_4172 (I75627,I75618,I75321);
DFFARX1 I_4173 (I75627,I515,I75123,I75654,);
nand I_4174 (I75663,I75618,I75222);
nand I_4175 (I75681,I75321,I75663);
nor I_4176 (I75699,I75681,I75285);
not I_4177 (I75717,I522);
DFFARX1 I_4178 (I75357,I515,I75717,I75744,);
and I_4179 (I75753,I75744,I75654);
DFFARX1 I_4180 (I75753,I515,I75717,I75780,);
DFFARX1 I_4181 (I75393,I515,I75717,I75798,);
not I_4182 (I75807,I75699);
not I_4183 (I75825,I75357);
nand I_4184 (I75843,I75825,I75807);
nor I_4185 (I75861,I75798,I75843);
DFFARX1 I_4186 (I75843,I515,I75717,I75888,);
not I_4187 (I75897,I75888);
not I_4188 (I75915,I75528);
nand I_4189 (I75933,I75825,I75915);
DFFARX1 I_4190 (I75933,I515,I75717,I75960,);
not I_4191 (I75969,I75960);
not I_4192 (I75987,I75492);
nand I_4193 (I76005,I75987,I75177);
and I_4194 (I76023,I75807,I76005);
nor I_4195 (I76041,I75933,I76023);
DFFARX1 I_4196 (I76041,I515,I75717,I76068,);
DFFARX1 I_4197 (I76023,I515,I75717,I76086,);
nor I_4198 (I76095,I75492,I75654);
nor I_4199 (I76113,I75933,I76095);
or I_4200 (I76131,I75492,I75654);
nor I_4201 (I76149,I75537,I75393);
DFFARX1 I_4202 (I76149,I515,I75717,I76176,);
not I_4203 (I76185,I76176);
nor I_4204 (I76203,I76185,I75969);
nand I_4205 (I76221,I76185,I75798);
not I_4206 (I76239,I75537);
nand I_4207 (I76257,I76239,I75915);
nand I_4208 (I76275,I76185,I76257);
nand I_4209 (I76293,I76275,I76221);
nand I_4210 (I76311,I76257,I76131);
not I_4211 (I76329,I522);
DFFARX1 I_4212 (I76068,I515,I76329,I76356,);
not I_4213 (I76365,I76356);
DFFARX1 I_4214 (I76311,I515,I76329,I76392,);
not I_4215 (I76401,I76068);
nand I_4216 (I76419,I76401,I75861);
not I_4217 (I76437,I76419);
nor I_4218 (I76455,I76437,I76086);
nor I_4219 (I76473,I76365,I76455);
DFFARX1 I_4220 (I76473,I515,I76329,I76500,);
not I_4221 (I76509,I76086);
nand I_4222 (I76527,I76509,I76437);
and I_4223 (I76545,I76509,I75897);
nand I_4224 (I76563,I76545,I75861);
nor I_4225 (I76581,I76563,I76509);
and I_4226 (I76599,I76392,I76563);
not I_4227 (I76617,I76563);
nand I_4228 (I76635,I76392,I76617);
nor I_4229 (I76653,I76356,I76563);
not I_4230 (I76671,I76293);
nor I_4231 (I76689,I76671,I75897);
nand I_4232 (I76707,I76689,I76509);
nor I_4233 (I76725,I76419,I76707);
nor I_4234 (I76743,I76671,I75780);
and I_4235 (I76761,I76743,I76113);
or I_4236 (I76779,I76761,I76203);
DFFARX1 I_4237 (I76779,I515,I76329,I76806,);
nor I_4238 (I76815,I76806,I76527);
DFFARX1 I_4239 (I76815,I515,I76329,I76842,);
DFFARX1 I_4240 (I76806,I515,I76329,I76860,);
not I_4241 (I76869,I76806);
nor I_4242 (I76887,I76869,I76392);
nor I_4243 (I76905,I76689,I76887);
DFFARX1 I_4244 (I76905,I515,I76329,I76932,);
not I_4245 (I76941,I522);
DFFARX1 I_4246 (I76635,I515,I76941,I76968,);
not I_4247 (I76977,I76968);
nand I_4248 (I76995,I76932,I76599);
and I_4249 (I77013,I76995,I76842);
DFFARX1 I_4250 (I77013,I515,I76941,I77040,);
DFFARX1 I_4251 (I76581,I515,I76941,I77058,);
and I_4252 (I77067,I77058,I76653);
nor I_4253 (I77085,I77040,I77067);
DFFARX1 I_4254 (I77085,I515,I76941,I77112,);
nand I_4255 (I77121,I77058,I76653);
nand I_4256 (I77139,I76977,I77121);
not I_4257 (I77157,I77139);
DFFARX1 I_4258 (I76725,I515,I76941,I77184,);
DFFARX1 I_4259 (I77184,I515,I76941,I77202,);
nand I_4260 (I77211,I76500,I76860);
and I_4261 (I77229,I77211,I76842);
DFFARX1 I_4262 (I77229,I515,I76941,I77256,);
DFFARX1 I_4263 (I77256,I515,I76941,I77274,);
not I_4264 (I77283,I77274);
not I_4265 (I77301,I77256);
nand I_4266 (I77319,I77301,I77121);
nor I_4267 (I77337,I76653,I76860);
not I_4268 (I77355,I77337);
nor I_4269 (I77373,I77301,I77355);
nor I_4270 (I77391,I76977,I77373);
DFFARX1 I_4271 (I77391,I515,I76941,I77418,);
nor I_4272 (I77427,I77040,I77355);
nor I_4273 (I77445,I77256,I77427);
nor I_4274 (I77463,I77184,I77337);
nor I_4275 (I77481,I77040,I77337);
not I_4276 (I77499,I522);
DFFARX1 I_4277 (I77283,I515,I77499,I77526,);
and I_4278 (I77535,I77526,I77112);
DFFARX1 I_4279 (I77535,I515,I77499,I77562,);
DFFARX1 I_4280 (I77418,I515,I77499,I77580,);
not I_4281 (I77589,I77445);
not I_4282 (I77607,I77481);
nand I_4283 (I77625,I77607,I77589);
nor I_4284 (I77643,I77580,I77625);
DFFARX1 I_4285 (I77625,I515,I77499,I77670,);
not I_4286 (I77679,I77670);
not I_4287 (I77697,I77157);
nand I_4288 (I77715,I77607,I77697);
DFFARX1 I_4289 (I77715,I515,I77499,I77742,);
not I_4290 (I77751,I77742);
not I_4291 (I77769,I77481);
nand I_4292 (I77787,I77769,I77202);
and I_4293 (I77805,I77589,I77787);
nor I_4294 (I77823,I77715,I77805);
DFFARX1 I_4295 (I77823,I515,I77499,I77850,);
DFFARX1 I_4296 (I77805,I515,I77499,I77868,);
nor I_4297 (I77877,I77481,I77463);
nor I_4298 (I77895,I77715,I77877);
or I_4299 (I77913,I77481,I77463);
nor I_4300 (I77931,I77319,I77112);
DFFARX1 I_4301 (I77931,I515,I77499,I77958,);
not I_4302 (I77967,I77958);
nor I_4303 (I77985,I77967,I77751);
nand I_4304 (I78003,I77967,I77580);
not I_4305 (I78021,I77319);
nand I_4306 (I78039,I78021,I77697);
nand I_4307 (I78057,I77967,I78039);
nand I_4308 (I78075,I78057,I78003);
nand I_4309 (I78093,I78039,I77913);
not I_4310 (I78111,I522);
DFFARX1 I_4311 (I77850,I515,I78111,I78138,);
DFFARX1 I_4312 (I78138,I515,I78111,I78156,);
not I_4313 (I78165,I78156);
not I_4314 (I78183,I78138);
DFFARX1 I_4315 (I77850,I515,I78111,I78210,);
not I_4316 (I78219,I78210);
and I_4317 (I78237,I78183,I77643);
not I_4318 (I78255,I77562);
nand I_4319 (I78273,I78255,I77643);
not I_4320 (I78291,I77868);
nor I_4321 (I78309,I78291,I77895);
nand I_4322 (I78327,I78309,I77985);
nor I_4323 (I78345,I78327,I78273);
DFFARX1 I_4324 (I78345,I515,I78111,I78372,);
not I_4325 (I78381,I78327);
not I_4326 (I78399,I77895);
nand I_4327 (I78417,I78399,I77643);
nor I_4328 (I78435,I77895,I77562);
nand I_4329 (I78453,I78237,I78435);
nand I_4330 (I78471,I78183,I77895);
nand I_4331 (I78489,I78291,I78075);
DFFARX1 I_4332 (I78489,I515,I78111,I78516,);
DFFARX1 I_4333 (I78489,I515,I78111,I78534,);
not I_4334 (I78543,I78075);
nor I_4335 (I78561,I78543,I78093);
and I_4336 (I78579,I78561,I77679);
or I_4337 (I78597,I78579,I77643);
DFFARX1 I_4338 (I78597,I515,I78111,I78624,);
nand I_4339 (I78633,I78624,I78255);
nor I_4340 (I78651,I78633,I78417);
nor I_4341 (I78669,I78624,I78219);
DFFARX1 I_4342 (I78624,I515,I78111,I78696,);
not I_4343 (I78705,I78696);
nor I_4344 (I78723,I78705,I78381);
not I_4345 (I78741,I522);
DFFARX1 I_4346 (I78372,I515,I78741,I78768,);
nand I_4347 (I78777,I78372,I78471);
and I_4348 (I78795,I78777,I78165);
DFFARX1 I_4349 (I78795,I515,I78741,I78822,);
nor I_4350 (I78831,I78822,I78768);
not I_4351 (I78849,I78822);
DFFARX1 I_4352 (I78453,I515,I78741,I78876,);
nand I_4353 (I78885,I78876,I78651);
not I_4354 (I78903,I78885);
DFFARX1 I_4355 (I78903,I515,I78741,I78930,);
not I_4356 (I78939,I78930);
nor I_4357 (I78957,I78768,I78885);
nor I_4358 (I78975,I78822,I78957);
DFFARX1 I_4359 (I78723,I515,I78741,I79002,);
DFFARX1 I_4360 (I79002,I515,I78741,I79020,);
not I_4361 (I79029,I79020);
not I_4362 (I79047,I79002);
nand I_4363 (I79065,I79047,I78849);
nand I_4364 (I79083,I78669,I78669);
and I_4365 (I79101,I79083,I78516);
DFFARX1 I_4366 (I79101,I515,I78741,I79128,);
nor I_4367 (I79137,I79128,I78768);
DFFARX1 I_4368 (I79137,I515,I78741,I79164,);
DFFARX1 I_4369 (I79128,I515,I78741,I79182,);
nor I_4370 (I79191,I78534,I78669);
not I_4371 (I79209,I79191);
nor I_4372 (I79227,I79029,I79209);
nand I_4373 (I79245,I79047,I79209);
nor I_4374 (I79263,I78768,I79191);
DFFARX1 I_4375 (I79191,I515,I78741,I79290,);
not I_4376 (I79299,I522);
DFFARX1 I_4377 (I79164,I515,I79299,I79326,);
DFFARX1 I_4378 (I79326,I515,I79299,I79344,);
not I_4379 (I79353,I79344);
not I_4380 (I79371,I79326);
DFFARX1 I_4381 (I79263,I515,I79299,I79398,);
not I_4382 (I79407,I79398);
and I_4383 (I79425,I79371,I79065);
not I_4384 (I79443,I79164);
nand I_4385 (I79461,I79443,I79065);
not I_4386 (I79479,I78975);
nor I_4387 (I79497,I79479,I79290);
nand I_4388 (I79515,I79497,I79227);
nor I_4389 (I79533,I79515,I79461);
DFFARX1 I_4390 (I79533,I515,I79299,I79560,);
not I_4391 (I79569,I79515);
not I_4392 (I79587,I79290);
nand I_4393 (I79605,I79587,I79065);
nor I_4394 (I79623,I79290,I79164);
nand I_4395 (I79641,I79425,I79623);
nand I_4396 (I79659,I79371,I79290);
nand I_4397 (I79677,I79479,I79182);
DFFARX1 I_4398 (I79677,I515,I79299,I79704,);
DFFARX1 I_4399 (I79677,I515,I79299,I79722,);
not I_4400 (I79731,I79182);
nor I_4401 (I79749,I79731,I79245);
and I_4402 (I79767,I79749,I78939);
or I_4403 (I79785,I79767,I78831);
DFFARX1 I_4404 (I79785,I515,I79299,I79812,);
nand I_4405 (I79821,I79812,I79443);
nor I_4406 (I79839,I79821,I79605);
nor I_4407 (I79857,I79812,I79407);
DFFARX1 I_4408 (I79812,I515,I79299,I79884,);
not I_4409 (I79893,I79884);
nor I_4410 (I79911,I79893,I79569);
not I_4411 (I79929,I522);
DFFARX1 I_4412 (I79560,I515,I79929,I79956,);
not I_4413 (I79965,I79956);
nand I_4414 (I79983,I79857,I79353);
and I_4415 (I80001,I79983,I79641);
DFFARX1 I_4416 (I80001,I515,I79929,I80028,);
not I_4417 (I80037,I79839);
DFFARX1 I_4418 (I79560,I515,I79929,I80064,);
not I_4419 (I80073,I80064);
nor I_4420 (I80091,I80073,I79965);
and I_4421 (I80109,I80091,I79839);
nor I_4422 (I80127,I80073,I80037);
nor I_4423 (I80145,I80028,I80127);
DFFARX1 I_4424 (I79911,I515,I79929,I80172,);
nor I_4425 (I80181,I80172,I80028);
not I_4426 (I80199,I80181);
not I_4427 (I80217,I80172);
nor I_4428 (I80235,I80217,I80109);
DFFARX1 I_4429 (I80235,I515,I79929,I80262,);
nand I_4430 (I80271,I79857,I79659);
and I_4431 (I80289,I80271,I79722);
DFFARX1 I_4432 (I80289,I515,I79929,I80316,);
nor I_4433 (I80325,I80316,I80172);
DFFARX1 I_4434 (I80325,I515,I79929,I80352,);
nand I_4435 (I80361,I80316,I80217);
nand I_4436 (I80379,I80199,I80361);
not I_4437 (I80397,I80316);
nor I_4438 (I80415,I80397,I80109);
DFFARX1 I_4439 (I80415,I515,I79929,I80442,);
nor I_4440 (I80451,I79704,I79659);
or I_4441 (I80469,I80172,I80451);
nor I_4442 (I80487,I80316,I80451);
or I_4443 (I80505,I80028,I80451);
DFFARX1 I_4444 (I80451,I515,I79929,I80532,);
not I_4445 (I80541,I522);
DFFARX1 I_4446 (I80487,I515,I80541,I80568,);
nand I_4447 (I80577,I80568,I80262);
DFFARX1 I_4448 (I80469,I515,I80541,I80604,);
DFFARX1 I_4449 (I80604,I515,I80541,I80622,);
not I_4450 (I80631,I80622);
not I_4451 (I80649,I80145);
nor I_4452 (I80667,I80145,I80442);
not I_4453 (I80685,I80487);
nand I_4454 (I80703,I80649,I80685);
nor I_4455 (I80721,I80487,I80145);
and I_4456 (I80739,I80721,I80577);
not I_4457 (I80757,I80352);
nand I_4458 (I80775,I80757,I80505);
nor I_4459 (I80793,I80352,I80352);
not I_4460 (I80811,I80793);
nand I_4461 (I80829,I80667,I80811);
DFFARX1 I_4462 (I80793,I515,I80541,I80856,);
nor I_4463 (I80865,I80379,I80487);
nor I_4464 (I80883,I80865,I80442);
and I_4465 (I80901,I80883,I80775);
DFFARX1 I_4466 (I80901,I515,I80541,I80928,);
nor I_4467 (I80937,I80865,I80703);
or I_4468 (I80955,I80793,I80865);
nor I_4469 (I80973,I80379,I80532);
DFFARX1 I_4470 (I80973,I515,I80541,I81000,);
not I_4471 (I81009,I81000);
nand I_4472 (I81027,I81009,I80649);
nor I_4473 (I81045,I81027,I80442);
DFFARX1 I_4474 (I81045,I515,I80541,I81072,);
nor I_4475 (I81081,I81009,I80703);
nor I_4476 (I81099,I80865,I81081);
not I_4477 (I81117,I522);
DFFARX1 I_4478 (I80955,I515,I81117,I81144,);
not I_4479 (I81153,I81144);
nand I_4480 (I81171,I80928,I81072);
and I_4481 (I81189,I81171,I81099);
DFFARX1 I_4482 (I81189,I515,I81117,I81216,);
DFFARX1 I_4483 (I81216,I515,I81117,I81234,);
DFFARX1 I_4484 (I80937,I515,I81117,I81252,);
nand I_4485 (I81261,I81252,I80739);
not I_4486 (I81279,I81261);
DFFARX1 I_4487 (I81279,I515,I81117,I81306,);
not I_4488 (I81315,I81306);
nor I_4489 (I81333,I81153,I81315);
DFFARX1 I_4490 (I80856,I515,I81117,I81360,);
nor I_4491 (I81369,I81360,I81216);
nor I_4492 (I81387,I81360,I81279);
nand I_4493 (I81405,I81072,I80829);
and I_4494 (I81423,I81405,I80631);
DFFARX1 I_4495 (I81423,I515,I81117,I81450,);
not I_4496 (I81459,I81450);
nand I_4497 (I81477,I81459,I81360);
nand I_4498 (I81495,I81459,I81261);
nor I_4499 (I81513,I80739,I80829);
and I_4500 (I81531,I81360,I81513);
nor I_4501 (I81549,I81459,I81531);
DFFARX1 I_4502 (I81549,I515,I81117,I81576,);
nor I_4503 (I81585,I81144,I81513);
DFFARX1 I_4504 (I81585,I515,I81117,I81612,);
nor I_4505 (I81621,I81450,I81513);
not I_4506 (I81639,I81621);
nand I_4507 (I81657,I81639,I81477);
not I_4508 (I81675,I522);
DFFARX1 I_4509 (I81495,I515,I81675,I81702,);
not I_4510 (I81711,I81702);
DFFARX1 I_4511 (I81495,I515,I81675,I81738,);
not I_4512 (I81747,I81387);
nand I_4513 (I81765,I81747,I81234);
not I_4514 (I81783,I81765);
nor I_4515 (I81801,I81783,I81369);
nor I_4516 (I81819,I81711,I81801);
DFFARX1 I_4517 (I81819,I515,I81675,I81846,);
not I_4518 (I81855,I81369);
nand I_4519 (I81873,I81855,I81783);
and I_4520 (I81891,I81855,I81657);
nand I_4521 (I81909,I81891,I81612);
nor I_4522 (I81927,I81909,I81855);
and I_4523 (I81945,I81738,I81909);
not I_4524 (I81963,I81909);
nand I_4525 (I81981,I81738,I81963);
nor I_4526 (I81999,I81702,I81909);
not I_4527 (I82017,I81333);
nor I_4528 (I82035,I82017,I81657);
nand I_4529 (I82053,I82035,I81855);
nor I_4530 (I82071,I81765,I82053);
nor I_4531 (I82089,I82017,I81612);
and I_4532 (I82107,I82089,I81387);
or I_4533 (I82125,I82107,I81576);
DFFARX1 I_4534 (I82125,I515,I81675,I82152,);
nor I_4535 (I82161,I82152,I81873);
DFFARX1 I_4536 (I82161,I515,I81675,I82188,);
DFFARX1 I_4537 (I82152,I515,I81675,I82206,);
not I_4538 (I82215,I82152);
nor I_4539 (I82233,I82215,I81738);
nor I_4540 (I82251,I82035,I82233);
DFFARX1 I_4541 (I82251,I515,I81675,I82278,);
not I_4542 (I82287,I522);
DFFARX1 I_4543 (I82278,I515,I82287,I82314,);
DFFARX1 I_4544 (I81927,I515,I82287,I82332,);
not I_4545 (I82341,I82332);
nor I_4546 (I82359,I82314,I82341);
DFFARX1 I_4547 (I82341,I515,I82287,I82386,);
nor I_4548 (I82395,I82071,I81999);
and I_4549 (I82413,I82395,I82188);
nor I_4550 (I82431,I82413,I82071);
not I_4551 (I82449,I82071);
and I_4552 (I82467,I82449,I81945);
nand I_4553 (I82485,I82467,I81846);
nor I_4554 (I82503,I82449,I82485);
DFFARX1 I_4555 (I82503,I515,I82287,I82530,);
not I_4556 (I82539,I82485);
nand I_4557 (I82557,I82341,I82539);
nand I_4558 (I82575,I82413,I82539);
DFFARX1 I_4559 (I82449,I515,I82287,I82602,);
not I_4560 (I82611,I82206);
nor I_4561 (I82629,I82611,I81945);
nor I_4562 (I82647,I82629,I82431);
DFFARX1 I_4563 (I82647,I515,I82287,I82674,);
not I_4564 (I82683,I82629);
DFFARX1 I_4565 (I82683,I515,I82287,I82710,);
not I_4566 (I82719,I82710);
nor I_4567 (I82737,I82719,I82629);
nor I_4568 (I82755,I82611,I81999);
and I_4569 (I82773,I82755,I81981);
or I_4570 (I82791,I82773,I82188);
DFFARX1 I_4571 (I82791,I515,I82287,I82818,);
not I_4572 (I82827,I82818);
nand I_4573 (I82845,I82827,I82539);
not I_4574 (I82863,I82845);
nand I_4575 (I82881,I82845,I82557);
nand I_4576 (I82899,I82827,I82413);
not I_4577 (I82917,I522);
DFFARX1 I_4578 (I82575,I515,I82917,I82944,);
not I_4579 (I82953,I82944);
nand I_4580 (I82971,I82899,I82602);
and I_4581 (I82989,I82971,I82359);
DFFARX1 I_4582 (I82989,I515,I82917,I83016,);
DFFARX1 I_4583 (I82674,I515,I82917,I83034,);
and I_4584 (I83043,I83034,I82737);
nor I_4585 (I83061,I83016,I83043);
DFFARX1 I_4586 (I83061,I515,I82917,I83088,);
nand I_4587 (I83097,I83034,I82737);
nand I_4588 (I83115,I82953,I83097);
not I_4589 (I83133,I83115);
DFFARX1 I_4590 (I82881,I515,I82917,I83160,);
DFFARX1 I_4591 (I83160,I515,I82917,I83178,);
nand I_4592 (I83187,I82386,I82863);
and I_4593 (I83205,I83187,I82530);
DFFARX1 I_4594 (I83205,I515,I82917,I83232,);
DFFARX1 I_4595 (I83232,I515,I82917,I83250,);
not I_4596 (I83259,I83250);
not I_4597 (I83277,I83232);
nand I_4598 (I83295,I83277,I83097);
nor I_4599 (I83313,I82530,I82863);
not I_4600 (I83331,I83313);
nor I_4601 (I83349,I83277,I83331);
nor I_4602 (I83367,I82953,I83349);
DFFARX1 I_4603 (I83367,I515,I82917,I83394,);
nor I_4604 (I83403,I83016,I83331);
nor I_4605 (I83421,I83232,I83403);
nor I_4606 (I83439,I83160,I83313);
nor I_4607 (I83457,I83016,I83313);
not I_4608 (I83475,I522);
DFFARX1 I_4609 (I83295,I515,I83475,I83502,);
DFFARX1 I_4610 (I83502,I515,I83475,I83520,);
not I_4611 (I83529,I83520);
not I_4612 (I83547,I83502);
DFFARX1 I_4613 (I83457,I515,I83475,I83574,);
not I_4614 (I83583,I83574);
and I_4615 (I83601,I83547,I83088);
not I_4616 (I83619,I83178);
nand I_4617 (I83637,I83619,I83088);
not I_4618 (I83655,I83439);
nor I_4619 (I83673,I83655,I83421);
nand I_4620 (I83691,I83673,I83133);
nor I_4621 (I83709,I83691,I83637);
DFFARX1 I_4622 (I83709,I515,I83475,I83736,);
not I_4623 (I83745,I83691);
not I_4624 (I83763,I83421);
nand I_4625 (I83781,I83763,I83088);
nor I_4626 (I83799,I83421,I83178);
nand I_4627 (I83817,I83601,I83799);
nand I_4628 (I83835,I83547,I83421);
nand I_4629 (I83853,I83655,I83088);
DFFARX1 I_4630 (I83853,I515,I83475,I83880,);
DFFARX1 I_4631 (I83853,I515,I83475,I83898,);
not I_4632 (I83907,I83088);
nor I_4633 (I83925,I83907,I83394);
and I_4634 (I83943,I83925,I83259);
or I_4635 (I83961,I83943,I83457);
DFFARX1 I_4636 (I83961,I515,I83475,I83988,);
nand I_4637 (I83997,I83988,I83619);
nor I_4638 (I84015,I83997,I83781);
nor I_4639 (I84033,I83988,I83583);
DFFARX1 I_4640 (I83988,I515,I83475,I84060,);
not I_4641 (I84069,I84060);
nor I_4642 (I84087,I84069,I83745);
not I_4643 (I84105,I522);
DFFARX1 I_4644 (I83736,I515,I84105,I84132,);
not I_4645 (I84141,I84132);
nand I_4646 (I84159,I84033,I83529);
and I_4647 (I84177,I84159,I83817);
DFFARX1 I_4648 (I84177,I515,I84105,I84204,);
not I_4649 (I84213,I84015);
DFFARX1 I_4650 (I83736,I515,I84105,I84240,);
not I_4651 (I84249,I84240);
nor I_4652 (I84267,I84249,I84141);
and I_4653 (I84285,I84267,I84015);
nor I_4654 (I84303,I84249,I84213);
nor I_4655 (I84321,I84204,I84303);
DFFARX1 I_4656 (I84087,I515,I84105,I84348,);
nor I_4657 (I84357,I84348,I84204);
not I_4658 (I84375,I84357);
not I_4659 (I84393,I84348);
nor I_4660 (I84411,I84393,I84285);
DFFARX1 I_4661 (I84411,I515,I84105,I84438,);
nand I_4662 (I84447,I84033,I83835);
and I_4663 (I84465,I84447,I83898);
DFFARX1 I_4664 (I84465,I515,I84105,I84492,);
nor I_4665 (I84501,I84492,I84348);
DFFARX1 I_4666 (I84501,I515,I84105,I84528,);
nand I_4667 (I84537,I84492,I84393);
nand I_4668 (I84555,I84375,I84537);
not I_4669 (I84573,I84492);
nor I_4670 (I84591,I84573,I84285);
DFFARX1 I_4671 (I84591,I515,I84105,I84618,);
nor I_4672 (I84627,I83880,I83835);
or I_4673 (I84645,I84348,I84627);
nor I_4674 (I84663,I84492,I84627);
or I_4675 (I84681,I84204,I84627);
DFFARX1 I_4676 (I84627,I515,I84105,I84708,);
not I_4677 (I84717,I522);
DFFARX1 I_4678 (I84528,I515,I84717,I84744,);
not I_4679 (I84753,I84744);
DFFARX1 I_4680 (I84645,I515,I84717,I84780,);
not I_4681 (I84789,I84663);
nand I_4682 (I84807,I84789,I84681);
not I_4683 (I84825,I84807);
nor I_4684 (I84843,I84825,I84555);
nor I_4685 (I84861,I84753,I84843);
DFFARX1 I_4686 (I84861,I515,I84717,I84888,);
not I_4687 (I84897,I84555);
nand I_4688 (I84915,I84897,I84825);
and I_4689 (I84933,I84897,I84663);
nand I_4690 (I84951,I84933,I84321);
nor I_4691 (I84969,I84951,I84897);
and I_4692 (I84987,I84780,I84951);
not I_4693 (I85005,I84951);
nand I_4694 (I85023,I84780,I85005);
nor I_4695 (I85041,I84744,I84951);
not I_4696 (I85059,I84618);
nor I_4697 (I85077,I85059,I84663);
nand I_4698 (I85095,I85077,I84897);
nor I_4699 (I85113,I84807,I85095);
nor I_4700 (I85131,I85059,I84528);
and I_4701 (I85149,I85131,I84438);
or I_4702 (I85167,I85149,I84708);
DFFARX1 I_4703 (I85167,I515,I84717,I85194,);
nor I_4704 (I85203,I85194,I84915);
DFFARX1 I_4705 (I85203,I515,I84717,I85230,);
DFFARX1 I_4706 (I85194,I515,I84717,I85248,);
not I_4707 (I85257,I85194);
nor I_4708 (I85275,I85257,I84780);
nor I_4709 (I85293,I85077,I85275);
DFFARX1 I_4710 (I85293,I515,I84717,I85320,);
not I_4711 (I85329,I522);
DFFARX1 I_4712 (I84969,I515,I85329,I85356,);
and I_4713 (I85365,I85356,I85041);
DFFARX1 I_4714 (I85365,I515,I85329,I85392,);
DFFARX1 I_4715 (I84888,I515,I85329,I85410,);
not I_4716 (I85419,I85023);
not I_4717 (I85437,I85230);
nand I_4718 (I85455,I85437,I85419);
nor I_4719 (I85473,I85410,I85455);
DFFARX1 I_4720 (I85455,I515,I85329,I85500,);
not I_4721 (I85509,I85500);
not I_4722 (I85527,I84987);
nand I_4723 (I85545,I85437,I85527);
DFFARX1 I_4724 (I85545,I515,I85329,I85572,);
not I_4725 (I85581,I85572);
not I_4726 (I85599,I85320);
nand I_4727 (I85617,I85599,I85248);
and I_4728 (I85635,I85419,I85617);
nor I_4729 (I85653,I85545,I85635);
DFFARX1 I_4730 (I85653,I515,I85329,I85680,);
DFFARX1 I_4731 (I85635,I515,I85329,I85698,);
nor I_4732 (I85707,I85320,I85230);
nor I_4733 (I85725,I85545,I85707);
or I_4734 (I85743,I85320,I85230);
nor I_4735 (I85761,I85113,I85041);
DFFARX1 I_4736 (I85761,I515,I85329,I85788,);
not I_4737 (I85797,I85788);
nor I_4738 (I85815,I85797,I85581);
nand I_4739 (I85833,I85797,I85410);
not I_4740 (I85851,I85113);
nand I_4741 (I85869,I85851,I85527);
nand I_4742 (I85887,I85797,I85869);
nand I_4743 (I85905,I85887,I85833);
nand I_4744 (I85923,I85869,I85743);
not I_4745 (I85941,I522);
DFFARX1 I_4746 (I85815,I515,I85941,I85968,);
not I_4747 (I85977,I85968);
nand I_4748 (I85995,I85680,I85725);
and I_4749 (I86013,I85995,I85392);
DFFARX1 I_4750 (I86013,I515,I85941,I86040,);
not I_4751 (I86049,I85905);
DFFARX1 I_4752 (I85923,I515,I85941,I86076,);
not I_4753 (I86085,I86076);
nor I_4754 (I86103,I86085,I85977);
and I_4755 (I86121,I86103,I85905);
nor I_4756 (I86139,I86085,I86049);
nor I_4757 (I86157,I86040,I86139);
DFFARX1 I_4758 (I85509,I515,I85941,I86184,);
nor I_4759 (I86193,I86184,I86040);
not I_4760 (I86211,I86193);
not I_4761 (I86229,I86184);
nor I_4762 (I86247,I86229,I86121);
DFFARX1 I_4763 (I86247,I515,I85941,I86274,);
nand I_4764 (I86283,I85473,I85473);
and I_4765 (I86301,I86283,I85680);
DFFARX1 I_4766 (I86301,I515,I85941,I86328,);
nor I_4767 (I86337,I86328,I86184);
DFFARX1 I_4768 (I86337,I515,I85941,I86364,);
nand I_4769 (I86373,I86328,I86229);
nand I_4770 (I86391,I86211,I86373);
not I_4771 (I86409,I86328);
nor I_4772 (I86427,I86409,I86121);
DFFARX1 I_4773 (I86427,I515,I85941,I86454,);
nor I_4774 (I86463,I85698,I85473);
or I_4775 (I86481,I86184,I86463);
nor I_4776 (I86499,I86328,I86463);
or I_4777 (I86517,I86040,I86463);
DFFARX1 I_4778 (I86463,I515,I85941,I86544,);
not I_4779 (I86553,I522);
DFFARX1 I_4780 (I86364,I515,I86553,I86580,);
not I_4781 (I86589,I86580);
nand I_4782 (I86607,I86499,I86364);
and I_4783 (I86625,I86607,I86481);
DFFARX1 I_4784 (I86625,I515,I86553,I86652,);
DFFARX1 I_4785 (I86652,I515,I86553,I86670,);
DFFARX1 I_4786 (I86391,I515,I86553,I86688,);
nand I_4787 (I86697,I86688,I86157);
not I_4788 (I86715,I86697);
DFFARX1 I_4789 (I86715,I515,I86553,I86742,);
not I_4790 (I86751,I86742);
nor I_4791 (I86769,I86589,I86751);
DFFARX1 I_4792 (I86544,I515,I86553,I86796,);
nor I_4793 (I86805,I86796,I86652);
nor I_4794 (I86823,I86796,I86715);
nand I_4795 (I86841,I86274,I86517);
and I_4796 (I86859,I86841,I86499);
DFFARX1 I_4797 (I86859,I515,I86553,I86886,);
not I_4798 (I86895,I86886);
nand I_4799 (I86913,I86895,I86796);
nand I_4800 (I86931,I86895,I86697);
nor I_4801 (I86949,I86454,I86517);
and I_4802 (I86967,I86796,I86949);
nor I_4803 (I86985,I86895,I86967);
DFFARX1 I_4804 (I86985,I515,I86553,I87012,);
nor I_4805 (I87021,I86580,I86949);
DFFARX1 I_4806 (I87021,I515,I86553,I87048,);
nor I_4807 (I87057,I86886,I86949);
not I_4808 (I87075,I87057);
nand I_4809 (I87093,I87075,I86913);
not I_4810 (I87111,I522);
DFFARX1 I_4811 (I87093,I515,I87111,I87138,);
DFFARX1 I_4812 (I87138,I515,I87111,I87156,);
not I_4813 (I87165,I87156);
nand I_4814 (I87183,I87048,I86769);
and I_4815 (I87201,I87183,I86823);
DFFARX1 I_4816 (I87201,I515,I87111,I87228,);
DFFARX1 I_4817 (I87228,I515,I87111,I87246,);
DFFARX1 I_4818 (I87228,I515,I87111,I87264,);
DFFARX1 I_4819 (I86823,I515,I87111,I87282,);
nand I_4820 (I87291,I87282,I86670);
not I_4821 (I87309,I87291);
nor I_4822 (I87327,I87138,I87309);
DFFARX1 I_4823 (I86805,I515,I87111,I87354,);
not I_4824 (I87363,I87354);
nor I_4825 (I87381,I87363,I87165);
nand I_4826 (I87399,I87363,I87291);
nand I_4827 (I87417,I86931,I87012);
and I_4828 (I87435,I87417,I87048);
DFFARX1 I_4829 (I87435,I515,I87111,I87462,);
nor I_4830 (I87471,I87462,I87138);
DFFARX1 I_4831 (I87471,I515,I87111,I87498,);
not I_4832 (I87507,I87462);
nor I_4833 (I87525,I86931,I87012);
not I_4834 (I87543,I87525);
nor I_4835 (I87561,I87291,I87543);
nor I_4836 (I87579,I87507,I87561);
DFFARX1 I_4837 (I87579,I515,I87111,I87606,);
nor I_4838 (I87615,I87462,I87543);
nor I_4839 (I87633,I87309,I87615);
nor I_4840 (I87651,I87462,I87525);
endmodule


