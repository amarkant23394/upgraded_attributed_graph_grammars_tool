module test_I15863(I11938,I1470,I13775,I15863);
input I11938,I1470,I13775;
output I15863;
wire I13908,I13743,I15832,I14162,I15628,I13749,I13891;
not I_0(I13908,I13891);
DFFARX1 I_1(I13891,I1470,I13775,,,I13743,);
nand I_2(I15832,I15628,I13749);
DFFARX1 I_3(I11938,I1470,I13775,,,I14162,);
not I_4(I15628,I13743);
nand I_5(I13749,I14162,I13908);
not I_6(I15863,I15832);
DFFARX1 I_7(I1470,I13775,,,I13891,);
endmodule


