module test_I2759_rst(I1477_rst,I2759_rst);
,I2759_rst);
input I1477_rst;
output I2759_rst;
wire ;
not I_0(I2759_rst,I1477_rst);
endmodule


