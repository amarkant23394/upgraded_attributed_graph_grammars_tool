module test_I16534(I1477,I1470,I16534);
input I1477,I1470;
output I16534;
wire I13361,I14901,I13162,I14335,I16240,I14808,I13248,I14370;
DFFARX1 I_0(I1470,,,I13361,);
DFFARX1 I_1(I14808,I1470,I14370,,,I14901,);
and I_2(I13162,I13248,I13361);
DFFARX1 I_3(I14335,I1470,I16240,,,I16534,);
and I_4(I14335,I14808,I14901);
not I_5(I16240,I1477);
DFFARX1 I_6(I13162,I1470,I14370,,,I14808,);
DFFARX1 I_7(I1470,,,I13248,);
not I_8(I14370,I1477);
endmodule


