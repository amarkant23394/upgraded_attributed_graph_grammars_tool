module test_I7173(I5266,I1477,I7105,I5070,I5368,I1470,I5642,I6924,I7173);
input I5266,I1477,I7105,I5070,I5368,I1470,I5642,I6924;
output I7173;
wire I5076,I7122,I7009,I7156,I6992,I5085,I6975,I6907,I5512,I5097,I7139;
nor I_0(I7173,I7156,I7009);
DFFARX1 I_1(I1470,,,I5076,);
and I_2(I7122,I7105,I5076);
not I_3(I7009,I6992);
DFFARX1 I_4(I7139,I1470,I6907,,,I7156,);
nand I_5(I6992,I6975,I5097);
nand I_6(I5085,I5512,I5266);
nor I_7(I6975,I6924,I5070);
not I_8(I6907,I1477);
DFFARX1 I_9(I1470,,,I5512,);
nand I_10(I5097,I5642,I5368);
or I_11(I7139,I7122,I5085);
endmodule


