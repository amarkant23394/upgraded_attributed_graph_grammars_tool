module test_final(IN_1_1_l_3,IN_2_1_l_3,IN_3_1_l_3,IN_1_8_l_3,IN_2_8_l_3,IN_3_8_l_3,IN_6_8_l_3,IN_1_10_l_3,IN_2_10_l_3,IN_3_10_l_3,IN_4_10_l_3,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1508_0_r_7,N6147_2_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7);
input IN_1_1_l_3,IN_2_1_l_3,IN_3_1_l_3,IN_1_8_l_3,IN_2_8_l_3,IN_3_8_l_3,IN_6_8_l_3,IN_1_10_l_3,IN_2_10_l_3,IN_3_10_l_3,IN_4_10_l_3,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1508_0_r_7,N6147_2_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7;
wire N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1372_10_r_3,N1508_10_r_3,N3_8_l_3,n39_3,n_431_5_r_3,n22_3,n23_3,n24_3,n25_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,N1371_0_r_7,N1507_6_r_7,N1508_6_r_7,n_431_5_r_7,n4_7,n19_7,n20_7,n21_7,n22_7,n23_7,n24_7,n25_7,n26_7,n27_7,n28_7,n29_7,n30_7,n31_7,n32_7;
nor I_0(N1371_0_r_3,n39_3,n37_3);
nor I_1(N1508_0_r_3,n25_3,n37_3);
nor I_2(N6147_3_r_3,N1372_10_r_3,n33_3);
nand I_3(n_429_or_0_5_r_3,N1372_10_r_3,n30_3);
DFFARX1 I_4(n_431_5_r_3,blif_clk_net_5_r_7,n4_7,G78_5_r_3,);
nand I_5(n_576_5_r_3,n22_3,n23_3);
not I_6(n_102_5_r_3,n39_3);
nand I_7(n_547_5_r_3,n26_3,n27_3);
not I_8(N1372_10_r_3,n36_3);
nor I_9(N1508_10_r_3,n35_3,n36_3);
and I_10(N3_8_l_3,IN_6_8_l_3,n34_3);
DFFARX1 I_11(N3_8_l_3,blif_clk_net_5_r_7,n4_7,n39_3,);
nand I_12(n_431_5_r_3,n29_3,n30_3);
nor I_13(n22_3,n24_3,n25_3);
nor I_14(n23_3,IN_3_1_l_3,n39_3);
not I_15(n24_3,n27_3);
nand I_16(n25_3,IN_1_1_l_3,IN_2_1_l_3);
nor I_17(n26_3,n39_3,n28_3);
nor I_18(n27_3,IN_1_8_l_3,IN_3_8_l_3);
not I_19(n28_3,n37_3);
nand I_20(n29_3,N1372_10_r_3,n39_3);
nand I_21(n30_3,n31_3,n32_3);
not I_22(n31_3,n25_3);
not I_23(n32_3,IN_3_1_l_3);
nand I_24(n33_3,n24_3,n25_3);
nand I_25(n34_3,IN_2_8_l_3,IN_3_8_l_3);
nor I_26(n35_3,n27_3,n31_3);
nand I_27(n36_3,n28_3,n38_3);
nand I_28(n37_3,IN_1_10_l_3,IN_2_10_l_3);
or I_29(n38_3,IN_3_10_l_3,IN_4_10_l_3);
nor I_30(N1371_0_r_7,n22_7,n24_7);
nor I_31(N1508_0_r_7,n24_7,n28_7);
nor I_32(N6147_2_r_7,n21_7,n26_7);
nand I_33(n_429_or_0_5_r_7,n19_7,n24_7);
DFFARX1 I_34(n_431_5_r_7,blif_clk_net_5_r_7,n4_7,G78_5_r_7,);
nand I_35(n_576_5_r_7,N1371_0_r_7,n19_7);
not I_36(n_102_5_r_7,n22_7);
nand I_37(n_547_5_r_7,n20_7,n21_7);
nor I_38(N1507_6_r_7,n22_7,n27_7);
nor I_39(N1508_6_r_7,n27_7,N6147_3_r_3);
nand I_40(n_431_5_r_7,n24_7,n25_7);
not I_41(n4_7,blif_reset_net_5_r_7);
nor I_42(n19_7,n30_7,n_547_5_r_3);
nor I_43(n20_7,n22_7,n23_7);
not I_44(n21_7,n29_7);
nor I_45(n22_7,n29_7,n31_7);
not I_46(n23_7,n27_7);
not I_47(n24_7,N1508_6_r_7);
nand I_48(n25_7,N1507_6_r_7,n19_7);
or I_49(n26_7,n19_7,n23_7);
nand I_50(n27_7,N1371_0_r_3,n_429_or_0_5_r_3);
nor I_51(n28_7,n19_7,n21_7);
nand I_52(n29_7,n_576_5_r_3,N1371_0_r_3);
or I_53(n30_7,G78_5_r_3,N1508_10_r_3);
nor I_54(n31_7,n32_7,n_102_5_r_3);
and I_55(n32_7,N1508_0_r_3,N6147_3_r_3);
endmodule


