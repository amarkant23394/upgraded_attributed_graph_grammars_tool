module test_I7088(I1477,I5546,I1470,I7088);
input I1477,I5546,I1470;
output I7088;
wire I5659,I5625,I5088,I5563,I5512,I5105,I5642;
or I_0(I5659,I5642,I5563);
DFFARX1 I_1(I1470,I5105,,,I5625,);
DFFARX1 I_2(I5659,I1470,I5105,,,I5088,);
and I_3(I5563,I5512,I5546);
DFFARX1 I_4(I1470,I5105,,,I5512,);
not I_5(I7088,I5088);
not I_6(I5105,I1477);
not I_7(I5642,I5625);
endmodule


