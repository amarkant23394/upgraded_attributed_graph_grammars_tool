module test_I11830(I1477,I1470,I6896,I11830);
input I1477,I1470,I6896;
output I11830;
wire I9320,I8854,I11813,I9303,I9179,I8862,I11310;
not I_0(I9320,I9303);
nor I_1(I8854,I9179,I9320);
DFFARX1 I_2(I8854,I1470,I11310,,,I11813,);
not I_3(I11830,I11813);
DFFARX1 I_4(I1470,I8862,,,I9303,);
DFFARX1 I_5(I6896,I1470,I8862,,,I9179,);
not I_6(I8862,I1477);
not I_7(I11310,I1477);
endmodule


