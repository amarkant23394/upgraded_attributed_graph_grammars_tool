module test_I15764(I1477,I11938,I1470,I13809,I14066,I15764);
input I1477,I11938,I1470,I13809,I14066;
output I15764;
wire I13826,I13908,I14004,I15747,I14162,I13737,I14114,I13749,I13775,I13891,I14131;
DFFARX1 I_0(I13809,I1470,I13775,,,I13826,);
not I_1(I13908,I13891);
DFFARX1 I_2(I1470,I13775,,,I14004,);
not I_3(I15747,I13749);
nor I_4(I15764,I15747,I13737);
DFFARX1 I_5(I11938,I1470,I13775,,,I14162,);
DFFARX1 I_6(I14131,I1470,I13775,,,I13737,);
nand I_7(I14114,I14066,I14004);
nand I_8(I13749,I14162,I13908);
not I_9(I13775,I1477);
DFFARX1 I_10(I1470,I13775,,,I13891,);
and I_11(I14131,I13826,I14114);
endmodule


