module test_I16086(I1477,I14278,I13987,I13809,I1470,I16086);
input I1477,I14278,I13987,I13809,I1470;
output I16086;
wire I15645,I14004,I13860,I15662,I13891,I16052,I13775,I15611,I13761,I13752,I13740,I13764,I16069,I13826,I14162;
nor I_0(I15645,I13761,I13740);
DFFARX1 I_1(I13987,I1470,I13775,,,I14004,);
nor I_2(I13860,I13826);
nand I_3(I15662,I15645,I13764);
DFFARX1 I_4(I1470,I13775,,,I13891,);
DFFARX1 I_5(I13752,I1470,I15611,,,I16052,);
not I_6(I13775,I1477);
not I_7(I15611,I1477);
nand I_8(I13761,I13891,I13860);
DFFARX1 I_9(I14278,I1470,I13775,,,I13752,);
DFFARX1 I_10(I14162,I1470,I13775,,,I13740,);
nor I_11(I13764,I14004,I13826);
not I_12(I16069,I16052);
DFFARX1 I_13(I13809,I1470,I13775,,,I13826,);
nor I_14(I16086,I16069,I15662);
DFFARX1 I_15(I1470,I13775,,,I14162,);
endmodule


