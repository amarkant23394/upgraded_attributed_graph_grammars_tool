module test_final(G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3,n4_1_l_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n4_1_r_3,blif_clk_net_1_r_4,n6_4,G42_1_r_3,);
nor I_1(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_2(n_573_1_r_3,n26_3,n27_3);
nor I_3(n_549_1_r_3,n40_3,n32_3);
nand I_4(n_569_1_r_3,n27_3,n31_3);
and I_5(n_452_1_r_3,G18_1_l_3,n26_3);
nor I_6(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_7(N3_2_r_3,blif_clk_net_1_r_4,n6_4,G199_2_r_3,);
DFFARX1 I_8(n_572_1_l_3,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_3,);
nor I_9(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_10(n4_1_l_3,G18_1_l_3,IN_1_1_l_3);
DFFARX1 I_11(n4_1_l_3,blif_clk_net_1_r_4,n6_4,G42_1_l_3,);
not I_12(n22_3,G42_1_l_3);
DFFARX1 I_13(IN_1_3_l_3,blif_clk_net_1_r_4,n6_4,n40_3,);
DFFARX1 I_14(IN_2_3_l_3,blif_clk_net_1_r_4,n6_4,n25_internal_3,);
not I_15(n25_3,n25_internal_3);
nor I_16(n4_1_r_3,n40_3,n36_3);
nor I_17(N3_2_r_3,n26_3,n37_3);
nor I_18(n_572_1_l_3,G15_1_l_3,IN_7_1_l_3);
DFFARX1 I_19(G42_1_l_3,blif_clk_net_1_r_4,n6_4,ACVQN1_3_r_3,);
nor I_20(n26_3,IN_5_1_l_3,IN_9_1_l_3);
not I_21(n27_3,IN_10_1_l_3);
nor I_22(n28_3,IN_10_1_l_3,n29_3);
nor I_23(n29_3,G15_1_l_3,n30_3);
not I_24(n30_3,IN_4_1_l_3);
nor I_25(n31_3,IN_9_1_l_3,n40_3);
nor I_26(n32_3,n25_3,n33_3);
nand I_27(n33_3,IN_4_3_l_3,n22_3);
or I_28(n34_3,IN_9_1_l_3,IN_10_1_l_3);
nand I_29(n35_3,IN_4_3_l_3,ACVQN1_3_r_3);
nor I_30(n36_3,G18_1_l_3,IN_5_1_l_3);
nor I_31(n37_3,n38_3,n39_3);
not I_32(n38_3,n_572_1_l_3);
nand I_33(n39_3,n27_3,n30_3);
DFFARX1 I_34(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_35(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_36(n_573_1_r_4,n16_4,G42_1_r_3);
nor I_37(n_549_1_r_4,n22_4,n23_4);
nand I_38(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_39(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_40(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_41(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_42(P6_5_r_4,P6_5_r_internal_4);
or I_43(n_431_0_l_4,n26_4,G42_1_r_3);
not I_44(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_45(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_46(n_452_1_r_3,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_47(n16_4,ACVQN1_5_l_4);
DFFARX1 I_48(n_572_1_r_3,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_49(n17_4,n17_internal_4);
nor I_50(n4_1_r_4,n30_4,n31_4);
nand I_51(n19_4,n33_4,n_549_1_r_3);
DFFARX1 I_52(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_53(n15_4,n15_internal_4);
DFFARX1 I_54(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_55(n20_4,n16_4,n_42_2_r_3);
nor I_56(n21_4,G199_2_r_3,G42_1_r_3);
nand I_57(n22_4,G78_0_l_4,n25_4);
nand I_58(n23_4,n24_4,n_42_2_r_3);
not I_59(n24_4,G42_1_r_3);
not I_60(n25_4,G199_2_r_3);
and I_61(n26_4,n27_4,n_569_1_r_3);
nor I_62(n27_4,n28_4,n_573_1_r_3);
not I_63(n28_4,n_549_1_r_3);
not I_64(n29_4,n30_4);
nand I_65(n30_4,n32_4,n_266_and_0_3_r_3);
nand I_66(n31_4,n25_4,n_42_2_r_3);
nor I_67(n32_4,n33_4,G42_1_r_3);
not I_68(n33_4,ACVQN2_3_r_3);
endmodule


