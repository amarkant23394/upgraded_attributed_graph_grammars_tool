module test_I6826(I2742,I4017,I2727,I1477,I1470,I6826);
input I2742,I4017,I2727,I1477,I1470;
output I6826;
wire I6781,I3975,I3954,I6442,I6329,I4113,I4308,I4068,I4034,I4130,I3957,I2724,I3983;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
nor I_1(I3975,I4308,I4034);
not I_2(I3954,I4068);
nand I_3(I6826,I6781,I6442);
nor I_4(I6442,I3975,I3954);
not I_5(I6329,I1477);
DFFARX1 I_6(I1470,I3983,,,I4113,);
DFFARX1 I_7(I2727,I1470,I3983,,,I4308,);
nor I_8(I4068,I2742,I2724);
DFFARX1 I_9(I4017,I1470,I3983,,,I4034,);
nor I_10(I4130,I4113,I4068);
nand I_11(I3957,I4308,I4130);
DFFARX1 I_12(I1470,,,I2724,);
not I_13(I3983,I1477);
endmodule


