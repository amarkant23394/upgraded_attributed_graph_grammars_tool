module test_I17696(I1477,I1470,I15573,I17611,I17696);
input I1477,I1470,I15573,I17611;
output I17696;
wire I15582,I17413,I17628,I17645,I17662,I15928;
not I_0(I15582,I15928);
not I_1(I17413,I1477);
and I_2(I17628,I17611,I15573);
or I_3(I17645,I17628,I15582);
DFFARX1 I_4(I17662,I1470,I17413,,,I17696,);
DFFARX1 I_5(I17645,I1470,I17413,,,I17662,);
DFFARX1 I_6(I1470,,,I15928,);
endmodule


