module test_final(IN_1_0_l,IN_2_0_l,IN_3_0_l,IN_4_0_l,IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,blif_clk_net_8_r,blif_reset_net_8_r,N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r,N1372_10_r,N1508_10_r);
input IN_1_0_l,IN_2_0_l,IN_3_0_l,IN_4_0_l,IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,blif_clk_net_8_r,blif_reset_net_8_r;
output N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r,N1372_10_r,N1508_10_r;
wire N1371_0_l,N1508_0_l,n3_0_l,n4_0_l,N1372_1_l,N1508_1_l,n4_1_l,N6147_2_l,n5_2_l,n6_2_l,N6138_2_l,n7_2_l,N6147_3_l,n3_3_l,N6138_3_l,n3_0_r,n4_0_r,n4_1_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,N3_8_r,n1_8_r,n3_8_r,N6150_9_r,n3_9_r,n5_10_r,n6_10_r;
nor I_0(N1371_0_l,IN_2_0_l,n4_0_l);
nor I_1(N1508_0_l,n3_0_l,n4_0_l);
nor I_2(n3_0_l,IN_3_0_l,IN_4_0_l);
not I_3(n4_0_l,IN_1_0_l);
not I_4(N1372_1_l,n4_1_l);
nor I_5(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_6(n4_1_l,IN_1_1_l,IN_2_1_l);
nor I_7(N6147_2_l,n5_2_l,n6_2_l);
nor I_8(n5_2_l,IN_5_2_l,n7_2_l);
not I_9(n6_2_l,N6138_2_l);
nor I_10(N6138_2_l,IN_1_2_l,IN_2_2_l);
nor I_11(n7_2_l,IN_3_2_l,IN_4_2_l);
nor I_12(N6147_3_l,IN_3_3_l,n3_3_l);
not I_13(n3_3_l,N6138_3_l);
nor I_14(N6138_3_l,IN_1_3_l,IN_2_3_l);
nor I_15(N1371_0_r,n4_0_r,N6147_2_l);
nor I_16(N1508_0_r,n3_0_r,n4_0_r);
nor I_17(n3_0_r,N1508_0_l,N6147_3_l);
not I_18(n4_0_r,N6147_3_l);
not I_19(N1372_1_r,n4_1_r);
nor I_20(N1508_1_r,n4_1_r,N1508_1_l);
nand I_21(n4_1_r,N1371_0_l,N1372_1_l);
nor I_22(N1507_6_r,n8_6_r,n9_6_r);
and I_23(N1508_6_r,n6_6_r,N1508_1_l);
nor I_24(n6_6_r,n7_6_r,n8_6_r);
not I_25(n7_6_r,N1508_0_l);
nor I_26(n8_6_r,n9_6_r,N1372_1_l);
and I_27(n9_6_r,N1508_1_l,N1371_0_l);
nor I_28(n_42_8_r,N6147_2_l,N6147_3_l);
DFFARX1 I_29(N3_8_r,blif_clk_net_8_r,n1_8_r,G199_8_r,);
and I_30(N3_8_r,n3_8_r,N1371_0_l);
not I_31(n1_8_r,blif_reset_net_8_r);
nand I_32(n3_8_r,N1371_0_l,N6147_2_l);
not I_33(N6150_9_r,N1508_1_l);
nor I_34(N6147_9_r,N6150_9_r,n3_9_r);
nor I_35(N6134_9_r,n3_9_r,N6147_2_l);
nor I_36(n3_9_r,N1508_0_l,N1371_0_l);
buf I_37(I_BUFF_1_9_r,N1372_1_l);
not I_38(N1372_10_r,n6_10_r);
nor I_39(N1508_10_r,n5_10_r,n6_10_r);
nor I_40(n5_10_r,N6147_3_l,N6147_2_l);
nand I_41(n6_10_r,N1508_0_l,N1372_1_l);
endmodule


