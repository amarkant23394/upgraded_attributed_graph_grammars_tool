module test_I7669(I3963,I6826,I6346,I1477,I1470,I7669);
input I3963,I6826,I6346,I1477,I1470;
output I7669;
wire I6606,I6297,I7652,I7587,I6380,I6843,I6329,I6318,I6363,I6493,I6300;
DFFARX1 I_0(I1470,I6329,,,I6606,);
DFFARX1 I_1(I6843,I1470,I6329,,,I6297,);
nor I_2(I7652,I7587,I6297);
not I_3(I7587,I6300);
DFFARX1 I_4(I6363,I1470,I6329,,,I6380,);
and I_5(I6843,I6493,I6826);
not I_6(I6329,I1477);
not I_7(I6318,I6380);
and I_8(I6363,I6346,I3963);
DFFARX1 I_9(I1470,I6329,,,I6493,);
DFFARX1 I_10(I6606,I1470,I6329,,,I6300,);
nand I_11(I7669,I7652,I6318);
endmodule


