module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_8,n8_8,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_8,n8_8,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_8,n8_8,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_8,n8_8,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_8,n8_8,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_8,n8_8,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_8,n8_8,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_32(n_572_1_r_8,n39_8,n23_8);
and I_33(n_549_1_r_8,n38_8,n23_8);
nand I_34(n_569_1_r_8,n38_8,n24_8);
nor I_35(n_452_1_r_8,n25_8,n26_8);
nor I_36(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_37(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_38(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_39(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_40(n_431_0_l_8,n29_8,n_549_1_r_14);
not I_41(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_42(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_43(n19_8,G78_0_l_8);
DFFARX1 I_44(P6_5_r_14,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_45(n22_8,n39_8);
DFFARX1 I_46(n_572_1_r_14,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_47(n4_1_r_8,G78_0_l_8,n33_8);
nor I_48(N3_2_r_8,n22_8,n35_8);
nor I_49(N1_4_r_8,n27_8,n37_8);
nand I_50(n23_8,n32_8,n_573_1_r_14);
not I_51(n24_8,n23_8);
nand I_52(n25_8,n36_8,n_572_1_r_14);
nand I_53(n26_8,n27_8,n28_8);
nor I_54(n27_8,n31_8,G42_1_r_14);
not I_55(n28_8,ACVQN1_5_r_14);
and I_56(n29_8,n30_8,G42_1_r_14);
nor I_57(n30_8,n31_8,n_42_2_r_14);
not I_58(n31_8,n_569_1_r_14);
and I_59(n32_8,n28_8,G42_1_r_14);
nand I_60(n33_8,n28_8,n34_8);
not I_61(n34_8,n25_8);
nor I_62(n35_8,n34_8,ACVQN1_5_r_14);
not I_63(n36_8,G199_2_r_14);
nor I_64(n37_8,n19_8,n38_8);
endmodule


