module test_I9114(I6975,I7427,I7026,I5097,I9114);
input I6975,I7427,I7026,I5097;
output I9114;
wire I6992,I7317,I7057,I6881,I8879,I6887,I9083;
nand I_0(I6992,I6975,I5097);
nor I_1(I7317,I7057);
not I_2(I9114,I9083);
not I_3(I7057,I7026);
nand I_4(I6881,I6992,I7057);
not I_5(I8879,I6887);
nand I_6(I6887,I7427,I7317);
nand I_7(I9083,I8879,I6881);
endmodule


