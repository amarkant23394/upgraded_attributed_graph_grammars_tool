module test_I16226(I14667,I1477,I16435,I14335,I1470,I14588,I16226);
input I14667,I1477,I16435,I14335,I1470,I14588;
output I16226;
wire I14362,I14344,I16469,I16644,I16551,I14715,I16452,I14537,I14370,I16568,I16534,I14347,I16240,I14777;
DFFARX1 I_0(I1470,I14370,,,I14362,);
nand I_1(I14344,I14537,I14715);
DFFARX1 I_2(I16452,I1470,I16240,,,I16469,);
DFFARX1 I_3(I14347,I1470,I16240,,,I16644,);
and I_4(I16551,I16534,I14344);
not I_5(I14715,I14667);
nand I_6(I16226,I16644,I16568);
and I_7(I16452,I16435,I14362);
DFFARX1 I_8(I1470,I14370,,,I14537,);
not I_9(I14370,I1477);
nor I_10(I16568,I16551,I16469);
DFFARX1 I_11(I14335,I1470,I16240,,,I16534,);
DFFARX1 I_12(I14777,I1470,I14370,,,I14347,);
not I_13(I16240,I1477);
or I_14(I14777,I14667,I14588);
endmodule


