module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_10,blif_reset_net_1_r_10,G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_10,blif_reset_net_1_r_10;
output G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_452_1_r_10,N3_2_l_10,n4_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_10,n4_10,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_10,n4_10,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_10,n4_10,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_10,n4_10,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_10,n4_10,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_10,n4_10,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_10,n4_10,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_10,n4_10,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_10,blif_clk_net_1_r_10,n4_10,G42_1_r_10,);
nor I_33(n_572_1_r_10,n26_10,n3_10);
nand I_34(n_573_1_r_10,n16_10,n18_10);
nand I_35(n_549_1_r_10,n19_10,n20_10);
nor I_36(n_452_1_r_10,n25_10,n21_10);
nor I_37(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_38(N3_2_r_10,blif_clk_net_1_r_10,n4_10,G199_2_r_10,);
DFFARX1 I_39(G199_4_l_10,blif_clk_net_1_r_10,n4_10,ACVQN2_3_r_10,);
nor I_40(n_266_and_0_3_r_10,n17_10,n13_10);
and I_41(N3_2_l_10,n23_10,n_572_1_r_16);
not I_42(n4_10,blif_reset_net_1_r_10);
DFFARX1 I_43(N3_2_l_10,blif_clk_net_1_r_10,n4_10,n25_10,);
not I_44(n16_10,n25_10);
DFFARX1 I_45(n_569_1_r_16,blif_clk_net_1_r_10,n4_10,n26_10,);
DFFARX1 I_46(P6_5_r_16,blif_clk_net_1_r_10,n4_10,ACVQN1_3_l_10,);
and I_47(N1_4_l_10,n24_10,n_573_1_r_16);
DFFARX1 I_48(N1_4_l_10,blif_clk_net_1_r_10,n4_10,G199_4_l_10,);
DFFARX1 I_49(n_452_1_r_16,blif_clk_net_1_r_10,n4_10,n27_10,);
not I_50(n17_10,n27_10);
nor I_51(n4_1_r_10,n27_10,n21_10);
nor I_52(N3_2_r_10,n16_10,n22_10);
not I_53(n3_10,n18_10);
DFFARX1 I_54(n3_10,blif_clk_net_1_r_10,n4_10,n13_internal_10,);
not I_55(n13_10,n13_internal_10);
nand I_56(n18_10,ACVQN1_3_l_10,G42_1_r_16);
not I_57(n19_10,n_452_1_r_10);
nand I_58(n20_10,n16_10,n26_10);
nor I_59(n21_10,G199_4_r_16,ACVQN1_5_r_16);
and I_60(n22_10,n26_10,n21_10);
nand I_61(n23_10,n_549_1_r_16,ACVQN1_5_r_16);
nand I_62(n24_10,G214_4_r_16,G42_1_r_16);
endmodule


