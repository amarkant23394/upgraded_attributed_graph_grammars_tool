module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_8_r_8,n8_8,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N1371_0_r_8,n46_8,n51_8);
not I_36(N1508_0_r_8,n46_8);
nor I_37(N1372_1_r_8,n37_8,n49_8);
and I_38(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_39(N1507_6_r_8,n47_8,n48_8);
nor I_40(N1508_6_r_8,n37_8,n38_8);
nor I_41(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_42(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_43(N6147_9_r_8,n29_8,n30_8);
nor I_44(N6134_9_r_8,n30_8,n31_8);
not I_45(I_BUFF_1_9_r_8,n35_8);
nor I_46(N1372_10_r_8,n46_8,n49_8);
nor I_47(N1508_10_r_8,n40_8,n41_8);
and I_48(N3_8_l_8,n36_8,N1508_6_r_4);
not I_49(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_50(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_51(n29_8,n53_8);
nor I_52(N3_8_r_8,n33_8,n34_8);
and I_53(n30_8,n32_8,n33_8);
nor I_54(n31_8,N1371_0_r_4,n_569_7_r_4);
nand I_55(n32_8,n42_8,N1508_6_r_4);
or I_56(n33_8,n46_8,N1507_6_r_4);
nor I_57(n34_8,n32_8,n35_8);
nand I_58(n35_8,n44_8,n_452_7_r_4);
nand I_59(n36_8,n_569_7_r_4,N1507_6_r_4);
not I_60(n37_8,n31_8);
nand I_61(n38_8,N1508_0_r_8,n39_8);
nand I_62(n39_8,n33_8,n50_8);
and I_63(n40_8,n32_8,n35_8);
not I_64(n41_8,N1372_10_r_8);
and I_65(n42_8,n43_8,n_572_7_r_4);
nand I_66(n43_8,n44_8,n45_8);
nand I_67(n44_8,n_572_7_r_4,G42_7_r_4);
not I_68(n45_8,n_452_7_r_4);
nand I_69(n46_8,G42_7_r_4,n_549_7_r_4);
not I_70(n47_8,n39_8);
nor I_71(n48_8,n35_8,n49_8);
not I_72(n49_8,n51_8);
nand I_73(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_74(n51_8,n52_8,N1371_0_r_4);
or I_75(n52_8,n_549_7_r_4,N6134_9_r_4);
endmodule


