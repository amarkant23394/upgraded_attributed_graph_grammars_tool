module test_final(IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_7_r_14,blif_reset_net_7_r_14,N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14);
input IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_7_r_14,blif_reset_net_7_r_14;
output N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14;
wire N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_102_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13,n4_7_l_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13,I_BUFF_1_9_r_14,N3_8_l_14,n8_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14;
nor I_0(N1371_0_r_13,n59_13,n61_13);
nor I_1(N1508_0_r_13,n59_13,n60_13);
not I_2(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_3(n_431_5_r_13,blif_clk_net_7_r_14,n8_14,G78_5_r_13,);
nand I_4(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_5(n_102_5_r_13,IN_9_7_l_13,IN_10_7_l_13);
nand I_6(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_7(n1_13,blif_clk_net_7_r_14,n8_14,G42_7_r_13,);
nor I_8(n_572_7_r_13,n40_13,n41_13);
nand I_9(n_573_7_r_13,n37_13,n38_13);
nor I_10(n_549_7_r_13,n46_13,n47_13);
nand I_11(n_569_7_r_13,n37_13,n43_13);
nand I_12(n_452_7_r_13,n52_13,n53_13);
nor I_13(n4_7_l_13,G18_7_l_13,IN_1_7_l_13);
DFFARX1 I_14(n4_7_l_13,blif_clk_net_7_r_14,n8_14,n62_13,);
not I_15(n33_13,n62_13);
nand I_16(n_431_5_r_13,n54_13,n55_13);
not I_17(n1_13,n52_13);
nor I_18(n34_13,n35_13,n36_13);
nor I_19(n35_13,G15_7_l_13,n42_13);
nand I_20(n36_13,n50_13,n58_13);
nand I_21(n37_13,n44_13,n45_13);
or I_22(n38_13,IN_3_1_l_13,n39_13);
nand I_23(n39_13,IN_1_1_l_13,IN_2_1_l_13);
not I_24(n40_13,n36_13);
nor I_25(n41_13,IN_10_7_l_13,n35_13);
not I_26(n42_13,IN_4_7_l_13);
or I_27(n43_13,G18_7_l_13,IN_5_7_l_13);
not I_28(n44_13,G15_7_l_13);
not I_29(n45_13,IN_7_7_l_13);
nor I_30(n46_13,n39_13,n40_13);
nor I_31(n47_13,G18_7_l_13,IN_5_7_l_13);
nor I_32(n48_13,n50_13,n51_13);
nor I_33(n49_13,G15_7_l_13,IN_7_7_l_13);
not I_34(n50_13,n59_13);
not I_35(n51_13,n_102_5_r_13);
nand I_36(n52_13,n33_13,n39_13);
nand I_37(n53_13,IN_3_1_l_13,n33_13);
nor I_38(n54_13,IN_5_7_l_13,IN_9_7_l_13);
nand I_39(n55_13,n62_13,n56_13);
nor I_40(n56_13,n39_13,n57_13);
not I_41(n57_13,G18_7_l_13);
or I_42(n58_13,IN_3_10_l_13,IN_4_10_l_13);
nand I_43(n59_13,IN_1_10_l_13,IN_2_10_l_13);
nor I_44(n60_13,IN_5_7_l_13,n51_13);
nor I_45(n61_13,IN_3_1_l_13,n39_13);
nor I_46(N1371_0_r_14,n47_14,n30_14);
nor I_47(N1508_0_r_14,n30_14,n41_14);
nor I_48(N1507_6_r_14,n37_14,n44_14);
nor I_49(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_50(n4_7_r_14,blif_clk_net_7_r_14,n8_14,G42_7_r_14,);
nor I_51(n_572_7_r_14,n28_14,n29_14);
nand I_52(n_573_7_r_14,n26_14,n27_14);
nor I_53(n_549_7_r_14,n31_14,n32_14);
nand I_54(n_569_7_r_14,n26_14,n30_14);
nor I_55(n_452_7_r_14,n47_14,n28_14);
nor I_56(N6147_9_r_14,n36_14,n37_14);
nor I_57(N6134_9_r_14,n28_14,n36_14);
not I_58(I_BUFF_1_9_r_14,n26_14);
and I_59(N3_8_l_14,n38_14,n_576_5_r_13);
not I_60(n8_14,blif_reset_net_7_r_14);
DFFARX1 I_61(N3_8_l_14,blif_clk_net_7_r_14,n8_14,n47_14,);
nor I_62(n4_7_r_14,n47_14,n35_14);
nand I_63(n26_14,G78_5_r_13,n_429_or_0_5_r_13);
not I_64(n27_14,n28_14);
nor I_65(n28_14,n43_14,n_569_7_r_13);
not I_66(n29_14,n33_14);
not I_67(n30_14,n31_14);
nor I_68(n31_14,n46_14,N1508_0_r_13);
and I_69(n32_14,n33_14,n34_14);
nand I_70(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_71(n34_14,n42_14,n43_14);
nor I_72(n35_14,n_547_5_r_13,G42_7_r_13);
nor I_73(n36_14,n47_14,n34_14);
not I_74(n37_14,n35_14);
nand I_75(n38_14,n_429_or_0_5_r_13,G42_7_r_13);
nand I_76(n39_14,n29_14,n40_14);
nand I_77(n40_14,n27_14,n37_14);
nor I_78(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_79(n42_14,n_573_7_r_13,n_549_7_r_13);
not I_80(n43_14,n_572_7_r_13);
nor I_81(n44_14,n27_14,n33_14);
or I_82(n45_14,N1371_0_r_13,N1508_0_r_13);
or I_83(n46_14,n_452_7_r_13,G78_5_r_13);
endmodule


