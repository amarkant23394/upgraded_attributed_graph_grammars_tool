module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_8_r_10,n11_10,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_8_r_10,n11_10,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N1371_0_r_10,n37_10,n38_10);
nor I_41(N1508_0_r_10,n37_10,n58_10);
nand I_42(N6147_2_r_10,n39_10,n40_10);
not I_43(N6147_3_r_10,n39_10);
nor I_44(N1372_4_r_10,n46_10,n49_10);
nor I_45(N1508_4_r_10,n51_10,n52_10);
nor I_46(N1507_6_r_10,n49_10,n60_10);
nor I_47(N1508_6_r_10,n49_10,n50_10);
nor I_48(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_49(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_50(N6147_9_r_10,n36_10,n37_10);
nor I_51(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_52(I_BUFF_1_9_r_10,n48_10);
nor I_53(N3_8_r_10,n44_10,n47_10);
not I_54(n11_10,blif_reset_net_8_r_10);
not I_55(n35_10,n49_10);
nor I_56(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_57(n37_10,N1371_0_r_16);
not I_58(n38_10,n46_10);
nand I_59(n39_10,n43_10,n44_10);
nand I_60(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_61(n41_10,n42_10,N1371_0_r_16);
not I_62(n42_10,n44_10);
nor I_63(n43_10,n45_10,N1371_0_r_16);
nand I_64(n44_10,n54_10,N1372_1_r_16);
nor I_65(n45_10,n59_10,N1508_1_r_16);
nand I_66(n46_10,n61_10,n_569_7_r_16);
nor I_67(n47_10,n46_10,n48_10);
nand I_68(n48_10,n62_10,n63_10);
nand I_69(n49_10,n56_10,N1508_6_r_16);
not I_70(n50_10,n45_10);
nor I_71(n51_10,n42_10,n53_10);
not I_72(n52_10,N1372_4_r_10);
nor I_73(n53_10,n48_10,n50_10);
and I_74(n54_10,n55_10,n_573_7_r_16);
nand I_75(n55_10,n56_10,n57_10);
nand I_76(n56_10,N1507_6_r_16,n_452_7_r_16);
not I_77(n57_10,N1508_6_r_16);
nor I_78(n58_10,n35_10,n45_10);
nor I_79(n59_10,G42_7_r_16,n_572_7_r_16);
nor I_80(n60_10,n37_10,n46_10);
or I_81(n61_10,G42_7_r_16,n_572_7_r_16);
nor I_82(n62_10,N1508_0_r_16,N1372_1_r_16);
or I_83(n63_10,n64_10,N1508_0_r_16);
nor I_84(n64_10,N6147_2_r_16,N1371_0_r_16);
endmodule


