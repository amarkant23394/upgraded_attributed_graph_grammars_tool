module test_I10026(I7562,I7547,I1477,I1470,I7731,I7669,I10026);
input I7562,I7547,I1477,I1470,I7731,I7669;
output I10026;
wire I10349,I7550,I10219,I7570,I10185,I10397,I7977,I7541,I10052,I10202,I7532,I10332;
and I_0(I10349,I10332,I7550);
nand I_1(I7550,I7977,I7731);
DFFARX1 I_2(I10202,I1470,I10052,,,I10219,);
not I_3(I7570,I1477);
nand I_4(I10185,I7547,I7562);
not I_5(I10397,I10349);
DFFARX1 I_6(I1470,I7570,,,I7977,);
DFFARX1 I_7(I7669,I1470,I7570,,,I7541,);
not I_8(I10052,I1477);
and I_9(I10202,I10185,I7541);
nand I_10(I10026,I10219,I10397);
DFFARX1 I_11(I1470,I7570,,,I7532,);
DFFARX1 I_12(I7532,I1470,I10052,,,I10332,);
endmodule


