module test_I6992(I5416,I5334,I3380,I3377,I5105,I3353,I1470,I6992);
input I5416,I5334,I3380,I3377,I5105,I3353,I1470;
output I6992;
wire I5368,I5249,I5097,I5481,I6975,I5204,I5073,I5187,I5625,I5070,I5642,I6924,I5450,I5351;
nor I_0(I5368,I5351,I5204);
not I_1(I5249,I3380);
nand I_2(I5097,I5642,I5368);
DFFARX1 I_3(I5416,I1470,I5105,,,I5481,);
nor I_4(I6975,I6924,I5070);
nand I_5(I5204,I5187,I3353);
DFFARX1 I_6(I5450,I1470,I5105,,,I5073,);
nand I_7(I6992,I6975,I5097);
nor I_8(I5187,I3380);
DFFARX1 I_9(I3377,I1470,I5105,,,I5625,);
and I_10(I5070,I5249,I5481);
not I_11(I5642,I5625);
not I_12(I6924,I5073);
and I_13(I5450,I5416);
DFFARX1 I_14(I5334,I1470,I5105,,,I5351,);
endmodule


