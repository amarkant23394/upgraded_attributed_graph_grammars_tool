module test_final(IN_1_0_l_4,IN_2_0_l_4,IN_4_0_l_4,G18_4_l_4,G15_4_l_4,IN_1_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_7_4_l_4,IN_9_4_l_4,IN_10_4_l_4,blif_clk_net_3_r_0,blif_reset_net_3_r_0,n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0);
input IN_1_0_l_4,IN_2_0_l_4,IN_4_0_l_4,G18_4_l_4,G15_4_l_4,IN_1_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_7_4_l_4,IN_9_4_l_4,IN_10_4_l_4,blif_clk_net_3_r_0,blif_reset_net_3_r_0;
output n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0;
wire ACVQN2_0_r_4,n_266_and_0_0_r_4,ACVQN1_2_r_4,P6_2_r_4,n_429_or_0_3_r_4,G78_3_r_4,n_576_3_r_4,n_102_3_r_4,n_547_3_r_4,n_42_5_r_4,G199_5_r_4,ACVQN2_0_l_4,n_266_and_0_0_l_4,ACVQN1_0_l_4,n4_4_l_4,G42_4_l_4,n_87_4_l_4,n_572_4_l_4,n_573_4_l_4,n_549_4_l_4,n7_4_l_4,n_569_4_l_4,n_452_4_l_4,ACVQN1_0_r_4,P6_internal_2_r_4,n12_3_r_4,n_431_3_r_4,n11_3_r_4,n13_3_r_4,n14_3_r_4,n15_3_r_4,n16_3_r_4,N3_5_r_4,n3_5_r_4,n2_3_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0;
DFFARX1 I_0(n_569_4_l_4,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_r_4,);
and I_1(n_266_and_0_0_r_4,ACVQN2_0_l_4,ACVQN1_0_r_4);
DFFARX1 I_2(n_266_and_0_0_l_4,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_2_r_4,);
not I_3(P6_2_r_4,P6_internal_2_r_4);
nand I_4(n_429_or_0_3_r_4,G42_4_l_4,n12_3_r_4);
DFFARX1 I_5(n_431_3_r_4,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_4,);
nand I_6(n_576_3_r_4,n_573_4_l_4,n11_3_r_4);
not I_7(n_102_3_r_4,n_569_4_l_4);
nand I_8(n_547_3_r_4,ACVQN2_0_l_4,n13_3_r_4);
nor I_9(n_42_5_r_4,G42_4_l_4,n_549_4_l_4);
DFFARX1 I_10(N3_5_r_4,blif_clk_net_3_r_0,n2_3_r_0,G199_5_r_4,);
DFFARX1 I_11(IN_1_0_l_4,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_4,);
and I_12(n_266_and_0_0_l_4,IN_4_0_l_4,ACVQN1_0_l_4);
DFFARX1 I_13(IN_2_0_l_4,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_4,);
nor I_14(n4_4_l_4,G18_4_l_4,IN_1_4_l_4);
DFFARX1 I_15(n4_4_l_4,blif_clk_net_3_r_0,n2_3_r_0,G42_4_l_4,);
not I_16(n_87_4_l_4,G15_4_l_4);
nor I_17(n_572_4_l_4,G15_4_l_4,IN_7_4_l_4);
or I_18(n_573_4_l_4,IN_5_4_l_4,IN_9_4_l_4);
nor I_19(n_549_4_l_4,IN_10_4_l_4,n7_4_l_4);
and I_20(n7_4_l_4,IN_4_4_l_4,n_87_4_l_4);
or I_21(n_569_4_l_4,IN_9_4_l_4,IN_10_4_l_4);
nor I_22(n_452_4_l_4,G18_4_l_4,IN_5_4_l_4);
DFFARX1 I_23(n_549_4_l_4,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_r_4,);
DFFARX1 I_24(ACVQN2_0_l_4,blif_clk_net_3_r_0,n2_3_r_0,P6_internal_2_r_4,);
not I_25(n12_3_r_4,n_266_and_0_0_l_4);
or I_26(n_431_3_r_4,n_572_4_l_4,n14_3_r_4);
nor I_27(n11_3_r_4,n_569_4_l_4,n12_3_r_4);
nor I_28(n13_3_r_4,n_572_4_l_4,n_569_4_l_4);
and I_29(n14_3_r_4,n_452_4_l_4,n15_3_r_4);
nor I_30(n15_3_r_4,n_266_and_0_0_l_4,n16_3_r_4);
not I_31(n16_3_r_4,G42_4_l_4);
and I_32(N3_5_r_4,n_573_4_l_4,n3_5_r_4);
nand I_33(n3_5_r_4,n_549_4_l_4,n_452_4_l_4);
nand I_34(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_35(n_431_3_r_0,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_0,);
nand I_36(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_37(n_102_3_r_0,n_42_5_l_0);
nand I_38(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_39(n4_4_r_0,blif_clk_net_3_r_0,n2_3_r_0,G42_4_r_0,);
nor I_40(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_41(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_42(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_43(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_44(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
not I_45(n2_3_r_0,blif_reset_net_3_r_0);
DFFARX1 I_46(P6_2_r_4,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_0,);
and I_47(n_266_and_0_0_l_0,ACVQN1_0_l_0,n_102_3_r_4);
DFFARX1 I_48(n_266_and_0_0_r_4,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_0,);
and I_49(N1_1_l_0,n3_1_l_0,G78_3_r_4);
DFFARX1 I_50(N1_1_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_1_l_0,);
DFFARX1 I_51(n_547_3_r_4,blif_clk_net_3_r_0,n2_3_r_0,G214_1_l_0,);
nand I_52(n3_1_l_0,n_576_3_r_4,G199_5_r_4);
nor I_53(n_42_5_l_0,ACVQN1_2_r_4,n_42_5_r_4);
and I_54(N3_5_l_0,n3_5_l_0,ACVQN2_0_r_4);
DFFARX1 I_55(N3_5_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_5_l_0,);
nand I_56(n3_5_l_0,ACVQN1_2_r_4,n_429_or_0_3_r_4);
not I_57(n12_3_r_0,G199_1_l_0);
or I_58(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_59(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_60(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_61(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_62(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_63(n16_3_r_0,ACVQN2_0_l_0);
nor I_64(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_65(n_87_4_r_0,G199_5_l_0);
and I_66(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
endmodule


