module test_I9672(I1477,I5743,I8298,I5731,I8250,I5737,I8360,I8445,I1470,I5740,I9672);
input I1477,I5743,I8298,I5731,I8250,I5737,I8360,I8445,I1470,I5740;
output I9672;
wire I8753,I8623,I8190,I8216,I9655,I8377,I8315,I8736,I8462,I8208,I8479,I8267,I8196;
not I_0(I8753,I8736);
DFFARX1 I_1(I5743,I1470,I8216,,,I8623,);
DFFARX1 I_2(I8267,I1470,I8216,,,I8190,);
not I_3(I8216,I1477);
nand I_4(I9655,I8190,I8196);
not I_5(I8377,I8360);
nand I_6(I8315,I8298,I5740);
and I_7(I9672,I9655,I8208);
DFFARX1 I_8(I5731,I1470,I8216,,,I8736,);
DFFARX1 I_9(I8445,I1470,I8216,,,I8462,);
nand I_10(I8208,I8753,I8479);
nor I_11(I8479,I8462,I8315);
nand I_12(I8267,I8250,I5737);
nand I_13(I8196,I8623,I8377);
endmodule


