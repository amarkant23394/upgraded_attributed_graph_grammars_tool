module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_0,blif_reset_net_1_r_0,G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_0,blif_reset_net_1_r_0;
output G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_569_1_r_0,n4_1_l_0,n6_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_0,n6_0,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_0,n6_0,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_0,n6_0,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_0,n6_0,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_0,n6_0,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_0,n6_0,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_0,n6_0,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_0,n6_0,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_0,n6_0,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_0,n6_0,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_0,blif_clk_net_1_r_0,n6_0,G42_1_r_0,);
nor I_32(n_572_1_r_0,n23_0,n_573_1_r_6);
nand I_33(n_573_1_r_0,n21_0,n22_0);
nand I_34(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_35(n_569_1_r_0,n21_0,n26_0);
nor I_36(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_37(N3_2_r_0,blif_clk_net_1_r_0,n6_0,G199_2_r_0,);
DFFARX1 I_38(N1_4_r_0,blif_clk_net_1_r_0,n6_0,G199_4_r_0,);
DFFARX1 I_39(n2_0,blif_clk_net_1_r_0,n6_0,G214_4_r_0,);
nor I_40(n4_1_l_0,G42_1_r_6,n_569_1_r_6);
not I_41(n6_0,blif_reset_net_1_r_0);
DFFARX1 I_42(n4_1_l_0,blif_clk_net_1_r_0,n6_0,n37_0,);
DFFARX1 I_43(n_452_1_r_6,blif_clk_net_1_r_0,n6_0,n38_0,);
not I_44(n20_0,n38_0);
DFFARX1 I_45(G214_4_r_6,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_0,);
nor I_46(n4_1_r_0,n23_0,G42_1_r_6);
nor I_47(N3_2_r_0,n31_0,n32_0);
nor I_48(N1_4_r_0,n29_0,n32_0);
not I_49(n2_0,n31_0);
nor I_50(n21_0,n37_0,n_549_1_r_6);
not I_51(n22_0,n_573_1_r_6);
nand I_52(n23_0,n20_0,n30_0);
nand I_53(n24_0,n38_0,n25_0);
nor I_54(n25_0,n_549_1_r_6,G42_1_r_6);
not I_55(n26_0,G42_1_r_6);
not I_56(n27_0,n29_0);
nor I_57(n28_0,G199_4_r_6,P6_5_r_6);
nand I_58(n29_0,n26_0,n33_0);
not I_59(n30_0,n_549_1_r_6);
nand I_60(n31_0,ACVQN1_3_l_0,n_572_1_r_6);
and I_61(n32_0,n35_0,n36_0);
nand I_62(n33_0,n34_0,ACVQN1_5_r_6);
not I_63(n34_0,G199_4_r_6);
nor I_64(n35_0,G42_1_r_6,G199_4_r_6);
nor I_65(n36_0,n_573_1_r_6,P6_5_r_6);
endmodule


