module test_I5204(I1492,I3504,I2103,I1383,I1832,I1504,I3685,I1470_clk,I1477_rst,I5204);
input I1492,I3504,I2103,I1383,I1832,I1504,I3685,I1470_clk,I1477_rst;
output I5204;
wire I3555,I3353,I1880,I5122,I3380,I3538,I3388_rst,I5187,I1518_rst,I1495,I3620,I3453,I1501,I1486,I1483,I3521,I3846,I3350,I3747,I3637;
DFFARX1 I_0 (I3538,I1470_clk,I3388_rst,I3555);
and I_1(I3353,I3453,I3637);
DFFARX1 I_2 (I1383,I1470_clk,I1518_rst,I1880);
not I_3(I5122,I3350);
nand I_4(I3380,I3521,I3846);
nor I_5(I3538,I1492);
not I_6(I3388_rst,I1477_rst);
nor I_7(I5187,I5122,I3380);
nand I_8(I5204,I5187,I3353);
not I_9(I1518_rst,I1477_rst);
DFFARX1 I_10 (I2103,I1470_clk,I1518_rst,I1495);
nor I_11(I3620,I1492,I1483);
nor I_12(I3453,I1486,I1501);
not I_13(I1501,I1880);
DFFARX1 I_14 (I1832,I1470_clk,I1518_rst,I1486);
DFFARX1 I_15 (I1880,I1470_clk,I1518_rst,I1483);
nor I_16(I3521,I3504,I1495);
nor I_17(I3846,I3747,I3555);
DFFARX1 I_18 (I3685,I1470_clk,I3388_rst,I3350);
DFFARX1 I_19 (I1504,I1470_clk,I3388_rst,I3747);
DFFARX1 I_20 (I3620,I1470_clk,I3388_rst,I3637);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule