module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_2,blif_reset_net_1_r_2,G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_2,blif_reset_net_1_r_2;
output G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n_573_1_r_2,N3_2_l_2,n5_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_2,n5_2,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_2,n5_2,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_2,n5_2,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_2,n5_2,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_2,n5_2,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_2,n5_2,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_2,n5_2,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_2,n5_2,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_2,n5_2,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_2,blif_clk_net_1_r_2,n5_2,G42_1_r_2,);
nor I_34(n_572_1_r_2,n26_2,n18_2);
nand I_35(n_573_1_r_2,n17_2,n19_2);
nor I_36(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_37(n_569_1_r_2,n13_2,n19_2);
not I_38(n_452_1_r_2,n_573_1_r_2);
nor I_39(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_40(N3_2_r_2,blif_clk_net_1_r_2,n5_2,G199_2_r_2,);
DFFARX1 I_41(ACVQN2_3_l_2,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_2,);
not I_42(P6_5_r_2,P6_5_r_internal_2);
and I_43(N3_2_l_2,n24_2,G199_2_r_9);
not I_44(n5_2,blif_reset_net_1_r_2);
DFFARX1 I_45(N3_2_l_2,blif_clk_net_1_r_2,n5_2,G199_2_l_2,);
not I_46(n13_2,G199_2_l_2);
DFFARX1 I_47(G199_4_r_9,blif_clk_net_1_r_2,n5_2,ACVQN2_3_l_2,);
DFFARX1 I_48(n_42_2_r_9,blif_clk_net_1_r_2,n5_2,n16_2,);
and I_49(N1_4_l_2,n25_2,G42_1_r_9);
DFFARX1 I_50(N1_4_l_2,blif_clk_net_1_r_2,n5_2,n26_2,);
DFFARX1 I_51(n_573_1_r_9,blif_clk_net_1_r_2,n5_2,n17_internal_2,);
not I_52(n17_2,n17_internal_2);
nor I_53(n4_1_r_2,n26_2,n22_2);
nor I_54(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_55(G199_2_l_2,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_2,);
nor I_56(n18_2,n_572_1_r_9,n_569_1_r_9);
nand I_57(n19_2,n16_2,G42_1_r_9);
nor I_58(n20_2,n26_2,n21_2);
not I_59(n21_2,n18_2);
and I_60(n22_2,n16_2,G42_1_r_9);
nor I_61(n23_2,n13_2,n21_2);
nand I_62(n24_2,n_569_1_r_9,n_572_1_r_9);
nand I_63(n25_2,n_549_1_r_9,G214_4_r_9);
endmodule


