module test_I2993(I1294,I1954,I1301,I2993);
input I1294,I1954,I1301;
output I2993;
wire I2172,I2733,I2583,I1902,I2203,I2234,I1908,I1937,I2039,I1304,I2945,I2702;
DFFARX1 I_0(I1294,I1937,,,I2172,);
not I_1(I2733,I2702);
not I_2(I2583,I1301);
and I_3(I1902,I2234,I2203);
DFFARX1 I_4(I2172,I1294,I1937,,,I2203,);
nand I_5(I2234,I1954,I1304);
not I_6(I1908,I2039);
not I_7(I1937,I1301);
nor I_8(I2993,I2945,I2733);
DFFARX1 I_9(I1294,I1937,,,I2039,);
DFFARX1 I_10(I1294,,,I1304,);
DFFARX1 I_11(I1902,I1294,I2583,,,I2945,);
not I_12(I2702,I1908);
endmodule


