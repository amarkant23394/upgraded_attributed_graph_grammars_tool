module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_8,n8_8,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_8,n8_8,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_8,n8_8,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_8,n8_8,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_8,n8_8,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_8,n8_8,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_8,n8_8,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_8,n8_8,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_8,n8_8,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_34(n_572_1_r_8,n39_8,n23_8);
and I_35(n_549_1_r_8,n38_8,n23_8);
nand I_36(n_569_1_r_8,n38_8,n24_8);
nor I_37(n_452_1_r_8,n25_8,n26_8);
nor I_38(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_39(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_40(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_41(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_42(n_431_0_l_8,n29_8,G199_4_r_9);
not I_43(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_44(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_45(n19_8,G78_0_l_8);
DFFARX1 I_46(n_572_1_r_9,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_47(n22_8,n39_8);
DFFARX1 I_48(G42_1_r_9,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_49(n4_1_r_8,G78_0_l_8,n33_8);
nor I_50(N3_2_r_8,n22_8,n35_8);
nor I_51(N1_4_r_8,n27_8,n37_8);
nand I_52(n23_8,n32_8,n_569_1_r_9);
not I_53(n24_8,n23_8);
nand I_54(n25_8,n36_8,G42_1_r_9);
nand I_55(n26_8,n27_8,n28_8);
nor I_56(n27_8,n31_8,n_573_1_r_9);
not I_57(n28_8,G199_2_r_9);
and I_58(n29_8,n30_8,G214_4_r_9);
nor I_59(n30_8,n31_8,n_549_1_r_9);
not I_60(n31_8,n_572_1_r_9);
and I_61(n32_8,n28_8,n_573_1_r_9);
nand I_62(n33_8,n28_8,n34_8);
not I_63(n34_8,n25_8);
nor I_64(n35_8,n34_8,G199_2_r_9);
not I_65(n36_8,n_42_2_r_9);
nor I_66(n37_8,n19_8,n38_8);
endmodule


