module test_I8190(I6265,I1477,I4518,I1470,I5881,I8190);
input I6265,I1477,I4518,I1470,I5881;
output I8190;
wire I5737,I8267,I5716,I8216,I6203,I5751,I5963,I5898,I5802,I5719,I8250;
nand I_0(I5737,I6203,I5898);
nand I_1(I8267,I8250,I5737);
and I_2(I5716,I5802,I5963);
not I_3(I8216,I1477);
DFFARX1 I_4(I4518,I1470,I5751,,,I6203,);
not I_5(I5751,I1477);
DFFARX1 I_6(I1470,I5751,,,I5963,);
nor I_7(I5898,I5802,I5881);
DFFARX1 I_8(I1470,I5751,,,I5802,);
DFFARX1 I_9(I6265,I1470,I5751,,,I5719,);
nor I_10(I8250,I5719,I5716);
DFFARX1 I_11(I8267,I1470,I8216,,,I8190,);
endmodule


