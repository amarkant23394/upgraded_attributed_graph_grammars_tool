module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,IN_1_3_l_7,IN_2_3_l_7,IN_3_3_l_7,IN_1_4_l_7,IN_2_4_l_7,IN_3_4_l_7,IN_4_4_l_7,IN_5_4_l_7,blif_clk_net_5_r_5,blif_reset_net_5_r_5,N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,IN_1_3_l_7,IN_2_3_l_7,IN_3_3_l_7,IN_1_4_l_7,IN_2_4_l_7,IN_3_4_l_7,IN_4_4_l_7,IN_5_4_l_7,blif_clk_net_5_r_5,blif_reset_net_5_r_5;
output N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5;
wire N1371_0_r_7,N1508_0_r_7,N6147_2_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,N1507_6_r_7,N1508_6_r_7,n_431_5_r_7,n19_7,n20_7,n21_7,n22_7,n23_7,n24_7,n25_7,n26_7,n27_7,n28_7,n29_7,n30_7,n31_7,n32_7,N1508_0_r_5,N1507_6_r_5,n_431_5_r_5,n6_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5;
nor I_0(N1371_0_r_7,n22_7,n24_7);
nor I_1(N1508_0_r_7,n24_7,n28_7);
nor I_2(N6147_2_r_7,n21_7,n26_7);
nand I_3(n_429_or_0_5_r_7,n19_7,n24_7);
DFFARX1 I_4(n_431_5_r_7,blif_clk_net_5_r_5,n6_5,G78_5_r_7,);
nand I_5(n_576_5_r_7,N1371_0_r_7,n19_7);
not I_6(n_102_5_r_7,n22_7);
nand I_7(n_547_5_r_7,n20_7,n21_7);
nor I_8(N1507_6_r_7,n22_7,n27_7);
nor I_9(N1508_6_r_7,IN_3_1_l_7,n27_7);
nand I_10(n_431_5_r_7,n24_7,n25_7);
nor I_11(n19_7,IN_1_3_l_7,n30_7);
nor I_12(n20_7,n22_7,n23_7);
not I_13(n21_7,n29_7);
nor I_14(n22_7,n29_7,n31_7);
not I_15(n23_7,n27_7);
not I_16(n24_7,N1508_6_r_7);
nand I_17(n25_7,N1507_6_r_7,n19_7);
or I_18(n26_7,n19_7,n23_7);
nand I_19(n27_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_20(n28_7,n19_7,n21_7);
nand I_21(n29_7,IN_1_4_l_7,IN_2_4_l_7);
or I_22(n30_7,IN_2_3_l_7,IN_3_3_l_7);
nor I_23(n31_7,IN_5_4_l_7,n32_7);
and I_24(n32_7,IN_3_4_l_7,IN_4_4_l_7);
nor I_25(N1371_0_r_5,n28_5,n39_5);
not I_26(N1508_0_r_5,n39_5);
nor I_27(N6147_2_r_5,n28_5,n37_5);
nand I_28(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_29(n_431_5_r_5,blif_clk_net_5_r_5,n6_5,G78_5_r_5,);
nand I_30(n_576_5_r_5,n26_5,n27_5);
not I_31(n_102_5_r_5,n28_5);
nand I_32(n_547_5_r_5,n31_5,n32_5);
nor I_33(N1507_6_r_5,n30_5,n32_5);
nor I_34(N1508_6_r_5,n39_5,n41_5);
nand I_35(n_431_5_r_5,n34_5,n35_5);
not I_36(n6_5,blif_reset_net_5_r_5);
nor I_37(n26_5,n29_5,n30_5);
nor I_38(n27_5,n28_5,N6147_2_r_7);
nor I_39(n28_5,n29_5,n44_5);
not I_40(n29_5,n_576_5_r_7);
nand I_41(n30_5,N1508_0_r_5,n43_5);
nor I_42(n31_5,n28_5,n33_5);
nor I_43(n32_5,n40_5,n_102_5_r_7);
nor I_44(n33_5,n29_5,N6147_2_r_7);
or I_45(n34_5,n29_5,N6147_2_r_7);
nand I_46(n35_5,n32_5,n36_5);
not I_47(n36_5,n30_5);
nor I_48(n37_5,N1507_6_r_5,n38_5);
and I_49(n38_5,n39_5,n40_5);
nand I_50(n39_5,n_429_or_0_5_r_7,G78_5_r_7);
nand I_51(n40_5,N1508_0_r_7,n_429_or_0_5_r_7);
nand I_52(n41_5,n28_5,n42_5);
or I_53(n42_5,n32_5,n36_5);
or I_54(n43_5,N6147_2_r_7,N1508_0_r_7);
nor I_55(n44_5,n_547_5_r_7,G78_5_r_7);
endmodule


