module test_I11672(I6896,I1477,I1470,I8930,I11672);
input I6896,I1477,I1470,I8930;
output I11672;
wire I9320,I6884,I6875,I8836,I9303,I9210,I9179,I8862,I11310,I8947;
not I_0(I9320,I9303);
DFFARX1 I_1(I8836,I1470,I11310,,,I11672,);
DFFARX1 I_2(I1470,,,I6884,);
DFFARX1 I_3(I1470,,,I6875,);
nand I_4(I8836,I9320,I9210);
DFFARX1 I_5(I6875,I1470,I8862,,,I9303,);
nor I_6(I9210,I9179,I8947);
DFFARX1 I_7(I6896,I1470,I8862,,,I9179,);
not I_8(I8862,I1477);
not I_9(I11310,I1477);
nand I_10(I8947,I8930,I6884);
endmodule


