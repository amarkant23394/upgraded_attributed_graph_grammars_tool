module test_I16223(I14667,I1477,I14520,I1470,I16223);
input I14667,I1477,I14520,I1470;
output I16223;
wire I14901,I14537,I14808,I14344,I16534,I16240,I14370,I16551,I14335,I14715;
DFFARX1 I_0(I14808,I1470,I14370,,,I14901,);
DFFARX1 I_1(I14520,I1470,I14370,,,I14537,);
DFFARX1 I_2(I1470,I14370,,,I14808,);
nand I_3(I14344,I14537,I14715);
DFFARX1 I_4(I14335,I1470,I16240,,,I16534,);
not I_5(I16240,I1477);
not I_6(I14370,I1477);
not I_7(I16223,I16551);
and I_8(I16551,I16534,I14344);
and I_9(I14335,I14808,I14901);
not I_10(I14715,I14667);
endmodule


