module test_I16789(I1477,I1470,I14954,I15310,I16789);
input I1477,I1470,I14954,I15310;
output I16789;
wire I14933,I17126,I17092,I16818,I14965,I17109;
DFFARX1 I_0(I15310,I1470,I14965,,,I14933,);
not I_1(I16789,I17126);
DFFARX1 I_2(I17109,I1470,I16818,,,I17126,);
DFFARX1 I_3(I14954,I1470,I16818,,,I17092,);
not I_4(I16818,I1477);
not I_5(I14965,I1477);
and I_6(I17109,I17092,I14933);
endmodule


