module test_I1928(I1477,I1215,I1470,I1383,I1928);
input I1477,I1215,I1470,I1383;
output I1928;
wire I1518,I1668,I1637,I1880;
not I_0(I1518,I1477);
not I_1(I1668,I1637);
not I_2(I1637,I1215);
nor I_3(I1928,I1880,I1668);
DFFARX1 I_4(I1383,I1470,I1518,,,I1880,);
endmodule


