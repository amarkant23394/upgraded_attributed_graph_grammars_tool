module test_I2742(I1447,I1391,I1477,I1263,I1470,I2912,I2742);
input I1447,I1391,I1477,I1263,I1470,I2912;
output I2742;
wire I2759,I2946,I2929,I3076,I2963;
not I_0(I2759,I1477);
or I_1(I2742,I3076,I2963);
or I_2(I2946,I2929,I1263);
and I_3(I2929,I2912,I1391);
DFFARX1 I_4(I1447,I1470,I2759,,,I3076,);
DFFARX1 I_5(I2946,I1470,I2759,,,I2963,);
endmodule


