module test_I15016(I10633,I11105,I1477,I1470,I12653,I15016);
input I10633,I11105,I1477,I1470,I12653;
output I15016;
wire I12619,I12670,I12590,I12584,I14999,I12930,I12783,I12752,I12913,I12735,I10647,I12581,I10609;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
not I_2(I12590,I12752);
nand I_3(I15016,I14999,I12581);
and I_4(I12584,I12670,I12783);
nor I_5(I14999,I12584,I12590);
and I_6(I12930,I12913,I10609);
DFFARX1 I_7(I12735,I1470,I12619,,,I12783,);
DFFARX1 I_8(I12735,I1470,I12619,,,I12752,);
DFFARX1 I_9(I10633,I1470,I12619,,,I12913,);
DFFARX1 I_10(I1470,I12619,,,I12735,);
not I_11(I10647,I1477);
DFFARX1 I_12(I12930,I1470,I12619,,,I12581,);
DFFARX1 I_13(I11105,I1470,I10647,,,I10609,);
endmodule


