module test_I9491_rst(I1477_rst,I9491_rst);
,I9491_rst);
input I1477_rst;
output I9491_rst;
wire ;
not I_0(I9491_rst,I1477_rst);
endmodule


