module test_I3512(I3137,I3430,I1294,I1301,I3512);
input I3137,I3430,I1294,I1301;
output I3512;
wire I3464,I3481,I2551,I2575,I2583,I3246,I3447;
or I_0(I3464,I3447,I2575);
DFFARX1 I_1(I3481,I1294,I3246,,,I3512,);
DFFARX1 I_2(I3464,I1294,I3246,,,I3481,);
DFFARX1 I_3(I1294,I2583,,,I2551,);
DFFARX1 I_4(I3137,I1294,I2583,,,I2575,);
not I_5(I2583,I1301);
not I_6(I3246,I1301);
and I_7(I3447,I3430,I2551);
endmodule


