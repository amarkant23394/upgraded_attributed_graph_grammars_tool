module test_I8216(I1477,I8216);
input I1477;
output I8216;
wire ;
not I_0(I8216,I1477);
endmodule


