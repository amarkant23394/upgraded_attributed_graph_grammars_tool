module test_I14359(I1477,I11299,I13296,I1470,I14359);
input I1477,I11299,I13296,I1470;
output I14359;
wire I14667,I13601,I13186,I14650,I13165,I14370,I13197,I13635,I13248,I13159,I13618,I14438,I13189,I11272,I13508,I13491;
and I_0(I14667,I14650,I13189);
DFFARX1 I_1(I11299,I1470,I13197,,,I13601,);
nor I_2(I13186,I13601,I13508);
DFFARX1 I_3(I13165,I1470,I14370,,,I14650,);
DFFARX1 I_4(I13248,I1470,I13197,,,I13165,);
nor I_5(I14359,I14667,I14438);
not I_6(I14370,I1477);
not I_7(I13197,I1477);
and I_8(I13635,I13296,I13618);
DFFARX1 I_9(I1470,I13197,,,I13248,);
DFFARX1 I_10(I13508,I1470,I13197,,,I13159,);
nand I_11(I13618,I13601);
nor I_12(I14438,I13159,I13186);
DFFARX1 I_13(I13635,I1470,I13197,,,I13189,);
DFFARX1 I_14(I1470,,,I11272,);
and I_15(I13508,I13491,I11272);
DFFARX1 I_16(I1470,I13197,,,I13491,);
endmodule


