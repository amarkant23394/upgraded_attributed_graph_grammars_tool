module test_I14370_rst(I1477_rst,I14370_rst);
,I14370_rst);
input I1477_rst;
output I14370_rst;
wire ;
not I_0(I14370_rst,I1477_rst);
endmodule


