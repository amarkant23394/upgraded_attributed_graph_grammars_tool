module test_I9396(I1477,I1470,I7221,I9396);
input I1477,I1470,I7221;
output I9396;
wire I9320,I6875,I9303,I8862,I6907;
not I_0(I9320,I9303);
not I_1(I9396,I9320);
DFFARX1 I_2(I7221,I1470,I6907,,,I6875,);
DFFARX1 I_3(I6875,I1470,I8862,,,I9303,);
not I_4(I8862,I1477);
not I_5(I6907,I1477);
endmodule


