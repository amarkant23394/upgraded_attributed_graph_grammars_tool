module test_I13843(I1477,I10041,I10397,I1470,I11990,I13843);
input I1477,I10041,I10397,I1470,I11990;
output I13843;
wire I12058,I12024,I12380,I10219,I12041,I11965,I10026,I12270,I12287,I12349,I12007,I10044,I12106,I12304,I10020,I11973,I11959;
nand I_0(I12058,I12041,I10026);
nand I_1(I12024,I12007,I10044);
nor I_2(I12380,I12349,I12024);
DFFARX1 I_3(I1470,,,I10219,);
nor I_4(I12041,I11990,I10020);
nor I_5(I13843,I11959,I11965);
DFFARX1 I_6(I12304,I1470,I11973,,,I11965,);
nand I_7(I10026,I10219,I10397);
nand I_8(I12270,I11990);
nand I_9(I12287,I12270,I12024);
DFFARX1 I_10(I10041,I1470,I11973,,,I12349,);
nor I_11(I12007,I10020);
DFFARX1 I_12(I1470,,,I10044,);
not I_13(I12106,I10020);
and I_14(I12304,I12106,I12287);
DFFARX1 I_15(I1470,,,I10020,);
not I_16(I11973,I1477);
nand I_17(I11959,I12058,I12380);
endmodule


