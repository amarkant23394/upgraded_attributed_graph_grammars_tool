module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_9,n5_9,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_9,n5_9,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_9,n5_9,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_9,n5_9,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_9,n5_9,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_9,n5_9,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_9,n5_9,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_32(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_33(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_34(n_549_1_r_9,n17_9,n18_9);
or I_35(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_36(n_452_1_r_9,n26_9,n25_9);
nor I_37(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_38(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_39(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_40(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_41(N3_2_l_9,n22_9,G199_2_r_14);
not I_42(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_43(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_44(n16_9,n27_9);
DFFARX1 I_45(n_572_1_r_14,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_46(n15_9,n26_9);
DFFARX1 I_47(n_573_1_r_14,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_48(n29_9,n29_internal_9);
and I_49(N1_4_l_9,n24_9,n_42_2_r_14);
DFFARX1 I_50(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_51(G42_1_r_14,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_52(n28_9,n28_internal_9);
nor I_53(n4_1_r_9,n27_9,n26_9);
nor I_54(N3_2_r_9,n15_9,n21_9);
nor I_55(N1_4_r_9,n16_9,n21_9);
nor I_56(n_42_2_l_9,G42_1_r_14,n_549_1_r_14);
not I_57(n17_9,n_452_1_r_9);
nand I_58(n18_9,n27_9,n15_9);
nor I_59(n19_9,n29_9,n20_9);
not I_60(n20_9,P6_5_r_14);
and I_61(n21_9,n23_9,P6_5_r_14);
nand I_62(n22_9,G42_1_r_14,ACVQN1_5_r_14);
nor I_63(n23_9,n29_9,n28_9);
nand I_64(n24_9,n_569_1_r_14,n_572_1_r_14);
endmodule


