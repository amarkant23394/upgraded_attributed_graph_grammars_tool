module Benchmark_testing100(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I2615,I2618,I2600,I2609,I2621,I2612,I2603,I2606,I2624);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458;
output I2615,I2618,I2600,I2609,I2621,I2612,I2603,I2606,I2624;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I1496,I3184,I1522,I1539,I1488,I1561,I1578,I3199,I3187,I1595,I3178,I1621,I1629,I3190,I1655,I1663,I3181,I1680,I1467,I3196,I1720,I1728,I1461,I1476,I1773,I3205,I3193,I1790,I3202,I1816,I1464,I1838,I1855,I1872,I1479,I1903,I1920,I1470,I1951,I1473,I1485,I1482,I2037,I2063,I2080,I2029,I2111,I2119,I2136,I2153,I2170,I2187,I2204,I2221,I2026,I2252,I2269,I2286,I2011,I2023,I2331,I2348,I2017,I2379,I2396,I2005,I2427,I2444,I2461,I2487,I2495,I2014,I2526,I2543,I2020,I2574,I2008,I2632,I2658,I2666,I2683,I2700,I2726,I2734,I2760,I2768,I2785,I2802,I2819,I2859,I2867,I2884,I2901,I2918,I2949,I2966,I2992,I3000,I3031,I3062,I3079,I3110,I3213,I3239,I3256,I3264,I3281,I3298,I3315,I3332,I3349,I3380,I3397,I3428,I3445,I3462,I3493,I3533,I3541,I3558,I3575,I3592,I3623,I3640,I3657,I3683,I3705,I3722,I3753,I3798;
not I_0 (I1496,I1458);
DFFARX1 I_1 (I3184,I1451,I1496,I1522,);
DFFARX1 I_2 (I1522,I1451,I1496,I1539,);
not I_3 (I1488,I1539);
not I_4 (I1561,I1522);
nand I_5 (I1578,I3199,I3187);
and I_6 (I1595,I1578,I3178);
DFFARX1 I_7 (I1595,I1451,I1496,I1621,);
not I_8 (I1629,I1621);
DFFARX1 I_9 (I3190,I1451,I1496,I1655,);
and I_10 (I1663,I1655,I3181);
nand I_11 (I1680,I1655,I3181);
nand I_12 (I1467,I1629,I1680);
DFFARX1 I_13 (I3196,I1451,I1496,I1720,);
nor I_14 (I1728,I1720,I1663);
DFFARX1 I_15 (I1728,I1451,I1496,I1461,);
nor I_16 (I1476,I1720,I1621);
nand I_17 (I1773,I3205,I3193);
and I_18 (I1790,I1773,I3202);
DFFARX1 I_19 (I1790,I1451,I1496,I1816,);
nor I_20 (I1464,I1816,I1720);
not I_21 (I1838,I1816);
nor I_22 (I1855,I1838,I1629);
nor I_23 (I1872,I1561,I1855);
DFFARX1 I_24 (I1872,I1451,I1496,I1479,);
nor I_25 (I1903,I1838,I1720);
nor I_26 (I1920,I3178,I3193);
nor I_27 (I1470,I1920,I1903);
not I_28 (I1951,I1920);
nand I_29 (I1473,I1680,I1951);
DFFARX1 I_30 (I1920,I1451,I1496,I1485,);
DFFARX1 I_31 (I1920,I1451,I1496,I1482,);
not I_32 (I2037,I1458);
DFFARX1 I_33 (I1404,I1451,I2037,I2063,);
DFFARX1 I_34 (I2063,I1451,I2037,I2080,);
not I_35 (I2029,I2080);
DFFARX1 I_36 (I1444,I1451,I2037,I2111,);
not I_37 (I2119,I1372);
nor I_38 (I2136,I2063,I2119);
not I_39 (I2153,I1420);
not I_40 (I2170,I1436);
nand I_41 (I2187,I2170,I1420);
nor I_42 (I2204,I2119,I2187);
nor I_43 (I2221,I2111,I2204);
DFFARX1 I_44 (I2170,I1451,I2037,I2026,);
nor I_45 (I2252,I1436,I1412);
nand I_46 (I2269,I2252,I1388);
nor I_47 (I2286,I2269,I2153);
nand I_48 (I2011,I2286,I1372);
DFFARX1 I_49 (I2269,I1451,I2037,I2023,);
nand I_50 (I2331,I2153,I1436);
nor I_51 (I2348,I2153,I1436);
nand I_52 (I2017,I2136,I2348);
not I_53 (I2379,I1428);
nor I_54 (I2396,I2379,I2331);
DFFARX1 I_55 (I2396,I1451,I2037,I2005,);
nor I_56 (I2427,I2379,I1396);
and I_57 (I2444,I2427,I1364);
or I_58 (I2461,I2444,I1380);
DFFARX1 I_59 (I2461,I1451,I2037,I2487,);
nor I_60 (I2495,I2487,I2111);
nor I_61 (I2014,I2063,I2495);
not I_62 (I2526,I2487);
nor I_63 (I2543,I2526,I2221);
DFFARX1 I_64 (I2543,I1451,I2037,I2020,);
nand I_65 (I2574,I2526,I2153);
nor I_66 (I2008,I2379,I2574);
not I_67 (I2632,I1458);
DFFARX1 I_68 (I1470,I1451,I2632,I2658,);
not I_69 (I2666,I2658);
nand I_70 (I2683,I1461,I1479);
and I_71 (I2700,I2683,I1482);
DFFARX1 I_72 (I2700,I1451,I2632,I2726,);
not I_73 (I2734,I1476);
DFFARX1 I_74 (I1464,I1451,I2632,I2760,);
not I_75 (I2768,I2760);
nor I_76 (I2785,I2768,I2666);
and I_77 (I2802,I2785,I1476);
nor I_78 (I2819,I2768,I2734);
nor I_79 (I2615,I2726,I2819);
DFFARX1 I_80 (I1473,I1451,I2632,I2859,);
nor I_81 (I2867,I2859,I2726);
not I_82 (I2884,I2867);
not I_83 (I2901,I2859);
nor I_84 (I2918,I2901,I2802);
DFFARX1 I_85 (I2918,I1451,I2632,I2618,);
nand I_86 (I2949,I1488,I1485);
and I_87 (I2966,I2949,I1467);
DFFARX1 I_88 (I2966,I1451,I2632,I2992,);
nor I_89 (I3000,I2992,I2859);
DFFARX1 I_90 (I3000,I1451,I2632,I2600,);
nand I_91 (I3031,I2992,I2901);
nand I_92 (I2609,I2884,I3031);
not I_93 (I3062,I2992);
nor I_94 (I3079,I3062,I2802);
DFFARX1 I_95 (I3079,I1451,I2632,I2621,);
nor I_96 (I3110,I1461,I1485);
or I_97 (I2612,I2859,I3110);
nor I_98 (I2603,I2992,I3110);
or I_99 (I2606,I2726,I3110);
DFFARX1 I_100 (I3110,I1451,I2632,I2624,);
not I_101 (I3213,I1458);
DFFARX1 I_102 (I2008,I1451,I3213,I3239,);
DFFARX1 I_103 (I2020,I1451,I3213,I3256,);
not I_104 (I3264,I3256);
not I_105 (I3281,I2005);
nor I_106 (I3298,I3281,I2023);
not I_107 (I3315,I2029);
nor I_108 (I3332,I3298,I2011);
nor I_109 (I3349,I3256,I3332);
DFFARX1 I_110 (I3349,I1451,I3213,I3199,);
nor I_111 (I3380,I2011,I2023);
nand I_112 (I3397,I3380,I2005);
DFFARX1 I_113 (I3397,I1451,I3213,I3202,);
nor I_114 (I3428,I3315,I2011);
nand I_115 (I3445,I3428,I2014);
nor I_116 (I3462,I3239,I3445);
DFFARX1 I_117 (I3462,I1451,I3213,I3178,);
not I_118 (I3493,I3445);
nand I_119 (I3190,I3256,I3493);
DFFARX1 I_120 (I3445,I1451,I3213,I3533,);
not I_121 (I3541,I3533);
not I_122 (I3558,I2011);
not I_123 (I3575,I2017);
nor I_124 (I3592,I3575,I2029);
nor I_125 (I3205,I3541,I3592);
nor I_126 (I3623,I3575,I2026);
and I_127 (I3640,I3623,I2005);
or I_128 (I3657,I3640,I2008);
DFFARX1 I_129 (I3657,I1451,I3213,I3683,);
nor I_130 (I3193,I3683,I3239);
not I_131 (I3705,I3683);
and I_132 (I3722,I3705,I3239);
nor I_133 (I3187,I3264,I3722);
nand I_134 (I3753,I3705,I3315);
nor I_135 (I3181,I3575,I3753);
nand I_136 (I3184,I3705,I3493);
nand I_137 (I3798,I3315,I2017);
nor I_138 (I3196,I3558,I3798);
endmodule


