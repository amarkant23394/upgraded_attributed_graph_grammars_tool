module test_I3969(I1477,I2980,I2810,I4017,I1470,I2844,I3969);
input I1477,I2980,I2810,I4017,I1470,I2844;
output I3969;
wire I2733,I3107,I3076,I3983,I3200,I4263,I4051,I3310,I4308,I4034,I2745,I3217,I4325,I3124,I2727,I4246;
nand I_0(I2733,I3217,I3107);
nor I_1(I3107,I3076,I2844);
DFFARX1 I_2(I1470,,,I3076,);
not I_3(I3983,I1477);
DFFARX1 I_4(I1470,,,I3200,);
and I_5(I4263,I4246,I2733);
not I_6(I4051,I4034);
and I_7(I3310,I2844);
DFFARX1 I_8(I2727,I1470,I3983,,,I4308,);
nor I_9(I3969,I4263,I4325);
DFFARX1 I_10(I4017,I1470,I3983,,,I4034,);
nor I_11(I2745,I2980,I3310);
not I_12(I3217,I3200);
and I_13(I4325,I4308,I4051);
nor I_14(I3124,I3076);
nand I_15(I2727,I2810,I3124);
DFFARX1 I_16(I2745,I1470,I3983,,,I4246,);
endmodule


