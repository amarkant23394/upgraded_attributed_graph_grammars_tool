module Benchmark_testing500(I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I982,I989,I2012,I2030,I2033,I2015,I2036,I2021,I2024,I2018,I2027,I2539,I2557,I2560,I2542,I2563,I2548,I2551,I2545,I2554,I5093,I5078,I5072,I5075,I5081,I5090,I5087,I5084,I8453,I8450,I8438,I8444,I8447,I8441,I8456);
input I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I982,I989;
output I2012,I2030,I2033,I2015,I2036,I2021,I2024,I2018,I2027,I2539,I2557,I2560,I2542,I2563,I2548,I2551,I2545,I2554,I5093,I5078,I5072,I5075,I5081,I5090,I5087,I5084,I8453,I8450,I8438,I8444,I8447,I8441,I8456;
wire I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I982,I989,I1024,I1041,I3090,I3069,I1058,I3078,I3087,I1075,I1092,I1109,I1126,I3084,I1143,I3075,I1169,I1177,I1194,I3066,I1211,I1228,I1245,I1004,I1276,I3081,I1293,I3072,I1310,I1013,I1016,I1355,I1007,I1001,I1400,I1417,I995,I998,I1010,I1476,I992,I1534,I1551,I1568,I1585,I1602,I1619,I1636,I1653,I1679,I1687,I1704,I1721,I1738,I1755,I1514,I1786,I1803,I1820,I1523,I1526,I1865,I1517,I1511,I1910,I1927,I1505,I1508,I1520,I1986,I1502,I2044,I2061,I6518,I6506,I2078,I6500,I2095,I2112,I2129,I2146,I6503,I2163,I6509,I2189,I2211,I2228,I2259,I6515,I2276,I2307,I6521,I2324,I2341,I6512,I2372,I2389,I2420,I2451,I2482,I2513,I2571,I2588,I6024,I6027,I2605,I6030,I6039,I2622,I2639,I2656,I2673,I6036,I6042,I2690,I2716,I2738,I2755,I2786,I2803,I2834,I6045,I2851,I2868,I6033,I2899,I2916,I2947,I2978,I3009,I3040,I3098,I3115,I3132,I3149,I3166,I3183,I3200,I3217,I3243,I3265,I3282,I3313,I3330,I3361,I3378,I3395,I3426,I3443,I3474,I3505,I3536,I3567,I3625,I3642,I4120,I4123,I3659,I4126,I4135,I3676,I3693,I3710,I3727,I4132,I4138,I3744,I3770,I3593,I3792,I3809,I3611,I3840,I3857,I3614,I3888,I4141,I3905,I3922,I4129,I3596,I3953,I3970,I3617,I4001,I3602,I4032,I3605,I4063,I3599,I4094,I3608,I4149,I4166,I7027,I7048,I4183,I7033,I4200,I7045,I4217,I7036,I4234,I7030,I4251,I4268,I4285,I4302,I4319,I7039,I7042,I4336,I4353,I4370,I4415,I4446,I4477,I4494,I4525,I4570,I4625,I4642,I4659,I4676,I4693,I4710,I4727,I4744,I4761,I4778,I4795,I4812,I4829,I4846,I4617,I4602,I4891,I4596,I4922,I4599,I4953,I4970,I4605,I5001,I4614,I4611,I5046,I4608,I5101,I5118,I7999,I8002,I5135,I5152,I7996,I8014,I5169,I5186,I8005,I5203,I5220,I5237,I5254,I5271,I8011,I8008,I5288,I5305,I5322,I5367,I5398,I5429,I5446,I5477,I5522,I5577,I5594,I5611,I5628,I5645,I5662,I5679,I5696,I5713,I5730,I5747,I5764,I5781,I5798,I5569,I5554,I5843,I5548,I5874,I5551,I5905,I5922,I5557,I5953,I5566,I5563,I5998,I5560,I6053,I6070,I7557,I7560,I6087,I6104,I7554,I7572,I6121,I6138,I7563,I6155,I6172,I6189,I6206,I6223,I7569,I7566,I6240,I6257,I6274,I6319,I6350,I6381,I6398,I6429,I6474,I6529,I6546,I6563,I6580,I6597,I6614,I6645,I6662,I6679,I6696,I6713,I6730,I6747,I6764,I6781,I6812,I6843,I6874,I6891,I6936,I6967,I6984,I7001,I7056,I7073,I7090,I7107,I7124,I7141,I7172,I7189,I7206,I7223,I7240,I7257,I7274,I7291,I7308,I7339,I7370,I7401,I7418,I7463,I7494,I7511,I7528,I7580,I7597,I7614,I7631,I7648,I7679,I7696,I7713,I7730,I7747,I7764,I7781,I7798,I7857,I7874,I7891,I7922,I7939,I7970,I8022,I8039,I8056,I8073,I8090,I8121,I8138,I8155,I8172,I8189,I8206,I8223,I8240,I8299,I8316,I8333,I8364,I8381,I8412,I8464,I8481,I8498,I8515,I8532,I8563,I8580,I8597,I8614,I8631,I8648,I8665,I8682,I8741,I8758,I8775,I8806,I8823,I8854;
not I_0 (I1024,I989);
or I_1 (I1041,I3090,I3069);
nand I_2 (I1058,I3078,I3087);
not I_3 (I1075,I1058);
nand I_4 (I1092,I1075,I1041);
not I_5 (I1109,I1092);
nand I_6 (I1126,I3084,I3069);
and I_7 (I1143,I1126,I3075);
DFFARX1 I_8 (I1143,I982,I1024,I1169,);
not I_9 (I1177,I1169);
nor I_10 (I1194,I3066,I3069);
nor I_11 (I1211,I1169,I1194);
and I_12 (I1228,I1169,I1194);
nor I_13 (I1245,I1228,I1092);
DFFARX1 I_14 (I1245,I982,I1024,I1004,);
nand I_15 (I1276,I3081,I3066);
nor I_16 (I1293,I1276,I3072);
nand I_17 (I1310,I1109,I1293);
not I_18 (I1013,I1310);
nor I_19 (I1016,I1211,I1310);
nor I_20 (I1355,I1293,I1075);
nor I_21 (I1007,I1177,I1355);
nor I_22 (I1001,I1293,I1194);
not I_23 (I1400,I1276);
nand I_24 (I1417,I1194,I1400);
not I_25 (I995,I1417);
nor I_26 (I998,I1058,I1417);
nor I_27 (I1010,I1400,I1058);
nand I_28 (I1476,I1177,I1276);
nor I_29 (I992,I1075,I1476);
not I_30 (I1534,I989);
or I_31 (I1551,I895,I967);
nand I_32 (I1568,I943,I951);
not I_33 (I1585,I1568);
nand I_34 (I1602,I1585,I1551);
not I_35 (I1619,I1602);
nand I_36 (I1636,I639,I679);
and I_37 (I1653,I1636,I703);
DFFARX1 I_38 (I1653,I982,I1534,I1679,);
not I_39 (I1687,I1679);
nor I_40 (I1704,I935,I679);
nor I_41 (I1721,I1679,I1704);
and I_42 (I1738,I1679,I1704);
nor I_43 (I1755,I1738,I1602);
DFFARX1 I_44 (I1755,I982,I1534,I1514,);
nand I_45 (I1786,I663,I807);
nor I_46 (I1803,I1786,I855);
nand I_47 (I1820,I1619,I1803);
not I_48 (I1523,I1820);
nor I_49 (I1526,I1721,I1820);
nor I_50 (I1865,I1803,I1585);
nor I_51 (I1517,I1687,I1865);
nor I_52 (I1511,I1803,I1704);
not I_53 (I1910,I1786);
nand I_54 (I1927,I1704,I1910);
not I_55 (I1505,I1927);
nor I_56 (I1508,I1568,I1927);
nor I_57 (I1520,I1910,I1568);
nand I_58 (I1986,I1687,I1786);
nor I_59 (I1502,I1585,I1986);
not I_60 (I2044,I989);
or I_61 (I2061,I6518,I6506);
nand I_62 (I2078,I6500,I6500);
not I_63 (I2095,I2078);
nand I_64 (I2112,I2095,I2061);
not I_65 (I2129,I2112);
nand I_66 (I2146,I6503,I6503);
and I_67 (I2163,I2146,I6509);
DFFARX1 I_68 (I2163,I982,I2044,I2189,);
nor I_69 (I2012,I2189,I2078);
nand I_70 (I2211,I2129,I2189);
nor I_71 (I2228,I2189,I2095);
not I_72 (I2030,I2189);
nor I_73 (I2259,I6515,I6503);
not I_74 (I2276,I2259);
nand I_75 (I2033,I2228,I2259);
not I_76 (I2307,I6521);
nor I_77 (I2324,I2189,I6521);
nand I_78 (I2341,I6506,I6512);
nor I_79 (I2015,I2341,I2078);
not I_80 (I2372,I2341);
nor I_81 (I2389,I2259,I2372);
nor I_82 (I2036,I2389,I2112);
nand I_83 (I2420,I2372,I2307);
nand I_84 (I2021,I2129,I2420);
nand I_85 (I2451,I2211,I2420);
DFFARX1 I_86 (I2451,I982,I2044,I2024,);
nand I_87 (I2482,I2276,I2341);
nor I_88 (I2018,I2129,I2482);
nor I_89 (I2513,I2276,I2341);
nand I_90 (I2027,I2513,I2324);
not I_91 (I2571,I989);
or I_92 (I2588,I6024,I6027);
nand I_93 (I2605,I6030,I6039);
not I_94 (I2622,I2605);
nand I_95 (I2639,I2622,I2588);
not I_96 (I2656,I2639);
nand I_97 (I2673,I6036,I6042);
and I_98 (I2690,I2673,I6024);
DFFARX1 I_99 (I2690,I982,I2571,I2716,);
nor I_100 (I2539,I2716,I2605);
nand I_101 (I2738,I2656,I2716);
nor I_102 (I2755,I2716,I2622);
not I_103 (I2557,I2716);
nor I_104 (I2786,I6027,I6042);
not I_105 (I2803,I2786);
nand I_106 (I2560,I2755,I2786);
not I_107 (I2834,I6045);
nor I_108 (I2851,I2716,I6045);
nand I_109 (I2868,I6033,I6030);
nor I_110 (I2542,I2868,I2605);
not I_111 (I2899,I2868);
nor I_112 (I2916,I2786,I2899);
nor I_113 (I2563,I2916,I2639);
nand I_114 (I2947,I2899,I2834);
nand I_115 (I2548,I2656,I2947);
nand I_116 (I2978,I2738,I2947);
DFFARX1 I_117 (I2978,I982,I2571,I2551,);
nand I_118 (I3009,I2803,I2868);
nor I_119 (I2545,I2656,I3009);
nor I_120 (I3040,I2803,I2868);
nand I_121 (I2554,I3040,I2851);
not I_122 (I3098,I989);
or I_123 (I3115,I775,I831);
nand I_124 (I3132,I815,I671);
not I_125 (I3149,I3132);
nand I_126 (I3166,I3149,I3115);
not I_127 (I3183,I3166);
nand I_128 (I3200,I919,I711);
and I_129 (I3217,I3200,I927);
DFFARX1 I_130 (I3217,I982,I3098,I3243,);
nor I_131 (I3066,I3243,I3132);
nand I_132 (I3265,I3183,I3243);
nor I_133 (I3282,I3243,I3149);
not I_134 (I3084,I3243);
nor I_135 (I3313,I887,I711);
not I_136 (I3330,I3313);
nand I_137 (I3087,I3282,I3313);
not I_138 (I3361,I631);
nor I_139 (I3378,I3243,I631);
nand I_140 (I3395,I751,I719);
nor I_141 (I3069,I3395,I3132);
not I_142 (I3426,I3395);
nor I_143 (I3443,I3313,I3426);
nor I_144 (I3090,I3443,I3166);
nand I_145 (I3474,I3426,I3361);
nand I_146 (I3075,I3183,I3474);
nand I_147 (I3505,I3265,I3474);
DFFARX1 I_148 (I3505,I982,I3098,I3078,);
nand I_149 (I3536,I3330,I3395);
nor I_150 (I3072,I3183,I3536);
nor I_151 (I3567,I3330,I3395);
nand I_152 (I3081,I3567,I3378);
not I_153 (I3625,I989);
or I_154 (I3642,I4120,I4123);
nand I_155 (I3659,I4126,I4135);
not I_156 (I3676,I3659);
nand I_157 (I3693,I3676,I3642);
not I_158 (I3710,I3693);
nand I_159 (I3727,I4132,I4138);
and I_160 (I3744,I3727,I4120);
DFFARX1 I_161 (I3744,I982,I3625,I3770,);
nor I_162 (I3593,I3770,I3659);
nand I_163 (I3792,I3710,I3770);
nor I_164 (I3809,I3770,I3676);
not I_165 (I3611,I3770);
nor I_166 (I3840,I4123,I4138);
not I_167 (I3857,I3840);
nand I_168 (I3614,I3809,I3840);
not I_169 (I3888,I4141);
nor I_170 (I3905,I3770,I4141);
nand I_171 (I3922,I4129,I4126);
nor I_172 (I3596,I3922,I3659);
not I_173 (I3953,I3922);
nor I_174 (I3970,I3840,I3953);
nor I_175 (I3617,I3970,I3693);
nand I_176 (I4001,I3953,I3888);
nand I_177 (I3602,I3710,I4001);
nand I_178 (I4032,I3792,I4001);
DFFARX1 I_179 (I4032,I982,I3625,I3605,);
nand I_180 (I4063,I3857,I3922);
nor I_181 (I3599,I3710,I4063);
nor I_182 (I4094,I3857,I3922);
nand I_183 (I3608,I4094,I3905);
not I_184 (I4149,I989);
or I_185 (I4166,I7027,I7048);
nor I_186 (I4183,I4166,I7033);
nor I_187 (I4200,I7027,I7045);
or I_188 (I4217,I4200,I7036);
nor I_189 (I4234,I7030,I7030);
nand I_190 (I4251,I4234,I4217);
not I_191 (I4268,I4251);
nand I_192 (I4285,I4183,I4268);
nor I_193 (I4302,I4183,I4268);
nand I_194 (I4319,I7039,I7042);
nor I_195 (I4336,I4319,I7033);
nor I_196 (I4353,I4319,I4336);
not I_197 (I4370,I4336);
nor I_198 (I4141,I4370,I4285);
or I_199 (I4126,I4183,I4370);
nor I_200 (I4415,I4183,I4336);
nor I_201 (I4120,I4319,I4415);
nor I_202 (I4446,I4353,I4415);
nor I_203 (I4123,I4268,I4446);
nand I_204 (I4477,I4183,I4336);
nand I_205 (I4494,I4251,I4477);
DFFARX1 I_206 (I4494,I982,I4149,I4129,);
not I_207 (I4525,I4319);
nor I_208 (I4138,I4525,I4370);
nand I_209 (I4135,I4302,I4525);
nor I_210 (I4570,I4268,I4319);
nand I_211 (I4132,I4570,I4183);
not I_212 (I4625,I989);
or I_213 (I4642,I1502,I1511);
nor I_214 (I4659,I4642,I1526);
nor I_215 (I4676,I1523,I1505);
or I_216 (I4693,I4676,I1505);
nor I_217 (I4710,I1502,I1508);
nand I_218 (I4727,I4710,I4693);
not I_219 (I4744,I4727);
nand I_220 (I4761,I4659,I4744);
nor I_221 (I4778,I4659,I4744);
nand I_222 (I4795,I1514,I1517);
nor I_223 (I4812,I4795,I1520);
nor I_224 (I4829,I4795,I4812);
not I_225 (I4846,I4812);
nor I_226 (I4617,I4846,I4761);
or I_227 (I4602,I4659,I4846);
nor I_228 (I4891,I4659,I4812);
nor I_229 (I4596,I4795,I4891);
nor I_230 (I4922,I4829,I4891);
nor I_231 (I4599,I4744,I4922);
nand I_232 (I4953,I4659,I4812);
nand I_233 (I4970,I4727,I4953);
DFFARX1 I_234 (I4970,I982,I4625,I4605,);
not I_235 (I5001,I4795);
nor I_236 (I4614,I5001,I4846);
nand I_237 (I4611,I4778,I5001);
nor I_238 (I5046,I4744,I4795);
nand I_239 (I4608,I5046,I4659);
not I_240 (I5101,I989);
or I_241 (I5118,I7999,I8002);
nor I_242 (I5135,I5118,I7999);
nor I_243 (I5152,I7996,I8014);
or I_244 (I5169,I5152,I8002);
nor I_245 (I5186,I8005,I7996);
nand I_246 (I5203,I5186,I5169);
not I_247 (I5220,I5203);
nand I_248 (I5237,I5135,I5220);
nor I_249 (I5254,I5135,I5220);
nand I_250 (I5271,I8011,I8008);
nor I_251 (I5288,I5271,I8005);
nor I_252 (I5305,I5271,I5288);
not I_253 (I5322,I5288);
nor I_254 (I5093,I5322,I5237);
or I_255 (I5078,I5135,I5322);
nor I_256 (I5367,I5135,I5288);
nor I_257 (I5072,I5271,I5367);
nor I_258 (I5398,I5305,I5367);
nor I_259 (I5075,I5220,I5398);
nand I_260 (I5429,I5135,I5288);
nand I_261 (I5446,I5203,I5429);
DFFARX1 I_262 (I5446,I982,I5101,I5081,);
not I_263 (I5477,I5271);
nor I_264 (I5090,I5477,I5322);
nand I_265 (I5087,I5254,I5477);
nor I_266 (I5522,I5220,I5271);
nand I_267 (I5084,I5522,I5135);
not I_268 (I5577,I989);
or I_269 (I5594,I975,I903);
nor I_270 (I5611,I5594,I727);
nor I_271 (I5628,I911,I783);
or I_272 (I5645,I5628,I871);
nor I_273 (I5662,I687,I863);
nand I_274 (I5679,I5662,I5645);
not I_275 (I5696,I5679);
nand I_276 (I5713,I5611,I5696);
nor I_277 (I5730,I5611,I5696);
nand I_278 (I5747,I655,I647);
nor I_279 (I5764,I5747,I959);
nor I_280 (I5781,I5747,I5764);
not I_281 (I5798,I5764);
nor I_282 (I5569,I5798,I5713);
or I_283 (I5554,I5611,I5798);
nor I_284 (I5843,I5611,I5764);
nor I_285 (I5548,I5747,I5843);
nor I_286 (I5874,I5781,I5843);
nor I_287 (I5551,I5696,I5874);
nand I_288 (I5905,I5611,I5764);
nand I_289 (I5922,I5679,I5905);
DFFARX1 I_290 (I5922,I982,I5577,I5557,);
not I_291 (I5953,I5747);
nor I_292 (I5566,I5953,I5798);
nand I_293 (I5563,I5730,I5953);
nor I_294 (I5998,I5696,I5747);
nand I_295 (I5560,I5998,I5611);
not I_296 (I6053,I989);
or I_297 (I6070,I7557,I7560);
nor I_298 (I6087,I6070,I7557);
nor I_299 (I6104,I7554,I7572);
or I_300 (I6121,I6104,I7560);
nor I_301 (I6138,I7563,I7554);
nand I_302 (I6155,I6138,I6121);
not I_303 (I6172,I6155);
nand I_304 (I6189,I6087,I6172);
nor I_305 (I6206,I6087,I6172);
nand I_306 (I6223,I7569,I7566);
nor I_307 (I6240,I6223,I7563);
nor I_308 (I6257,I6223,I6240);
not I_309 (I6274,I6240);
nor I_310 (I6045,I6274,I6189);
or I_311 (I6030,I6087,I6274);
nor I_312 (I6319,I6087,I6240);
nor I_313 (I6024,I6223,I6319);
nor I_314 (I6350,I6257,I6319);
nor I_315 (I6027,I6172,I6350);
nand I_316 (I6381,I6087,I6240);
nand I_317 (I6398,I6155,I6381);
DFFARX1 I_318 (I6398,I982,I6053,I6033,);
not I_319 (I6429,I6223);
nor I_320 (I6042,I6429,I6274);
nand I_321 (I6039,I6206,I6429);
nor I_322 (I6474,I6172,I6223);
nand I_323 (I6036,I6474,I6087);
not I_324 (I6529,I989);
nor I_325 (I6546,I995,I992);
not I_326 (I6563,I1010);
not I_327 (I6580,I1001);
nor I_328 (I6597,I6580,I6546);
nand I_329 (I6614,I6597,I1010);
not I_330 (I6503,I6614);
nor I_331 (I6645,I6580,I6563);
and I_332 (I6662,I6614,I1016);
nor I_333 (I6679,I6645,I1016);
nand I_334 (I6696,I1013,I1004);
not I_335 (I6713,I6696);
nand I_336 (I6730,I6713,I6679);
nor I_337 (I6747,I992,I995);
not I_338 (I6764,I1007);
nor I_339 (I6781,I6764,I998);
nor I_340 (I6500,I6781,I6614);
not I_341 (I6812,I6781);
or I_342 (I6515,I6730,I6781);
nor I_343 (I6843,I6781,I6696);
nand I_344 (I6512,I6645,I6843);
nor I_345 (I6874,I6747,I6764);
nand I_346 (I6891,I6713,I6874);
not I_347 (I6518,I6891);
nor I_348 (I6521,I6662,I6891);
or I_349 (I6936,I6781,I6874);
nor I_350 (I6506,I6713,I6936);
nor I_351 (I6967,I6874,I1016);
nand I_352 (I6984,I6967,I6713);
nand I_353 (I7001,I6812,I6984);
DFFARX1 I_354 (I7001,I982,I6529,I6509,);
not I_355 (I7056,I989);
nor I_356 (I7073,I879,I839);
not I_357 (I7090,I759);
not I_358 (I7107,I743);
nor I_359 (I7124,I7107,I7073);
nand I_360 (I7141,I7124,I759);
not I_361 (I7030,I7141);
nor I_362 (I7172,I7107,I7090);
and I_363 (I7189,I7141,I823);
nor I_364 (I7206,I7172,I823);
nand I_365 (I7223,I791,I767);
not I_366 (I7240,I7223);
nand I_367 (I7257,I7240,I7206);
nor I_368 (I7274,I847,I695);
not I_369 (I7291,I735);
nor I_370 (I7308,I7291,I799);
nor I_371 (I7027,I7308,I7141);
not I_372 (I7339,I7308);
or I_373 (I7042,I7257,I7308);
nor I_374 (I7370,I7308,I7223);
nand I_375 (I7039,I7172,I7370);
nor I_376 (I7401,I7274,I7291);
nand I_377 (I7418,I7240,I7401);
not I_378 (I7045,I7418);
nor I_379 (I7048,I7189,I7418);
or I_380 (I7463,I7308,I7401);
nor I_381 (I7033,I7240,I7463);
nor I_382 (I7494,I7401,I823);
nand I_383 (I7511,I7494,I7240);
nand I_384 (I7528,I7339,I7511);
DFFARX1 I_385 (I7528,I982,I7056,I7036,);
not I_386 (I7580,I989);
and I_387 (I7597,I5560,I5566);
nor I_388 (I7614,I7597,I5554);
nand I_389 (I7631,I5551,I5548);
nor I_390 (I7648,I7631,I7614);
not I_391 (I7569,I7648);
not I_392 (I7679,I7631);
or I_393 (I7696,I5557,I5569);
nor I_394 (I7713,I7696,I5551);
nor I_395 (I7730,I7713,I7679);
nand I_396 (I7747,I5548,I5563);
nor I_397 (I7764,I7747,I5554);
not I_398 (I7781,I7764);
nor I_399 (I7798,I7648,I7781);
nand I_400 (I7566,I7798,I7713);
nor I_401 (I7554,I7781,I7730);
nand I_402 (I7560,I7713,I7781);
nor I_403 (I7857,I7648,I7747);
nand I_404 (I7874,I7857,I7713);
nand I_405 (I7891,I7781,I7874);
DFFARX1 I_406 (I7891,I982,I7580,I7563,);
not I_407 (I7922,I7747);
or I_408 (I7939,I7713,I7922);
nor I_409 (I7557,I7679,I7939);
nor I_410 (I7970,I7648,I7922);
nand I_411 (I7572,I7970,I7679);
not I_412 (I8022,I989);
and I_413 (I8039,I4608,I4614);
nor I_414 (I8056,I8039,I4602);
nand I_415 (I8073,I4599,I4596);
nor I_416 (I8090,I8073,I8056);
not I_417 (I8011,I8090);
not I_418 (I8121,I8073);
or I_419 (I8138,I4605,I4617);
nor I_420 (I8155,I8138,I4599);
nor I_421 (I8172,I8155,I8121);
nand I_422 (I8189,I4596,I4611);
nor I_423 (I8206,I8189,I4602);
not I_424 (I8223,I8206);
nor I_425 (I8240,I8090,I8223);
nand I_426 (I8008,I8240,I8155);
nor I_427 (I7996,I8223,I8172);
nand I_428 (I8002,I8155,I8223);
nor I_429 (I8299,I8090,I8189);
nand I_430 (I8316,I8299,I8155);
nand I_431 (I8333,I8223,I8316);
DFFARX1 I_432 (I8333,I982,I8022,I8005,);
not I_433 (I8364,I8189);
or I_434 (I8381,I8155,I8364);
nor I_435 (I7999,I8121,I8381);
nor I_436 (I8412,I8090,I8364);
nand I_437 (I8014,I8412,I8121);
not I_438 (I8464,I989);
and I_439 (I8481,I3593,I3593);
nor I_440 (I8498,I8481,I3617);
nand I_441 (I8515,I3614,I3602);
nor I_442 (I8532,I8515,I8498);
not I_443 (I8453,I8532);
not I_444 (I8563,I8515);
or I_445 (I8580,I3596,I3596);
nor I_446 (I8597,I8580,I3599);
nor I_447 (I8614,I8597,I8563);
nand I_448 (I8631,I3608,I3611);
nor I_449 (I8648,I8631,I3605);
not I_450 (I8665,I8648);
nor I_451 (I8682,I8532,I8665);
nand I_452 (I8450,I8682,I8597);
nor I_453 (I8438,I8665,I8614);
nand I_454 (I8444,I8597,I8665);
nor I_455 (I8741,I8532,I8631);
nand I_456 (I8758,I8741,I8597);
nand I_457 (I8775,I8665,I8758);
DFFARX1 I_458 (I8775,I982,I8464,I8447,);
not I_459 (I8806,I8631);
or I_460 (I8823,I8597,I8806);
nor I_461 (I8441,I8563,I8823);
nor I_462 (I8854,I8532,I8806);
nand I_463 (I8456,I8854,I8563);
endmodule


