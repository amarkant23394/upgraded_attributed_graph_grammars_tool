module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_5,blif_reset_net_7_r_5,N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_5,blif_reset_net_7_r_5;
output N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,n_549_7_r_5,n4_7_r_5,n7_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_7_r_5,n7_5,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_7_r_5,n7_5,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
nor I_40(N1371_0_r_5,n28_5,n46_5);
nand I_41(N1508_0_r_5,n26_5,n43_5);
not I_42(N1372_1_r_5,n43_5);
nor I_43(N1508_1_r_5,n30_5,n43_5);
nor I_44(N6147_2_r_5,n29_5,n32_5);
nor I_45(N1507_6_r_5,n26_5,n44_5);
nor I_46(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_47(n4_7_r_5,blif_clk_net_7_r_5,n7_5,G42_7_r_5,);
and I_48(n_572_7_r_5,n27_5,n28_5);
nand I_49(n_573_7_r_5,n26_5,n27_5);
nand I_50(n_549_7_r_5,n_42_8_r_8,G199_8_r_8);
nand I_51(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_52(n_452_7_r_5,n29_5);
nor I_53(n4_7_r_5,n30_5,n31_5);
not I_54(n7_5,blif_reset_net_7_r_5);
not I_55(n26_5,n35_5);
nand I_56(n27_5,n40_5,n41_5);
nand I_57(n28_5,N6134_9_r_8,G199_8_r_8);
nand I_58(n29_5,n27_5,n33_5);
nor I_59(n30_5,n45_5,N1508_6_r_8);
not I_60(n31_5,n_549_7_r_5);
nor I_61(n32_5,n34_5,n35_5);
not I_62(n33_5,n30_5);
nor I_63(n34_5,n31_5,n36_5);
nor I_64(n35_5,n28_5,n_42_8_r_8);
not I_65(n36_5,n28_5);
nand I_66(n37_5,n36_5,n38_5);
nand I_67(n38_5,n26_5,n39_5);
nand I_68(n39_5,n30_5,n31_5);
nor I_69(n40_5,N1508_1_r_8,N1508_10_r_8);
or I_70(n41_5,n42_5,N1507_6_r_8);
nor I_71(n42_5,N6147_9_r_8,N1371_0_r_8);
nand I_72(n43_5,n36_5,n46_5);
nor I_73(n44_5,n_549_7_r_5,n33_5);
or I_74(n45_5,N1371_0_r_8,N1508_6_r_8);
and I_75(n46_5,n31_5,n47_5);
or I_76(n47_5,N1507_6_r_8,N1508_1_r_8);
endmodule


