module test_I13197(I1477,I13197);
input I1477;
output I13197;
wire ;
not I_0(I13197,I1477);
endmodule


