module test_I1971(I1410,I1492,I1543,I1294,I1207,I1301,I1971);
input I1410,I1492,I1543,I1294,I1207,I1301;
output I1971;
wire I1444,I1319,I1560,I1622,I1749,I1342,I1427,I1509,I1639,I1310,I1577;
nand I_0(I1444,I1427,I1410);
DFFARX1 I_1(I1749,I1294,I1342,,,I1319,);
and I_2(I1560,I1410,I1543);
DFFARX1 I_3(I1294,I1342,,,I1622,);
or I_4(I1749,I1639,I1560);
nor I_5(I1971,I1310,I1319);
not I_6(I1342,I1301);
DFFARX1 I_7(I1294,I1342,,,I1427,);
DFFARX1 I_8(I1492,I1294,I1342,,,I1509,);
and I_9(I1639,I1622,I1207);
DFFARX1 I_10(I1577,I1294,I1342,,,I1310,);
and I_11(I1577,I1509,I1444);
endmodule


