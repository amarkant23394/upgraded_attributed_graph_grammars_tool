module test_I14332(I13697,I13180,I1477,I13168,I1470,I14332);
input I13697,I13180,I1477,I13168,I1470;
output I14332;
wire I13197,I14503,I14520,I13174,I14537,I14370;
not I_0(I13197,I1477);
nand I_1(I14503,I13180,I13168);
and I_2(I14520,I14503,I13174);
DFFARX1 I_3(I13697,I1470,I13197,,,I13174,);
DFFARX1 I_4(I14520,I1470,I14370,,,I14537,);
not I_5(I14370,I1477);
DFFARX1 I_6(I14537,I1470,I14370,,,I14332,);
endmodule


