module test_I15603(I1477,I14066,I1470,I15603);
input I1477,I14066,I1470;
output I15603;
wire I14083,I13752,I13746,I16052,I13775,I15611,I14278,I15928,I16069;
DFFARX1 I_0(I14066,I1470,I13775,,,I14083,);
DFFARX1 I_1(I14278,I1470,I13775,,,I13752,);
not I_2(I13746,I14083);
nor I_3(I15603,I15928,I16069);
DFFARX1 I_4(I13752,I1470,I15611,,,I16052,);
not I_5(I13775,I1477);
not I_6(I15611,I1477);
or I_7(I14278,I14066);
DFFARX1 I_8(I13746,I1470,I15611,,,I15928,);
not I_9(I16069,I16052);
endmodule


