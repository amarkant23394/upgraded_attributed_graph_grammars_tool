module test_final(G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_14,blif_reset_net_1_r_14,G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14);
input G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_14,blif_reset_net_1_r_14;
output G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14;
wire G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12,n_431_0_l_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n_452_1_r_14,n4_1_l_14,n3_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14;
DFFARX1 I_0(n4_1_r_12,blif_clk_net_1_r_14,n3_14,G42_1_r_12,);
nor I_1(n_572_1_r_12,n29_12,n30_12);
nand I_2(n_573_1_r_12,n26_12,n27_12);
nor I_3(n_549_1_r_12,n33_12,n34_12);
and I_4(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_5(N3_2_r_12,blif_clk_net_1_r_14,n3_14,G199_2_r_12,);
DFFARX1 I_6(n3_12,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_12,);
not I_7(P6_5_r_12,P6_5_r_internal_12);
or I_8(n_431_0_l_12,IN_8_0_l_12,n36_12);
DFFARX1 I_9(n_431_0_l_12,blif_clk_net_1_r_14,n3_14,n41_12,);
DFFARX1 I_10(IN_2_5_l_12,blif_clk_net_1_r_14,n3_14,ACVQN1_5_l_12,);
not I_11(n22_12,ACVQN1_5_l_12);
DFFARX1 I_12(IN_1_5_l_12,blif_clk_net_1_r_14,n3_14,n42_12,);
nor I_13(n4_1_r_12,n41_12,n31_12);
nor I_14(N3_2_r_12,n22_12,n40_12);
not I_15(n3_12,n39_12);
DFFARX1 I_16(ACVQN1_5_l_12,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_12,);
and I_17(n26_12,IN_5_0_l_12,IN_7_0_l_12);
nor I_18(n27_12,n28_12,n29_12);
not I_19(n28_12,IN_11_0_l_12);
nand I_20(n29_12,n31_12,n32_12);
nand I_21(n30_12,IN_11_0_l_12,n42_12);
not I_22(n31_12,G2_0_l_12);
not I_23(n32_12,IN_10_0_l_12);
nand I_24(n33_12,n31_12,n35_12);
nand I_25(n34_12,IN_5_0_l_12,IN_7_0_l_12);
nand I_26(n35_12,n41_12,n42_12);
and I_27(n36_12,IN_2_0_l_12,n37_12);
nor I_28(n37_12,IN_4_0_l_12,n38_12);
not I_29(n38_12,G1_0_l_12);
nor I_30(n39_12,IN_5_0_l_12,n38_12);
nor I_31(n40_12,G2_0_l_12,n39_12);
DFFARX1 I_32(n_452_1_r_14,blif_clk_net_1_r_14,n3_14,G42_1_r_14,);
and I_33(n_572_1_r_14,n18_14,n19_14);
nand I_34(n_573_1_r_14,n16_14,n17_14);
nor I_35(n_549_1_r_14,n20_14,n21_14);
or I_36(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_37(n_452_1_r_14,n23_14,n_42_2_r_12);
nor I_38(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_39(N3_2_r_14,blif_clk_net_1_r_14,n3_14,G199_2_r_14,);
DFFARX1 I_40(n_572_1_l_14,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_14,);
not I_41(P6_5_r_14,P6_5_r_internal_14);
nor I_42(n4_1_l_14,n_572_1_r_12,n_573_1_r_12);
not I_43(n3_14,blif_reset_net_1_r_14);
DFFARX1 I_44(n4_1_l_14,blif_clk_net_1_r_14,n3_14,n15_internal_14,);
not I_45(n15_14,n15_internal_14);
DFFARX1 I_46(G42_1_r_12,blif_clk_net_1_r_14,n3_14,ACVQN2_3_l_14,);
DFFARX1 I_47(ACVQN1_5_r_12,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_14,);
and I_48(N3_2_r_14,n26_14,n27_14);
nor I_49(n_572_1_l_14,n_572_1_r_12,P6_5_r_12);
DFFARX1 I_50(ACVQN2_3_l_14,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_14,);
nor I_51(n16_14,G42_1_r_12,n_42_2_r_12);
not I_52(n17_14,n_572_1_l_14);
nor I_53(n18_14,G42_1_r_12,n_549_1_r_12);
nand I_54(n19_14,ACVQN1_3_l_14,n_573_1_r_12);
nor I_55(n20_14,n_549_1_r_12,n_573_1_r_12);
nor I_56(n21_14,n15_14,n22_14);
nand I_57(n22_14,n24_14,n25_14);
nand I_58(n23_14,n15_14,n24_14);
not I_59(n24_14,G42_1_r_12);
not I_60(n25_14,n_549_1_r_12);
nor I_61(n26_14,n20_14,n_42_2_r_12);
nand I_62(n27_14,n28_14,G199_2_r_12);
not I_63(n28_14,n_572_1_r_12);
endmodule


