module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_5_r_15,n9_15,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
and I_42(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_43(N1508_0_r_15,n55_15,N1508_6_r_11);
nor I_44(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_45(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_46(N1372_4_r_15,n39_15);
nor I_47(N1508_4_r_15,n39_15,n43_15);
nand I_48(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_49(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_50(n_576_5_r_15,n31_15,n32_15);
not I_51(n_102_5_r_15,n33_15);
nand I_52(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_53(N1507_6_r_15,n42_15,n46_15);
nand I_54(N1508_6_r_15,n39_15,n40_15);
nand I_55(n_431_5_r_15,n36_15,n37_15);
not I_56(n9_15,blif_reset_net_5_r_15);
nor I_57(n31_15,n33_15,n34_15);
nor I_58(n32_15,n44_15,N1372_1_r_11);
nor I_59(n33_15,n54_15,n55_15);
nand I_60(n34_15,n49_15,n_429_or_0_5_r_11);
nand I_61(n35_15,N1508_1_r_11,N1507_6_r_11);
not I_62(n36_15,n32_15);
nand I_63(n37_15,n34_15,n38_15);
not I_64(n38_15,n46_15);
nand I_65(n39_15,n38_15,n41_15);
nand I_66(n40_15,n41_15,n42_15);
and I_67(n41_15,n51_15,N1372_1_r_11);
and I_68(n42_15,n47_15,N1507_6_r_11);
and I_69(n43_15,n34_15,n36_15);
or I_70(n44_15,N6147_2_r_11,N6147_3_r_11);
not I_71(n45_15,N1372_1_r_15);
nand I_72(n46_15,n53_15,N1507_6_r_11);
nor I_73(n47_15,n34_15,n48_15);
not I_74(n48_15,N1508_1_r_11);
and I_75(n49_15,n50_15,N1508_10_r_11);
nand I_76(n50_15,n51_15,n52_15);
nand I_77(n51_15,N6147_3_r_11,n_576_5_r_11);
not I_78(n52_15,N1372_1_r_11);
nor I_79(n53_15,n48_15,N6147_2_r_11);
nor I_80(n54_15,G78_5_r_11,n_547_5_r_11);
not I_81(n55_15,N1508_1_r_11);
endmodule


