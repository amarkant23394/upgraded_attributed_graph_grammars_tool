module test_I2005_rst(I1301_rst,I2005_rst);
,I2005_rst);
input I1301_rst;
output I2005_rst;
wire ;
not I_0(I2005_rst,I1301_rst);
endmodule


