module test_I5512(I1477,I1470,I1501,I1897,I5512);
input I1477,I1470,I1501,I1897;
output I5512;
wire I3388,I1486,I3368,I3470,I1504,I3453,I3747,I5105,I1767;
not I_0(I3388,I1477);
DFFARX1 I_1(I1470,,,I1486,);
nand I_2(I3368,I3747,I3470);
not I_3(I3470,I3453);
nand I_4(I1504,I1767,I1897);
nor I_5(I3453,I1486,I1501);
DFFARX1 I_6(I3368,I1470,I5105,,,I5512,);
DFFARX1 I_7(I1504,I1470,I3388,,,I3747,);
not I_8(I5105,I1477);
DFFARX1 I_9(I1470,,,I1767,);
endmodule


