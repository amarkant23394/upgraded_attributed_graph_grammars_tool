module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_17,n6_17,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_17,n6_17,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_17,n6_17,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_17,n6_17,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_17,n6_17,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_17,n6_17,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_17,n6_17,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_32(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_33(n_573_1_r_17,n20_17,n21_17);
nand I_34(n_549_1_r_17,n23_17,n24_17);
nand I_35(n_569_1_r_17,n21_17,n22_17);
not I_36(n_452_1_r_17,n23_17);
DFFARX1 I_37(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_38(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_39(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_40(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_41(n_431_0_l_17,n26_17,G199_2_r_14);
not I_42(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_43(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_44(n20_17,n20_internal_17);
DFFARX1 I_45(n_569_1_r_14,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_46(n_549_1_r_14,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_47(n19_17,n19_internal_17);
nor I_48(n4_1_r_17,n5_17,n25_17);
not I_49(n2_17,n29_17);
DFFARX1 I_50(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_51(n17_17,n17_internal_17);
nor I_52(N1_4_r_17,n29_17,n31_17);
not I_53(n5_17,G42_1_r_14);
and I_54(n21_17,n32_17,n_572_1_r_14);
not I_55(n22_17,n25_17);
nand I_56(n23_17,n20_17,n22_17);
nand I_57(n24_17,n19_17,n22_17);
nand I_58(n25_17,n30_17,ACVQN1_5_r_14);
and I_59(n26_17,n27_17,n_42_2_r_14);
nor I_60(n27_17,n28_17,n_573_1_r_14);
not I_61(n28_17,G42_1_r_14);
nor I_62(n29_17,n28_17,P6_5_r_14);
and I_63(n30_17,n5_17,P6_5_r_14);
nor I_64(n31_17,n21_17,G42_1_r_14);
nor I_65(n32_17,G42_1_r_14,n_572_1_r_14);
endmodule


