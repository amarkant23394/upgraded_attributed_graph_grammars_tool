module test_I9456(I8202,I8181,I8753,I1477,I1470,I9909,I9456);
input I8202,I8181,I8753,I1477,I1470,I9909;
output I9456;
wire I9926,I8187,I9576,I8216,I9754,I9689,I9771,I9960,I8178,I9943,I9491;
nor I_0(I9926,I9689,I9909);
DFFARX1 I_1(I1470,I8216,,,I8187,);
nor I_2(I9576,I8181,I8202);
not I_3(I8216,I1477);
DFFARX1 I_4(I8187,I1470,I9491,,,I9754,);
DFFARX1 I_5(I1470,I9491,,,I9689,);
and I_6(I9771,I9754,I8178);
or I_7(I9960,I9771,I9943);
DFFARX1 I_8(I8753,I1470,I8216,,,I8178,);
and I_9(I9943,I9576,I9926);
DFFARX1 I_10(I9960,I1470,I9491,,,I9456,);
not I_11(I9491,I1477);
endmodule


