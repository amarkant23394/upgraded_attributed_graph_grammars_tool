module test_I2505(I1223,I1207,I1294,I1239,I1301,I2505);
input I1223,I1207,I1294,I1239,I1301;
output I2505;
wire I1410,I1328,I1622,I2313,I1937,I1331,I2389,I1639,I2406,I2488;
nor I_0(I1410,I1223,I1239);
nand I_1(I1328,I1639);
DFFARX1 I_2(I1294,,,I1622,);
DFFARX1 I_3(I1331,I1294,I1937,,,I2313,);
not I_4(I1937,I1301);
nor I_5(I2505,I2313,I2488);
nor I_6(I1331,I1639,I1410);
DFFARX1 I_7(I1328,I1294,I1937,,,I2389,);
and I_8(I1639,I1622,I1207);
not I_9(I2406,I2389);
not I_10(I2488,I2406);
endmodule


