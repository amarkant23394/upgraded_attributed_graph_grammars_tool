module test_I9413(I7238,I1477,I7427,I1470,I7286,I9413);
input I7238,I1477,I7427,I1470,I7286;
output I9413;
wire I9320,I9396,I6884,I6893,I6875,I7156,I9303,I8930,I6907,I8879,I8862,I6887,I7492,I8947;
not I_0(I9320,I9303);
not I_1(I9396,I9320);
DFFARX1 I_2(I7492,I1470,I6907,,,I6884,);
nand I_3(I6893,I7156,I7286);
DFFARX1 I_4(I1470,I6907,,,I6875,);
DFFARX1 I_5(I1470,I6907,,,I7156,);
DFFARX1 I_6(I6875,I1470,I8862,,,I9303,);
nor I_7(I8930,I8879,I6893);
not I_8(I6907,I1477);
not I_9(I8879,I6887);
not I_10(I8862,I1477);
nand I_11(I6887,I7427);
or I_12(I7492,I7427,I7238);
and I_13(I9413,I8947,I9396);
nand I_14(I8947,I8930,I6884);
endmodule


