module test_I7559(I6843,I6329,I1470,I6363,I7559);
input I6843,I6329,I1470,I6363;
output I7559;
wire I6297,I7652,I7587,I6380,I6318,I6300,I7669;
DFFARX1 I_0(I6843,I1470,I6329,,,I6297,);
nor I_1(I7652,I7587,I6297);
not I_2(I7559,I7669);
not I_3(I7587,I6300);
DFFARX1 I_4(I6363,I1470,I6329,,,I6380,);
not I_5(I6318,I6380);
DFFARX1 I_6(I1470,I6329,,,I6300,);
nand I_7(I7669,I7652,I6318);
endmodule


