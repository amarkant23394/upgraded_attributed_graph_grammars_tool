module test_I12191(I7556,I1477,I8124,I1470,I12191);
input I7556,I1477,I8124,I1470;
output I12191;
wire I12140,I10583,I7570,I10014,I10023,I10052,I10137,I7553,I12157,I10490,I10017,I12174,I10035;
not I_0(I12140,I10014);
DFFARX1 I_1(I10490,I1470,I10052,,,I10583,);
not I_2(I7570,I1477);
DFFARX1 I_3(I1470,I10052,,,I10014,);
DFFARX1 I_4(I10137,I1470,I10052,,,I10023,);
not I_5(I10052,I1477);
DFFARX1 I_6(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_7(I8124,I1470,I7570,,,I7553,);
nor I_8(I12157,I12140,I10035);
DFFARX1 I_9(I7556,I1470,I10052,,,I10490,);
and I_10(I10017,I10490,I10583);
and I_11(I12174,I12157,I10017);
or I_12(I12191,I12174,I10023);
not I_13(I10035,I10490);
endmodule


