module test_final(IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_1_8_l_0,IN_2_8_l_0,IN_3_8_l_0,IN_6_8_l_0,IN_1_10_l_0,IN_2_10_l_0,IN_3_10_l_0,IN_4_10_l_0,blif_clk_net_8_r_1,blif_reset_net_8_r_1,N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1);
input IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_1_8_l_0,IN_2_8_l_0,IN_3_8_l_0,IN_6_8_l_0,IN_1_10_l_0,IN_2_10_l_0,IN_3_10_l_0,IN_4_10_l_0,blif_clk_net_8_r_1,blif_reset_net_8_r_1;
output N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1;
wire N1371_0_r_0,N1508_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0,N3_8_l_0,n40_0,n4_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,I_BUFF_1_9_r_1,N3_8_l_1,n7_1,n38_1,n22_1,N3_8_r_1,n23_1,n24_1,n25_1,n26_1,n27_1,n28_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1;
nor I_0(N1371_0_r_0,n24_0,n25_0);
not I_1(N1508_0_r_0,n25_0);
nor I_2(N6147_2_r_0,n28_0,n29_0);
nand I_3(n_429_or_0_5_r_0,n4_0,n25_0);
DFFARX1 I_4(n4_0,blif_clk_net_8_r_1,n7_1,G78_5_r_0,);
nand I_5(n_576_5_r_0,n23_0,n24_0);
not I_6(n_102_5_r_0,n40_0);
nand I_7(n_547_5_r_0,n26_0,n27_0);
nor I_8(N1507_6_r_0,n_102_5_r_0,n37_0);
nor I_9(N1508_6_r_0,n25_0,n33_0);
and I_10(N3_8_l_0,IN_6_8_l_0,n32_0);
DFFARX1 I_11(N3_8_l_0,blif_clk_net_8_r_1,n7_1,n40_0,);
not I_12(n4_0,n31_0);
nor I_13(n23_0,n40_0,n25_0);
and I_14(n24_0,n4_0,n39_0);
nand I_15(n25_0,IN_1_1_l_0,IN_2_1_l_0);
nor I_16(n26_0,n40_0,n24_0);
nor I_17(n27_0,IN_1_8_l_0,IN_3_8_l_0);
nor I_18(n28_0,IN_3_1_l_0,n25_0);
nand I_19(n29_0,n_102_5_r_0,n30_0);
nand I_20(n30_0,n27_0,n31_0);
nand I_21(n31_0,IN_1_10_l_0,IN_2_10_l_0);
nand I_22(n32_0,IN_2_8_l_0,IN_3_8_l_0);
nand I_23(n33_0,n34_0,n35_0);
nand I_24(n34_0,n_102_5_r_0,n36_0);
not I_25(n35_0,IN_3_1_l_0);
not I_26(n36_0,n27_0);
nor I_27(n37_0,n36_0,n38_0);
nand I_28(n38_0,N1508_0_r_0,n35_0);
or I_29(n39_0,IN_3_10_l_0,IN_4_10_l_0);
nor I_30(N6147_3_r_1,n26_1,n27_1);
not I_31(N1372_4_r_1,n34_1);
nor I_32(N1508_4_r_1,n30_1,n34_1);
nor I_33(n_42_8_r_1,n23_1,n24_1);
DFFARX1 I_34(N3_8_r_1,blif_clk_net_8_r_1,n7_1,G199_8_r_1,);
nor I_35(N6147_9_r_1,n22_1,n25_1);
nor I_36(N6134_9_r_1,n29_1,n30_1);
not I_37(I_BUFF_1_9_r_1,n32_1);
not I_38(N1372_10_r_1,n36_1);
nor I_39(N1508_10_r_1,n35_1,n36_1);
and I_40(N3_8_l_1,n33_1,G78_5_r_0);
not I_41(n7_1,blif_reset_net_8_r_1);
DFFARX1 I_42(N3_8_l_1,blif_clk_net_8_r_1,n7_1,n38_1,);
not I_43(n22_1,n38_1);
nor I_44(N3_8_r_1,n31_1,n32_1);
nor I_45(n23_1,n28_1,N1507_6_r_0);
nor I_46(n24_1,N1508_6_r_0,G78_5_r_0);
nor I_47(n25_1,n23_1,n26_1);
not I_48(n26_1,n30_1);
nand I_49(n27_1,n22_1,n28_1);
nand I_50(n28_1,n_576_5_r_0,n_429_or_0_5_r_0);
not I_51(n29_1,n28_1);
nand I_52(n30_1,N6147_2_r_0,n_429_or_0_5_r_0);
and I_53(n31_1,n38_1,n24_1);
nand I_54(n32_1,n26_1,n37_1);
nand I_55(n33_1,n_547_5_r_0,N1508_6_r_0);
nand I_56(n34_1,n24_1,n29_1);
nor I_57(n35_1,n38_1,n24_1);
nand I_58(n36_1,I_BUFF_1_9_r_1,n23_1);
or I_59(n37_1,N1371_0_r_0,N6147_2_r_0);
endmodule


