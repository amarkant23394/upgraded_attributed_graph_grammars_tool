module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_15,n4_15,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_15,n4_15,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_15,n4_15,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_15,n4_15,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_15,n4_15,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_15,n4_15,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_15,n4_15,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_15,n4_15,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_15,n4_15,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_34(n_572_1_r_15,n17_15,n19_15);
nand I_35(n_573_1_r_15,n15_15,n18_15);
nor I_36(n_549_1_r_15,n21_15,n22_15);
nand I_37(n_569_1_r_15,n15_15,n20_15);
nor I_38(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_39(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_40(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_41(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_42(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_43(n4_1_l_15,n_569_1_r_9,G214_4_r_9);
not I_44(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_45(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_46(n15_15,G42_1_l_15);
DFFARX1 I_47(n_42_2_r_9,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_48(n17_15,n17_internal_15);
DFFARX1 I_49(G42_1_r_9,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_50(n_572_1_l_15,n_573_1_r_9,G199_4_r_9);
DFFARX1 I_51(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_52(n14_15,n14_internal_15);
nand I_53(N1_4_r_15,n25_15,n26_15);
or I_54(n_573_1_l_15,n_549_1_r_9,G199_2_r_9);
nor I_55(n18_15,n_549_1_r_9,G42_1_r_9);
nand I_56(n19_15,n27_15,n28_15);
nand I_57(n20_15,n30_15,n_572_1_r_9);
not I_58(n21_15,n20_15);
and I_59(n22_15,n17_15,n_572_1_l_15);
nor I_60(n23_15,n_569_1_r_9,G199_2_r_9);
or I_61(n24_15,n_549_1_r_9,G42_1_r_9);
or I_62(n25_15,n_573_1_l_15,n_569_1_r_9);
nand I_63(n26_15,n19_15,n23_15);
not I_64(n27_15,G42_1_r_9);
nand I_65(n28_15,n29_15,n_572_1_r_9);
not I_66(n29_15,G199_4_r_9);
endmodule


