module test_I1328(I1231,I1255,I1215,I1359,I1294,I1207,I1301,I1328);
input I1231,I1255,I1215,I1359,I1294,I1207,I1301;
output I1328;
wire I1622,I1376,I1342,I1393,I1828,I1639,I1780;
nand I_0(I1328,I1639,I1828);
DFFARX1 I_1(I1255,I1294,I1342,,,I1622,);
and I_2(I1376,I1359,I1231);
not I_3(I1342,I1301);
DFFARX1 I_4(I1376,I1294,I1342,,,I1393,);
nor I_5(I1828,I1780,I1393);
and I_6(I1639,I1622,I1207);
DFFARX1 I_7(I1215,I1294,I1342,,,I1780,);
endmodule


