module test_I1784(I1716,I1423,I1215,I1279,I1439,I1535,I1470_clk,I1477_rst,I1784);
input I1716,I1423,I1215,I1279,I1439,I1535,I1470_clk,I1477_rst;
output I1784;
wire I1733,I1767,I1620,I1603,I1750,I1586,I1518_rst;
and I_0(I1733,I1716,I1439);
nor I_1(I1784,I1767,I1620);
DFFARX1 I_2 (I1750,I1470_clk,I1518_rst,I1767);
not I_3(I1620,I1603);
nand I_4(I1603,I1586,I1423);
or I_5(I1750,I1733,I1279);
nor I_6(I1586,I1535,I1215);
not I_7(I1518_rst,I1477_rst);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule