module test_I2158(I1477,I1470,I2198,I1271,I2158);
input I1477,I1470,I2198,I1271;
output I2158;
wire I2181,I2232,I2263,I2215;
not I_0(I2181,I1477);
DFFARX1 I_1(I2215,I1470,I2181,,,I2232,);
DFFARX1 I_2(I2232,I1470,I2181,,,I2263,);
not I_3(I2158,I2263);
and I_4(I2215,I2198,I1271);
endmodule


