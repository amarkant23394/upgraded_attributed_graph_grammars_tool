module test_final(G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7,n_431_0_l_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_7,blif_clk_net_1_r_17,n6_17,G42_1_r_7,);
nor I_1(n_572_1_r_7,n30_7,n31_7);
nand I_2(n_573_1_r_7,IN_7_0_l_7,n28_7);
nor I_3(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_4(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_5(N1_4_r_7,blif_clk_net_1_r_17,n6_17,G199_4_r_7,);
DFFARX1 I_6(n26_7,blif_clk_net_1_r_17,n6_17,G214_4_r_7,);
DFFARX1 I_7(n5_7,blif_clk_net_1_r_17,n6_17,ACVQN1_5_r_7,);
not I_8(P6_5_r_7,P6_5_r_internal_7);
or I_9(n_431_0_l_7,IN_8_0_l_7,n36_7);
DFFARX1 I_10(n_431_0_l_7,blif_clk_net_1_r_17,n6_17,n43_7,);
not I_11(n27_7,n43_7);
DFFARX1 I_12(IN_2_5_l_7,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_7,);
DFFARX1 I_13(IN_1_5_l_7,blif_clk_net_1_r_17,n6_17,n44_7,);
nor I_14(n4_1_r_7,n30_7,n38_7);
nor I_15(N1_4_r_7,n27_7,n40_7);
nand I_16(n26_7,IN_11_0_l_7,n39_7);
not I_17(n5_7,G2_0_l_7);
DFFARX1 I_18(ACVQN1_5_l_7,blif_clk_net_1_r_17,n6_17,P6_5_r_internal_7,);
nor I_19(n28_7,n26_7,n29_7);
not I_20(n29_7,IN_5_0_l_7);
not I_21(n30_7,G1_0_l_7);
nand I_22(n31_7,n27_7,n29_7);
nor I_23(n32_7,ACVQN1_5_l_7,n34_7);
nor I_24(n33_7,G2_0_l_7,n29_7);
not I_25(n34_7,IN_7_0_l_7);
nor I_26(n35_7,n43_7,n44_7);
and I_27(n36_7,IN_2_0_l_7,n37_7);
nor I_28(n37_7,IN_4_0_l_7,n30_7);
nand I_29(n38_7,G2_0_l_7,n29_7);
nor I_30(n39_7,G2_0_l_7,IN_10_0_l_7);
nor I_31(n40_7,n44_7,n41_7);
nor I_32(n41_7,n34_7,n42_7);
nand I_33(n42_7,IN_5_0_l_7,n5_7);
DFFARX1 I_34(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_35(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_36(n_573_1_r_17,n20_17,n21_17);
nand I_37(n_549_1_r_17,n23_17,n24_17);
nand I_38(n_569_1_r_17,n21_17,n22_17);
not I_39(n_452_1_r_17,n23_17);
DFFARX1 I_40(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_41(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_42(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_43(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_44(n_431_0_l_17,n26_17,G42_1_r_7);
not I_45(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_46(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_47(n20_17,n20_internal_17);
DFFARX1 I_48(G214_4_r_7,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_49(n_549_1_r_7,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_50(n19_17,n19_internal_17);
nor I_51(n4_1_r_17,n5_17,n25_17);
not I_52(n2_17,n29_17);
DFFARX1 I_53(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_54(n17_17,n17_internal_17);
nor I_55(N1_4_r_17,n29_17,n31_17);
not I_56(n5_17,G199_4_r_7);
and I_57(n21_17,n32_17,P6_5_r_7);
not I_58(n22_17,n25_17);
nand I_59(n23_17,n20_17,n22_17);
nand I_60(n24_17,n19_17,n22_17);
nand I_61(n25_17,n30_17,n_572_1_r_7);
and I_62(n26_17,n27_17,n_572_1_r_7);
nor I_63(n27_17,n28_17,n_573_1_r_7);
not I_64(n28_17,G42_1_r_7);
nor I_65(n29_17,n28_17,n_569_1_r_7);
and I_66(n30_17,n5_17,n_569_1_r_7);
nor I_67(n31_17,n21_17,G199_4_r_7);
nor I_68(n32_17,G199_4_r_7,ACVQN1_5_r_7);
endmodule


