module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_5_r_13,n9_13,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_5_r_13,n9_13,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N1371_0_r_13,n59_13,n61_13);
nor I_41(N1508_0_r_13,n59_13,n60_13);
not I_42(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_43(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_44(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_45(n_102_5_r_13,N1372_1_r_16,n_452_7_r_16);
nand I_46(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_47(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_48(n_572_7_r_13,n40_13,n41_13);
nand I_49(n_573_7_r_13,n37_13,n38_13);
nor I_50(n_549_7_r_13,n46_13,n47_13);
nand I_51(n_569_7_r_13,n37_13,n43_13);
nand I_52(n_452_7_r_13,n52_13,n53_13);
nor I_53(n4_7_l_13,N1508_1_r_16,N6147_2_r_16);
not I_54(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_55(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_56(n33_13,n62_13);
nand I_57(n_431_5_r_13,n54_13,n55_13);
not I_58(n1_13,n52_13);
nor I_59(n34_13,n35_13,n36_13);
nor I_60(n35_13,n42_13,N1508_6_r_16);
nand I_61(n36_13,n50_13,n58_13);
nand I_62(n37_13,n44_13,n45_13);
or I_63(n38_13,n39_13,N1372_1_r_16);
nand I_64(n39_13,N1371_0_r_16,N1508_0_r_16);
not I_65(n40_13,n36_13);
nor I_66(n41_13,n35_13,n_452_7_r_16);
not I_67(n42_13,N1507_6_r_16);
or I_68(n43_13,n_572_7_r_16,N1508_1_r_16);
not I_69(n44_13,N1508_6_r_16);
not I_70(n45_13,N1508_0_r_16);
nor I_71(n46_13,n39_13,n40_13);
nor I_72(n47_13,n_572_7_r_16,N1508_1_r_16);
nor I_73(n48_13,n50_13,n51_13);
nor I_74(n49_13,N1508_0_r_16,N1508_6_r_16);
not I_75(n50_13,n59_13);
not I_76(n51_13,n_102_5_r_13);
nand I_77(n52_13,n33_13,n39_13);
nand I_78(n53_13,n33_13,N1372_1_r_16);
nor I_79(n54_13,N1372_1_r_16,n_572_7_r_16);
nand I_80(n55_13,n62_13,n56_13);
nor I_81(n56_13,n39_13,n57_13);
not I_82(n57_13,N1508_1_r_16);
or I_83(n58_13,N6147_2_r_16,n_569_7_r_16);
nand I_84(n59_13,G42_7_r_16,n_573_7_r_16);
nor I_85(n60_13,n51_13,n_572_7_r_16);
nor I_86(n61_13,n39_13,N1372_1_r_16);
endmodule


