module test_final(G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7,n_431_0_l_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_7,blif_clk_net_1_r_15,n4_15,G42_1_r_7,);
nor I_1(n_572_1_r_7,n30_7,n31_7);
nand I_2(n_573_1_r_7,IN_7_0_l_7,n28_7);
nor I_3(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_4(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_5(N1_4_r_7,blif_clk_net_1_r_15,n4_15,G199_4_r_7,);
DFFARX1 I_6(n26_7,blif_clk_net_1_r_15,n4_15,G214_4_r_7,);
DFFARX1 I_7(n5_7,blif_clk_net_1_r_15,n4_15,ACVQN1_5_r_7,);
not I_8(P6_5_r_7,P6_5_r_internal_7);
or I_9(n_431_0_l_7,IN_8_0_l_7,n36_7);
DFFARX1 I_10(n_431_0_l_7,blif_clk_net_1_r_15,n4_15,n43_7,);
not I_11(n27_7,n43_7);
DFFARX1 I_12(IN_2_5_l_7,blif_clk_net_1_r_15,n4_15,ACVQN1_5_l_7,);
DFFARX1 I_13(IN_1_5_l_7,blif_clk_net_1_r_15,n4_15,n44_7,);
nor I_14(n4_1_r_7,n30_7,n38_7);
nor I_15(N1_4_r_7,n27_7,n40_7);
nand I_16(n26_7,IN_11_0_l_7,n39_7);
not I_17(n5_7,G2_0_l_7);
DFFARX1 I_18(ACVQN1_5_l_7,blif_clk_net_1_r_15,n4_15,P6_5_r_internal_7,);
nor I_19(n28_7,n26_7,n29_7);
not I_20(n29_7,IN_5_0_l_7);
not I_21(n30_7,G1_0_l_7);
nand I_22(n31_7,n27_7,n29_7);
nor I_23(n32_7,ACVQN1_5_l_7,n34_7);
nor I_24(n33_7,G2_0_l_7,n29_7);
not I_25(n34_7,IN_7_0_l_7);
nor I_26(n35_7,n43_7,n44_7);
and I_27(n36_7,IN_2_0_l_7,n37_7);
nor I_28(n37_7,IN_4_0_l_7,n30_7);
nand I_29(n38_7,G2_0_l_7,n29_7);
nor I_30(n39_7,G2_0_l_7,IN_10_0_l_7);
nor I_31(n40_7,n44_7,n41_7);
nor I_32(n41_7,n34_7,n42_7);
nand I_33(n42_7,IN_5_0_l_7,n5_7);
DFFARX1 I_34(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_35(n_572_1_r_15,n17_15,n19_15);
nand I_36(n_573_1_r_15,n15_15,n18_15);
nor I_37(n_549_1_r_15,n21_15,n22_15);
nand I_38(n_569_1_r_15,n15_15,n20_15);
nor I_39(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_40(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_41(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_42(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_43(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_44(n4_1_l_15,n_549_1_r_7,G42_1_r_7);
not I_45(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_46(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_47(n15_15,G42_1_l_15);
DFFARX1 I_48(n_572_1_r_7,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_49(n17_15,n17_internal_15);
DFFARX1 I_50(G42_1_r_7,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_51(n_572_1_l_15,n_573_1_r_7,P6_5_r_7);
DFFARX1 I_52(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_53(n14_15,n14_internal_15);
nand I_54(N1_4_r_15,n25_15,n26_15);
or I_55(n_573_1_l_15,G199_4_r_7,ACVQN1_5_r_7);
nor I_56(n18_15,n_572_1_r_7,G199_4_r_7);
nand I_57(n19_15,n27_15,n28_15);
nand I_58(n20_15,n30_15,G214_4_r_7);
not I_59(n21_15,n20_15);
and I_60(n22_15,n17_15,n_572_1_l_15);
nor I_61(n23_15,ACVQN1_5_r_7,G42_1_r_7);
or I_62(n24_15,n_572_1_r_7,G199_4_r_7);
or I_63(n25_15,n_573_1_l_15,G42_1_r_7);
nand I_64(n26_15,n19_15,n23_15);
not I_65(n27_15,n_572_1_r_7);
nand I_66(n28_15,n29_15,n_569_1_r_7);
not I_67(n29_15,n_573_1_r_7);
endmodule


