module test_I6363(I2733,I1477,I2748,I2742,I2730,I4147,I1470,I6363);
input I2733,I1477,I2748,I2742,I2730,I4147,I1470;
output I6363;
wire I3983,I3954,I6346,I4164,I4068,I4263,I2724,I4000,I4308,I3969,I4034,I3963,I4325,I4017,I4181,I4051,I4246;
not I_0(I3983,I1477);
not I_1(I3954,I4068);
nand I_2(I6346,I3969,I3954);
and I_3(I6363,I6346,I3963);
and I_4(I4164,I4147,I2748);
nor I_5(I4068,I2742,I2724);
and I_6(I4263,I4246,I2733);
DFFARX1 I_7(I1470,,,I2724,);
nand I_8(I4000,I2724);
DFFARX1 I_9(I1470,I3983,,,I4308,);
nor I_10(I3969,I4263,I4325);
DFFARX1 I_11(I4017,I1470,I3983,,,I4034,);
nor I_12(I3963,I4181,I4034);
and I_13(I4325,I4308,I4051);
and I_14(I4017,I4000,I2730);
DFFARX1 I_15(I4164,I1470,I3983,,,I4181,);
not I_16(I4051,I4034);
DFFARX1 I_17(I1470,I3983,,,I4246,);
endmodule


