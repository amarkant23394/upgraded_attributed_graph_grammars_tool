module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_1,n5_1,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_1,n5_1,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_1,n5_1,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_1,n5_1,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_1,n5_1,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_1,n5_1,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_1,n5_1,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_1,n5_1,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_1,n5_1,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_34(n_572_1_r_1,n26_1,n19_1);
nand I_35(n_573_1_r_1,n16_1,n18_1);
nor I_36(n_549_1_r_1,n20_1,n21_1);
nor I_37(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_38(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_39(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_40(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_41(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_42(N3_2_l_1,n23_1,n_569_1_r_9);
not I_43(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_44(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_45(n17_1,n26_1);
DFFARX1 I_46(n_572_1_r_9,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_47(n16_1,n16_internal_1);
DFFARX1 I_48(n_549_1_r_9,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_49(N1_4_l_1,n25_1,n_573_1_r_9);
DFFARX1 I_50(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_51(n_573_1_r_9,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_52(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_53(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_54(n14_1,n14_internal_1);
nor I_55(N1_4_r_1,n17_1,n24_1);
nand I_56(n18_1,ACVQN1_3_l_1,n_42_2_r_9);
nor I_57(n19_1,G42_1_r_9,n_572_1_r_9);
not I_58(n20_1,n18_1);
nor I_59(n21_1,n26_1,n22_1);
not I_60(n22_1,n19_1);
nand I_61(n23_1,G42_1_r_9,G199_2_r_9);
nor I_62(n24_1,n18_1,n22_1);
nand I_63(n25_1,G199_4_r_9,G214_4_r_9);
endmodule


