module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_5_r_15,n9_15,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
and I_35(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_36(N1508_0_r_15,n55_15,N1508_6_r_4);
nor I_37(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_38(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_39(N1372_4_r_15,n39_15);
nor I_40(N1508_4_r_15,n39_15,n43_15);
nand I_41(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_42(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_43(n_576_5_r_15,n31_15,n32_15);
not I_44(n_102_5_r_15,n33_15);
nand I_45(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_46(N1507_6_r_15,n42_15,n46_15);
nand I_47(N1508_6_r_15,n39_15,n40_15);
nand I_48(n_431_5_r_15,n36_15,n37_15);
not I_49(n9_15,blif_reset_net_5_r_15);
nor I_50(n31_15,n33_15,n34_15);
nor I_51(n32_15,n44_15,N1508_6_r_4);
nor I_52(n33_15,n54_15,n55_15);
nand I_53(n34_15,n49_15,n_549_7_r_4);
nand I_54(n35_15,G42_7_r_4,N6134_9_r_4);
not I_55(n36_15,n32_15);
nand I_56(n37_15,n34_15,n38_15);
not I_57(n38_15,n46_15);
nand I_58(n39_15,n38_15,n41_15);
nand I_59(n40_15,n41_15,n42_15);
and I_60(n41_15,n51_15,n_572_7_r_4);
and I_61(n42_15,n47_15,G42_7_r_4);
and I_62(n43_15,n34_15,n36_15);
or I_63(n44_15,n_569_7_r_4,N1371_0_r_4);
not I_64(n45_15,N1372_1_r_15);
nand I_65(n46_15,n53_15,G42_7_r_4);
nor I_66(n47_15,n34_15,n48_15);
not I_67(n48_15,N6134_9_r_4);
and I_68(n49_15,n50_15,G42_7_r_4);
nand I_69(n50_15,n51_15,n52_15);
nand I_70(n51_15,N1371_0_r_4,n_452_7_r_4);
not I_71(n52_15,n_572_7_r_4);
nor I_72(n53_15,n48_15,n_572_7_r_4);
nor I_73(n54_15,N1507_6_r_4,n_549_7_r_4);
not I_74(n55_15,N1507_6_r_4);
endmodule


