module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_5,blif_reset_net_7_r_5,N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_5,blif_reset_net_7_r_5;
output N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,n_549_7_r_5,n4_7_r_5,n7_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_7_r_5,n7_5,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
nor I_34(N1371_0_r_5,n28_5,n46_5);
nand I_35(N1508_0_r_5,n26_5,n43_5);
not I_36(N1372_1_r_5,n43_5);
nor I_37(N1508_1_r_5,n30_5,n43_5);
nor I_38(N6147_2_r_5,n29_5,n32_5);
nor I_39(N1507_6_r_5,n26_5,n44_5);
nor I_40(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_41(n4_7_r_5,blif_clk_net_7_r_5,n7_5,G42_7_r_5,);
and I_42(n_572_7_r_5,n27_5,n28_5);
nand I_43(n_573_7_r_5,n26_5,n27_5);
nand I_44(n_549_7_r_5,N1508_0_r_12,N1508_6_r_12);
nand I_45(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_46(n_452_7_r_5,n29_5);
nor I_47(n4_7_r_5,n30_5,n31_5);
not I_48(n7_5,blif_reset_net_7_r_5);
not I_49(n26_5,n35_5);
nand I_50(n27_5,n40_5,n41_5);
nand I_51(n28_5,N6147_9_r_12,N1507_6_r_12);
nand I_52(n29_5,n27_5,n33_5);
nor I_53(n30_5,n45_5,n_572_7_r_12);
not I_54(n31_5,n_549_7_r_5);
nor I_55(n32_5,n34_5,n35_5);
not I_56(n33_5,n30_5);
nor I_57(n34_5,n31_5,n36_5);
nor I_58(n35_5,n28_5,G42_7_r_12);
not I_59(n36_5,n28_5);
nand I_60(n37_5,n36_5,n38_5);
nand I_61(n38_5,n26_5,n39_5);
nand I_62(n39_5,n30_5,n31_5);
nor I_63(n40_5,N1371_0_r_12,n_549_7_r_12);
or I_64(n41_5,n42_5,n_572_7_r_12);
nor I_65(n42_5,N1507_6_r_12,G42_7_r_12);
nand I_66(n43_5,n36_5,n46_5);
nor I_67(n44_5,n_549_7_r_5,n33_5);
or I_68(n45_5,N1508_6_r_12,N1508_0_r_12);
and I_69(n46_5,n31_5,n47_5);
or I_70(n47_5,n_569_7_r_12,N1371_0_r_12);
endmodule


