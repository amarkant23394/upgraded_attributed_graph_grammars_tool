module test_I8947(I1477,I7221,I7139,I6992,I1470,I8947);
input I1477,I7221,I7139,I6992,I1470;
output I8947;
wire I7173,I6893,I7317,I6907,I6887,I7238,I8930,I7410,I7269,I7492,I6884,I7286,I7156,I7427,I8879;
nor I_0(I7173,I7156);
nand I_1(I6893,I7156,I7286);
nor I_2(I7317,I7269);
not I_3(I6907,I1477);
nand I_4(I6887,I7427,I7317);
and I_5(I7238,I7221,I7173);
nor I_6(I8930,I8879,I6893);
DFFARX1 I_7(I1470,I6907,,,I7410,);
DFFARX1 I_8(I1470,I6907,,,I7269,);
or I_9(I7492,I7427,I7238);
DFFARX1 I_10(I7492,I1470,I6907,,,I6884,);
nor I_11(I7286,I7269,I6992);
nand I_12(I8947,I8930,I6884);
DFFARX1 I_13(I7139,I1470,I6907,,,I7156,);
not I_14(I7427,I7410);
not I_15(I8879,I6887);
endmodule


