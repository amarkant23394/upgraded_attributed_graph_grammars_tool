module test_I12380(I1477,I7535,I7550,I1470,I10287,I12380);
input I1477,I7535,I7550,I1470,I10287;
output I12380;
wire I10507,I12024,I10120,I7538,I10029,I10041,I10490,I10052,I10366,I10349,I12349,I12007,I10044,I10332,I10459,I10020,I11973;
and I_0(I10507,I10490,I10366);
nand I_1(I12024,I12007,I10044);
nor I_2(I12380,I12349,I12024);
nor I_3(I10120,I7538,I7535);
DFFARX1 I_4(I1470,,,I7538,);
DFFARX1 I_5(I10459,I1470,I10052,,,I10029,);
nor I_6(I10041,I10349,I10120);
DFFARX1 I_7(I1470,I10052,,,I10490,);
not I_8(I10052,I1477);
nand I_9(I10366,I10349);
and I_10(I10349,I10332,I7550);
DFFARX1 I_11(I10041,I1470,I11973,,,I12349,);
nor I_12(I12007,I10020,I10029);
DFFARX1 I_13(I10507,I1470,I10052,,,I10044,);
DFFARX1 I_14(I1470,I10052,,,I10332,);
or I_15(I10459,I10349);
DFFARX1 I_16(I10287,I1470,I10052,,,I10020,);
not I_17(I11973,I1477);
endmodule


