module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14,I_BUFF_1_9_r_14,N3_8_l_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_14,n47_14,n30_14);
nor I_1(N1508_0_r_14,n30_14,n41_14);
nor I_2(N1507_6_r_14,n37_14,n44_14);
nor I_3(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_4(n4_7_r_14,blif_clk_net_7_r_3,n10_3,G42_7_r_14,);
nor I_5(n_572_7_r_14,n28_14,n29_14);
nand I_6(n_573_7_r_14,n26_14,n27_14);
nor I_7(n_549_7_r_14,n31_14,n32_14);
nand I_8(n_569_7_r_14,n26_14,n30_14);
nor I_9(n_452_7_r_14,n47_14,n28_14);
nor I_10(N6147_9_r_14,n36_14,n37_14);
nor I_11(N6134_9_r_14,n28_14,n36_14);
not I_12(I_BUFF_1_9_r_14,n26_14);
and I_13(N3_8_l_14,IN_6_8_l_14,n38_14);
DFFARX1 I_14(N3_8_l_14,blif_clk_net_7_r_3,n10_3,n47_14,);
nor I_15(n4_7_r_14,n47_14,n35_14);
nand I_16(n26_14,IN_1_10_l_14,IN_2_10_l_14);
not I_17(n27_14,n28_14);
nor I_18(n28_14,IN_2_0_l_14,n43_14);
not I_19(n29_14,n33_14);
not I_20(n30_14,n31_14);
nor I_21(n31_14,IN_1_3_l_14,n46_14);
and I_22(n32_14,n33_14,n34_14);
nand I_23(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_24(n34_14,n42_14,n43_14);
nor I_25(n35_14,IN_1_8_l_14,IN_3_8_l_14);
nor I_26(n36_14,n47_14,n34_14);
not I_27(n37_14,n35_14);
nand I_28(n38_14,IN_2_8_l_14,IN_3_8_l_14);
nand I_29(n39_14,n29_14,n40_14);
nand I_30(n40_14,n27_14,n37_14);
nor I_31(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_32(n42_14,IN_3_0_l_14,IN_4_0_l_14);
not I_33(n43_14,IN_1_0_l_14);
nor I_34(n44_14,n27_14,n33_14);
or I_35(n45_14,IN_3_10_l_14,IN_4_10_l_14);
or I_36(n46_14,IN_2_3_l_14,IN_3_3_l_14);
not I_37(N1372_1_r_3,n40_3);
nor I_38(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_39(N1507_6_r_3,n31_3,n42_3);
nor I_40(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_41(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_42(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_43(n_573_7_r_3,n30_3,n31_3);
nor I_44(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_45(n_569_7_r_3,n30_3,n32_3);
nor I_46(n_452_7_r_3,n35_3,n_549_7_r_14);
not I_47(N6147_9_r_3,n32_3);
nor I_48(N6134_9_r_3,n36_3,n37_3);
not I_49(I_BUFF_1_9_r_3,n45_3);
nor I_50(n4_7_r_3,I_BUFF_1_9_r_3,n_549_7_r_14);
not I_51(n10_3,blif_reset_net_7_r_3);
not I_52(n30_3,n39_3);
not I_53(n31_3,n35_3);
nand I_54(n32_3,n41_3,n_573_7_r_14);
nor I_55(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_56(n34_3,n46_3,N1507_6_r_14);
nor I_57(n35_3,n43_3,n44_3);
not I_58(n36_3,n34_3);
nor I_59(n37_3,N6147_9_r_3,n_549_7_r_14);
or I_60(n38_3,n_572_7_r_3,n34_3);
nor I_61(n39_3,n44_3,N6147_9_r_14);
nand I_62(n40_3,n39_3,n_549_7_r_14);
nand I_63(n41_3,N1371_0_r_14,N1508_0_r_14);
nor I_64(n42_3,n34_3,n45_3);
not I_65(n43_3,n_452_7_r_14);
nor I_66(n44_3,n_572_7_r_14,N1371_0_r_14);
nand I_67(n45_3,n49_3,n50_3);
and I_68(n46_3,n47_3,N1508_0_r_14);
nand I_69(n47_3,n41_3,n48_3);
not I_70(n48_3,n_573_7_r_14);
nor I_71(n49_3,G42_7_r_14,n_569_7_r_14);
or I_72(n50_3,n51_3,N1507_6_r_14);
nor I_73(n51_3,N1508_6_r_14,N6134_9_r_14);
endmodule


