module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_5,blif_reset_net_7_r_5,N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_5,blif_reset_net_7_r_5;
output N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,n_549_7_r_5,n4_7_r_5,n7_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_7_r_5,n7_5,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N1371_0_r_5,n28_5,n46_5);
nand I_36(N1508_0_r_5,n26_5,n43_5);
not I_37(N1372_1_r_5,n43_5);
nor I_38(N1508_1_r_5,n30_5,n43_5);
nor I_39(N6147_2_r_5,n29_5,n32_5);
nor I_40(N1507_6_r_5,n26_5,n44_5);
nor I_41(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_42(n4_7_r_5,blif_clk_net_7_r_5,n7_5,G42_7_r_5,);
and I_43(n_572_7_r_5,n27_5,n28_5);
nand I_44(n_573_7_r_5,n26_5,n27_5);
nand I_45(n_549_7_r_5,G42_7_r_4,N1507_6_r_4);
nand I_46(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_47(n_452_7_r_5,n29_5);
nor I_48(n4_7_r_5,n30_5,n31_5);
not I_49(n7_5,blif_reset_net_7_r_5);
not I_50(n26_5,n35_5);
nand I_51(n27_5,n40_5,n41_5);
nand I_52(n28_5,n_452_7_r_4,n_569_7_r_4);
nand I_53(n29_5,n27_5,n33_5);
nor I_54(n30_5,n45_5,n_572_7_r_4);
not I_55(n31_5,n_549_7_r_5);
nor I_56(n32_5,n34_5,n35_5);
not I_57(n33_5,n30_5);
nor I_58(n34_5,n31_5,n36_5);
nor I_59(n35_5,n28_5,N6134_9_r_4);
not I_60(n36_5,n28_5);
nand I_61(n37_5,n36_5,n38_5);
nand I_62(n38_5,n26_5,n39_5);
nand I_63(n39_5,n30_5,n31_5);
nor I_64(n40_5,N1371_0_r_4,n_572_7_r_4);
or I_65(n41_5,n42_5,N1507_6_r_4);
nor I_66(n42_5,N1508_6_r_4,G42_7_r_4);
nand I_67(n43_5,n36_5,n46_5);
nor I_68(n44_5,n_549_7_r_5,n33_5);
or I_69(n45_5,N1371_0_r_4,n_549_7_r_4);
and I_70(n46_5,n31_5,n47_5);
or I_71(n47_5,n_569_7_r_4,n_549_7_r_4);
endmodule


