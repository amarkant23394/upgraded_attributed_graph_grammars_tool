module test_I15600(I15764,I1477,I1470,I11938,I13755,I14196,I15600);
input I15764,I1477,I1470,I11938,I13755,I14196;
output I15600;
wire I13908,I13767,I13743,I15832,I15815,I14162,I15628,I13749,I13891,I15611,I13775,I15781,I15798;
not I_0(I13908,I13891);
DFFARX1 I_1(I14196,I1470,I13775,,,I13767,);
DFFARX1 I_2(I13891,I1470,I13775,,,I13743,);
or I_3(I15600,I15832,I15815);
nand I_4(I15832,I15628,I13749);
DFFARX1 I_5(I15798,I1470,I15611,,,I15815,);
DFFARX1 I_6(I11938,I1470,I13775,,,I14162,);
not I_7(I15628,I13743);
nand I_8(I13749,I14162,I13908);
DFFARX1 I_9(I1470,I13775,,,I13891,);
not I_10(I15611,I1477);
not I_11(I13775,I1477);
and I_12(I15781,I15764,I13755);
or I_13(I15798,I15781,I13767);
endmodule


