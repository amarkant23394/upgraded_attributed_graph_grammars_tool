module test_I1492(I1215,I1423,I1455,I1492);
input I1215,I1423,I1455;
output I1492;
wire I1668,I1637,I1586,I1603,I1535;
not I_0(I1668,I1637);
not I_1(I1637,I1215);
nor I_2(I1586,I1535,I1215);
nand I_3(I1603,I1586,I1423);
not I_4(I1535,I1455);
nand I_5(I1492,I1603,I1668);
endmodule


