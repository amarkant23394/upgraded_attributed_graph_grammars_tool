module test_I7915(I1477,I1470,I7782,I3972,I6306,I7915);
input I1477,I1470,I7782,I3972,I6306;
output I7915;
wire I6606,I7898,I6300,I7799,I7816,I7881,I7570,I7587,I6329,I6688,I6705,I6291;
DFFARX1 I_0(I1470,I6329,,,I6606,);
nand I_1(I7898,I7881,I7816);
DFFARX1 I_2(I6606,I1470,I6329,,,I6300,);
or I_3(I7799,I7782,I6306);
DFFARX1 I_4(I7799,I1470,I7570,,,I7816,);
nand I_5(I7881,I7587,I6291);
not I_6(I7570,I1477);
not I_7(I7587,I6300);
not I_8(I6329,I1477);
DFFARX1 I_9(I1470,I6329,,,I6688,);
and I_10(I6705,I6688,I3972);
and I_11(I7915,I7881,I7898);
DFFARX1 I_12(I6705,I1470,I6329,,,I6291,);
endmodule


