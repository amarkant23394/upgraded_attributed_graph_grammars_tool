module Benchmark_testing500(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1539,I1546,I1573,I1564,I1561,I1567,I1555,I1549,I1570,I1558,I1552,I6993,I6996,I6972,I6984,I6999,I6987,I6981,I6975,I6978,I6990);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1539,I1546;
output I1573,I1564,I1561,I1567,I1555,I1549,I1570,I1558,I1552,I6993,I6996,I6972,I6984,I6999,I6987,I6981,I6975,I6978,I6990;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1539,I1546,I1581,I10559,I1607,I1624,I1632,I1649,I10562,I10568,I1666,I10577,I1692,I10580,I1737,I1745,I10571,I1762,I1802,I1810,I1855,I10586,I10565,I1872,I10574,I1898,I1906,I1937,I1954,I10583,I1971,I1988,I2005,I2036,I2108,I2134,I2142,I2159,I2176,I2202,I2219,I2227,I2244,I2076,I2275,I2292,I2088,I2332,I2097,I2354,I2371,I2397,I2414,I2100,I2436,I2085,I2467,I2484,I2501,I2518,I2094,I2549,I2082,I2091,I2079,I2635,I11166,I2661,I2669,I2686,I11160,I11181,I2703,I11157,I2729,I11178,I2746,I2754,I11175,I2771,I2603,I2802,I2819,I2615,I11163,I2859,I2624,I2881,I11172,I11169,I2898,I11154,I2924,I2941,I2627,I2963,I2612,I2994,I3011,I3028,I3045,I2621,I3076,I2609,I2618,I2606,I3162,I3188,I3196,I3213,I3230,I3256,I3273,I3281,I3298,I3130,I3329,I3346,I3142,I3386,I3151,I3408,I3425,I3451,I3468,I3154,I3490,I3139,I3521,I3538,I3555,I3572,I3148,I3603,I3136,I3145,I3133,I3692,I3718,I3726,I3743,I3769,I3660,I3791,I3817,I3825,I3842,I3868,I3684,I3890,I3666,I3930,I3947,I3955,I3972,I3669,I4003,I4020,I4046,I4054,I3657,I3675,I4099,I4116,I3678,I3663,I3672,I3681,I4216,I8825,I4242,I4250,I8831,I4276,I4284,I4301,I8828,I4318,I4335,I8846,I4352,I4202,I4383,I4400,I4417,I8849,I4434,I4199,I4190,I4479,I4193,I4187,I4524,I8834,I4541,I4558,I4196,I4589,I8840,I4606,I8837,I4623,I8843,I4649,I4657,I4184,I4208,I4702,I4719,I4736,I4205,I4794,I4820,I4828,I4845,I4862,I4888,I4896,I4922,I4930,I4947,I4964,I4981,I4777,I5021,I5029,I5046,I5063,I5080,I4780,I5111,I5128,I5154,I5162,I4762,I5193,I4771,I5224,I5241,I4783,I5272,I4774,I4765,I4768,I4786,I5372,I8270,I5398,I5406,I5423,I8267,I8285,I5440,I8282,I5466,I5474,I8264,I5500,I5508,I5525,I5542,I5559,I5355,I8276,I5599,I5607,I5624,I5641,I5658,I5358,I5689,I8279,I5706,I5732,I5740,I5340,I5771,I5349,I5802,I5819,I5361,I5850,I8273,I5352,I5343,I5346,I5364,I5947,I5973,I5981,I5998,I6015,I6041,I5936,I6072,I6080,I6097,I6123,I6131,I5939,I6171,I5930,I5921,I6207,I6224,I6250,I6258,I6275,I5924,I6306,I6323,I6340,I5933,I6371,I5918,I6402,I6419,I5927,I6474,I6500,I6508,I6525,I6542,I6568,I6463,I6599,I6607,I6624,I6650,I6658,I6466,I6698,I6457,I6448,I6734,I6751,I6777,I6785,I6802,I6451,I6833,I6850,I6867,I6460,I6898,I6445,I6929,I6946,I6454,I7007,I7033,I7050,I7058,I7075,I7092,I7109,I7126,I7143,I7174,I7191,I7222,I7239,I7256,I7287,I7327,I7335,I7352,I7369,I7386,I7417,I7434,I7451,I7477,I7499,I7516,I7547,I7592,I7653,I7679,I7696,I7704,I7721,I7738,I7755,I7772,I7789,I7639,I7820,I7837,I7642,I7868,I7885,I7902,I7618,I7933,I7630,I7973,I7981,I7998,I8015,I8032,I7645,I8063,I8080,I8097,I8123,I7633,I8145,I8162,I7627,I8193,I7621,I7624,I8238,I7636,I8293,I8319,I8336,I8358,I8384,I8392,I8409,I8426,I8443,I8460,I8477,I8494,I8525,I8556,I8573,I8590,I8607,I8638,I8683,I8700,I8717,I8743,I8751,I8782,I8799,I8857,I8883,I8891,I8931,I8939,I8956,I8973,I9013,I9035,I9052,I9078,I9086,I9103,I9120,I9137,I9154,I9199,I9230,I9247,I9273,I9281,I9312,I9329,I9346,I9363,I9435,I9461,I9469,I9418,I9509,I9517,I9534,I9551,I9406,I9591,I9427,I9613,I9630,I9656,I9664,I9681,I9698,I9715,I9732,I9403,I9424,I9777,I9415,I9808,I9825,I9851,I9859,I9421,I9890,I9907,I9924,I9941,I9412,I9409,I10013,I10039,I10047,I9996,I10087,I10095,I10112,I10129,I9984,I10169,I10005,I10191,I10208,I10234,I10242,I10259,I10276,I10293,I10310,I9981,I10002,I10355,I9993,I10386,I10403,I10429,I10437,I9999,I10468,I10485,I10502,I10519,I9990,I9987,I10594,I10620,I10637,I10645,I10690,I10707,I10724,I10741,I10758,I10775,I10792,I10823,I10840,I10885,I10902,I10919,I10950,I10976,I10984,I11015,I11032,I11049,I11075,I11083,I11100,I11189,I11215,I11232,I11240,I11285,I11302,I11319,I11336,I11353,I11370,I11387,I11418,I11435,I11480,I11497,I11514,I11545,I11571,I11579,I11610,I11627,I11644,I11670,I11678,I11695;
not I_0 (I1581,I1546);
DFFARX1 I_1 (I10559,I1539,I1581,I1607,);
DFFARX1 I_2 (I1607,I1539,I1581,I1624,);
not I_3 (I1632,I1624);
nand I_4 (I1649,I10562,I10568);
and I_5 (I1666,I1649,I10577);
DFFARX1 I_6 (I1666,I1539,I1581,I1692,);
DFFARX1 I_7 (I1692,I1539,I1581,I1573,);
DFFARX1 I_8 (I1692,I1539,I1581,I1564,);
DFFARX1 I_9 (I10580,I1539,I1581,I1737,);
nand I_10 (I1745,I1737,I10571);
not I_11 (I1762,I1745);
nor I_12 (I1561,I1607,I1762);
DFFARX1 I_13 (I10559,I1539,I1581,I1802,);
not I_14 (I1810,I1802);
nor I_15 (I1567,I1810,I1632);
nand I_16 (I1555,I1810,I1745);
nand I_17 (I1855,I10586,I10565);
and I_18 (I1872,I1855,I10574);
DFFARX1 I_19 (I1872,I1539,I1581,I1898,);
nor I_20 (I1906,I1898,I1607);
DFFARX1 I_21 (I1906,I1539,I1581,I1549,);
not I_22 (I1937,I1898);
nor I_23 (I1954,I10583,I10565);
not I_24 (I1971,I1954);
nor I_25 (I1988,I1745,I1971);
nor I_26 (I2005,I1937,I1988);
DFFARX1 I_27 (I2005,I1539,I1581,I1570,);
nor I_28 (I2036,I1898,I1971);
nor I_29 (I1558,I1762,I2036);
nor I_30 (I1552,I1898,I1954);
not I_31 (I2108,I1546);
DFFARX1 I_32 (I1532,I1539,I2108,I2134,);
not I_33 (I2142,I2134);
nand I_34 (I2159,I1364,I1444);
and I_35 (I2176,I2159,I1516);
DFFARX1 I_36 (I2176,I1539,I2108,I2202,);
DFFARX1 I_37 (I1460,I1539,I2108,I2219,);
and I_38 (I2227,I2219,I1524);
nor I_39 (I2244,I2202,I2227);
DFFARX1 I_40 (I2244,I1539,I2108,I2076,);
nand I_41 (I2275,I2219,I1524);
nand I_42 (I2292,I2142,I2275);
not I_43 (I2088,I2292);
DFFARX1 I_44 (I1492,I1539,I2108,I2332,);
DFFARX1 I_45 (I2332,I1539,I2108,I2097,);
nand I_46 (I2354,I1476,I1468);
and I_47 (I2371,I2354,I1412);
DFFARX1 I_48 (I2371,I1539,I2108,I2397,);
DFFARX1 I_49 (I2397,I1539,I2108,I2414,);
not I_50 (I2100,I2414);
not I_51 (I2436,I2397);
nand I_52 (I2085,I2436,I2275);
nor I_53 (I2467,I1388,I1468);
not I_54 (I2484,I2467);
nor I_55 (I2501,I2436,I2484);
nor I_56 (I2518,I2142,I2501);
DFFARX1 I_57 (I2518,I1539,I2108,I2094,);
nor I_58 (I2549,I2202,I2484);
nor I_59 (I2082,I2397,I2549);
nor I_60 (I2091,I2332,I2467);
nor I_61 (I2079,I2202,I2467);
not I_62 (I2635,I1546);
DFFARX1 I_63 (I11166,I1539,I2635,I2661,);
not I_64 (I2669,I2661);
nand I_65 (I2686,I11160,I11181);
and I_66 (I2703,I2686,I11157);
DFFARX1 I_67 (I2703,I1539,I2635,I2729,);
DFFARX1 I_68 (I11178,I1539,I2635,I2746,);
and I_69 (I2754,I2746,I11175);
nor I_70 (I2771,I2729,I2754);
DFFARX1 I_71 (I2771,I1539,I2635,I2603,);
nand I_72 (I2802,I2746,I11175);
nand I_73 (I2819,I2669,I2802);
not I_74 (I2615,I2819);
DFFARX1 I_75 (I11163,I1539,I2635,I2859,);
DFFARX1 I_76 (I2859,I1539,I2635,I2624,);
nand I_77 (I2881,I11172,I11169);
and I_78 (I2898,I2881,I11154);
DFFARX1 I_79 (I2898,I1539,I2635,I2924,);
DFFARX1 I_80 (I2924,I1539,I2635,I2941,);
not I_81 (I2627,I2941);
not I_82 (I2963,I2924);
nand I_83 (I2612,I2963,I2802);
nor I_84 (I2994,I11154,I11169);
not I_85 (I3011,I2994);
nor I_86 (I3028,I2963,I3011);
nor I_87 (I3045,I2669,I3028);
DFFARX1 I_88 (I3045,I1539,I2635,I2621,);
nor I_89 (I3076,I2729,I3011);
nor I_90 (I2609,I2924,I3076);
nor I_91 (I2618,I2859,I2994);
nor I_92 (I2606,I2729,I2994);
not I_93 (I3162,I1546);
DFFARX1 I_94 (I1500,I1539,I3162,I3188,);
not I_95 (I3196,I3188);
nand I_96 (I3213,I1404,I1420);
and I_97 (I3230,I3213,I1508);
DFFARX1 I_98 (I3230,I1539,I3162,I3256,);
DFFARX1 I_99 (I1396,I1539,I3162,I3273,);
and I_100 (I3281,I3273,I1484);
nor I_101 (I3298,I3256,I3281);
DFFARX1 I_102 (I3298,I1539,I3162,I3130,);
nand I_103 (I3329,I3273,I1484);
nand I_104 (I3346,I3196,I3329);
not I_105 (I3142,I3346);
DFFARX1 I_106 (I1436,I1539,I3162,I3386,);
DFFARX1 I_107 (I3386,I1539,I3162,I3151,);
nand I_108 (I3408,I1372,I1380);
and I_109 (I3425,I3408,I1452);
DFFARX1 I_110 (I3425,I1539,I3162,I3451,);
DFFARX1 I_111 (I3451,I1539,I3162,I3468,);
not I_112 (I3154,I3468);
not I_113 (I3490,I3451);
nand I_114 (I3139,I3490,I3329);
nor I_115 (I3521,I1428,I1380);
not I_116 (I3538,I3521);
nor I_117 (I3555,I3490,I3538);
nor I_118 (I3572,I3196,I3555);
DFFARX1 I_119 (I3572,I1539,I3162,I3148,);
nor I_120 (I3603,I3256,I3538);
nor I_121 (I3136,I3451,I3603);
nor I_122 (I3145,I3386,I3521);
nor I_123 (I3133,I3256,I3521);
not I_124 (I3692,I1546);
DFFARX1 I_125 (I3133,I1539,I3692,I3718,);
nand I_126 (I3726,I3145,I3154);
and I_127 (I3743,I3726,I3133);
DFFARX1 I_128 (I3743,I1539,I3692,I3769,);
nor I_129 (I3660,I3769,I3718);
not I_130 (I3791,I3769);
DFFARX1 I_131 (I3148,I1539,I3692,I3817,);
nand I_132 (I3825,I3817,I3136);
not I_133 (I3842,I3825);
DFFARX1 I_134 (I3842,I1539,I3692,I3868,);
not I_135 (I3684,I3868);
nor I_136 (I3890,I3718,I3825);
nor I_137 (I3666,I3769,I3890);
DFFARX1 I_138 (I3139,I1539,I3692,I3930,);
DFFARX1 I_139 (I3930,I1539,I3692,I3947,);
not I_140 (I3955,I3947);
not I_141 (I3972,I3930);
nand I_142 (I3669,I3972,I3791);
nand I_143 (I4003,I3130,I3130);
and I_144 (I4020,I4003,I3142);
DFFARX1 I_145 (I4020,I1539,I3692,I4046,);
nor I_146 (I4054,I4046,I3718);
DFFARX1 I_147 (I4054,I1539,I3692,I3657,);
DFFARX1 I_148 (I4046,I1539,I3692,I3675,);
nor I_149 (I4099,I3151,I3130);
not I_150 (I4116,I4099);
nor I_151 (I3678,I3955,I4116);
nand I_152 (I3663,I3972,I4116);
nor I_153 (I3672,I3718,I4099);
DFFARX1 I_154 (I4099,I1539,I3692,I3681,);
not I_155 (I4216,I1546);
DFFARX1 I_156 (I8825,I1539,I4216,I4242,);
not I_157 (I4250,I4242);
DFFARX1 I_158 (I8831,I1539,I4216,I4276,);
not I_159 (I4284,I8825);
nand I_160 (I4301,I4284,I8828);
not I_161 (I4318,I4301);
nor I_162 (I4335,I4318,I8846);
nor I_163 (I4352,I4250,I4335);
DFFARX1 I_164 (I4352,I1539,I4216,I4202,);
not I_165 (I4383,I8846);
nand I_166 (I4400,I4383,I4318);
and I_167 (I4417,I4383,I8849);
nand I_168 (I4434,I4417,I8828);
nor I_169 (I4199,I4434,I4383);
and I_170 (I4190,I4276,I4434);
not I_171 (I4479,I4434);
nand I_172 (I4193,I4276,I4479);
nor I_173 (I4187,I4242,I4434);
not I_174 (I4524,I8834);
nor I_175 (I4541,I4524,I8849);
nand I_176 (I4558,I4541,I4383);
nor I_177 (I4196,I4301,I4558);
nor I_178 (I4589,I4524,I8840);
and I_179 (I4606,I4589,I8837);
or I_180 (I4623,I4606,I8843);
DFFARX1 I_181 (I4623,I1539,I4216,I4649,);
nor I_182 (I4657,I4649,I4400);
DFFARX1 I_183 (I4657,I1539,I4216,I4184,);
DFFARX1 I_184 (I4649,I1539,I4216,I4208,);
not I_185 (I4702,I4649);
nor I_186 (I4719,I4702,I4276);
nor I_187 (I4736,I4541,I4719);
DFFARX1 I_188 (I4736,I1539,I4216,I4205,);
not I_189 (I4794,I1546);
DFFARX1 I_190 (I3681,I1539,I4794,I4820,);
not I_191 (I4828,I4820);
nand I_192 (I4845,I3684,I3660);
and I_193 (I4862,I4845,I3657);
DFFARX1 I_194 (I4862,I1539,I4794,I4888,);
not I_195 (I4896,I3663);
DFFARX1 I_196 (I3657,I1539,I4794,I4922,);
not I_197 (I4930,I4922);
nor I_198 (I4947,I4930,I4828);
and I_199 (I4964,I4947,I3663);
nor I_200 (I4981,I4930,I4896);
nor I_201 (I4777,I4888,I4981);
DFFARX1 I_202 (I3666,I1539,I4794,I5021,);
nor I_203 (I5029,I5021,I4888);
not I_204 (I5046,I5029);
not I_205 (I5063,I5021);
nor I_206 (I5080,I5063,I4964);
DFFARX1 I_207 (I5080,I1539,I4794,I4780,);
nand I_208 (I5111,I3669,I3678);
and I_209 (I5128,I5111,I3675);
DFFARX1 I_210 (I5128,I1539,I4794,I5154,);
nor I_211 (I5162,I5154,I5021);
DFFARX1 I_212 (I5162,I1539,I4794,I4762,);
nand I_213 (I5193,I5154,I5063);
nand I_214 (I4771,I5046,I5193);
not I_215 (I5224,I5154);
nor I_216 (I5241,I5224,I4964);
DFFARX1 I_217 (I5241,I1539,I4794,I4783,);
nor I_218 (I5272,I3672,I3678);
or I_219 (I4774,I5021,I5272);
nor I_220 (I4765,I5154,I5272);
or I_221 (I4768,I4888,I5272);
DFFARX1 I_222 (I5272,I1539,I4794,I4786,);
not I_223 (I5372,I1546);
DFFARX1 I_224 (I8270,I1539,I5372,I5398,);
not I_225 (I5406,I5398);
nand I_226 (I5423,I8267,I8285);
and I_227 (I5440,I5423,I8282);
DFFARX1 I_228 (I5440,I1539,I5372,I5466,);
not I_229 (I5474,I8264);
DFFARX1 I_230 (I8267,I1539,I5372,I5500,);
not I_231 (I5508,I5500);
nor I_232 (I5525,I5508,I5406);
and I_233 (I5542,I5525,I8264);
nor I_234 (I5559,I5508,I5474);
nor I_235 (I5355,I5466,I5559);
DFFARX1 I_236 (I8276,I1539,I5372,I5599,);
nor I_237 (I5607,I5599,I5466);
not I_238 (I5624,I5607);
not I_239 (I5641,I5599);
nor I_240 (I5658,I5641,I5542);
DFFARX1 I_241 (I5658,I1539,I5372,I5358,);
nand I_242 (I5689,I8279,I8264);
and I_243 (I5706,I5689,I8270);
DFFARX1 I_244 (I5706,I1539,I5372,I5732,);
nor I_245 (I5740,I5732,I5599);
DFFARX1 I_246 (I5740,I1539,I5372,I5340,);
nand I_247 (I5771,I5732,I5641);
nand I_248 (I5349,I5624,I5771);
not I_249 (I5802,I5732);
nor I_250 (I5819,I5802,I5542);
DFFARX1 I_251 (I5819,I1539,I5372,I5361,);
nor I_252 (I5850,I8273,I8264);
or I_253 (I5352,I5599,I5850);
nor I_254 (I5343,I5732,I5850);
or I_255 (I5346,I5466,I5850);
DFFARX1 I_256 (I5850,I1539,I5372,I5364,);
not I_257 (I5947,I1546);
DFFARX1 I_258 (I5340,I1539,I5947,I5973,);
not I_259 (I5981,I5973);
nand I_260 (I5998,I5343,I5340);
and I_261 (I6015,I5998,I5352);
DFFARX1 I_262 (I6015,I1539,I5947,I6041,);
DFFARX1 I_263 (I6041,I1539,I5947,I5936,);
DFFARX1 I_264 (I5349,I1539,I5947,I6072,);
nand I_265 (I6080,I6072,I5355);
not I_266 (I6097,I6080);
DFFARX1 I_267 (I6097,I1539,I5947,I6123,);
not I_268 (I6131,I6123);
nor I_269 (I5939,I5981,I6131);
DFFARX1 I_270 (I5364,I1539,I5947,I6171,);
nor I_271 (I5930,I6171,I6041);
nor I_272 (I5921,I6171,I6097);
nand I_273 (I6207,I5358,I5346);
and I_274 (I6224,I6207,I5343);
DFFARX1 I_275 (I6224,I1539,I5947,I6250,);
not I_276 (I6258,I6250);
nand I_277 (I6275,I6258,I6171);
nand I_278 (I5924,I6258,I6080);
nor I_279 (I6306,I5361,I5346);
and I_280 (I6323,I6171,I6306);
nor I_281 (I6340,I6258,I6323);
DFFARX1 I_282 (I6340,I1539,I5947,I5933,);
nor I_283 (I6371,I5973,I6306);
DFFARX1 I_284 (I6371,I1539,I5947,I5918,);
nor I_285 (I6402,I6250,I6306);
not I_286 (I6419,I6402);
nand I_287 (I5927,I6419,I6275);
not I_288 (I6474,I1546);
DFFARX1 I_289 (I2627,I1539,I6474,I6500,);
not I_290 (I6508,I6500);
nand I_291 (I6525,I2603,I2612);
and I_292 (I6542,I6525,I2606);
DFFARX1 I_293 (I6542,I1539,I6474,I6568,);
DFFARX1 I_294 (I6568,I1539,I6474,I6463,);
DFFARX1 I_295 (I2624,I1539,I6474,I6599,);
nand I_296 (I6607,I6599,I2615);
not I_297 (I6624,I6607);
DFFARX1 I_298 (I6624,I1539,I6474,I6650,);
not I_299 (I6658,I6650);
nor I_300 (I6466,I6508,I6658);
DFFARX1 I_301 (I2609,I1539,I6474,I6698,);
nor I_302 (I6457,I6698,I6568);
nor I_303 (I6448,I6698,I6624);
nand I_304 (I6734,I2621,I2618);
and I_305 (I6751,I6734,I2606);
DFFARX1 I_306 (I6751,I1539,I6474,I6777,);
not I_307 (I6785,I6777);
nand I_308 (I6802,I6785,I6698);
nand I_309 (I6451,I6785,I6607);
nor I_310 (I6833,I2603,I2618);
and I_311 (I6850,I6698,I6833);
nor I_312 (I6867,I6785,I6850);
DFFARX1 I_313 (I6867,I1539,I6474,I6460,);
nor I_314 (I6898,I6500,I6833);
DFFARX1 I_315 (I6898,I1539,I6474,I6445,);
nor I_316 (I6929,I6777,I6833);
not I_317 (I6946,I6929);
nand I_318 (I6454,I6946,I6802);
not I_319 (I7007,I1546);
DFFARX1 I_320 (I5924,I1539,I7007,I7033,);
DFFARX1 I_321 (I5921,I1539,I7007,I7050,);
not I_322 (I7058,I7050);
not I_323 (I7075,I5921);
nor I_324 (I7092,I7075,I5924);
not I_325 (I7109,I5936);
nor I_326 (I7126,I7092,I5930);
nor I_327 (I7143,I7050,I7126);
DFFARX1 I_328 (I7143,I1539,I7007,I6993,);
nor I_329 (I7174,I5930,I5924);
nand I_330 (I7191,I7174,I5921);
DFFARX1 I_331 (I7191,I1539,I7007,I6996,);
nor I_332 (I7222,I7109,I5930);
nand I_333 (I7239,I7222,I5918);
nor I_334 (I7256,I7033,I7239);
DFFARX1 I_335 (I7256,I1539,I7007,I6972,);
not I_336 (I7287,I7239);
nand I_337 (I6984,I7050,I7287);
DFFARX1 I_338 (I7239,I1539,I7007,I7327,);
not I_339 (I7335,I7327);
not I_340 (I7352,I5930);
not I_341 (I7369,I5927);
nor I_342 (I7386,I7369,I5936);
nor I_343 (I6999,I7335,I7386);
nor I_344 (I7417,I7369,I5933);
and I_345 (I7434,I7417,I5939);
or I_346 (I7451,I7434,I5918);
DFFARX1 I_347 (I7451,I1539,I7007,I7477,);
nor I_348 (I6987,I7477,I7033);
not I_349 (I7499,I7477);
and I_350 (I7516,I7499,I7033);
nor I_351 (I6981,I7058,I7516);
nand I_352 (I7547,I7499,I7109);
nor I_353 (I6975,I7369,I7547);
nand I_354 (I6978,I7499,I7287);
nand I_355 (I7592,I7109,I5927);
nor I_356 (I6990,I7352,I7592);
not I_357 (I7653,I1546);
DFFARX1 I_358 (I2076,I1539,I7653,I7679,);
DFFARX1 I_359 (I2082,I1539,I7653,I7696,);
not I_360 (I7704,I7696);
not I_361 (I7721,I2100);
nor I_362 (I7738,I7721,I2079);
not I_363 (I7755,I2085);
nor I_364 (I7772,I7738,I2091);
nor I_365 (I7789,I7696,I7772);
DFFARX1 I_366 (I7789,I1539,I7653,I7639,);
nor I_367 (I7820,I2091,I2079);
nand I_368 (I7837,I7820,I2100);
DFFARX1 I_369 (I7837,I1539,I7653,I7642,);
nor I_370 (I7868,I7755,I2091);
nand I_371 (I7885,I7868,I2097);
nor I_372 (I7902,I7679,I7885);
DFFARX1 I_373 (I7902,I1539,I7653,I7618,);
not I_374 (I7933,I7885);
nand I_375 (I7630,I7696,I7933);
DFFARX1 I_376 (I7885,I1539,I7653,I7973,);
not I_377 (I7981,I7973);
not I_378 (I7998,I2091);
not I_379 (I8015,I2079);
nor I_380 (I8032,I8015,I2085);
nor I_381 (I7645,I7981,I8032);
nor I_382 (I8063,I8015,I2088);
and I_383 (I8080,I8063,I2076);
or I_384 (I8097,I8080,I2094);
DFFARX1 I_385 (I8097,I1539,I7653,I8123,);
nor I_386 (I7633,I8123,I7679);
not I_387 (I8145,I8123);
and I_388 (I8162,I8145,I7679);
nor I_389 (I7627,I7704,I8162);
nand I_390 (I8193,I8145,I7755);
nor I_391 (I7621,I8015,I8193);
nand I_392 (I7624,I8145,I7933);
nand I_393 (I8238,I7755,I2079);
nor I_394 (I7636,I7998,I8238);
not I_395 (I8293,I1546);
DFFARX1 I_396 (I4184,I1539,I8293,I8319,);
DFFARX1 I_397 (I8319,I1539,I8293,I8336,);
not I_398 (I8285,I8336);
not I_399 (I8358,I8319);
DFFARX1 I_400 (I4199,I1539,I8293,I8384,);
nand I_401 (I8392,I8384,I4190);
not I_402 (I8409,I4190);
not I_403 (I8426,I4196);
nand I_404 (I8443,I4193,I4202);
and I_405 (I8460,I4193,I4202);
not I_406 (I8477,I4187);
nand I_407 (I8494,I8477,I8426);
nor I_408 (I8267,I8494,I8392);
nor I_409 (I8525,I8409,I8494);
nand I_410 (I8270,I8460,I8525);
not I_411 (I8556,I4184);
nor I_412 (I8573,I8556,I4193);
nor I_413 (I8590,I8573,I4187);
nor I_414 (I8607,I8358,I8590);
DFFARX1 I_415 (I8607,I1539,I8293,I8279,);
not I_416 (I8638,I8573);
DFFARX1 I_417 (I8638,I1539,I8293,I8282,);
and I_418 (I8276,I8384,I8573);
nor I_419 (I8683,I8556,I4208);
and I_420 (I8700,I8683,I4187);
or I_421 (I8717,I8700,I4205);
DFFARX1 I_422 (I8717,I1539,I8293,I8743,);
nor I_423 (I8751,I8743,I8477);
DFFARX1 I_424 (I8751,I1539,I8293,I8264,);
nand I_425 (I8782,I8743,I8384);
nand I_426 (I8799,I8477,I8782);
nor I_427 (I8273,I8799,I8443);
not I_428 (I8857,I1546);
DFFARX1 I_429 (I4777,I1539,I8857,I8883,);
and I_430 (I8891,I8883,I4765);
DFFARX1 I_431 (I8891,I1539,I8857,I8840,);
DFFARX1 I_432 (I4768,I1539,I8857,I8931,);
not I_433 (I8939,I4762);
not I_434 (I8956,I4786);
nand I_435 (I8973,I8956,I8939);
nor I_436 (I8828,I8931,I8973);
DFFARX1 I_437 (I8973,I1539,I8857,I9013,);
not I_438 (I8849,I9013);
not I_439 (I9035,I4774);
nand I_440 (I9052,I8956,I9035);
DFFARX1 I_441 (I9052,I1539,I8857,I9078,);
not I_442 (I9086,I9078);
not I_443 (I9103,I4783);
nand I_444 (I9120,I9103,I4780);
and I_445 (I9137,I8939,I9120);
nor I_446 (I9154,I9052,I9137);
DFFARX1 I_447 (I9154,I1539,I8857,I8825,);
DFFARX1 I_448 (I9137,I1539,I8857,I8846,);
nor I_449 (I9199,I4783,I4771);
nor I_450 (I8837,I9052,I9199);
or I_451 (I9230,I4783,I4771);
nor I_452 (I9247,I4762,I4765);
DFFARX1 I_453 (I9247,I1539,I8857,I9273,);
not I_454 (I9281,I9273);
nor I_455 (I8843,I9281,I9086);
nand I_456 (I9312,I9281,I8931);
not I_457 (I9329,I4762);
nand I_458 (I9346,I9329,I9035);
nand I_459 (I9363,I9281,I9346);
nand I_460 (I8834,I9363,I9312);
nand I_461 (I8831,I9346,I9230);
not I_462 (I9435,I1546);
DFFARX1 I_463 (I7624,I1539,I9435,I9461,);
and I_464 (I9469,I9461,I7618);
DFFARX1 I_465 (I9469,I1539,I9435,I9418,);
DFFARX1 I_466 (I7636,I1539,I9435,I9509,);
not I_467 (I9517,I7627);
not I_468 (I9534,I7639);
nand I_469 (I9551,I9534,I9517);
nor I_470 (I9406,I9509,I9551);
DFFARX1 I_471 (I9551,I1539,I9435,I9591,);
not I_472 (I9427,I9591);
not I_473 (I9613,I7645);
nand I_474 (I9630,I9534,I9613);
DFFARX1 I_475 (I9630,I1539,I9435,I9656,);
not I_476 (I9664,I9656);
not I_477 (I9681,I7621);
nand I_478 (I9698,I9681,I7642);
and I_479 (I9715,I9517,I9698);
nor I_480 (I9732,I9630,I9715);
DFFARX1 I_481 (I9732,I1539,I9435,I9403,);
DFFARX1 I_482 (I9715,I1539,I9435,I9424,);
nor I_483 (I9777,I7621,I7633);
nor I_484 (I9415,I9630,I9777);
or I_485 (I9808,I7621,I7633);
nor I_486 (I9825,I7618,I7630);
DFFARX1 I_487 (I9825,I1539,I9435,I9851,);
not I_488 (I9859,I9851);
nor I_489 (I9421,I9859,I9664);
nand I_490 (I9890,I9859,I9509);
not I_491 (I9907,I7618);
nand I_492 (I9924,I9907,I9613);
nand I_493 (I9941,I9859,I9924);
nand I_494 (I9412,I9941,I9890);
nand I_495 (I9409,I9924,I9808);
not I_496 (I10013,I1546);
DFFARX1 I_497 (I6448,I1539,I10013,I10039,);
and I_498 (I10047,I10039,I6454);
DFFARX1 I_499 (I10047,I1539,I10013,I9996,);
DFFARX1 I_500 (I6460,I1539,I10013,I10087,);
not I_501 (I10095,I6445);
not I_502 (I10112,I6445);
nand I_503 (I10129,I10112,I10095);
nor I_504 (I9984,I10087,I10129);
DFFARX1 I_505 (I10129,I1539,I10013,I10169,);
not I_506 (I10005,I10169);
not I_507 (I10191,I6463);
nand I_508 (I10208,I10112,I10191);
DFFARX1 I_509 (I10208,I1539,I10013,I10234,);
not I_510 (I10242,I10234);
not I_511 (I10259,I6457);
nand I_512 (I10276,I10259,I6448);
and I_513 (I10293,I10095,I10276);
nor I_514 (I10310,I10208,I10293);
DFFARX1 I_515 (I10310,I1539,I10013,I9981,);
DFFARX1 I_516 (I10293,I1539,I10013,I10002,);
nor I_517 (I10355,I6457,I6466);
nor I_518 (I9993,I10208,I10355);
or I_519 (I10386,I6457,I6466);
nor I_520 (I10403,I6451,I6451);
DFFARX1 I_521 (I10403,I1539,I10013,I10429,);
not I_522 (I10437,I10429);
nor I_523 (I9999,I10437,I10242);
nand I_524 (I10468,I10437,I10087);
not I_525 (I10485,I6451);
nand I_526 (I10502,I10485,I10191);
nand I_527 (I10519,I10437,I10502);
nand I_528 (I9990,I10519,I10468);
nand I_529 (I9987,I10502,I10386);
not I_530 (I10594,I1546);
DFFARX1 I_531 (I9984,I1539,I10594,I10620,);
DFFARX1 I_532 (I9996,I1539,I10594,I10637,);
not I_533 (I10645,I10637);
nor I_534 (I10562,I10620,I10645);
DFFARX1 I_535 (I10645,I1539,I10594,I10577,);
nor I_536 (I10690,I9993,I9987);
and I_537 (I10707,I10690,I9981);
nor I_538 (I10724,I10707,I9993);
not I_539 (I10741,I9993);
and I_540 (I10758,I10741,I9990);
nand I_541 (I10775,I10758,I9981);
nor I_542 (I10792,I10741,I10775);
DFFARX1 I_543 (I10792,I1539,I10594,I10559,);
not I_544 (I10823,I10775);
nand I_545 (I10840,I10645,I10823);
nand I_546 (I10571,I10707,I10823);
DFFARX1 I_547 (I10741,I1539,I10594,I10586,);
not I_548 (I10885,I10005);
nor I_549 (I10902,I10885,I9990);
nor I_550 (I10919,I10902,I10724);
DFFARX1 I_551 (I10919,I1539,I10594,I10583,);
not I_552 (I10950,I10902);
DFFARX1 I_553 (I10950,I1539,I10594,I10976,);
not I_554 (I10984,I10976);
nor I_555 (I10580,I10984,I10902);
nor I_556 (I11015,I10885,I9999);
and I_557 (I11032,I11015,I10002);
or I_558 (I11049,I11032,I9984);
DFFARX1 I_559 (I11049,I1539,I10594,I11075,);
not I_560 (I11083,I11075);
nand I_561 (I11100,I11083,I10823);
not I_562 (I10574,I11100);
nand I_563 (I10568,I11100,I10840);
nand I_564 (I10565,I11083,I10707);
not I_565 (I11189,I1546);
DFFARX1 I_566 (I9406,I1539,I11189,I11215,);
DFFARX1 I_567 (I9418,I1539,I11189,I11232,);
not I_568 (I11240,I11232);
nor I_569 (I11157,I11215,I11240);
DFFARX1 I_570 (I11240,I1539,I11189,I11172,);
nor I_571 (I11285,I9415,I9409);
and I_572 (I11302,I11285,I9403);
nor I_573 (I11319,I11302,I9415);
not I_574 (I11336,I9415);
and I_575 (I11353,I11336,I9412);
nand I_576 (I11370,I11353,I9403);
nor I_577 (I11387,I11336,I11370);
DFFARX1 I_578 (I11387,I1539,I11189,I11154,);
not I_579 (I11418,I11370);
nand I_580 (I11435,I11240,I11418);
nand I_581 (I11166,I11302,I11418);
DFFARX1 I_582 (I11336,I1539,I11189,I11181,);
not I_583 (I11480,I9427);
nor I_584 (I11497,I11480,I9412);
nor I_585 (I11514,I11497,I11319);
DFFARX1 I_586 (I11514,I1539,I11189,I11178,);
not I_587 (I11545,I11497);
DFFARX1 I_588 (I11545,I1539,I11189,I11571,);
not I_589 (I11579,I11571);
nor I_590 (I11175,I11579,I11497);
nor I_591 (I11610,I11480,I9421);
and I_592 (I11627,I11610,I9424);
or I_593 (I11644,I11627,I9406);
DFFARX1 I_594 (I11644,I1539,I11189,I11670,);
not I_595 (I11678,I11670);
nand I_596 (I11695,I11678,I11418);
not I_597 (I11169,I11695);
nand I_598 (I11163,I11695,I11435);
nand I_599 (I11160,I11678,I11302);
endmodule


