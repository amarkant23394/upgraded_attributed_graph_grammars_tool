module test_I12653(I10961,I1477,I9474,I1470,I10766,I12653);
input I10961,I1477,I9474,I1470,I10766;
output I12653;
wire I11009,I10612,I10647,I10797,I11167,I11057,I11184,I10627,I10639,I9468,I11201,I11150,I12636;
DFFARX1 I_0(I9468,I1470,I10647,,,I11009,);
DFFARX1 I_1(I11009,I1470,I10647,,,I10612,);
not I_2(I10647,I1477);
not I_3(I10797,I10766);
not I_4(I11167,I11150);
nor I_5(I11057,I11009,I10797);
nand I_6(I11184,I11167);
nand I_7(I10627,I11167,I11057);
DFFARX1 I_8(I11201,I1470,I10647,,,I10639,);
DFFARX1 I_9(I1470,,,I9468,);
and I_10(I11201,I10961,I11184);
DFFARX1 I_11(I9474,I1470,I10647,,,I11150,);
nand I_12(I12636,I10612,I10639);
and I_13(I12653,I12636,I10627);
endmodule


