module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14,I_BUFF_1_9_r_14,N3_8_l_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
nor I_0(N1371_0_r_14,n47_14,n30_14);
nor I_1(N1508_0_r_14,n30_14,n41_14);
nor I_2(N1507_6_r_14,n37_14,n44_14);
nor I_3(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_4(n4_7_r_14,blif_clk_net_5_r_7,n6_7,G42_7_r_14,);
nor I_5(n_572_7_r_14,n28_14,n29_14);
nand I_6(n_573_7_r_14,n26_14,n27_14);
nor I_7(n_549_7_r_14,n31_14,n32_14);
nand I_8(n_569_7_r_14,n26_14,n30_14);
nor I_9(n_452_7_r_14,n47_14,n28_14);
nor I_10(N6147_9_r_14,n36_14,n37_14);
nor I_11(N6134_9_r_14,n28_14,n36_14);
not I_12(I_BUFF_1_9_r_14,n26_14);
and I_13(N3_8_l_14,IN_6_8_l_14,n38_14);
DFFARX1 I_14(N3_8_l_14,blif_clk_net_5_r_7,n6_7,n47_14,);
nor I_15(n4_7_r_14,n47_14,n35_14);
nand I_16(n26_14,IN_1_10_l_14,IN_2_10_l_14);
not I_17(n27_14,n28_14);
nor I_18(n28_14,IN_2_0_l_14,n43_14);
not I_19(n29_14,n33_14);
not I_20(n30_14,n31_14);
nor I_21(n31_14,IN_1_3_l_14,n46_14);
and I_22(n32_14,n33_14,n34_14);
nand I_23(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_24(n34_14,n42_14,n43_14);
nor I_25(n35_14,IN_1_8_l_14,IN_3_8_l_14);
nor I_26(n36_14,n47_14,n34_14);
not I_27(n37_14,n35_14);
nand I_28(n38_14,IN_2_8_l_14,IN_3_8_l_14);
nand I_29(n39_14,n29_14,n40_14);
nand I_30(n40_14,n27_14,n37_14);
nor I_31(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_32(n42_14,IN_3_0_l_14,IN_4_0_l_14);
not I_33(n43_14,IN_1_0_l_14);
nor I_34(n44_14,n27_14,n33_14);
or I_35(n45_14,IN_3_10_l_14,IN_4_10_l_14);
or I_36(n46_14,IN_2_3_l_14,IN_3_3_l_14);
nor I_37(N1371_0_r_7,n53_7,n52_7);
nor I_38(N1508_0_r_7,n51_7,n52_7);
nand I_39(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_40(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_41(n_576_5_r_7,n31_7,n32_7);
nor I_42(n_102_5_r_7,N1371_0_r_14,N1508_0_r_14);
nand I_43(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_44(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_45(n_572_7_r_7,n54_7,n33_7);
nand I_46(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_47(n_549_7_r_7,n53_7,n36_7);
nand I_48(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_49(n_452_7_r_7,N6147_9_r_14,N1507_6_r_14);
nor I_50(n4_7_l_7,N1508_6_r_14,n_569_7_r_14);
not I_51(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_52(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_53(n30_7,n53_7);
and I_54(N3_8_l_7,n50_7,N1371_0_r_14);
DFFARX1 I_55(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_56(n_431_5_r_7,n40_7,n41_7);
nor I_57(n4_7_r_7,n54_7,n49_7);
and I_58(n31_7,n_102_5_r_7,n39_7);
not I_59(n32_7,N1508_6_r_14);
nor I_60(n33_7,n34_7,G42_7_r_14);
and I_61(n34_7,n35_7,n_573_7_r_14);
not I_62(n35_7,N6134_9_r_14);
nor I_63(n36_7,n37_7,N1508_6_r_14);
or I_64(n37_7,n54_7,N1371_0_r_14);
or I_65(n38_7,N1508_0_r_14,n_452_7_r_14);
nor I_66(n39_7,n_452_7_r_7,n_549_7_r_14);
nand I_67(n40_7,n46_7,n47_7);
nand I_68(n41_7,n42_7,n43_7);
nor I_69(n42_7,n44_7,n45_7);
nor I_70(n43_7,N1508_0_r_14,n_452_7_r_14);
nor I_71(n44_7,N1507_6_r_14,N6134_9_r_14);
nor I_72(n45_7,G42_7_r_14,N1508_0_r_14);
nand I_73(n46_7,n35_7,n_573_7_r_14);
not I_74(n47_7,G42_7_r_14);
or I_75(n48_7,n_452_7_r_7,n_549_7_r_14);
not I_76(n49_7,n_452_7_r_7);
nand I_77(n50_7,N1508_0_r_14,n_572_7_r_14);
and I_78(n51_7,n_452_7_r_7,n45_7);
not I_79(n52_7,n44_7);
endmodule


