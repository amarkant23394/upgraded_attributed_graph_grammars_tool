module test_I17823(I15696,I1477,I15832,I1470,I17823);
input I15696,I1477,I15832,I1470;
output I17823;
wire I17563,I17413,I15597,I17775,I17532,I16052,I15585,I15959,I16162,I15928,I16069;
not I_0(I17563,I17532);
not I_1(I17413,I1477);
nor I_2(I15597,I15832,I16162);
DFFARX1 I_3(I15585,I1470,I17413,,,I17775,);
not I_4(I17532,I15597);
DFFARX1 I_5(I1470,,,I16052,);
nand I_6(I15585,I16069,I15959);
nor I_7(I15959,I15928,I15696);
nor I_8(I17823,I17775,I17563);
and I_9(I16162,I15696);
DFFARX1 I_10(I1470,,,I15928,);
not I_11(I16069,I16052);
endmodule


