module test_I9508(I1477,I5898,I5716,I8657,I8445,I1470,I9508);
input I1477,I5898,I5716,I8657,I8445,I1470;
output I9508;
wire I8202,I8753,I8496,I8623,I8770,I8674,I8216,I5719,I8377,I8250,I5737,I8360,I6203,I8736,I8462,I8267,I8199;
nand I_0(I8202,I8267,I8496);
not I_1(I8753,I8736);
nor I_2(I8496,I8462,I8377);
DFFARX1 I_3(I1470,I8216,,,I8623,);
nand I_4(I9508,I8199,I8202);
or I_5(I8770,I8753,I8674);
and I_6(I8674,I8623,I8657);
not I_7(I8216,I1477);
DFFARX1 I_8(I1470,,,I5719,);
not I_9(I8377,I8360);
nor I_10(I8250,I5719,I5716);
nand I_11(I5737,I6203,I5898);
not I_12(I8360,I5719);
DFFARX1 I_13(I1470,,,I6203,);
DFFARX1 I_14(I1470,I8216,,,I8736,);
DFFARX1 I_15(I8445,I1470,I8216,,,I8462,);
nand I_16(I8267,I8250,I5737);
DFFARX1 I_17(I8770,I1470,I8216,,,I8199,);
endmodule


