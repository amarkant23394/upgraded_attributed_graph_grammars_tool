module test_I8196(I6265,I1477,I1470,I4533,I8196);
input I6265,I1477,I1470,I4533;
output I8196;
wire I8216,I8360,I5751,I6110,I8623,I5743,I6028,I6127,I6079,I5802,I5719,I8377;
not I_0(I8216,I1477);
not I_1(I8360,I5719);
not I_2(I5751,I1477);
DFFARX1 I_3(I1470,I5751,,,I6110,);
DFFARX1 I_4(I5743,I1470,I8216,,,I8623,);
nand I_5(I5743,I6127,I6079);
DFFARX1 I_6(I1470,I5751,,,I6028,);
and I_7(I6127,I6110,I4533);
nand I_8(I8196,I8623,I8377);
nor I_9(I6079,I6028,I5802);
DFFARX1 I_10(I1470,I5751,,,I5802,);
DFFARX1 I_11(I6265,I1470,I5751,,,I5719,);
not I_12(I8377,I8360);
endmodule


