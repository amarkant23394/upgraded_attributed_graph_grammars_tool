module test_final(IN_1_0_l_6,IN_2_0_l_6,IN_3_0_l_6,IN_4_0_l_6,IN_1_1_l_6,IN_2_1_l_6,IN_3_1_l_6,IN_1_10_l_6,IN_2_10_l_6,IN_3_10_l_6,IN_4_10_l_6,blif_clk_net_5_r_4,blif_reset_net_5_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4);
input IN_1_0_l_6,IN_2_0_l_6,IN_3_0_l_6,IN_4_0_l_6,IN_1_1_l_6,IN_2_1_l_6,IN_3_1_l_6,IN_1_10_l_6,IN_2_10_l_6,IN_3_10_l_6,IN_4_10_l_6,blif_clk_net_5_r_4,blif_reset_net_5_r_4;
output N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4;
wire N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,n_429_or_0_5_r_6,G78_5_r_6,n_576_5_r_6,n_102_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6,n_431_5_r_6,n24_6,n25_6,n26_6,n27_6,n28_6,n29_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,N1371_0_r_4,n_102_5_r_4,n_431_5_r_4,n4_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4;
nor I_0(N1371_0_r_6,n26_6,n38_6);
not I_1(N1508_0_r_6,n38_6);
nor I_2(N6147_3_r_6,n30_6,n35_6);
nand I_3(n_429_or_0_5_r_6,n30_6,n32_6);
DFFARX1 I_4(n_431_5_r_6,blif_clk_net_5_r_4,n4_4,G78_5_r_6,);
nand I_5(n_576_5_r_6,n24_6,n25_6);
not I_6(n_102_5_r_6,n26_6);
or I_7(n_547_5_r_6,n_429_or_0_5_r_6,n26_6);
not I_8(N1372_10_r_6,n37_6);
nor I_9(N1508_10_r_6,n36_6,n37_6);
nand I_10(n_431_5_r_6,n_102_5_r_6,n28_6);
nor I_11(n24_6,n33_6,n34_6);
nor I_12(n25_6,n26_6,n27_6);
nor I_13(n26_6,IN_2_0_l_6,n40_6);
nand I_14(n27_6,IN_1_1_l_6,IN_2_1_l_6);
nand I_15(n28_6,n29_6,n30_6);
nor I_16(n29_6,IN_3_1_l_6,n31_6);
not I_17(n30_6,n27_6);
nor I_18(n31_6,n39_6,n40_6);
nor I_19(n32_6,IN_3_1_l_6,n24_6);
not I_20(n33_6,IN_1_10_l_6);
not I_21(n34_6,IN_2_10_l_6);
or I_22(n35_6,n26_6,n31_6);
and I_23(n36_6,IN_3_1_l_6,n38_6);
nand I_24(n37_6,n30_6,n31_6);
nand I_25(n38_6,IN_2_10_l_6,n41_6);
nor I_26(n39_6,IN_3_0_l_6,IN_4_0_l_6);
not I_27(n40_6,IN_1_0_l_6);
nor I_28(n41_6,n33_6,n42_6);
nor I_29(n42_6,IN_3_10_l_6,IN_4_10_l_6);
nor I_30(N1371_0_r_4,n25_4,n29_4);
nor I_31(N1508_0_r_4,n25_4,n32_4);
nor I_32(N6147_2_r_4,n24_4,n31_4);
or I_33(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_34(n_431_5_r_4,blif_clk_net_5_r_4,n4_4,G78_5_r_4,);
nand I_35(n_576_5_r_4,n22_4,n23_4);
nand I_36(n_102_5_r_4,n34_4,n35_4);
nand I_37(n_547_5_r_4,n26_4,n27_4);
nor I_38(N1507_6_r_4,n27_4,n30_4);
nor I_39(N1508_6_r_4,n30_4,n33_4);
nand I_40(n_431_5_r_4,n_102_5_r_4,n28_4);
not I_41(n4_4,blif_reset_net_5_r_4);
nor I_42(n22_4,n24_4,n25_4);
nor I_43(n23_4,n37_4,G78_5_r_6);
not I_44(n24_4,n_102_5_r_4);
nand I_45(n25_4,n_576_5_r_6,n_547_5_r_6);
nor I_46(n26_4,n23_4,n24_4);
not I_47(n27_4,n25_4);
nand I_48(n28_4,n23_4,n29_4);
nor I_49(n29_4,n25_4,N6147_3_r_6);
not I_50(n30_4,n29_4);
nor I_51(n31_4,N1371_0_r_4,n32_4);
nor I_52(n32_4,n23_4,n29_4);
nand I_53(n33_4,n23_4,n24_4);
nor I_54(n34_4,N1508_0_r_6,N6147_3_r_6);
or I_55(n35_4,n36_4,G78_5_r_6);
nor I_56(n36_4,N1371_0_r_6,N1372_10_r_6);
or I_57(n37_4,N1508_10_r_6,N1371_0_r_6);
endmodule


