module test_I11941(I1477,I1470,I12157,I10017,I11941);
input I1477,I1470,I12157,I10017;
output I11941;
wire I12208,I10023,I10052,I10137,I11973,I12174,I12191;
DFFARX1 I_0(I12191,I1470,I11973,,,I12208,);
DFFARX1 I_1(I10137,I1470,I10052,,,I10023,);
not I_2(I10052,I1477);
DFFARX1 I_3(I1470,I10052,,,I10137,);
not I_4(I11973,I1477);
and I_5(I12174,I12157,I10017);
or I_6(I12191,I12174,I10023);
DFFARX1 I_7(I12208,I1470,I11973,,,I11941,);
endmodule


