module test_I4246(I1415,I3217,I1477,I1470,I1359,I1407,I4246);
input I1415,I3217,I1477,I1470,I1359,I1407;
output I4246;
wire I3293,I3983,I3310,I2745,I2844,I2827,I2980,I2776;
not I_0(I3293,I3217);
not I_1(I3983,I1477);
and I_2(I3310,I2844,I3293);
nor I_3(I2745,I2980,I3310);
nand I_4(I2844,I2827,I1359);
nor I_5(I2827,I2776);
nand I_6(I2980,I2776,I1415);
not I_7(I2776,I1407);
DFFARX1 I_8(I2745,I1470,I3983,,,I4246,);
endmodule


