module test_I11327(I6893,I1470,I8862,I6896,I11327);
input I6893,I1470,I8862,I6896;
output I11327;
wire I7190,I8830,I8896,I8913,I6872,I8964,I8981,I9227,I9179,I6878;
DFFARX1 I_0(I1470,,,I7190,);
nand I_1(I8830,I8913,I9227);
nor I_2(I8896,I6893,I6872);
nand I_3(I8913,I8896,I6878);
DFFARX1 I_4(I1470,,,I6872,);
not I_5(I8964,I6893);
not I_6(I8981,I8964);
nor I_7(I9227,I9179,I8981);
DFFARX1 I_8(I6896,I1470,I8862,,,I9179,);
not I_9(I11327,I8830);
not I_10(I6878,I7190);
endmodule


