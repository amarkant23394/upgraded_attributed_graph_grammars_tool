module test_I3877(I1750,I1477,I1603,I1470,I1832,I3877);
input I1750,I1477,I1603,I1470,I1832;
output I3877;
wire I1518,I3388,I1486,I1504,I3470,I1880,I3453,I1501,I3747,I1897,I1767;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
DFFARX1 I_2(I1832,I1470,I1518,,,I1486,);
nand I_3(I1504,I1767,I1897);
not I_4(I3470,I3453);
DFFARX1 I_5(I1470,I1518,,,I1880,);
nor I_6(I3877,I3747,I3470);
nor I_7(I3453,I1486,I1501);
not I_8(I1501,I1880);
DFFARX1 I_9(I1504,I1470,I3388,,,I3747,);
nor I_10(I1897,I1880,I1603);
DFFARX1 I_11(I1750,I1470,I1518,,,I1767,);
endmodule


