module test_I11973(I1477,I11973);
input I1477;
output I11973;
wire ;
not I_0(I11973,I1477);
endmodule


