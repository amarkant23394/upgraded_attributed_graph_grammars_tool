module test_I12459(I10349,I1477,I10538,I1470,I10287,I12459);
input I10349,I1477,I10538,I1470,I10287;
output I12459;
wire I10038,I12425,I10020,I12106,I11973,I12442,I10052,I12123;
nand I_0(I10038,I10349,I10538);
DFFARX1 I_1(I10038,I1470,I11973,,,I12425,);
DFFARX1 I_2(I10287,I1470,I10052,,,I10020,);
not I_3(I12106,I10020);
not I_4(I11973,I1477);
not I_5(I12442,I12425);
not I_6(I10052,I1477);
not I_7(I12123,I12106);
nor I_8(I12459,I12442,I12123);
endmodule


