module test_I5300(I1477,I3521,I3572,I1668,I1504,I1603,I3453,I1470,I5300);
input I1477,I3521,I3572,I1668,I1504,I1603,I3453,I1470;
output I5300;
wire I3470,I3747,I3356,I1483,I3388,I5283,I1492,I1518,I3620,I1880,I3589,I3877,I3374;
not I_0(I3470,I3453);
DFFARX1 I_1(I1504,I1470,I3388,,,I3747,);
DFFARX1 I_2(I3589,I1470,I3388,,,I3356,);
DFFARX1 I_3(I1880,I1470,I1518,,,I1483,);
nor I_4(I5300,I5283,I3374);
not I_5(I3388,I1477);
not I_6(I5283,I3356);
nand I_7(I1492,I1603,I1668);
not I_8(I1518,I1477);
nor I_9(I3620,I1492,I1483);
DFFARX1 I_10(I1470,I1518,,,I1880,);
and I_11(I3589,I3521,I3572);
nor I_12(I3877,I3747,I3470);
nand I_13(I3374,I3620,I3877);
endmodule


