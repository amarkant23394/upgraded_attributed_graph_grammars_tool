module test_I12140(I1477,I10185,I1470,I12140);
input I1477,I10185,I1470;
output I12140;
wire I10219,I10014,I7541,I10052,I10202;
not I_0(I12140,I10014);
DFFARX1 I_1(I10202,I1470,I10052,,,I10219,);
DFFARX1 I_2(I10219,I1470,I10052,,,I10014,);
DFFARX1 I_3(I1470,,,I7541,);
not I_4(I10052,I1477);
and I_5(I10202,I10185,I7541);
endmodule


