module test_I3238(I3263,I2563,I1294,I1301,I3238);
input I3263,I2563,I1294,I1301;
output I3238;
wire I3297,I3560,I3379,I2548,I2583,I3280,I3577,I3246,I2566,I2945,I3543;
DFFARX1 I_0(I3577,I1294,I3246,,,I3238,);
nand I_1(I3297,I3280,I2563);
nand I_2(I3560,I3543,I3297);
not I_3(I3379,I2548);
DFFARX1 I_4(I2945,I1294,I2583,,,I2548,);
not I_5(I2583,I1301);
nor I_6(I3280,I2548);
and I_7(I3577,I3379,I3560);
not I_8(I3246,I1301);
not I_9(I2566,I2945);
DFFARX1 I_10(I1294,I2583,,,I2945,);
nand I_11(I3543,I3263,I2566);
endmodule


