module test_I1510(I1477,I1423,I1470,I1207,I1455,I1510);
input I1477,I1423,I1470,I1207,I1455;
output I1510;
wire I1518,I2038,I2072,I2021,I1586,I1603,I1832,I1535,I2055;
not I_0(I1518,I1477);
not I_1(I2038,I2021);
and I_2(I2072,I1832,I2055);
DFFARX1 I_3(I1470,I1518,,,I2021,);
nor I_4(I1586,I1535);
DFFARX1 I_5(I2072,I1470,I1518,,,I1510,);
nand I_6(I1603,I1586,I1423);
nand I_7(I1832,I1535,I1207);
not I_8(I1535,I1455);
nand I_9(I2055,I2038,I1603);
endmodule


