module test_I8193(I1477,I6127,I6079,I1470,I8193);
input I1477,I6127,I6079,I1470;
output I8193;
wire I8216,I8623,I8705,I5743;
not I_0(I8216,I1477);
DFFARX1 I_1(I5743,I1470,I8216,,,I8623,);
DFFARX1 I_2(I8623,I1470,I8216,,,I8705,);
nand I_3(I5743,I6127,I6079);
not I_4(I8193,I8705);
endmodule


