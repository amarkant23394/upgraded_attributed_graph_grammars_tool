module test_I12287(I1477,I10202,I10414,I10459,I1470,I12287);
input I1477,I10202,I10414,I10459,I1470;
output I12287;
wire I10507,I12024,I10032,I10029,I10219,I10014,I10490,I10052,I10366,I12270,I12007,I10044,I10020,I11990,I10137,I10287;
and I_0(I10507,I10490,I10366);
nand I_1(I12024,I12007,I10044);
nand I_2(I10032,I10137,I10414);
DFFARX1 I_3(I10459,I1470,I10052,,,I10029,);
DFFARX1 I_4(I10202,I1470,I10052,,,I10219,);
DFFARX1 I_5(I10219,I1470,I10052,,,I10014,);
DFFARX1 I_6(I1470,I10052,,,I10490,);
not I_7(I10052,I1477);
nand I_8(I10366,I10219);
nand I_9(I12270,I11990,I10014);
nand I_10(I12287,I12270,I12024);
nor I_11(I12007,I10020,I10029);
DFFARX1 I_12(I10507,I1470,I10052,,,I10044,);
DFFARX1 I_13(I10287,I1470,I10052,,,I10020,);
not I_14(I11990,I10032);
DFFARX1 I_15(I1470,I10052,,,I10137,);
and I_16(I10287,I10219);
endmodule


