module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_5_r_11,n9_11,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_5_r_11,n9_11,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
not I_40(N1372_1_r_11,n53_11);
nor I_41(N1508_1_r_11,n39_11,n53_11);
nor I_42(N6147_2_r_11,n48_11,n49_11);
nor I_43(N6147_3_r_11,n44_11,n45_11);
nand I_44(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_45(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_46(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_47(n_102_5_r_11,n39_11);
nand I_48(n_547_5_r_11,n36_11,n37_11);
nor I_49(N1507_6_r_11,n52_11,n57_11);
nor I_50(N1508_6_r_11,n46_11,n51_11);
nor I_51(N1372_10_r_11,n43_11,n47_11);
nor I_52(N1508_10_r_11,n55_11,n56_11);
nand I_53(n_431_5_r_11,n40_11,n41_11);
not I_54(n9_11,blif_reset_net_5_r_11);
nor I_55(n36_11,n38_11,n39_11);
not I_56(n37_11,n40_11);
nor I_57(n38_11,n60_11,N1371_0_r_8);
nor I_58(n39_11,n54_11,N6147_9_r_8);
nand I_59(n40_11,N1508_10_r_8,n_42_8_r_8);
nand I_60(n41_11,n_102_5_r_11,n42_11);
and I_61(n42_11,n58_11,G199_8_r_8);
not I_62(n43_11,n44_11);
nor I_63(n44_11,n40_11,N1371_0_r_8);
nand I_64(n45_11,n46_11,n47_11);
not I_65(n46_11,n38_11);
nand I_66(n47_11,n59_11,n62_11);
and I_67(n48_11,n37_11,n47_11);
or I_68(n49_11,n44_11,n50_11);
nor I_69(n50_11,n60_11,n61_11);
or I_70(n51_11,n_102_5_r_11,n52_11);
nor I_71(n52_11,n42_11,n57_11);
nand I_72(n53_11,n37_11,n50_11);
or I_73(n54_11,N1508_1_r_8,N1507_6_r_8);
nor I_74(n55_11,n38_11,n42_11);
not I_75(n56_11,N1372_10_r_11);
and I_76(n57_11,n38_11,n50_11);
and I_77(n58_11,n59_11,N1507_6_r_8);
or I_78(n59_11,n63_11,N1508_6_r_8);
not I_79(n60_11,G199_8_r_8);
nor I_80(n61_11,N1508_6_r_8,n_42_8_r_8);
nand I_81(n62_11,N6147_9_r_8,N6134_9_r_8);
and I_82(n63_11,N6147_9_r_8,N6134_9_r_8);
endmodule


