module test_I12619_rst(I1477_rst,I12619_rst);
,I12619_rst);
input I1477_rst;
output I12619_rst;
wire ;
not I_0(I12619_rst,I1477_rst);
endmodule


