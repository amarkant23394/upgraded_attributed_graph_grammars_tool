module test_I9258(I1477,I5097,I9049,I5070,I9083,I1470,I9258);
input I1477,I5097,I9049,I5070,I9083,I1470;
output I9258;
wire I6893,I9179,I9148,I9131,I6975,I6992,I7026,I9114,I8862,I7286,I6896,I9066,I7156,I8964;
nand I_0(I6893,I7156,I7286);
DFFARX1 I_1(I6896,I1470,I8862,,,I9179,);
and I_2(I9148,I8964,I9131);
nor I_3(I9131,I9066,I9114);
nor I_4(I6975,I5070);
nand I_5(I6992,I6975,I5097);
not I_6(I7026,I5070);
not I_7(I9114,I9083);
not I_8(I8862,I1477);
or I_9(I9258,I9179,I9148);
nor I_10(I7286,I6992);
nor I_11(I6896,I6992,I7026);
DFFARX1 I_12(I9049,I1470,I8862,,,I9066,);
DFFARX1 I_13(I1470,,,I7156,);
not I_14(I8964,I6893);
endmodule


