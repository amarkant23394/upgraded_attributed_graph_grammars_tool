module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_14,blif_reset_net_7_r_14,N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_14,blif_reset_net_7_r_14;
output N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,I_BUFF_1_9_r_14,N3_8_l_14,n8_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_7_r_14,n8_14,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_14,n47_14,n30_14);
nor I_37(N1508_0_r_14,n30_14,n41_14);
nor I_38(N1507_6_r_14,n37_14,n44_14);
nor I_39(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_40(n4_7_r_14,blif_clk_net_7_r_14,n8_14,G42_7_r_14,);
nor I_41(n_572_7_r_14,n28_14,n29_14);
nand I_42(n_573_7_r_14,n26_14,n27_14);
nor I_43(n_549_7_r_14,n31_14,n32_14);
nand I_44(n_569_7_r_14,n26_14,n30_14);
nor I_45(n_452_7_r_14,n47_14,n28_14);
nor I_46(N6147_9_r_14,n36_14,n37_14);
nor I_47(N6134_9_r_14,n28_14,n36_14);
not I_48(I_BUFF_1_9_r_14,n26_14);
and I_49(N3_8_l_14,n38_14,N6134_9_r_3);
not I_50(n8_14,blif_reset_net_7_r_14);
DFFARX1 I_51(N3_8_l_14,blif_clk_net_7_r_14,n8_14,n47_14,);
nor I_52(n4_7_r_14,n47_14,n35_14);
nand I_53(n26_14,G42_7_r_3,n_569_7_r_3);
not I_54(n27_14,n28_14);
nor I_55(n28_14,n43_14,N1372_1_r_3);
not I_56(n29_14,n33_14);
not I_57(n30_14,n31_14);
nor I_58(n31_14,n46_14,n_549_7_r_3);
and I_59(n32_14,n33_14,n34_14);
nand I_60(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_61(n34_14,n42_14,n43_14);
nor I_62(n35_14,N1508_1_r_3,N1507_6_r_3);
nor I_63(n36_14,n47_14,n34_14);
not I_64(n37_14,n35_14);
nand I_65(n38_14,N1508_1_r_3,G42_7_r_3);
nand I_66(n39_14,n29_14,n40_14);
nand I_67(n40_14,n27_14,n37_14);
nor I_68(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_69(n42_14,N1507_6_r_3,n_452_7_r_3);
not I_70(n43_14,N1508_6_r_3);
nor I_71(n44_14,n27_14,n33_14);
or I_72(n45_14,N1372_1_r_3,n_573_7_r_3);
or I_73(n46_14,N1508_6_r_3,n_573_7_r_3);
endmodule


