module test_final(IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_102_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13,n4_7_l_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_13,n59_13,n61_13);
nor I_1(N1508_0_r_13,n59_13,n60_13);
not I_2(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_3(n_431_5_r_13,blif_clk_net_8_r_10,n11_10,G78_5_r_13,);
nand I_4(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_5(n_102_5_r_13,IN_9_7_l_13,IN_10_7_l_13);
nand I_6(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_7(n1_13,blif_clk_net_8_r_10,n11_10,G42_7_r_13,);
nor I_8(n_572_7_r_13,n40_13,n41_13);
nand I_9(n_573_7_r_13,n37_13,n38_13);
nor I_10(n_549_7_r_13,n46_13,n47_13);
nand I_11(n_569_7_r_13,n37_13,n43_13);
nand I_12(n_452_7_r_13,n52_13,n53_13);
nor I_13(n4_7_l_13,G18_7_l_13,IN_1_7_l_13);
DFFARX1 I_14(n4_7_l_13,blif_clk_net_8_r_10,n11_10,n62_13,);
not I_15(n33_13,n62_13);
nand I_16(n_431_5_r_13,n54_13,n55_13);
not I_17(n1_13,n52_13);
nor I_18(n34_13,n35_13,n36_13);
nor I_19(n35_13,G15_7_l_13,n42_13);
nand I_20(n36_13,n50_13,n58_13);
nand I_21(n37_13,n44_13,n45_13);
or I_22(n38_13,IN_3_1_l_13,n39_13);
nand I_23(n39_13,IN_1_1_l_13,IN_2_1_l_13);
not I_24(n40_13,n36_13);
nor I_25(n41_13,IN_10_7_l_13,n35_13);
not I_26(n42_13,IN_4_7_l_13);
or I_27(n43_13,G18_7_l_13,IN_5_7_l_13);
not I_28(n44_13,G15_7_l_13);
not I_29(n45_13,IN_7_7_l_13);
nor I_30(n46_13,n39_13,n40_13);
nor I_31(n47_13,G18_7_l_13,IN_5_7_l_13);
nor I_32(n48_13,n50_13,n51_13);
nor I_33(n49_13,G15_7_l_13,IN_7_7_l_13);
not I_34(n50_13,n59_13);
not I_35(n51_13,n_102_5_r_13);
nand I_36(n52_13,n33_13,n39_13);
nand I_37(n53_13,IN_3_1_l_13,n33_13);
nor I_38(n54_13,IN_5_7_l_13,IN_9_7_l_13);
nand I_39(n55_13,n62_13,n56_13);
nor I_40(n56_13,n39_13,n57_13);
not I_41(n57_13,G18_7_l_13);
or I_42(n58_13,IN_3_10_l_13,IN_4_10_l_13);
nand I_43(n59_13,IN_1_10_l_13,IN_2_10_l_13);
nor I_44(n60_13,IN_5_7_l_13,n51_13);
nor I_45(n61_13,IN_3_1_l_13,n39_13);
nor I_46(N1371_0_r_10,n37_10,n38_10);
nor I_47(N1508_0_r_10,n37_10,n58_10);
nand I_48(N6147_2_r_10,n39_10,n40_10);
not I_49(N6147_3_r_10,n39_10);
nor I_50(N1372_4_r_10,n46_10,n49_10);
nor I_51(N1508_4_r_10,n51_10,n52_10);
nor I_52(N1507_6_r_10,n49_10,n60_10);
nor I_53(N1508_6_r_10,n49_10,n50_10);
nor I_54(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_55(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_56(N6147_9_r_10,n36_10,n37_10);
nor I_57(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_58(I_BUFF_1_9_r_10,n48_10);
nor I_59(N3_8_r_10,n44_10,n47_10);
not I_60(n11_10,blif_reset_net_8_r_10);
not I_61(n35_10,n49_10);
nor I_62(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_63(n37_10,n_576_5_r_13);
not I_64(n38_10,n46_10);
nand I_65(n39_10,n43_10,n44_10);
nand I_66(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_67(n41_10,n42_10,n_576_5_r_13);
not I_68(n42_10,n44_10);
nor I_69(n43_10,n45_10,n_576_5_r_13);
nand I_70(n44_10,n54_10,G78_5_r_13);
nor I_71(n45_10,n59_10,n_573_7_r_13);
nand I_72(n46_10,n61_10,n_549_7_r_13);
nor I_73(n47_10,n46_10,n48_10);
nand I_74(n48_10,n62_10,n63_10);
nand I_75(n49_10,n56_10,N1508_0_r_13);
not I_76(n50_10,n45_10);
nor I_77(n51_10,n42_10,n53_10);
not I_78(n52_10,N1372_4_r_10);
nor I_79(n53_10,n48_10,n50_10);
and I_80(n54_10,n55_10,N1371_0_r_13);
nand I_81(n55_10,n56_10,n57_10);
nand I_82(n56_10,n_452_7_r_13,n_429_or_0_5_r_13);
not I_83(n57_10,N1508_0_r_13);
nor I_84(n58_10,n35_10,n45_10);
nor I_85(n59_10,n_429_or_0_5_r_13,G42_7_r_13);
nor I_86(n60_10,n37_10,n46_10);
or I_87(n61_10,n_429_or_0_5_r_13,G42_7_r_13);
nor I_88(n62_10,N1371_0_r_13,N1508_0_r_13);
or I_89(n63_10,n64_10,n_569_7_r_13);
nor I_90(n64_10,n_547_5_r_13,n_572_7_r_13);
endmodule


