module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_8_r_6,n9_6,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N1371_0_r_6,n30_6,n33_6);
nor I_37(N1508_0_r_6,n33_6,n44_6);
not I_38(N1372_1_r_6,n41_6);
nor I_39(N1508_1_r_6,n40_6,n41_6);
nor I_40(N1507_6_r_6,n39_6,n45_6);
nor I_41(N1508_6_r_6,n37_6,n38_6);
nor I_42(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_43(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_44(N6147_9_r_6,n32_6,n33_6);
nor I_45(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_46(I_BUFF_1_9_r_6,n37_6);
not I_47(N1372_10_r_6,n43_6);
nor I_48(N1508_10_r_6,n42_6,n43_6);
nor I_49(N3_8_r_6,n36_6,n_573_7_r_5);
not I_50(n9_6,blif_reset_net_8_r_6);
nor I_51(n30_6,n53_6,N1372_1_r_5);
not I_52(n31_6,n36_6);
nor I_53(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_54(n33_6,n_573_7_r_5);
not I_55(n34_6,n35_6);
nand I_56(n35_6,n49_6,G42_7_r_5);
nand I_57(n36_6,n51_6,N1508_6_r_5);
nand I_58(n37_6,n54_6,n_572_7_r_5);
or I_59(n38_6,n35_6,n39_6);
nor I_60(n39_6,n40_6,n45_6);
and I_61(n40_6,n46_6,n47_6);
nand I_62(n41_6,n30_6,n31_6);
nor I_63(n42_6,n34_6,n40_6);
nand I_64(n43_6,n30_6,n_573_7_r_5);
nor I_65(n44_6,n31_6,n40_6);
nor I_66(n45_6,n35_6,n36_6);
nor I_67(n46_6,N1508_0_r_5,N1372_1_r_5);
or I_68(n47_6,n48_6,n_569_7_r_5);
nor I_69(n48_6,N1507_6_r_5,N1371_0_r_5);
and I_70(n49_6,n50_6,N6147_2_r_5);
nand I_71(n50_6,n51_6,n52_6);
nand I_72(n51_6,N1371_0_r_5,N1508_1_r_5);
not I_73(n52_6,N1508_6_r_5);
nor I_74(n53_6,n_452_7_r_5,N1508_1_r_5);
or I_75(n54_6,n_452_7_r_5,N1508_1_r_5);
endmodule


