module test_I2702(I1316,I2005,I1294,I1301,I2702);
input I1316,I2005,I1294,I1301;
output I2702;
wire I1937,I2022,I2039,I1908;
not I_0(I1937,I1301);
nand I_1(I2022,I2005,I1316);
DFFARX1 I_2(I2022,I1294,I1937,,,I2039,);
not I_3(I1908,I2039);
not I_4(I2702,I1908);
endmodule


