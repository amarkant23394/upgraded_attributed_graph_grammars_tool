module test_I2849(I2600,I2781,I1908,I1294,I2505,I2457,I2406,I1301,I2849);
input I2600,I2781,I1908,I1294,I2505,I2457,I2406,I1301;
output I2849;
wire I2815,I2668,I2798,I1917,I1914,I2583,I2651,I1899,I1937,I2685,I2832;
or I_0(I2815,I2798,I1917);
nand I_1(I2668,I2651,I1914);
and I_2(I2798,I2781,I1899);
nand I_3(I1917,I2406,I2505);
DFFARX1 I_4(I2457,I1294,I1937,,,I1914,);
not I_5(I2583,I1301);
nor I_6(I2651,I2600,I1908);
DFFARX1 I_7(I1294,I1937,,,I1899,);
not I_8(I1937,I1301);
nor I_9(I2849,I2832,I2685);
not I_10(I2685,I2668);
DFFARX1 I_11(I2815,I1294,I2583,,,I2832,);
endmodule


