module test_I2733(I1937,I2022,I1294,I2733);
input I1937,I2022,I1294;
output I2733;
wire I2039,I1908,I2702;
not I_0(I2733,I2702);
DFFARX1 I_1(I2022,I1294,I1937,,,I2039,);
not I_2(I1908,I2039);
not I_3(I2702,I1908);
endmodule


