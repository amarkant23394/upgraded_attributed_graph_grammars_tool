module test_I13214(I9320,I1477,I11830,I1470,I9210,I11395,I11327,I13214);
input I9320,I1477,I11830,I1470,I9210,I11395,I11327;
output I13214;
wire I11672,I8827,I8836,I11275,I11302,I11847,I11310,I11864,I11624;
nand I_0(I13214,I11275,I11302);
DFFARX1 I_1(I8836,I1470,I11310,,,I11672,);
DFFARX1 I_2(I1470,,,I8827,);
nand I_3(I8836,I9320,I9210);
DFFARX1 I_4(I11672,I1470,I11310,,,I11275,);
DFFARX1 I_5(I11864,I1470,I11310,,,I11302,);
nand I_6(I11847,I11830,I11395);
not I_7(I11310,I1477);
and I_8(I11864,I11624,I11847);
nand I_9(I11624,I11327,I8827);
endmodule


