module test_I1313(I1263,I1294,I1301,I1313);
input I1263,I1294,I1301;
output I1313;
wire I1342,I1427;
not I_0(I1342,I1301);
DFFARX1 I_1(I1263,I1294,I1342,,,I1427,);
DFFARX1 I_2(I1427,I1294,I1342,,,I1313,);
endmodule


