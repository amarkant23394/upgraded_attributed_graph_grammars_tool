module test_I5156(I3781,I1477,I3504,I3685,I1504,I1470,I5156);
input I3781,I1477,I3504,I3685,I1504,I1470;
output I5156;
wire I3521,I1495,I3815,I3747,I3388,I3846,I3405,I1480,I3371,I3380,I5139,I3359,I3798,I3555;
nor I_0(I3521,I3504,I1495);
DFFARX1 I_1(I1470,,,I1495,);
or I_2(I3815,I3405,I3798);
DFFARX1 I_3(I1504,I1470,I3388,,,I3747,);
nand I_4(I5156,I5139,I3371);
not I_5(I3388,I1477);
nor I_6(I3846,I3747,I3555);
or I_7(I3405,I1480,I1495);
DFFARX1 I_8(I1470,,,I1480,);
DFFARX1 I_9(I3815,I1470,I3388,,,I3371,);
nand I_10(I3380,I3521,I3846);
nor I_11(I5139,I3380,I3359);
DFFARX1 I_12(I3747,I1470,I3388,,,I3359,);
and I_13(I3798,I3685,I3781);
DFFARX1 I_14(I1470,I3388,,,I3555,);
endmodule


