module Benchmark_testing5000(I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I983,I991,I999,I1007,I1015,I1023,I1031,I1039,I1047,I1055,I1063,I1071,I1079,I1087,I1095,I1103,I1111,I1119,I1127,I1135,I1143,I1151,I1159,I1167,I1175,I1183,I1191,I1199,I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1598,I1605,I3725,I3731,I3716,I3734,I3737,I3719,I3722,I3728,I15033,I15042,I15045,I15036,I15030,I15024,I15027,I15039,I15021,I23589,I23604,I23607,I23592,I23595,I23601,I23598,I36666,I36651,I36645,I36648,I36654,I36663,I36660,I36657,I40474,I40459,I40453,I40456,I40462,I40471,I40468,I40465,I45710,I45695,I45689,I45692,I45698,I45707,I45704,I45701,I47614,I47599,I47593,I47596,I47602,I47611,I47608,I47605,I51898,I51883,I51877,I51880,I51886,I51895,I51892,I51889,I52359,I52353,I52374,I52356,I52368,I52362,I52371,I52365,I57626,I57623,I57638,I57635,I57641,I57644,I57629,I57632,I62369,I62366,I62381,I62378,I62384,I62387,I62372,I62375);
input I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I983,I991,I999,I1007,I1015,I1023,I1031,I1039,I1047,I1055,I1063,I1071,I1079,I1087,I1095,I1103,I1111,I1119,I1127,I1135,I1143,I1151,I1159,I1167,I1175,I1183,I1191,I1199,I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1598,I1605;
output I3725,I3731,I3716,I3734,I3737,I3719,I3722,I3728,I15033,I15042,I15045,I15036,I15030,I15024,I15027,I15039,I15021,I23589,I23604,I23607,I23592,I23595,I23601,I23598,I36666,I36651,I36645,I36648,I36654,I36663,I36660,I36657,I40474,I40459,I40453,I40456,I40462,I40471,I40468,I40465,I45710,I45695,I45689,I45692,I45698,I45707,I45704,I45701,I47614,I47599,I47593,I47596,I47602,I47611,I47608,I47605,I51898,I51883,I51877,I51880,I51886,I51895,I51892,I51889,I52359,I52353,I52374,I52356,I52368,I52362,I52371,I52365,I57626,I57623,I57638,I57635,I57641,I57644,I57629,I57632,I62369,I62366,I62381,I62378,I62384,I62387,I62372,I62375;
wire I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I983,I991,I999,I1007,I1015,I1023,I1031,I1039,I1047,I1055,I1063,I1071,I1079,I1087,I1095,I1103,I1111,I1119,I1127,I1135,I1143,I1151,I1159,I1167,I1175,I1183,I1191,I1199,I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1598,I1605,I1637,I1654,I21153,I21156,I1671,I21141,I21150,I1688,I1705,I1617,I1736,I21159,I1753,I1779,I1787,I1804,I1821,I21144,I1838,I1855,I1872,I1889,I1623,I1920,I1937,I1954,I21147,I1608,I1985,I2002,I2019,I1626,I1629,I2064,I1611,I1614,I2109,I1620,I2164,I2181,I51419,I51401,I2198,I51407,I51422,I2215,I2232,I2144,I2263,I51404,I51410,I2280,I2306,I2314,I2331,I2348,I51413,I2365,I2382,I2399,I2416,I2150,I2447,I2464,I2481,I51416,I2135,I2512,I2529,I2546,I2153,I2156,I2591,I2138,I2141,I2636,I2147,I2691,I2708,I2725,I2742,I2759,I2671,I2790,I2807,I2833,I2841,I2858,I2875,I2892,I2909,I2926,I2943,I2677,I2974,I2991,I3008,I2662,I3039,I3056,I3073,I2680,I2683,I3118,I2665,I2668,I3163,I2674,I3218,I3235,I7884,I3252,I7905,I7902,I3269,I3286,I3198,I3317,I7881,I7893,I3334,I7890,I3360,I3368,I3385,I3402,I7899,I3419,I3436,I3453,I3470,I3204,I3501,I3518,I3535,I7896,I7887,I3189,I3566,I3583,I3600,I3207,I3210,I3645,I3192,I3195,I3690,I3201,I3745,I3762,I48563,I48545,I3779,I48551,I48566,I3796,I3813,I3844,I48548,I48554,I3861,I3887,I3895,I3912,I3929,I48557,I3946,I3963,I3980,I3997,I4028,I4045,I4062,I48560,I4093,I4110,I4127,I4172,I4217,I4272,I4289,I13494,I4306,I13515,I13512,I4323,I4340,I4252,I4371,I13491,I13503,I4388,I13500,I4414,I4422,I4439,I4456,I13509,I4473,I4490,I4507,I4524,I4258,I4555,I4572,I4589,I13506,I13497,I4243,I4620,I4637,I4654,I4261,I4264,I4699,I4246,I4249,I4744,I4255,I4799,I4816,I38567,I38549,I4833,I38555,I38570,I4850,I4867,I4779,I4898,I38552,I38558,I4915,I4941,I4949,I4966,I4983,I38561,I5000,I5017,I5034,I5051,I4785,I5082,I5099,I5116,I38564,I4770,I5147,I5164,I5181,I4788,I4791,I5226,I4773,I4776,I5271,I4782,I5326,I5343,I8904,I5360,I8925,I8922,I5377,I5394,I5306,I5425,I8901,I8913,I5442,I8910,I5468,I5476,I5493,I5510,I8919,I5527,I5544,I5561,I5578,I5312,I5609,I5626,I5643,I8916,I8907,I5297,I5674,I5691,I5708,I5315,I5318,I5753,I5300,I5303,I5798,I5309,I5853,I5870,I67648,I67642,I5887,I67639,I5904,I5921,I5833,I5952,I67645,I67651,I5969,I5995,I6003,I6020,I6037,I67636,I6054,I6071,I6088,I6105,I5839,I6136,I6153,I6170,I67654,I5824,I6201,I6218,I6235,I5842,I5845,I6280,I5827,I5830,I6325,I5836,I6383,I6400,I70288,I6417,I70303,I70306,I6434,I6451,I6468,I6485,I70294,I70297,I6502,I70291,I6528,I6536,I6553,I6570,I6587,I6604,I6363,I6635,I70300,I6652,I6669,I6372,I6375,I6714,I6366,I6360,I6759,I6776,I6354,I6357,I6369,I6835,I6351,I6893,I6910,I69846,I6927,I69861,I69864,I6944,I6961,I6978,I6995,I69852,I69855,I7012,I69849,I7038,I7046,I7063,I7080,I7097,I7114,I6873,I7145,I69858,I7162,I7179,I6882,I6885,I7224,I6876,I6870,I7269,I7286,I6864,I6867,I6879,I7345,I6861,I7403,I7420,I63953,I63947,I7437,I63956,I63959,I7454,I7471,I7488,I7505,I63950,I7522,I7548,I7556,I7573,I63965,I7590,I7607,I7624,I7383,I7655,I63962,I7672,I63968,I7689,I7392,I7395,I7734,I7386,I7380,I7779,I7796,I7374,I7377,I7389,I7855,I7371,I7913,I7930,I74266,I7947,I74281,I74284,I7964,I7981,I7998,I8015,I74272,I74275,I8032,I74269,I8058,I8066,I8083,I8100,I8117,I8134,I8165,I74278,I8182,I8199,I8244,I8289,I8306,I8365,I8423,I8440,I61318,I61312,I8457,I61321,I61324,I8474,I8491,I8508,I8525,I61315,I8542,I8568,I8576,I8593,I61330,I8610,I8627,I8644,I8403,I8675,I61327,I8692,I61333,I8709,I8412,I8415,I8754,I8406,I8400,I8799,I8816,I8394,I8397,I8409,I8875,I8391,I8933,I8950,I21963,I21957,I8967,I21975,I8984,I9001,I9018,I9035,I21969,I21960,I9052,I9078,I9086,I9103,I21972,I9120,I9137,I9154,I9185,I21966,I9202,I9219,I9264,I9309,I9326,I9385,I9443,I9460,I25602,I25581,I9477,I25590,I25599,I9494,I9511,I9528,I9545,I25596,I9562,I25587,I9588,I9596,I9613,I25578,I9630,I9647,I9664,I9423,I9695,I25593,I9712,I25584,I9729,I9432,I9435,I9774,I9426,I9420,I9819,I9836,I9414,I9417,I9429,I9895,I9411,I9953,I9970,I35088,I35067,I9987,I35076,I35085,I10004,I10021,I10038,I10055,I35082,I10072,I35073,I10098,I10106,I10123,I35064,I10140,I10157,I10174,I9933,I10205,I35079,I10222,I35070,I10239,I9942,I9945,I10284,I9936,I9930,I10329,I10346,I9924,I9927,I9939,I10405,I9921,I10463,I10480,I10497,I10514,I10531,I10548,I10565,I10582,I10608,I10616,I10633,I10650,I10667,I10684,I10443,I10715,I10732,I10749,I10452,I10455,I10794,I10446,I10440,I10839,I10856,I10434,I10437,I10449,I10915,I10431,I10973,I10990,I11007,I11024,I11041,I11058,I11075,I11092,I11118,I11126,I11143,I11160,I11177,I11194,I10953,I11225,I11242,I11259,I10962,I10965,I11304,I10956,I10950,I11349,I11366,I10944,I10947,I10959,I11425,I10941,I11483,I11500,I31399,I31378,I11517,I31387,I31396,I11534,I11551,I11568,I11585,I31393,I11602,I31384,I11628,I11636,I11653,I31375,I11670,I11687,I11704,I11463,I11735,I31390,I11752,I31381,I11769,I11472,I11475,I11814,I11466,I11460,I11859,I11876,I11454,I11457,I11469,I11935,I11451,I11993,I12010,I72498,I12027,I72513,I72516,I12044,I12061,I12078,I12095,I72504,I72507,I12112,I72501,I12138,I12146,I12163,I12180,I12197,I12214,I11973,I12245,I72510,I12262,I12279,I11982,I11985,I12324,I11976,I11970,I12369,I12386,I11964,I11967,I11979,I12445,I11961,I12503,I12520,I35615,I35594,I12537,I35603,I35612,I12554,I12571,I12588,I12605,I35609,I12622,I35600,I12648,I12656,I12673,I35591,I12690,I12707,I12724,I12483,I12755,I35606,I12772,I35597,I12789,I12492,I12495,I12834,I12486,I12480,I12879,I12896,I12474,I12477,I12489,I12955,I12471,I13013,I13030,I13047,I13064,I13081,I13098,I13115,I13132,I13158,I13166,I13183,I13200,I13217,I13234,I12993,I13265,I13282,I13299,I13002,I13005,I13344,I12996,I12990,I13389,I13406,I12984,I12987,I12999,I13465,I12981,I13523,I13540,I58683,I58677,I13557,I58686,I58689,I13574,I13591,I13608,I13625,I58680,I13642,I13668,I13676,I13693,I58695,I13710,I13727,I13744,I13775,I58692,I13792,I58698,I13809,I13854,I13899,I13916,I13975,I14033,I14050,I46644,I46647,I14067,I46653,I46641,I14084,I14101,I14118,I14135,I46659,I46662,I14152,I46656,I14178,I14186,I14203,I14220,I14237,I14254,I14013,I14285,I46650,I14302,I14319,I14022,I14025,I14364,I14016,I14010,I14409,I14426,I14004,I14007,I14019,I14485,I14001,I14543,I14560,I68078,I14577,I68093,I68096,I14594,I14611,I14628,I14645,I68084,I68087,I14662,I68081,I14688,I14696,I14713,I14730,I14747,I14764,I14523,I14795,I68090,I14812,I14829,I14532,I14535,I14874,I14526,I14520,I14919,I14936,I14514,I14517,I14529,I14995,I14511,I15053,I15070,I61845,I61839,I15087,I61848,I61851,I15104,I15121,I15138,I15155,I61842,I15172,I15198,I15206,I15223,I61857,I15240,I15257,I15274,I15305,I61854,I15322,I61860,I15339,I15384,I15429,I15446,I15505,I15563,I15580,I46168,I46171,I15597,I46177,I46165,I15614,I15631,I15648,I15665,I46183,I46186,I15682,I46180,I15708,I15716,I15733,I15750,I15767,I15784,I15543,I15815,I46174,I15832,I15849,I15552,I15555,I15894,I15546,I15540,I15939,I15956,I15534,I15537,I15549,I16015,I15531,I16073,I16090,I70730,I16107,I70745,I70748,I16124,I16141,I16158,I16175,I70736,I70739,I16192,I70733,I16218,I16226,I16243,I16260,I16277,I16294,I16053,I16325,I70742,I16342,I16359,I16062,I16065,I16404,I16056,I16050,I16449,I16466,I16044,I16047,I16059,I16525,I16041,I16583,I16600,I74708,I16617,I74723,I74726,I16634,I16651,I16668,I16685,I74714,I74717,I16702,I74711,I16728,I16736,I16753,I16770,I16787,I16804,I16563,I16835,I74720,I16852,I16869,I16572,I16575,I16914,I16566,I16560,I16959,I16976,I16554,I16557,I16569,I17035,I16551,I17093,I17110,I54464,I54461,I17127,I54467,I54479,I17144,I17161,I17178,I17195,I54470,I17212,I54476,I17238,I17246,I17263,I54482,I17280,I17297,I17314,I17073,I17345,I54473,I17362,I17379,I17082,I17085,I17424,I17076,I17070,I17469,I17486,I17064,I17067,I17079,I17545,I17061,I17603,I17620,I17637,I17654,I17671,I17688,I17705,I17722,I17748,I17756,I17773,I17790,I17807,I17824,I17583,I17855,I17872,I17889,I17592,I17595,I17934,I17586,I17580,I17979,I17996,I17574,I17577,I17589,I18055,I17571,I18113,I18130,I18147,I18164,I18181,I18198,I18215,I18232,I18258,I18266,I18283,I18300,I18317,I18334,I18093,I18365,I18382,I18399,I18102,I18105,I18444,I18096,I18090,I18489,I18506,I18084,I18087,I18099,I18565,I18081,I18623,I18640,I39980,I39983,I18657,I39989,I39977,I18674,I18691,I18708,I18725,I39995,I39998,I18742,I39992,I18768,I18776,I18793,I18810,I18827,I18844,I18603,I18875,I39986,I18892,I18909,I18612,I18615,I18954,I18606,I18600,I18999,I19016,I18594,I18597,I18609,I19075,I18591,I19133,I19150,I26129,I26108,I19167,I26117,I26126,I19184,I19201,I19218,I19235,I26123,I19252,I26114,I19278,I19286,I19303,I26105,I19320,I19337,I19354,I19113,I19385,I26120,I19402,I26111,I19419,I19122,I19125,I19464,I19116,I19110,I19509,I19526,I19104,I19107,I19119,I19585,I19101,I19643,I19660,I77360,I19677,I77375,I77378,I19694,I19711,I19728,I19745,I77366,I77369,I19762,I77363,I19788,I19796,I19813,I19830,I19847,I19864,I19623,I19895,I77372,I19912,I19929,I19632,I19635,I19974,I19626,I19620,I20019,I20036,I19614,I19617,I19629,I20095,I19611,I20153,I20170,I41884,I41887,I20187,I41893,I41881,I20204,I20221,I20238,I20255,I41899,I41902,I20272,I41896,I20298,I20306,I20323,I20340,I20357,I20374,I20133,I20405,I41890,I20422,I20439,I20142,I20145,I20484,I20136,I20130,I20529,I20546,I20124,I20127,I20139,I20605,I20121,I20663,I20680,I20697,I20714,I20731,I20748,I20765,I20782,I20808,I20816,I20833,I20850,I20867,I20884,I20643,I20915,I20932,I20949,I20652,I20655,I20994,I20646,I20640,I21039,I21056,I20634,I20637,I20649,I21115,I20631,I21167,I21184,I32450,I32432,I21201,I32453,I21218,I32429,I32444,I21235,I21266,I21283,I21300,I32447,I21317,I32435,I21334,I21365,I32441,I21382,I32438,I21399,I21444,I21461,I21478,I21495,I21575,I21592,I68977,I68971,I21609,I68974,I21626,I68968,I21643,I21549,I21674,I21691,I21708,I68965,I68962,I21725,I21742,I21564,I21773,I21790,I68980,I21807,I21567,I21552,I21852,I21869,I21886,I21903,I21555,I21561,I21558,I21983,I22000,I22017,I22034,I22051,I22082,I22099,I22116,I22133,I22150,I22181,I22198,I22215,I22260,I22277,I22294,I22311,I22391,I22408,I49021,I22425,I49042,I22442,I49024,I49027,I22459,I22365,I22490,I22507,I22524,I49030,I49039,I22541,I49036,I22558,I22380,I22589,I22606,I49033,I22623,I22383,I22368,I22668,I22685,I22702,I22719,I22371,I22377,I22374,I22799,I22816,I22833,I22850,I22867,I22773,I22898,I22915,I22932,I22949,I22966,I22788,I22997,I23014,I23031,I22791,I22776,I23076,I23093,I23110,I23127,I22779,I22785,I22782,I23207,I23224,I57114,I57099,I23241,I57102,I23258,I57096,I57111,I23275,I23181,I23306,I23323,I23340,I23357,I23374,I23196,I23405,I57117,I23422,I57108,I57105,I23439,I23199,I23184,I23484,I23501,I23518,I23535,I23187,I23193,I23190,I23615,I23632,I59222,I59207,I23649,I59210,I23666,I59204,I59219,I23683,I23714,I23731,I23748,I23765,I23782,I23813,I59225,I23830,I59216,I59213,I23847,I23892,I23909,I23926,I23943,I24029,I24046,I37121,I37124,I24063,I37127,I37136,I24080,I24097,I24114,I24131,I37133,I37139,I24148,I24174,I23997,I24196,I24213,I24015,I24244,I24261,I24018,I24292,I37142,I24309,I24326,I37130,I24000,I24357,I24374,I24021,I24405,I24006,I24436,I24009,I24467,I24003,I24498,I24012,I24556,I24573,I24590,I24607,I24624,I24641,I24658,I24675,I24701,I24524,I24723,I24740,I24542,I24771,I24788,I24545,I24819,I24836,I24853,I24527,I24884,I24901,I24548,I24932,I24533,I24963,I24536,I24994,I24530,I25025,I24539,I25083,I25100,I44261,I44264,I25117,I44267,I44276,I25134,I25151,I25168,I25185,I44273,I44279,I25202,I25228,I25051,I25250,I25267,I25069,I25298,I25315,I25072,I25346,I44282,I25363,I25380,I44270,I25054,I25411,I25428,I25075,I25459,I25060,I25490,I25063,I25521,I25057,I25552,I25066,I25610,I25627,I71620,I71617,I25644,I71629,I71632,I25661,I25678,I25695,I25712,I71623,I71614,I25729,I25755,I25777,I25794,I25825,I25842,I25873,I25890,I25907,I71626,I25938,I25955,I25986,I26017,I26048,I26079,I26137,I26154,I67127,I67115,I26171,I67109,I26188,I26205,I26222,I26239,I67112,I26256,I67118,I26282,I26304,I26321,I26352,I67124,I26369,I26400,I67130,I26417,I26434,I67121,I26465,I26482,I26513,I26544,I26575,I26606,I26664,I26681,I26698,I26715,I26732,I26749,I26766,I26783,I26809,I26632,I26831,I26848,I26650,I26879,I26896,I26653,I26927,I26944,I26961,I26635,I26992,I27009,I26656,I27040,I26641,I27071,I26644,I27102,I26638,I27133,I26647,I27191,I27208,I59749,I59737,I27225,I59731,I27242,I27259,I27276,I27293,I59734,I27310,I59740,I27336,I27159,I27358,I27375,I27177,I27406,I59746,I27423,I27180,I27454,I59752,I27471,I27488,I59743,I27162,I27519,I27536,I27183,I27567,I27168,I27598,I27171,I27629,I27165,I27660,I27174,I27718,I27735,I71178,I71175,I27752,I71187,I71190,I27769,I27786,I27803,I27820,I71181,I71172,I27837,I27863,I27686,I27885,I27902,I27704,I27933,I27950,I27707,I27981,I27998,I28015,I71184,I27689,I28046,I28063,I27710,I28094,I27695,I28125,I27698,I28156,I27692,I28187,I27701,I28245,I28262,I28279,I28296,I28313,I28330,I28347,I28364,I28390,I28213,I28412,I28429,I28231,I28460,I28477,I28234,I28508,I28525,I28542,I28216,I28573,I28590,I28237,I28621,I28222,I28652,I28225,I28683,I28219,I28714,I28228,I28772,I28789,I28806,I28823,I28840,I28857,I28874,I28891,I28917,I28740,I28939,I28956,I28758,I28987,I29004,I28761,I29035,I29052,I29069,I28743,I29100,I29117,I28764,I29148,I28749,I29179,I28752,I29210,I28746,I29241,I28755,I29299,I29316,I58168,I58156,I29333,I58150,I29350,I29367,I29384,I29401,I58153,I29418,I58159,I29444,I29267,I29466,I29483,I29285,I29514,I58165,I29531,I29288,I29562,I58171,I29579,I29596,I58162,I29270,I29627,I29644,I29291,I29675,I29276,I29706,I29279,I29737,I29273,I29768,I29282,I29826,I29843,I29860,I29877,I29894,I29911,I29928,I29945,I29971,I29794,I29993,I30010,I29812,I30041,I30058,I29815,I30089,I30106,I30123,I29797,I30154,I30171,I29818,I30202,I29803,I30233,I29806,I30264,I29800,I30295,I29809,I30353,I30370,I42357,I42360,I30387,I42363,I42372,I30404,I30421,I30438,I30455,I42369,I42375,I30472,I30498,I30321,I30520,I30537,I30339,I30568,I30585,I30342,I30616,I42378,I30633,I30650,I42366,I30324,I30681,I30698,I30345,I30729,I30330,I30760,I30333,I30791,I30327,I30822,I30336,I30880,I30897,I56063,I56051,I30914,I56054,I56048,I30931,I30948,I30965,I30982,I56045,I30999,I56042,I31025,I30848,I31047,I31064,I30866,I31095,I31112,I30869,I31143,I31160,I31177,I56060,I56057,I30851,I31208,I31225,I30872,I31256,I30857,I31287,I30860,I31318,I30854,I31349,I30863,I31407,I31424,I72946,I72943,I31441,I72955,I72958,I31458,I31475,I31492,I31509,I72949,I72940,I31526,I31552,I31574,I31591,I31622,I31639,I31670,I31687,I31704,I72952,I31735,I31752,I31783,I31814,I31845,I31876,I31934,I31951,I31968,I31985,I32002,I32019,I32036,I32053,I32079,I31902,I32101,I32118,I31920,I32149,I32166,I31923,I32197,I32214,I32231,I31905,I32262,I32279,I31926,I32310,I31911,I32341,I31914,I32372,I31908,I32403,I31917,I32461,I32478,I42833,I42836,I32495,I42839,I42848,I32512,I32529,I32546,I32563,I42845,I42851,I32580,I32606,I32628,I32645,I32676,I32693,I32724,I42854,I32741,I32758,I42842,I32789,I32806,I32837,I32868,I32899,I32930,I32988,I33005,I33022,I33039,I33056,I33073,I33090,I33107,I33133,I32956,I33155,I33172,I32974,I33203,I33220,I32977,I33251,I33268,I33285,I32959,I33316,I33333,I32980,I33364,I32965,I33395,I32968,I33426,I32962,I33457,I32971,I33515,I33532,I49497,I49500,I33549,I49503,I49512,I33566,I33583,I33600,I33617,I49509,I49515,I33634,I33660,I33483,I33682,I33699,I33501,I33730,I33747,I33504,I33778,I49518,I33795,I33812,I49506,I33486,I33843,I33860,I33507,I33891,I33492,I33922,I33495,I33953,I33489,I33984,I33498,I34042,I34059,I50925,I50928,I34076,I50931,I50940,I34093,I34110,I34127,I34144,I50937,I50943,I34161,I34187,I34010,I34209,I34226,I34028,I34257,I34274,I34031,I34305,I50946,I34322,I34339,I50934,I34013,I34370,I34387,I34034,I34418,I34019,I34449,I34022,I34480,I34016,I34511,I34025,I34569,I34586,I66600,I66588,I34603,I66582,I34620,I34637,I34654,I34671,I66585,I34688,I66591,I34714,I34537,I34736,I34753,I34555,I34784,I66597,I34801,I34558,I34832,I66603,I34849,I34866,I66594,I34540,I34897,I34914,I34561,I34945,I34546,I34976,I34549,I35007,I34543,I35038,I34552,I35096,I35113,I35130,I35147,I35164,I35181,I35198,I35215,I35241,I35263,I35280,I35311,I35328,I35359,I35376,I35393,I35424,I35441,I35472,I35503,I35534,I35565,I35623,I35640,I50449,I50452,I35657,I50455,I50464,I35674,I35691,I35708,I35725,I50461,I50467,I35742,I35768,I35790,I35807,I35838,I35855,I35886,I50470,I35903,I35920,I50458,I35951,I35968,I35999,I36030,I36061,I36092,I36150,I36167,I36184,I36201,I36218,I36235,I36252,I36269,I36295,I36118,I36317,I36334,I36136,I36365,I36382,I36139,I36413,I36430,I36447,I36121,I36478,I36495,I36142,I36526,I36127,I36557,I36130,I36588,I36124,I36619,I36133,I36674,I36691,I36708,I36725,I36742,I36759,I36776,I36793,I36810,I36827,I36844,I36861,I36878,I36895,I36940,I36971,I37002,I37019,I37050,I37095,I37150,I37167,I73385,I73388,I37184,I37201,I73382,I73400,I37218,I37235,I73391,I37252,I37269,I37286,I37303,I37320,I73397,I73394,I37337,I37354,I37371,I37416,I37447,I37478,I37495,I37526,I37571,I37626,I37643,I56569,I56590,I37660,I56575,I37677,I56587,I37694,I56578,I37711,I56572,I37728,I37745,I37762,I37779,I37796,I56581,I56584,I37813,I37830,I37847,I37618,I37603,I37892,I37597,I37923,I37600,I37954,I37971,I37606,I38002,I37615,I37612,I38047,I37609,I38102,I38119,I38136,I38153,I38170,I38187,I38204,I38221,I38238,I38255,I38272,I38289,I38306,I38323,I38094,I38079,I38368,I38073,I38399,I38076,I38430,I38447,I38082,I38478,I38091,I38088,I38523,I38085,I38578,I38595,I38612,I38629,I38646,I38663,I38680,I38697,I38714,I38731,I38748,I38765,I38782,I38799,I38844,I38875,I38906,I38923,I38954,I38999,I39054,I39071,I39088,I39105,I39122,I39139,I39156,I39173,I39190,I39207,I39224,I39241,I39258,I39275,I39046,I39031,I39320,I39025,I39351,I39028,I39382,I39399,I39034,I39430,I39043,I39040,I39475,I39037,I39530,I39547,I39564,I39581,I39598,I39615,I39632,I39649,I39666,I39683,I39700,I39717,I39734,I39751,I39522,I39507,I39796,I39501,I39827,I39504,I39858,I39875,I39510,I39906,I39519,I39516,I39951,I39513,I40006,I40023,I60785,I60806,I40040,I60791,I40057,I60803,I40074,I60794,I40091,I60788,I40108,I40125,I40142,I40159,I40176,I60797,I60800,I40193,I40210,I40227,I40272,I40303,I40334,I40351,I40382,I40427,I40482,I40499,I40516,I40533,I40550,I40567,I40584,I40601,I40618,I40635,I40652,I40669,I40686,I40703,I40748,I40779,I40810,I40827,I40858,I40903,I40958,I40975,I40992,I41009,I41026,I41043,I41060,I41077,I41094,I41111,I41128,I41145,I41162,I41179,I40950,I40935,I41224,I40929,I41255,I40932,I41286,I41303,I40938,I41334,I40947,I40944,I41379,I40941,I41434,I41451,I41468,I41485,I41502,I41519,I41536,I41553,I41570,I41587,I41604,I41621,I41638,I41655,I41426,I41411,I41700,I41405,I41731,I41408,I41762,I41779,I41414,I41810,I41423,I41420,I41855,I41417,I41910,I41927,I41944,I41961,I41978,I41995,I42012,I42029,I42046,I42063,I42080,I42097,I42114,I42131,I42176,I42207,I42238,I42255,I42286,I42331,I42386,I42403,I42420,I42437,I42454,I42471,I42488,I42505,I42522,I42539,I42556,I42573,I42590,I42607,I42652,I42683,I42714,I42731,I42762,I42807,I42862,I42879,I72059,I72062,I42896,I42913,I72056,I72074,I42930,I42947,I72065,I42964,I42981,I42998,I43015,I43032,I72071,I72068,I43049,I43066,I43083,I43128,I43159,I43190,I43207,I43238,I43283,I43338,I43355,I66055,I66076,I43372,I66061,I43389,I66073,I43406,I66064,I43423,I66058,I43440,I43457,I43474,I43491,I43508,I66067,I66070,I43525,I43542,I43559,I43330,I43315,I43604,I43309,I43635,I43312,I43666,I43683,I43318,I43714,I43327,I43324,I43759,I43321,I43814,I43831,I76037,I76040,I43848,I43865,I76034,I76052,I43882,I43899,I76043,I43916,I43933,I43950,I43967,I43984,I76049,I76046,I44001,I44018,I44035,I43806,I43791,I44080,I43785,I44111,I43788,I44142,I44159,I43794,I44190,I43803,I43800,I44235,I43797,I44290,I44307,I44324,I44341,I44358,I44375,I44392,I44409,I44426,I44443,I44460,I44477,I44494,I44511,I44556,I44587,I44618,I44635,I44666,I44711,I44766,I44783,I75595,I75598,I44800,I44817,I75592,I75610,I44834,I44851,I75601,I44868,I44885,I44902,I44919,I44936,I75607,I75604,I44953,I44970,I44987,I44758,I44743,I45032,I44737,I45063,I44740,I45094,I45111,I44746,I45142,I44755,I44752,I45187,I44749,I45242,I45259,I45276,I45293,I45310,I45327,I45344,I45361,I45378,I45395,I45412,I45429,I45446,I45463,I45234,I45219,I45508,I45213,I45539,I45216,I45570,I45587,I45222,I45618,I45231,I45228,I45663,I45225,I45718,I45735,I45752,I45769,I45786,I45803,I45820,I45837,I45854,I45871,I45888,I45905,I45922,I45939,I45984,I46015,I46046,I46063,I46094,I46139,I46194,I46211,I53937,I53934,I46228,I53943,I46245,I53955,I53940,I46262,I46279,I53946,I46296,I46313,I46330,I46347,I46364,I53952,I46381,I53949,I46398,I46415,I46460,I46491,I46522,I46539,I46570,I46615,I46670,I46687,I46704,I46721,I46738,I46755,I46772,I46789,I46806,I46823,I46840,I46857,I46874,I46891,I46936,I46967,I46998,I47015,I47046,I47091,I47146,I47163,I76921,I76924,I47180,I47197,I76918,I76936,I47214,I47231,I76927,I47248,I47265,I47282,I47299,I47316,I76933,I76930,I47333,I47350,I47367,I47138,I47123,I47412,I47117,I47443,I47120,I47474,I47491,I47126,I47522,I47135,I47132,I47567,I47129,I47622,I47639,I65001,I65022,I47656,I65007,I47673,I65019,I47690,I65010,I47707,I65004,I47724,I47741,I47758,I47775,I47792,I65013,I65016,I47809,I47826,I47843,I47888,I47919,I47950,I47967,I47998,I48043,I48098,I48115,I54991,I54988,I48132,I54997,I48149,I55009,I54994,I48166,I48183,I55000,I48200,I48217,I48234,I48251,I48268,I55006,I48285,I55003,I48302,I48319,I48090,I48075,I48364,I48069,I48395,I48072,I48426,I48443,I48078,I48474,I48087,I48084,I48519,I48081,I48574,I48591,I62893,I62914,I48608,I62899,I48625,I62911,I48642,I62902,I48659,I62896,I48676,I48693,I48710,I48727,I48744,I62905,I62908,I48761,I48778,I48795,I48840,I48871,I48902,I48919,I48950,I48995,I49050,I49067,I49084,I49101,I49118,I49135,I49152,I49169,I49186,I49203,I49220,I49237,I49254,I49271,I49316,I49347,I49378,I49395,I49426,I49471,I49526,I49543,I49560,I49577,I49594,I49611,I49628,I49645,I49662,I49679,I49696,I49713,I49730,I49747,I49792,I49823,I49854,I49871,I49902,I49947,I50002,I50019,I76479,I76482,I50036,I50053,I76476,I76494,I50070,I50087,I76485,I50104,I50121,I50138,I50155,I50172,I76491,I76488,I50189,I50206,I50223,I49994,I49979,I50268,I49973,I50299,I49976,I50330,I50347,I49982,I50378,I49991,I49988,I50423,I49985,I50478,I50495,I50512,I50529,I50546,I50563,I50580,I50597,I50614,I50631,I50648,I50665,I50682,I50699,I50744,I50775,I50806,I50823,I50854,I50899,I50954,I50971,I50988,I51005,I51022,I51039,I51056,I51073,I51090,I51107,I51124,I51141,I51158,I51175,I51220,I51251,I51282,I51299,I51330,I51375,I51430,I51447,I52883,I52880,I51464,I52889,I51481,I52901,I52886,I51498,I51515,I52892,I51532,I51549,I51566,I51583,I51600,I52898,I51617,I52895,I51634,I51651,I51696,I51727,I51758,I51775,I51806,I51851,I51906,I51923,I51940,I51957,I51974,I51991,I52008,I52025,I52042,I52059,I52076,I52093,I52110,I52127,I52172,I52203,I52234,I52251,I52282,I52327,I52382,I52399,I52416,I52433,I52450,I52467,I52484,I52501,I52518,I52535,I52566,I52583,I52600,I52617,I52634,I52651,I52682,I52741,I52758,I52775,I52806,I52823,I52854,I52909,I52926,I52943,I52960,I52977,I52994,I53011,I53028,I53045,I53062,I53093,I53110,I53127,I53144,I53161,I53178,I53209,I53268,I53285,I53302,I53333,I53350,I53381,I53436,I53453,I53470,I53487,I53504,I53521,I53538,I53555,I53572,I53589,I53413,I53620,I53637,I53654,I53671,I53688,I53705,I53407,I53736,I53428,I53410,I53422,I53795,I53812,I53829,I53416,I53860,I53877,I53425,I53908,I53419,I53963,I53980,I60258,I60270,I53997,I60273,I60276,I54014,I54031,I54048,I54065,I60261,I54082,I60264,I54099,I54116,I54147,I54164,I54181,I54198,I60267,I54215,I60279,I54232,I54263,I54322,I54339,I54356,I54387,I54404,I54435,I54490,I54507,I54524,I54541,I54558,I54575,I54592,I54609,I54626,I54643,I54674,I54691,I54708,I54725,I54742,I54759,I54790,I54849,I54866,I54883,I54914,I54931,I54962,I55017,I55034,I55051,I55068,I55085,I55102,I55119,I55136,I55153,I55170,I55201,I55218,I55235,I55252,I55269,I55286,I55317,I55376,I55393,I55410,I55441,I55458,I55489,I55544,I55561,I55578,I55595,I55612,I55629,I55646,I55663,I55680,I55697,I55521,I55728,I55745,I55762,I55779,I55796,I55813,I55515,I55844,I55536,I55518,I55530,I55903,I55920,I55937,I55524,I55968,I55985,I55533,I56016,I55527,I56071,I56088,I56105,I56122,I56139,I56156,I56173,I56190,I56207,I56224,I56255,I56272,I56289,I56306,I56323,I56340,I56371,I56430,I56447,I56464,I56495,I56512,I56543,I56598,I56615,I56632,I56649,I56666,I56683,I56714,I56731,I56748,I56765,I56782,I56799,I56816,I56833,I56850,I56881,I56912,I56943,I56960,I57005,I57036,I57053,I57070,I57125,I57142,I57159,I57176,I57193,I57210,I57241,I57258,I57275,I57292,I57309,I57326,I57343,I57360,I57377,I57408,I57439,I57470,I57487,I57532,I57563,I57580,I57597,I57652,I57669,I57686,I57703,I57720,I57737,I57768,I57785,I57802,I57819,I57836,I57853,I57870,I57887,I57904,I57935,I57966,I57997,I58014,I58059,I58090,I58107,I58124,I58179,I58196,I69404,I69407,I58213,I69419,I58230,I69410,I58247,I58264,I58295,I58312,I69413,I58329,I58346,I69416,I58363,I58380,I58397,I69422,I58414,I58431,I58462,I58493,I58524,I58541,I58586,I58617,I58634,I58651,I58706,I58723,I58740,I58757,I58774,I58791,I58822,I58839,I58856,I58873,I58890,I58907,I58924,I58941,I58958,I58989,I59020,I59051,I59068,I59113,I59144,I59161,I59178,I59233,I59250,I59267,I59284,I59301,I59318,I59349,I59366,I59383,I59400,I59417,I59434,I59451,I59468,I59485,I59516,I59547,I59578,I59595,I59640,I59671,I59688,I59705,I59760,I59777,I59794,I59811,I59828,I59845,I59876,I59893,I59910,I59927,I59944,I59961,I59978,I59995,I60012,I60043,I60074,I60105,I60122,I60167,I60198,I60215,I60232,I60287,I60304,I75150,I75153,I60321,I75165,I60338,I75156,I60355,I60372,I60403,I60420,I75159,I60437,I60454,I75162,I60471,I60488,I60505,I75168,I60522,I60539,I60570,I60601,I60632,I60649,I60694,I60725,I60742,I60759,I60814,I60831,I60848,I60865,I60882,I60899,I60930,I60947,I60964,I60981,I60998,I61015,I61032,I61049,I61066,I61097,I61128,I61159,I61176,I61221,I61252,I61269,I61286,I61341,I61358,I73824,I73827,I61375,I73839,I61392,I73830,I61409,I61426,I61457,I61474,I73833,I61491,I61508,I73836,I61525,I61542,I61559,I73842,I61576,I61593,I61624,I61655,I61686,I61703,I61748,I61779,I61796,I61813,I61868,I61885,I68520,I68523,I61902,I68535,I61919,I68526,I61936,I61953,I61984,I62001,I68529,I62018,I62035,I68532,I62052,I62069,I62086,I68538,I62103,I62120,I62151,I62182,I62213,I62230,I62275,I62306,I62323,I62340,I62395,I62412,I62429,I62446,I62463,I62480,I62511,I62528,I62545,I62562,I62579,I62596,I62613,I62630,I62647,I62678,I62709,I62740,I62757,I62802,I62833,I62850,I62867,I62922,I62939,I62956,I62973,I62990,I63007,I63038,I63055,I63072,I63089,I63106,I63123,I63140,I63157,I63174,I63205,I63236,I63267,I63284,I63329,I63360,I63377,I63394,I63449,I63466,I63483,I63500,I63517,I63534,I63423,I63565,I63582,I63599,I63616,I63633,I63650,I63667,I63684,I63701,I63420,I63732,I63435,I63763,I63432,I63794,I63811,I63438,I63441,I63856,I63426,I63887,I63904,I63921,I63429,I63976,I63993,I64010,I64027,I64044,I64061,I64092,I64109,I64126,I64143,I64160,I64177,I64194,I64211,I64228,I64259,I64290,I64321,I64338,I64383,I64414,I64431,I64448,I64503,I64520,I64537,I64554,I64571,I64588,I64477,I64619,I64636,I64653,I64670,I64687,I64704,I64721,I64738,I64755,I64474,I64786,I64489,I64817,I64486,I64848,I64865,I64492,I64495,I64910,I64480,I64941,I64958,I64975,I64483,I65030,I65047,I65064,I65081,I65098,I65115,I65146,I65163,I65180,I65197,I65214,I65231,I65248,I65265,I65282,I65313,I65344,I65375,I65392,I65437,I65468,I65485,I65502,I65557,I65574,I65591,I65608,I65625,I65642,I65531,I65673,I65690,I65707,I65724,I65741,I65758,I65775,I65792,I65809,I65528,I65840,I65543,I65871,I65540,I65902,I65919,I65546,I65549,I65964,I65534,I65995,I66012,I66029,I65537,I66084,I66101,I66118,I66135,I66152,I66169,I66200,I66217,I66234,I66251,I66268,I66285,I66302,I66319,I66336,I66367,I66398,I66429,I66446,I66491,I66522,I66539,I66556,I66611,I66628,I66645,I66662,I66679,I66696,I66727,I66744,I66761,I66778,I66795,I66812,I66829,I66846,I66863,I66894,I66925,I66956,I66973,I67018,I67049,I67066,I67083,I67138,I67155,I67172,I67189,I67206,I67223,I67254,I67271,I67288,I67305,I67322,I67339,I67356,I67373,I67390,I67421,I67452,I67483,I67500,I67545,I67576,I67593,I67610,I67662,I67679,I67696,I67713,I67730,I67761,I67778,I67795,I67812,I67829,I67846,I67863,I67880,I67939,I67956,I67973,I68004,I68021,I68052,I68104,I68121,I68138,I68155,I68172,I68203,I68220,I68237,I68254,I68271,I68288,I68305,I68322,I68381,I68398,I68415,I68446,I68463,I68494,I68546,I68563,I68580,I68597,I68614,I68645,I68662,I68679,I68696,I68713,I68730,I68747,I68764,I68823,I68840,I68857,I68888,I68905,I68936,I68988,I69005,I69022,I69039,I69056,I69087,I69104,I69121,I69138,I69155,I69172,I69189,I69206,I69265,I69282,I69299,I69330,I69347,I69378,I69430,I69447,I69464,I69481,I69498,I69529,I69546,I69563,I69580,I69597,I69614,I69631,I69648,I69707,I69724,I69741,I69772,I69789,I69820,I69872,I69889,I69906,I69923,I69940,I69971,I69988,I70005,I70022,I70039,I70056,I70073,I70090,I70149,I70166,I70183,I70214,I70231,I70262,I70314,I70331,I70348,I70365,I70382,I70413,I70430,I70447,I70464,I70481,I70498,I70515,I70532,I70591,I70608,I70625,I70656,I70673,I70704,I70756,I70773,I70790,I70807,I70824,I70855,I70872,I70889,I70906,I70923,I70940,I70957,I70974,I71033,I71050,I71067,I71098,I71115,I71146,I71198,I71215,I71232,I71249,I71266,I71297,I71314,I71331,I71348,I71365,I71382,I71399,I71416,I71475,I71492,I71509,I71540,I71557,I71588,I71640,I71657,I71674,I71691,I71708,I71739,I71756,I71773,I71790,I71807,I71824,I71841,I71858,I71917,I71934,I71951,I71982,I71999,I72030,I72082,I72099,I72116,I72133,I72150,I72181,I72198,I72215,I72232,I72249,I72266,I72283,I72300,I72359,I72376,I72393,I72424,I72441,I72472,I72524,I72541,I72558,I72575,I72592,I72623,I72640,I72657,I72674,I72691,I72708,I72725,I72742,I72801,I72818,I72835,I72866,I72883,I72914,I72966,I72983,I73000,I73017,I73034,I73065,I73082,I73099,I73116,I73133,I73150,I73167,I73184,I73243,I73260,I73277,I73308,I73325,I73356,I73408,I73425,I73442,I73459,I73476,I73507,I73524,I73541,I73558,I73575,I73592,I73609,I73626,I73685,I73702,I73719,I73750,I73767,I73798,I73850,I73867,I73884,I73901,I73918,I73949,I73966,I73983,I74000,I74017,I74034,I74051,I74068,I74127,I74144,I74161,I74192,I74209,I74240,I74292,I74309,I74326,I74343,I74360,I74391,I74408,I74425,I74442,I74459,I74476,I74493,I74510,I74569,I74586,I74603,I74634,I74651,I74682,I74734,I74751,I74768,I74785,I74802,I74833,I74850,I74867,I74884,I74901,I74918,I74935,I74952,I75011,I75028,I75045,I75076,I75093,I75124,I75176,I75193,I75210,I75227,I75244,I75275,I75292,I75309,I75326,I75343,I75360,I75377,I75394,I75453,I75470,I75487,I75518,I75535,I75566,I75618,I75635,I75652,I75669,I75686,I75717,I75734,I75751,I75768,I75785,I75802,I75819,I75836,I75895,I75912,I75929,I75960,I75977,I76008,I76060,I76077,I76094,I76111,I76128,I76159,I76176,I76193,I76210,I76227,I76244,I76261,I76278,I76337,I76354,I76371,I76402,I76419,I76450,I76502,I76519,I76536,I76553,I76570,I76601,I76618,I76635,I76652,I76669,I76686,I76703,I76720,I76779,I76796,I76813,I76844,I76861,I76892,I76944,I76961,I76978,I76995,I77012,I77043,I77060,I77077,I77094,I77111,I77128,I77145,I77162,I77221,I77238,I77255,I77286,I77303,I77334,I77386,I77403,I77420,I77437,I77454,I77485,I77502,I77519,I77536,I77553,I77570,I77587,I77604,I77663,I77680,I77697,I77728,I77745,I77776;
not I_0 (I1637,I1605);
or I_1 (I1654,I21153,I21156);
nand I_2 (I1671,I21141,I21150);
not I_3 (I1688,I1671);
and I_4 (I1705,I1688,I1654);
DFFARX1 I_5 (I1688,I1598,I1637,I1617,);
nand I_6 (I1736,I21141,I21159);
and I_7 (I1753,I1736,I21150);
DFFARX1 I_8 (I1753,I1598,I1637,I1779,);
nor I_9 (I1787,I1779,I1705);
not I_10 (I1804,I1779);
nor I_11 (I1821,I21144,I21159);
not I_12 (I1838,I1821);
nand I_13 (I1855,I1804,I1838);
nand I_14 (I1872,I1821,I1671);
nand I_15 (I1889,I1804,I1872);
nand I_16 (I1623,I1787,I1821);
not I_17 (I1920,I21144);
nand I_18 (I1937,I1855,I1920);
nand I_19 (I1954,I21147,I21147);
nor I_20 (I1608,I1705,I1954);
not I_21 (I1985,I1954);
nand I_22 (I2002,I1985,I1920);
nor I_23 (I2019,I1838,I2002);
nor I_24 (I1626,I1804,I2019);
nor I_25 (I1629,I1954,I1937);
nor I_26 (I2064,I1954,I21144);
nor I_27 (I1611,I2064,I1889);
nand I_28 (I1614,I1688,I1954);
nor I_29 (I2109,I1779,I1954);
nand I_30 (I1620,I2109,I1705);
not I_31 (I2164,I1605);
or I_32 (I2181,I51419,I51401);
nand I_33 (I2198,I51407,I51422);
not I_34 (I2215,I2198);
and I_35 (I2232,I2215,I2181);
DFFARX1 I_36 (I2215,I1598,I2164,I2144,);
nand I_37 (I2263,I51404,I51410);
and I_38 (I2280,I2263,I51407);
DFFARX1 I_39 (I2280,I1598,I2164,I2306,);
nor I_40 (I2314,I2306,I2232);
not I_41 (I2331,I2306);
nor I_42 (I2348,I51413,I51410);
not I_43 (I2365,I2348);
nand I_44 (I2382,I2331,I2365);
nand I_45 (I2399,I2348,I2198);
nand I_46 (I2416,I2331,I2399);
nand I_47 (I2150,I2314,I2348);
not I_48 (I2447,I51404);
nand I_49 (I2464,I2382,I2447);
nand I_50 (I2481,I51416,I51401);
nor I_51 (I2135,I2232,I2481);
not I_52 (I2512,I2481);
nand I_53 (I2529,I2512,I2447);
nor I_54 (I2546,I2365,I2529);
nor I_55 (I2153,I2331,I2546);
nor I_56 (I2156,I2481,I2464);
nor I_57 (I2591,I2481,I51404);
nor I_58 (I2138,I2591,I2416);
nand I_59 (I2141,I2215,I2481);
nor I_60 (I2636,I2306,I2481);
nand I_61 (I2147,I2636,I2232);
not I_62 (I2691,I1605);
or I_63 (I2708,I1231,I823);
nand I_64 (I2725,I1327,I647);
not I_65 (I2742,I2725);
and I_66 (I2759,I2742,I2708);
DFFARX1 I_67 (I2742,I1598,I2691,I2671,);
nand I_68 (I2790,I863,I1575);
and I_69 (I2807,I2790,I799);
DFFARX1 I_70 (I2807,I1598,I2691,I2833,);
nor I_71 (I2841,I2833,I2759);
not I_72 (I2858,I2833);
nor I_73 (I2875,I1079,I1575);
not I_74 (I2892,I2875);
nand I_75 (I2909,I2858,I2892);
nand I_76 (I2926,I2875,I2725);
nand I_77 (I2943,I2858,I2926);
nand I_78 (I2677,I2841,I2875);
not I_79 (I2974,I639);
nand I_80 (I2991,I2909,I2974);
nand I_81 (I3008,I783,I943);
nor I_82 (I2662,I2759,I3008);
not I_83 (I3039,I3008);
nand I_84 (I3056,I3039,I2974);
nor I_85 (I3073,I2892,I3056);
nor I_86 (I2680,I2858,I3073);
nor I_87 (I2683,I3008,I2991);
nor I_88 (I3118,I3008,I639);
nor I_89 (I2665,I3118,I2943);
nand I_90 (I2668,I2742,I3008);
nor I_91 (I3163,I2833,I3008);
nand I_92 (I2674,I3163,I2759);
not I_93 (I3218,I1605);
or I_94 (I3235,I7884,I7884);
nand I_95 (I3252,I7905,I7902);
not I_96 (I3269,I3252);
and I_97 (I3286,I3269,I3235);
DFFARX1 I_98 (I3269,I1598,I3218,I3198,);
nand I_99 (I3317,I7881,I7893);
and I_100 (I3334,I3317,I7890);
DFFARX1 I_101 (I3334,I1598,I3218,I3360,);
nor I_102 (I3368,I3360,I3286);
not I_103 (I3385,I3360);
nor I_104 (I3402,I7899,I7893);
not I_105 (I3419,I3402);
nand I_106 (I3436,I3385,I3419);
nand I_107 (I3453,I3402,I3252);
nand I_108 (I3470,I3385,I3453);
nand I_109 (I3204,I3368,I3402);
not I_110 (I3501,I7881);
nand I_111 (I3518,I3436,I3501);
nand I_112 (I3535,I7896,I7887);
nor I_113 (I3189,I3286,I3535);
not I_114 (I3566,I3535);
nand I_115 (I3583,I3566,I3501);
nor I_116 (I3600,I3419,I3583);
nor I_117 (I3207,I3385,I3600);
nor I_118 (I3210,I3535,I3518);
nor I_119 (I3645,I3535,I7881);
nor I_120 (I3192,I3645,I3470);
nand I_121 (I3195,I3269,I3535);
nor I_122 (I3690,I3360,I3535);
nand I_123 (I3201,I3690,I3286);
not I_124 (I3745,I1605);
or I_125 (I3762,I48563,I48545);
nand I_126 (I3779,I48551,I48566);
not I_127 (I3796,I3779);
and I_128 (I3813,I3796,I3762);
DFFARX1 I_129 (I3796,I1598,I3745,I3725,);
nand I_130 (I3844,I48548,I48554);
and I_131 (I3861,I3844,I48551);
DFFARX1 I_132 (I3861,I1598,I3745,I3887,);
nor I_133 (I3895,I3887,I3813);
not I_134 (I3912,I3887);
nor I_135 (I3929,I48557,I48554);
not I_136 (I3946,I3929);
nand I_137 (I3963,I3912,I3946);
nand I_138 (I3980,I3929,I3779);
nand I_139 (I3997,I3912,I3980);
nand I_140 (I3731,I3895,I3929);
not I_141 (I4028,I48548);
nand I_142 (I4045,I3963,I4028);
nand I_143 (I4062,I48560,I48545);
nor I_144 (I3716,I3813,I4062);
not I_145 (I4093,I4062);
nand I_146 (I4110,I4093,I4028);
nor I_147 (I4127,I3946,I4110);
nor I_148 (I3734,I3912,I4127);
nor I_149 (I3737,I4062,I4045);
nor I_150 (I4172,I4062,I48548);
nor I_151 (I3719,I4172,I3997);
nand I_152 (I3722,I3796,I4062);
nor I_153 (I4217,I3887,I4062);
nand I_154 (I3728,I4217,I3813);
not I_155 (I4272,I1605);
or I_156 (I4289,I13494,I13494);
nand I_157 (I4306,I13515,I13512);
not I_158 (I4323,I4306);
and I_159 (I4340,I4323,I4289);
DFFARX1 I_160 (I4323,I1598,I4272,I4252,);
nand I_161 (I4371,I13491,I13503);
and I_162 (I4388,I4371,I13500);
DFFARX1 I_163 (I4388,I1598,I4272,I4414,);
nor I_164 (I4422,I4414,I4340);
not I_165 (I4439,I4414);
nor I_166 (I4456,I13509,I13503);
not I_167 (I4473,I4456);
nand I_168 (I4490,I4439,I4473);
nand I_169 (I4507,I4456,I4306);
nand I_170 (I4524,I4439,I4507);
nand I_171 (I4258,I4422,I4456);
not I_172 (I4555,I13491);
nand I_173 (I4572,I4490,I4555);
nand I_174 (I4589,I13506,I13497);
nor I_175 (I4243,I4340,I4589);
not I_176 (I4620,I4589);
nand I_177 (I4637,I4620,I4555);
nor I_178 (I4654,I4473,I4637);
nor I_179 (I4261,I4439,I4654);
nor I_180 (I4264,I4589,I4572);
nor I_181 (I4699,I4589,I13491);
nor I_182 (I4246,I4699,I4524);
nand I_183 (I4249,I4323,I4589);
nor I_184 (I4744,I4414,I4589);
nand I_185 (I4255,I4744,I4340);
not I_186 (I4799,I1605);
or I_187 (I4816,I38567,I38549);
nand I_188 (I4833,I38555,I38570);
not I_189 (I4850,I4833);
and I_190 (I4867,I4850,I4816);
DFFARX1 I_191 (I4850,I1598,I4799,I4779,);
nand I_192 (I4898,I38552,I38558);
and I_193 (I4915,I4898,I38555);
DFFARX1 I_194 (I4915,I1598,I4799,I4941,);
nor I_195 (I4949,I4941,I4867);
not I_196 (I4966,I4941);
nor I_197 (I4983,I38561,I38558);
not I_198 (I5000,I4983);
nand I_199 (I5017,I4966,I5000);
nand I_200 (I5034,I4983,I4833);
nand I_201 (I5051,I4966,I5034);
nand I_202 (I4785,I4949,I4983);
not I_203 (I5082,I38552);
nand I_204 (I5099,I5017,I5082);
nand I_205 (I5116,I38564,I38549);
nor I_206 (I4770,I4867,I5116);
not I_207 (I5147,I5116);
nand I_208 (I5164,I5147,I5082);
nor I_209 (I5181,I5000,I5164);
nor I_210 (I4788,I4966,I5181);
nor I_211 (I4791,I5116,I5099);
nor I_212 (I5226,I5116,I38552);
nor I_213 (I4773,I5226,I5051);
nand I_214 (I4776,I4850,I5116);
nor I_215 (I5271,I4941,I5116);
nand I_216 (I4782,I5271,I4867);
not I_217 (I5326,I1605);
or I_218 (I5343,I8904,I8904);
nand I_219 (I5360,I8925,I8922);
not I_220 (I5377,I5360);
and I_221 (I5394,I5377,I5343);
DFFARX1 I_222 (I5377,I1598,I5326,I5306,);
nand I_223 (I5425,I8901,I8913);
and I_224 (I5442,I5425,I8910);
DFFARX1 I_225 (I5442,I1598,I5326,I5468,);
nor I_226 (I5476,I5468,I5394);
not I_227 (I5493,I5468);
nor I_228 (I5510,I8919,I8913);
not I_229 (I5527,I5510);
nand I_230 (I5544,I5493,I5527);
nand I_231 (I5561,I5510,I5360);
nand I_232 (I5578,I5493,I5561);
nand I_233 (I5312,I5476,I5510);
not I_234 (I5609,I8901);
nand I_235 (I5626,I5544,I5609);
nand I_236 (I5643,I8916,I8907);
nor I_237 (I5297,I5394,I5643);
not I_238 (I5674,I5643);
nand I_239 (I5691,I5674,I5609);
nor I_240 (I5708,I5527,I5691);
nor I_241 (I5315,I5493,I5708);
nor I_242 (I5318,I5643,I5626);
nor I_243 (I5753,I5643,I8901);
nor I_244 (I5300,I5753,I5578);
nand I_245 (I5303,I5377,I5643);
nor I_246 (I5798,I5468,I5643);
nand I_247 (I5309,I5798,I5394);
not I_248 (I5853,I1605);
or I_249 (I5870,I67648,I67642);
nand I_250 (I5887,I67639,I67639);
not I_251 (I5904,I5887);
and I_252 (I5921,I5904,I5870);
DFFARX1 I_253 (I5904,I1598,I5853,I5833,);
nand I_254 (I5952,I67645,I67651);
and I_255 (I5969,I5952,I67645);
DFFARX1 I_256 (I5969,I1598,I5853,I5995,);
nor I_257 (I6003,I5995,I5921);
not I_258 (I6020,I5995);
nor I_259 (I6037,I67636,I67651);
not I_260 (I6054,I6037);
nand I_261 (I6071,I6020,I6054);
nand I_262 (I6088,I6037,I5887);
nand I_263 (I6105,I6020,I6088);
nand I_264 (I5839,I6003,I6037);
not I_265 (I6136,I67636);
nand I_266 (I6153,I6071,I6136);
nand I_267 (I6170,I67654,I67642);
nor I_268 (I5824,I5921,I6170);
not I_269 (I6201,I6170);
nand I_270 (I6218,I6201,I6136);
nor I_271 (I6235,I6054,I6218);
nor I_272 (I5842,I6020,I6235);
nor I_273 (I5845,I6170,I6153);
nor I_274 (I6280,I6170,I67636);
nor I_275 (I5827,I6280,I6105);
nand I_276 (I5830,I5904,I6170);
nor I_277 (I6325,I5995,I6170);
nand I_278 (I5836,I6325,I5921);
not I_279 (I6383,I1605);
or I_280 (I6400,I70288,I70288);
nand I_281 (I6417,I70303,I70306);
not I_282 (I6434,I6417);
nand I_283 (I6451,I6434,I6400);
not I_284 (I6468,I6451);
nand I_285 (I6485,I70294,I70297);
and I_286 (I6502,I6485,I70291);
DFFARX1 I_287 (I6502,I1598,I6383,I6528,);
not I_288 (I6536,I6528);
nor I_289 (I6553,I70297,I70297);
nor I_290 (I6570,I6528,I6553);
and I_291 (I6587,I6528,I6553);
nor I_292 (I6604,I6587,I6451);
DFFARX1 I_293 (I6604,I1598,I6383,I6363,);
nand I_294 (I6635,I70300,I70294);
nor I_295 (I6652,I6635,I70291);
nand I_296 (I6669,I6468,I6652);
not I_297 (I6372,I6669);
nor I_298 (I6375,I6570,I6669);
nor I_299 (I6714,I6652,I6434);
nor I_300 (I6366,I6536,I6714);
nor I_301 (I6360,I6652,I6553);
not I_302 (I6759,I6635);
nand I_303 (I6776,I6553,I6759);
not I_304 (I6354,I6776);
nor I_305 (I6357,I6417,I6776);
nor I_306 (I6369,I6759,I6417);
nand I_307 (I6835,I6536,I6635);
nor I_308 (I6351,I6434,I6835);
not I_309 (I6893,I1605);
or I_310 (I6910,I69846,I69846);
nand I_311 (I6927,I69861,I69864);
not I_312 (I6944,I6927);
nand I_313 (I6961,I6944,I6910);
not I_314 (I6978,I6961);
nand I_315 (I6995,I69852,I69855);
and I_316 (I7012,I6995,I69849);
DFFARX1 I_317 (I7012,I1598,I6893,I7038,);
not I_318 (I7046,I7038);
nor I_319 (I7063,I69855,I69855);
nor I_320 (I7080,I7038,I7063);
and I_321 (I7097,I7038,I7063);
nor I_322 (I7114,I7097,I6961);
DFFARX1 I_323 (I7114,I1598,I6893,I6873,);
nand I_324 (I7145,I69858,I69852);
nor I_325 (I7162,I7145,I69849);
nand I_326 (I7179,I6978,I7162);
not I_327 (I6882,I7179);
nor I_328 (I6885,I7080,I7179);
nor I_329 (I7224,I7162,I6944);
nor I_330 (I6876,I7046,I7224);
nor I_331 (I6870,I7162,I7063);
not I_332 (I7269,I7145);
nand I_333 (I7286,I7063,I7269);
not I_334 (I6864,I7286);
nor I_335 (I6867,I6927,I7286);
nor I_336 (I6879,I7269,I6927);
nand I_337 (I7345,I7046,I7145);
nor I_338 (I6861,I6944,I7345);
not I_339 (I7403,I1605);
or I_340 (I7420,I63953,I63947);
nand I_341 (I7437,I63956,I63959);
not I_342 (I7454,I7437);
nand I_343 (I7471,I7454,I7420);
not I_344 (I7488,I7471);
nand I_345 (I7505,I63950,I63953);
and I_346 (I7522,I7505,I63947);
DFFARX1 I_347 (I7522,I1598,I7403,I7548,);
not I_348 (I7556,I7548);
nor I_349 (I7573,I63965,I63953);
nor I_350 (I7590,I7548,I7573);
and I_351 (I7607,I7548,I7573);
nor I_352 (I7624,I7607,I7471);
DFFARX1 I_353 (I7624,I1598,I7403,I7383,);
nand I_354 (I7655,I63962,I63950);
nor I_355 (I7672,I7655,I63968);
nand I_356 (I7689,I7488,I7672);
not I_357 (I7392,I7689);
nor I_358 (I7395,I7590,I7689);
nor I_359 (I7734,I7672,I7454);
nor I_360 (I7386,I7556,I7734);
nor I_361 (I7380,I7672,I7573);
not I_362 (I7779,I7655);
nand I_363 (I7796,I7573,I7779);
not I_364 (I7374,I7796);
nor I_365 (I7377,I7437,I7796);
nor I_366 (I7389,I7779,I7437);
nand I_367 (I7855,I7556,I7655);
nor I_368 (I7371,I7454,I7855);
not I_369 (I7913,I1605);
or I_370 (I7930,I74266,I74266);
nand I_371 (I7947,I74281,I74284);
not I_372 (I7964,I7947);
nand I_373 (I7981,I7964,I7930);
not I_374 (I7998,I7981);
nand I_375 (I8015,I74272,I74275);
and I_376 (I8032,I8015,I74269);
DFFARX1 I_377 (I8032,I1598,I7913,I8058,);
not I_378 (I8066,I8058);
nor I_379 (I8083,I74275,I74275);
nor I_380 (I8100,I8058,I8083);
and I_381 (I8117,I8058,I8083);
nor I_382 (I8134,I8117,I7981);
DFFARX1 I_383 (I8134,I1598,I7913,I7893,);
nand I_384 (I8165,I74278,I74272);
nor I_385 (I8182,I8165,I74269);
nand I_386 (I8199,I7998,I8182);
not I_387 (I7902,I8199);
nor I_388 (I7905,I8100,I8199);
nor I_389 (I8244,I8182,I7964);
nor I_390 (I7896,I8066,I8244);
nor I_391 (I7890,I8182,I8083);
not I_392 (I8289,I8165);
nand I_393 (I8306,I8083,I8289);
not I_394 (I7884,I8306);
nor I_395 (I7887,I7947,I8306);
nor I_396 (I7899,I8289,I7947);
nand I_397 (I8365,I8066,I8165);
nor I_398 (I7881,I7964,I8365);
not I_399 (I8423,I1605);
or I_400 (I8440,I61318,I61312);
nand I_401 (I8457,I61321,I61324);
not I_402 (I8474,I8457);
nand I_403 (I8491,I8474,I8440);
not I_404 (I8508,I8491);
nand I_405 (I8525,I61315,I61318);
and I_406 (I8542,I8525,I61312);
DFFARX1 I_407 (I8542,I1598,I8423,I8568,);
not I_408 (I8576,I8568);
nor I_409 (I8593,I61330,I61318);
nor I_410 (I8610,I8568,I8593);
and I_411 (I8627,I8568,I8593);
nor I_412 (I8644,I8627,I8491);
DFFARX1 I_413 (I8644,I1598,I8423,I8403,);
nand I_414 (I8675,I61327,I61315);
nor I_415 (I8692,I8675,I61333);
nand I_416 (I8709,I8508,I8692);
not I_417 (I8412,I8709);
nor I_418 (I8415,I8610,I8709);
nor I_419 (I8754,I8692,I8474);
nor I_420 (I8406,I8576,I8754);
nor I_421 (I8400,I8692,I8593);
not I_422 (I8799,I8675);
nand I_423 (I8816,I8593,I8799);
not I_424 (I8394,I8816);
nor I_425 (I8397,I8457,I8816);
nor I_426 (I8409,I8799,I8457);
nand I_427 (I8875,I8576,I8675);
nor I_428 (I8391,I8474,I8875);
not I_429 (I8933,I1605);
or I_430 (I8950,I21963,I21957);
nand I_431 (I8967,I21963,I21975);
not I_432 (I8984,I8967);
nand I_433 (I9001,I8984,I8950);
not I_434 (I9018,I9001);
nand I_435 (I9035,I21969,I21960);
and I_436 (I9052,I9035,I21957);
DFFARX1 I_437 (I9052,I1598,I8933,I9078,);
not I_438 (I9086,I9078);
nor I_439 (I9103,I21972,I21960);
nor I_440 (I9120,I9078,I9103);
and I_441 (I9137,I9078,I9103);
nor I_442 (I9154,I9137,I9001);
DFFARX1 I_443 (I9154,I1598,I8933,I8913,);
nand I_444 (I9185,I21966,I21966);
nor I_445 (I9202,I9185,I21960);
nand I_446 (I9219,I9018,I9202);
not I_447 (I8922,I9219);
nor I_448 (I8925,I9120,I9219);
nor I_449 (I9264,I9202,I8984);
nor I_450 (I8916,I9086,I9264);
nor I_451 (I8910,I9202,I9103);
not I_452 (I9309,I9185);
nand I_453 (I9326,I9103,I9309);
not I_454 (I8904,I9326);
nor I_455 (I8907,I8967,I9326);
nor I_456 (I8919,I9309,I8967);
nand I_457 (I9385,I9086,I9185);
nor I_458 (I8901,I8984,I9385);
not I_459 (I9443,I1605);
or I_460 (I9460,I25602,I25581);
nand I_461 (I9477,I25590,I25599);
not I_462 (I9494,I9477);
nand I_463 (I9511,I9494,I9460);
not I_464 (I9528,I9511);
nand I_465 (I9545,I25596,I25581);
and I_466 (I9562,I9545,I25587);
DFFARX1 I_467 (I9562,I1598,I9443,I9588,);
not I_468 (I9596,I9588);
nor I_469 (I9613,I25578,I25581);
nor I_470 (I9630,I9588,I9613);
and I_471 (I9647,I9588,I9613);
nor I_472 (I9664,I9647,I9511);
DFFARX1 I_473 (I9664,I1598,I9443,I9423,);
nand I_474 (I9695,I25593,I25578);
nor I_475 (I9712,I9695,I25584);
nand I_476 (I9729,I9528,I9712);
not I_477 (I9432,I9729);
nor I_478 (I9435,I9630,I9729);
nor I_479 (I9774,I9712,I9494);
nor I_480 (I9426,I9596,I9774);
nor I_481 (I9420,I9712,I9613);
not I_482 (I9819,I9695);
nand I_483 (I9836,I9613,I9819);
not I_484 (I9414,I9836);
nor I_485 (I9417,I9477,I9836);
nor I_486 (I9429,I9819,I9477);
nand I_487 (I9895,I9596,I9695);
nor I_488 (I9411,I9494,I9895);
not I_489 (I9953,I1605);
or I_490 (I9970,I35088,I35067);
nand I_491 (I9987,I35076,I35085);
not I_492 (I10004,I9987);
nand I_493 (I10021,I10004,I9970);
not I_494 (I10038,I10021);
nand I_495 (I10055,I35082,I35067);
and I_496 (I10072,I10055,I35073);
DFFARX1 I_497 (I10072,I1598,I9953,I10098,);
not I_498 (I10106,I10098);
nor I_499 (I10123,I35064,I35067);
nor I_500 (I10140,I10098,I10123);
and I_501 (I10157,I10098,I10123);
nor I_502 (I10174,I10157,I10021);
DFFARX1 I_503 (I10174,I1598,I9953,I9933,);
nand I_504 (I10205,I35079,I35064);
nor I_505 (I10222,I10205,I35070);
nand I_506 (I10239,I10038,I10222);
not I_507 (I9942,I10239);
nor I_508 (I9945,I10140,I10239);
nor I_509 (I10284,I10222,I10004);
nor I_510 (I9936,I10106,I10284);
nor I_511 (I9930,I10222,I10123);
not I_512 (I10329,I10205);
nand I_513 (I10346,I10123,I10329);
not I_514 (I9924,I10346);
nor I_515 (I9927,I9987,I10346);
nor I_516 (I9939,I10329,I9987);
nand I_517 (I10405,I10106,I10205);
nor I_518 (I9921,I10004,I10405);
not I_519 (I10463,I1605);
or I_520 (I10480,I3189,I3189);
nand I_521 (I10497,I3192,I3195);
not I_522 (I10514,I10497);
nand I_523 (I10531,I10514,I10480);
not I_524 (I10548,I10531);
nand I_525 (I10565,I3204,I3210);
and I_526 (I10582,I10565,I3198);
DFFARX1 I_527 (I10582,I1598,I10463,I10608,);
not I_528 (I10616,I10608);
nor I_529 (I10633,I3195,I3210);
nor I_530 (I10650,I10608,I10633);
and I_531 (I10667,I10608,I10633);
nor I_532 (I10684,I10667,I10531);
DFFARX1 I_533 (I10684,I1598,I10463,I10443,);
nand I_534 (I10715,I3192,I3201);
nor I_535 (I10732,I10715,I3207);
nand I_536 (I10749,I10548,I10732);
not I_537 (I10452,I10749);
nor I_538 (I10455,I10650,I10749);
nor I_539 (I10794,I10732,I10514);
nor I_540 (I10446,I10616,I10794);
nor I_541 (I10440,I10732,I10633);
not I_542 (I10839,I10715);
nand I_543 (I10856,I10633,I10839);
not I_544 (I10434,I10856);
nor I_545 (I10437,I10497,I10856);
nor I_546 (I10449,I10839,I10497);
nand I_547 (I10915,I10616,I10715);
nor I_548 (I10431,I10514,I10915);
not I_549 (I10973,I1605);
or I_550 (I10990,I1567,I1295);
nand I_551 (I11007,I991,I671);
not I_552 (I11024,I11007);
nand I_553 (I11041,I11024,I10990);
not I_554 (I11058,I11041);
nand I_555 (I11075,I751,I1175);
and I_556 (I11092,I11075,I831);
DFFARX1 I_557 (I11092,I1598,I10973,I11118,);
not I_558 (I11126,I11118);
nor I_559 (I11143,I1391,I1175);
nor I_560 (I11160,I11118,I11143);
and I_561 (I11177,I11118,I11143);
nor I_562 (I11194,I11177,I11041);
DFFARX1 I_563 (I11194,I1598,I10973,I10953,);
nand I_564 (I11225,I663,I967);
nor I_565 (I11242,I11225,I1263);
nand I_566 (I11259,I11058,I11242);
not I_567 (I10962,I11259);
nor I_568 (I10965,I11160,I11259);
nor I_569 (I11304,I11242,I11024);
nor I_570 (I10956,I11126,I11304);
nor I_571 (I10950,I11242,I11143);
not I_572 (I11349,I11225);
nand I_573 (I11366,I11143,I11349);
not I_574 (I10944,I11366);
nor I_575 (I10947,I11007,I11366);
nor I_576 (I10959,I11349,I11007);
nand I_577 (I11425,I11126,I11225);
nor I_578 (I10941,I11024,I11425);
not I_579 (I11483,I1605);
or I_580 (I11500,I31399,I31378);
nand I_581 (I11517,I31387,I31396);
not I_582 (I11534,I11517);
nand I_583 (I11551,I11534,I11500);
not I_584 (I11568,I11551);
nand I_585 (I11585,I31393,I31378);
and I_586 (I11602,I11585,I31384);
DFFARX1 I_587 (I11602,I1598,I11483,I11628,);
not I_588 (I11636,I11628);
nor I_589 (I11653,I31375,I31378);
nor I_590 (I11670,I11628,I11653);
and I_591 (I11687,I11628,I11653);
nor I_592 (I11704,I11687,I11551);
DFFARX1 I_593 (I11704,I1598,I11483,I11463,);
nand I_594 (I11735,I31390,I31375);
nor I_595 (I11752,I11735,I31381);
nand I_596 (I11769,I11568,I11752);
not I_597 (I11472,I11769);
nor I_598 (I11475,I11670,I11769);
nor I_599 (I11814,I11752,I11534);
nor I_600 (I11466,I11636,I11814);
nor I_601 (I11460,I11752,I11653);
not I_602 (I11859,I11735);
nand I_603 (I11876,I11653,I11859);
not I_604 (I11454,I11876);
nor I_605 (I11457,I11517,I11876);
nor I_606 (I11469,I11859,I11517);
nand I_607 (I11935,I11636,I11735);
nor I_608 (I11451,I11534,I11935);
not I_609 (I11993,I1605);
or I_610 (I12010,I72498,I72498);
nand I_611 (I12027,I72513,I72516);
not I_612 (I12044,I12027);
nand I_613 (I12061,I12044,I12010);
not I_614 (I12078,I12061);
nand I_615 (I12095,I72504,I72507);
and I_616 (I12112,I12095,I72501);
DFFARX1 I_617 (I12112,I1598,I11993,I12138,);
not I_618 (I12146,I12138);
nor I_619 (I12163,I72507,I72507);
nor I_620 (I12180,I12138,I12163);
and I_621 (I12197,I12138,I12163);
nor I_622 (I12214,I12197,I12061);
DFFARX1 I_623 (I12214,I1598,I11993,I11973,);
nand I_624 (I12245,I72510,I72504);
nor I_625 (I12262,I12245,I72501);
nand I_626 (I12279,I12078,I12262);
not I_627 (I11982,I12279);
nor I_628 (I11985,I12180,I12279);
nor I_629 (I12324,I12262,I12044);
nor I_630 (I11976,I12146,I12324);
nor I_631 (I11970,I12262,I12163);
not I_632 (I12369,I12245);
nand I_633 (I12386,I12163,I12369);
not I_634 (I11964,I12386);
nor I_635 (I11967,I12027,I12386);
nor I_636 (I11979,I12369,I12027);
nand I_637 (I12445,I12146,I12245);
nor I_638 (I11961,I12044,I12445);
not I_639 (I12503,I1605);
or I_640 (I12520,I35615,I35594);
nand I_641 (I12537,I35603,I35612);
not I_642 (I12554,I12537);
nand I_643 (I12571,I12554,I12520);
not I_644 (I12588,I12571);
nand I_645 (I12605,I35609,I35594);
and I_646 (I12622,I12605,I35600);
DFFARX1 I_647 (I12622,I1598,I12503,I12648,);
not I_648 (I12656,I12648);
nor I_649 (I12673,I35591,I35594);
nor I_650 (I12690,I12648,I12673);
and I_651 (I12707,I12648,I12673);
nor I_652 (I12724,I12707,I12571);
DFFARX1 I_653 (I12724,I1598,I12503,I12483,);
nand I_654 (I12755,I35606,I35591);
nor I_655 (I12772,I12755,I35597);
nand I_656 (I12789,I12588,I12772);
not I_657 (I12492,I12789);
nor I_658 (I12495,I12690,I12789);
nor I_659 (I12834,I12772,I12554);
nor I_660 (I12486,I12656,I12834);
nor I_661 (I12480,I12772,I12673);
not I_662 (I12879,I12755);
nand I_663 (I12896,I12673,I12879);
not I_664 (I12474,I12896);
nor I_665 (I12477,I12537,I12896);
nor I_666 (I12489,I12879,I12537);
nand I_667 (I12955,I12656,I12755);
nor I_668 (I12471,I12554,I12955);
not I_669 (I13013,I1605);
or I_670 (I13030,I4770,I4770);
nand I_671 (I13047,I4773,I4776);
not I_672 (I13064,I13047);
nand I_673 (I13081,I13064,I13030);
not I_674 (I13098,I13081);
nand I_675 (I13115,I4785,I4791);
and I_676 (I13132,I13115,I4779);
DFFARX1 I_677 (I13132,I1598,I13013,I13158,);
not I_678 (I13166,I13158);
nor I_679 (I13183,I4776,I4791);
nor I_680 (I13200,I13158,I13183);
and I_681 (I13217,I13158,I13183);
nor I_682 (I13234,I13217,I13081);
DFFARX1 I_683 (I13234,I1598,I13013,I12993,);
nand I_684 (I13265,I4773,I4782);
nor I_685 (I13282,I13265,I4788);
nand I_686 (I13299,I13098,I13282);
not I_687 (I13002,I13299);
nor I_688 (I13005,I13200,I13299);
nor I_689 (I13344,I13282,I13064);
nor I_690 (I12996,I13166,I13344);
nor I_691 (I12990,I13282,I13183);
not I_692 (I13389,I13265);
nand I_693 (I13406,I13183,I13389);
not I_694 (I12984,I13406);
nor I_695 (I12987,I13047,I13406);
nor I_696 (I12999,I13389,I13047);
nand I_697 (I13465,I13166,I13265);
nor I_698 (I12981,I13064,I13465);
not I_699 (I13523,I1605);
or I_700 (I13540,I58683,I58677);
nand I_701 (I13557,I58686,I58689);
not I_702 (I13574,I13557);
nand I_703 (I13591,I13574,I13540);
not I_704 (I13608,I13591);
nand I_705 (I13625,I58680,I58683);
and I_706 (I13642,I13625,I58677);
DFFARX1 I_707 (I13642,I1598,I13523,I13668,);
not I_708 (I13676,I13668);
nor I_709 (I13693,I58695,I58683);
nor I_710 (I13710,I13668,I13693);
and I_711 (I13727,I13668,I13693);
nor I_712 (I13744,I13727,I13591);
DFFARX1 I_713 (I13744,I1598,I13523,I13503,);
nand I_714 (I13775,I58692,I58680);
nor I_715 (I13792,I13775,I58698);
nand I_716 (I13809,I13608,I13792);
not I_717 (I13512,I13809);
nor I_718 (I13515,I13710,I13809);
nor I_719 (I13854,I13792,I13574);
nor I_720 (I13506,I13676,I13854);
nor I_721 (I13500,I13792,I13693);
not I_722 (I13899,I13775);
nand I_723 (I13916,I13693,I13899);
not I_724 (I13494,I13916);
nor I_725 (I13497,I13557,I13916);
nor I_726 (I13509,I13899,I13557);
nand I_727 (I13975,I13676,I13775);
nor I_728 (I13491,I13574,I13975);
not I_729 (I14033,I1605);
or I_730 (I14050,I46644,I46647);
nand I_731 (I14067,I46653,I46641);
not I_732 (I14084,I14067);
nand I_733 (I14101,I14084,I14050);
not I_734 (I14118,I14101);
nand I_735 (I14135,I46659,I46662);
and I_736 (I14152,I14135,I46656);
DFFARX1 I_737 (I14152,I1598,I14033,I14178,);
not I_738 (I14186,I14178);
nor I_739 (I14203,I46644,I46662);
nor I_740 (I14220,I14178,I14203);
and I_741 (I14237,I14178,I14203);
nor I_742 (I14254,I14237,I14101);
DFFARX1 I_743 (I14254,I1598,I14033,I14013,);
nand I_744 (I14285,I46647,I46650);
nor I_745 (I14302,I14285,I46641);
nand I_746 (I14319,I14118,I14302);
not I_747 (I14022,I14319);
nor I_748 (I14025,I14220,I14319);
nor I_749 (I14364,I14302,I14084);
nor I_750 (I14016,I14186,I14364);
nor I_751 (I14010,I14302,I14203);
not I_752 (I14409,I14285);
nand I_753 (I14426,I14203,I14409);
not I_754 (I14004,I14426);
nor I_755 (I14007,I14067,I14426);
nor I_756 (I14019,I14409,I14067);
nand I_757 (I14485,I14186,I14285);
nor I_758 (I14001,I14084,I14485);
not I_759 (I14543,I1605);
or I_760 (I14560,I68078,I68078);
nand I_761 (I14577,I68093,I68096);
not I_762 (I14594,I14577);
nand I_763 (I14611,I14594,I14560);
not I_764 (I14628,I14611);
nand I_765 (I14645,I68084,I68087);
and I_766 (I14662,I14645,I68081);
DFFARX1 I_767 (I14662,I1598,I14543,I14688,);
not I_768 (I14696,I14688);
nor I_769 (I14713,I68087,I68087);
nor I_770 (I14730,I14688,I14713);
and I_771 (I14747,I14688,I14713);
nor I_772 (I14764,I14747,I14611);
DFFARX1 I_773 (I14764,I1598,I14543,I14523,);
nand I_774 (I14795,I68090,I68084);
nor I_775 (I14812,I14795,I68081);
nand I_776 (I14829,I14628,I14812);
not I_777 (I14532,I14829);
nor I_778 (I14535,I14730,I14829);
nor I_779 (I14874,I14812,I14594);
nor I_780 (I14526,I14696,I14874);
nor I_781 (I14520,I14812,I14713);
not I_782 (I14919,I14795);
nand I_783 (I14936,I14713,I14919);
not I_784 (I14514,I14936);
nor I_785 (I14517,I14577,I14936);
nor I_786 (I14529,I14919,I14577);
nand I_787 (I14995,I14696,I14795);
nor I_788 (I14511,I14594,I14995);
not I_789 (I15053,I1605);
or I_790 (I15070,I61845,I61839);
nand I_791 (I15087,I61848,I61851);
not I_792 (I15104,I15087);
nand I_793 (I15121,I15104,I15070);
not I_794 (I15138,I15121);
nand I_795 (I15155,I61842,I61845);
and I_796 (I15172,I15155,I61839);
DFFARX1 I_797 (I15172,I1598,I15053,I15198,);
not I_798 (I15206,I15198);
nor I_799 (I15223,I61857,I61845);
nor I_800 (I15240,I15198,I15223);
and I_801 (I15257,I15198,I15223);
nor I_802 (I15274,I15257,I15121);
DFFARX1 I_803 (I15274,I1598,I15053,I15033,);
nand I_804 (I15305,I61854,I61842);
nor I_805 (I15322,I15305,I61860);
nand I_806 (I15339,I15138,I15322);
not I_807 (I15042,I15339);
nor I_808 (I15045,I15240,I15339);
nor I_809 (I15384,I15322,I15104);
nor I_810 (I15036,I15206,I15384);
nor I_811 (I15030,I15322,I15223);
not I_812 (I15429,I15305);
nand I_813 (I15446,I15223,I15429);
not I_814 (I15024,I15446);
nor I_815 (I15027,I15087,I15446);
nor I_816 (I15039,I15429,I15087);
nand I_817 (I15505,I15206,I15305);
nor I_818 (I15021,I15104,I15505);
not I_819 (I15563,I1605);
or I_820 (I15580,I46168,I46171);
nand I_821 (I15597,I46177,I46165);
not I_822 (I15614,I15597);
nand I_823 (I15631,I15614,I15580);
not I_824 (I15648,I15631);
nand I_825 (I15665,I46183,I46186);
and I_826 (I15682,I15665,I46180);
DFFARX1 I_827 (I15682,I1598,I15563,I15708,);
not I_828 (I15716,I15708);
nor I_829 (I15733,I46168,I46186);
nor I_830 (I15750,I15708,I15733);
and I_831 (I15767,I15708,I15733);
nor I_832 (I15784,I15767,I15631);
DFFARX1 I_833 (I15784,I1598,I15563,I15543,);
nand I_834 (I15815,I46171,I46174);
nor I_835 (I15832,I15815,I46165);
nand I_836 (I15849,I15648,I15832);
not I_837 (I15552,I15849);
nor I_838 (I15555,I15750,I15849);
nor I_839 (I15894,I15832,I15614);
nor I_840 (I15546,I15716,I15894);
nor I_841 (I15540,I15832,I15733);
not I_842 (I15939,I15815);
nand I_843 (I15956,I15733,I15939);
not I_844 (I15534,I15956);
nor I_845 (I15537,I15597,I15956);
nor I_846 (I15549,I15939,I15597);
nand I_847 (I16015,I15716,I15815);
nor I_848 (I15531,I15614,I16015);
not I_849 (I16073,I1605);
or I_850 (I16090,I70730,I70730);
nand I_851 (I16107,I70745,I70748);
not I_852 (I16124,I16107);
nand I_853 (I16141,I16124,I16090);
not I_854 (I16158,I16141);
nand I_855 (I16175,I70736,I70739);
and I_856 (I16192,I16175,I70733);
DFFARX1 I_857 (I16192,I1598,I16073,I16218,);
not I_858 (I16226,I16218);
nor I_859 (I16243,I70739,I70739);
nor I_860 (I16260,I16218,I16243);
and I_861 (I16277,I16218,I16243);
nor I_862 (I16294,I16277,I16141);
DFFARX1 I_863 (I16294,I1598,I16073,I16053,);
nand I_864 (I16325,I70742,I70736);
nor I_865 (I16342,I16325,I70733);
nand I_866 (I16359,I16158,I16342);
not I_867 (I16062,I16359);
nor I_868 (I16065,I16260,I16359);
nor I_869 (I16404,I16342,I16124);
nor I_870 (I16056,I16226,I16404);
nor I_871 (I16050,I16342,I16243);
not I_872 (I16449,I16325);
nand I_873 (I16466,I16243,I16449);
not I_874 (I16044,I16466);
nor I_875 (I16047,I16107,I16466);
nor I_876 (I16059,I16449,I16107);
nand I_877 (I16525,I16226,I16325);
nor I_878 (I16041,I16124,I16525);
not I_879 (I16583,I1605);
or I_880 (I16600,I74708,I74708);
nand I_881 (I16617,I74723,I74726);
not I_882 (I16634,I16617);
nand I_883 (I16651,I16634,I16600);
not I_884 (I16668,I16651);
nand I_885 (I16685,I74714,I74717);
and I_886 (I16702,I16685,I74711);
DFFARX1 I_887 (I16702,I1598,I16583,I16728,);
not I_888 (I16736,I16728);
nor I_889 (I16753,I74717,I74717);
nor I_890 (I16770,I16728,I16753);
and I_891 (I16787,I16728,I16753);
nor I_892 (I16804,I16787,I16651);
DFFARX1 I_893 (I16804,I1598,I16583,I16563,);
nand I_894 (I16835,I74720,I74714);
nor I_895 (I16852,I16835,I74711);
nand I_896 (I16869,I16668,I16852);
not I_897 (I16572,I16869);
nor I_898 (I16575,I16770,I16869);
nor I_899 (I16914,I16852,I16634);
nor I_900 (I16566,I16736,I16914);
nor I_901 (I16560,I16852,I16753);
not I_902 (I16959,I16835);
nand I_903 (I16976,I16753,I16959);
not I_904 (I16554,I16976);
nor I_905 (I16557,I16617,I16976);
nor I_906 (I16569,I16959,I16617);
nand I_907 (I17035,I16736,I16835);
nor I_908 (I16551,I16634,I17035);
not I_909 (I17093,I1605);
or I_910 (I17110,I54464,I54461);
nand I_911 (I17127,I54467,I54479);
not I_912 (I17144,I17127);
nand I_913 (I17161,I17144,I17110);
not I_914 (I17178,I17161);
nand I_915 (I17195,I54464,I54470);
and I_916 (I17212,I17195,I54476);
DFFARX1 I_917 (I17212,I1598,I17093,I17238,);
not I_918 (I17246,I17238);
nor I_919 (I17263,I54482,I54470);
nor I_920 (I17280,I17238,I17263);
and I_921 (I17297,I17238,I17263);
nor I_922 (I17314,I17297,I17161);
DFFARX1 I_923 (I17314,I1598,I17093,I17073,);
nand I_924 (I17345,I54473,I54467);
nor I_925 (I17362,I17345,I54461);
nand I_926 (I17379,I17178,I17362);
not I_927 (I17082,I17379);
nor I_928 (I17085,I17280,I17379);
nor I_929 (I17424,I17362,I17144);
nor I_930 (I17076,I17246,I17424);
nor I_931 (I17070,I17362,I17263);
not I_932 (I17469,I17345);
nand I_933 (I17486,I17263,I17469);
not I_934 (I17064,I17486);
nor I_935 (I17067,I17127,I17486);
nor I_936 (I17079,I17469,I17127);
nand I_937 (I17545,I17246,I17345);
nor I_938 (I17061,I17144,I17545);
not I_939 (I17603,I1605);
or I_940 (I17620,I1207,I1055);
nand I_941 (I17637,I1359,I775);
not I_942 (I17654,I17637);
nand I_943 (I17671,I17654,I17620);
not I_944 (I17688,I17671);
nand I_945 (I17705,I1431,I1423);
and I_946 (I17722,I17705,I1335);
DFFARX1 I_947 (I17722,I1598,I17603,I17748,);
not I_948 (I17756,I17748);
nor I_949 (I17773,I1063,I1423);
nor I_950 (I17790,I17748,I17773);
and I_951 (I17807,I17748,I17773);
nor I_952 (I17824,I17807,I17671);
DFFARX1 I_953 (I17824,I1598,I17603,I17583,);
nand I_954 (I17855,I983,I1183);
nor I_955 (I17872,I17855,I1447);
nand I_956 (I17889,I17688,I17872);
not I_957 (I17592,I17889);
nor I_958 (I17595,I17790,I17889);
nor I_959 (I17934,I17872,I17654);
nor I_960 (I17586,I17756,I17934);
nor I_961 (I17580,I17872,I17773);
not I_962 (I17979,I17855);
nand I_963 (I17996,I17773,I17979);
not I_964 (I17574,I17996);
nor I_965 (I17577,I17637,I17996);
nor I_966 (I17589,I17979,I17637);
nand I_967 (I18055,I17756,I17855);
nor I_968 (I17571,I17654,I18055);
not I_969 (I18113,I1605);
or I_970 (I18130,I1167,I1215);
nand I_971 (I18147,I1271,I1255);
not I_972 (I18164,I18147);
nand I_973 (I18181,I18164,I18130);
not I_974 (I18198,I18181);
nand I_975 (I18215,I727,I655);
and I_976 (I18232,I18215,I1031);
DFFARX1 I_977 (I18232,I1598,I18113,I18258,);
not I_978 (I18266,I18258);
nor I_979 (I18283,I1535,I655);
nor I_980 (I18300,I18258,I18283);
and I_981 (I18317,I18258,I18283);
nor I_982 (I18334,I18317,I18181);
DFFARX1 I_983 (I18334,I1598,I18113,I18093,);
nand I_984 (I18365,I1343,I1415);
nor I_985 (I18382,I18365,I1511);
nand I_986 (I18399,I18198,I18382);
not I_987 (I18102,I18399);
nor I_988 (I18105,I18300,I18399);
nor I_989 (I18444,I18382,I18164);
nor I_990 (I18096,I18266,I18444);
nor I_991 (I18090,I18382,I18283);
not I_992 (I18489,I18365);
nand I_993 (I18506,I18283,I18489);
not I_994 (I18084,I18506);
nor I_995 (I18087,I18147,I18506);
nor I_996 (I18099,I18489,I18147);
nand I_997 (I18565,I18266,I18365);
nor I_998 (I18081,I18164,I18565);
not I_999 (I18623,I1605);
or I_1000 (I18640,I39980,I39983);
nand I_1001 (I18657,I39989,I39977);
not I_1002 (I18674,I18657);
nand I_1003 (I18691,I18674,I18640);
not I_1004 (I18708,I18691);
nand I_1005 (I18725,I39995,I39998);
and I_1006 (I18742,I18725,I39992);
DFFARX1 I_1007 (I18742,I1598,I18623,I18768,);
not I_1008 (I18776,I18768);
nor I_1009 (I18793,I39980,I39998);
nor I_1010 (I18810,I18768,I18793);
and I_1011 (I18827,I18768,I18793);
nor I_1012 (I18844,I18827,I18691);
DFFARX1 I_1013 (I18844,I1598,I18623,I18603,);
nand I_1014 (I18875,I39983,I39986);
nor I_1015 (I18892,I18875,I39977);
nand I_1016 (I18909,I18708,I18892);
not I_1017 (I18612,I18909);
nor I_1018 (I18615,I18810,I18909);
nor I_1019 (I18954,I18892,I18674);
nor I_1020 (I18606,I18776,I18954);
nor I_1021 (I18600,I18892,I18793);
not I_1022 (I18999,I18875);
nand I_1023 (I19016,I18793,I18999);
not I_1024 (I18594,I19016);
nor I_1025 (I18597,I18657,I19016);
nor I_1026 (I18609,I18999,I18657);
nand I_1027 (I19075,I18776,I18875);
nor I_1028 (I18591,I18674,I19075);
not I_1029 (I19133,I1605);
or I_1030 (I19150,I26129,I26108);
nand I_1031 (I19167,I26117,I26126);
not I_1032 (I19184,I19167);
nand I_1033 (I19201,I19184,I19150);
not I_1034 (I19218,I19201);
nand I_1035 (I19235,I26123,I26108);
and I_1036 (I19252,I19235,I26114);
DFFARX1 I_1037 (I19252,I1598,I19133,I19278,);
not I_1038 (I19286,I19278);
nor I_1039 (I19303,I26105,I26108);
nor I_1040 (I19320,I19278,I19303);
and I_1041 (I19337,I19278,I19303);
nor I_1042 (I19354,I19337,I19201);
DFFARX1 I_1043 (I19354,I1598,I19133,I19113,);
nand I_1044 (I19385,I26120,I26105);
nor I_1045 (I19402,I19385,I26111);
nand I_1046 (I19419,I19218,I19402);
not I_1047 (I19122,I19419);
nor I_1048 (I19125,I19320,I19419);
nor I_1049 (I19464,I19402,I19184);
nor I_1050 (I19116,I19286,I19464);
nor I_1051 (I19110,I19402,I19303);
not I_1052 (I19509,I19385);
nand I_1053 (I19526,I19303,I19509);
not I_1054 (I19104,I19526);
nor I_1055 (I19107,I19167,I19526);
nor I_1056 (I19119,I19509,I19167);
nand I_1057 (I19585,I19286,I19385);
nor I_1058 (I19101,I19184,I19585);
not I_1059 (I19643,I1605);
or I_1060 (I19660,I77360,I77360);
nand I_1061 (I19677,I77375,I77378);
not I_1062 (I19694,I19677);
nand I_1063 (I19711,I19694,I19660);
not I_1064 (I19728,I19711);
nand I_1065 (I19745,I77366,I77369);
and I_1066 (I19762,I19745,I77363);
DFFARX1 I_1067 (I19762,I1598,I19643,I19788,);
not I_1068 (I19796,I19788);
nor I_1069 (I19813,I77369,I77369);
nor I_1070 (I19830,I19788,I19813);
and I_1071 (I19847,I19788,I19813);
nor I_1072 (I19864,I19847,I19711);
DFFARX1 I_1073 (I19864,I1598,I19643,I19623,);
nand I_1074 (I19895,I77372,I77366);
nor I_1075 (I19912,I19895,I77363);
nand I_1076 (I19929,I19728,I19912);
not I_1077 (I19632,I19929);
nor I_1078 (I19635,I19830,I19929);
nor I_1079 (I19974,I19912,I19694);
nor I_1080 (I19626,I19796,I19974);
nor I_1081 (I19620,I19912,I19813);
not I_1082 (I20019,I19895);
nand I_1083 (I20036,I19813,I20019);
not I_1084 (I19614,I20036);
nor I_1085 (I19617,I19677,I20036);
nor I_1086 (I19629,I20019,I19677);
nand I_1087 (I20095,I19796,I19895);
nor I_1088 (I19611,I19694,I20095);
not I_1089 (I20153,I1605);
or I_1090 (I20170,I41884,I41887);
nand I_1091 (I20187,I41893,I41881);
not I_1092 (I20204,I20187);
nand I_1093 (I20221,I20204,I20170);
not I_1094 (I20238,I20221);
nand I_1095 (I20255,I41899,I41902);
and I_1096 (I20272,I20255,I41896);
DFFARX1 I_1097 (I20272,I1598,I20153,I20298,);
not I_1098 (I20306,I20298);
nor I_1099 (I20323,I41884,I41902);
nor I_1100 (I20340,I20298,I20323);
and I_1101 (I20357,I20298,I20323);
nor I_1102 (I20374,I20357,I20221);
DFFARX1 I_1103 (I20374,I1598,I20153,I20133,);
nand I_1104 (I20405,I41887,I41890);
nor I_1105 (I20422,I20405,I41881);
nand I_1106 (I20439,I20238,I20422);
not I_1107 (I20142,I20439);
nor I_1108 (I20145,I20340,I20439);
nor I_1109 (I20484,I20422,I20204);
nor I_1110 (I20136,I20306,I20484);
nor I_1111 (I20130,I20422,I20323);
not I_1112 (I20529,I20405);
nand I_1113 (I20546,I20323,I20529);
not I_1114 (I20124,I20546);
nor I_1115 (I20127,I20187,I20546);
nor I_1116 (I20139,I20529,I20187);
nand I_1117 (I20605,I20306,I20405);
nor I_1118 (I20121,I20204,I20605);
not I_1119 (I20663,I1605);
or I_1120 (I20680,I2135,I2135);
nand I_1121 (I20697,I2138,I2141);
not I_1122 (I20714,I20697);
nand I_1123 (I20731,I20714,I20680);
not I_1124 (I20748,I20731);
nand I_1125 (I20765,I2150,I2156);
and I_1126 (I20782,I20765,I2144);
DFFARX1 I_1127 (I20782,I1598,I20663,I20808,);
not I_1128 (I20816,I20808);
nor I_1129 (I20833,I2141,I2156);
nor I_1130 (I20850,I20808,I20833);
and I_1131 (I20867,I20808,I20833);
nor I_1132 (I20884,I20867,I20731);
DFFARX1 I_1133 (I20884,I1598,I20663,I20643,);
nand I_1134 (I20915,I2138,I2147);
nor I_1135 (I20932,I20915,I2153);
nand I_1136 (I20949,I20748,I20932);
not I_1137 (I20652,I20949);
nor I_1138 (I20655,I20850,I20949);
nor I_1139 (I20994,I20932,I20714);
nor I_1140 (I20646,I20816,I20994);
nor I_1141 (I20640,I20932,I20833);
not I_1142 (I21039,I20915);
nand I_1143 (I21056,I20833,I21039);
not I_1144 (I20634,I21056);
nor I_1145 (I20637,I20697,I21056);
nor I_1146 (I20649,I21039,I20697);
nand I_1147 (I21115,I20816,I20915);
nor I_1148 (I20631,I20714,I21115);
not I_1149 (I21167,I1605);
and I_1150 (I21184,I32450,I32432);
nor I_1151 (I21201,I21184,I32453);
nand I_1152 (I21218,I32429,I32444);
nor I_1153 (I21235,I21218,I21201);
nor I_1154 (I21141,I21235,I21218);
not I_1155 (I21266,I21235);
not I_1156 (I21283,I21218);
or I_1157 (I21300,I32447,I32429);
nor I_1158 (I21317,I21300,I32435);
nand I_1159 (I21334,I21283,I21317);
not I_1160 (I21156,I21334);
nor I_1161 (I21365,I21235,I32441);
and I_1162 (I21382,I32438,I32432);
nor I_1163 (I21399,I21382,I21235);
nor I_1164 (I21159,I21399,I21334);
nor I_1165 (I21144,I21382,I21317);
nand I_1166 (I21444,I21382,I32441);
not I_1167 (I21461,I21444);
nand I_1168 (I21478,I21317,I21461);
nand I_1169 (I21495,I21266,I21478);
DFFARX1 I_1170 (I21495,I1598,I21167,I21147,);
nand I_1171 (I21153,I21382,I21218);
nand I_1172 (I21150,I21365,I21382);
not I_1173 (I21575,I1605);
and I_1174 (I21592,I68977,I68971);
nor I_1175 (I21609,I21592,I68974);
nand I_1176 (I21626,I68968,I68968);
nor I_1177 (I21643,I21626,I21609);
nor I_1178 (I21549,I21643,I21626);
not I_1179 (I21674,I21643);
not I_1180 (I21691,I21626);
or I_1181 (I21708,I68965,I68962);
nor I_1182 (I21725,I21708,I68965);
nand I_1183 (I21742,I21691,I21725);
not I_1184 (I21564,I21742);
nor I_1185 (I21773,I21643,I68962);
and I_1186 (I21790,I68971,I68980);
nor I_1187 (I21807,I21790,I21643);
nor I_1188 (I21567,I21807,I21742);
nor I_1189 (I21552,I21790,I21725);
nand I_1190 (I21852,I21790,I68962);
not I_1191 (I21869,I21852);
nand I_1192 (I21886,I21725,I21869);
nand I_1193 (I21903,I21674,I21886);
DFFARX1 I_1194 (I21903,I1598,I21575,I21555,);
nand I_1195 (I21561,I21790,I21626);
nand I_1196 (I21558,I21773,I21790);
not I_1197 (I21983,I1605);
and I_1198 (I22000,I887,I1095);
nor I_1199 (I22017,I22000,I1551);
nand I_1200 (I22034,I719,I927);
nor I_1201 (I22051,I22034,I22017);
nor I_1202 (I21957,I22051,I22034);
not I_1203 (I22082,I22051);
not I_1204 (I22099,I22034);
or I_1205 (I22116,I695,I1519);
nor I_1206 (I22133,I22116,I1071);
nand I_1207 (I22150,I22099,I22133);
not I_1208 (I21972,I22150);
nor I_1209 (I22181,I22051,I1047);
and I_1210 (I22198,I1319,I951);
nor I_1211 (I22215,I22198,I22051);
nor I_1212 (I21975,I22215,I22150);
nor I_1213 (I21960,I22198,I22133);
nand I_1214 (I22260,I22198,I1047);
not I_1215 (I22277,I22260);
nand I_1216 (I22294,I22133,I22277);
nand I_1217 (I22311,I22082,I22294);
DFFARX1 I_1218 (I22311,I1598,I21983,I21963,);
nand I_1219 (I21969,I22198,I22034);
nand I_1220 (I21966,I22181,I22198);
not I_1221 (I22391,I1605);
and I_1222 (I22408,I49021,I49021);
nor I_1223 (I22425,I22408,I49042);
nand I_1224 (I22442,I49024,I49027);
nor I_1225 (I22459,I22442,I22425);
nor I_1226 (I22365,I22459,I22442);
not I_1227 (I22490,I22459);
not I_1228 (I22507,I22442);
or I_1229 (I22524,I49030,I49039);
nor I_1230 (I22541,I22524,I49036);
nand I_1231 (I22558,I22507,I22541);
not I_1232 (I22380,I22558);
nor I_1233 (I22589,I22459,I49027);
and I_1234 (I22606,I49024,I49033);
nor I_1235 (I22623,I22606,I22459);
nor I_1236 (I22383,I22623,I22558);
nor I_1237 (I22368,I22606,I22541);
nand I_1238 (I22668,I22606,I49027);
not I_1239 (I22685,I22668);
nand I_1240 (I22702,I22541,I22685);
nand I_1241 (I22719,I22490,I22702);
DFFARX1 I_1242 (I22719,I1598,I22391,I22371,);
nand I_1243 (I22377,I22606,I22442);
nand I_1244 (I22374,I22589,I22606);
not I_1245 (I22799,I1605);
and I_1246 (I22816,I1375,I959);
nor I_1247 (I22833,I22816,I1311);
nand I_1248 (I22850,I1495,I1399);
nor I_1249 (I22867,I22850,I22833);
nor I_1250 (I22773,I22867,I22850);
not I_1251 (I22898,I22867);
not I_1252 (I22915,I22850);
or I_1253 (I22932,I1151,I1559);
nor I_1254 (I22949,I22932,I1383);
nand I_1255 (I22966,I22915,I22949);
not I_1256 (I22788,I22966);
nor I_1257 (I22997,I22867,I935);
and I_1258 (I23014,I1119,I855);
nor I_1259 (I23031,I23014,I22867);
nor I_1260 (I22791,I23031,I22966);
nor I_1261 (I22776,I23014,I22949);
nand I_1262 (I23076,I23014,I935);
not I_1263 (I23093,I23076);
nand I_1264 (I23110,I22949,I23093);
nand I_1265 (I23127,I22898,I23110);
DFFARX1 I_1266 (I23127,I1598,I22799,I22779,);
nand I_1267 (I22785,I23014,I22850);
nand I_1268 (I22782,I22997,I23014);
not I_1269 (I23207,I1605);
and I_1270 (I23224,I57114,I57099);
nor I_1271 (I23241,I23224,I57102);
nand I_1272 (I23258,I57096,I57111);
nor I_1273 (I23275,I23258,I23241);
nor I_1274 (I23181,I23275,I23258);
not I_1275 (I23306,I23275);
not I_1276 (I23323,I23258);
or I_1277 (I23340,I57099,I57102);
nor I_1278 (I23357,I23340,I57096);
nand I_1279 (I23374,I23323,I23357);
not I_1280 (I23196,I23374);
nor I_1281 (I23405,I23275,I57117);
and I_1282 (I23422,I57108,I57105);
nor I_1283 (I23439,I23422,I23275);
nor I_1284 (I23199,I23439,I23374);
nor I_1285 (I23184,I23422,I23357);
nand I_1286 (I23484,I23422,I57117);
not I_1287 (I23501,I23484);
nand I_1288 (I23518,I23357,I23501);
nand I_1289 (I23535,I23306,I23518);
DFFARX1 I_1290 (I23535,I1598,I23207,I23187,);
nand I_1291 (I23193,I23422,I23258);
nand I_1292 (I23190,I23405,I23422);
not I_1293 (I23615,I1605);
and I_1294 (I23632,I59222,I59207);
nor I_1295 (I23649,I23632,I59210);
nand I_1296 (I23666,I59204,I59219);
nor I_1297 (I23683,I23666,I23649);
nor I_1298 (I23589,I23683,I23666);
not I_1299 (I23714,I23683);
not I_1300 (I23731,I23666);
or I_1301 (I23748,I59207,I59210);
nor I_1302 (I23765,I23748,I59204);
nand I_1303 (I23782,I23731,I23765);
not I_1304 (I23604,I23782);
nor I_1305 (I23813,I23683,I59225);
and I_1306 (I23830,I59216,I59213);
nor I_1307 (I23847,I23830,I23683);
nor I_1308 (I23607,I23847,I23782);
nor I_1309 (I23592,I23830,I23765);
nand I_1310 (I23892,I23830,I59225);
not I_1311 (I23909,I23892);
nand I_1312 (I23926,I23765,I23909);
nand I_1313 (I23943,I23714,I23926);
DFFARX1 I_1314 (I23943,I1598,I23615,I23595,);
nand I_1315 (I23601,I23830,I23666);
nand I_1316 (I23598,I23813,I23830);
not I_1317 (I24029,I1605);
or I_1318 (I24046,I37121,I37124);
nand I_1319 (I24063,I37127,I37136);
not I_1320 (I24080,I24063);
nand I_1321 (I24097,I24080,I24046);
not I_1322 (I24114,I24097);
nand I_1323 (I24131,I37133,I37139);
and I_1324 (I24148,I24131,I37121);
DFFARX1 I_1325 (I24148,I1598,I24029,I24174,);
nor I_1326 (I23997,I24174,I24063);
nand I_1327 (I24196,I24114,I24174);
nor I_1328 (I24213,I24174,I24080);
not I_1329 (I24015,I24174);
nor I_1330 (I24244,I37124,I37139);
not I_1331 (I24261,I24244);
nand I_1332 (I24018,I24213,I24244);
not I_1333 (I24292,I37142);
nor I_1334 (I24309,I24174,I37142);
nand I_1335 (I24326,I37130,I37127);
nor I_1336 (I24000,I24326,I24063);
not I_1337 (I24357,I24326);
nor I_1338 (I24374,I24244,I24357);
nor I_1339 (I24021,I24374,I24097);
nand I_1340 (I24405,I24357,I24292);
nand I_1341 (I24006,I24114,I24405);
nand I_1342 (I24436,I24196,I24405);
DFFARX1 I_1343 (I24436,I1598,I24029,I24009,);
nand I_1344 (I24467,I24261,I24326);
nor I_1345 (I24003,I24114,I24467);
nor I_1346 (I24498,I24261,I24326);
nand I_1347 (I24012,I24498,I24309);
not I_1348 (I24556,I1605);
or I_1349 (I24573,I9414,I9411);
nand I_1350 (I24590,I9417,I9414);
not I_1351 (I24607,I24590);
nand I_1352 (I24624,I24607,I24573);
not I_1353 (I24641,I24624);
nand I_1354 (I24658,I9432,I9435);
and I_1355 (I24675,I24658,I9411);
DFFARX1 I_1356 (I24675,I1598,I24556,I24701,);
nor I_1357 (I24524,I24701,I24590);
nand I_1358 (I24723,I24641,I24701);
nor I_1359 (I24740,I24701,I24607);
not I_1360 (I24542,I24701);
nor I_1361 (I24771,I9429,I9435);
not I_1362 (I24788,I24771);
nand I_1363 (I24545,I24740,I24771);
not I_1364 (I24819,I9420);
nor I_1365 (I24836,I24701,I9420);
nand I_1366 (I24853,I9423,I9426);
nor I_1367 (I24527,I24853,I24590);
not I_1368 (I24884,I24853);
nor I_1369 (I24901,I24771,I24884);
nor I_1370 (I24548,I24901,I24624);
nand I_1371 (I24932,I24884,I24819);
nand I_1372 (I24533,I24641,I24932);
nand I_1373 (I24963,I24723,I24932);
DFFARX1 I_1374 (I24963,I1598,I24556,I24536,);
nand I_1375 (I24994,I24788,I24853);
nor I_1376 (I24530,I24641,I24994);
nor I_1377 (I25025,I24788,I24853);
nand I_1378 (I24539,I25025,I24836);
not I_1379 (I25083,I1605);
or I_1380 (I25100,I44261,I44264);
nand I_1381 (I25117,I44267,I44276);
not I_1382 (I25134,I25117);
nand I_1383 (I25151,I25134,I25100);
not I_1384 (I25168,I25151);
nand I_1385 (I25185,I44273,I44279);
and I_1386 (I25202,I25185,I44261);
DFFARX1 I_1387 (I25202,I1598,I25083,I25228,);
nor I_1388 (I25051,I25228,I25117);
nand I_1389 (I25250,I25168,I25228);
nor I_1390 (I25267,I25228,I25134);
not I_1391 (I25069,I25228);
nor I_1392 (I25298,I44264,I44279);
not I_1393 (I25315,I25298);
nand I_1394 (I25072,I25267,I25298);
not I_1395 (I25346,I44282);
nor I_1396 (I25363,I25228,I44282);
nand I_1397 (I25380,I44270,I44267);
nor I_1398 (I25054,I25380,I25117);
not I_1399 (I25411,I25380);
nor I_1400 (I25428,I25298,I25411);
nor I_1401 (I25075,I25428,I25151);
nand I_1402 (I25459,I25411,I25346);
nand I_1403 (I25060,I25168,I25459);
nand I_1404 (I25490,I25250,I25459);
DFFARX1 I_1405 (I25490,I1598,I25083,I25063,);
nand I_1406 (I25521,I25315,I25380);
nor I_1407 (I25057,I25168,I25521);
nor I_1408 (I25552,I25315,I25380);
nand I_1409 (I25066,I25552,I25363);
not I_1410 (I25610,I1605);
or I_1411 (I25627,I71620,I71617);
nand I_1412 (I25644,I71629,I71632);
not I_1413 (I25661,I25644);
nand I_1414 (I25678,I25661,I25627);
not I_1415 (I25695,I25678);
nand I_1416 (I25712,I71623,I71614);
and I_1417 (I25729,I25712,I71614);
DFFARX1 I_1418 (I25729,I1598,I25610,I25755,);
nor I_1419 (I25578,I25755,I25644);
nand I_1420 (I25777,I25695,I25755);
nor I_1421 (I25794,I25755,I25661);
not I_1422 (I25596,I25755);
nor I_1423 (I25825,I71617,I71614);
not I_1424 (I25842,I25825);
nand I_1425 (I25599,I25794,I25825);
not I_1426 (I25873,I71620);
nor I_1427 (I25890,I25755,I71620);
nand I_1428 (I25907,I71623,I71626);
nor I_1429 (I25581,I25907,I25644);
not I_1430 (I25938,I25907);
nor I_1431 (I25955,I25825,I25938);
nor I_1432 (I25602,I25955,I25678);
nand I_1433 (I25986,I25938,I25873);
nand I_1434 (I25587,I25695,I25986);
nand I_1435 (I26017,I25777,I25986);
DFFARX1 I_1436 (I26017,I1598,I25610,I25590,);
nand I_1437 (I26048,I25842,I25907);
nor I_1438 (I25584,I25695,I26048);
nor I_1439 (I26079,I25842,I25907);
nand I_1440 (I25593,I26079,I25890);
not I_1441 (I26137,I1605);
or I_1442 (I26154,I67127,I67115);
nand I_1443 (I26171,I67109,I67109);
not I_1444 (I26188,I26171);
nand I_1445 (I26205,I26188,I26154);
not I_1446 (I26222,I26205);
nand I_1447 (I26239,I67112,I67112);
and I_1448 (I26256,I26239,I67118);
DFFARX1 I_1449 (I26256,I1598,I26137,I26282,);
nor I_1450 (I26105,I26282,I26171);
nand I_1451 (I26304,I26222,I26282);
nor I_1452 (I26321,I26282,I26188);
not I_1453 (I26123,I26282);
nor I_1454 (I26352,I67124,I67112);
not I_1455 (I26369,I26352);
nand I_1456 (I26126,I26321,I26352);
not I_1457 (I26400,I67130);
nor I_1458 (I26417,I26282,I67130);
nand I_1459 (I26434,I67115,I67121);
nor I_1460 (I26108,I26434,I26171);
not I_1461 (I26465,I26434);
nor I_1462 (I26482,I26352,I26465);
nor I_1463 (I26129,I26482,I26205);
nand I_1464 (I26513,I26465,I26400);
nand I_1465 (I26114,I26222,I26513);
nand I_1466 (I26544,I26304,I26513);
DFFARX1 I_1467 (I26544,I1598,I26137,I26117,);
nand I_1468 (I26575,I26369,I26434);
nor I_1469 (I26111,I26222,I26575);
nor I_1470 (I26606,I26369,I26434);
nand I_1471 (I26120,I26606,I26417);
not I_1472 (I26664,I1605);
or I_1473 (I26681,I703,I1543);
nand I_1474 (I26698,I631,I1007);
not I_1475 (I26715,I26698);
nand I_1476 (I26732,I26715,I26681);
not I_1477 (I26749,I26732);
nand I_1478 (I26766,I687,I1191);
and I_1479 (I26783,I26766,I1111);
DFFARX1 I_1480 (I26783,I1598,I26664,I26809,);
nor I_1481 (I26632,I26809,I26698);
nand I_1482 (I26831,I26749,I26809);
nor I_1483 (I26848,I26809,I26715);
not I_1484 (I26650,I26809);
nor I_1485 (I26879,I1455,I1191);
not I_1486 (I26896,I26879);
nand I_1487 (I26653,I26848,I26879);
not I_1488 (I26927,I903);
nor I_1489 (I26944,I26809,I903);
nand I_1490 (I26961,I1199,I679);
nor I_1491 (I26635,I26961,I26698);
not I_1492 (I26992,I26961);
nor I_1493 (I27009,I26879,I26992);
nor I_1494 (I26656,I27009,I26732);
nand I_1495 (I27040,I26992,I26927);
nand I_1496 (I26641,I26749,I27040);
nand I_1497 (I27071,I26831,I27040);
DFFARX1 I_1498 (I27071,I1598,I26664,I26644,);
nand I_1499 (I27102,I26896,I26961);
nor I_1500 (I26638,I26749,I27102);
nor I_1501 (I27133,I26896,I26961);
nand I_1502 (I26647,I27133,I26944);
not I_1503 (I27191,I1605);
or I_1504 (I27208,I59749,I59737);
nand I_1505 (I27225,I59731,I59731);
not I_1506 (I27242,I27225);
nand I_1507 (I27259,I27242,I27208);
not I_1508 (I27276,I27259);
nand I_1509 (I27293,I59734,I59734);
and I_1510 (I27310,I27293,I59740);
DFFARX1 I_1511 (I27310,I1598,I27191,I27336,);
nor I_1512 (I27159,I27336,I27225);
nand I_1513 (I27358,I27276,I27336);
nor I_1514 (I27375,I27336,I27242);
not I_1515 (I27177,I27336);
nor I_1516 (I27406,I59746,I59734);
not I_1517 (I27423,I27406);
nand I_1518 (I27180,I27375,I27406);
not I_1519 (I27454,I59752);
nor I_1520 (I27471,I27336,I59752);
nand I_1521 (I27488,I59737,I59743);
nor I_1522 (I27162,I27488,I27225);
not I_1523 (I27519,I27488);
nor I_1524 (I27536,I27406,I27519);
nor I_1525 (I27183,I27536,I27259);
nand I_1526 (I27567,I27519,I27454);
nand I_1527 (I27168,I27276,I27567);
nand I_1528 (I27598,I27358,I27567);
DFFARX1 I_1529 (I27598,I1598,I27191,I27171,);
nand I_1530 (I27629,I27423,I27488);
nor I_1531 (I27165,I27276,I27629);
nor I_1532 (I27660,I27423,I27488);
nand I_1533 (I27174,I27660,I27471);
not I_1534 (I27718,I1605);
or I_1535 (I27735,I71178,I71175);
nand I_1536 (I27752,I71187,I71190);
not I_1537 (I27769,I27752);
nand I_1538 (I27786,I27769,I27735);
not I_1539 (I27803,I27786);
nand I_1540 (I27820,I71181,I71172);
and I_1541 (I27837,I27820,I71172);
DFFARX1 I_1542 (I27837,I1598,I27718,I27863,);
nor I_1543 (I27686,I27863,I27752);
nand I_1544 (I27885,I27803,I27863);
nor I_1545 (I27902,I27863,I27769);
not I_1546 (I27704,I27863);
nor I_1547 (I27933,I71175,I71172);
not I_1548 (I27950,I27933);
nand I_1549 (I27707,I27902,I27933);
not I_1550 (I27981,I71178);
nor I_1551 (I27998,I27863,I71178);
nand I_1552 (I28015,I71181,I71184);
nor I_1553 (I27689,I28015,I27752);
not I_1554 (I28046,I28015);
nor I_1555 (I28063,I27933,I28046);
nor I_1556 (I27710,I28063,I27786);
nand I_1557 (I28094,I28046,I27981);
nand I_1558 (I27695,I27803,I28094);
nand I_1559 (I28125,I27885,I28094);
DFFARX1 I_1560 (I28125,I1598,I27718,I27698,);
nand I_1561 (I28156,I27950,I28015);
nor I_1562 (I27692,I27803,I28156);
nor I_1563 (I28187,I27950,I28015);
nand I_1564 (I27701,I28187,I27998);
not I_1565 (I28245,I1605);
or I_1566 (I28262,I14514,I14511);
nand I_1567 (I28279,I14517,I14514);
not I_1568 (I28296,I28279);
nand I_1569 (I28313,I28296,I28262);
not I_1570 (I28330,I28313);
nand I_1571 (I28347,I14532,I14535);
and I_1572 (I28364,I28347,I14511);
DFFARX1 I_1573 (I28364,I1598,I28245,I28390,);
nor I_1574 (I28213,I28390,I28279);
nand I_1575 (I28412,I28330,I28390);
nor I_1576 (I28429,I28390,I28296);
not I_1577 (I28231,I28390);
nor I_1578 (I28460,I14529,I14535);
not I_1579 (I28477,I28460);
nand I_1580 (I28234,I28429,I28460);
not I_1581 (I28508,I14520);
nor I_1582 (I28525,I28390,I14520);
nand I_1583 (I28542,I14523,I14526);
nor I_1584 (I28216,I28542,I28279);
not I_1585 (I28573,I28542);
nor I_1586 (I28590,I28460,I28573);
nor I_1587 (I28237,I28590,I28313);
nand I_1588 (I28621,I28573,I28508);
nand I_1589 (I28222,I28330,I28621);
nand I_1590 (I28652,I28412,I28621);
DFFARX1 I_1591 (I28652,I1598,I28245,I28225,);
nand I_1592 (I28683,I28477,I28542);
nor I_1593 (I28219,I28330,I28683);
nor I_1594 (I28714,I28477,I28542);
nand I_1595 (I28228,I28714,I28525);
not I_1596 (I28772,I1605);
or I_1597 (I28789,I4243,I4243);
nand I_1598 (I28806,I4249,I4252);
not I_1599 (I28823,I28806);
nand I_1600 (I28840,I28823,I28789);
not I_1601 (I28857,I28840);
nand I_1602 (I28874,I4261,I4264);
and I_1603 (I28891,I28874,I4246);
DFFARX1 I_1604 (I28891,I1598,I28772,I28917,);
nor I_1605 (I28740,I28917,I28806);
nand I_1606 (I28939,I28857,I28917);
nor I_1607 (I28956,I28917,I28823);
not I_1608 (I28758,I28917);
nor I_1609 (I28987,I4258,I4264);
not I_1610 (I29004,I28987);
nand I_1611 (I28761,I28956,I28987);
not I_1612 (I29035,I4246);
nor I_1613 (I29052,I28917,I4246);
nand I_1614 (I29069,I4249,I4255);
nor I_1615 (I28743,I29069,I28806);
not I_1616 (I29100,I29069);
nor I_1617 (I29117,I28987,I29100);
nor I_1618 (I28764,I29117,I28840);
nand I_1619 (I29148,I29100,I29035);
nand I_1620 (I28749,I28857,I29148);
nand I_1621 (I29179,I28939,I29148);
DFFARX1 I_1622 (I29179,I1598,I28772,I28752,);
nand I_1623 (I29210,I29004,I29069);
nor I_1624 (I28746,I28857,I29210);
nor I_1625 (I29241,I29004,I29069);
nand I_1626 (I28755,I29241,I29052);
not I_1627 (I29299,I1605);
or I_1628 (I29316,I58168,I58156);
nand I_1629 (I29333,I58150,I58150);
not I_1630 (I29350,I29333);
nand I_1631 (I29367,I29350,I29316);
not I_1632 (I29384,I29367);
nand I_1633 (I29401,I58153,I58153);
and I_1634 (I29418,I29401,I58159);
DFFARX1 I_1635 (I29418,I1598,I29299,I29444,);
nor I_1636 (I29267,I29444,I29333);
nand I_1637 (I29466,I29384,I29444);
nor I_1638 (I29483,I29444,I29350);
not I_1639 (I29285,I29444);
nor I_1640 (I29514,I58165,I58153);
not I_1641 (I29531,I29514);
nand I_1642 (I29288,I29483,I29514);
not I_1643 (I29562,I58171);
nor I_1644 (I29579,I29444,I58171);
nand I_1645 (I29596,I58156,I58162);
nor I_1646 (I29270,I29596,I29333);
not I_1647 (I29627,I29596);
nor I_1648 (I29644,I29514,I29627);
nor I_1649 (I29291,I29644,I29367);
nand I_1650 (I29675,I29627,I29562);
nand I_1651 (I29276,I29384,I29675);
nand I_1652 (I29706,I29466,I29675);
DFFARX1 I_1653 (I29706,I1598,I29299,I29279,);
nand I_1654 (I29737,I29531,I29596);
nor I_1655 (I29273,I29384,I29737);
nor I_1656 (I29768,I29531,I29596);
nand I_1657 (I29282,I29768,I29579);
not I_1658 (I29826,I1605);
or I_1659 (I29843,I16044,I16041);
nand I_1660 (I29860,I16047,I16044);
not I_1661 (I29877,I29860);
nand I_1662 (I29894,I29877,I29843);
not I_1663 (I29911,I29894);
nand I_1664 (I29928,I16062,I16065);
and I_1665 (I29945,I29928,I16041);
DFFARX1 I_1666 (I29945,I1598,I29826,I29971,);
nor I_1667 (I29794,I29971,I29860);
nand I_1668 (I29993,I29911,I29971);
nor I_1669 (I30010,I29971,I29877);
not I_1670 (I29812,I29971);
nor I_1671 (I30041,I16059,I16065);
not I_1672 (I30058,I30041);
nand I_1673 (I29815,I30010,I30041);
not I_1674 (I30089,I16050);
nor I_1675 (I30106,I29971,I16050);
nand I_1676 (I30123,I16053,I16056);
nor I_1677 (I29797,I30123,I29860);
not I_1678 (I30154,I30123);
nor I_1679 (I30171,I30041,I30154);
nor I_1680 (I29818,I30171,I29894);
nand I_1681 (I30202,I30154,I30089);
nand I_1682 (I29803,I29911,I30202);
nand I_1683 (I30233,I29993,I30202);
DFFARX1 I_1684 (I30233,I1598,I29826,I29806,);
nand I_1685 (I30264,I30058,I30123);
nor I_1686 (I29800,I29911,I30264);
nor I_1687 (I30295,I30058,I30123);
nand I_1688 (I29809,I30295,I30106);
not I_1689 (I30353,I1605);
or I_1690 (I30370,I42357,I42360);
nand I_1691 (I30387,I42363,I42372);
not I_1692 (I30404,I30387);
nand I_1693 (I30421,I30404,I30370);
not I_1694 (I30438,I30421);
nand I_1695 (I30455,I42369,I42375);
and I_1696 (I30472,I30455,I42357);
DFFARX1 I_1697 (I30472,I1598,I30353,I30498,);
nor I_1698 (I30321,I30498,I30387);
nand I_1699 (I30520,I30438,I30498);
nor I_1700 (I30537,I30498,I30404);
not I_1701 (I30339,I30498);
nor I_1702 (I30568,I42360,I42375);
not I_1703 (I30585,I30568);
nand I_1704 (I30342,I30537,I30568);
not I_1705 (I30616,I42378);
nor I_1706 (I30633,I30498,I42378);
nand I_1707 (I30650,I42366,I42363);
nor I_1708 (I30324,I30650,I30387);
not I_1709 (I30681,I30650);
nor I_1710 (I30698,I30568,I30681);
nor I_1711 (I30345,I30698,I30421);
nand I_1712 (I30729,I30681,I30616);
nand I_1713 (I30330,I30438,I30729);
nand I_1714 (I30760,I30520,I30729);
DFFARX1 I_1715 (I30760,I1598,I30353,I30333,);
nand I_1716 (I30791,I30585,I30650);
nor I_1717 (I30327,I30438,I30791);
nor I_1718 (I30822,I30585,I30650);
nand I_1719 (I30336,I30822,I30633);
not I_1720 (I30880,I1605);
or I_1721 (I30897,I56063,I56051);
nand I_1722 (I30914,I56054,I56048);
not I_1723 (I30931,I30914);
nand I_1724 (I30948,I30931,I30897);
not I_1725 (I30965,I30948);
nand I_1726 (I30982,I56045,I56048);
and I_1727 (I30999,I30982,I56042);
DFFARX1 I_1728 (I30999,I1598,I30880,I31025,);
nor I_1729 (I30848,I31025,I30914);
nand I_1730 (I31047,I30965,I31025);
nor I_1731 (I31064,I31025,I30931);
not I_1732 (I30866,I31025);
nor I_1733 (I31095,I56042,I56048);
not I_1734 (I31112,I31095);
nand I_1735 (I30869,I31064,I31095);
not I_1736 (I31143,I56045);
nor I_1737 (I31160,I31025,I56045);
nand I_1738 (I31177,I56060,I56057);
nor I_1739 (I30851,I31177,I30914);
not I_1740 (I31208,I31177);
nor I_1741 (I31225,I31095,I31208);
nor I_1742 (I30872,I31225,I30948);
nand I_1743 (I31256,I31208,I31143);
nand I_1744 (I30857,I30965,I31256);
nand I_1745 (I31287,I31047,I31256);
DFFARX1 I_1746 (I31287,I1598,I30880,I30860,);
nand I_1747 (I31318,I31112,I31177);
nor I_1748 (I30854,I30965,I31318);
nor I_1749 (I31349,I31112,I31177);
nand I_1750 (I30863,I31349,I31160);
not I_1751 (I31407,I1605);
or I_1752 (I31424,I72946,I72943);
nand I_1753 (I31441,I72955,I72958);
not I_1754 (I31458,I31441);
nand I_1755 (I31475,I31458,I31424);
not I_1756 (I31492,I31475);
nand I_1757 (I31509,I72949,I72940);
and I_1758 (I31526,I31509,I72940);
DFFARX1 I_1759 (I31526,I1598,I31407,I31552,);
nor I_1760 (I31375,I31552,I31441);
nand I_1761 (I31574,I31492,I31552);
nor I_1762 (I31591,I31552,I31458);
not I_1763 (I31393,I31552);
nor I_1764 (I31622,I72943,I72940);
not I_1765 (I31639,I31622);
nand I_1766 (I31396,I31591,I31622);
not I_1767 (I31670,I72946);
nor I_1768 (I31687,I31552,I72946);
nand I_1769 (I31704,I72949,I72952);
nor I_1770 (I31378,I31704,I31441);
not I_1771 (I31735,I31704);
nor I_1772 (I31752,I31622,I31735);
nor I_1773 (I31399,I31752,I31475);
nand I_1774 (I31783,I31735,I31670);
nand I_1775 (I31384,I31492,I31783);
nand I_1776 (I31814,I31574,I31783);
DFFARX1 I_1777 (I31814,I1598,I31407,I31387,);
nand I_1778 (I31845,I31639,I31704);
nor I_1779 (I31381,I31492,I31845);
nor I_1780 (I31876,I31639,I31704);
nand I_1781 (I31390,I31876,I31687);
not I_1782 (I31934,I1605);
or I_1783 (I31951,I6864,I6861);
nand I_1784 (I31968,I6867,I6864);
not I_1785 (I31985,I31968);
nand I_1786 (I32002,I31985,I31951);
not I_1787 (I32019,I32002);
nand I_1788 (I32036,I6882,I6885);
and I_1789 (I32053,I32036,I6861);
DFFARX1 I_1790 (I32053,I1598,I31934,I32079,);
nor I_1791 (I31902,I32079,I31968);
nand I_1792 (I32101,I32019,I32079);
nor I_1793 (I32118,I32079,I31985);
not I_1794 (I31920,I32079);
nor I_1795 (I32149,I6879,I6885);
not I_1796 (I32166,I32149);
nand I_1797 (I31923,I32118,I32149);
not I_1798 (I32197,I6870);
nor I_1799 (I32214,I32079,I6870);
nand I_1800 (I32231,I6873,I6876);
nor I_1801 (I31905,I32231,I31968);
not I_1802 (I32262,I32231);
nor I_1803 (I32279,I32149,I32262);
nor I_1804 (I31926,I32279,I32002);
nand I_1805 (I32310,I32262,I32197);
nand I_1806 (I31911,I32019,I32310);
nand I_1807 (I32341,I32101,I32310);
DFFARX1 I_1808 (I32341,I1598,I31934,I31914,);
nand I_1809 (I32372,I32166,I32231);
nor I_1810 (I31908,I32019,I32372);
nor I_1811 (I32403,I32166,I32231);
nand I_1812 (I31917,I32403,I32214);
not I_1813 (I32461,I1605);
or I_1814 (I32478,I42833,I42836);
nand I_1815 (I32495,I42839,I42848);
not I_1816 (I32512,I32495);
nand I_1817 (I32529,I32512,I32478);
not I_1818 (I32546,I32529);
nand I_1819 (I32563,I42845,I42851);
and I_1820 (I32580,I32563,I42833);
DFFARX1 I_1821 (I32580,I1598,I32461,I32606,);
nor I_1822 (I32429,I32606,I32495);
nand I_1823 (I32628,I32546,I32606);
nor I_1824 (I32645,I32606,I32512);
not I_1825 (I32447,I32606);
nor I_1826 (I32676,I42836,I42851);
not I_1827 (I32693,I32676);
nand I_1828 (I32450,I32645,I32676);
not I_1829 (I32724,I42854);
nor I_1830 (I32741,I32606,I42854);
nand I_1831 (I32758,I42842,I42839);
nor I_1832 (I32432,I32758,I32495);
not I_1833 (I32789,I32758);
nor I_1834 (I32806,I32676,I32789);
nor I_1835 (I32453,I32806,I32529);
nand I_1836 (I32837,I32789,I32724);
nand I_1837 (I32438,I32546,I32837);
nand I_1838 (I32868,I32628,I32837);
DFFARX1 I_1839 (I32868,I1598,I32461,I32441,);
nand I_1840 (I32899,I32693,I32758);
nor I_1841 (I32435,I32546,I32899);
nor I_1842 (I32930,I32693,I32758);
nand I_1843 (I32444,I32930,I32741);
not I_1844 (I32988,I1605);
or I_1845 (I33005,I11454,I11451);
nand I_1846 (I33022,I11457,I11454);
not I_1847 (I33039,I33022);
nand I_1848 (I33056,I33039,I33005);
not I_1849 (I33073,I33056);
nand I_1850 (I33090,I11472,I11475);
and I_1851 (I33107,I33090,I11451);
DFFARX1 I_1852 (I33107,I1598,I32988,I33133,);
nor I_1853 (I32956,I33133,I33022);
nand I_1854 (I33155,I33073,I33133);
nor I_1855 (I33172,I33133,I33039);
not I_1856 (I32974,I33133);
nor I_1857 (I33203,I11469,I11475);
not I_1858 (I33220,I33203);
nand I_1859 (I32977,I33172,I33203);
not I_1860 (I33251,I11460);
nor I_1861 (I33268,I33133,I11460);
nand I_1862 (I33285,I11463,I11466);
nor I_1863 (I32959,I33285,I33022);
not I_1864 (I33316,I33285);
nor I_1865 (I33333,I33203,I33316);
nor I_1866 (I32980,I33333,I33056);
nand I_1867 (I33364,I33316,I33251);
nand I_1868 (I32965,I33073,I33364);
nand I_1869 (I33395,I33155,I33364);
DFFARX1 I_1870 (I33395,I1598,I32988,I32968,);
nand I_1871 (I33426,I33220,I33285);
nor I_1872 (I32962,I33073,I33426);
nor I_1873 (I33457,I33220,I33285);
nand I_1874 (I32971,I33457,I33268);
not I_1875 (I33515,I1605);
or I_1876 (I33532,I49497,I49500);
nand I_1877 (I33549,I49503,I49512);
not I_1878 (I33566,I33549);
nand I_1879 (I33583,I33566,I33532);
not I_1880 (I33600,I33583);
nand I_1881 (I33617,I49509,I49515);
and I_1882 (I33634,I33617,I49497);
DFFARX1 I_1883 (I33634,I1598,I33515,I33660,);
nor I_1884 (I33483,I33660,I33549);
nand I_1885 (I33682,I33600,I33660);
nor I_1886 (I33699,I33660,I33566);
not I_1887 (I33501,I33660);
nor I_1888 (I33730,I49500,I49515);
not I_1889 (I33747,I33730);
nand I_1890 (I33504,I33699,I33730);
not I_1891 (I33778,I49518);
nor I_1892 (I33795,I33660,I49518);
nand I_1893 (I33812,I49506,I49503);
nor I_1894 (I33486,I33812,I33549);
not I_1895 (I33843,I33812);
nor I_1896 (I33860,I33730,I33843);
nor I_1897 (I33507,I33860,I33583);
nand I_1898 (I33891,I33843,I33778);
nand I_1899 (I33492,I33600,I33891);
nand I_1900 (I33922,I33682,I33891);
DFFARX1 I_1901 (I33922,I1598,I33515,I33495,);
nand I_1902 (I33953,I33747,I33812);
nor I_1903 (I33489,I33600,I33953);
nor I_1904 (I33984,I33747,I33812);
nand I_1905 (I33498,I33984,I33795);
not I_1906 (I34042,I1605);
or I_1907 (I34059,I50925,I50928);
nand I_1908 (I34076,I50931,I50940);
not I_1909 (I34093,I34076);
nand I_1910 (I34110,I34093,I34059);
not I_1911 (I34127,I34110);
nand I_1912 (I34144,I50937,I50943);
and I_1913 (I34161,I34144,I50925);
DFFARX1 I_1914 (I34161,I1598,I34042,I34187,);
nor I_1915 (I34010,I34187,I34076);
nand I_1916 (I34209,I34127,I34187);
nor I_1917 (I34226,I34187,I34093);
not I_1918 (I34028,I34187);
nor I_1919 (I34257,I50928,I50943);
not I_1920 (I34274,I34257);
nand I_1921 (I34031,I34226,I34257);
not I_1922 (I34305,I50946);
nor I_1923 (I34322,I34187,I50946);
nand I_1924 (I34339,I50934,I50931);
nor I_1925 (I34013,I34339,I34076);
not I_1926 (I34370,I34339);
nor I_1927 (I34387,I34257,I34370);
nor I_1928 (I34034,I34387,I34110);
nand I_1929 (I34418,I34370,I34305);
nand I_1930 (I34019,I34127,I34418);
nand I_1931 (I34449,I34209,I34418);
DFFARX1 I_1932 (I34449,I1598,I34042,I34022,);
nand I_1933 (I34480,I34274,I34339);
nor I_1934 (I34016,I34127,I34480);
nor I_1935 (I34511,I34274,I34339);
nand I_1936 (I34025,I34511,I34322);
not I_1937 (I34569,I1605);
or I_1938 (I34586,I66600,I66588);
nand I_1939 (I34603,I66582,I66582);
not I_1940 (I34620,I34603);
nand I_1941 (I34637,I34620,I34586);
not I_1942 (I34654,I34637);
nand I_1943 (I34671,I66585,I66585);
and I_1944 (I34688,I34671,I66591);
DFFARX1 I_1945 (I34688,I1598,I34569,I34714,);
nor I_1946 (I34537,I34714,I34603);
nand I_1947 (I34736,I34654,I34714);
nor I_1948 (I34753,I34714,I34620);
not I_1949 (I34555,I34714);
nor I_1950 (I34784,I66597,I66585);
not I_1951 (I34801,I34784);
nand I_1952 (I34558,I34753,I34784);
not I_1953 (I34832,I66603);
nor I_1954 (I34849,I34714,I66603);
nand I_1955 (I34866,I66588,I66594);
nor I_1956 (I34540,I34866,I34603);
not I_1957 (I34897,I34866);
nor I_1958 (I34914,I34784,I34897);
nor I_1959 (I34561,I34914,I34637);
nand I_1960 (I34945,I34897,I34832);
nand I_1961 (I34546,I34654,I34945);
nand I_1962 (I34976,I34736,I34945);
DFFARX1 I_1963 (I34976,I1598,I34569,I34549,);
nand I_1964 (I35007,I34801,I34866);
nor I_1965 (I34543,I34654,I35007);
nor I_1966 (I35038,I34801,I34866);
nand I_1967 (I34552,I35038,I34849);
not I_1968 (I35096,I1605);
or I_1969 (I35113,I1287,I1463);
nand I_1970 (I35130,I1159,I999);
not I_1971 (I35147,I35130);
nand I_1972 (I35164,I35147,I35113);
not I_1973 (I35181,I35164);
nand I_1974 (I35198,I1247,I1303);
and I_1975 (I35215,I35198,I1407);
DFFARX1 I_1976 (I35215,I1598,I35096,I35241,);
nor I_1977 (I35064,I35241,I35130);
nand I_1978 (I35263,I35181,I35241);
nor I_1979 (I35280,I35241,I35147);
not I_1980 (I35082,I35241);
nor I_1981 (I35311,I807,I1303);
not I_1982 (I35328,I35311);
nand I_1983 (I35085,I35280,I35311);
not I_1984 (I35359,I1279);
nor I_1985 (I35376,I35241,I1279);
nand I_1986 (I35393,I711,I1351);
nor I_1987 (I35067,I35393,I35130);
not I_1988 (I35424,I35393);
nor I_1989 (I35441,I35311,I35424);
nor I_1990 (I35088,I35441,I35164);
nand I_1991 (I35472,I35424,I35359);
nand I_1992 (I35073,I35181,I35472);
nand I_1993 (I35503,I35263,I35472);
DFFARX1 I_1994 (I35503,I1598,I35096,I35076,);
nand I_1995 (I35534,I35328,I35393);
nor I_1996 (I35070,I35181,I35534);
nor I_1997 (I35565,I35328,I35393);
nand I_1998 (I35079,I35565,I35376);
not I_1999 (I35623,I1605);
or I_2000 (I35640,I50449,I50452);
nand I_2001 (I35657,I50455,I50464);
not I_2002 (I35674,I35657);
nand I_2003 (I35691,I35674,I35640);
not I_2004 (I35708,I35691);
nand I_2005 (I35725,I50461,I50467);
and I_2006 (I35742,I35725,I50449);
DFFARX1 I_2007 (I35742,I1598,I35623,I35768,);
nor I_2008 (I35591,I35768,I35657);
nand I_2009 (I35790,I35708,I35768);
nor I_2010 (I35807,I35768,I35674);
not I_2011 (I35609,I35768);
nor I_2012 (I35838,I50452,I50467);
not I_2013 (I35855,I35838);
nand I_2014 (I35612,I35807,I35838);
not I_2015 (I35886,I50470);
nor I_2016 (I35903,I35768,I50470);
nand I_2017 (I35920,I50458,I50455);
nor I_2018 (I35594,I35920,I35657);
not I_2019 (I35951,I35920);
nor I_2020 (I35968,I35838,I35951);
nor I_2021 (I35615,I35968,I35691);
nand I_2022 (I35999,I35951,I35886);
nand I_2023 (I35600,I35708,I35999);
nand I_2024 (I36030,I35790,I35999);
DFFARX1 I_2025 (I36030,I1598,I35623,I35603,);
nand I_2026 (I36061,I35855,I35920);
nor I_2027 (I35597,I35708,I36061);
nor I_2028 (I36092,I35855,I35920);
nand I_2029 (I35606,I36092,I35903);
not I_2030 (I36150,I1605);
or I_2031 (I36167,I1471,I1015);
nand I_2032 (I36184,I911,I919);
not I_2033 (I36201,I36184);
nand I_2034 (I36218,I36201,I36167);
not I_2035 (I36235,I36218);
nand I_2036 (I36252,I1239,I1479);
and I_2037 (I36269,I36252,I759);
DFFARX1 I_2038 (I36269,I1598,I36150,I36295,);
nor I_2039 (I36118,I36295,I36184);
nand I_2040 (I36317,I36235,I36295);
nor I_2041 (I36334,I36295,I36201);
not I_2042 (I36136,I36295);
nor I_2043 (I36365,I1103,I1479);
not I_2044 (I36382,I36365);
nand I_2045 (I36139,I36334,I36365);
not I_2046 (I36413,I1223);
nor I_2047 (I36430,I36295,I1223);
nand I_2048 (I36447,I1127,I1135);
nor I_2049 (I36121,I36447,I36184);
not I_2050 (I36478,I36447);
nor I_2051 (I36495,I36365,I36478);
nor I_2052 (I36142,I36495,I36218);
nand I_2053 (I36526,I36478,I36413);
nand I_2054 (I36127,I36235,I36526);
nand I_2055 (I36557,I36317,I36526);
DFFARX1 I_2056 (I36557,I1598,I36150,I36130,);
nand I_2057 (I36588,I36382,I36447);
nor I_2058 (I36124,I36235,I36588);
nor I_2059 (I36619,I36382,I36447);
nand I_2060 (I36133,I36619,I36430);
not I_2061 (I36674,I1605);
or I_2062 (I36691,I24021,I24006);
nor I_2063 (I36708,I36691,I24000);
nor I_2064 (I36725,I23997,I24018);
or I_2065 (I36742,I36725,I24015);
nor I_2066 (I36759,I24003,I24000);
nand I_2067 (I36776,I36759,I36742);
not I_2068 (I36793,I36776);
nand I_2069 (I36810,I36708,I36793);
nor I_2070 (I36827,I36708,I36793);
nand I_2071 (I36844,I24009,I24012);
nor I_2072 (I36861,I36844,I23997);
nor I_2073 (I36878,I36844,I36861);
not I_2074 (I36895,I36861);
nor I_2075 (I36666,I36895,I36810);
or I_2076 (I36651,I36708,I36895);
nor I_2077 (I36940,I36708,I36861);
nor I_2078 (I36645,I36844,I36940);
nor I_2079 (I36971,I36878,I36940);
nor I_2080 (I36648,I36793,I36971);
nand I_2081 (I37002,I36708,I36861);
nand I_2082 (I37019,I36776,I37002);
DFFARX1 I_2083 (I37019,I1598,I36674,I36654,);
not I_2084 (I37050,I36844);
nor I_2085 (I36663,I37050,I36895);
nand I_2086 (I36660,I36827,I37050);
nor I_2087 (I37095,I36793,I36844);
nand I_2088 (I36657,I37095,I36708);
not I_2089 (I37150,I1605);
or I_2090 (I37167,I73385,I73388);
nor I_2091 (I37184,I37167,I73385);
nor I_2092 (I37201,I73382,I73400);
or I_2093 (I37218,I37201,I73388);
nor I_2094 (I37235,I73391,I73382);
nand I_2095 (I37252,I37235,I37218);
not I_2096 (I37269,I37252);
nand I_2097 (I37286,I37184,I37269);
nor I_2098 (I37303,I37184,I37269);
nand I_2099 (I37320,I73397,I73394);
nor I_2100 (I37337,I37320,I73391);
nor I_2101 (I37354,I37320,I37337);
not I_2102 (I37371,I37337);
nor I_2103 (I37142,I37371,I37286);
or I_2104 (I37127,I37184,I37371);
nor I_2105 (I37416,I37184,I37337);
nor I_2106 (I37121,I37320,I37416);
nor I_2107 (I37447,I37354,I37416);
nor I_2108 (I37124,I37269,I37447);
nand I_2109 (I37478,I37184,I37337);
nand I_2110 (I37495,I37252,I37478);
DFFARX1 I_2111 (I37495,I1598,I37150,I37130,);
not I_2112 (I37526,I37320);
nor I_2113 (I37139,I37526,I37371);
nand I_2114 (I37136,I37303,I37526);
nor I_2115 (I37571,I37269,I37320);
nand I_2116 (I37133,I37571,I37184);
not I_2117 (I37626,I1605);
or I_2118 (I37643,I56569,I56590);
nor I_2119 (I37660,I37643,I56575);
nor I_2120 (I37677,I56569,I56587);
or I_2121 (I37694,I37677,I56578);
nor I_2122 (I37711,I56572,I56572);
nand I_2123 (I37728,I37711,I37694);
not I_2124 (I37745,I37728);
nand I_2125 (I37762,I37660,I37745);
nor I_2126 (I37779,I37660,I37745);
nand I_2127 (I37796,I56581,I56584);
nor I_2128 (I37813,I37796,I56575);
nor I_2129 (I37830,I37796,I37813);
not I_2130 (I37847,I37813);
nor I_2131 (I37618,I37847,I37762);
or I_2132 (I37603,I37660,I37847);
nor I_2133 (I37892,I37660,I37813);
nor I_2134 (I37597,I37796,I37892);
nor I_2135 (I37923,I37830,I37892);
nor I_2136 (I37600,I37745,I37923);
nand I_2137 (I37954,I37660,I37813);
nand I_2138 (I37971,I37728,I37954);
DFFARX1 I_2139 (I37971,I1598,I37626,I37606,);
not I_2140 (I38002,I37796);
nor I_2141 (I37615,I38002,I37847);
nand I_2142 (I37612,I37779,I38002);
nor I_2143 (I38047,I37745,I37796);
nand I_2144 (I37609,I38047,I37660);
not I_2145 (I38102,I1605);
or I_2146 (I38119,I23184,I23181);
nor I_2147 (I38136,I38119,I23181);
nor I_2148 (I38153,I23190,I23187);
or I_2149 (I38170,I38153,I23196);
nor I_2150 (I38187,I23199,I23184);
nand I_2151 (I38204,I38187,I38170);
not I_2152 (I38221,I38204);
nand I_2153 (I38238,I38136,I38221);
nor I_2154 (I38255,I38136,I38221);
nand I_2155 (I38272,I23187,I23193);
nor I_2156 (I38289,I38272,I23190);
nor I_2157 (I38306,I38272,I38289);
not I_2158 (I38323,I38289);
nor I_2159 (I38094,I38323,I38238);
or I_2160 (I38079,I38136,I38323);
nor I_2161 (I38368,I38136,I38289);
nor I_2162 (I38073,I38272,I38368);
nor I_2163 (I38399,I38306,I38368);
nor I_2164 (I38076,I38221,I38399);
nand I_2165 (I38430,I38136,I38289);
nand I_2166 (I38447,I38204,I38430);
DFFARX1 I_2167 (I38447,I1598,I38102,I38082,);
not I_2168 (I38478,I38272);
nor I_2169 (I38091,I38478,I38323);
nand I_2170 (I38088,I38255,I38478);
nor I_2171 (I38523,I38221,I38272);
nand I_2172 (I38085,I38523,I38136);
not I_2173 (I38578,I1605);
or I_2174 (I38595,I10431,I10440);
nor I_2175 (I38612,I38595,I10455);
nor I_2176 (I38629,I10452,I10434);
or I_2177 (I38646,I38629,I10434);
nor I_2178 (I38663,I10431,I10437);
nand I_2179 (I38680,I38663,I38646);
not I_2180 (I38697,I38680);
nand I_2181 (I38714,I38612,I38697);
nor I_2182 (I38731,I38612,I38697);
nand I_2183 (I38748,I10443,I10446);
nor I_2184 (I38765,I38748,I10449);
nor I_2185 (I38782,I38748,I38765);
not I_2186 (I38799,I38765);
nor I_2187 (I38570,I38799,I38714);
or I_2188 (I38555,I38612,I38799);
nor I_2189 (I38844,I38612,I38765);
nor I_2190 (I38549,I38748,I38844);
nor I_2191 (I38875,I38782,I38844);
nor I_2192 (I38552,I38697,I38875);
nand I_2193 (I38906,I38612,I38765);
nand I_2194 (I38923,I38680,I38906);
DFFARX1 I_2195 (I38923,I1598,I38578,I38558,);
not I_2196 (I38954,I38748);
nor I_2197 (I38567,I38954,I38799);
nand I_2198 (I38564,I38731,I38954);
nor I_2199 (I38999,I38697,I38748);
nand I_2200 (I38561,I38999,I38612);
not I_2201 (I39054,I1605);
or I_2202 (I39071,I20631,I20640);
nor I_2203 (I39088,I39071,I20655);
nor I_2204 (I39105,I20652,I20634);
or I_2205 (I39122,I39105,I20634);
nor I_2206 (I39139,I20631,I20637);
nand I_2207 (I39156,I39139,I39122);
not I_2208 (I39173,I39156);
nand I_2209 (I39190,I39088,I39173);
nor I_2210 (I39207,I39088,I39173);
nand I_2211 (I39224,I20643,I20646);
nor I_2212 (I39241,I39224,I20649);
nor I_2213 (I39258,I39224,I39241);
not I_2214 (I39275,I39241);
nor I_2215 (I39046,I39275,I39190);
or I_2216 (I39031,I39088,I39275);
nor I_2217 (I39320,I39088,I39241);
nor I_2218 (I39025,I39224,I39320);
nor I_2219 (I39351,I39258,I39320);
nor I_2220 (I39028,I39173,I39351);
nand I_2221 (I39382,I39088,I39241);
nand I_2222 (I39399,I39156,I39382);
DFFARX1 I_2223 (I39399,I1598,I39054,I39034,);
not I_2224 (I39430,I39224);
nor I_2225 (I39043,I39430,I39275);
nand I_2226 (I39040,I39207,I39430);
nor I_2227 (I39475,I39173,I39224);
nand I_2228 (I39037,I39475,I39088);
not I_2229 (I39530,I1605);
or I_2230 (I39547,I1527,I815);
nor I_2231 (I39564,I39547,I1591);
nor I_2232 (I39581,I1487,I1439);
or I_2233 (I39598,I39581,I879);
nor I_2234 (I39615,I735,I847);
nand I_2235 (I39632,I39615,I39598);
not I_2236 (I39649,I39632);
nand I_2237 (I39666,I39564,I39649);
nor I_2238 (I39683,I39564,I39649);
nand I_2239 (I39700,I975,I1503);
nor I_2240 (I39717,I39700,I791);
nor I_2241 (I39734,I39700,I39717);
not I_2242 (I39751,I39717);
nor I_2243 (I39522,I39751,I39666);
or I_2244 (I39507,I39564,I39751);
nor I_2245 (I39796,I39564,I39717);
nor I_2246 (I39501,I39700,I39796);
nor I_2247 (I39827,I39734,I39796);
nor I_2248 (I39504,I39649,I39827);
nand I_2249 (I39858,I39564,I39717);
nand I_2250 (I39875,I39632,I39858);
DFFARX1 I_2251 (I39875,I1598,I39530,I39510,);
not I_2252 (I39906,I39700);
nor I_2253 (I39519,I39906,I39751);
nand I_2254 (I39516,I39683,I39906);
nor I_2255 (I39951,I39649,I39700);
nand I_2256 (I39513,I39951,I39564);
not I_2257 (I40006,I1605);
or I_2258 (I40023,I60785,I60806);
nor I_2259 (I40040,I40023,I60791);
nor I_2260 (I40057,I60785,I60803);
or I_2261 (I40074,I40057,I60794);
nor I_2262 (I40091,I60788,I60788);
nand I_2263 (I40108,I40091,I40074);
not I_2264 (I40125,I40108);
nand I_2265 (I40142,I40040,I40125);
nor I_2266 (I40159,I40040,I40125);
nand I_2267 (I40176,I60797,I60800);
nor I_2268 (I40193,I40176,I60791);
nor I_2269 (I40210,I40176,I40193);
not I_2270 (I40227,I40193);
nor I_2271 (I39998,I40227,I40142);
or I_2272 (I39983,I40040,I40227);
nor I_2273 (I40272,I40040,I40193);
nor I_2274 (I39977,I40176,I40272);
nor I_2275 (I40303,I40210,I40272);
nor I_2276 (I39980,I40125,I40303);
nand I_2277 (I40334,I40040,I40193);
nand I_2278 (I40351,I40108,I40334);
DFFARX1 I_2279 (I40351,I1598,I40006,I39986,);
not I_2280 (I40382,I40176);
nor I_2281 (I39995,I40382,I40227);
nand I_2282 (I39992,I40159,I40382);
nor I_2283 (I40427,I40125,I40176);
nand I_2284 (I39989,I40427,I40040);
not I_2285 (I40482,I1605);
or I_2286 (I40499,I31926,I31911);
nor I_2287 (I40516,I40499,I31905);
nor I_2288 (I40533,I31902,I31923);
or I_2289 (I40550,I40533,I31920);
nor I_2290 (I40567,I31908,I31905);
nand I_2291 (I40584,I40567,I40550);
not I_2292 (I40601,I40584);
nand I_2293 (I40618,I40516,I40601);
nor I_2294 (I40635,I40516,I40601);
nand I_2295 (I40652,I31914,I31917);
nor I_2296 (I40669,I40652,I31902);
nor I_2297 (I40686,I40652,I40669);
not I_2298 (I40703,I40669);
nor I_2299 (I40474,I40703,I40618);
or I_2300 (I40459,I40516,I40703);
nor I_2301 (I40748,I40516,I40669);
nor I_2302 (I40453,I40652,I40748);
nor I_2303 (I40779,I40686,I40748);
nor I_2304 (I40456,I40601,I40779);
nand I_2305 (I40810,I40516,I40669);
nand I_2306 (I40827,I40584,I40810);
DFFARX1 I_2307 (I40827,I1598,I40482,I40462,);
not I_2308 (I40858,I40652);
nor I_2309 (I40471,I40858,I40703);
nand I_2310 (I40468,I40635,I40858);
nor I_2311 (I40903,I40601,I40652);
nand I_2312 (I40465,I40903,I40516);
not I_2313 (I40958,I1605);
or I_2314 (I40975,I21552,I21549);
nor I_2315 (I40992,I40975,I21549);
nor I_2316 (I41009,I21558,I21555);
or I_2317 (I41026,I41009,I21564);
nor I_2318 (I41043,I21567,I21552);
nand I_2319 (I41060,I41043,I41026);
not I_2320 (I41077,I41060);
nand I_2321 (I41094,I40992,I41077);
nor I_2322 (I41111,I40992,I41077);
nand I_2323 (I41128,I21555,I21561);
nor I_2324 (I41145,I41128,I21558);
nor I_2325 (I41162,I41128,I41145);
not I_2326 (I41179,I41145);
nor I_2327 (I40950,I41179,I41094);
or I_2328 (I40935,I40992,I41179);
nor I_2329 (I41224,I40992,I41145);
nor I_2330 (I40929,I41128,I41224);
nor I_2331 (I41255,I41162,I41224);
nor I_2332 (I40932,I41077,I41255);
nand I_2333 (I41286,I40992,I41145);
nand I_2334 (I41303,I41060,I41286);
DFFARX1 I_2335 (I41303,I1598,I40958,I40938,);
not I_2336 (I41334,I41128);
nor I_2337 (I40947,I41334,I41179);
nand I_2338 (I40944,I41111,I41334);
nor I_2339 (I41379,I41077,I41128);
nand I_2340 (I40941,I41379,I40992);
not I_2341 (I41434,I1605);
or I_2342 (I41451,I18591,I18600);
nor I_2343 (I41468,I41451,I18615);
nor I_2344 (I41485,I18612,I18594);
or I_2345 (I41502,I41485,I18594);
nor I_2346 (I41519,I18591,I18597);
nand I_2347 (I41536,I41519,I41502);
not I_2348 (I41553,I41536);
nand I_2349 (I41570,I41468,I41553);
nor I_2350 (I41587,I41468,I41553);
nand I_2351 (I41604,I18603,I18606);
nor I_2352 (I41621,I41604,I18609);
nor I_2353 (I41638,I41604,I41621);
not I_2354 (I41655,I41621);
nor I_2355 (I41426,I41655,I41570);
or I_2356 (I41411,I41468,I41655);
nor I_2357 (I41700,I41468,I41621);
nor I_2358 (I41405,I41604,I41700);
nor I_2359 (I41731,I41638,I41700);
nor I_2360 (I41408,I41553,I41731);
nand I_2361 (I41762,I41468,I41621);
nand I_2362 (I41779,I41536,I41762);
DFFARX1 I_2363 (I41779,I1598,I41434,I41414,);
not I_2364 (I41810,I41604);
nor I_2365 (I41423,I41810,I41655);
nand I_2366 (I41420,I41587,I41810);
nor I_2367 (I41855,I41553,I41604);
nand I_2368 (I41417,I41855,I41468);
not I_2369 (I41910,I1605);
or I_2370 (I41927,I14001,I14010);
nor I_2371 (I41944,I41927,I14025);
nor I_2372 (I41961,I14022,I14004);
or I_2373 (I41978,I41961,I14004);
nor I_2374 (I41995,I14001,I14007);
nand I_2375 (I42012,I41995,I41978);
not I_2376 (I42029,I42012);
nand I_2377 (I42046,I41944,I42029);
nor I_2378 (I42063,I41944,I42029);
nand I_2379 (I42080,I14013,I14016);
nor I_2380 (I42097,I42080,I14019);
nor I_2381 (I42114,I42080,I42097);
not I_2382 (I42131,I42097);
nor I_2383 (I41902,I42131,I42046);
or I_2384 (I41887,I41944,I42131);
nor I_2385 (I42176,I41944,I42097);
nor I_2386 (I41881,I42080,I42176);
nor I_2387 (I42207,I42114,I42176);
nor I_2388 (I41884,I42029,I42207);
nand I_2389 (I42238,I41944,I42097);
nand I_2390 (I42255,I42012,I42238);
DFFARX1 I_2391 (I42255,I1598,I41910,I41890,);
not I_2392 (I42286,I42080);
nor I_2393 (I41899,I42286,I42131);
nand I_2394 (I41896,I42063,I42286);
nor I_2395 (I42331,I42029,I42080);
nand I_2396 (I41893,I42331,I41944);
not I_2397 (I42386,I1605);
or I_2398 (I42403,I29291,I29276);
nor I_2399 (I42420,I42403,I29270);
nor I_2400 (I42437,I29267,I29288);
or I_2401 (I42454,I42437,I29285);
nor I_2402 (I42471,I29273,I29270);
nand I_2403 (I42488,I42471,I42454);
not I_2404 (I42505,I42488);
nand I_2405 (I42522,I42420,I42505);
nor I_2406 (I42539,I42420,I42505);
nand I_2407 (I42556,I29279,I29282);
nor I_2408 (I42573,I42556,I29267);
nor I_2409 (I42590,I42556,I42573);
not I_2410 (I42607,I42573);
nor I_2411 (I42378,I42607,I42522);
or I_2412 (I42363,I42420,I42607);
nor I_2413 (I42652,I42420,I42573);
nor I_2414 (I42357,I42556,I42652);
nor I_2415 (I42683,I42590,I42652);
nor I_2416 (I42360,I42505,I42683);
nand I_2417 (I42714,I42420,I42573);
nand I_2418 (I42731,I42488,I42714);
DFFARX1 I_2419 (I42731,I1598,I42386,I42366,);
not I_2420 (I42762,I42556);
nor I_2421 (I42375,I42762,I42607);
nand I_2422 (I42372,I42539,I42762);
nor I_2423 (I42807,I42505,I42556);
nand I_2424 (I42369,I42807,I42420);
not I_2425 (I42862,I1605);
or I_2426 (I42879,I72059,I72062);
nor I_2427 (I42896,I42879,I72059);
nor I_2428 (I42913,I72056,I72074);
or I_2429 (I42930,I42913,I72062);
nor I_2430 (I42947,I72065,I72056);
nand I_2431 (I42964,I42947,I42930);
not I_2432 (I42981,I42964);
nand I_2433 (I42998,I42896,I42981);
nor I_2434 (I43015,I42896,I42981);
nand I_2435 (I43032,I72071,I72068);
nor I_2436 (I43049,I43032,I72065);
nor I_2437 (I43066,I43032,I43049);
not I_2438 (I43083,I43049);
nor I_2439 (I42854,I43083,I42998);
or I_2440 (I42839,I42896,I43083);
nor I_2441 (I43128,I42896,I43049);
nor I_2442 (I42833,I43032,I43128);
nor I_2443 (I43159,I43066,I43128);
nor I_2444 (I42836,I42981,I43159);
nand I_2445 (I43190,I42896,I43049);
nand I_2446 (I43207,I42964,I43190);
DFFARX1 I_2447 (I43207,I1598,I42862,I42842,);
not I_2448 (I43238,I43032);
nor I_2449 (I42851,I43238,I43083);
nand I_2450 (I42848,I43015,I43238);
nor I_2451 (I43283,I42981,I43032);
nand I_2452 (I42845,I43283,I42896);
not I_2453 (I43338,I1605);
or I_2454 (I43355,I66055,I66076);
nor I_2455 (I43372,I43355,I66061);
nor I_2456 (I43389,I66055,I66073);
or I_2457 (I43406,I43389,I66064);
nor I_2458 (I43423,I66058,I66058);
nand I_2459 (I43440,I43423,I43406);
not I_2460 (I43457,I43440);
nand I_2461 (I43474,I43372,I43457);
nor I_2462 (I43491,I43372,I43457);
nand I_2463 (I43508,I66067,I66070);
nor I_2464 (I43525,I43508,I66061);
nor I_2465 (I43542,I43508,I43525);
not I_2466 (I43559,I43525);
nor I_2467 (I43330,I43559,I43474);
or I_2468 (I43315,I43372,I43559);
nor I_2469 (I43604,I43372,I43525);
nor I_2470 (I43309,I43508,I43604);
nor I_2471 (I43635,I43542,I43604);
nor I_2472 (I43312,I43457,I43635);
nand I_2473 (I43666,I43372,I43525);
nand I_2474 (I43683,I43440,I43666);
DFFARX1 I_2475 (I43683,I1598,I43338,I43318,);
not I_2476 (I43714,I43508);
nor I_2477 (I43327,I43714,I43559);
nand I_2478 (I43324,I43491,I43714);
nor I_2479 (I43759,I43457,I43508);
nand I_2480 (I43321,I43759,I43372);
not I_2481 (I43814,I1605);
or I_2482 (I43831,I76037,I76040);
nor I_2483 (I43848,I43831,I76037);
nor I_2484 (I43865,I76034,I76052);
or I_2485 (I43882,I43865,I76040);
nor I_2486 (I43899,I76043,I76034);
nand I_2487 (I43916,I43899,I43882);
not I_2488 (I43933,I43916);
nand I_2489 (I43950,I43848,I43933);
nor I_2490 (I43967,I43848,I43933);
nand I_2491 (I43984,I76049,I76046);
nor I_2492 (I44001,I43984,I76043);
nor I_2493 (I44018,I43984,I44001);
not I_2494 (I44035,I44001);
nor I_2495 (I43806,I44035,I43950);
or I_2496 (I43791,I43848,I44035);
nor I_2497 (I44080,I43848,I44001);
nor I_2498 (I43785,I43984,I44080);
nor I_2499 (I44111,I44018,I44080);
nor I_2500 (I43788,I43933,I44111);
nand I_2501 (I44142,I43848,I44001);
nand I_2502 (I44159,I43916,I44142);
DFFARX1 I_2503 (I44159,I1598,I43814,I43794,);
not I_2504 (I44190,I43984);
nor I_2505 (I43803,I44190,I44035);
nand I_2506 (I43800,I43967,I44190);
nor I_2507 (I44235,I43933,I43984);
nand I_2508 (I43797,I44235,I43848);
not I_2509 (I44290,I1605);
or I_2510 (I44307,I12471,I12480);
nor I_2511 (I44324,I44307,I12495);
nor I_2512 (I44341,I12492,I12474);
or I_2513 (I44358,I44341,I12474);
nor I_2514 (I44375,I12471,I12477);
nand I_2515 (I44392,I44375,I44358);
not I_2516 (I44409,I44392);
nand I_2517 (I44426,I44324,I44409);
nor I_2518 (I44443,I44324,I44409);
nand I_2519 (I44460,I12483,I12486);
nor I_2520 (I44477,I44460,I12489);
nor I_2521 (I44494,I44460,I44477);
not I_2522 (I44511,I44477);
nor I_2523 (I44282,I44511,I44426);
or I_2524 (I44267,I44324,I44511);
nor I_2525 (I44556,I44324,I44477);
nor I_2526 (I44261,I44460,I44556);
nor I_2527 (I44587,I44494,I44556);
nor I_2528 (I44264,I44409,I44587);
nand I_2529 (I44618,I44324,I44477);
nand I_2530 (I44635,I44392,I44618);
DFFARX1 I_2531 (I44635,I1598,I44290,I44270,);
not I_2532 (I44666,I44460);
nor I_2533 (I44279,I44666,I44511);
nand I_2534 (I44276,I44443,I44666);
nor I_2535 (I44711,I44409,I44460);
nand I_2536 (I44273,I44711,I44324);
not I_2537 (I44766,I1605);
or I_2538 (I44783,I75595,I75598);
nor I_2539 (I44800,I44783,I75595);
nor I_2540 (I44817,I75592,I75610);
or I_2541 (I44834,I44817,I75598);
nor I_2542 (I44851,I75601,I75592);
nand I_2543 (I44868,I44851,I44834);
not I_2544 (I44885,I44868);
nand I_2545 (I44902,I44800,I44885);
nor I_2546 (I44919,I44800,I44885);
nand I_2547 (I44936,I75607,I75604);
nor I_2548 (I44953,I44936,I75601);
nor I_2549 (I44970,I44936,I44953);
not I_2550 (I44987,I44953);
nor I_2551 (I44758,I44987,I44902);
or I_2552 (I44743,I44800,I44987);
nor I_2553 (I45032,I44800,I44953);
nor I_2554 (I44737,I44936,I45032);
nor I_2555 (I45063,I44970,I45032);
nor I_2556 (I44740,I44885,I45063);
nand I_2557 (I45094,I44800,I44953);
nand I_2558 (I45111,I44868,I45094);
DFFARX1 I_2559 (I45111,I1598,I44766,I44746,);
not I_2560 (I45142,I44936);
nor I_2561 (I44755,I45142,I44987);
nand I_2562 (I44752,I44919,I45142);
nor I_2563 (I45187,I44885,I44936);
nand I_2564 (I44749,I45187,I44800);
not I_2565 (I45242,I1605);
or I_2566 (I45259,I17061,I17070);
nor I_2567 (I45276,I45259,I17085);
nor I_2568 (I45293,I17082,I17064);
or I_2569 (I45310,I45293,I17064);
nor I_2570 (I45327,I17061,I17067);
nand I_2571 (I45344,I45327,I45310);
not I_2572 (I45361,I45344);
nand I_2573 (I45378,I45276,I45361);
nor I_2574 (I45395,I45276,I45361);
nand I_2575 (I45412,I17073,I17076);
nor I_2576 (I45429,I45412,I17079);
nor I_2577 (I45446,I45412,I45429);
not I_2578 (I45463,I45429);
nor I_2579 (I45234,I45463,I45378);
or I_2580 (I45219,I45276,I45463);
nor I_2581 (I45508,I45276,I45429);
nor I_2582 (I45213,I45412,I45508);
nor I_2583 (I45539,I45446,I45508);
nor I_2584 (I45216,I45361,I45539);
nand I_2585 (I45570,I45276,I45429);
nand I_2586 (I45587,I45344,I45570);
DFFARX1 I_2587 (I45587,I1598,I45242,I45222,);
not I_2588 (I45618,I45412);
nor I_2589 (I45231,I45618,I45463);
nand I_2590 (I45228,I45395,I45618);
nor I_2591 (I45663,I45361,I45412);
nand I_2592 (I45225,I45663,I45276);
not I_2593 (I45718,I1605);
or I_2594 (I45735,I11961,I11970);
nor I_2595 (I45752,I45735,I11985);
nor I_2596 (I45769,I11982,I11964);
or I_2597 (I45786,I45769,I11964);
nor I_2598 (I45803,I11961,I11967);
nand I_2599 (I45820,I45803,I45786);
not I_2600 (I45837,I45820);
nand I_2601 (I45854,I45752,I45837);
nor I_2602 (I45871,I45752,I45837);
nand I_2603 (I45888,I11973,I11976);
nor I_2604 (I45905,I45888,I11979);
nor I_2605 (I45922,I45888,I45905);
not I_2606 (I45939,I45905);
nor I_2607 (I45710,I45939,I45854);
or I_2608 (I45695,I45752,I45939);
nor I_2609 (I45984,I45752,I45905);
nor I_2610 (I45689,I45888,I45984);
nor I_2611 (I46015,I45922,I45984);
nor I_2612 (I45692,I45837,I46015);
nand I_2613 (I46046,I45752,I45905);
nand I_2614 (I46063,I45820,I46046);
DFFARX1 I_2615 (I46063,I1598,I45718,I45698,);
not I_2616 (I46094,I45888);
nor I_2617 (I45707,I46094,I45939);
nand I_2618 (I45704,I45871,I46094);
nor I_2619 (I46139,I45837,I45888);
nand I_2620 (I45701,I46139,I45752);
not I_2621 (I46194,I1605);
or I_2622 (I46211,I53937,I53934);
nor I_2623 (I46228,I46211,I53943);
nor I_2624 (I46245,I53955,I53940);
or I_2625 (I46262,I46245,I53934);
nor I_2626 (I46279,I53946,I53937);
nand I_2627 (I46296,I46279,I46262);
not I_2628 (I46313,I46296);
nand I_2629 (I46330,I46228,I46313);
nor I_2630 (I46347,I46228,I46313);
nand I_2631 (I46364,I53940,I53952);
nor I_2632 (I46381,I46364,I53949);
nor I_2633 (I46398,I46364,I46381);
not I_2634 (I46415,I46381);
nor I_2635 (I46186,I46415,I46330);
or I_2636 (I46171,I46228,I46415);
nor I_2637 (I46460,I46228,I46381);
nor I_2638 (I46165,I46364,I46460);
nor I_2639 (I46491,I46398,I46460);
nor I_2640 (I46168,I46313,I46491);
nand I_2641 (I46522,I46228,I46381);
nand I_2642 (I46539,I46296,I46522);
DFFARX1 I_2643 (I46539,I1598,I46194,I46174,);
not I_2644 (I46570,I46364);
nor I_2645 (I46183,I46570,I46415);
nand I_2646 (I46180,I46347,I46570);
nor I_2647 (I46615,I46313,I46364);
nand I_2648 (I46177,I46615,I46228);
not I_2649 (I46670,I1605);
or I_2650 (I46687,I19611,I19620);
nor I_2651 (I46704,I46687,I19635);
nor I_2652 (I46721,I19632,I19614);
or I_2653 (I46738,I46721,I19614);
nor I_2654 (I46755,I19611,I19617);
nand I_2655 (I46772,I46755,I46738);
not I_2656 (I46789,I46772);
nand I_2657 (I46806,I46704,I46789);
nor I_2658 (I46823,I46704,I46789);
nand I_2659 (I46840,I19623,I19626);
nor I_2660 (I46857,I46840,I19629);
nor I_2661 (I46874,I46840,I46857);
not I_2662 (I46891,I46857);
nor I_2663 (I46662,I46891,I46806);
or I_2664 (I46647,I46704,I46891);
nor I_2665 (I46936,I46704,I46857);
nor I_2666 (I46641,I46840,I46936);
nor I_2667 (I46967,I46874,I46936);
nor I_2668 (I46644,I46789,I46967);
nand I_2669 (I46998,I46704,I46857);
nand I_2670 (I47015,I46772,I46998);
DFFARX1 I_2671 (I47015,I1598,I46670,I46650,);
not I_2672 (I47046,I46840);
nor I_2673 (I46659,I47046,I46891);
nand I_2674 (I46656,I46823,I47046);
nor I_2675 (I47091,I46789,I46840);
nand I_2676 (I46653,I47091,I46704);
not I_2677 (I47146,I1605);
or I_2678 (I47163,I76921,I76924);
nor I_2679 (I47180,I47163,I76921);
nor I_2680 (I47197,I76918,I76936);
or I_2681 (I47214,I47197,I76924);
nor I_2682 (I47231,I76927,I76918);
nand I_2683 (I47248,I47231,I47214);
not I_2684 (I47265,I47248);
nand I_2685 (I47282,I47180,I47265);
nor I_2686 (I47299,I47180,I47265);
nand I_2687 (I47316,I76933,I76930);
nor I_2688 (I47333,I47316,I76927);
nor I_2689 (I47350,I47316,I47333);
not I_2690 (I47367,I47333);
nor I_2691 (I47138,I47367,I47282);
or I_2692 (I47123,I47180,I47367);
nor I_2693 (I47412,I47180,I47333);
nor I_2694 (I47117,I47316,I47412);
nor I_2695 (I47443,I47350,I47412);
nor I_2696 (I47120,I47265,I47443);
nand I_2697 (I47474,I47180,I47333);
nand I_2698 (I47491,I47248,I47474);
DFFARX1 I_2699 (I47491,I1598,I47146,I47126,);
not I_2700 (I47522,I47316);
nor I_2701 (I47135,I47522,I47367);
nand I_2702 (I47132,I47299,I47522);
nor I_2703 (I47567,I47265,I47316);
nand I_2704 (I47129,I47567,I47180);
not I_2705 (I47622,I1605);
or I_2706 (I47639,I65001,I65022);
nor I_2707 (I47656,I47639,I65007);
nor I_2708 (I47673,I65001,I65019);
or I_2709 (I47690,I47673,I65010);
nor I_2710 (I47707,I65004,I65004);
nand I_2711 (I47724,I47707,I47690);
not I_2712 (I47741,I47724);
nand I_2713 (I47758,I47656,I47741);
nor I_2714 (I47775,I47656,I47741);
nand I_2715 (I47792,I65013,I65016);
nor I_2716 (I47809,I47792,I65007);
nor I_2717 (I47826,I47792,I47809);
not I_2718 (I47843,I47809);
nor I_2719 (I47614,I47843,I47758);
or I_2720 (I47599,I47656,I47843);
nor I_2721 (I47888,I47656,I47809);
nor I_2722 (I47593,I47792,I47888);
nor I_2723 (I47919,I47826,I47888);
nor I_2724 (I47596,I47741,I47919);
nand I_2725 (I47950,I47656,I47809);
nand I_2726 (I47967,I47724,I47950);
DFFARX1 I_2727 (I47967,I1598,I47622,I47602,);
not I_2728 (I47998,I47792);
nor I_2729 (I47611,I47998,I47843);
nand I_2730 (I47608,I47775,I47998);
nor I_2731 (I48043,I47741,I47792);
nand I_2732 (I47605,I48043,I47656);
not I_2733 (I48098,I1605);
or I_2734 (I48115,I54991,I54988);
nor I_2735 (I48132,I48115,I54997);
nor I_2736 (I48149,I55009,I54994);
or I_2737 (I48166,I48149,I54988);
nor I_2738 (I48183,I55000,I54991);
nand I_2739 (I48200,I48183,I48166);
not I_2740 (I48217,I48200);
nand I_2741 (I48234,I48132,I48217);
nor I_2742 (I48251,I48132,I48217);
nand I_2743 (I48268,I54994,I55006);
nor I_2744 (I48285,I48268,I55003);
nor I_2745 (I48302,I48268,I48285);
not I_2746 (I48319,I48285);
nor I_2747 (I48090,I48319,I48234);
or I_2748 (I48075,I48132,I48319);
nor I_2749 (I48364,I48132,I48285);
nor I_2750 (I48069,I48268,I48364);
nor I_2751 (I48395,I48302,I48364);
nor I_2752 (I48072,I48217,I48395);
nand I_2753 (I48426,I48132,I48285);
nand I_2754 (I48443,I48200,I48426);
DFFARX1 I_2755 (I48443,I1598,I48098,I48078,);
not I_2756 (I48474,I48268);
nor I_2757 (I48087,I48474,I48319);
nand I_2758 (I48084,I48251,I48474);
nor I_2759 (I48519,I48217,I48268);
nand I_2760 (I48081,I48519,I48132);
not I_2761 (I48574,I1605);
or I_2762 (I48591,I62893,I62914);
nor I_2763 (I48608,I48591,I62899);
nor I_2764 (I48625,I62893,I62911);
or I_2765 (I48642,I48625,I62902);
nor I_2766 (I48659,I62896,I62896);
nand I_2767 (I48676,I48659,I48642);
not I_2768 (I48693,I48676);
nand I_2769 (I48710,I48608,I48693);
nor I_2770 (I48727,I48608,I48693);
nand I_2771 (I48744,I62905,I62908);
nor I_2772 (I48761,I48744,I62899);
nor I_2773 (I48778,I48744,I48761);
not I_2774 (I48795,I48761);
nor I_2775 (I48566,I48795,I48710);
or I_2776 (I48551,I48608,I48795);
nor I_2777 (I48840,I48608,I48761);
nor I_2778 (I48545,I48744,I48840);
nor I_2779 (I48871,I48778,I48840);
nor I_2780 (I48548,I48693,I48871);
nand I_2781 (I48902,I48608,I48761);
nand I_2782 (I48919,I48676,I48902);
DFFARX1 I_2783 (I48919,I1598,I48574,I48554,);
not I_2784 (I48950,I48744);
nor I_2785 (I48563,I48950,I48795);
nand I_2786 (I48560,I48727,I48950);
nor I_2787 (I48995,I48693,I48744);
nand I_2788 (I48557,I48995,I48608);
not I_2789 (I49050,I1605);
or I_2790 (I49067,I28764,I28749);
nor I_2791 (I49084,I49067,I28743);
nor I_2792 (I49101,I28740,I28761);
or I_2793 (I49118,I49101,I28758);
nor I_2794 (I49135,I28746,I28743);
nand I_2795 (I49152,I49135,I49118);
not I_2796 (I49169,I49152);
nand I_2797 (I49186,I49084,I49169);
nor I_2798 (I49203,I49084,I49169);
nand I_2799 (I49220,I28752,I28755);
nor I_2800 (I49237,I49220,I28740);
nor I_2801 (I49254,I49220,I49237);
not I_2802 (I49271,I49237);
nor I_2803 (I49042,I49271,I49186);
or I_2804 (I49027,I49084,I49271);
nor I_2805 (I49316,I49084,I49237);
nor I_2806 (I49021,I49220,I49316);
nor I_2807 (I49347,I49254,I49316);
nor I_2808 (I49024,I49169,I49347);
nand I_2809 (I49378,I49084,I49237);
nand I_2810 (I49395,I49152,I49378);
DFFARX1 I_2811 (I49395,I1598,I49050,I49030,);
not I_2812 (I49426,I49220);
nor I_2813 (I49039,I49426,I49271);
nand I_2814 (I49036,I49203,I49426);
nor I_2815 (I49471,I49169,I49220);
nand I_2816 (I49033,I49471,I49084);
not I_2817 (I49526,I1605);
or I_2818 (I49543,I22368,I22365);
nor I_2819 (I49560,I49543,I22365);
nor I_2820 (I49577,I22374,I22371);
or I_2821 (I49594,I49577,I22380);
nor I_2822 (I49611,I22383,I22368);
nand I_2823 (I49628,I49611,I49594);
not I_2824 (I49645,I49628);
nand I_2825 (I49662,I49560,I49645);
nor I_2826 (I49679,I49560,I49645);
nand I_2827 (I49696,I22371,I22377);
nor I_2828 (I49713,I49696,I22374);
nor I_2829 (I49730,I49696,I49713);
not I_2830 (I49747,I49713);
nor I_2831 (I49518,I49747,I49662);
or I_2832 (I49503,I49560,I49747);
nor I_2833 (I49792,I49560,I49713);
nor I_2834 (I49497,I49696,I49792);
nor I_2835 (I49823,I49730,I49792);
nor I_2836 (I49500,I49645,I49823);
nand I_2837 (I49854,I49560,I49713);
nand I_2838 (I49871,I49628,I49854);
DFFARX1 I_2839 (I49871,I1598,I49526,I49506,);
not I_2840 (I49902,I49696);
nor I_2841 (I49515,I49902,I49747);
nand I_2842 (I49512,I49679,I49902);
nor I_2843 (I49947,I49645,I49696);
nand I_2844 (I49509,I49947,I49560);
not I_2845 (I50002,I1605);
or I_2846 (I50019,I76479,I76482);
nor I_2847 (I50036,I50019,I76479);
nor I_2848 (I50053,I76476,I76494);
or I_2849 (I50070,I50053,I76482);
nor I_2850 (I50087,I76485,I76476);
nand I_2851 (I50104,I50087,I50070);
not I_2852 (I50121,I50104);
nand I_2853 (I50138,I50036,I50121);
nor I_2854 (I50155,I50036,I50121);
nand I_2855 (I50172,I76491,I76488);
nor I_2856 (I50189,I50172,I76485);
nor I_2857 (I50206,I50172,I50189);
not I_2858 (I50223,I50189);
nor I_2859 (I49994,I50223,I50138);
or I_2860 (I49979,I50036,I50223);
nor I_2861 (I50268,I50036,I50189);
nor I_2862 (I49973,I50172,I50268);
nor I_2863 (I50299,I50206,I50268);
nor I_2864 (I49976,I50121,I50299);
nand I_2865 (I50330,I50036,I50189);
nand I_2866 (I50347,I50104,I50330);
DFFARX1 I_2867 (I50347,I1598,I50002,I49982,);
not I_2868 (I50378,I50172);
nor I_2869 (I49991,I50378,I50223);
nand I_2870 (I49988,I50155,I50378);
nor I_2871 (I50423,I50121,I50172);
nand I_2872 (I49985,I50423,I50036);
not I_2873 (I50478,I1605);
or I_2874 (I50495,I32980,I32965);
nor I_2875 (I50512,I50495,I32959);
nor I_2876 (I50529,I32956,I32977);
or I_2877 (I50546,I50529,I32974);
nor I_2878 (I50563,I32962,I32959);
nand I_2879 (I50580,I50563,I50546);
not I_2880 (I50597,I50580);
nand I_2881 (I50614,I50512,I50597);
nor I_2882 (I50631,I50512,I50597);
nand I_2883 (I50648,I32968,I32971);
nor I_2884 (I50665,I50648,I32956);
nor I_2885 (I50682,I50648,I50665);
not I_2886 (I50699,I50665);
nor I_2887 (I50470,I50699,I50614);
or I_2888 (I50455,I50512,I50699);
nor I_2889 (I50744,I50512,I50665);
nor I_2890 (I50449,I50648,I50744);
nor I_2891 (I50775,I50682,I50744);
nor I_2892 (I50452,I50597,I50775);
nand I_2893 (I50806,I50512,I50665);
nand I_2894 (I50823,I50580,I50806);
DFFARX1 I_2895 (I50823,I1598,I50478,I50458,);
not I_2896 (I50854,I50648);
nor I_2897 (I50467,I50854,I50699);
nand I_2898 (I50464,I50631,I50854);
nor I_2899 (I50899,I50597,I50648);
nand I_2900 (I50461,I50899,I50512);
not I_2901 (I50954,I1605);
or I_2902 (I50971,I22776,I22773);
nor I_2903 (I50988,I50971,I22773);
nor I_2904 (I51005,I22782,I22779);
or I_2905 (I51022,I51005,I22788);
nor I_2906 (I51039,I22791,I22776);
nand I_2907 (I51056,I51039,I51022);
not I_2908 (I51073,I51056);
nand I_2909 (I51090,I50988,I51073);
nor I_2910 (I51107,I50988,I51073);
nand I_2911 (I51124,I22779,I22785);
nor I_2912 (I51141,I51124,I22782);
nor I_2913 (I51158,I51124,I51141);
not I_2914 (I51175,I51141);
nor I_2915 (I50946,I51175,I51090);
or I_2916 (I50931,I50988,I51175);
nor I_2917 (I51220,I50988,I51141);
nor I_2918 (I50925,I51124,I51220);
nor I_2919 (I51251,I51158,I51220);
nor I_2920 (I50928,I51073,I51251);
nand I_2921 (I51282,I50988,I51141);
nand I_2922 (I51299,I51056,I51282);
DFFARX1 I_2923 (I51299,I1598,I50954,I50934,);
not I_2924 (I51330,I51124);
nor I_2925 (I50943,I51330,I51175);
nand I_2926 (I50940,I51107,I51330);
nor I_2927 (I51375,I51073,I51124);
nand I_2928 (I50937,I51375,I50988);
not I_2929 (I51430,I1605);
or I_2930 (I51447,I52883,I52880);
nor I_2931 (I51464,I51447,I52889);
nor I_2932 (I51481,I52901,I52886);
or I_2933 (I51498,I51481,I52880);
nor I_2934 (I51515,I52892,I52883);
nand I_2935 (I51532,I51515,I51498);
not I_2936 (I51549,I51532);
nand I_2937 (I51566,I51464,I51549);
nor I_2938 (I51583,I51464,I51549);
nand I_2939 (I51600,I52886,I52898);
nor I_2940 (I51617,I51600,I52895);
nor I_2941 (I51634,I51600,I51617);
not I_2942 (I51651,I51617);
nor I_2943 (I51422,I51651,I51566);
or I_2944 (I51407,I51464,I51651);
nor I_2945 (I51696,I51464,I51617);
nor I_2946 (I51401,I51600,I51696);
nor I_2947 (I51727,I51634,I51696);
nor I_2948 (I51404,I51549,I51727);
nand I_2949 (I51758,I51464,I51617);
nand I_2950 (I51775,I51532,I51758);
DFFARX1 I_2951 (I51775,I1598,I51430,I51410,);
not I_2952 (I51806,I51600);
nor I_2953 (I51419,I51806,I51651);
nand I_2954 (I51416,I51583,I51806);
nor I_2955 (I51851,I51549,I51600);
nand I_2956 (I51413,I51851,I51464);
not I_2957 (I51906,I1605);
or I_2958 (I51923,I33507,I33492);
nor I_2959 (I51940,I51923,I33486);
nor I_2960 (I51957,I33483,I33504);
or I_2961 (I51974,I51957,I33501);
nor I_2962 (I51991,I33489,I33486);
nand I_2963 (I52008,I51991,I51974);
not I_2964 (I52025,I52008);
nand I_2965 (I52042,I51940,I52025);
nor I_2966 (I52059,I51940,I52025);
nand I_2967 (I52076,I33495,I33498);
nor I_2968 (I52093,I52076,I33483);
nor I_2969 (I52110,I52076,I52093);
not I_2970 (I52127,I52093);
nor I_2971 (I51898,I52127,I52042);
or I_2972 (I51883,I51940,I52127);
nor I_2973 (I52172,I51940,I52093);
nor I_2974 (I51877,I52076,I52172);
nor I_2975 (I52203,I52110,I52172);
nor I_2976 (I51880,I52025,I52203);
nand I_2977 (I52234,I51940,I52093);
nand I_2978 (I52251,I52008,I52234);
DFFARX1 I_2979 (I52251,I1598,I51906,I51886,);
not I_2980 (I52282,I52076);
nor I_2981 (I51895,I52282,I52127);
nand I_2982 (I51892,I52059,I52282);
nor I_2983 (I52327,I52025,I52076);
nand I_2984 (I51889,I52327,I51940);
not I_2985 (I52382,I1605);
or I_2986 (I52399,I25054,I25072);
nand I_2987 (I52416,I25069,I25063);
not I_2988 (I52433,I52416);
nand I_2989 (I52450,I52433,I52399);
not I_2990 (I52467,I52450);
nand I_2991 (I52484,I25060,I25051);
nor I_2992 (I52501,I52484,I25075);
nor I_2993 (I52518,I52450,I52501);
or I_2994 (I52535,I52501,I52467);
nand I_2995 (I52359,I52450,I52501);
nand I_2996 (I52566,I52501,I52467);
and I_2997 (I52583,I52416,I52484);
nor I_2998 (I52600,I52518,I52583);
nor I_2999 (I52617,I25057,I25051);
not I_3000 (I52634,I25066);
nor I_3001 (I52651,I52634,I52617);
nor I_3002 (I52353,I52651,I52416);
nand I_3003 (I52682,I52651,I52535);
nor I_3004 (I52374,I52416,I52682);
nor I_3005 (I52356,I52651,I52600);
not I_3006 (I52368,I52651);
nor I_3007 (I52741,I52651,I25054);
or I_3008 (I52758,I52634,I25054);
nand I_3009 (I52775,I52758,I52566);
DFFARX1 I_3010 (I52775,I1598,I52382,I52362,);
nor I_3011 (I52806,I52634,I25054);
nor I_3012 (I52823,I52651,I52806);
nand I_3013 (I52371,I52823,I52501);
nor I_3014 (I52854,I52634,I52450);
nand I_3015 (I52365,I52854,I52741);
not I_3016 (I52909,I1605);
or I_3017 (I52926,I40950,I40932);
nand I_3018 (I52943,I40944,I40935);
not I_3019 (I52960,I52943);
nand I_3020 (I52977,I52960,I52926);
not I_3021 (I52994,I52977);
nand I_3022 (I53011,I40941,I40932);
nor I_3023 (I53028,I53011,I40929);
nor I_3024 (I53045,I52977,I53028);
or I_3025 (I53062,I53028,I52994);
nand I_3026 (I52886,I52977,I53028);
nand I_3027 (I53093,I53028,I52994);
and I_3028 (I53110,I52943,I53011);
nor I_3029 (I53127,I53045,I53110);
nor I_3030 (I53144,I40947,I40938);
not I_3031 (I53161,I40929);
nor I_3032 (I53178,I53161,I53144);
nor I_3033 (I52880,I53178,I52943);
nand I_3034 (I53209,I53178,I53062);
nor I_3035 (I52901,I52943,I53209);
nor I_3036 (I52883,I53178,I53127);
not I_3037 (I52895,I53178);
nor I_3038 (I53268,I53178,I40935);
or I_3039 (I53285,I53161,I40935);
nand I_3040 (I53302,I53285,I53093);
DFFARX1 I_3041 (I53302,I1598,I52909,I52889,);
nor I_3042 (I53333,I53161,I40935);
nor I_3043 (I53350,I53178,I53333);
nand I_3044 (I52898,I53350,I53028);
nor I_3045 (I53381,I53161,I52977);
nand I_3046 (I52892,I53381,I53268);
not I_3047 (I53436,I1605);
or I_3048 (I53453,I36121,I36139);
nand I_3049 (I53470,I36136,I36130);
not I_3050 (I53487,I53470);
nand I_3051 (I53504,I53487,I53453);
not I_3052 (I53521,I53504);
nand I_3053 (I53538,I36127,I36118);
nor I_3054 (I53555,I53538,I36142);
nor I_3055 (I53572,I53504,I53555);
or I_3056 (I53589,I53555,I53521);
nand I_3057 (I53413,I53504,I53555);
nand I_3058 (I53620,I53555,I53521);
and I_3059 (I53637,I53470,I53538);
nor I_3060 (I53654,I53572,I53637);
nor I_3061 (I53671,I36124,I36118);
not I_3062 (I53688,I36133);
nor I_3063 (I53705,I53688,I53671);
nor I_3064 (I53407,I53705,I53470);
nand I_3065 (I53736,I53705,I53589);
nor I_3066 (I53428,I53470,I53736);
nor I_3067 (I53410,I53705,I53654);
not I_3068 (I53422,I53705);
nor I_3069 (I53795,I53705,I36121);
or I_3070 (I53812,I53688,I36121);
nand I_3071 (I53829,I53812,I53620);
DFFARX1 I_3072 (I53829,I1598,I53436,I53416,);
nor I_3073 (I53860,I53688,I36121);
nor I_3074 (I53877,I53705,I53860);
nand I_3075 (I53425,I53877,I53555);
nor I_3076 (I53908,I53688,I53504);
nand I_3077 (I53419,I53908,I53795);
not I_3078 (I53963,I1605);
or I_3079 (I53980,I60258,I60270);
nand I_3080 (I53997,I60273,I60276);
not I_3081 (I54014,I53997);
nand I_3082 (I54031,I54014,I53980);
not I_3083 (I54048,I54031);
nand I_3084 (I54065,I60258,I60261);
nor I_3085 (I54082,I54065,I60264);
nor I_3086 (I54099,I54031,I54082);
or I_3087 (I54116,I54082,I54048);
nand I_3088 (I53940,I54031,I54082);
nand I_3089 (I54147,I54082,I54048);
and I_3090 (I54164,I53997,I54065);
nor I_3091 (I54181,I54099,I54164);
nor I_3092 (I54198,I60267,I60264);
not I_3093 (I54215,I60279);
nor I_3094 (I54232,I54215,I54198);
nor I_3095 (I53934,I54232,I53997);
nand I_3096 (I54263,I54232,I54116);
nor I_3097 (I53955,I53997,I54263);
nor I_3098 (I53937,I54232,I54181);
not I_3099 (I53949,I54232);
nor I_3100 (I54322,I54232,I60261);
or I_3101 (I54339,I54215,I60261);
nand I_3102 (I54356,I54339,I54147);
DFFARX1 I_3103 (I54356,I1598,I53963,I53943,);
nor I_3104 (I54387,I54215,I60261);
nor I_3105 (I54404,I54232,I54387);
nand I_3106 (I53952,I54404,I54082);
nor I_3107 (I54435,I54215,I54031);
nand I_3108 (I53946,I54435,I54322);
not I_3109 (I54490,I1605);
or I_3110 (I54507,I9921,I9942);
nand I_3111 (I54524,I9936,I9924);
not I_3112 (I54541,I54524);
nand I_3113 (I54558,I54541,I54507);
not I_3114 (I54575,I54558);
nand I_3115 (I54592,I9927,I9933);
nor I_3116 (I54609,I54592,I9939);
nor I_3117 (I54626,I54558,I54609);
or I_3118 (I54643,I54609,I54575);
nand I_3119 (I54467,I54558,I54609);
nand I_3120 (I54674,I54609,I54575);
and I_3121 (I54691,I54524,I54592);
nor I_3122 (I54708,I54626,I54691);
nor I_3123 (I54725,I9924,I9930);
not I_3124 (I54742,I9945);
nor I_3125 (I54759,I54742,I54725);
nor I_3126 (I54461,I54759,I54524);
nand I_3127 (I54790,I54759,I54643);
nor I_3128 (I54482,I54524,I54790);
nor I_3129 (I54464,I54759,I54708);
not I_3130 (I54476,I54759);
nor I_3131 (I54849,I54759,I9921);
or I_3132 (I54866,I54742,I9921);
nand I_3133 (I54883,I54866,I54674);
DFFARX1 I_3134 (I54883,I1598,I54490,I54470,);
nor I_3135 (I54914,I54742,I9921);
nor I_3136 (I54931,I54759,I54914);
nand I_3137 (I54479,I54931,I54609);
nor I_3138 (I54962,I54742,I54558);
nand I_3139 (I54473,I54962,I54849);
not I_3140 (I55017,I1605);
or I_3141 (I55034,I17571,I17592);
nand I_3142 (I55051,I17586,I17574);
not I_3143 (I55068,I55051);
nand I_3144 (I55085,I55068,I55034);
not I_3145 (I55102,I55085);
nand I_3146 (I55119,I17577,I17583);
nor I_3147 (I55136,I55119,I17589);
nor I_3148 (I55153,I55085,I55136);
or I_3149 (I55170,I55136,I55102);
nand I_3150 (I54994,I55085,I55136);
nand I_3151 (I55201,I55136,I55102);
and I_3152 (I55218,I55051,I55119);
nor I_3153 (I55235,I55153,I55218);
nor I_3154 (I55252,I17574,I17580);
not I_3155 (I55269,I17595);
nor I_3156 (I55286,I55269,I55252);
nor I_3157 (I54988,I55286,I55051);
nand I_3158 (I55317,I55286,I55170);
nor I_3159 (I55009,I55051,I55317);
nor I_3160 (I54991,I55286,I55235);
not I_3161 (I55003,I55286);
nor I_3162 (I55376,I55286,I17571);
or I_3163 (I55393,I55269,I17571);
nand I_3164 (I55410,I55393,I55201);
DFFARX1 I_3165 (I55410,I1598,I55017,I54997,);
nor I_3166 (I55441,I55269,I17571);
nor I_3167 (I55458,I55286,I55441);
nand I_3168 (I55006,I55458,I55136);
nor I_3169 (I55489,I55269,I55085);
nand I_3170 (I55000,I55489,I55376);
not I_3171 (I55544,I1605);
or I_3172 (I55561,I2665,I2680);
nand I_3173 (I55578,I2668,I2668);
not I_3174 (I55595,I55578);
nand I_3175 (I55612,I55595,I55561);
not I_3176 (I55629,I55612);
nand I_3177 (I55646,I2671,I2674);
nor I_3178 (I55663,I55646,I2683);
nor I_3179 (I55680,I55612,I55663);
or I_3180 (I55697,I55663,I55629);
nand I_3181 (I55521,I55612,I55663);
nand I_3182 (I55728,I55663,I55629);
and I_3183 (I55745,I55578,I55646);
nor I_3184 (I55762,I55680,I55745);
nor I_3185 (I55779,I2665,I2662);
not I_3186 (I55796,I2677);
nor I_3187 (I55813,I55796,I55779);
nor I_3188 (I55515,I55813,I55578);
nand I_3189 (I55844,I55813,I55697);
nor I_3190 (I55536,I55578,I55844);
nor I_3191 (I55518,I55813,I55762);
not I_3192 (I55530,I55813);
nor I_3193 (I55903,I55813,I2662);
or I_3194 (I55920,I55796,I2662);
nand I_3195 (I55937,I55920,I55728);
DFFARX1 I_3196 (I55937,I1598,I55544,I55524,);
nor I_3197 (I55968,I55796,I2662);
nor I_3198 (I55985,I55813,I55968);
nand I_3199 (I55533,I55985,I55663);
nor I_3200 (I56016,I55796,I55612);
nand I_3201 (I55527,I56016,I55903);
not I_3202 (I56071,I1605);
or I_3203 (I56088,I29797,I29815);
nand I_3204 (I56105,I29812,I29806);
not I_3205 (I56122,I56105);
nand I_3206 (I56139,I56122,I56088);
not I_3207 (I56156,I56139);
nand I_3208 (I56173,I29803,I29794);
nor I_3209 (I56190,I56173,I29818);
nor I_3210 (I56207,I56139,I56190);
or I_3211 (I56224,I56190,I56156);
nand I_3212 (I56048,I56139,I56190);
nand I_3213 (I56255,I56190,I56156);
and I_3214 (I56272,I56105,I56173);
nor I_3215 (I56289,I56207,I56272);
nor I_3216 (I56306,I29800,I29794);
not I_3217 (I56323,I29809);
nor I_3218 (I56340,I56323,I56306);
nor I_3219 (I56042,I56340,I56105);
nand I_3220 (I56371,I56340,I56224);
nor I_3221 (I56063,I56105,I56371);
nor I_3222 (I56045,I56340,I56289);
not I_3223 (I56057,I56340);
nor I_3224 (I56430,I56340,I29797);
or I_3225 (I56447,I56323,I29797);
nand I_3226 (I56464,I56447,I56255);
DFFARX1 I_3227 (I56464,I1598,I56071,I56051,);
nor I_3228 (I56495,I56323,I29797);
nor I_3229 (I56512,I56340,I56495);
nand I_3230 (I56060,I56512,I56190);
nor I_3231 (I56543,I56323,I56139);
nand I_3232 (I56054,I56543,I56430);
not I_3233 (I56598,I1605);
nor I_3234 (I56615,I47135,I47123);
not I_3235 (I56632,I47120);
not I_3236 (I56649,I47117);
nor I_3237 (I56666,I56649,I56615);
nand I_3238 (I56683,I56666,I47120);
not I_3239 (I56572,I56683);
nor I_3240 (I56714,I56649,I56632);
and I_3241 (I56731,I56683,I47120);
nor I_3242 (I56748,I56714,I47120);
nand I_3243 (I56765,I47123,I47129);
not I_3244 (I56782,I56765);
nand I_3245 (I56799,I56782,I56748);
nor I_3246 (I56816,I47138,I47132);
not I_3247 (I56833,I47126);
nor I_3248 (I56850,I56833,I47117);
nor I_3249 (I56569,I56850,I56683);
not I_3250 (I56881,I56850);
or I_3251 (I56584,I56799,I56850);
nor I_3252 (I56912,I56850,I56765);
nand I_3253 (I56581,I56714,I56912);
nor I_3254 (I56943,I56816,I56833);
nand I_3255 (I56960,I56782,I56943);
not I_3256 (I56587,I56960);
nor I_3257 (I56590,I56731,I56960);
or I_3258 (I57005,I56850,I56943);
nor I_3259 (I56575,I56782,I57005);
nor I_3260 (I57036,I56943,I47120);
nand I_3261 (I57053,I57036,I56782);
nand I_3262 (I57070,I56881,I57053);
DFFARX1 I_3263 (I57070,I1598,I56598,I56578,);
not I_3264 (I57125,I1605);
nor I_3265 (I57142,I1143,I1367);
not I_3266 (I57159,I1583);
not I_3267 (I57176,I767);
nor I_3268 (I57193,I57176,I57142);
nand I_3269 (I57210,I57193,I1583);
not I_3270 (I57099,I57210);
nor I_3271 (I57241,I57176,I57159);
and I_3272 (I57258,I57210,I871);
nor I_3273 (I57275,I57241,I871);
nand I_3274 (I57292,I1087,I895);
not I_3275 (I57309,I57292);
nand I_3276 (I57326,I57309,I57275);
nor I_3277 (I57343,I1039,I1023);
not I_3278 (I57360,I839);
nor I_3279 (I57377,I57360,I743);
nor I_3280 (I57096,I57377,I57210);
not I_3281 (I57408,I57377);
or I_3282 (I57111,I57326,I57377);
nor I_3283 (I57439,I57377,I57292);
nand I_3284 (I57108,I57241,I57439);
nor I_3285 (I57470,I57343,I57360);
nand I_3286 (I57487,I57309,I57470);
not I_3287 (I57114,I57487);
nor I_3288 (I57117,I57258,I57487);
or I_3289 (I57532,I57377,I57470);
nor I_3290 (I57102,I57309,I57532);
nor I_3291 (I57563,I57470,I871);
nand I_3292 (I57580,I57563,I57309);
nand I_3293 (I57597,I57408,I57580);
DFFARX1 I_3294 (I57597,I1598,I57125,I57105,);
not I_3295 (I57652,I1605);
nor I_3296 (I57669,I30848,I30872);
not I_3297 (I57686,I30857);
not I_3298 (I57703,I30851);
nor I_3299 (I57720,I57703,I57669);
nand I_3300 (I57737,I57720,I30857);
not I_3301 (I57626,I57737);
nor I_3302 (I57768,I57703,I57686);
and I_3303 (I57785,I57737,I30854);
nor I_3304 (I57802,I57768,I30854);
nand I_3305 (I57819,I30848,I30863);
not I_3306 (I57836,I57819);
nand I_3307 (I57853,I57836,I57802);
nor I_3308 (I57870,I30860,I30851);
not I_3309 (I57887,I30869);
nor I_3310 (I57904,I57887,I30866);
nor I_3311 (I57623,I57904,I57737);
not I_3312 (I57935,I57904);
or I_3313 (I57638,I57853,I57904);
nor I_3314 (I57966,I57904,I57819);
nand I_3315 (I57635,I57768,I57966);
nor I_3316 (I57997,I57870,I57887);
nand I_3317 (I58014,I57836,I57997);
not I_3318 (I57641,I58014);
nor I_3319 (I57644,I57785,I58014);
or I_3320 (I58059,I57904,I57997);
nor I_3321 (I57629,I57836,I58059);
nor I_3322 (I58090,I57997,I30854);
nand I_3323 (I58107,I58090,I57836);
nand I_3324 (I58124,I57935,I58107);
DFFARX1 I_3325 (I58124,I1598,I57652,I57632,);
not I_3326 (I58179,I1605);
nor I_3327 (I58196,I69404,I69407);
not I_3328 (I58213,I69419);
not I_3329 (I58230,I69410);
nor I_3330 (I58247,I58230,I58196);
nand I_3331 (I58264,I58247,I69419);
not I_3332 (I58153,I58264);
nor I_3333 (I58295,I58230,I58213);
and I_3334 (I58312,I58264,I69413);
nor I_3335 (I58329,I58295,I69413);
nand I_3336 (I58346,I69410,I69416);
not I_3337 (I58363,I58346);
nand I_3338 (I58380,I58363,I58329);
nor I_3339 (I58397,I69407,I69422);
not I_3340 (I58414,I69413);
nor I_3341 (I58431,I58414,I69404);
nor I_3342 (I58150,I58431,I58264);
not I_3343 (I58462,I58431);
or I_3344 (I58165,I58380,I58431);
nor I_3345 (I58493,I58431,I58346);
nand I_3346 (I58162,I58295,I58493);
nor I_3347 (I58524,I58397,I58414);
nand I_3348 (I58541,I58363,I58524);
not I_3349 (I58168,I58541);
nor I_3350 (I58171,I58312,I58541);
or I_3351 (I58586,I58431,I58524);
nor I_3352 (I58156,I58363,I58586);
nor I_3353 (I58617,I58524,I69413);
nand I_3354 (I58634,I58617,I58363);
nand I_3355 (I58651,I58462,I58634);
DFFARX1 I_3356 (I58651,I1598,I58179,I58159,);
not I_3357 (I58706,I1605);
nor I_3358 (I58723,I45231,I45219);
not I_3359 (I58740,I45216);
not I_3360 (I58757,I45213);
nor I_3361 (I58774,I58757,I58723);
nand I_3362 (I58791,I58774,I45216);
not I_3363 (I58680,I58791);
nor I_3364 (I58822,I58757,I58740);
and I_3365 (I58839,I58791,I45216);
nor I_3366 (I58856,I58822,I45216);
nand I_3367 (I58873,I45219,I45225);
not I_3368 (I58890,I58873);
nand I_3369 (I58907,I58890,I58856);
nor I_3370 (I58924,I45234,I45228);
not I_3371 (I58941,I45222);
nor I_3372 (I58958,I58941,I45213);
nor I_3373 (I58677,I58958,I58791);
not I_3374 (I58989,I58958);
or I_3375 (I58692,I58907,I58958);
nor I_3376 (I59020,I58958,I58873);
nand I_3377 (I58689,I58822,I59020);
nor I_3378 (I59051,I58924,I58941);
nand I_3379 (I59068,I58890,I59051);
not I_3380 (I58695,I59068);
nor I_3381 (I58698,I58839,I59068);
or I_3382 (I59113,I58958,I59051);
nor I_3383 (I58683,I58890,I59113);
nor I_3384 (I59144,I59051,I45216);
nand I_3385 (I59161,I59144,I58890);
nand I_3386 (I59178,I58989,I59161);
DFFARX1 I_3387 (I59178,I1598,I58706,I58686,);
not I_3388 (I59233,I1605);
nor I_3389 (I59250,I27159,I27183);
not I_3390 (I59267,I27168);
not I_3391 (I59284,I27162);
nor I_3392 (I59301,I59284,I59250);
nand I_3393 (I59318,I59301,I27168);
not I_3394 (I59207,I59318);
nor I_3395 (I59349,I59284,I59267);
and I_3396 (I59366,I59318,I27165);
nor I_3397 (I59383,I59349,I27165);
nand I_3398 (I59400,I27159,I27174);
not I_3399 (I59417,I59400);
nand I_3400 (I59434,I59417,I59383);
nor I_3401 (I59451,I27171,I27162);
not I_3402 (I59468,I27180);
nor I_3403 (I59485,I59468,I27177);
nor I_3404 (I59204,I59485,I59318);
not I_3405 (I59516,I59485);
or I_3406 (I59219,I59434,I59485);
nor I_3407 (I59547,I59485,I59400);
nand I_3408 (I59216,I59349,I59547);
nor I_3409 (I59578,I59451,I59468);
nand I_3410 (I59595,I59417,I59578);
not I_3411 (I59222,I59595);
nor I_3412 (I59225,I59366,I59595);
or I_3413 (I59640,I59485,I59578);
nor I_3414 (I59210,I59417,I59640);
nor I_3415 (I59671,I59578,I27165);
nand I_3416 (I59688,I59671,I59417);
nand I_3417 (I59705,I59516,I59688);
DFFARX1 I_3418 (I59705,I1598,I59233,I59213,);
not I_3419 (I59760,I1605);
nor I_3420 (I59777,I5824,I5827);
not I_3421 (I59794,I5839);
not I_3422 (I59811,I5830);
nor I_3423 (I59828,I59811,I59777);
nand I_3424 (I59845,I59828,I5839);
not I_3425 (I59734,I59845);
nor I_3426 (I59876,I59811,I59794);
and I_3427 (I59893,I59845,I5827);
nor I_3428 (I59910,I59876,I5827);
nand I_3429 (I59927,I5833,I5830);
not I_3430 (I59944,I59927);
nand I_3431 (I59961,I59944,I59910);
nor I_3432 (I59978,I5845,I5842);
not I_3433 (I59995,I5836);
nor I_3434 (I60012,I59995,I5824);
nor I_3435 (I59731,I60012,I59845);
not I_3436 (I60043,I60012);
or I_3437 (I59746,I59961,I60012);
nor I_3438 (I60074,I60012,I59927);
nand I_3439 (I59743,I59876,I60074);
nor I_3440 (I60105,I59978,I59995);
nand I_3441 (I60122,I59944,I60105);
not I_3442 (I59749,I60122);
nor I_3443 (I59752,I59893,I60122);
or I_3444 (I60167,I60012,I60105);
nor I_3445 (I59737,I59944,I60167);
nor I_3446 (I60198,I60105,I5827);
nand I_3447 (I60215,I60198,I59944);
nand I_3448 (I60232,I60043,I60215);
DFFARX1 I_3449 (I60232,I1598,I59760,I59740,);
not I_3450 (I60287,I1605);
nor I_3451 (I60304,I75150,I75153);
not I_3452 (I60321,I75165);
not I_3453 (I60338,I75156);
nor I_3454 (I60355,I60338,I60304);
nand I_3455 (I60372,I60355,I75165);
not I_3456 (I60261,I60372);
nor I_3457 (I60403,I60338,I60321);
and I_3458 (I60420,I60372,I75159);
nor I_3459 (I60437,I60403,I75159);
nand I_3460 (I60454,I75156,I75162);
not I_3461 (I60471,I60454);
nand I_3462 (I60488,I60471,I60437);
nor I_3463 (I60505,I75153,I75168);
not I_3464 (I60522,I75159);
nor I_3465 (I60539,I60522,I75150);
nor I_3466 (I60258,I60539,I60372);
not I_3467 (I60570,I60539);
or I_3468 (I60273,I60488,I60539);
nor I_3469 (I60601,I60539,I60454);
nand I_3470 (I60270,I60403,I60601);
nor I_3471 (I60632,I60505,I60522);
nand I_3472 (I60649,I60471,I60632);
not I_3473 (I60276,I60649);
nor I_3474 (I60279,I60420,I60649);
or I_3475 (I60694,I60539,I60632);
nor I_3476 (I60264,I60471,I60694);
nor I_3477 (I60725,I60632,I75159);
nand I_3478 (I60742,I60725,I60471);
nand I_3479 (I60759,I60570,I60742);
DFFARX1 I_3480 (I60759,I1598,I60287,I60267,);
not I_3481 (I60814,I1605);
nor I_3482 (I60831,I44755,I44743);
not I_3483 (I60848,I44740);
not I_3484 (I60865,I44737);
nor I_3485 (I60882,I60865,I60831);
nand I_3486 (I60899,I60882,I44740);
not I_3487 (I60788,I60899);
nor I_3488 (I60930,I60865,I60848);
and I_3489 (I60947,I60899,I44740);
nor I_3490 (I60964,I60930,I44740);
nand I_3491 (I60981,I44743,I44749);
not I_3492 (I60998,I60981);
nand I_3493 (I61015,I60998,I60964);
nor I_3494 (I61032,I44758,I44752);
not I_3495 (I61049,I44746);
nor I_3496 (I61066,I61049,I44737);
nor I_3497 (I60785,I61066,I60899);
not I_3498 (I61097,I61066);
or I_3499 (I60800,I61015,I61066);
nor I_3500 (I61128,I61066,I60981);
nand I_3501 (I60797,I60930,I61128);
nor I_3502 (I61159,I61032,I61049);
nand I_3503 (I61176,I60998,I61159);
not I_3504 (I60803,I61176);
nor I_3505 (I60806,I60947,I61176);
or I_3506 (I61221,I61066,I61159);
nor I_3507 (I60791,I60998,I61221);
nor I_3508 (I61252,I61159,I44740);
nand I_3509 (I61269,I61252,I60998);
nand I_3510 (I61286,I61097,I61269);
DFFARX1 I_3511 (I61286,I1598,I60814,I60794,);
not I_3512 (I61341,I1605);
nor I_3513 (I61358,I73824,I73827);
not I_3514 (I61375,I73839);
not I_3515 (I61392,I73830);
nor I_3516 (I61409,I61392,I61358);
nand I_3517 (I61426,I61409,I73839);
not I_3518 (I61315,I61426);
nor I_3519 (I61457,I61392,I61375);
and I_3520 (I61474,I61426,I73833);
nor I_3521 (I61491,I61457,I73833);
nand I_3522 (I61508,I73830,I73836);
not I_3523 (I61525,I61508);
nand I_3524 (I61542,I61525,I61491);
nor I_3525 (I61559,I73827,I73842);
not I_3526 (I61576,I73833);
nor I_3527 (I61593,I61576,I73824);
nor I_3528 (I61312,I61593,I61426);
not I_3529 (I61624,I61593);
or I_3530 (I61327,I61542,I61593);
nor I_3531 (I61655,I61593,I61508);
nand I_3532 (I61324,I61457,I61655);
nor I_3533 (I61686,I61559,I61576);
nand I_3534 (I61703,I61525,I61686);
not I_3535 (I61330,I61703);
nor I_3536 (I61333,I61474,I61703);
or I_3537 (I61748,I61593,I61686);
nor I_3538 (I61318,I61525,I61748);
nor I_3539 (I61779,I61686,I73833);
nand I_3540 (I61796,I61779,I61525);
nand I_3541 (I61813,I61624,I61796);
DFFARX1 I_3542 (I61813,I1598,I61341,I61321,);
not I_3543 (I61868,I1605);
nor I_3544 (I61885,I68520,I68523);
not I_3545 (I61902,I68535);
not I_3546 (I61919,I68526);
nor I_3547 (I61936,I61919,I61885);
nand I_3548 (I61953,I61936,I68535);
not I_3549 (I61842,I61953);
nor I_3550 (I61984,I61919,I61902);
and I_3551 (I62001,I61953,I68529);
nor I_3552 (I62018,I61984,I68529);
nand I_3553 (I62035,I68526,I68532);
not I_3554 (I62052,I62035);
nand I_3555 (I62069,I62052,I62018);
nor I_3556 (I62086,I68523,I68538);
not I_3557 (I62103,I68529);
nor I_3558 (I62120,I62103,I68520);
nor I_3559 (I61839,I62120,I61953);
not I_3560 (I62151,I62120);
or I_3561 (I61854,I62069,I62120);
nor I_3562 (I62182,I62120,I62035);
nand I_3563 (I61851,I61984,I62182);
nor I_3564 (I62213,I62086,I62103);
nand I_3565 (I62230,I62052,I62213);
not I_3566 (I61857,I62230);
nor I_3567 (I61860,I62001,I62230);
or I_3568 (I62275,I62120,I62213);
nor I_3569 (I61845,I62052,I62275);
nor I_3570 (I62306,I62213,I68529);
nand I_3571 (I62323,I62306,I62052);
nand I_3572 (I62340,I62151,I62323);
DFFARX1 I_3573 (I62340,I1598,I61868,I61848,);
not I_3574 (I62395,I1605);
nor I_3575 (I62412,I12984,I12981);
not I_3576 (I62429,I12999);
not I_3577 (I62446,I12990);
nor I_3578 (I62463,I62446,I62412);
nand I_3579 (I62480,I62463,I12999);
not I_3580 (I62369,I62480);
nor I_3581 (I62511,I62446,I62429);
and I_3582 (I62528,I62480,I13005);
nor I_3583 (I62545,I62511,I13005);
nand I_3584 (I62562,I13002,I12993);
not I_3585 (I62579,I62562);
nand I_3586 (I62596,I62579,I62545);
nor I_3587 (I62613,I12981,I12984);
not I_3588 (I62630,I12996);
nor I_3589 (I62647,I62630,I12987);
nor I_3590 (I62366,I62647,I62480);
not I_3591 (I62678,I62647);
or I_3592 (I62381,I62596,I62647);
nor I_3593 (I62709,I62647,I62562);
nand I_3594 (I62378,I62511,I62709);
nor I_3595 (I62740,I62613,I62630);
nand I_3596 (I62757,I62579,I62740);
not I_3597 (I62384,I62757);
nor I_3598 (I62387,I62528,I62757);
or I_3599 (I62802,I62647,I62740);
nor I_3600 (I62372,I62579,I62802);
nor I_3601 (I62833,I62740,I13005);
nand I_3602 (I62850,I62833,I62579);
nand I_3603 (I62867,I62678,I62850);
DFFARX1 I_3604 (I62867,I1598,I62395,I62375,);
not I_3605 (I62922,I1605);
nor I_3606 (I62939,I1608,I1611);
not I_3607 (I62956,I1623);
not I_3608 (I62973,I1614);
nor I_3609 (I62990,I62973,I62939);
nand I_3610 (I63007,I62990,I1623);
not I_3611 (I62896,I63007);
nor I_3612 (I63038,I62973,I62956);
and I_3613 (I63055,I63007,I1611);
nor I_3614 (I63072,I63038,I1611);
nand I_3615 (I63089,I1617,I1614);
not I_3616 (I63106,I63089);
nand I_3617 (I63123,I63106,I63072);
nor I_3618 (I63140,I1629,I1626);
not I_3619 (I63157,I1620);
nor I_3620 (I63174,I63157,I1608);
nor I_3621 (I62893,I63174,I63007);
not I_3622 (I63205,I63174);
or I_3623 (I62908,I63123,I63174);
nor I_3624 (I63236,I63174,I63089);
nand I_3625 (I62905,I63038,I63236);
nor I_3626 (I63267,I63140,I63157);
nand I_3627 (I63284,I63106,I63267);
not I_3628 (I62911,I63284);
nor I_3629 (I62914,I63055,I63284);
or I_3630 (I63329,I63174,I63267);
nor I_3631 (I62899,I63106,I63329);
nor I_3632 (I63360,I63267,I1611);
nand I_3633 (I63377,I63360,I63106);
nand I_3634 (I63394,I63205,I63377);
DFFARX1 I_3635 (I63394,I1598,I62922,I62902,);
not I_3636 (I63449,I1605);
nor I_3637 (I63466,I34010,I34034);
not I_3638 (I63483,I34019);
not I_3639 (I63500,I34013);
nor I_3640 (I63517,I63500,I63466);
nand I_3641 (I63534,I63517,I34019);
not I_3642 (I63423,I63534);
nor I_3643 (I63565,I63500,I63483);
and I_3644 (I63582,I63534,I34016);
nor I_3645 (I63599,I63565,I34016);
nand I_3646 (I63616,I34010,I34025);
not I_3647 (I63633,I63616);
nand I_3648 (I63650,I63633,I63599);
nor I_3649 (I63667,I34022,I34013);
not I_3650 (I63684,I34031);
nor I_3651 (I63701,I63684,I34028);
nor I_3652 (I63420,I63701,I63534);
not I_3653 (I63732,I63701);
or I_3654 (I63435,I63650,I63701);
nor I_3655 (I63763,I63701,I63616);
nand I_3656 (I63432,I63565,I63763);
nor I_3657 (I63794,I63667,I63684);
nand I_3658 (I63811,I63633,I63794);
not I_3659 (I63438,I63811);
nor I_3660 (I63441,I63582,I63811);
or I_3661 (I63856,I63701,I63794);
nor I_3662 (I63426,I63633,I63856);
nor I_3663 (I63887,I63794,I34016);
nand I_3664 (I63904,I63887,I63633);
nand I_3665 (I63921,I63732,I63904);
DFFARX1 I_3666 (I63921,I1598,I63449,I63429,);
not I_3667 (I63976,I1605);
nor I_3668 (I63993,I43803,I43791);
not I_3669 (I64010,I43788);
not I_3670 (I64027,I43785);
nor I_3671 (I64044,I64027,I63993);
nand I_3672 (I64061,I64044,I43788);
not I_3673 (I63950,I64061);
nor I_3674 (I64092,I64027,I64010);
and I_3675 (I64109,I64061,I43788);
nor I_3676 (I64126,I64092,I43788);
nand I_3677 (I64143,I43791,I43797);
not I_3678 (I64160,I64143);
nand I_3679 (I64177,I64160,I64126);
nor I_3680 (I64194,I43806,I43800);
not I_3681 (I64211,I43794);
nor I_3682 (I64228,I64211,I43785);
nor I_3683 (I63947,I64228,I64061);
not I_3684 (I64259,I64228);
or I_3685 (I63962,I64177,I64228);
nor I_3686 (I64290,I64228,I64143);
nand I_3687 (I63959,I64092,I64290);
nor I_3688 (I64321,I64194,I64211);
nand I_3689 (I64338,I64160,I64321);
not I_3690 (I63965,I64338);
nor I_3691 (I63968,I64109,I64338);
or I_3692 (I64383,I64228,I64321);
nor I_3693 (I63953,I64160,I64383);
nor I_3694 (I64414,I64321,I43788);
nand I_3695 (I64431,I64414,I64160);
nand I_3696 (I64448,I64259,I64431);
DFFARX1 I_3697 (I64448,I1598,I63976,I63956,);
not I_3698 (I64503,I1605);
nor I_3699 (I64520,I55518,I55515);
not I_3700 (I64537,I55524);
not I_3701 (I64554,I55521);
nor I_3702 (I64571,I64554,I64520);
nand I_3703 (I64588,I64571,I55524);
not I_3704 (I64477,I64588);
nor I_3705 (I64619,I64554,I64537);
and I_3706 (I64636,I64588,I55527);
nor I_3707 (I64653,I64619,I55527);
nand I_3708 (I64670,I55530,I55521);
not I_3709 (I64687,I64670);
nand I_3710 (I64704,I64687,I64653);
nor I_3711 (I64721,I55536,I55533);
not I_3712 (I64738,I55515);
nor I_3713 (I64755,I64738,I55518);
nor I_3714 (I64474,I64755,I64588);
not I_3715 (I64786,I64755);
or I_3716 (I64489,I64704,I64755);
nor I_3717 (I64817,I64755,I64670);
nand I_3718 (I64486,I64619,I64817);
nor I_3719 (I64848,I64721,I64738);
nand I_3720 (I64865,I64687,I64848);
not I_3721 (I64492,I64865);
nor I_3722 (I64495,I64636,I64865);
or I_3723 (I64910,I64755,I64848);
nor I_3724 (I64480,I64687,I64910);
nor I_3725 (I64941,I64848,I55527);
nand I_3726 (I64958,I64941,I64687);
nand I_3727 (I64975,I64786,I64958);
DFFARX1 I_3728 (I64975,I1598,I64503,I64483,);
not I_3729 (I65030,I1605);
nor I_3730 (I65047,I41423,I41411);
not I_3731 (I65064,I41408);
not I_3732 (I65081,I41405);
nor I_3733 (I65098,I65081,I65047);
nand I_3734 (I65115,I65098,I41408);
not I_3735 (I65004,I65115);
nor I_3736 (I65146,I65081,I65064);
and I_3737 (I65163,I65115,I41408);
nor I_3738 (I65180,I65146,I41408);
nand I_3739 (I65197,I41411,I41417);
not I_3740 (I65214,I65197);
nand I_3741 (I65231,I65214,I65180);
nor I_3742 (I65248,I41426,I41420);
not I_3743 (I65265,I41414);
nor I_3744 (I65282,I65265,I41405);
nor I_3745 (I65001,I65282,I65115);
not I_3746 (I65313,I65282);
or I_3747 (I65016,I65231,I65282);
nor I_3748 (I65344,I65282,I65197);
nand I_3749 (I65013,I65146,I65344);
nor I_3750 (I65375,I65248,I65265);
nand I_3751 (I65392,I65214,I65375);
not I_3752 (I65019,I65392);
nor I_3753 (I65022,I65163,I65392);
or I_3754 (I65437,I65282,I65375);
nor I_3755 (I65007,I65214,I65437);
nor I_3756 (I65468,I65375,I41408);
nand I_3757 (I65485,I65468,I65214);
nand I_3758 (I65502,I65313,I65485);
DFFARX1 I_3759 (I65502,I1598,I65030,I65010,);
not I_3760 (I65557,I1605);
nor I_3761 (I65574,I7374,I7371);
not I_3762 (I65591,I7389);
not I_3763 (I65608,I7380);
nor I_3764 (I65625,I65608,I65574);
nand I_3765 (I65642,I65625,I7389);
not I_3766 (I65531,I65642);
nor I_3767 (I65673,I65608,I65591);
and I_3768 (I65690,I65642,I7395);
nor I_3769 (I65707,I65673,I7395);
nand I_3770 (I65724,I7392,I7383);
not I_3771 (I65741,I65724);
nand I_3772 (I65758,I65741,I65707);
nor I_3773 (I65775,I7371,I7374);
not I_3774 (I65792,I7386);
nor I_3775 (I65809,I65792,I7377);
nor I_3776 (I65528,I65809,I65642);
not I_3777 (I65840,I65809);
or I_3778 (I65543,I65758,I65809);
nor I_3779 (I65871,I65809,I65724);
nand I_3780 (I65540,I65673,I65871);
nor I_3781 (I65902,I65775,I65792);
nand I_3782 (I65919,I65741,I65902);
not I_3783 (I65546,I65919);
nor I_3784 (I65549,I65690,I65919);
or I_3785 (I65964,I65809,I65902);
nor I_3786 (I65534,I65741,I65964);
nor I_3787 (I65995,I65902,I7395);
nand I_3788 (I66012,I65995,I65741);
nand I_3789 (I66029,I65840,I66012);
DFFARX1 I_3790 (I66029,I1598,I65557,I65537,);
not I_3791 (I66084,I1605);
nor I_3792 (I66101,I16554,I16551);
not I_3793 (I66118,I16569);
not I_3794 (I66135,I16560);
nor I_3795 (I66152,I66135,I66101);
nand I_3796 (I66169,I66152,I16569);
not I_3797 (I66058,I66169);
nor I_3798 (I66200,I66135,I66118);
and I_3799 (I66217,I66169,I16575);
nor I_3800 (I66234,I66200,I16575);
nand I_3801 (I66251,I16572,I16563);
not I_3802 (I66268,I66251);
nand I_3803 (I66285,I66268,I66234);
nor I_3804 (I66302,I16551,I16554);
not I_3805 (I66319,I16566);
nor I_3806 (I66336,I66319,I16557);
nor I_3807 (I66055,I66336,I66169);
not I_3808 (I66367,I66336);
or I_3809 (I66070,I66285,I66336);
nor I_3810 (I66398,I66336,I66251);
nand I_3811 (I66067,I66200,I66398);
nor I_3812 (I66429,I66302,I66319);
nand I_3813 (I66446,I66268,I66429);
not I_3814 (I66073,I66446);
nor I_3815 (I66076,I66217,I66446);
or I_3816 (I66491,I66336,I66429);
nor I_3817 (I66061,I66268,I66491);
nor I_3818 (I66522,I66429,I16575);
nand I_3819 (I66539,I66522,I66268);
nand I_3820 (I66556,I66367,I66539);
DFFARX1 I_3821 (I66556,I1598,I66084,I66064,);
not I_3822 (I66611,I1605);
nor I_3823 (I66628,I39519,I39507);
not I_3824 (I66645,I39504);
not I_3825 (I66662,I39501);
nor I_3826 (I66679,I66662,I66628);
nand I_3827 (I66696,I66679,I39504);
not I_3828 (I66585,I66696);
nor I_3829 (I66727,I66662,I66645);
and I_3830 (I66744,I66696,I39504);
nor I_3831 (I66761,I66727,I39504);
nand I_3832 (I66778,I39507,I39513);
not I_3833 (I66795,I66778);
nand I_3834 (I66812,I66795,I66761);
nor I_3835 (I66829,I39522,I39516);
not I_3836 (I66846,I39510);
nor I_3837 (I66863,I66846,I39501);
nor I_3838 (I66582,I66863,I66696);
not I_3839 (I66894,I66863);
or I_3840 (I66597,I66812,I66863);
nor I_3841 (I66925,I66863,I66778);
nand I_3842 (I66594,I66727,I66925);
nor I_3843 (I66956,I66829,I66846);
nand I_3844 (I66973,I66795,I66956);
not I_3845 (I66600,I66973);
nor I_3846 (I66603,I66744,I66973);
or I_3847 (I67018,I66863,I66956);
nor I_3848 (I66588,I66795,I67018);
nor I_3849 (I67049,I66956,I39504);
nand I_3850 (I67066,I67049,I66795);
nand I_3851 (I67083,I66894,I67066);
DFFARX1 I_3852 (I67083,I1598,I66611,I66591,);
not I_3853 (I67138,I1605);
nor I_3854 (I67155,I38091,I38079);
not I_3855 (I67172,I38076);
not I_3856 (I67189,I38073);
nor I_3857 (I67206,I67189,I67155);
nand I_3858 (I67223,I67206,I38076);
not I_3859 (I67112,I67223);
nor I_3860 (I67254,I67189,I67172);
and I_3861 (I67271,I67223,I38076);
nor I_3862 (I67288,I67254,I38076);
nand I_3863 (I67305,I38079,I38085);
not I_3864 (I67322,I67305);
nand I_3865 (I67339,I67322,I67288);
nor I_3866 (I67356,I38094,I38088);
not I_3867 (I67373,I38082);
nor I_3868 (I67390,I67373,I38073);
nor I_3869 (I67109,I67390,I67223);
not I_3870 (I67421,I67390);
or I_3871 (I67124,I67339,I67390);
nor I_3872 (I67452,I67390,I67305);
nand I_3873 (I67121,I67254,I67452);
nor I_3874 (I67483,I67356,I67373);
nand I_3875 (I67500,I67322,I67483);
not I_3876 (I67127,I67500);
nor I_3877 (I67130,I67271,I67500);
or I_3878 (I67545,I67390,I67483);
nor I_3879 (I67115,I67322,I67545);
nor I_3880 (I67576,I67483,I38076);
nand I_3881 (I67593,I67576,I67322);
nand I_3882 (I67610,I67421,I67593);
DFFARX1 I_3883 (I67610,I1598,I67138,I67118,);
not I_3884 (I67662,I1605);
and I_3885 (I67679,I30321,I30321);
nor I_3886 (I67696,I67679,I30345);
nand I_3887 (I67713,I30342,I30330);
nor I_3888 (I67730,I67713,I67696);
not I_3889 (I67651,I67730);
not I_3890 (I67761,I67713);
or I_3891 (I67778,I30324,I30324);
nor I_3892 (I67795,I67778,I30327);
nor I_3893 (I67812,I67795,I67761);
nand I_3894 (I67829,I30336,I30339);
nor I_3895 (I67846,I67829,I30333);
not I_3896 (I67863,I67846);
nor I_3897 (I67880,I67730,I67863);
nand I_3898 (I67648,I67880,I67795);
nor I_3899 (I67636,I67863,I67812);
nand I_3900 (I67642,I67795,I67863);
nor I_3901 (I67939,I67730,I67829);
nand I_3902 (I67956,I67939,I67795);
nand I_3903 (I67973,I67863,I67956);
DFFARX1 I_3904 (I67973,I1598,I67662,I67645,);
not I_3905 (I68004,I67829);
or I_3906 (I68021,I67795,I68004);
nor I_3907 (I67639,I67761,I68021);
nor I_3908 (I68052,I67730,I68004);
nand I_3909 (I67654,I68052,I67761);
not I_3910 (I68104,I1605);
and I_3911 (I68121,I37609,I37615);
nor I_3912 (I68138,I68121,I37603);
nand I_3913 (I68155,I37600,I37597);
nor I_3914 (I68172,I68155,I68138);
not I_3915 (I68093,I68172);
not I_3916 (I68203,I68155);
or I_3917 (I68220,I37606,I37618);
nor I_3918 (I68237,I68220,I37600);
nor I_3919 (I68254,I68237,I68203);
nand I_3920 (I68271,I37597,I37612);
nor I_3921 (I68288,I68271,I37603);
not I_3922 (I68305,I68288);
nor I_3923 (I68322,I68172,I68305);
nand I_3924 (I68090,I68322,I68237);
nor I_3925 (I68078,I68305,I68254);
nand I_3926 (I68084,I68237,I68305);
nor I_3927 (I68381,I68172,I68271);
nand I_3928 (I68398,I68381,I68237);
nand I_3929 (I68415,I68305,I68398);
DFFARX1 I_3930 (I68415,I1598,I68104,I68087,);
not I_3931 (I68446,I68271);
or I_3932 (I68463,I68237,I68446);
nor I_3933 (I68081,I68203,I68463);
nor I_3934 (I68494,I68172,I68446);
nand I_3935 (I68096,I68494,I68203);
not I_3936 (I68546,I1605);
and I_3937 (I68563,I39037,I39043);
nor I_3938 (I68580,I68563,I39031);
nand I_3939 (I68597,I39028,I39025);
nor I_3940 (I68614,I68597,I68580);
not I_3941 (I68535,I68614);
not I_3942 (I68645,I68597);
or I_3943 (I68662,I39034,I39046);
nor I_3944 (I68679,I68662,I39028);
nor I_3945 (I68696,I68679,I68645);
nand I_3946 (I68713,I39025,I39040);
nor I_3947 (I68730,I68713,I39031);
not I_3948 (I68747,I68730);
nor I_3949 (I68764,I68614,I68747);
nand I_3950 (I68532,I68764,I68679);
nor I_3951 (I68520,I68747,I68696);
nand I_3952 (I68526,I68679,I68747);
nor I_3953 (I68823,I68614,I68713);
nand I_3954 (I68840,I68823,I68679);
nand I_3955 (I68857,I68747,I68840);
DFFARX1 I_3956 (I68857,I1598,I68546,I68529,);
not I_3957 (I68888,I68713);
or I_3958 (I68905,I68679,I68888);
nor I_3959 (I68523,I68645,I68905);
nor I_3960 (I68936,I68614,I68888);
nand I_3961 (I68538,I68936,I68645);
not I_3962 (I68988,I1605);
and I_3963 (I69005,I27686,I27686);
nor I_3964 (I69022,I69005,I27710);
nand I_3965 (I69039,I27707,I27695);
nor I_3966 (I69056,I69039,I69022);
not I_3967 (I68977,I69056);
not I_3968 (I69087,I69039);
or I_3969 (I69104,I27689,I27689);
nor I_3970 (I69121,I69104,I27692);
nor I_3971 (I69138,I69121,I69087);
nand I_3972 (I69155,I27701,I27704);
nor I_3973 (I69172,I69155,I27698);
not I_3974 (I69189,I69172);
nor I_3975 (I69206,I69056,I69189);
nand I_3976 (I68974,I69206,I69121);
nor I_3977 (I68962,I69189,I69138);
nand I_3978 (I68968,I69121,I69189);
nor I_3979 (I69265,I69056,I69155);
nand I_3980 (I69282,I69265,I69121);
nand I_3981 (I69299,I69189,I69282);
DFFARX1 I_3982 (I69299,I1598,I68988,I68971,);
not I_3983 (I69330,I69155);
or I_3984 (I69347,I69121,I69330);
nor I_3985 (I68965,I69087,I69347);
nor I_3986 (I69378,I69056,I69330);
nand I_3987 (I68980,I69378,I69087);
not I_3988 (I69430,I1605);
and I_3989 (I69447,I64492,I64477);
nor I_3990 (I69464,I69447,I64480);
nand I_3991 (I69481,I64474,I64474);
nor I_3992 (I69498,I69481,I69464);
not I_3993 (I69419,I69498);
not I_3994 (I69529,I69481);
or I_3995 (I69546,I64477,I64495);
nor I_3996 (I69563,I69546,I64486);
nor I_3997 (I69580,I69563,I69529);
nand I_3998 (I69597,I64489,I64483);
nor I_3999 (I69614,I69597,I64480);
not I_4000 (I69631,I69614);
nor I_4001 (I69648,I69498,I69631);
nand I_4002 (I69416,I69648,I69563);
nor I_4003 (I69404,I69631,I69580);
nand I_4004 (I69410,I69563,I69631);
nor I_4005 (I69707,I69498,I69597);
nand I_4006 (I69724,I69707,I69563);
nand I_4007 (I69741,I69631,I69724);
DFFARX1 I_4008 (I69741,I1598,I69430,I69413,);
not I_4009 (I69772,I69597);
or I_4010 (I69789,I69563,I69772);
nor I_4011 (I69407,I69529,I69789);
nor I_4012 (I69820,I69498,I69772);
nand I_4013 (I69422,I69820,I69529);
not I_4014 (I69872,I1605);
and I_4015 (I69889,I8415,I8391);
nor I_4016 (I69906,I69889,I8397);
nand I_4017 (I69923,I8412,I8394);
nor I_4018 (I69940,I69923,I69906);
not I_4019 (I69861,I69940);
not I_4020 (I69971,I69923);
or I_4021 (I69988,I8391,I8394);
nor I_4022 (I70005,I69988,I8406);
nor I_4023 (I70022,I70005,I69971);
nand I_4024 (I70039,I8400,I8403);
nor I_4025 (I70056,I70039,I8409);
not I_4026 (I70073,I70056);
nor I_4027 (I70090,I69940,I70073);
nand I_4028 (I69858,I70090,I70005);
nor I_4029 (I69846,I70073,I70022);
nand I_4030 (I69852,I70005,I70073);
nor I_4031 (I70149,I69940,I70039);
nand I_4032 (I70166,I70149,I70005);
nand I_4033 (I70183,I70073,I70166);
DFFARX1 I_4034 (I70183,I1598,I69872,I69855,);
not I_4035 (I70214,I70039);
or I_4036 (I70231,I70005,I70214);
nor I_4037 (I69849,I69971,I70231);
nor I_4038 (I70262,I69940,I70214);
nand I_4039 (I69864,I70262,I69971);
not I_4040 (I70314,I1605);
and I_4041 (I70331,I53428,I53410);
nor I_4042 (I70348,I70331,I53425);
nand I_4043 (I70365,I53422,I53413);
nor I_4044 (I70382,I70365,I70348);
not I_4045 (I70303,I70382);
not I_4046 (I70413,I70365);
or I_4047 (I70430,I53407,I53413);
nor I_4048 (I70447,I70430,I53407);
nor I_4049 (I70464,I70447,I70413);
nand I_4050 (I70481,I53416,I53419);
nor I_4051 (I70498,I70481,I53410);
not I_4052 (I70515,I70498);
nor I_4053 (I70532,I70382,I70515);
nand I_4054 (I70300,I70532,I70447);
nor I_4055 (I70288,I70515,I70464);
nand I_4056 (I70294,I70447,I70515);
nor I_4057 (I70591,I70382,I70481);
nand I_4058 (I70608,I70591,I70447);
nand I_4059 (I70625,I70515,I70608);
DFFARX1 I_4060 (I70625,I1598,I70314,I70297,);
not I_4061 (I70656,I70481);
or I_4062 (I70673,I70447,I70656);
nor I_4063 (I70291,I70413,I70673);
nor I_4064 (I70704,I70382,I70656);
nand I_4065 (I70306,I70704,I70413);
not I_4066 (I70756,I1605);
and I_4067 (I70773,I65546,I65531);
nor I_4068 (I70790,I70773,I65534);
nand I_4069 (I70807,I65528,I65528);
nor I_4070 (I70824,I70807,I70790);
not I_4071 (I70745,I70824);
not I_4072 (I70855,I70807);
or I_4073 (I70872,I65531,I65549);
nor I_4074 (I70889,I70872,I65540);
nor I_4075 (I70906,I70889,I70855);
nand I_4076 (I70923,I65543,I65537);
nor I_4077 (I70940,I70923,I65534);
not I_4078 (I70957,I70940);
nor I_4079 (I70974,I70824,I70957);
nand I_4080 (I70742,I70974,I70889);
nor I_4081 (I70730,I70957,I70906);
nand I_4082 (I70736,I70889,I70957);
nor I_4083 (I71033,I70824,I70923);
nand I_4084 (I71050,I71033,I70889);
nand I_4085 (I71067,I70957,I71050);
DFFARX1 I_4086 (I71067,I1598,I70756,I70739,);
not I_4087 (I71098,I70923);
or I_4088 (I71115,I70889,I71098);
nor I_4089 (I70733,I70855,I71115);
nor I_4090 (I71146,I70824,I71098);
nand I_4091 (I70748,I71146,I70855);
not I_4092 (I71198,I1605);
and I_4093 (I71215,I18105,I18081);
nor I_4094 (I71232,I71215,I18087);
nand I_4095 (I71249,I18102,I18084);
nor I_4096 (I71266,I71249,I71232);
not I_4097 (I71187,I71266);
not I_4098 (I71297,I71249);
or I_4099 (I71314,I18081,I18084);
nor I_4100 (I71331,I71314,I18096);
nor I_4101 (I71348,I71331,I71297);
nand I_4102 (I71365,I18090,I18093);
nor I_4103 (I71382,I71365,I18099);
not I_4104 (I71399,I71382);
nor I_4105 (I71416,I71266,I71399);
nand I_4106 (I71184,I71416,I71331);
nor I_4107 (I71172,I71399,I71348);
nand I_4108 (I71178,I71331,I71399);
nor I_4109 (I71475,I71266,I71365);
nand I_4110 (I71492,I71475,I71331);
nand I_4111 (I71509,I71399,I71492);
DFFARX1 I_4112 (I71509,I1598,I71198,I71181,);
not I_4113 (I71540,I71365);
or I_4114 (I71557,I71331,I71540);
nor I_4115 (I71175,I71297,I71557);
nor I_4116 (I71588,I71266,I71540);
nand I_4117 (I71190,I71588,I71297);
not I_4118 (I71640,I1605);
and I_4119 (I71657,I34537,I34537);
nor I_4120 (I71674,I71657,I34561);
nand I_4121 (I71691,I34558,I34546);
nor I_4122 (I71708,I71691,I71674);
not I_4123 (I71629,I71708);
not I_4124 (I71739,I71691);
or I_4125 (I71756,I34540,I34540);
nor I_4126 (I71773,I71756,I34543);
nor I_4127 (I71790,I71773,I71739);
nand I_4128 (I71807,I34552,I34555);
nor I_4129 (I71824,I71807,I34549);
not I_4130 (I71841,I71824);
nor I_4131 (I71858,I71708,I71841);
nand I_4132 (I71626,I71858,I71773);
nor I_4133 (I71614,I71841,I71790);
nand I_4134 (I71620,I71773,I71841);
nor I_4135 (I71917,I71708,I71807);
nand I_4136 (I71934,I71917,I71773);
nand I_4137 (I71951,I71841,I71934);
DFFARX1 I_4138 (I71951,I1598,I71640,I71623,);
not I_4139 (I71982,I71807);
or I_4140 (I71999,I71773,I71982);
nor I_4141 (I71617,I71739,I71999);
nor I_4142 (I72030,I71708,I71982);
nand I_4143 (I71632,I72030,I71739);
not I_4144 (I72082,I1605);
and I_4145 (I72099,I49985,I49991);
nor I_4146 (I72116,I72099,I49979);
nand I_4147 (I72133,I49976,I49973);
nor I_4148 (I72150,I72133,I72116);
not I_4149 (I72071,I72150);
not I_4150 (I72181,I72133);
or I_4151 (I72198,I49982,I49994);
nor I_4152 (I72215,I72198,I49976);
nor I_4153 (I72232,I72215,I72181);
nand I_4154 (I72249,I49973,I49988);
nor I_4155 (I72266,I72249,I49979);
not I_4156 (I72283,I72266);
nor I_4157 (I72300,I72150,I72283);
nand I_4158 (I72068,I72300,I72215);
nor I_4159 (I72056,I72283,I72232);
nand I_4160 (I72062,I72215,I72283);
nor I_4161 (I72359,I72150,I72249);
nand I_4162 (I72376,I72359,I72215);
nand I_4163 (I72393,I72283,I72376);
DFFARX1 I_4164 (I72393,I1598,I72082,I72065,);
not I_4165 (I72424,I72249);
or I_4166 (I72441,I72215,I72424);
nor I_4167 (I72059,I72181,I72441);
nor I_4168 (I72472,I72150,I72424);
nand I_4169 (I72074,I72472,I72181);
not I_4170 (I72524,I1605);
and I_4171 (I72541,I20145,I20121);
nor I_4172 (I72558,I72541,I20127);
nand I_4173 (I72575,I20142,I20124);
nor I_4174 (I72592,I72575,I72558);
not I_4175 (I72513,I72592);
not I_4176 (I72623,I72575);
or I_4177 (I72640,I20121,I20124);
nor I_4178 (I72657,I72640,I20136);
nor I_4179 (I72674,I72657,I72623);
nand I_4180 (I72691,I20130,I20133);
nor I_4181 (I72708,I72691,I20139);
not I_4182 (I72725,I72708);
nor I_4183 (I72742,I72592,I72725);
nand I_4184 (I72510,I72742,I72657);
nor I_4185 (I72498,I72725,I72674);
nand I_4186 (I72504,I72657,I72725);
nor I_4187 (I72801,I72592,I72691);
nand I_4188 (I72818,I72801,I72657);
nand I_4189 (I72835,I72725,I72818);
DFFARX1 I_4190 (I72835,I1598,I72524,I72507,);
not I_4191 (I72866,I72691);
or I_4192 (I72883,I72657,I72866);
nor I_4193 (I72501,I72623,I72883);
nor I_4194 (I72914,I72592,I72866);
nand I_4195 (I72516,I72914,I72623);
not I_4196 (I72966,I1605);
and I_4197 (I72983,I6375,I6351);
nor I_4198 (I73000,I72983,I6357);
nand I_4199 (I73017,I6372,I6354);
nor I_4200 (I73034,I73017,I73000);
not I_4201 (I72955,I73034);
not I_4202 (I73065,I73017);
or I_4203 (I73082,I6351,I6354);
nor I_4204 (I73099,I73082,I6366);
nor I_4205 (I73116,I73099,I73065);
nand I_4206 (I73133,I6360,I6363);
nor I_4207 (I73150,I73133,I6369);
not I_4208 (I73167,I73150);
nor I_4209 (I73184,I73034,I73167);
nand I_4210 (I72952,I73184,I73099);
nor I_4211 (I72940,I73167,I73116);
nand I_4212 (I72946,I73099,I73167);
nor I_4213 (I73243,I73034,I73133);
nand I_4214 (I73260,I73243,I73099);
nand I_4215 (I73277,I73167,I73260);
DFFARX1 I_4216 (I73277,I1598,I72966,I72949,);
not I_4217 (I73308,I73133);
or I_4218 (I73325,I73099,I73308);
nor I_4219 (I72943,I73065,I73325);
nor I_4220 (I73356,I73034,I73308);
nand I_4221 (I72958,I73356,I73065);
not I_4222 (I73408,I1605);
and I_4223 (I73425,I28213,I28213);
nor I_4224 (I73442,I73425,I28237);
nand I_4225 (I73459,I28234,I28222);
nor I_4226 (I73476,I73459,I73442);
not I_4227 (I73397,I73476);
not I_4228 (I73507,I73459);
or I_4229 (I73524,I28216,I28216);
nor I_4230 (I73541,I73524,I28219);
nor I_4231 (I73558,I73541,I73507);
nand I_4232 (I73575,I28228,I28231);
nor I_4233 (I73592,I73575,I28225);
not I_4234 (I73609,I73592);
nor I_4235 (I73626,I73476,I73609);
nand I_4236 (I73394,I73626,I73541);
nor I_4237 (I73382,I73609,I73558);
nand I_4238 (I73388,I73541,I73609);
nor I_4239 (I73685,I73476,I73575);
nand I_4240 (I73702,I73685,I73541);
nand I_4241 (I73719,I73609,I73702);
DFFARX1 I_4242 (I73719,I1598,I73408,I73391,);
not I_4243 (I73750,I73575);
or I_4244 (I73767,I73541,I73750);
nor I_4245 (I73385,I73507,I73767);
nor I_4246 (I73798,I73476,I73750);
nand I_4247 (I73400,I73798,I73507);
not I_4248 (I73850,I1605);
and I_4249 (I73867,I24524,I24524);
nor I_4250 (I73884,I73867,I24548);
nand I_4251 (I73901,I24545,I24533);
nor I_4252 (I73918,I73901,I73884);
not I_4253 (I73839,I73918);
not I_4254 (I73949,I73901);
or I_4255 (I73966,I24527,I24527);
nor I_4256 (I73983,I73966,I24530);
nor I_4257 (I74000,I73983,I73949);
nand I_4258 (I74017,I24539,I24542);
nor I_4259 (I74034,I74017,I24536);
not I_4260 (I74051,I74034);
nor I_4261 (I74068,I73918,I74051);
nand I_4262 (I73836,I74068,I73983);
nor I_4263 (I73824,I74051,I74000);
nand I_4264 (I73830,I73983,I74051);
nor I_4265 (I74127,I73918,I74017);
nand I_4266 (I74144,I74127,I73983);
nand I_4267 (I74161,I74051,I74144);
DFFARX1 I_4268 (I74161,I1598,I73850,I73833,);
not I_4269 (I74192,I74017);
or I_4270 (I74209,I73983,I74192);
nor I_4271 (I73827,I73949,I74209);
nor I_4272 (I74240,I73918,I74192);
nand I_4273 (I73842,I74240,I73949);
not I_4274 (I74292,I1605);
and I_4275 (I74309,I15555,I15531);
nor I_4276 (I74326,I74309,I15537);
nand I_4277 (I74343,I15552,I15534);
nor I_4278 (I74360,I74343,I74326);
not I_4279 (I74281,I74360);
not I_4280 (I74391,I74343);
or I_4281 (I74408,I15531,I15534);
nor I_4282 (I74425,I74408,I15546);
nor I_4283 (I74442,I74425,I74391);
nand I_4284 (I74459,I15540,I15543);
nor I_4285 (I74476,I74459,I15549);
not I_4286 (I74493,I74476);
nor I_4287 (I74510,I74360,I74493);
nand I_4288 (I74278,I74510,I74425);
nor I_4289 (I74266,I74493,I74442);
nand I_4290 (I74272,I74425,I74493);
nor I_4291 (I74569,I74360,I74459);
nand I_4292 (I74586,I74569,I74425);
nand I_4293 (I74603,I74493,I74586);
DFFARX1 I_4294 (I74603,I1598,I74292,I74275,);
not I_4295 (I74634,I74459);
or I_4296 (I74651,I74425,I74634);
nor I_4297 (I74269,I74391,I74651);
nor I_4298 (I74682,I74360,I74634);
nand I_4299 (I74284,I74682,I74391);
not I_4300 (I74734,I1605);
and I_4301 (I74751,I26632,I26632);
nor I_4302 (I74768,I74751,I26656);
nand I_4303 (I74785,I26653,I26641);
nor I_4304 (I74802,I74785,I74768);
not I_4305 (I74723,I74802);
not I_4306 (I74833,I74785);
or I_4307 (I74850,I26635,I26635);
nor I_4308 (I74867,I74850,I26638);
nor I_4309 (I74884,I74867,I74833);
nand I_4310 (I74901,I26647,I26650);
nor I_4311 (I74918,I74901,I26644);
not I_4312 (I74935,I74918);
nor I_4313 (I74952,I74802,I74935);
nand I_4314 (I74720,I74952,I74867);
nor I_4315 (I74708,I74935,I74884);
nand I_4316 (I74714,I74867,I74935);
nor I_4317 (I75011,I74802,I74901);
nand I_4318 (I75028,I75011,I74867);
nand I_4319 (I75045,I74935,I75028);
DFFARX1 I_4320 (I75045,I1598,I74734,I74717,);
not I_4321 (I75076,I74901);
or I_4322 (I75093,I74867,I75076);
nor I_4323 (I74711,I74833,I75093);
nor I_4324 (I75124,I74802,I75076);
nand I_4325 (I74726,I75124,I74833);
not I_4326 (I75176,I1605);
and I_4327 (I75193,I10965,I10941);
nor I_4328 (I75210,I75193,I10947);
nand I_4329 (I75227,I10962,I10944);
nor I_4330 (I75244,I75227,I75210);
not I_4331 (I75165,I75244);
not I_4332 (I75275,I75227);
or I_4333 (I75292,I10941,I10944);
nor I_4334 (I75309,I75292,I10956);
nor I_4335 (I75326,I75309,I75275);
nand I_4336 (I75343,I10950,I10953);
nor I_4337 (I75360,I75343,I10959);
not I_4338 (I75377,I75360);
nor I_4339 (I75394,I75244,I75377);
nand I_4340 (I75162,I75394,I75309);
nor I_4341 (I75150,I75377,I75326);
nand I_4342 (I75156,I75309,I75377);
nor I_4343 (I75453,I75244,I75343);
nand I_4344 (I75470,I75453,I75309);
nand I_4345 (I75487,I75377,I75470);
DFFARX1 I_4346 (I75487,I1598,I75176,I75159,);
not I_4347 (I75518,I75343);
or I_4348 (I75535,I75309,I75518);
nor I_4349 (I75153,I75275,I75535);
nor I_4350 (I75566,I75244,I75518);
nand I_4351 (I75168,I75566,I75275);
not I_4352 (I75618,I1605);
and I_4353 (I75635,I19125,I19101);
nor I_4354 (I75652,I75635,I19107);
nand I_4355 (I75669,I19122,I19104);
nor I_4356 (I75686,I75669,I75652);
not I_4357 (I75607,I75686);
not I_4358 (I75717,I75669);
or I_4359 (I75734,I19101,I19104);
nor I_4360 (I75751,I75734,I19116);
nor I_4361 (I75768,I75751,I75717);
nand I_4362 (I75785,I19110,I19113);
nor I_4363 (I75802,I75785,I19119);
not I_4364 (I75819,I75802);
nor I_4365 (I75836,I75686,I75819);
nand I_4366 (I75604,I75836,I75751);
nor I_4367 (I75592,I75819,I75768);
nand I_4368 (I75598,I75751,I75819);
nor I_4369 (I75895,I75686,I75785);
nand I_4370 (I75912,I75895,I75751);
nand I_4371 (I75929,I75819,I75912);
DFFARX1 I_4372 (I75929,I1598,I75618,I75601,);
not I_4373 (I75960,I75785);
or I_4374 (I75977,I75751,I75960);
nor I_4375 (I75595,I75717,I75977);
nor I_4376 (I76008,I75686,I75960);
nand I_4377 (I75610,I76008,I75717);
not I_4378 (I76060,I1605);
and I_4379 (I76077,I48081,I48087);
nor I_4380 (I76094,I76077,I48075);
nand I_4381 (I76111,I48072,I48069);
nor I_4382 (I76128,I76111,I76094);
not I_4383 (I76049,I76128);
not I_4384 (I76159,I76111);
or I_4385 (I76176,I48078,I48090);
nor I_4386 (I76193,I76176,I48072);
nor I_4387 (I76210,I76193,I76159);
nand I_4388 (I76227,I48069,I48084);
nor I_4389 (I76244,I76227,I48075);
not I_4390 (I76261,I76244);
nor I_4391 (I76278,I76128,I76261);
nand I_4392 (I76046,I76278,I76193);
nor I_4393 (I76034,I76261,I76210);
nand I_4394 (I76040,I76193,I76261);
nor I_4395 (I76337,I76128,I76227);
nand I_4396 (I76354,I76337,I76193);
nand I_4397 (I76371,I76261,I76354);
DFFARX1 I_4398 (I76371,I1598,I76060,I76043,);
not I_4399 (I76402,I76227);
or I_4400 (I76419,I76193,I76402);
nor I_4401 (I76037,I76159,I76419);
nor I_4402 (I76450,I76128,I76402);
nand I_4403 (I76052,I76450,I76159);
not I_4404 (I76502,I1605);
and I_4405 (I76519,I63438,I63423);
nor I_4406 (I76536,I76519,I63426);
nand I_4407 (I76553,I63420,I63420);
nor I_4408 (I76570,I76553,I76536);
not I_4409 (I76491,I76570);
not I_4410 (I76601,I76553);
or I_4411 (I76618,I63423,I63441);
nor I_4412 (I76635,I76618,I63432);
nor I_4413 (I76652,I76635,I76601);
nand I_4414 (I76669,I63435,I63429);
nor I_4415 (I76686,I76669,I63426);
not I_4416 (I76703,I76686);
nor I_4417 (I76720,I76570,I76703);
nand I_4418 (I76488,I76720,I76635);
nor I_4419 (I76476,I76703,I76652);
nand I_4420 (I76482,I76635,I76703);
nor I_4421 (I76779,I76570,I76669);
nand I_4422 (I76796,I76779,I76635);
nand I_4423 (I76813,I76703,I76796);
DFFARX1 I_4424 (I76813,I1598,I76502,I76485,);
not I_4425 (I76844,I76669);
or I_4426 (I76861,I76635,I76844);
nor I_4427 (I76479,I76601,I76861);
nor I_4428 (I76892,I76570,I76844);
nand I_4429 (I76494,I76892,I76601);
not I_4430 (I76944,I1605);
and I_4431 (I76961,I5312,I5300);
nor I_4432 (I76978,I76961,I5318);
nand I_4433 (I76995,I5306,I5303);
nor I_4434 (I77012,I76995,I76978);
not I_4435 (I76933,I77012);
not I_4436 (I77043,I76995);
or I_4437 (I77060,I5300,I5297);
nor I_4438 (I77077,I77060,I5297);
nor I_4439 (I77094,I77077,I77043);
nand I_4440 (I77111,I5309,I5303);
nor I_4441 (I77128,I77111,I5315);
not I_4442 (I77145,I77128);
nor I_4443 (I77162,I77012,I77145);
nand I_4444 (I76930,I77162,I77077);
nor I_4445 (I76918,I77145,I77094);
nand I_4446 (I76924,I77077,I77145);
nor I_4447 (I77221,I77012,I77111);
nand I_4448 (I77238,I77221,I77077);
nand I_4449 (I77255,I77145,I77238);
DFFARX1 I_4450 (I77255,I1598,I76944,I76927,);
not I_4451 (I77286,I77111);
or I_4452 (I77303,I77077,I77286);
nor I_4453 (I76921,I77043,I77303);
nor I_4454 (I77334,I77012,I77286);
nand I_4455 (I76936,I77334,I77043);
not I_4456 (I77386,I1605);
and I_4457 (I77403,I43321,I43327);
nor I_4458 (I77420,I77403,I43315);
nand I_4459 (I77437,I43312,I43309);
nor I_4460 (I77454,I77437,I77420);
not I_4461 (I77375,I77454);
not I_4462 (I77485,I77437);
or I_4463 (I77502,I43318,I43330);
nor I_4464 (I77519,I77502,I43312);
nor I_4465 (I77536,I77519,I77485);
nand I_4466 (I77553,I43309,I43324);
nor I_4467 (I77570,I77553,I43315);
not I_4468 (I77587,I77570);
nor I_4469 (I77604,I77454,I77587);
nand I_4470 (I77372,I77604,I77519);
nor I_4471 (I77360,I77587,I77536);
nand I_4472 (I77366,I77519,I77587);
nor I_4473 (I77663,I77454,I77553);
nand I_4474 (I77680,I77663,I77519);
nand I_4475 (I77697,I77587,I77680);
DFFARX1 I_4476 (I77697,I1598,I77386,I77369,);
not I_4477 (I77728,I77553);
or I_4478 (I77745,I77519,I77728);
nor I_4479 (I77363,I77485,I77745);
nor I_4480 (I77776,I77454,I77728);
nand I_4481 (I77378,I77776,I77485);
endmodule


