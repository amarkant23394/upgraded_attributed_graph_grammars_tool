module test_I8561(I8428,I5728,I1477,I4533,I1470,I8561);
input I8428,I5728,I1477,I4533,I1470;
output I8561;
wire I8527,I8233,I8216,I5751,I5713,I6028,I6110,I8445,I8544,I6127,I5722,I8462;
nand I_0(I8527,I8233,I5713);
not I_1(I8233,I5722);
not I_2(I8216,I1477);
not I_3(I5751,I1477);
DFFARX1 I_4(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_5(I1470,I5751,,,I6028,);
DFFARX1 I_6(I1470,I5751,,,I6110,);
or I_7(I8445,I8428,I5728);
nand I_8(I8544,I8527,I8462);
and I_9(I6127,I6110,I4533);
and I_10(I8561,I8527,I8544);
DFFARX1 I_11(I6028,I1470,I5751,,,I5722,);
DFFARX1 I_12(I8445,I1470,I8216,,,I8462,);
endmodule


