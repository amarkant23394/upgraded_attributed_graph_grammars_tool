module test_I7547(I1477,I1470,I6705,I6657,I7547);
input I1477,I1470,I6705,I6657;
output I7547;
wire I6321,I7570,I8059,I7977;
nand I_0(I6321,I6705,I6657);
not I_1(I7547,I8059);
not I_2(I7570,I1477);
DFFARX1 I_3(I7977,I1470,I7570,,,I8059,);
DFFARX1 I_4(I6321,I1470,I7570,,,I7977,);
endmodule


