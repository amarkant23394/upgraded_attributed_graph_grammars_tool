module test_final(G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_13,blif_reset_net_1_r_13,G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13);
input G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_13,blif_reset_net_1_r_13;
output G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13;
wire G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4,n_431_0_l_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n_569_1_r_13,n4_1_l_13,n7_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13;
DFFARX1 I_0(n4_1_r_4,blif_clk_net_1_r_13,n7_13,G42_1_r_4,);
nor I_1(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_2(n_573_1_r_4,G2_0_l_4,n16_4);
nor I_3(n_549_1_r_4,n22_4,n23_4);
nand I_4(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_5(n19_4,blif_clk_net_1_r_13,n7_13,ACVQN2_3_r_4,);
nor I_6(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_7(n19_4,blif_clk_net_1_r_13,n7_13,ACVQN1_5_r_4,);
not I_8(P6_5_r_4,P6_5_r_internal_4);
or I_9(n_431_0_l_4,IN_8_0_l_4,n26_4);
DFFARX1 I_10(n_431_0_l_4,blif_clk_net_1_r_13,n7_13,G78_0_l_4,);
DFFARX1 I_11(IN_2_5_l_4,blif_clk_net_1_r_13,n7_13,ACVQN1_5_l_4,);
not I_12(n16_4,ACVQN1_5_l_4);
DFFARX1 I_13(IN_1_5_l_4,blif_clk_net_1_r_13,n7_13,n17_internal_4,);
not I_14(n17_4,n17_internal_4);
nor I_15(n4_1_r_4,n30_4,n31_4);
nand I_16(n19_4,G1_0_l_4,n33_4);
DFFARX1 I_17(G78_0_l_4,blif_clk_net_1_r_13,n7_13,n15_internal_4,);
not I_18(n15_4,n15_internal_4);
DFFARX1 I_19(ACVQN1_5_l_4,blif_clk_net_1_r_13,n7_13,P6_5_r_internal_4,);
and I_20(n20_4,IN_11_0_l_4,n16_4);
nor I_21(n21_4,G2_0_l_4,IN_10_0_l_4);
nand I_22(n22_4,G78_0_l_4,n25_4);
nand I_23(n23_4,IN_11_0_l_4,n24_4);
not I_24(n24_4,G2_0_l_4);
not I_25(n25_4,IN_10_0_l_4);
and I_26(n26_4,IN_2_0_l_4,n27_4);
nor I_27(n27_4,IN_4_0_l_4,n28_4);
not I_28(n28_4,G1_0_l_4);
not I_29(n29_4,n30_4);
nand I_30(n30_4,IN_7_0_l_4,n32_4);
nand I_31(n31_4,IN_11_0_l_4,n25_4);
nor I_32(n32_4,G2_0_l_4,n33_4);
not I_33(n33_4,IN_5_0_l_4);
DFFARX1 I_34(n4_1_r_13,blif_clk_net_1_r_13,n7_13,G42_1_r_13,);
nor I_35(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_36(n_573_1_r_13,n18_13,n19_13);
nand I_37(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_38(n_569_1_r_13,n17_13,n18_13);
nor I_39(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_40(n_266_and_0_3_l_13,blif_clk_net_1_r_13,n7_13,ACVQN2_3_r_13,);
nor I_41(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_42(n_549_1_l_13,blif_clk_net_1_r_13,n7_13,ACVQN1_5_r_13,);
not I_43(P6_5_r_13,P6_5_r_internal_13);
nor I_44(n4_1_l_13,n_266_and_0_3_r_4,G42_1_r_4);
not I_45(n7_13,blif_reset_net_1_r_13);
DFFARX1 I_46(n4_1_l_13,blif_clk_net_1_r_13,n7_13,n17_internal_13,);
not I_47(n17_13,n17_internal_13);
DFFARX1 I_48(P6_5_r_4,blif_clk_net_1_r_13,n7_13,n28_13,);
DFFARX1 I_49(ACVQN1_5_r_4,blif_clk_net_1_r_13,n7_13,ACVQN1_3_l_13,);
nor I_50(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_51(n_266_and_0_3_l_13,ACVQN1_3_l_13,n_569_1_r_4);
nand I_52(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_53(n_573_1_l_13,blif_clk_net_1_r_13,n7_13,n14_internal_13,);
not I_54(n14_13,n14_internal_13);
and I_55(n_549_1_l_13,n21_13,n26_13);
nand I_56(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_57(n_569_1_l_13,blif_clk_net_1_r_13,n7_13,P6_5_r_internal_13,);
nand I_58(n18_13,n23_13,n24_13);
or I_59(n19_13,G42_1_r_4,n_549_1_r_4);
not I_60(n20_13,n_573_1_r_4);
not I_61(n21_13,n_572_1_r_4);
nand I_62(n22_13,n17_13,n28_13);
not I_63(n23_13,G42_1_r_4);
not I_64(n24_13,n_572_1_r_4);
nor I_65(n25_13,G42_1_r_4,n_549_1_r_4);
nand I_66(n26_13,n27_13,ACVQN2_3_r_4);
not I_67(n27_13,n_549_1_r_4);
endmodule


