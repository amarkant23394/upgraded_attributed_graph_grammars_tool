module test_I6884(I7009,I1477,I1470,I5082,I6924,I6884);
input I7009,I1477,I1470,I5082,I6924;
output I6884;
wire I7173,I7156,I7238,I7427,I5088,I6907,I7410,I7221,I7492;
nor I_0(I7173,I7156,I7009);
DFFARX1 I_1(I7492,I1470,I6907,,,I6884,);
DFFARX1 I_2(I1470,I6907,,,I7156,);
and I_3(I7238,I7221,I7173);
not I_4(I7427,I7410);
DFFARX1 I_5(I1470,,,I5088,);
not I_6(I6907,I1477);
DFFARX1 I_7(I5082,I1470,I6907,,,I7410,);
nand I_8(I7221,I6924,I5088);
or I_9(I7492,I7427,I7238);
endmodule


