module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_7_r_2,n10_2,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N1371_0_r_2,n32_2,n35_2);
nor I_40(N1508_0_r_2,n32_2,n55_2);
not I_41(N1372_1_r_2,n54_2);
nor I_42(N1508_1_r_2,n59_2,n54_2);
nor I_43(N6147_2_r_2,n42_2,n43_2);
nor I_44(N1507_6_r_2,n40_2,n53_2);
nor I_45(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_46(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_47(n_572_7_r_2,n36_2,n37_2);
or I_48(n_573_7_r_2,n34_2,n35_2);
nor I_49(n_549_7_r_2,n40_2,n41_2);
nand I_50(n_569_7_r_2,n38_2,n39_2);
nor I_51(n_452_7_r_2,n59_2,n35_2);
nor I_52(n4_7_l_2,n_429_or_0_5_r_15,N1508_4_r_15);
not I_53(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_54(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_55(n33_2,n59_2);
and I_56(N3_8_l_2,n49_2,n_576_5_r_15);
DFFARX1 I_57(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_58(n32_2,n32_internal_2);
nor I_59(n4_7_r_2,n59_2,n36_2);
not I_60(n34_2,n39_2);
nor I_61(n35_2,N1508_4_r_15,n_429_or_0_5_r_15);
nor I_62(n36_2,N1508_1_r_15,n_429_or_0_5_r_15);
or I_63(n37_2,n_576_5_r_15,N1372_4_r_15);
not I_64(n38_2,n40_2);
nand I_65(n39_2,n45_2,n57_2);
nor I_66(n40_2,n47_2,n_547_5_r_15);
nor I_67(n41_2,n32_2,n36_2);
not I_68(n42_2,n53_2);
nand I_69(n43_2,n44_2,n45_2);
nand I_70(n44_2,n38_2,n46_2);
not I_71(n45_2,n_576_5_r_15);
nand I_72(n46_2,n47_2,n48_2);
nand I_73(n47_2,G78_5_r_15,N1508_6_r_15);
or I_74(n48_2,N1508_1_r_15,G78_5_r_15);
nand I_75(n49_2,N1508_4_r_15,N1507_6_r_15);
nand I_76(n50_2,n51_2,n52_2);
not I_77(n51_2,n47_2);
nand I_78(n52_2,n38_2,n53_2);
nor I_79(n53_2,N1508_1_r_15,N1372_4_r_15);
nand I_80(n54_2,n42_2,n56_2);
nor I_81(n55_2,n34_2,n56_2);
nor I_82(n56_2,N1508_1_r_15,G78_5_r_15);
nand I_83(n57_2,n58_2,N1372_4_r_15);
not I_84(n58_2,G78_5_r_15);
endmodule


