module test_I15798(I13908,I1477,I13987,I13843,I1470,I15798);
input I13908,I1477,I13987,I13843,I1470;
output I15798;
wire I14004,I13749,I15781,I14131,I13737,I13775,I13755,I14196,I14179,I15747,I13826,I13767,I15764,I14162,I13925;
DFFARX1 I_0(I13987,I1470,I13775,,,I14004,);
nand I_1(I13749,I14162,I13908);
and I_2(I15781,I15764,I13755);
and I_3(I14131,I13826);
DFFARX1 I_4(I14131,I1470,I13775,,,I13737,);
not I_5(I13775,I1477);
or I_6(I15798,I15781,I13767);
nand I_7(I13755,I14004,I13925);
and I_8(I14196,I14004,I14179);
nand I_9(I14179,I14162,I13826);
not I_10(I15747,I13749);
DFFARX1 I_11(I1470,I13775,,,I13826,);
DFFARX1 I_12(I14196,I1470,I13775,,,I13767,);
nor I_13(I15764,I15747,I13737);
DFFARX1 I_14(I1470,I13775,,,I14162,);
nor I_15(I13925,I13843,I13908);
endmodule


