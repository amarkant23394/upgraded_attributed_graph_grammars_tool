module test_I12636(I1477,I10664,I11167,I9459,I1470,I10732,I9864,I12636);
input I1477,I10664,I11167,I9459,I1470,I10732,I9864;
output I12636;
wire I10612,I10647,I9491,I10961,I11184,I10639,I9468,I11201,I11009;
DFFARX1 I_0(I11009,I1470,I10647,,,I10612,);
not I_1(I10647,I1477);
not I_2(I9491,I1477);
nand I_3(I10961,I10664,I9459);
nand I_4(I11184,I11167,I10732);
DFFARX1 I_5(I11201,I1470,I10647,,,I10639,);
DFFARX1 I_6(I9864,I1470,I9491,,,I9468,);
and I_7(I11201,I10961,I11184);
nand I_8(I12636,I10612,I10639);
DFFARX1 I_9(I9468,I1470,I10647,,,I11009,);
endmodule


